
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  G42,
  G43,
  G44,
  G45,
  G46,
  G47,
  G48,
  G49,
  G50,
  n1836_lo,
  n1872_lo,
  n1884_lo,
  n1911_lo,
  n1914_lo,
  n1917_lo,
  n1923_lo,
  n1926_lo,
  n1929_lo,
  n1935_lo,
  n1938_lo,
  n1947_lo,
  n1950_lo,
  n1959_lo,
  n1962_lo,
  n1971_lo,
  n1974_lo,
  n1983_lo,
  n1995_lo,
  n2007_lo,
  n2019_lo,
  n2031_lo,
  n2043_lo,
  n2055_lo,
  n2064_lo,
  n2067_lo,
  n2100_lo,
  n2112_lo,
  n2124_lo,
  n2136_lo,
  n2148_lo,
  n2160_lo,
  n2163_lo,
  n2172_lo,
  n2175_lo,
  n2184_lo,
  n2223_lo,
  n2235_lo,
  n2238_lo,
  n2247_lo,
  n2250_lo,
  n2259_lo,
  n2262_lo,
  n2271_lo,
  n2274_lo,
  n2283_lo,
  n2286_lo,
  n2295_lo,
  n2298_lo,
  n2304_lo,
  n2307_lo,
  n2331_lo,
  n2334_lo,
  n2337_lo,
  n2340_lo,
  n3241_o2,
  n3242_o2,
  n3610_o2,
  n3980_o2,
  n3968_o2,
  n4298_o2,
  n4371_o2,
  n4413_o2,
  n4418_o2,
  n4628_o2,
  n4629_o2,
  n4633_o2,
  n4634_o2,
  n4732_o2,
  n4733_o2,
  n4884_o2,
  n4886_o2,
  n4890_o2,
  n5011_o2,
  n5012_o2,
  n5013_o2,
  n5014_o2,
  n5015_o2,
  n5021_o2,
  n5016_o2,
  n5026_o2,
  n4377_o2,
  n4378_o2,
  n4389_o2,
  n327_inv,
  n330_inv,
  n4398_o2,
  n4401_o2,
  n5117_o2,
  n5115_o2,
  n5122_o2,
  n5121_o2,
  n5119_o2,
  n5116_o2,
  n5123_o2,
  n5156_o2,
  n5167_o2,
  n4454_o2,
  n4455_o2,
  n4456_o2,
  n4505_o2,
  G742_o2,
  G727_o2,
  n4567_o2,
  n4568_o2,
  n4569_o2,
  n4571_o2,
  n4572_o2,
  n399_inv,
  n4539_o2,
  n4651_o2,
  n4652_o2,
  n4653_o2,
  G1514_o2,
  G1823_o2,
  n4783_o2,
  n4787_o2,
  n426_inv,
  n429_inv,
  n4816_o2,
  n435_inv,
  G572_o2,
  n4919_o2,
  n4920_o2,
  n4921_o2,
  G1048_o2,
  n5041_o2,
  n5094_o2,
  n5278_o2,
  n5301_o2,
  G2610_o2,
  G3174_o2,
  G3146_o2,
  G3217_o2,
  G3220_o2,
  G2839_o2,
  G3251_o2,
  G3042_o2,
  G3045_o2,
  G3262_o2,
  G2845_o2,
  G2929_o2,
  G2848_o2,
  G2851_o2,
  G3291_o2,
  G3254_o2,
  G2666_o2,
  n5099_o2,
  n5100_o2,
  n5101_o2,
  G2558_o2,
  n5266_o2,
  n5267_o2,
  G2759_o2,
  n537_inv,
  n540_inv,
  n543_inv,
  n5292_o2,
  n5293_o2,
  n5294_o2,
  n5295_o2,
  G618_o2,
  G621_o2,
  G384_o2,
  G377_o2,
  n570_inv,
  G3171_o2,
  G2552_o2,
  G3272_o2,
  G2015_o2,
  G3294_o2,
  G3281_o2,
  G3320_o2,
  G3275_o2,
  G3140_o2,
  G2836_o2,
  G2926_o2,
  G2842_o2,
  G3302_o2,
  G3288_o2,
  G3143_o2,
  G3100_o2,
  G2512_o2,
  n5325_o2,
  n5326_o2,
  n5327_o2,
  n1857_lo_buf_o2,
  n2097_lo_buf_o2,
  G2669_o2,
  n642_inv,
  G568_o2,
  n648_inv,
  G565_o2,
  G559_o2,
  n1821_lo_buf_o2,
  n1905_lo_buf_o2,
  n2133_lo_buf_o2,
  n2145_lo_buf_o2,
  n2157_lo_buf_o2,
  n2205_lo_buf_o2,
  n2217_lo_buf_o2,
  G447_o2,
  G434_o2,
  G422_o2,
  G461_o2,
  G3312_o2,
  G3332_o2,
  G3195_o2,
  G2607_o2,
  n702_inv,
  G1005_o2,
  G1008_o2,
  n2001_lo_buf_o2,
  n2169_lo_buf_o2,
  n2229_lo_buf_o2,
  n2301_lo_buf_o2,
  n723_inv,
  G2947_o2,
  n2013_lo_buf_o2,
  n2025_lo_buf_o2,
  n2037_lo_buf_o2,
  n2049_lo_buf_o2,
  n2181_lo_buf_o2,
  n744_inv,
  n747_inv,
  n750_inv,
  n753_inv,
  G3350_o2,
  G3360_o2,
  G3373_o2,
  G3237_o2,
  G2773_o2,
  G1733_o2,
  G1738_o2,
  G1751_o2,
  G2216_o2,
  G2219_o2,
  n786_inv,
  n789_inv,
  G787_o2,
  G2823_o2,
  G2796_o2,
  G875_o2,
  G2208_o2,
  G2211_o2,
  n1989_lo_buf_o2,
  n2061_lo_buf_o2,
  n2313_lo_buf_o2,
  G2232_o2,
  G1725_o2,
  G1764_o2,
  G2356_o2,
  G2359_o2,
  G1180_o2,
  G1756_o2,
  G2441_o2,
  G2887_o2,
  G2991_o2,
  n849_inv,
  n852_inv,
  n855_inv,
  n858_inv,
  n861_inv,
  G2805_o2,
  G2906_o2,
  G2833_o2,
  n873_inv,
  G3353_o2,
  G3367_o2,
  G3346_o2,
  G3340_o2,
  G3376_o2,
  G3359_o2,
  G3240_o2,
  G3344_o2,
  G2880_o2,
  G2939_o2,
  G2248_o2,
  G2251_o2,
  G2021_o2,
  G3383_o2,
  G3399_o2,
  G3404_o2,
  G3265_o2,
  G2866_o2,
  G2999_o2,
  G736_o2,
  G739_o2,
  G1200_o2,
  G1203_o2,
  G3027_o2,
  G1463_o2,
  G1460_o2,
  G3012_o2,
  G1574_o2,
  G1646_o2,
  G1592_o2,
  G1664_o2,
  G1547_o2,
  G1619_o2,
  G1556_o2,
  G1628_o2,
  G1583_o2,
  G1655_o2,
  G1529_o2,
  G1601_o2,
  G1538_o2,
  G1610_o2,
  G1565_o2,
  G1637_o2,
  G2437_o2,
  n1008_inv,
  n1785_lo_buf_o2,
  n1845_lo_buf_o2,
  n1893_lo_buf_o2,
  n1941_lo_buf_o2,
  n1953_lo_buf_o2,
  n1965_lo_buf_o2,
  n1977_lo_buf_o2,
  n2241_lo_buf_o2,
  n2253_lo_buf_o2,
  n2265_lo_buf_o2,
  n2277_lo_buf_o2,
  n2289_lo_buf_o2,
  G519_o2,
  n1050_inv,
  n1053_inv,
  n1056_inv,
  G1318_o2,
  n1062_inv,
  G593_o2,
  n1068_inv,
  n1071_inv,
  n1074_inv,
  G2284_o2,
  G2580_o2,
  G2302_o2,
  G2598_o2,
  G2497_o2,
  G2651_o2,
  G2296_o2,
  G2308_o2,
  G2592_o2,
  G2604_o2,
  G2902_o2,
  G2975_o2,
  G2962_o2,
  G3069_o2,
  G2018_o2,
  G1176_o2,
  G1189_o2,
  G3066_o2,
  G3137_o2,
  G3038_o2,
  G3117_o2,
  G2384_o2,
  G2472_o2,
  G772_o2,
  G935_o2,
  G2923_o2,
  G2971_o2,
  G2980_o2,
  G3039_o2,
  G2388_o2,
  G2287_o2,
  G3024_o2,
  G2916_o2,
  n1176_inv,
  G3035_o2,
  G3107_o2,
  G1023_o2,
  G1024_o2,
  G1311_o2,
  G1312_o2,
  G3063_o2,
  G1520_o2,
  G1519_o2,
  G3078_o2,
  G2038_o2,
  G1848_o2,
  G1864_o2,
  G1872_o2,
  G1880_o2,
  G1888_o2,
  G1912_o2,
  G1928_o2,
  G1936_o2,
  G1944_o2,
  G1952_o2,
  G1850_o2,
  G1866_o2,
  G1874_o2,
  G1882_o2,
  G1890_o2,
  G1914_o2,
  G1930_o2,
  G1938_o2,
  G1946_o2,
  G1954_o2,
  G1845_o2,
  G1861_o2,
  G1869_o2,
  G1877_o2,
  G1885_o2,
  G1909_o2,
  G1925_o2,
  G1933_o2,
  G1941_o2,
  G1949_o2,
  G1846_o2,
  G1862_o2,
  G1870_o2,
  G1878_o2,
  G1886_o2,
  G1910_o2,
  G1926_o2,
  G1934_o2,
  G1942_o2,
  G1950_o2,
  G1849_o2,
  G1865_o2,
  G1873_o2,
  G1881_o2,
  G1889_o2,
  G1913_o2,
  G1929_o2,
  G1937_o2,
  G1945_o2,
  G1953_o2,
  G1843_o2,
  G1859_o2,
  G1867_o2,
  G1875_o2,
  G1883_o2,
  G1907_o2,
  G1923_o2,
  G1931_o2,
  G1939_o2,
  G1947_o2,
  G1844_o2,
  G1860_o2,
  G1868_o2,
  G1876_o2,
  G1884_o2,
  G1908_o2,
  G1924_o2,
  G1932_o2,
  G1940_o2,
  G1948_o2,
  G1847_o2,
  G1863_o2,
  G1871_o2,
  G1879_o2,
  G1887_o2,
  G1911_o2,
  G1927_o2,
  G1935_o2,
  G1943_o2,
  G1951_o2,
  G2444_o2,
  G2451_o2,
  G2502_o2,
  G2507_o2,
  n1464_inv,
  G2583_o2,
  n1797_lo_buf_o2,
  n1833_lo_buf_o2,
  n1881_lo_buf_o2,
  n1479_inv,
  n1482_inv,
  n1485_inv,
  G615_o2,
  G2254_o2,
  G2255_o2,
  G2027_o2,
  G2393_o2,
  G527_o2,
  G594_o2,
  G1689_o2,
  G1693_o2,
  G2281_o2,
  G2014_o2,
  G2459_o2,
  G2561_o2,
  G2533_o2,
  n1749_lo_buf_o2,
  n1761_lo_buf_o2,
  n1773_lo_buf_o2,
  n1809_lo_buf_o2,
  G1955_o2,
  G1958_o2,
  G2562_o2,
  G2398_o2,
  n1554_inv,
  n1557_inv,
  G2577_o2,
  G2627_o2,
  G654_o2,
  G660_o2,
  G831_o2,
  G919_o2,
  G925_o2,
  n1815_lo_buf_o2,
  n1899_lo_buf_o2,
  n2079_lo_buf_o2,
  n2127_lo_buf_o2,
  n2139_lo_buf_o2,
  n2151_lo_buf_o2,
  n2187_lo_buf_o2,
  n2199_lo_buf_o2,
  n2211_lo_buf_o2,
  G533_o2,
  n1854_lo_buf_o2,
  n2094_lo_buf_o2,
  G667_o2,
  G874_o2,
  G851_o2,
  G1127_o2,
  n1869_lo_buf_o2,
  n2109_lo_buf_o2,
  n2121_lo_buf_o2,
  G477_o2,
  G491_o2,
  G501_o2,
  G786_o2,
  G791_o2,
  G1126_o2,
  G1052_o2,
  G1054_o2,
  G3519,
  G3520,
  G3521,
  G3522,
  G3523,
  G3524,
  G3525,
  G3526,
  G3527,
  G3528,
  G3529,
  G3530,
  G3531,
  G3532,
  G3533,
  G3534,
  G3535,
  G3536,
  G3537,
  G3538,
  G3539,
  G3540,
  n1836_li,
  n1872_li,
  n1884_li,
  n1911_li,
  n1914_li,
  n1917_li,
  n1923_li,
  n1926_li,
  n1929_li,
  n1935_li,
  n1938_li,
  n1947_li,
  n1950_li,
  n1959_li,
  n1962_li,
  n1971_li,
  n1974_li,
  n1983_li,
  n1995_li,
  n2007_li,
  n2019_li,
  n2031_li,
  n2043_li,
  n2055_li,
  n2064_li,
  n2067_li,
  n2100_li,
  n2112_li,
  n2124_li,
  n2136_li,
  n2148_li,
  n2160_li,
  n2163_li,
  n2172_li,
  n2175_li,
  n2184_li,
  n2223_li,
  n2235_li,
  n2238_li,
  n2247_li,
  n2250_li,
  n2259_li,
  n2262_li,
  n2271_li,
  n2274_li,
  n2283_li,
  n2286_li,
  n2295_li,
  n2298_li,
  n2304_li,
  n2307_li,
  n2331_li,
  n2334_li,
  n2337_li,
  n2340_li,
  n3241_i2,
  n3242_i2,
  n3610_i2,
  n3980_i2,
  n3968_i2,
  n4298_i2,
  n4371_i2,
  n4413_i2,
  n4418_i2,
  n4628_i2,
  n4629_i2,
  n4633_i2,
  n4634_i2,
  n4732_i2,
  n4733_i2,
  n4884_i2,
  n4886_i2,
  n4890_i2,
  n5011_i2,
  n5012_i2,
  n5013_i2,
  n5014_i2,
  n5015_i2,
  n5021_i2,
  n5016_i2,
  n5026_i2,
  n4377_i2,
  n4378_i2,
  n4389_i2,
  n4390_i2,
  n4391_i2,
  n4398_i2,
  n4401_i2,
  n5117_i2,
  n5115_i2,
  n5122_i2,
  n5121_i2,
  n5119_i2,
  n5116_i2,
  n5123_i2,
  n5156_i2,
  n5167_i2,
  n4454_i2,
  n4455_i2,
  n4456_i2,
  n4505_i2,
  G742_i2,
  G727_i2,
  n4567_i2,
  n4568_i2,
  n4569_i2,
  n4571_i2,
  n4572_i2,
  n4537_i2,
  n4539_i2,
  n4651_i2,
  n4652_i2,
  n4653_i2,
  G1514_i2,
  G1823_i2,
  n4783_i2,
  n4787_i2,
  n4808_i2,
  n4815_i2,
  n4816_i2,
  n4822_i2,
  G572_i2,
  n4919_i2,
  n4920_i2,
  n4921_i2,
  G1048_i2,
  n5041_i2,
  n5094_i2,
  n5278_i2,
  n5301_i2,
  G2610_i2,
  G3174_i2,
  G3146_i2,
  G3217_i2,
  G3220_i2,
  G2839_i2,
  G3251_i2,
  G3042_i2,
  G3045_i2,
  G3262_i2,
  G2845_i2,
  G2929_i2,
  G2848_i2,
  G2851_i2,
  G3291_i2,
  G3254_i2,
  G2666_i2,
  n5099_i2,
  n5100_i2,
  n5101_i2,
  G2558_i2,
  n5266_i2,
  n5267_i2,
  G2759_i2,
  n5269_i2,
  n5270_i2,
  n5271_i2,
  n5292_i2,
  n5293_i2,
  n5294_i2,
  n5295_i2,
  G618_i2,
  G621_i2,
  G384_i2,
  G377_i2,
  G400_i2,
  G3171_i2,
  G2552_i2,
  G3272_i2,
  G2015_i2,
  G3294_i2,
  G3281_i2,
  G3320_i2,
  G3275_i2,
  G3140_i2,
  G2836_i2,
  G2926_i2,
  G2842_i2,
  G3302_i2,
  G3288_i2,
  G3143_i2,
  G3100_i2,
  G2512_i2,
  n5325_i2,
  n5326_i2,
  n5327_i2,
  n1857_lo_buf_i2,
  n2097_lo_buf_i2,
  G2669_i2,
  G552_i2,
  G568_i2,
  G530_i2,
  G565_i2,
  G559_i2,
  n1821_lo_buf_i2,
  n1905_lo_buf_i2,
  n2133_lo_buf_i2,
  n2145_lo_buf_i2,
  n2157_lo_buf_i2,
  n2205_lo_buf_i2,
  n2217_lo_buf_i2,
  G447_i2,
  G434_i2,
  G422_i2,
  G461_i2,
  G3312_i2,
  G3332_i2,
  G3195_i2,
  G2607_i2,
  G2799_i2,
  G1005_i2,
  G1008_i2,
  n2001_lo_buf_i2,
  n2169_lo_buf_i2,
  n2229_lo_buf_i2,
  n2301_lo_buf_i2,
  G2816_i2,
  G2947_i2,
  n2013_lo_buf_i2,
  n2025_lo_buf_i2,
  n2037_lo_buf_i2,
  n2049_lo_buf_i2,
  n2181_lo_buf_i2,
  G546_i2,
  G480_i2,
  G492_i2,
  G540_i2,
  G3350_i2,
  G3360_i2,
  G3373_i2,
  G3237_i2,
  G2773_i2,
  G1733_i2,
  G1738_i2,
  G1751_i2,
  G2216_i2,
  G2219_i2,
  G381_i2,
  G397_i2,
  G787_i2,
  G2823_i2,
  G2796_i2,
  G875_i2,
  G2208_i2,
  G2211_i2,
  n1989_lo_buf_i2,
  n2061_lo_buf_i2,
  n2313_lo_buf_i2,
  G2232_i2,
  G1725_i2,
  G1764_i2,
  G2356_i2,
  G2359_i2,
  G1180_i2,
  G1756_i2,
  G2441_i2,
  G2887_i2,
  G2991_i2,
  G470_i2,
  G484_i2,
  G496_i2,
  G353_i2,
  G363_i2,
  G2805_i2,
  G2906_i2,
  G2833_i2,
  G1012_i2,
  G3353_i2,
  G3367_i2,
  G3346_i2,
  G3340_i2,
  G3376_i2,
  G3359_i2,
  G3240_i2,
  G3344_i2,
  G2880_i2,
  G2939_i2,
  G2248_i2,
  G2251_i2,
  G2021_i2,
  G3383_i2,
  G3399_i2,
  G3404_i2,
  G3265_i2,
  G2866_i2,
  G2999_i2,
  G736_i2,
  G739_i2,
  G1200_i2,
  G1203_i2,
  G3027_i2,
  G1463_i2,
  G1460_i2,
  G3012_i2,
  G1574_i2,
  G1646_i2,
  G1592_i2,
  G1664_i2,
  G1547_i2,
  G1619_i2,
  G1556_i2,
  G1628_i2,
  G1583_i2,
  G1655_i2,
  G1529_i2,
  G1601_i2,
  G1538_i2,
  G1610_i2,
  G1565_i2,
  G1637_i2,
  G2437_i2,
  G2518_i2,
  n1785_lo_buf_i2,
  n1845_lo_buf_i2,
  n1893_lo_buf_i2,
  n1941_lo_buf_i2,
  n1953_lo_buf_i2,
  n1965_lo_buf_i2,
  n1977_lo_buf_i2,
  n2241_lo_buf_i2,
  n2253_lo_buf_i2,
  n2265_lo_buf_i2,
  n2277_lo_buf_i2,
  n2289_lo_buf_i2,
  G519_i2,
  G388_i2,
  G438_i2,
  G368_i2,
  G1318_i2,
  G425_i2,
  G593_i2,
  G413_i2,
  G404_i2,
  G451_i2,
  G2284_i2,
  G2580_i2,
  G2302_i2,
  G2598_i2,
  G2497_i2,
  G2651_i2,
  G2296_i2,
  G2308_i2,
  G2592_i2,
  G2604_i2,
  G2902_i2,
  G2975_i2,
  G2962_i2,
  G3069_i2,
  G2018_i2,
  G1176_i2,
  G1189_i2,
  G3066_i2,
  G3137_i2,
  G3038_i2,
  G3117_i2,
  G2384_i2,
  G2472_i2,
  G772_i2,
  G935_i2,
  G2923_i2,
  G2971_i2,
  G2980_i2,
  G3039_i2,
  G2388_i2,
  G2287_i2,
  G3024_i2,
  G2916_i2,
  G1819_i2,
  G3035_i2,
  G3107_i2,
  G1023_i2,
  G1024_i2,
  G1311_i2,
  G1312_i2,
  G3063_i2,
  G1520_i2,
  G1519_i2,
  G3078_i2,
  G2038_i2,
  G1848_i2,
  G1864_i2,
  G1872_i2,
  G1880_i2,
  G1888_i2,
  G1912_i2,
  G1928_i2,
  G1936_i2,
  G1944_i2,
  G1952_i2,
  G1850_i2,
  G1866_i2,
  G1874_i2,
  G1882_i2,
  G1890_i2,
  G1914_i2,
  G1930_i2,
  G1938_i2,
  G1946_i2,
  G1954_i2,
  G1845_i2,
  G1861_i2,
  G1869_i2,
  G1877_i2,
  G1885_i2,
  G1909_i2,
  G1925_i2,
  G1933_i2,
  G1941_i2,
  G1949_i2,
  G1846_i2,
  G1862_i2,
  G1870_i2,
  G1878_i2,
  G1886_i2,
  G1910_i2,
  G1926_i2,
  G1934_i2,
  G1942_i2,
  G1950_i2,
  G1849_i2,
  G1865_i2,
  G1873_i2,
  G1881_i2,
  G1889_i2,
  G1913_i2,
  G1929_i2,
  G1937_i2,
  G1945_i2,
  G1953_i2,
  G1843_i2,
  G1859_i2,
  G1867_i2,
  G1875_i2,
  G1883_i2,
  G1907_i2,
  G1923_i2,
  G1931_i2,
  G1939_i2,
  G1947_i2,
  G1844_i2,
  G1860_i2,
  G1868_i2,
  G1876_i2,
  G1884_i2,
  G1908_i2,
  G1924_i2,
  G1932_i2,
  G1940_i2,
  G1948_i2,
  G1847_i2,
  G1863_i2,
  G1871_i2,
  G1879_i2,
  G1887_i2,
  G1911_i2,
  G1927_i2,
  G1935_i2,
  G1943_i2,
  G1951_i2,
  G2444_i2,
  G2451_i2,
  G2502_i2,
  G2507_i2,
  G2515_i2,
  G2583_i2,
  n1797_lo_buf_i2,
  n1833_lo_buf_i2,
  n1881_lo_buf_i2,
  G523_i2,
  G575_i2,
  G578_i2,
  G615_i2,
  G2254_i2,
  G2255_i2,
  G2027_i2,
  G2393_i2,
  G527_i2,
  G594_i2,
  G1689_i2,
  G1693_i2,
  G2281_i2,
  G2014_i2,
  G2459_i2,
  G2561_i2,
  G2533_i2,
  n1749_lo_buf_i2,
  n1761_lo_buf_i2,
  n1773_lo_buf_i2,
  n1809_lo_buf_i2,
  G1955_i2,
  G1958_i2,
  G2562_i2,
  G2398_i2,
  G2524_i2,
  G2563_i2,
  G2577_i2,
  G2627_i2,
  G654_i2,
  G660_i2,
  G831_i2,
  G919_i2,
  G925_i2,
  n1815_lo_buf_i2,
  n1899_lo_buf_i2,
  n2079_lo_buf_i2,
  n2127_lo_buf_i2,
  n2139_lo_buf_i2,
  n2151_lo_buf_i2,
  n2187_lo_buf_i2,
  n2199_lo_buf_i2,
  n2211_lo_buf_i2,
  G533_i2,
  n1854_lo_buf_i2,
  n2094_lo_buf_i2,
  G667_i2,
  G874_i2,
  G851_i2,
  G1127_i2,
  n1869_lo_buf_i2,
  n2109_lo_buf_i2,
  n2121_lo_buf_i2,
  G477_i2,
  G491_i2,
  G501_i2,
  G786_i2,
  G791_i2,
  G1126_i2,
  G1052_i2,
  G1054_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input G42;input G43;input G44;input G45;input G46;input G47;input G48;input G49;input G50;input n1836_lo;input n1872_lo;input n1884_lo;input n1911_lo;input n1914_lo;input n1917_lo;input n1923_lo;input n1926_lo;input n1929_lo;input n1935_lo;input n1938_lo;input n1947_lo;input n1950_lo;input n1959_lo;input n1962_lo;input n1971_lo;input n1974_lo;input n1983_lo;input n1995_lo;input n2007_lo;input n2019_lo;input n2031_lo;input n2043_lo;input n2055_lo;input n2064_lo;input n2067_lo;input n2100_lo;input n2112_lo;input n2124_lo;input n2136_lo;input n2148_lo;input n2160_lo;input n2163_lo;input n2172_lo;input n2175_lo;input n2184_lo;input n2223_lo;input n2235_lo;input n2238_lo;input n2247_lo;input n2250_lo;input n2259_lo;input n2262_lo;input n2271_lo;input n2274_lo;input n2283_lo;input n2286_lo;input n2295_lo;input n2298_lo;input n2304_lo;input n2307_lo;input n2331_lo;input n2334_lo;input n2337_lo;input n2340_lo;input n3241_o2;input n3242_o2;input n3610_o2;input n3980_o2;input n3968_o2;input n4298_o2;input n4371_o2;input n4413_o2;input n4418_o2;input n4628_o2;input n4629_o2;input n4633_o2;input n4634_o2;input n4732_o2;input n4733_o2;input n4884_o2;input n4886_o2;input n4890_o2;input n5011_o2;input n5012_o2;input n5013_o2;input n5014_o2;input n5015_o2;input n5021_o2;input n5016_o2;input n5026_o2;input n4377_o2;input n4378_o2;input n4389_o2;input n327_inv;input n330_inv;input n4398_o2;input n4401_o2;input n5117_o2;input n5115_o2;input n5122_o2;input n5121_o2;input n5119_o2;input n5116_o2;input n5123_o2;input n5156_o2;input n5167_o2;input n4454_o2;input n4455_o2;input n4456_o2;input n4505_o2;input G742_o2;input G727_o2;input n4567_o2;input n4568_o2;input n4569_o2;input n4571_o2;input n4572_o2;input n399_inv;input n4539_o2;input n4651_o2;input n4652_o2;input n4653_o2;input G1514_o2;input G1823_o2;input n4783_o2;input n4787_o2;input n426_inv;input n429_inv;input n4816_o2;input n435_inv;input G572_o2;input n4919_o2;input n4920_o2;input n4921_o2;input G1048_o2;input n5041_o2;input n5094_o2;input n5278_o2;input n5301_o2;input G2610_o2;input G3174_o2;input G3146_o2;input G3217_o2;input G3220_o2;input G2839_o2;input G3251_o2;input G3042_o2;input G3045_o2;input G3262_o2;input G2845_o2;input G2929_o2;input G2848_o2;input G2851_o2;input G3291_o2;input G3254_o2;input G2666_o2;input n5099_o2;input n5100_o2;input n5101_o2;input G2558_o2;input n5266_o2;input n5267_o2;input G2759_o2;input n537_inv;input n540_inv;input n543_inv;input n5292_o2;input n5293_o2;input n5294_o2;input n5295_o2;input G618_o2;input G621_o2;input G384_o2;input G377_o2;input n570_inv;input G3171_o2;input G2552_o2;input G3272_o2;input G2015_o2;input G3294_o2;input G3281_o2;input G3320_o2;input G3275_o2;input G3140_o2;input G2836_o2;input G2926_o2;input G2842_o2;input G3302_o2;input G3288_o2;input G3143_o2;input G3100_o2;input G2512_o2;input n5325_o2;input n5326_o2;input n5327_o2;input n1857_lo_buf_o2;input n2097_lo_buf_o2;input G2669_o2;input n642_inv;input G568_o2;input n648_inv;input G565_o2;input G559_o2;input n1821_lo_buf_o2;input n1905_lo_buf_o2;input n2133_lo_buf_o2;input n2145_lo_buf_o2;input n2157_lo_buf_o2;input n2205_lo_buf_o2;input n2217_lo_buf_o2;input G447_o2;input G434_o2;input G422_o2;input G461_o2;input G3312_o2;input G3332_o2;input G3195_o2;input G2607_o2;input n702_inv;input G1005_o2;input G1008_o2;input n2001_lo_buf_o2;input n2169_lo_buf_o2;input n2229_lo_buf_o2;input n2301_lo_buf_o2;input n723_inv;input G2947_o2;input n2013_lo_buf_o2;input n2025_lo_buf_o2;input n2037_lo_buf_o2;input n2049_lo_buf_o2;input n2181_lo_buf_o2;input n744_inv;input n747_inv;input n750_inv;input n753_inv;input G3350_o2;input G3360_o2;input G3373_o2;input G3237_o2;input G2773_o2;input G1733_o2;input G1738_o2;input G1751_o2;input G2216_o2;input G2219_o2;input n786_inv;input n789_inv;input G787_o2;input G2823_o2;input G2796_o2;input G875_o2;input G2208_o2;input G2211_o2;input n1989_lo_buf_o2;input n2061_lo_buf_o2;input n2313_lo_buf_o2;input G2232_o2;input G1725_o2;input G1764_o2;input G2356_o2;input G2359_o2;input G1180_o2;input G1756_o2;input G2441_o2;input G2887_o2;input G2991_o2;input n849_inv;input n852_inv;input n855_inv;input n858_inv;input n861_inv;input G2805_o2;input G2906_o2;input G2833_o2;input n873_inv;input G3353_o2;input G3367_o2;input G3346_o2;input G3340_o2;input G3376_o2;input G3359_o2;input G3240_o2;input G3344_o2;input G2880_o2;input G2939_o2;input G2248_o2;input G2251_o2;input G2021_o2;input G3383_o2;input G3399_o2;input G3404_o2;input G3265_o2;input G2866_o2;input G2999_o2;input G736_o2;input G739_o2;input G1200_o2;input G1203_o2;input G3027_o2;input G1463_o2;input G1460_o2;input G3012_o2;input G1574_o2;input G1646_o2;input G1592_o2;input G1664_o2;input G1547_o2;input G1619_o2;input G1556_o2;input G1628_o2;input G1583_o2;input G1655_o2;input G1529_o2;input G1601_o2;input G1538_o2;input G1610_o2;input G1565_o2;input G1637_o2;input G2437_o2;input n1008_inv;input n1785_lo_buf_o2;input n1845_lo_buf_o2;input n1893_lo_buf_o2;input n1941_lo_buf_o2;input n1953_lo_buf_o2;input n1965_lo_buf_o2;input n1977_lo_buf_o2;input n2241_lo_buf_o2;input n2253_lo_buf_o2;input n2265_lo_buf_o2;input n2277_lo_buf_o2;input n2289_lo_buf_o2;input G519_o2;input n1050_inv;input n1053_inv;input n1056_inv;input G1318_o2;input n1062_inv;input G593_o2;input n1068_inv;input n1071_inv;input n1074_inv;input G2284_o2;input G2580_o2;input G2302_o2;input G2598_o2;input G2497_o2;input G2651_o2;input G2296_o2;input G2308_o2;input G2592_o2;input G2604_o2;input G2902_o2;input G2975_o2;input G2962_o2;input G3069_o2;input G2018_o2;input G1176_o2;input G1189_o2;input G3066_o2;input G3137_o2;input G3038_o2;input G3117_o2;input G2384_o2;input G2472_o2;input G772_o2;input G935_o2;input G2923_o2;input G2971_o2;input G2980_o2;input G3039_o2;input G2388_o2;input G2287_o2;input G3024_o2;input G2916_o2;input n1176_inv;input G3035_o2;input G3107_o2;input G1023_o2;input G1024_o2;input G1311_o2;input G1312_o2;input G3063_o2;input G1520_o2;input G1519_o2;input G3078_o2;input G2038_o2;input G1848_o2;input G1864_o2;input G1872_o2;input G1880_o2;input G1888_o2;input G1912_o2;input G1928_o2;input G1936_o2;input G1944_o2;input G1952_o2;input G1850_o2;input G1866_o2;input G1874_o2;input G1882_o2;input G1890_o2;input G1914_o2;input G1930_o2;input G1938_o2;input G1946_o2;input G1954_o2;input G1845_o2;input G1861_o2;input G1869_o2;input G1877_o2;input G1885_o2;input G1909_o2;input G1925_o2;input G1933_o2;input G1941_o2;input G1949_o2;input G1846_o2;input G1862_o2;input G1870_o2;input G1878_o2;input G1886_o2;input G1910_o2;input G1926_o2;input G1934_o2;input G1942_o2;input G1950_o2;input G1849_o2;input G1865_o2;input G1873_o2;input G1881_o2;input G1889_o2;input G1913_o2;input G1929_o2;input G1937_o2;input G1945_o2;input G1953_o2;input G1843_o2;input G1859_o2;input G1867_o2;input G1875_o2;input G1883_o2;input G1907_o2;input G1923_o2;input G1931_o2;input G1939_o2;input G1947_o2;input G1844_o2;input G1860_o2;input G1868_o2;input G1876_o2;input G1884_o2;input G1908_o2;input G1924_o2;input G1932_o2;input G1940_o2;input G1948_o2;input G1847_o2;input G1863_o2;input G1871_o2;input G1879_o2;input G1887_o2;input G1911_o2;input G1927_o2;input G1935_o2;input G1943_o2;input G1951_o2;input G2444_o2;input G2451_o2;input G2502_o2;input G2507_o2;input n1464_inv;input G2583_o2;input n1797_lo_buf_o2;input n1833_lo_buf_o2;input n1881_lo_buf_o2;input n1479_inv;input n1482_inv;input n1485_inv;input G615_o2;input G2254_o2;input G2255_o2;input G2027_o2;input G2393_o2;input G527_o2;input G594_o2;input G1689_o2;input G1693_o2;input G2281_o2;input G2014_o2;input G2459_o2;input G2561_o2;input G2533_o2;input n1749_lo_buf_o2;input n1761_lo_buf_o2;input n1773_lo_buf_o2;input n1809_lo_buf_o2;input G1955_o2;input G1958_o2;input G2562_o2;input G2398_o2;input n1554_inv;input n1557_inv;input G2577_o2;input G2627_o2;input G654_o2;input G660_o2;input G831_o2;input G919_o2;input G925_o2;input n1815_lo_buf_o2;input n1899_lo_buf_o2;input n2079_lo_buf_o2;input n2127_lo_buf_o2;input n2139_lo_buf_o2;input n2151_lo_buf_o2;input n2187_lo_buf_o2;input n2199_lo_buf_o2;input n2211_lo_buf_o2;input G533_o2;input n1854_lo_buf_o2;input n2094_lo_buf_o2;input G667_o2;input G874_o2;input G851_o2;input G1127_o2;input n1869_lo_buf_o2;input n2109_lo_buf_o2;input n2121_lo_buf_o2;input G477_o2;input G491_o2;input G501_o2;input G786_o2;input G791_o2;input G1126_o2;input G1052_o2;input G1054_o2;
  output G3519;output G3520;output G3521;output G3522;output G3523;output G3524;output G3525;output G3526;output G3527;output G3528;output G3529;output G3530;output G3531;output G3532;output G3533;output G3534;output G3535;output G3536;output G3537;output G3538;output G3539;output G3540;output n1836_li;output n1872_li;output n1884_li;output n1911_li;output n1914_li;output n1917_li;output n1923_li;output n1926_li;output n1929_li;output n1935_li;output n1938_li;output n1947_li;output n1950_li;output n1959_li;output n1962_li;output n1971_li;output n1974_li;output n1983_li;output n1995_li;output n2007_li;output n2019_li;output n2031_li;output n2043_li;output n2055_li;output n2064_li;output n2067_li;output n2100_li;output n2112_li;output n2124_li;output n2136_li;output n2148_li;output n2160_li;output n2163_li;output n2172_li;output n2175_li;output n2184_li;output n2223_li;output n2235_li;output n2238_li;output n2247_li;output n2250_li;output n2259_li;output n2262_li;output n2271_li;output n2274_li;output n2283_li;output n2286_li;output n2295_li;output n2298_li;output n2304_li;output n2307_li;output n2331_li;output n2334_li;output n2337_li;output n2340_li;output n3241_i2;output n3242_i2;output n3610_i2;output n3980_i2;output n3968_i2;output n4298_i2;output n4371_i2;output n4413_i2;output n4418_i2;output n4628_i2;output n4629_i2;output n4633_i2;output n4634_i2;output n4732_i2;output n4733_i2;output n4884_i2;output n4886_i2;output n4890_i2;output n5011_i2;output n5012_i2;output n5013_i2;output n5014_i2;output n5015_i2;output n5021_i2;output n5016_i2;output n5026_i2;output n4377_i2;output n4378_i2;output n4389_i2;output n4390_i2;output n4391_i2;output n4398_i2;output n4401_i2;output n5117_i2;output n5115_i2;output n5122_i2;output n5121_i2;output n5119_i2;output n5116_i2;output n5123_i2;output n5156_i2;output n5167_i2;output n4454_i2;output n4455_i2;output n4456_i2;output n4505_i2;output G742_i2;output G727_i2;output n4567_i2;output n4568_i2;output n4569_i2;output n4571_i2;output n4572_i2;output n4537_i2;output n4539_i2;output n4651_i2;output n4652_i2;output n4653_i2;output G1514_i2;output G1823_i2;output n4783_i2;output n4787_i2;output n4808_i2;output n4815_i2;output n4816_i2;output n4822_i2;output G572_i2;output n4919_i2;output n4920_i2;output n4921_i2;output G1048_i2;output n5041_i2;output n5094_i2;output n5278_i2;output n5301_i2;output G2610_i2;output G3174_i2;output G3146_i2;output G3217_i2;output G3220_i2;output G2839_i2;output G3251_i2;output G3042_i2;output G3045_i2;output G3262_i2;output G2845_i2;output G2929_i2;output G2848_i2;output G2851_i2;output G3291_i2;output G3254_i2;output G2666_i2;output n5099_i2;output n5100_i2;output n5101_i2;output G2558_i2;output n5266_i2;output n5267_i2;output G2759_i2;output n5269_i2;output n5270_i2;output n5271_i2;output n5292_i2;output n5293_i2;output n5294_i2;output n5295_i2;output G618_i2;output G621_i2;output G384_i2;output G377_i2;output G400_i2;output G3171_i2;output G2552_i2;output G3272_i2;output G2015_i2;output G3294_i2;output G3281_i2;output G3320_i2;output G3275_i2;output G3140_i2;output G2836_i2;output G2926_i2;output G2842_i2;output G3302_i2;output G3288_i2;output G3143_i2;output G3100_i2;output G2512_i2;output n5325_i2;output n5326_i2;output n5327_i2;output n1857_lo_buf_i2;output n2097_lo_buf_i2;output G2669_i2;output G552_i2;output G568_i2;output G530_i2;output G565_i2;output G559_i2;output n1821_lo_buf_i2;output n1905_lo_buf_i2;output n2133_lo_buf_i2;output n2145_lo_buf_i2;output n2157_lo_buf_i2;output n2205_lo_buf_i2;output n2217_lo_buf_i2;output G447_i2;output G434_i2;output G422_i2;output G461_i2;output G3312_i2;output G3332_i2;output G3195_i2;output G2607_i2;output G2799_i2;output G1005_i2;output G1008_i2;output n2001_lo_buf_i2;output n2169_lo_buf_i2;output n2229_lo_buf_i2;output n2301_lo_buf_i2;output G2816_i2;output G2947_i2;output n2013_lo_buf_i2;output n2025_lo_buf_i2;output n2037_lo_buf_i2;output n2049_lo_buf_i2;output n2181_lo_buf_i2;output G546_i2;output G480_i2;output G492_i2;output G540_i2;output G3350_i2;output G3360_i2;output G3373_i2;output G3237_i2;output G2773_i2;output G1733_i2;output G1738_i2;output G1751_i2;output G2216_i2;output G2219_i2;output G381_i2;output G397_i2;output G787_i2;output G2823_i2;output G2796_i2;output G875_i2;output G2208_i2;output G2211_i2;output n1989_lo_buf_i2;output n2061_lo_buf_i2;output n2313_lo_buf_i2;output G2232_i2;output G1725_i2;output G1764_i2;output G2356_i2;output G2359_i2;output G1180_i2;output G1756_i2;output G2441_i2;output G2887_i2;output G2991_i2;output G470_i2;output G484_i2;output G496_i2;output G353_i2;output G363_i2;output G2805_i2;output G2906_i2;output G2833_i2;output G1012_i2;output G3353_i2;output G3367_i2;output G3346_i2;output G3340_i2;output G3376_i2;output G3359_i2;output G3240_i2;output G3344_i2;output G2880_i2;output G2939_i2;output G2248_i2;output G2251_i2;output G2021_i2;output G3383_i2;output G3399_i2;output G3404_i2;output G3265_i2;output G2866_i2;output G2999_i2;output G736_i2;output G739_i2;output G1200_i2;output G1203_i2;output G3027_i2;output G1463_i2;output G1460_i2;output G3012_i2;output G1574_i2;output G1646_i2;output G1592_i2;output G1664_i2;output G1547_i2;output G1619_i2;output G1556_i2;output G1628_i2;output G1583_i2;output G1655_i2;output G1529_i2;output G1601_i2;output G1538_i2;output G1610_i2;output G1565_i2;output G1637_i2;output G2437_i2;output G2518_i2;output n1785_lo_buf_i2;output n1845_lo_buf_i2;output n1893_lo_buf_i2;output n1941_lo_buf_i2;output n1953_lo_buf_i2;output n1965_lo_buf_i2;output n1977_lo_buf_i2;output n2241_lo_buf_i2;output n2253_lo_buf_i2;output n2265_lo_buf_i2;output n2277_lo_buf_i2;output n2289_lo_buf_i2;output G519_i2;output G388_i2;output G438_i2;output G368_i2;output G1318_i2;output G425_i2;output G593_i2;output G413_i2;output G404_i2;output G451_i2;output G2284_i2;output G2580_i2;output G2302_i2;output G2598_i2;output G2497_i2;output G2651_i2;output G2296_i2;output G2308_i2;output G2592_i2;output G2604_i2;output G2902_i2;output G2975_i2;output G2962_i2;output G3069_i2;output G2018_i2;output G1176_i2;output G1189_i2;output G3066_i2;output G3137_i2;output G3038_i2;output G3117_i2;output G2384_i2;output G2472_i2;output G772_i2;output G935_i2;output G2923_i2;output G2971_i2;output G2980_i2;output G3039_i2;output G2388_i2;output G2287_i2;output G3024_i2;output G2916_i2;output G1819_i2;output G3035_i2;output G3107_i2;output G1023_i2;output G1024_i2;output G1311_i2;output G1312_i2;output G3063_i2;output G1520_i2;output G1519_i2;output G3078_i2;output G2038_i2;output G1848_i2;output G1864_i2;output G1872_i2;output G1880_i2;output G1888_i2;output G1912_i2;output G1928_i2;output G1936_i2;output G1944_i2;output G1952_i2;output G1850_i2;output G1866_i2;output G1874_i2;output G1882_i2;output G1890_i2;output G1914_i2;output G1930_i2;output G1938_i2;output G1946_i2;output G1954_i2;output G1845_i2;output G1861_i2;output G1869_i2;output G1877_i2;output G1885_i2;output G1909_i2;output G1925_i2;output G1933_i2;output G1941_i2;output G1949_i2;output G1846_i2;output G1862_i2;output G1870_i2;output G1878_i2;output G1886_i2;output G1910_i2;output G1926_i2;output G1934_i2;output G1942_i2;output G1950_i2;output G1849_i2;output G1865_i2;output G1873_i2;output G1881_i2;output G1889_i2;output G1913_i2;output G1929_i2;output G1937_i2;output G1945_i2;output G1953_i2;output G1843_i2;output G1859_i2;output G1867_i2;output G1875_i2;output G1883_i2;output G1907_i2;output G1923_i2;output G1931_i2;output G1939_i2;output G1947_i2;output G1844_i2;output G1860_i2;output G1868_i2;output G1876_i2;output G1884_i2;output G1908_i2;output G1924_i2;output G1932_i2;output G1940_i2;output G1948_i2;output G1847_i2;output G1863_i2;output G1871_i2;output G1879_i2;output G1887_i2;output G1911_i2;output G1927_i2;output G1935_i2;output G1943_i2;output G1951_i2;output G2444_i2;output G2451_i2;output G2502_i2;output G2507_i2;output G2515_i2;output G2583_i2;output n1797_lo_buf_i2;output n1833_lo_buf_i2;output n1881_lo_buf_i2;output G523_i2;output G575_i2;output G578_i2;output G615_i2;output G2254_i2;output G2255_i2;output G2027_i2;output G2393_i2;output G527_i2;output G594_i2;output G1689_i2;output G1693_i2;output G2281_i2;output G2014_i2;output G2459_i2;output G2561_i2;output G2533_i2;output n1749_lo_buf_i2;output n1761_lo_buf_i2;output n1773_lo_buf_i2;output n1809_lo_buf_i2;output G1955_i2;output G1958_i2;output G2562_i2;output G2398_i2;output G2524_i2;output G2563_i2;output G2577_i2;output G2627_i2;output G654_i2;output G660_i2;output G831_i2;output G919_i2;output G925_i2;output n1815_lo_buf_i2;output n1899_lo_buf_i2;output n2079_lo_buf_i2;output n2127_lo_buf_i2;output n2139_lo_buf_i2;output n2151_lo_buf_i2;output n2187_lo_buf_i2;output n2199_lo_buf_i2;output n2211_lo_buf_i2;output G533_i2;output n1854_lo_buf_i2;output n2094_lo_buf_i2;output G667_i2;output G874_i2;output G851_i2;output G1127_i2;output n1869_lo_buf_i2;output n2109_lo_buf_i2;output n2121_lo_buf_i2;output G477_i2;output G491_i2;output G501_i2;output G786_i2;output G791_i2;output G1126_i2;output G1052_i2;output G1054_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire n1836_lo_p;
  wire n1836_lo_n;
  wire n1872_lo_p;
  wire n1872_lo_n;
  wire n1884_lo_p;
  wire n1884_lo_n;
  wire n1911_lo_p;
  wire n1911_lo_n;
  wire n1914_lo_p;
  wire n1914_lo_n;
  wire n1917_lo_p;
  wire n1917_lo_n;
  wire n1923_lo_p;
  wire n1923_lo_n;
  wire n1926_lo_p;
  wire n1926_lo_n;
  wire n1929_lo_p;
  wire n1929_lo_n;
  wire n1935_lo_p;
  wire n1935_lo_n;
  wire n1938_lo_p;
  wire n1938_lo_n;
  wire n1947_lo_p;
  wire n1947_lo_n;
  wire n1950_lo_p;
  wire n1950_lo_n;
  wire n1959_lo_p;
  wire n1959_lo_n;
  wire n1962_lo_p;
  wire n1962_lo_n;
  wire n1971_lo_p;
  wire n1971_lo_n;
  wire n1974_lo_p;
  wire n1974_lo_n;
  wire n1983_lo_p;
  wire n1983_lo_n;
  wire n1995_lo_p;
  wire n1995_lo_n;
  wire n2007_lo_p;
  wire n2007_lo_n;
  wire n2019_lo_p;
  wire n2019_lo_n;
  wire n2031_lo_p;
  wire n2031_lo_n;
  wire n2043_lo_p;
  wire n2043_lo_n;
  wire n2055_lo_p;
  wire n2055_lo_n;
  wire n2064_lo_p;
  wire n2064_lo_n;
  wire n2067_lo_p;
  wire n2067_lo_n;
  wire n2100_lo_p;
  wire n2100_lo_n;
  wire n2112_lo_p;
  wire n2112_lo_n;
  wire n2124_lo_p;
  wire n2124_lo_n;
  wire n2136_lo_p;
  wire n2136_lo_n;
  wire n2148_lo_p;
  wire n2148_lo_n;
  wire n2160_lo_p;
  wire n2160_lo_n;
  wire n2163_lo_p;
  wire n2163_lo_n;
  wire n2172_lo_p;
  wire n2172_lo_n;
  wire n2175_lo_p;
  wire n2175_lo_n;
  wire n2184_lo_p;
  wire n2184_lo_n;
  wire n2223_lo_p;
  wire n2223_lo_n;
  wire n2235_lo_p;
  wire n2235_lo_n;
  wire n2238_lo_p;
  wire n2238_lo_n;
  wire n2247_lo_p;
  wire n2247_lo_n;
  wire n2250_lo_p;
  wire n2250_lo_n;
  wire n2259_lo_p;
  wire n2259_lo_n;
  wire n2262_lo_p;
  wire n2262_lo_n;
  wire n2271_lo_p;
  wire n2271_lo_n;
  wire n2274_lo_p;
  wire n2274_lo_n;
  wire n2283_lo_p;
  wire n2283_lo_n;
  wire n2286_lo_p;
  wire n2286_lo_n;
  wire n2295_lo_p;
  wire n2295_lo_n;
  wire n2298_lo_p;
  wire n2298_lo_n;
  wire n2304_lo_p;
  wire n2304_lo_n;
  wire n2307_lo_p;
  wire n2307_lo_n;
  wire n2331_lo_p;
  wire n2331_lo_n;
  wire n2334_lo_p;
  wire n2334_lo_n;
  wire n2337_lo_p;
  wire n2337_lo_n;
  wire n2340_lo_p;
  wire n2340_lo_n;
  wire n3241_o2_p;
  wire n3241_o2_n;
  wire n3242_o2_p;
  wire n3242_o2_n;
  wire n3610_o2_p;
  wire n3610_o2_n;
  wire n3980_o2_p;
  wire n3980_o2_n;
  wire n3968_o2_p;
  wire n3968_o2_n;
  wire n4298_o2_p;
  wire n4298_o2_n;
  wire n4371_o2_p;
  wire n4371_o2_n;
  wire n4413_o2_p;
  wire n4413_o2_n;
  wire n4418_o2_p;
  wire n4418_o2_n;
  wire n4628_o2_p;
  wire n4628_o2_n;
  wire n4629_o2_p;
  wire n4629_o2_n;
  wire n4633_o2_p;
  wire n4633_o2_n;
  wire n4634_o2_p;
  wire n4634_o2_n;
  wire n4732_o2_p;
  wire n4732_o2_n;
  wire n4733_o2_p;
  wire n4733_o2_n;
  wire n4884_o2_p;
  wire n4884_o2_n;
  wire n4886_o2_p;
  wire n4886_o2_n;
  wire n4890_o2_p;
  wire n4890_o2_n;
  wire n5011_o2_p;
  wire n5011_o2_n;
  wire n5012_o2_p;
  wire n5012_o2_n;
  wire n5013_o2_p;
  wire n5013_o2_n;
  wire n5014_o2_p;
  wire n5014_o2_n;
  wire n5015_o2_p;
  wire n5015_o2_n;
  wire n5021_o2_p;
  wire n5021_o2_n;
  wire n5016_o2_p;
  wire n5016_o2_n;
  wire n5026_o2_p;
  wire n5026_o2_n;
  wire n4377_o2_p;
  wire n4377_o2_n;
  wire n4378_o2_p;
  wire n4378_o2_n;
  wire n4389_o2_p;
  wire n4389_o2_n;
  wire n327_inv_p;
  wire n327_inv_n;
  wire n330_inv_p;
  wire n330_inv_n;
  wire n4398_o2_p;
  wire n4398_o2_n;
  wire n4401_o2_p;
  wire n4401_o2_n;
  wire n5117_o2_p;
  wire n5117_o2_n;
  wire n5115_o2_p;
  wire n5115_o2_n;
  wire n5122_o2_p;
  wire n5122_o2_n;
  wire n5121_o2_p;
  wire n5121_o2_n;
  wire n5119_o2_p;
  wire n5119_o2_n;
  wire n5116_o2_p;
  wire n5116_o2_n;
  wire n5123_o2_p;
  wire n5123_o2_n;
  wire n5156_o2_p;
  wire n5156_o2_n;
  wire n5167_o2_p;
  wire n5167_o2_n;
  wire n4454_o2_p;
  wire n4454_o2_n;
  wire n4455_o2_p;
  wire n4455_o2_n;
  wire n4456_o2_p;
  wire n4456_o2_n;
  wire n4505_o2_p;
  wire n4505_o2_n;
  wire G742_o2_p;
  wire G742_o2_n;
  wire G727_o2_p;
  wire G727_o2_n;
  wire n4567_o2_p;
  wire n4567_o2_n;
  wire n4568_o2_p;
  wire n4568_o2_n;
  wire n4569_o2_p;
  wire n4569_o2_n;
  wire n4571_o2_p;
  wire n4571_o2_n;
  wire n4572_o2_p;
  wire n4572_o2_n;
  wire n399_inv_p;
  wire n399_inv_n;
  wire n4539_o2_p;
  wire n4539_o2_n;
  wire n4651_o2_p;
  wire n4651_o2_n;
  wire n4652_o2_p;
  wire n4652_o2_n;
  wire n4653_o2_p;
  wire n4653_o2_n;
  wire G1514_o2_p;
  wire G1514_o2_n;
  wire G1823_o2_p;
  wire G1823_o2_n;
  wire n4783_o2_p;
  wire n4783_o2_n;
  wire n4787_o2_p;
  wire n4787_o2_n;
  wire n426_inv_p;
  wire n426_inv_n;
  wire n429_inv_p;
  wire n429_inv_n;
  wire n4816_o2_p;
  wire n4816_o2_n;
  wire n435_inv_p;
  wire n435_inv_n;
  wire G572_o2_p;
  wire G572_o2_n;
  wire n4919_o2_p;
  wire n4919_o2_n;
  wire n4920_o2_p;
  wire n4920_o2_n;
  wire n4921_o2_p;
  wire n4921_o2_n;
  wire G1048_o2_p;
  wire G1048_o2_n;
  wire n5041_o2_p;
  wire n5041_o2_n;
  wire n5094_o2_p;
  wire n5094_o2_n;
  wire n5278_o2_p;
  wire n5278_o2_n;
  wire n5301_o2_p;
  wire n5301_o2_n;
  wire G2610_o2_p;
  wire G2610_o2_n;
  wire G3174_o2_p;
  wire G3174_o2_n;
  wire G3146_o2_p;
  wire G3146_o2_n;
  wire G3217_o2_p;
  wire G3217_o2_n;
  wire G3220_o2_p;
  wire G3220_o2_n;
  wire G2839_o2_p;
  wire G2839_o2_n;
  wire G3251_o2_p;
  wire G3251_o2_n;
  wire G3042_o2_p;
  wire G3042_o2_n;
  wire G3045_o2_p;
  wire G3045_o2_n;
  wire G3262_o2_p;
  wire G3262_o2_n;
  wire G2845_o2_p;
  wire G2845_o2_n;
  wire G2929_o2_p;
  wire G2929_o2_n;
  wire G2848_o2_p;
  wire G2848_o2_n;
  wire G2851_o2_p;
  wire G2851_o2_n;
  wire G3291_o2_p;
  wire G3291_o2_n;
  wire G3254_o2_p;
  wire G3254_o2_n;
  wire G2666_o2_p;
  wire G2666_o2_n;
  wire n5099_o2_p;
  wire n5099_o2_n;
  wire n5100_o2_p;
  wire n5100_o2_n;
  wire n5101_o2_p;
  wire n5101_o2_n;
  wire G2558_o2_p;
  wire G2558_o2_n;
  wire n5266_o2_p;
  wire n5266_o2_n;
  wire n5267_o2_p;
  wire n5267_o2_n;
  wire G2759_o2_p;
  wire G2759_o2_n;
  wire n537_inv_p;
  wire n537_inv_n;
  wire n540_inv_p;
  wire n540_inv_n;
  wire n543_inv_p;
  wire n543_inv_n;
  wire n5292_o2_p;
  wire n5292_o2_n;
  wire n5293_o2_p;
  wire n5293_o2_n;
  wire n5294_o2_p;
  wire n5294_o2_n;
  wire n5295_o2_p;
  wire n5295_o2_n;
  wire G618_o2_p;
  wire G618_o2_n;
  wire G621_o2_p;
  wire G621_o2_n;
  wire G384_o2_p;
  wire G384_o2_n;
  wire G377_o2_p;
  wire G377_o2_n;
  wire n570_inv_p;
  wire n570_inv_n;
  wire G3171_o2_p;
  wire G3171_o2_n;
  wire G2552_o2_p;
  wire G2552_o2_n;
  wire G3272_o2_p;
  wire G3272_o2_n;
  wire G2015_o2_p;
  wire G2015_o2_n;
  wire G3294_o2_p;
  wire G3294_o2_n;
  wire G3281_o2_p;
  wire G3281_o2_n;
  wire G3320_o2_p;
  wire G3320_o2_n;
  wire G3275_o2_p;
  wire G3275_o2_n;
  wire G3140_o2_p;
  wire G3140_o2_n;
  wire G2836_o2_p;
  wire G2836_o2_n;
  wire G2926_o2_p;
  wire G2926_o2_n;
  wire G2842_o2_p;
  wire G2842_o2_n;
  wire G3302_o2_p;
  wire G3302_o2_n;
  wire G3288_o2_p;
  wire G3288_o2_n;
  wire G3143_o2_p;
  wire G3143_o2_n;
  wire G3100_o2_p;
  wire G3100_o2_n;
  wire G2512_o2_p;
  wire G2512_o2_n;
  wire n5325_o2_p;
  wire n5325_o2_n;
  wire n5326_o2_p;
  wire n5326_o2_n;
  wire n5327_o2_p;
  wire n5327_o2_n;
  wire n1857_lo_buf_o2_p;
  wire n1857_lo_buf_o2_n;
  wire n2097_lo_buf_o2_p;
  wire n2097_lo_buf_o2_n;
  wire G2669_o2_p;
  wire G2669_o2_n;
  wire n642_inv_p;
  wire n642_inv_n;
  wire G568_o2_p;
  wire G568_o2_n;
  wire n648_inv_p;
  wire n648_inv_n;
  wire G565_o2_p;
  wire G565_o2_n;
  wire G559_o2_p;
  wire G559_o2_n;
  wire n1821_lo_buf_o2_p;
  wire n1821_lo_buf_o2_n;
  wire n1905_lo_buf_o2_p;
  wire n1905_lo_buf_o2_n;
  wire n2133_lo_buf_o2_p;
  wire n2133_lo_buf_o2_n;
  wire n2145_lo_buf_o2_p;
  wire n2145_lo_buf_o2_n;
  wire n2157_lo_buf_o2_p;
  wire n2157_lo_buf_o2_n;
  wire n2205_lo_buf_o2_p;
  wire n2205_lo_buf_o2_n;
  wire n2217_lo_buf_o2_p;
  wire n2217_lo_buf_o2_n;
  wire G447_o2_p;
  wire G447_o2_n;
  wire G434_o2_p;
  wire G434_o2_n;
  wire G422_o2_p;
  wire G422_o2_n;
  wire G461_o2_p;
  wire G461_o2_n;
  wire G3312_o2_p;
  wire G3312_o2_n;
  wire G3332_o2_p;
  wire G3332_o2_n;
  wire G3195_o2_p;
  wire G3195_o2_n;
  wire G2607_o2_p;
  wire G2607_o2_n;
  wire n702_inv_p;
  wire n702_inv_n;
  wire G1005_o2_p;
  wire G1005_o2_n;
  wire G1008_o2_p;
  wire G1008_o2_n;
  wire n2001_lo_buf_o2_p;
  wire n2001_lo_buf_o2_n;
  wire n2169_lo_buf_o2_p;
  wire n2169_lo_buf_o2_n;
  wire n2229_lo_buf_o2_p;
  wire n2229_lo_buf_o2_n;
  wire n2301_lo_buf_o2_p;
  wire n2301_lo_buf_o2_n;
  wire n723_inv_p;
  wire n723_inv_n;
  wire G2947_o2_p;
  wire G2947_o2_n;
  wire n2013_lo_buf_o2_p;
  wire n2013_lo_buf_o2_n;
  wire n2025_lo_buf_o2_p;
  wire n2025_lo_buf_o2_n;
  wire n2037_lo_buf_o2_p;
  wire n2037_lo_buf_o2_n;
  wire n2049_lo_buf_o2_p;
  wire n2049_lo_buf_o2_n;
  wire n2181_lo_buf_o2_p;
  wire n2181_lo_buf_o2_n;
  wire n744_inv_p;
  wire n744_inv_n;
  wire n747_inv_p;
  wire n747_inv_n;
  wire n750_inv_p;
  wire n750_inv_n;
  wire n753_inv_p;
  wire n753_inv_n;
  wire G3350_o2_p;
  wire G3350_o2_n;
  wire G3360_o2_p;
  wire G3360_o2_n;
  wire G3373_o2_p;
  wire G3373_o2_n;
  wire G3237_o2_p;
  wire G3237_o2_n;
  wire G2773_o2_p;
  wire G2773_o2_n;
  wire G1733_o2_p;
  wire G1733_o2_n;
  wire G1738_o2_p;
  wire G1738_o2_n;
  wire G1751_o2_p;
  wire G1751_o2_n;
  wire G2216_o2_p;
  wire G2216_o2_n;
  wire G2219_o2_p;
  wire G2219_o2_n;
  wire n786_inv_p;
  wire n786_inv_n;
  wire n789_inv_p;
  wire n789_inv_n;
  wire G787_o2_p;
  wire G787_o2_n;
  wire G2823_o2_p;
  wire G2823_o2_n;
  wire G2796_o2_p;
  wire G2796_o2_n;
  wire G875_o2_p;
  wire G875_o2_n;
  wire G2208_o2_p;
  wire G2208_o2_n;
  wire G2211_o2_p;
  wire G2211_o2_n;
  wire n1989_lo_buf_o2_p;
  wire n1989_lo_buf_o2_n;
  wire n2061_lo_buf_o2_p;
  wire n2061_lo_buf_o2_n;
  wire n2313_lo_buf_o2_p;
  wire n2313_lo_buf_o2_n;
  wire G2232_o2_p;
  wire G2232_o2_n;
  wire G1725_o2_p;
  wire G1725_o2_n;
  wire G1764_o2_p;
  wire G1764_o2_n;
  wire G2356_o2_p;
  wire G2356_o2_n;
  wire G2359_o2_p;
  wire G2359_o2_n;
  wire G1180_o2_p;
  wire G1180_o2_n;
  wire G1756_o2_p;
  wire G1756_o2_n;
  wire G2441_o2_p;
  wire G2441_o2_n;
  wire G2887_o2_p;
  wire G2887_o2_n;
  wire G2991_o2_p;
  wire G2991_o2_n;
  wire n849_inv_p;
  wire n849_inv_n;
  wire n852_inv_p;
  wire n852_inv_n;
  wire n855_inv_p;
  wire n855_inv_n;
  wire n858_inv_p;
  wire n858_inv_n;
  wire n861_inv_p;
  wire n861_inv_n;
  wire G2805_o2_p;
  wire G2805_o2_n;
  wire G2906_o2_p;
  wire G2906_o2_n;
  wire G2833_o2_p;
  wire G2833_o2_n;
  wire n873_inv_p;
  wire n873_inv_n;
  wire G3353_o2_p;
  wire G3353_o2_n;
  wire G3367_o2_p;
  wire G3367_o2_n;
  wire G3346_o2_p;
  wire G3346_o2_n;
  wire G3340_o2_p;
  wire G3340_o2_n;
  wire G3376_o2_p;
  wire G3376_o2_n;
  wire G3359_o2_p;
  wire G3359_o2_n;
  wire G3240_o2_p;
  wire G3240_o2_n;
  wire G3344_o2_p;
  wire G3344_o2_n;
  wire G2880_o2_p;
  wire G2880_o2_n;
  wire G2939_o2_p;
  wire G2939_o2_n;
  wire G2248_o2_p;
  wire G2248_o2_n;
  wire G2251_o2_p;
  wire G2251_o2_n;
  wire G2021_o2_p;
  wire G2021_o2_n;
  wire G3383_o2_p;
  wire G3383_o2_n;
  wire G3399_o2_p;
  wire G3399_o2_n;
  wire G3404_o2_p;
  wire G3404_o2_n;
  wire G3265_o2_p;
  wire G3265_o2_n;
  wire G2866_o2_p;
  wire G2866_o2_n;
  wire G2999_o2_p;
  wire G2999_o2_n;
  wire G736_o2_p;
  wire G736_o2_n;
  wire G739_o2_p;
  wire G739_o2_n;
  wire G1200_o2_p;
  wire G1200_o2_n;
  wire G1203_o2_p;
  wire G1203_o2_n;
  wire G3027_o2_p;
  wire G3027_o2_n;
  wire G1463_o2_p;
  wire G1463_o2_n;
  wire G1460_o2_p;
  wire G1460_o2_n;
  wire G3012_o2_p;
  wire G3012_o2_n;
  wire G1574_o2_p;
  wire G1574_o2_n;
  wire G1646_o2_p;
  wire G1646_o2_n;
  wire G1592_o2_p;
  wire G1592_o2_n;
  wire G1664_o2_p;
  wire G1664_o2_n;
  wire G1547_o2_p;
  wire G1547_o2_n;
  wire G1619_o2_p;
  wire G1619_o2_n;
  wire G1556_o2_p;
  wire G1556_o2_n;
  wire G1628_o2_p;
  wire G1628_o2_n;
  wire G1583_o2_p;
  wire G1583_o2_n;
  wire G1655_o2_p;
  wire G1655_o2_n;
  wire G1529_o2_p;
  wire G1529_o2_n;
  wire G1601_o2_p;
  wire G1601_o2_n;
  wire G1538_o2_p;
  wire G1538_o2_n;
  wire G1610_o2_p;
  wire G1610_o2_n;
  wire G1565_o2_p;
  wire G1565_o2_n;
  wire G1637_o2_p;
  wire G1637_o2_n;
  wire G2437_o2_p;
  wire G2437_o2_n;
  wire n1008_inv_p;
  wire n1008_inv_n;
  wire n1785_lo_buf_o2_p;
  wire n1785_lo_buf_o2_n;
  wire n1845_lo_buf_o2_p;
  wire n1845_lo_buf_o2_n;
  wire n1893_lo_buf_o2_p;
  wire n1893_lo_buf_o2_n;
  wire n1941_lo_buf_o2_p;
  wire n1941_lo_buf_o2_n;
  wire n1953_lo_buf_o2_p;
  wire n1953_lo_buf_o2_n;
  wire n1965_lo_buf_o2_p;
  wire n1965_lo_buf_o2_n;
  wire n1977_lo_buf_o2_p;
  wire n1977_lo_buf_o2_n;
  wire n2241_lo_buf_o2_p;
  wire n2241_lo_buf_o2_n;
  wire n2253_lo_buf_o2_p;
  wire n2253_lo_buf_o2_n;
  wire n2265_lo_buf_o2_p;
  wire n2265_lo_buf_o2_n;
  wire n2277_lo_buf_o2_p;
  wire n2277_lo_buf_o2_n;
  wire n2289_lo_buf_o2_p;
  wire n2289_lo_buf_o2_n;
  wire G519_o2_p;
  wire G519_o2_n;
  wire n1050_inv_p;
  wire n1050_inv_n;
  wire n1053_inv_p;
  wire n1053_inv_n;
  wire n1056_inv_p;
  wire n1056_inv_n;
  wire G1318_o2_p;
  wire G1318_o2_n;
  wire n1062_inv_p;
  wire n1062_inv_n;
  wire G593_o2_p;
  wire G593_o2_n;
  wire n1068_inv_p;
  wire n1068_inv_n;
  wire n1071_inv_p;
  wire n1071_inv_n;
  wire n1074_inv_p;
  wire n1074_inv_n;
  wire G2284_o2_p;
  wire G2284_o2_n;
  wire G2580_o2_p;
  wire G2580_o2_n;
  wire G2302_o2_p;
  wire G2302_o2_n;
  wire G2598_o2_p;
  wire G2598_o2_n;
  wire G2497_o2_p;
  wire G2497_o2_n;
  wire G2651_o2_p;
  wire G2651_o2_n;
  wire G2296_o2_p;
  wire G2296_o2_n;
  wire G2308_o2_p;
  wire G2308_o2_n;
  wire G2592_o2_p;
  wire G2592_o2_n;
  wire G2604_o2_p;
  wire G2604_o2_n;
  wire G2902_o2_p;
  wire G2902_o2_n;
  wire G2975_o2_p;
  wire G2975_o2_n;
  wire G2962_o2_p;
  wire G2962_o2_n;
  wire G3069_o2_p;
  wire G3069_o2_n;
  wire G2018_o2_p;
  wire G2018_o2_n;
  wire G1176_o2_p;
  wire G1176_o2_n;
  wire G1189_o2_p;
  wire G1189_o2_n;
  wire G3066_o2_p;
  wire G3066_o2_n;
  wire G3137_o2_p;
  wire G3137_o2_n;
  wire G3038_o2_p;
  wire G3038_o2_n;
  wire G3117_o2_p;
  wire G3117_o2_n;
  wire G2384_o2_p;
  wire G2384_o2_n;
  wire G2472_o2_p;
  wire G2472_o2_n;
  wire G772_o2_p;
  wire G772_o2_n;
  wire G935_o2_p;
  wire G935_o2_n;
  wire G2923_o2_p;
  wire G2923_o2_n;
  wire G2971_o2_p;
  wire G2971_o2_n;
  wire G2980_o2_p;
  wire G2980_o2_n;
  wire G3039_o2_p;
  wire G3039_o2_n;
  wire G2388_o2_p;
  wire G2388_o2_n;
  wire G2287_o2_p;
  wire G2287_o2_n;
  wire G3024_o2_p;
  wire G3024_o2_n;
  wire G2916_o2_p;
  wire G2916_o2_n;
  wire n1176_inv_p;
  wire n1176_inv_n;
  wire G3035_o2_p;
  wire G3035_o2_n;
  wire G3107_o2_p;
  wire G3107_o2_n;
  wire G1023_o2_p;
  wire G1023_o2_n;
  wire G1024_o2_p;
  wire G1024_o2_n;
  wire G1311_o2_p;
  wire G1311_o2_n;
  wire G1312_o2_p;
  wire G1312_o2_n;
  wire G3063_o2_p;
  wire G3063_o2_n;
  wire G1520_o2_p;
  wire G1520_o2_n;
  wire G1519_o2_p;
  wire G1519_o2_n;
  wire G3078_o2_p;
  wire G3078_o2_n;
  wire G2038_o2_p;
  wire G2038_o2_n;
  wire G1848_o2_p;
  wire G1848_o2_n;
  wire G1864_o2_p;
  wire G1864_o2_n;
  wire G1872_o2_p;
  wire G1872_o2_n;
  wire G1880_o2_p;
  wire G1880_o2_n;
  wire G1888_o2_p;
  wire G1888_o2_n;
  wire G1912_o2_p;
  wire G1912_o2_n;
  wire G1928_o2_p;
  wire G1928_o2_n;
  wire G1936_o2_p;
  wire G1936_o2_n;
  wire G1944_o2_p;
  wire G1944_o2_n;
  wire G1952_o2_p;
  wire G1952_o2_n;
  wire G1850_o2_p;
  wire G1850_o2_n;
  wire G1866_o2_p;
  wire G1866_o2_n;
  wire G1874_o2_p;
  wire G1874_o2_n;
  wire G1882_o2_p;
  wire G1882_o2_n;
  wire G1890_o2_p;
  wire G1890_o2_n;
  wire G1914_o2_p;
  wire G1914_o2_n;
  wire G1930_o2_p;
  wire G1930_o2_n;
  wire G1938_o2_p;
  wire G1938_o2_n;
  wire G1946_o2_p;
  wire G1946_o2_n;
  wire G1954_o2_p;
  wire G1954_o2_n;
  wire G1845_o2_p;
  wire G1845_o2_n;
  wire G1861_o2_p;
  wire G1861_o2_n;
  wire G1869_o2_p;
  wire G1869_o2_n;
  wire G1877_o2_p;
  wire G1877_o2_n;
  wire G1885_o2_p;
  wire G1885_o2_n;
  wire G1909_o2_p;
  wire G1909_o2_n;
  wire G1925_o2_p;
  wire G1925_o2_n;
  wire G1933_o2_p;
  wire G1933_o2_n;
  wire G1941_o2_p;
  wire G1941_o2_n;
  wire G1949_o2_p;
  wire G1949_o2_n;
  wire G1846_o2_p;
  wire G1846_o2_n;
  wire G1862_o2_p;
  wire G1862_o2_n;
  wire G1870_o2_p;
  wire G1870_o2_n;
  wire G1878_o2_p;
  wire G1878_o2_n;
  wire G1886_o2_p;
  wire G1886_o2_n;
  wire G1910_o2_p;
  wire G1910_o2_n;
  wire G1926_o2_p;
  wire G1926_o2_n;
  wire G1934_o2_p;
  wire G1934_o2_n;
  wire G1942_o2_p;
  wire G1942_o2_n;
  wire G1950_o2_p;
  wire G1950_o2_n;
  wire G1849_o2_p;
  wire G1849_o2_n;
  wire G1865_o2_p;
  wire G1865_o2_n;
  wire G1873_o2_p;
  wire G1873_o2_n;
  wire G1881_o2_p;
  wire G1881_o2_n;
  wire G1889_o2_p;
  wire G1889_o2_n;
  wire G1913_o2_p;
  wire G1913_o2_n;
  wire G1929_o2_p;
  wire G1929_o2_n;
  wire G1937_o2_p;
  wire G1937_o2_n;
  wire G1945_o2_p;
  wire G1945_o2_n;
  wire G1953_o2_p;
  wire G1953_o2_n;
  wire G1843_o2_p;
  wire G1843_o2_n;
  wire G1859_o2_p;
  wire G1859_o2_n;
  wire G1867_o2_p;
  wire G1867_o2_n;
  wire G1875_o2_p;
  wire G1875_o2_n;
  wire G1883_o2_p;
  wire G1883_o2_n;
  wire G1907_o2_p;
  wire G1907_o2_n;
  wire G1923_o2_p;
  wire G1923_o2_n;
  wire G1931_o2_p;
  wire G1931_o2_n;
  wire G1939_o2_p;
  wire G1939_o2_n;
  wire G1947_o2_p;
  wire G1947_o2_n;
  wire G1844_o2_p;
  wire G1844_o2_n;
  wire G1860_o2_p;
  wire G1860_o2_n;
  wire G1868_o2_p;
  wire G1868_o2_n;
  wire G1876_o2_p;
  wire G1876_o2_n;
  wire G1884_o2_p;
  wire G1884_o2_n;
  wire G1908_o2_p;
  wire G1908_o2_n;
  wire G1924_o2_p;
  wire G1924_o2_n;
  wire G1932_o2_p;
  wire G1932_o2_n;
  wire G1940_o2_p;
  wire G1940_o2_n;
  wire G1948_o2_p;
  wire G1948_o2_n;
  wire G1847_o2_p;
  wire G1847_o2_n;
  wire G1863_o2_p;
  wire G1863_o2_n;
  wire G1871_o2_p;
  wire G1871_o2_n;
  wire G1879_o2_p;
  wire G1879_o2_n;
  wire G1887_o2_p;
  wire G1887_o2_n;
  wire G1911_o2_p;
  wire G1911_o2_n;
  wire G1927_o2_p;
  wire G1927_o2_n;
  wire G1935_o2_p;
  wire G1935_o2_n;
  wire G1943_o2_p;
  wire G1943_o2_n;
  wire G1951_o2_p;
  wire G1951_o2_n;
  wire G2444_o2_p;
  wire G2444_o2_n;
  wire G2451_o2_p;
  wire G2451_o2_n;
  wire G2502_o2_p;
  wire G2502_o2_n;
  wire G2507_o2_p;
  wire G2507_o2_n;
  wire n1464_inv_p;
  wire n1464_inv_n;
  wire G2583_o2_p;
  wire G2583_o2_n;
  wire n1797_lo_buf_o2_p;
  wire n1797_lo_buf_o2_n;
  wire n1833_lo_buf_o2_p;
  wire n1833_lo_buf_o2_n;
  wire n1881_lo_buf_o2_p;
  wire n1881_lo_buf_o2_n;
  wire n1479_inv_p;
  wire n1479_inv_n;
  wire n1482_inv_p;
  wire n1482_inv_n;
  wire n1485_inv_p;
  wire n1485_inv_n;
  wire G615_o2_p;
  wire G615_o2_n;
  wire G2254_o2_p;
  wire G2254_o2_n;
  wire G2255_o2_p;
  wire G2255_o2_n;
  wire G2027_o2_p;
  wire G2027_o2_n;
  wire G2393_o2_p;
  wire G2393_o2_n;
  wire G527_o2_p;
  wire G527_o2_n;
  wire G594_o2_p;
  wire G594_o2_n;
  wire G1689_o2_p;
  wire G1689_o2_n;
  wire G1693_o2_p;
  wire G1693_o2_n;
  wire G2281_o2_p;
  wire G2281_o2_n;
  wire G2014_o2_p;
  wire G2014_o2_n;
  wire G2459_o2_p;
  wire G2459_o2_n;
  wire G2561_o2_p;
  wire G2561_o2_n;
  wire G2533_o2_p;
  wire G2533_o2_n;
  wire n1749_lo_buf_o2_p;
  wire n1749_lo_buf_o2_n;
  wire n1761_lo_buf_o2_p;
  wire n1761_lo_buf_o2_n;
  wire n1773_lo_buf_o2_p;
  wire n1773_lo_buf_o2_n;
  wire n1809_lo_buf_o2_p;
  wire n1809_lo_buf_o2_n;
  wire G1955_o2_p;
  wire G1955_o2_n;
  wire G1958_o2_p;
  wire G1958_o2_n;
  wire G2562_o2_p;
  wire G2562_o2_n;
  wire G2398_o2_p;
  wire G2398_o2_n;
  wire n1554_inv_p;
  wire n1554_inv_n;
  wire n1557_inv_p;
  wire n1557_inv_n;
  wire G2577_o2_p;
  wire G2577_o2_n;
  wire G2627_o2_p;
  wire G2627_o2_n;
  wire G654_o2_p;
  wire G654_o2_n;
  wire G660_o2_p;
  wire G660_o2_n;
  wire G831_o2_p;
  wire G831_o2_n;
  wire G919_o2_p;
  wire G919_o2_n;
  wire G925_o2_p;
  wire G925_o2_n;
  wire n1815_lo_buf_o2_p;
  wire n1815_lo_buf_o2_n;
  wire n1899_lo_buf_o2_p;
  wire n1899_lo_buf_o2_n;
  wire n2079_lo_buf_o2_p;
  wire n2079_lo_buf_o2_n;
  wire n2127_lo_buf_o2_p;
  wire n2127_lo_buf_o2_n;
  wire n2139_lo_buf_o2_p;
  wire n2139_lo_buf_o2_n;
  wire n2151_lo_buf_o2_p;
  wire n2151_lo_buf_o2_n;
  wire n2187_lo_buf_o2_p;
  wire n2187_lo_buf_o2_n;
  wire n2199_lo_buf_o2_p;
  wire n2199_lo_buf_o2_n;
  wire n2211_lo_buf_o2_p;
  wire n2211_lo_buf_o2_n;
  wire G533_o2_p;
  wire G533_o2_n;
  wire n1854_lo_buf_o2_p;
  wire n1854_lo_buf_o2_n;
  wire n2094_lo_buf_o2_p;
  wire n2094_lo_buf_o2_n;
  wire G667_o2_p;
  wire G667_o2_n;
  wire G874_o2_p;
  wire G874_o2_n;
  wire G851_o2_p;
  wire G851_o2_n;
  wire G1127_o2_p;
  wire G1127_o2_n;
  wire n1869_lo_buf_o2_p;
  wire n1869_lo_buf_o2_n;
  wire n2109_lo_buf_o2_p;
  wire n2109_lo_buf_o2_n;
  wire n2121_lo_buf_o2_p;
  wire n2121_lo_buf_o2_n;
  wire G477_o2_p;
  wire G477_o2_n;
  wire G491_o2_p;
  wire G491_o2_n;
  wire G501_o2_p;
  wire G501_o2_n;
  wire G786_o2_p;
  wire G786_o2_n;
  wire G791_o2_p;
  wire G791_o2_n;
  wire G1126_o2_p;
  wire G1126_o2_n;
  wire G1052_o2_p;
  wire G1052_o2_n;
  wire G1054_o2_p;
  wire G1054_o2_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire g693_p;
  wire g693_n;
  wire g694_p;
  wire g694_n;
  wire g695_p;
  wire g695_n;
  wire g696_p;
  wire g696_n;
  wire g697_p;
  wire g697_n;
  wire g698_p;
  wire g698_n;
  wire g699_p;
  wire g699_n;
  wire g700_p;
  wire g700_n;
  wire g701_p;
  wire g701_n;
  wire g702_p;
  wire g702_n;
  wire g703_p;
  wire g703_n;
  wire g704_p;
  wire g704_n;
  wire g705_p;
  wire g705_n;
  wire g706_p;
  wire g706_n;
  wire g707_p;
  wire g707_n;
  wire g708_p;
  wire g708_n;
  wire g709_p;
  wire g709_n;
  wire g710_p;
  wire g710_n;
  wire g711_p;
  wire g711_n;
  wire g712_p;
  wire g712_n;
  wire g713_p;
  wire g713_n;
  wire g714_p;
  wire g714_n;
  wire g715_p;
  wire g715_n;
  wire g716_p;
  wire g716_n;
  wire g717_p;
  wire g717_n;
  wire g718_p;
  wire g718_n;
  wire g719_p;
  wire g719_n;
  wire g720_p;
  wire g720_n;
  wire g721_p;
  wire g721_n;
  wire g722_p;
  wire g722_n;
  wire g723_p;
  wire g723_n;
  wire g724_p;
  wire g724_n;
  wire g725_p;
  wire g725_n;
  wire g726_p;
  wire g726_n;
  wire g727_p;
  wire g727_n;
  wire g728_p;
  wire g728_n;
  wire g729_p;
  wire g729_n;
  wire g730_p;
  wire g730_n;
  wire g731_p;
  wire g731_n;
  wire g732_p;
  wire g732_n;
  wire g733_p;
  wire g733_n;
  wire g734_p;
  wire g734_n;
  wire g735_p;
  wire g735_n;
  wire g736_p;
  wire g736_n;
  wire g737_p;
  wire g737_n;
  wire g738_p;
  wire g738_n;
  wire g739_p;
  wire g739_n;
  wire g740_p;
  wire g740_n;
  wire g741_p;
  wire g741_n;
  wire g742_p;
  wire g742_n;
  wire g743_p;
  wire g743_n;
  wire g744_p;
  wire g744_n;
  wire g745_p;
  wire g745_n;
  wire g746_p;
  wire g746_n;
  wire g747_p;
  wire g747_n;
  wire g748_p;
  wire g748_n;
  wire g749_p;
  wire g749_n;
  wire g750_p;
  wire g750_n;
  wire g751_p;
  wire g751_n;
  wire g752_p;
  wire g752_n;
  wire g753_p;
  wire g753_n;
  wire g754_p;
  wire g754_n;
  wire g755_p;
  wire g755_n;
  wire g756_p;
  wire g756_n;
  wire g757_p;
  wire g757_n;
  wire g758_p;
  wire g758_n;
  wire g759_p;
  wire g759_n;
  wire g760_p;
  wire g760_n;
  wire g761_p;
  wire g761_n;
  wire g762_p;
  wire g762_n;
  wire g763_p;
  wire g763_n;
  wire g764_p;
  wire g764_n;
  wire g765_p;
  wire g765_n;
  wire g766_p;
  wire g766_n;
  wire g767_p;
  wire g767_n;
  wire g768_p;
  wire g768_n;
  wire g769_p;
  wire g769_n;
  wire g770_p;
  wire g770_n;
  wire g771_p;
  wire g771_n;
  wire g772_p;
  wire g772_n;
  wire g773_p;
  wire g773_n;
  wire g774_p;
  wire g774_n;
  wire g775_p;
  wire g775_n;
  wire g776_p;
  wire g776_n;
  wire g777_p;
  wire g777_n;
  wire g778_p;
  wire g778_n;
  wire g779_p;
  wire g779_n;
  wire g780_p;
  wire g780_n;
  wire g781_p;
  wire g781_n;
  wire g782_p;
  wire g782_n;
  wire g783_p;
  wire g783_n;
  wire g784_p;
  wire g784_n;
  wire g785_p;
  wire g785_n;
  wire g786_p;
  wire g786_n;
  wire g787_p;
  wire g787_n;
  wire g788_p;
  wire g788_n;
  wire g789_p;
  wire g789_n;
  wire g790_p;
  wire g790_n;
  wire g791_p;
  wire g791_n;
  wire g792_p;
  wire g792_n;
  wire g793_p;
  wire g793_n;
  wire g794_p;
  wire g794_n;
  wire g795_p;
  wire g795_n;
  wire g796_p;
  wire g796_n;
  wire g797_p;
  wire g797_n;
  wire g798_p;
  wire g798_n;
  wire g799_p;
  wire g799_n;
  wire g800_p;
  wire g800_n;
  wire g801_p;
  wire g801_n;
  wire g802_p;
  wire g802_n;
  wire g803_p;
  wire g803_n;
  wire g804_p;
  wire g804_n;
  wire g805_p;
  wire g805_n;
  wire g806_p;
  wire g806_n;
  wire g807_p;
  wire g807_n;
  wire g808_p;
  wire g808_n;
  wire g809_p;
  wire g809_n;
  wire g810_p;
  wire g810_n;
  wire g811_p;
  wire g811_n;
  wire g812_p;
  wire g812_n;
  wire g813_p;
  wire g813_n;
  wire g814_p;
  wire g814_n;
  wire g815_p;
  wire g815_n;
  wire g816_p;
  wire g816_n;
  wire g817_p;
  wire g817_n;
  wire g818_p;
  wire g818_n;
  wire g819_p;
  wire g819_n;
  wire g820_p;
  wire g820_n;
  wire g821_p;
  wire g821_n;
  wire g822_p;
  wire g822_n;
  wire g823_p;
  wire g823_n;
  wire g824_p;
  wire g824_n;
  wire g825_p;
  wire g825_n;
  wire g826_p;
  wire g826_n;
  wire g827_p;
  wire g827_n;
  wire g828_p;
  wire g828_n;
  wire g829_p;
  wire g829_n;
  wire g830_p;
  wire g830_n;
  wire g831_p;
  wire g831_n;
  wire g832_p;
  wire g832_n;
  wire g833_p;
  wire g833_n;
  wire g834_p;
  wire g834_n;
  wire g835_p;
  wire g835_n;
  wire g836_p;
  wire g836_n;
  wire g837_p;
  wire g837_n;
  wire g838_p;
  wire g838_n;
  wire g839_p;
  wire g839_n;
  wire g840_p;
  wire g840_n;
  wire g841_p;
  wire g841_n;
  wire g842_p;
  wire g842_n;
  wire g843_p;
  wire g843_n;
  wire g844_p;
  wire g844_n;
  wire g845_p;
  wire g845_n;
  wire g846_p;
  wire g846_n;
  wire g847_p;
  wire g847_n;
  wire g848_p;
  wire g848_n;
  wire g849_p;
  wire g849_n;
  wire g850_p;
  wire g850_n;
  wire g851_p;
  wire g851_n;
  wire g852_p;
  wire g852_n;
  wire g853_p;
  wire g853_n;
  wire g854_p;
  wire g854_n;
  wire g855_p;
  wire g855_n;
  wire g856_p;
  wire g856_n;
  wire g857_p;
  wire g857_n;
  wire g858_p;
  wire g858_n;
  wire g859_p;
  wire g859_n;
  wire g860_p;
  wire g860_n;
  wire g861_p;
  wire g861_n;
  wire g862_p;
  wire g862_n;
  wire g863_p;
  wire g863_n;
  wire g864_p;
  wire g864_n;
  wire g865_p;
  wire g865_n;
  wire g866_p;
  wire g866_n;
  wire g867_p;
  wire g867_n;
  wire g868_p;
  wire g868_n;
  wire g869_p;
  wire g869_n;
  wire g870_p;
  wire g870_n;
  wire g871_p;
  wire g871_n;
  wire g872_p;
  wire g872_n;
  wire g873_p;
  wire g873_n;
  wire g874_p;
  wire g874_n;
  wire g875_p;
  wire g875_n;
  wire g876_p;
  wire g876_n;
  wire g877_p;
  wire g877_n;
  wire g878_p;
  wire g878_n;
  wire g879_p;
  wire g879_n;
  wire g880_p;
  wire g880_n;
  wire g881_p;
  wire g881_n;
  wire g882_p;
  wire g882_n;
  wire g883_p;
  wire g883_n;
  wire g884_p;
  wire g884_n;
  wire g885_p;
  wire g885_n;
  wire g886_p;
  wire g886_n;
  wire g887_p;
  wire g887_n;
  wire g888_p;
  wire g888_n;
  wire g889_p;
  wire g889_n;
  wire g890_p;
  wire g890_n;
  wire g891_p;
  wire g891_n;
  wire g892_p;
  wire g892_n;
  wire g893_p;
  wire g893_n;
  wire g894_p;
  wire g894_n;
  wire g895_p;
  wire g895_n;
  wire g896_p;
  wire g896_n;
  wire g897_p;
  wire g897_n;
  wire g898_p;
  wire g898_n;
  wire g899_p;
  wire g899_n;
  wire g900_p;
  wire g900_n;
  wire g901_p;
  wire g901_n;
  wire g902_p;
  wire g902_n;
  wire g903_p;
  wire g903_n;
  wire g904_p;
  wire g904_n;
  wire g905_p;
  wire g905_n;
  wire g906_p;
  wire g906_n;
  wire g907_p;
  wire g907_n;
  wire g908_p;
  wire g908_n;
  wire g909_p;
  wire g909_n;
  wire g910_p;
  wire g910_n;
  wire g911_p;
  wire g911_n;
  wire g912_p;
  wire g912_n;
  wire g913_p;
  wire g913_n;
  wire g914_p;
  wire g914_n;
  wire g915_p;
  wire g915_n;
  wire g916_p;
  wire g916_n;
  wire g917_p;
  wire g917_n;
  wire g918_p;
  wire g918_n;
  wire g919_p;
  wire g919_n;
  wire g920_p;
  wire g920_n;
  wire g921_p;
  wire g921_n;
  wire g922_p;
  wire g922_n;
  wire g923_p;
  wire g923_n;
  wire g924_p;
  wire g924_n;
  wire g925_p;
  wire g925_n;
  wire g926_p;
  wire g926_n;
  wire g927_p;
  wire g927_n;
  wire g928_p;
  wire g928_n;
  wire g929_p;
  wire g929_n;
  wire g930_p;
  wire g930_n;
  wire g931_p;
  wire g931_n;
  wire g932_p;
  wire g932_n;
  wire g933_p;
  wire g933_n;
  wire g934_p;
  wire g934_n;
  wire g935_p;
  wire g935_n;
  wire g936_p;
  wire g936_n;
  wire g937_p;
  wire g937_n;
  wire g938_p;
  wire g938_n;
  wire g939_p;
  wire g939_n;
  wire g940_p;
  wire g940_n;
  wire g941_p;
  wire g941_n;
  wire g942_p;
  wire g942_n;
  wire g943_p;
  wire g943_n;
  wire g944_p;
  wire g944_n;
  wire g945_p;
  wire g945_n;
  wire g946_p;
  wire g946_n;
  wire g947_p;
  wire g947_n;
  wire g948_p;
  wire g948_n;
  wire g949_p;
  wire g949_n;
  wire g950_p;
  wire g950_n;
  wire g951_p;
  wire g951_n;
  wire g952_p;
  wire g952_n;
  wire g953_p;
  wire g953_n;
  wire g954_p;
  wire g954_n;
  wire g955_p;
  wire g955_n;
  wire g956_p;
  wire g956_n;
  wire g957_p;
  wire g957_n;
  wire g958_p;
  wire g958_n;
  wire g959_p;
  wire g959_n;
  wire g960_p;
  wire g960_n;
  wire g961_p;
  wire g961_n;
  wire g962_p;
  wire g962_n;
  wire g963_p;
  wire g963_n;
  wire g964_p;
  wire g964_n;
  wire g965_p;
  wire g965_n;
  wire g966_p;
  wire g966_n;
  wire g967_p;
  wire g967_n;
  wire g968_p;
  wire g968_n;
  wire g969_p;
  wire g969_n;
  wire g970_p;
  wire g970_n;
  wire g971_p;
  wire g971_n;
  wire g972_p;
  wire g972_n;
  wire g973_p;
  wire g973_n;
  wire g974_p;
  wire g974_n;
  wire g975_p;
  wire g975_n;
  wire g976_p;
  wire g976_n;
  wire g977_p;
  wire g977_n;
  wire g978_p;
  wire g978_n;
  wire g979_p;
  wire g979_n;
  wire g980_p;
  wire g980_n;
  wire g981_p;
  wire g981_n;
  wire g982_p;
  wire g982_n;
  wire g983_p;
  wire g983_n;
  wire g984_p;
  wire g984_n;
  wire g985_p;
  wire g985_n;
  wire g986_p;
  wire g986_n;
  wire g987_p;
  wire g987_n;
  wire g988_p;
  wire g988_n;
  wire g989_p;
  wire g989_n;
  wire g990_p;
  wire g990_n;
  wire g991_p;
  wire g991_n;
  wire g992_p;
  wire g992_n;
  wire g993_p;
  wire g993_n;
  wire g994_p;
  wire g994_n;
  wire g995_p;
  wire g995_n;
  wire g996_p;
  wire g996_n;
  wire g997_p;
  wire g997_n;
  wire g998_p;
  wire g998_n;
  wire g999_p;
  wire g999_n;
  wire g1000_p;
  wire g1000_n;
  wire g1001_p;
  wire g1001_n;
  wire g1002_p;
  wire g1002_n;
  wire g1003_p;
  wire g1003_n;
  wire g1004_p;
  wire g1004_n;
  wire g1005_p;
  wire g1005_n;
  wire g1006_p;
  wire g1006_n;
  wire g1007_p;
  wire g1007_n;
  wire g1008_p;
  wire g1008_n;
  wire g1009_p;
  wire g1009_n;
  wire g1010_p;
  wire g1010_n;
  wire g1011_p;
  wire g1011_n;
  wire g1012_p;
  wire g1012_n;
  wire g1013_p;
  wire g1013_n;
  wire g1014_p;
  wire g1014_n;
  wire g1015_p;
  wire g1015_n;
  wire g1016_p;
  wire g1016_n;
  wire g1017_p;
  wire g1017_n;
  wire g1018_p;
  wire g1018_n;
  wire g1019_p;
  wire g1019_n;
  wire g1020_p;
  wire g1020_n;
  wire g1021_p;
  wire g1021_n;
  wire g1022_p;
  wire g1022_n;
  wire g1023_p;
  wire g1023_n;
  wire g1024_p;
  wire g1024_n;
  wire g1025_p;
  wire g1025_n;
  wire g1026_p;
  wire g1026_n;
  wire g1027_p;
  wire g1027_n;
  wire g1028_p;
  wire g1028_n;
  wire g1029_p;
  wire g1029_n;
  wire g1030_p;
  wire g1030_n;
  wire g1031_p;
  wire g1031_n;
  wire g1032_p;
  wire g1032_n;
  wire g1033_p;
  wire g1033_n;
  wire g1034_p;
  wire g1034_n;
  wire g1035_p;
  wire g1035_n;
  wire g1036_p;
  wire g1036_n;
  wire g1037_p;
  wire g1037_n;
  wire g1038_p;
  wire g1038_n;
  wire g1039_p;
  wire g1039_n;
  wire g1040_p;
  wire g1040_n;
  wire g1041_p;
  wire g1041_n;
  wire g1042_p;
  wire g1042_n;
  wire g1043_p;
  wire g1043_n;
  wire g1044_p;
  wire g1044_n;
  wire g1045_p;
  wire g1045_n;
  wire g1046_p;
  wire g1046_n;
  wire g1047_p;
  wire g1047_n;
  wire g1048_p;
  wire g1048_n;
  wire g1049_p;
  wire g1049_n;
  wire g1050_p;
  wire g1050_n;
  wire g1051_p;
  wire g1051_n;
  wire g1052_p;
  wire g1052_n;
  wire g1053_p;
  wire g1053_n;
  wire g1054_p;
  wire g1054_n;
  wire g1055_p;
  wire g1055_n;
  wire g1056_p;
  wire g1056_n;
  wire g1057_p;
  wire g1057_n;
  wire g1058_p;
  wire g1058_n;
  wire g1059_p;
  wire g1059_n;
  wire g1060_p;
  wire g1060_n;
  wire g1061_p;
  wire g1061_n;
  wire g1062_p;
  wire g1062_n;
  wire g1063_p;
  wire g1063_n;
  wire g1064_p;
  wire g1064_n;
  wire g1065_p;
  wire g1065_n;
  wire g1066_p;
  wire g1066_n;
  wire g1067_p;
  wire g1067_n;
  wire g1068_p;
  wire g1068_n;
  wire g1069_p;
  wire g1069_n;
  wire g1070_p;
  wire g1070_n;
  wire g1071_p;
  wire g1071_n;
  wire g1072_p;
  wire g1072_n;
  wire g1073_p;
  wire g1073_n;
  wire g1074_p;
  wire g1074_n;
  wire g1075_p;
  wire g1075_n;
  wire g1076_p;
  wire g1076_n;
  wire g1077_p;
  wire g1077_n;
  wire g1078_p;
  wire g1078_n;
  wire g1079_p;
  wire g1079_n;
  wire g1080_p;
  wire g1080_n;
  wire g1081_p;
  wire g1081_n;
  wire g1082_p;
  wire g1082_n;
  wire g1083_p;
  wire g1083_n;
  wire g1084_p;
  wire g1084_n;
  wire g1085_p;
  wire g1085_n;
  wire g1086_p;
  wire g1086_n;
  wire g1087_p;
  wire g1087_n;
  wire g1088_p;
  wire g1088_n;
  wire g1089_p;
  wire g1089_n;
  wire g1090_p;
  wire g1090_n;
  wire g1091_p;
  wire g1091_n;
  wire g1092_p;
  wire g1092_n;
  wire g1093_p;
  wire g1093_n;
  wire g1094_p;
  wire g1094_n;
  wire g1095_p;
  wire g1095_n;
  wire g1096_p;
  wire g1096_n;
  wire g1097_p;
  wire g1097_n;
  wire g1098_p;
  wire g1098_n;
  wire g1099_p;
  wire g1099_n;
  wire g1100_p;
  wire g1100_n;
  wire g1101_p;
  wire g1101_n;
  wire g1102_p;
  wire g1102_n;
  wire g1103_p;
  wire g1103_n;
  wire g1104_p;
  wire g1104_n;
  wire g1105_p;
  wire g1105_n;
  wire g1106_p;
  wire g1106_n;
  wire g1107_p;
  wire g1107_n;
  wire g1108_p;
  wire g1108_n;
  wire g1109_p;
  wire g1109_n;
  wire g1110_p;
  wire g1110_n;
  wire g1111_p;
  wire g1111_n;
  wire g1112_p;
  wire g1112_n;
  wire g1113_p;
  wire g1113_n;
  wire g1114_p;
  wire g1114_n;
  wire g1115_p;
  wire g1115_n;
  wire g1116_p;
  wire g1116_n;
  wire g1117_p;
  wire g1117_n;
  wire g1118_p;
  wire g1118_n;
  wire g1119_p;
  wire g1119_n;
  wire g1120_p;
  wire g1120_n;
  wire g1121_p;
  wire g1121_n;
  wire g1122_p;
  wire g1122_n;
  wire g1123_p;
  wire g1123_n;
  wire g1124_p;
  wire g1124_n;
  wire g1125_p;
  wire g1125_n;
  wire g1126_p;
  wire g1126_n;
  wire g1127_p;
  wire g1127_n;
  wire g1128_p;
  wire g1128_n;
  wire g1129_p;
  wire g1129_n;
  wire g1130_p;
  wire g1130_n;
  wire g1131_p;
  wire g1131_n;
  wire g1132_p;
  wire g1132_n;
  wire g1133_p;
  wire g1133_n;
  wire g1134_p;
  wire g1134_n;
  wire g1135_p;
  wire g1135_n;
  wire g1136_p;
  wire g1136_n;
  wire g1137_p;
  wire g1137_n;
  wire g1138_p;
  wire g1138_n;
  wire g1139_p;
  wire g1139_n;
  wire g1140_p;
  wire g1140_n;
  wire g1141_p;
  wire g1141_n;
  wire g1142_p;
  wire g1142_n;
  wire g1143_p;
  wire g1143_n;
  wire g1144_p;
  wire g1144_n;
  wire g1145_p;
  wire g1145_n;
  wire g1146_p;
  wire g1146_n;
  wire g1147_p;
  wire g1147_n;
  wire g1148_p;
  wire g1148_n;
  wire g1149_p;
  wire g1149_n;
  wire g1150_p;
  wire g1150_n;
  wire g1151_p;
  wire g1151_n;
  wire g1152_p;
  wire g1152_n;
  wire g1153_p;
  wire g1153_n;
  wire g1154_p;
  wire g1154_n;
  wire g1155_p;
  wire g1155_n;
  wire g1156_p;
  wire g1156_n;
  wire g1157_p;
  wire g1157_n;
  wire g1158_p;
  wire g1158_n;
  wire g1159_p;
  wire g1159_n;
  wire g1160_p;
  wire g1160_n;
  wire g1161_p;
  wire g1161_n;
  wire g1162_p;
  wire g1162_n;
  wire g1163_p;
  wire g1163_n;
  wire g1164_p;
  wire g1164_n;
  wire g1165_p;
  wire g1165_n;
  wire g1166_p;
  wire g1166_n;
  wire g1167_p;
  wire g1167_n;
  wire g1168_p;
  wire g1168_n;
  wire g1169_p;
  wire g1169_n;
  wire g1170_p;
  wire g1170_n;
  wire g1171_p;
  wire g1171_n;
  wire g1172_p;
  wire g1172_n;
  wire g1173_p;
  wire g1173_n;
  wire g1174_p;
  wire g1174_n;
  wire g1175_p;
  wire g1175_n;
  wire g1176_p;
  wire g1176_n;
  wire g1177_p;
  wire g1177_n;
  wire g1178_p;
  wire g1178_n;
  wire g1179_p;
  wire g1179_n;
  wire g1180_p;
  wire g1180_n;
  wire g1181_p;
  wire g1181_n;
  wire g1182_p;
  wire g1182_n;
  wire g1183_p;
  wire g1183_n;
  wire g1184_p;
  wire g1184_n;
  wire g1185_p;
  wire g1185_n;
  wire g1186_p;
  wire g1186_n;
  wire g1187_p;
  wire g1187_n;
  wire g1188_p;
  wire g1188_n;
  wire g1189_p;
  wire g1189_n;
  wire g1190_p;
  wire g1190_n;
  wire g1191_p;
  wire g1191_n;
  wire g1192_p;
  wire g1192_n;
  wire g1193_p;
  wire g1193_n;
  wire g1194_p;
  wire g1194_n;
  wire g1195_p;
  wire g1195_n;
  wire g1196_p;
  wire g1196_n;
  wire g1197_p;
  wire g1197_n;
  wire g1198_p;
  wire g1198_n;
  wire g1199_p;
  wire g1199_n;
  wire g1200_p;
  wire g1200_n;
  wire g1201_p;
  wire g1201_n;
  wire g1202_p;
  wire g1202_n;
  wire g1203_p;
  wire g1203_n;
  wire g1204_p;
  wire g1204_n;
  wire g1205_p;
  wire g1205_n;
  wire g1206_p;
  wire g1206_n;
  wire g1207_p;
  wire g1207_n;
  wire g1208_p;
  wire g1208_n;
  wire g1209_p;
  wire g1209_n;
  wire g1210_p;
  wire g1210_n;
  wire g1211_p;
  wire g1211_n;
  wire g1212_p;
  wire g1212_n;
  wire g1213_p;
  wire g1213_n;
  wire g1214_p;
  wire g1214_n;
  wire g1215_p;
  wire g1215_n;
  wire g1216_p;
  wire g1216_n;
  wire g1217_p;
  wire g1217_n;
  wire g1218_p;
  wire g1218_n;
  wire g1219_p;
  wire g1219_n;
  wire g1220_p;
  wire g1220_n;
  wire g1221_p;
  wire g1221_n;
  wire g1222_p;
  wire g1222_n;
  wire g1223_p;
  wire g1223_n;
  wire g1224_p;
  wire g1224_n;
  wire g1225_p;
  wire g1225_n;
  wire g1226_p;
  wire g1226_n;
  wire g1227_p;
  wire g1227_n;
  wire g1228_p;
  wire g1228_n;
  wire g1229_p;
  wire g1229_n;
  wire g1230_p;
  wire g1230_n;
  wire g1231_p;
  wire g1231_n;
  wire g1232_p;
  wire g1232_n;
  wire g1233_p;
  wire g1233_n;
  wire g1234_p;
  wire g1234_n;
  wire g1235_p;
  wire g1235_n;
  wire g1236_p;
  wire g1236_n;
  wire g1237_p;
  wire g1237_n;
  wire g1238_p;
  wire g1238_n;
  wire g1239_p;
  wire g1239_n;
  wire g1240_p;
  wire g1240_n;
  wire g1241_p;
  wire g1241_n;
  wire g1242_p;
  wire g1242_n;
  wire g1243_p;
  wire g1243_n;
  wire g1244_p;
  wire g1244_n;
  wire g1245_p;
  wire g1245_n;
  wire g1246_p;
  wire g1246_n;
  wire g1247_p;
  wire g1247_n;
  wire g1248_p;
  wire g1248_n;
  wire g1249_p;
  wire g1249_n;
  wire g1250_p;
  wire g1250_n;
  wire g1251_p;
  wire g1251_n;
  wire g1252_p;
  wire g1252_n;
  wire g1253_p;
  wire g1253_n;
  wire g1254_p;
  wire g1254_n;
  wire g1255_p;
  wire g1255_n;
  wire g1256_p;
  wire g1256_n;
  wire g1257_p;
  wire g1257_n;
  wire g1258_p;
  wire g1258_n;
  wire g1259_p;
  wire g1259_n;
  wire g1260_p;
  wire g1260_n;
  wire g1261_p;
  wire g1261_n;
  wire g1262_p;
  wire g1262_n;
  wire g1263_p;
  wire g1263_n;
  wire g1264_p;
  wire g1264_n;
  wire g1265_p;
  wire g1265_n;
  wire g1266_p;
  wire g1266_n;
  wire g1267_p;
  wire g1267_n;
  wire g1268_p;
  wire g1268_n;
  wire g1269_p;
  wire g1269_n;
  wire g1270_p;
  wire g1270_n;
  wire g1271_p;
  wire g1271_n;
  wire g1272_p;
  wire g1272_n;
  wire g1273_p;
  wire g1273_n;
  wire g1274_p;
  wire g1274_n;
  wire g1275_p;
  wire g1275_n;
  wire g1276_p;
  wire g1276_n;
  wire g1277_p;
  wire g1277_n;
  wire g1278_p;
  wire g1278_n;
  wire g1279_p;
  wire g1279_n;
  wire g1280_p;
  wire g1280_n;
  wire g1281_p;
  wire g1281_n;
  wire g1282_p;
  wire g1282_n;
  wire g1283_p;
  wire g1283_n;
  wire g1284_p;
  wire g1284_n;
  wire g1285_p;
  wire g1285_n;
  wire g1286_p;
  wire g1286_n;
  wire g1287_p;
  wire g1287_n;
  wire g1288_p;
  wire g1288_n;
  wire g1289_p;
  wire g1289_n;
  wire g1290_p;
  wire g1290_n;
  wire g1291_p;
  wire g1291_n;
  wire g1292_p;
  wire g1292_n;
  wire g1293_p;
  wire g1293_n;
  wire g1294_p;
  wire g1294_n;
  wire g1295_p;
  wire g1295_n;
  wire g1296_p;
  wire g1296_n;
  wire g1297_p;
  wire g1297_n;
  wire g1298_p;
  wire g1298_n;
  wire g1299_p;
  wire g1299_n;
  wire g1300_p;
  wire g1300_n;
  wire g1301_p;
  wire g1301_n;
  wire g1302_p;
  wire g1302_n;
  wire g1303_p;
  wire g1303_n;
  wire g1304_p;
  wire g1304_n;
  wire g1305_p;
  wire g1305_n;
  wire g1306_p;
  wire g1306_n;
  wire g1307_p;
  wire g1307_n;
  wire g1308_p;
  wire g1308_n;
  wire g1309_p;
  wire g1309_n;
  wire g1310_p;
  wire g1310_n;
  wire g1311_p;
  wire g1311_n;
  wire g1312_p;
  wire g1312_n;
  wire g1313_p;
  wire g1313_n;
  wire g1314_p;
  wire g1314_n;
  wire g1315_p;
  wire g1315_n;
  wire g1316_p;
  wire g1316_n;
  wire g1317_p;
  wire g1317_n;
  wire g1318_p;
  wire g1318_n;
  wire g1319_p;
  wire g1319_n;
  wire g1320_p;
  wire g1320_n;
  wire g1321_p;
  wire g1321_n;
  wire g1322_p;
  wire g1322_n;
  wire g1323_p;
  wire g1323_n;
  wire g1324_p;
  wire g1324_n;
  wire g1325_p;
  wire g1325_n;
  wire g1326_p;
  wire g1326_n;
  wire g1327_p;
  wire g1327_n;
  wire g1328_p;
  wire g1328_n;
  wire g1329_p;
  wire g1329_n;
  wire g1330_p;
  wire g1330_n;
  wire g1331_p;
  wire g1331_n;
  wire g1332_p;
  wire g1332_n;
  wire g1333_p;
  wire g1333_n;
  wire g1334_p;
  wire g1334_n;
  wire g1335_p;
  wire g1335_n;
  wire g1336_p;
  wire g1336_n;
  wire g1337_p;
  wire g1337_n;
  wire g1338_p;
  wire g1338_n;
  wire g1339_p;
  wire g1339_n;
  wire g1340_p;
  wire g1340_n;
  wire g1341_p;
  wire g1341_n;
  wire g1342_p;
  wire g1342_n;
  wire g1343_p;
  wire g1343_n;
  wire g1344_p;
  wire g1344_n;
  wire g1345_p;
  wire g1345_n;
  wire g1346_p;
  wire g1346_n;
  wire g1347_p;
  wire g1347_n;
  wire g1348_p;
  wire g1348_n;
  wire g1349_p;
  wire g1349_n;
  wire g1350_p;
  wire g1350_n;
  wire g1351_p;
  wire g1351_n;
  wire g1352_p;
  wire g1352_n;
  wire g1353_p;
  wire g1353_n;
  wire g1354_p;
  wire g1354_n;
  wire g1355_p;
  wire g1355_n;
  wire g1356_p;
  wire g1356_n;
  wire g1357_p;
  wire g1357_n;
  wire g1358_p;
  wire g1358_n;
  wire g1359_p;
  wire g1359_n;
  wire g1360_p;
  wire g1360_n;
  wire g1361_p;
  wire g1361_n;
  wire g1362_p;
  wire g1362_n;
  wire g1363_p;
  wire g1363_n;
  wire g1364_p;
  wire g1364_n;
  wire g1365_p;
  wire g1365_n;
  wire g1366_p;
  wire g1366_n;
  wire g1367_p;
  wire g1367_n;
  wire g1368_p;
  wire g1368_n;
  wire g1369_p;
  wire g1369_n;
  wire g1370_p;
  wire g1370_n;
  wire g1371_p;
  wire g1371_n;
  wire g1372_p;
  wire g1372_n;
  wire g1373_p;
  wire g1373_n;
  wire g1374_p;
  wire g1374_n;
  wire g1375_p;
  wire g1375_n;
  wire g1376_p;
  wire g1376_n;
  wire g1377_p;
  wire g1377_n;
  wire g1378_p;
  wire g1378_n;
  wire g1379_p;
  wire g1379_n;
  wire g1380_p;
  wire g1380_n;
  wire g1381_p;
  wire g1381_n;
  wire g1382_p;
  wire g1382_n;
  wire g1383_p;
  wire g1383_n;
  wire g1384_p;
  wire g1384_n;
  wire g1385_p;
  wire g1385_n;
  wire g1386_p;
  wire g1386_n;
  wire g1387_p;
  wire g1387_n;
  wire g1388_p;
  wire g1388_n;
  wire g1389_p;
  wire g1389_n;
  wire g1390_p;
  wire g1390_n;
  wire g1391_p;
  wire g1391_n;
  wire g1392_p;
  wire g1392_n;
  wire g1393_p;
  wire g1393_n;
  wire g1394_p;
  wire g1394_n;
  wire g1395_p;
  wire g1395_n;
  wire g1396_p;
  wire g1396_n;
  wire g1397_p;
  wire g1397_n;
  wire g1398_p;
  wire g1398_n;
  wire g1399_p;
  wire g1399_n;
  wire g1400_p;
  wire g1400_n;
  wire g1401_p;
  wire g1401_n;
  wire g1402_p;
  wire g1402_n;
  wire g1403_p;
  wire g1403_n;
  wire g1404_p;
  wire g1404_n;
  wire g1405_p;
  wire g1405_n;
  wire g1406_p;
  wire g1406_n;
  wire g1407_p;
  wire g1407_n;
  wire g1408_p;
  wire g1408_n;
  wire g1409_p;
  wire g1409_n;
  wire g1410_p;
  wire g1410_n;
  wire g1411_p;
  wire g1411_n;
  wire g1412_p;
  wire g1412_n;
  wire g1413_p;
  wire g1413_n;
  wire g1414_p;
  wire g1414_n;
  wire g1415_p;
  wire g1415_n;
  wire g1416_p;
  wire g1416_n;
  wire g1417_p;
  wire g1417_n;
  wire g1418_p;
  wire g1418_n;
  wire g1419_p;
  wire g1419_n;
  wire g1420_p;
  wire g1420_n;
  wire g1421_p;
  wire g1421_n;
  wire g1422_p;
  wire g1422_n;
  wire g1423_p;
  wire g1423_n;
  wire g1424_p;
  wire g1424_n;
  wire g1425_p;
  wire g1425_n;
  wire g1426_p;
  wire g1426_n;
  wire g1427_p;
  wire g1427_n;
  wire g1428_p;
  wire g1428_n;
  wire g1429_p;
  wire g1429_n;
  wire g1430_p;
  wire g1430_n;
  wire g1431_p;
  wire g1431_n;
  wire g1432_p;
  wire g1432_n;
  wire g1433_p;
  wire g1433_n;
  wire g1434_p;
  wire g1434_n;
  wire g1435_p;
  wire g1435_n;
  wire g1436_p;
  wire g1436_n;
  wire g1437_p;
  wire g1437_n;
  wire g1438_p;
  wire g1438_n;
  wire g1439_p;
  wire g1439_n;
  wire g1440_p;
  wire g1440_n;
  wire g1441_p;
  wire g1441_n;
  wire g1442_p;
  wire g1442_n;
  wire g1443_p;
  wire g1443_n;
  wire g1444_p;
  wire g1444_n;
  wire g1445_p;
  wire g1445_n;
  wire g1446_p;
  wire g1446_n;
  wire g1447_p;
  wire g1447_n;
  wire g1448_p;
  wire g1448_n;
  wire g1449_p;
  wire g1449_n;
  wire g1450_p;
  wire g1450_n;
  wire g1451_p;
  wire g1451_n;
  wire g1452_p;
  wire g1452_n;
  wire g1453_p;
  wire g1453_n;
  wire g1454_p;
  wire g1454_n;
  wire g1455_p;
  wire g1455_n;
  wire g1456_p;
  wire g1456_n;
  wire g1457_p;
  wire g1457_n;
  wire g1458_p;
  wire g1458_n;
  wire g1459_p;
  wire g1459_n;
  wire g1460_p;
  wire g1460_n;
  wire g1461_p;
  wire g1461_n;
  wire g1462_p;
  wire g1462_n;
  wire g1463_p;
  wire g1463_n;
  wire g1464_p;
  wire g1464_n;
  wire g1465_p;
  wire g1465_n;
  wire g1466_p;
  wire g1466_n;
  wire g1467_p;
  wire g1467_n;
  wire g1468_p;
  wire g1468_n;
  wire g1469_p;
  wire g1469_n;
  wire g1470_p;
  wire g1470_n;
  wire g1471_p;
  wire g1471_n;
  wire g1472_p;
  wire g1472_n;
  wire g1473_p;
  wire g1473_n;
  wire g1474_p;
  wire g1474_n;
  wire g1475_p;
  wire g1475_n;
  wire g1476_p;
  wire g1476_n;
  wire g1477_p;
  wire g1477_n;
  wire g1478_p;
  wire g1478_n;
  wire g1479_p;
  wire g1479_n;
  wire g1480_p;
  wire g1480_n;
  wire g1481_p;
  wire g1481_n;
  wire g1482_p;
  wire g1482_n;
  wire g1483_p;
  wire g1483_n;
  wire g1484_p;
  wire g1484_n;
  wire g1485_p;
  wire g1485_n;
  wire g1486_p;
  wire g1486_n;
  wire g1487_p;
  wire g1487_n;
  wire g1488_p;
  wire g1488_n;
  wire g1489_p;
  wire g1489_n;
  wire g1490_p;
  wire g1490_n;
  wire g1491_p;
  wire g1491_n;
  wire g1492_p;
  wire g1492_n;
  wire g1493_p;
  wire g1493_n;
  wire g1494_p;
  wire g1494_n;
  wire g1495_p;
  wire g1495_n;
  wire g1496_p;
  wire g1496_n;
  wire g1497_p;
  wire g1497_n;
  wire g1498_p;
  wire g1498_n;
  wire g1499_p;
  wire g1499_n;
  wire g1500_p;
  wire g1500_n;
  wire g1501_p;
  wire g1501_n;
  wire g1502_p;
  wire g1502_n;
  wire g1503_p;
  wire g1503_n;
  wire g1504_p;
  wire g1504_n;
  wire g1505_p;
  wire g1505_n;
  wire g1506_p;
  wire g1506_n;
  wire g1507_p;
  wire g1507_n;
  wire g1508_p;
  wire g1508_n;
  wire g1509_p;
  wire g1509_n;
  wire g1510_p;
  wire g1510_n;
  wire g1511_p;
  wire g1511_n;
  wire g1512_p;
  wire g1512_n;
  wire g1513_p;
  wire g1513_n;
  wire g1514_p;
  wire g1514_n;
  wire g1515_p;
  wire g1515_n;
  wire g1516_p;
  wire g1516_n;
  wire g1517_p;
  wire g1517_n;
  wire g1518_p;
  wire g1518_n;
  wire g1519_p;
  wire g1519_n;
  wire g1520_p;
  wire g1520_n;
  wire g1521_p;
  wire g1521_n;
  wire g1522_p;
  wire g1522_n;
  wire g1523_p;
  wire g1523_n;
  wire g1524_p;
  wire g1524_n;
  wire g1525_p;
  wire g1525_n;
  wire g1526_p;
  wire g1526_n;
  wire g1527_p;
  wire g1527_n;
  wire g1528_p;
  wire g1528_n;
  wire g1529_p;
  wire g1529_n;
  wire g1530_p;
  wire g1530_n;
  wire g1531_p;
  wire g1531_n;
  wire g1532_p;
  wire g1532_n;
  wire g1533_p;
  wire g1533_n;
  wire g1534_p;
  wire g1534_n;
  wire g1535_p;
  wire g1535_n;
  wire g1536_p;
  wire g1536_n;
  wire g1537_p;
  wire g1537_n;
  wire g1538_p;
  wire g1538_n;
  wire g1539_p;
  wire g1539_n;
  wire g1540_p;
  wire g1540_n;
  wire g1541_p;
  wire g1541_n;
  wire g1542_p;
  wire g1542_n;
  wire g1543_p;
  wire g1543_n;
  wire g1544_p;
  wire g1544_n;
  wire g1545_p;
  wire g1545_n;
  wire g1546_p;
  wire g1546_n;
  wire g1547_p;
  wire g1547_n;
  wire g1548_p;
  wire g1548_n;
  wire g1549_p;
  wire g1549_n;
  wire g1550_p;
  wire g1550_n;
  wire g1551_p;
  wire g1551_n;
  wire g1552_p;
  wire g1552_n;
  wire g1553_p;
  wire g1553_n;
  wire g1554_p;
  wire g1554_n;
  wire g1555_p;
  wire g1555_n;
  wire g1556_p;
  wire g1556_n;
  wire g1557_p;
  wire g1557_n;
  wire g1558_p;
  wire g1558_n;
  wire g1559_p;
  wire g1559_n;
  wire g1560_p;
  wire g1560_n;
  wire g1561_p;
  wire g1561_n;
  wire g1562_p;
  wire g1562_n;
  wire g1563_p;
  wire g1563_n;
  wire g1564_p;
  wire g1564_n;
  wire g1565_p;
  wire g1565_n;
  wire g1566_p;
  wire g1566_n;
  wire g1567_p;
  wire g1567_n;
  wire g1568_p;
  wire g1568_n;
  wire g1569_p;
  wire g1569_n;
  wire g1570_p;
  wire g1570_n;
  wire g1571_p;
  wire g1571_n;
  wire g1572_p;
  wire g1572_n;
  wire g1573_p;
  wire g1573_n;
  wire g1574_p;
  wire g1574_n;
  wire g1575_p;
  wire g1575_n;
  wire g1576_p;
  wire g1576_n;
  wire g1577_p;
  wire g1577_n;
  wire g1578_p;
  wire g1578_n;
  wire g1579_p;
  wire g1579_n;
  wire g1580_p;
  wire g1580_n;
  wire g1581_p;
  wire g1581_n;
  wire g1582_p;
  wire g1582_n;
  wire g1583_p;
  wire g1583_n;
  wire g1584_p;
  wire g1584_n;
  wire g1585_p;
  wire g1585_n;
  wire g1586_p;
  wire g1586_n;
  wire g1587_p;
  wire g1587_n;
  wire g1588_p;
  wire g1588_n;
  wire g1589_p;
  wire g1589_n;
  wire g1590_p;
  wire g1590_n;
  wire g1591_p;
  wire g1591_n;
  wire g1592_p;
  wire g1592_n;
  wire g1593_p;
  wire g1593_n;
  wire g1594_p;
  wire g1594_n;
  wire g1595_p;
  wire g1595_n;
  wire g1596_p;
  wire g1596_n;
  wire g1597_p;
  wire g1597_n;
  wire g1598_p;
  wire g1598_n;
  wire g1599_p;
  wire g1599_n;
  wire g1600_p;
  wire g1600_n;
  wire g1601_p;
  wire g1601_n;
  wire g1602_p;
  wire g1602_n;
  wire g1603_p;
  wire g1603_n;
  wire g1604_p;
  wire g1604_n;
  wire g1605_p;
  wire g1605_n;
  wire g1606_p;
  wire g1606_n;
  wire g1607_p;
  wire g1607_n;
  wire g1608_p;
  wire g1608_n;
  wire g1609_p;
  wire g1609_n;
  wire g1610_p;
  wire g1610_n;
  wire g1611_p;
  wire g1611_n;
  wire g1612_p;
  wire g1612_n;
  wire g1613_p;
  wire g1613_n;
  wire g1614_p;
  wire g1614_n;
  wire g1615_p;
  wire g1615_n;
  wire g1616_p;
  wire g1616_n;
  wire g1617_p;
  wire g1617_n;
  wire g1618_p;
  wire g1618_n;
  wire g1619_p;
  wire g1619_n;
  wire g1620_p;
  wire g1620_n;
  wire g1621_p;
  wire g1621_n;
  wire g1622_p;
  wire g1622_n;
  wire g1623_p;
  wire g1623_n;
  wire g1624_p;
  wire g1624_n;
  wire g1625_p;
  wire g1625_n;
  wire g1626_p;
  wire g1626_n;
  wire g1627_p;
  wire g1627_n;
  wire g1628_p;
  wire g1628_n;
  wire g1629_p;
  wire g1629_n;
  wire g1630_p;
  wire g1630_n;
  wire g1631_p;
  wire g1631_n;
  wire g1632_p;
  wire g1632_n;
  wire g1633_p;
  wire g1633_n;
  wire g1634_p;
  wire g1634_n;
  wire g1635_p;
  wire g1635_n;
  wire g1636_p;
  wire g1636_n;
  wire g1637_p;
  wire g1637_n;
  wire g1638_p;
  wire g1638_n;
  wire g1639_p;
  wire g1639_n;
  wire g1640_p;
  wire g1640_n;
  wire g1641_p;
  wire g1641_n;
  wire g1642_p;
  wire g1642_n;
  wire g1643_p;
  wire g1643_n;
  wire g1644_p;
  wire g1644_n;
  wire g1645_p;
  wire g1645_n;
  wire g1646_p;
  wire g1646_n;
  wire g1647_p;
  wire g1647_n;
  wire g1648_p;
  wire g1648_n;
  wire g1649_p;
  wire g1649_n;
  wire g1650_p;
  wire g1650_n;
  wire g1651_p;
  wire g1651_n;
  wire g1652_p;
  wire g1652_n;
  wire g1653_p;
  wire g1653_n;
  wire g1654_p;
  wire g1654_n;
  wire g1655_p;
  wire g1655_n;
  wire g1656_p;
  wire g1656_n;
  wire g1657_p;
  wire g1657_n;
  wire g1658_p;
  wire g1658_n;
  wire g1659_p;
  wire g1659_n;
  wire g1660_p;
  wire g1660_n;
  wire g1661_p;
  wire g1661_n;
  wire g1662_p;
  wire g1662_n;
  wire g1663_p;
  wire g1663_n;
  wire g1664_p;
  wire g1664_n;
  wire g1665_p;
  wire g1665_n;
  wire g1666_p;
  wire g1666_n;
  wire g1667_p;
  wire g1667_n;
  wire g1668_p;
  wire g1668_n;
  wire g1669_p;
  wire g1669_n;
  wire g1670_p;
  wire g1670_n;
  wire g1671_p;
  wire g1671_n;
  wire g1672_p;
  wire g1672_n;
  wire g1673_p;
  wire g1673_n;
  wire g1674_p;
  wire g1674_n;
  wire g1675_p;
  wire g1675_n;
  wire g1676_p;
  wire g1676_n;
  wire g1677_p;
  wire g1677_n;
  wire g1678_p;
  wire g1678_n;
  wire g1679_p;
  wire g1679_n;
  wire g1680_p;
  wire g1680_n;
  wire g1681_p;
  wire g1681_n;
  wire g1682_p;
  wire g1682_n;
  wire g1683_p;
  wire g1683_n;
  wire g1684_p;
  wire g1684_n;
  wire g1685_p;
  wire g1685_n;
  wire g1686_p;
  wire g1686_n;
  wire g1687_p;
  wire g1687_n;
  wire g1688_p;
  wire g1688_n;
  wire g1689_p;
  wire g1689_n;
  wire g1690_p;
  wire g1690_n;
  wire g1691_p;
  wire g1691_n;
  wire g1692_p;
  wire g1692_n;
  wire g1693_p;
  wire g1693_n;
  wire g1694_p;
  wire g1694_n;
  wire g1695_p;
  wire g1695_n;
  wire g1696_p;
  wire g1696_n;
  wire g1697_p;
  wire g1697_n;
  wire g1698_p;
  wire g1698_n;
  wire g1699_p;
  wire g1699_n;
  wire g1700_p;
  wire g1700_n;
  wire g1701_p;
  wire g1701_n;
  wire g1702_p;
  wire g1702_n;
  wire g1703_p;
  wire g1703_n;
  wire g1704_p;
  wire g1704_n;
  wire g1705_p;
  wire g1705_n;
  wire g1706_p;
  wire g1706_n;
  wire g1707_p;
  wire g1707_n;
  wire g1708_p;
  wire g1708_n;
  wire g1709_p;
  wire g1709_n;
  wire g1710_p;
  wire g1710_n;
  wire g1711_p;
  wire g1711_n;
  wire g1712_p;
  wire g1712_n;
  wire g1713_p;
  wire g1713_n;
  wire g1714_p;
  wire g1714_n;
  wire g1715_p;
  wire g1715_n;
  wire g1716_p;
  wire g1716_n;
  wire g1717_p;
  wire g1717_n;
  wire g1718_p;
  wire g1718_n;
  wire g1719_p;
  wire g1719_n;
  wire g1720_p;
  wire g1720_n;
  wire g1721_p;
  wire g1721_n;
  wire g1722_p;
  wire g1722_n;
  wire g1723_p;
  wire g1723_n;
  wire g1724_p;
  wire g1724_n;
  wire g1725_p;
  wire g1725_n;
  wire g1726_p;
  wire g1726_n;
  wire n5011_o2_n_spl_;
  wire n5011_o2_p_spl_;
  wire n5013_o2_n_spl_;
  wire n5013_o2_p_spl_;
  wire g585_n_spl_;
  wire n2172_lo_n_spl_;
  wire n2160_lo_n_spl_;
  wire n2148_lo_n_spl_;
  wire g589_p_spl_;
  wire g589_n_spl_;
  wire g585_p_spl_;
  wire n4634_o2_n_spl_;
  wire n4633_o2_p_spl_;
  wire n4634_o2_p_spl_;
  wire n4633_o2_n_spl_;
  wire n4418_o2_p_spl_;
  wire n2304_lo_p_spl_;
  wire g633_n_spl_;
  wire g636_n_spl_;
  wire G2991_o2_n_spl_;
  wire G2887_o2_p_spl_;
  wire G2991_o2_p_spl_;
  wire G2887_o2_n_spl_;
  wire n4733_o2_p_spl_;
  wire n4732_o2_p_spl_;
  wire n4733_o2_n_spl_;
  wire n4732_o2_n_spl_;
  wire g666_n_spl_;
  wire g669_n_spl_;
  wire g672_n_spl_;
  wire g675_n_spl_;
  wire g681_n_spl_;
  wire g683_n_spl_;
  wire g688_n_spl_;
  wire g687_n_spl_;
  wire g694_n_spl_;
  wire g693_p_spl_;
  wire g694_p_spl_;
  wire g693_n_spl_;
  wire G3360_o2_p_spl_;
  wire G3350_o2_n_spl_;
  wire G3360_o2_n_spl_;
  wire G3350_o2_p_spl_;
  wire g703_n_spl_;
  wire g700_n_spl_;
  wire g700_n_spl_0;
  wire g700_n_spl_1;
  wire g703_p_spl_;
  wire g700_p_spl_;
  wire g700_p_spl_0;
  wire g700_p_spl_1;
  wire g704_p_spl_;
  wire g704_p_spl_0;
  wire g704_p_spl_1;
  wire g704_n_spl_;
  wire g704_n_spl_0;
  wire g704_n_spl_1;
  wire G3399_o2_p_spl_;
  wire G3383_o2_n_spl_;
  wire G3399_o2_n_spl_;
  wire G3383_o2_p_spl_;
  wire g709_p_spl_;
  wire g709_n_spl_;
  wire G3240_o2_p_spl_;
  wire G3376_o2_p_spl_;
  wire G3240_o2_n_spl_;
  wire G3376_o2_n_spl_;
  wire g714_p_spl_;
  wire g714_n_spl_;
  wire g697_n_spl_;
  wire g697_p_spl_;
  wire G3367_o2_n_spl_;
  wire G3353_o2_p_spl_;
  wire G3367_o2_p_spl_;
  wire G3353_o2_n_spl_;
  wire g727_n_spl_;
  wire g727_p_spl_;
  wire G434_o2_p_spl_;
  wire n852_inv_n_spl_;
  wire n852_inv_n_spl_0;
  wire n849_inv_n_spl_;
  wire n852_inv_p_spl_;
  wire n852_inv_p_spl_0;
  wire n852_inv_p_spl_1;
  wire n849_inv_p_spl_;
  wire n849_inv_p_spl_0;
  wire n855_inv_p_spl_;
  wire n4539_o2_p_spl_;
  wire n4539_o2_p_spl_0;
  wire n4539_o2_n_spl_;
  wire n4539_o2_n_spl_0;
  wire n4816_o2_n_spl_;
  wire n429_inv_n_spl_;
  wire n4816_o2_p_spl_;
  wire n429_inv_p_spl_;
  wire n429_inv_p_spl_0;
  wire n4398_o2_p_spl_;
  wire g752_n_spl_;
  wire g752_n_spl_0;
  wire g749_n_spl_;
  wire g756_p_spl_;
  wire g756_p_spl_0;
  wire g752_p_spl_;
  wire g752_p_spl_0;
  wire g752_p_spl_00;
  wire g752_p_spl_01;
  wire g752_p_spl_1;
  wire g752_p_spl_10;
  wire G3069_o2_n_spl_;
  wire G2962_o2_n_spl_;
  wire G3069_o2_p_spl_;
  wire G2962_o2_p_spl_;
  wire g760_p_spl_;
  wire g760_p_spl_0;
  wire g764_p_spl_;
  wire n1941_lo_buf_o2_n_spl_;
  wire n1941_lo_buf_o2_n_spl_0;
  wire n1056_inv_p_spl_;
  wire n1056_inv_p_spl_0;
  wire n1056_inv_p_spl_00;
  wire n1056_inv_p_spl_01;
  wire n1056_inv_p_spl_1;
  wire n858_inv_p_spl_;
  wire n858_inv_p_spl_0;
  wire n858_inv_p_spl_00;
  wire n858_inv_p_spl_01;
  wire n858_inv_p_spl_1;
  wire n4651_o2_n_spl_;
  wire n4651_o2_n_spl_0;
  wire n4651_o2_n_spl_00;
  wire n4651_o2_n_spl_01;
  wire n4651_o2_n_spl_1;
  wire n4919_o2_n_spl_;
  wire n4919_o2_n_spl_0;
  wire n4919_o2_n_spl_00;
  wire n4919_o2_n_spl_01;
  wire n4919_o2_n_spl_1;
  wire n1977_lo_buf_o2_n_spl_;
  wire n1977_lo_buf_o2_n_spl_0;
  wire n1977_lo_buf_o2_n_spl_00;
  wire n1977_lo_buf_o2_n_spl_1;
  wire n1965_lo_buf_o2_n_spl_;
  wire n1965_lo_buf_o2_n_spl_0;
  wire n1965_lo_buf_o2_n_spl_00;
  wire n1965_lo_buf_o2_n_spl_1;
  wire n1953_lo_buf_o2_n_spl_;
  wire n1953_lo_buf_o2_n_spl_0;
  wire n1953_lo_buf_o2_n_spl_1;
  wire G519_o2_n_spl_;
  wire G519_o2_n_spl_0;
  wire G519_o2_n_spl_00;
  wire G519_o2_n_spl_000;
  wire G519_o2_n_spl_01;
  wire G519_o2_n_spl_1;
  wire G519_o2_n_spl_10;
  wire G519_o2_n_spl_11;
  wire n4653_o2_n_spl_;
  wire n4653_o2_n_spl_0;
  wire n4653_o2_n_spl_1;
  wire n1071_inv_p_spl_;
  wire n1071_inv_p_spl_0;
  wire n1071_inv_p_spl_00;
  wire n1071_inv_p_spl_01;
  wire n1071_inv_p_spl_1;
  wire n1068_inv_p_spl_;
  wire n1068_inv_p_spl_0;
  wire n1068_inv_p_spl_00;
  wire n1068_inv_p_spl_01;
  wire n1068_inv_p_spl_1;
  wire n1062_inv_p_spl_;
  wire n1062_inv_p_spl_0;
  wire n1062_inv_p_spl_00;
  wire n1062_inv_p_spl_01;
  wire n1062_inv_p_spl_1;
  wire n1062_inv_p_spl_10;
  wire n1053_inv_p_spl_;
  wire n1053_inv_p_spl_0;
  wire n1053_inv_p_spl_00;
  wire n1053_inv_p_spl_01;
  wire n1053_inv_p_spl_1;
  wire n1074_inv_p_spl_;
  wire n1074_inv_p_spl_0;
  wire n1074_inv_p_spl_00;
  wire n1074_inv_p_spl_01;
  wire n1074_inv_p_spl_1;
  wire n1074_inv_p_spl_10;
  wire n4571_o2_n_spl_;
  wire n4571_o2_n_spl_0;
  wire n4571_o2_n_spl_00;
  wire n4571_o2_n_spl_01;
  wire n4571_o2_n_spl_1;
  wire n4572_o2_n_spl_;
  wire n4572_o2_n_spl_0;
  wire n4572_o2_n_spl_00;
  wire n4572_o2_n_spl_1;
  wire G519_o2_p_spl_;
  wire G519_o2_p_spl_0;
  wire G519_o2_p_spl_00;
  wire G519_o2_p_spl_000;
  wire G519_o2_p_spl_01;
  wire G519_o2_p_spl_1;
  wire G519_o2_p_spl_10;
  wire G519_o2_p_spl_11;
  wire g801_n_spl_;
  wire g801_n_spl_0;
  wire g801_n_spl_00;
  wire g801_n_spl_01;
  wire g801_n_spl_1;
  wire g801_n_spl_10;
  wire n4389_o2_p_spl_;
  wire n4389_o2_p_spl_0;
  wire n4389_o2_p_spl_1;
  wire n4389_o2_n_spl_;
  wire n4389_o2_n_spl_0;
  wire n4389_o2_n_spl_1;
  wire g806_p_spl_;
  wire g806_p_spl_0;
  wire g806_p_spl_1;
  wire g801_p_spl_;
  wire g801_p_spl_0;
  wire g801_p_spl_1;
  wire g808_p_spl_;
  wire g808_p_spl_0;
  wire g808_p_spl_1;
  wire g743_p_spl_;
  wire g743_p_spl_0;
  wire g743_p_spl_00;
  wire g743_p_spl_01;
  wire g743_p_spl_1;
  wire g743_p_spl_10;
  wire g743_p_spl_11;
  wire g743_n_spl_;
  wire g743_n_spl_0;
  wire g812_n_spl_;
  wire g812_n_spl_0;
  wire g812_n_spl_00;
  wire g812_n_spl_01;
  wire g812_n_spl_1;
  wire G2923_o2_p_spl_;
  wire G2923_o2_p_spl_0;
  wire g749_p_spl_;
  wire G2923_o2_n_spl_;
  wire G2923_o2_n_spl_0;
  wire n2301_lo_buf_o2_p_spl_;
  wire n2301_lo_buf_o2_p_spl_0;
  wire n2301_lo_buf_o2_n_spl_;
  wire g825_n_spl_;
  wire n1050_inv_p_spl_;
  wire n1050_inv_p_spl_0;
  wire n1050_inv_p_spl_00;
  wire n1050_inv_p_spl_01;
  wire n1050_inv_p_spl_1;
  wire n2253_lo_buf_o2_n_spl_;
  wire n2241_lo_buf_o2_n_spl_;
  wire n2241_lo_buf_o2_n_spl_0;
  wire g871_p_spl_;
  wire g871_p_spl_0;
  wire G772_o2_n_spl_;
  wire G772_o2_p_spl_;
  wire g873_p_spl_;
  wire g873_p_spl_0;
  wire g737_n_spl_;
  wire g875_n_spl_;
  wire g875_n_spl_0;
  wire g873_n_spl_;
  wire g873_n_spl_0;
  wire g875_p_spl_;
  wire g875_p_spl_0;
  wire g876_p_spl_;
  wire g871_n_spl_;
  wire g871_n_spl_0;
  wire g880_p_spl_;
  wire n1068_inv_n_spl_;
  wire n1071_inv_n_spl_;
  wire n1050_inv_n_spl_;
  wire n1056_inv_n_spl_;
  wire n858_inv_n_spl_;
  wire n4651_o2_p_spl_;
  wire n2265_lo_buf_o2_p_spl_;
  wire n1053_inv_n_spl_;
  wire n4571_o2_p_spl_;
  wire n4572_o2_p_spl_;
  wire n4653_o2_p_spl_;
  wire n2241_lo_buf_o2_p_spl_;
  wire n2253_lo_buf_o2_p_spl_;
  wire g740_p_spl_;
  wire g876_n_spl_;
  wire g880_n_spl_;
  wire g812_p_spl_;
  wire G461_o2_p_spl_;
  wire G935_o2_p_spl_;
  wire g734_n_spl_;
  wire n4454_o2_p_spl_;
  wire G3039_o2_n_spl_;
  wire G3039_o2_n_spl_0;
  wire G3039_o2_p_spl_;
  wire G3039_o2_p_spl_0;
  wire n2061_lo_buf_o2_p_spl_;
  wire g1043_p_spl_;
  wire n2313_lo_buf_o2_p_spl_;
  wire g1043_n_spl_;
  wire g1044_n_spl_;
  wire g1044_n_spl_0;
  wire g1044_n_spl_00;
  wire g1044_n_spl_01;
  wire g1044_n_spl_1;
  wire g1044_n_spl_10;
  wire g1044_n_spl_11;
  wire g746_n_spl_;
  wire g1044_p_spl_;
  wire g1044_p_spl_0;
  wire g1044_p_spl_00;
  wire g1044_p_spl_01;
  wire g1044_p_spl_1;
  wire g1044_p_spl_10;
  wire g1044_p_spl_11;
  wire G2507_o2_p_spl_;
  wire G2507_o2_p_spl_0;
  wire G2507_o2_p_spl_1;
  wire G2444_o2_p_spl_;
  wire G2444_o2_p_spl_0;
  wire G2444_o2_p_spl_1;
  wire G2507_o2_n_spl_;
  wire G2507_o2_n_spl_0;
  wire G2444_o2_n_spl_;
  wire G2444_o2_n_spl_0;
  wire g1049_p_spl_;
  wire g1049_p_spl_0;
  wire g1049_p_spl_1;
  wire g1049_n_spl_;
  wire g1049_n_spl_0;
  wire G3024_o2_n_spl_;
  wire G2902_o2_p_spl_;
  wire G3024_o2_p_spl_;
  wire G2902_o2_n_spl_;
  wire g1058_p_spl_;
  wire g1058_p_spl_0;
  wire G1689_o2_p_spl_;
  wire G1689_o2_p_spl_0;
  wire n2013_lo_buf_o2_p_spl_;
  wire G1689_o2_n_spl_;
  wire G1689_o2_n_spl_0;
  wire G1955_o2_n_spl_;
  wire G1955_o2_p_spl_;
  wire n2025_lo_buf_o2_p_spl_;
  wire n2025_lo_buf_o2_n_spl_;
  wire G1958_o2_n_spl_;
  wire G1958_o2_p_spl_;
  wire G1693_o2_n_spl_;
  wire G1693_o2_n_spl_0;
  wire n2037_lo_buf_o2_p_spl_;
  wire G1693_o2_p_spl_;
  wire G1693_o2_p_spl_0;
  wire n2037_lo_buf_o2_n_spl_;
  wire n2049_lo_buf_o2_p_spl_;
  wire n2049_lo_buf_o2_n_spl_;
  wire n2049_lo_buf_o2_n_spl_0;
  wire g1064_n_spl_;
  wire g1071_p_spl_;
  wire g1071_p_spl_0;
  wire g1071_p_spl_00;
  wire g1071_p_spl_01;
  wire g1071_p_spl_1;
  wire G2502_o2_p_spl_;
  wire g1071_n_spl_;
  wire g1071_n_spl_0;
  wire g1077_p_spl_;
  wire g1077_p_spl_0;
  wire g832_p_spl_;
  wire g753_p_spl_;
  wire g930_p_spl_;
  wire g1042_n_spl_;
  wire g757_n_spl_;
  wire g981_n_spl_;
  wire g1037_n_spl_;
  wire g761_n_spl_;
  wire g813_n_spl_;
  wire g822_n_spl_;
  wire g765_n_spl_;
  wire g884_n_spl_;
  wire G2759_o2_n_spl_;
  wire G2666_o2_p_spl_;
  wire G2759_o2_p_spl_;
  wire G2666_o2_n_spl_;
  wire g1094_p_spl_;
  wire G1529_o2_p_spl_;
  wire G1529_o2_p_spl_0;
  wire G1538_o2_p_spl_;
  wire G1538_o2_p_spl_0;
  wire G1547_o2_n_spl_;
  wire G1547_o2_n_spl_0;
  wire G1556_o2_p_spl_;
  wire G1556_o2_p_spl_0;
  wire G1565_o2_p_spl_;
  wire G1565_o2_p_spl_0;
  wire G1574_o2_p_spl_;
  wire G1574_o2_p_spl_0;
  wire G1583_o2_n_spl_;
  wire G1583_o2_n_spl_0;
  wire G1592_o2_p_spl_;
  wire G1592_o2_p_spl_0;
  wire n1929_lo_n_spl_;
  wire G1601_o2_p_spl_;
  wire G1601_o2_p_spl_0;
  wire G1610_o2_p_spl_;
  wire G1610_o2_p_spl_0;
  wire G1619_o2_n_spl_;
  wire G1619_o2_n_spl_0;
  wire G1628_o2_p_spl_;
  wire G1628_o2_p_spl_0;
  wire G1637_o2_p_spl_;
  wire G1637_o2_p_spl_0;
  wire G1646_o2_p_spl_;
  wire G1646_o2_p_spl_0;
  wire G1655_o2_n_spl_;
  wire G1655_o2_n_spl_0;
  wire G1664_o2_p_spl_;
  wire G1664_o2_p_spl_0;
  wire n861_inv_n_spl_;
  wire g827_p_spl_;
  wire g826_p_spl_;
  wire g1032_p_spl_;
  wire G1738_o2_p_spl_;
  wire G1733_o2_p_spl_;
  wire G1738_o2_n_spl_;
  wire G1733_o2_n_spl_;
  wire G1751_o2_p_spl_;
  wire G1751_o2_n_spl_;
  wire G1764_o2_p_spl_;
  wire G1764_o2_n_spl_;
  wire G615_o2_p_spl_;
  wire G615_o2_n_spl_;
  wire g1052_p_spl_;
  wire g1237_n_spl_;
  wire g1059_n_spl_;
  wire g1184_n_spl_;
  wire g1232_n_spl_;
  wire g1078_n_spl_;
  wire g1142_n_spl_;
  wire g1238_n_spl_;
  wire g1095_n_spl_;
  wire g1226_n_spl_;
  wire g1259_n_spl_;
  wire g1261_n_spl_;
  wire g1263_n_spl_;
  wire n1554_inv_n_spl_;
  wire G2027_o2_n_spl_;
  wire n1554_inv_p_spl_;
  wire n1554_inv_p_spl_0;
  wire G2027_o2_p_spl_;
  wire G2027_o2_p_spl_0;
  wire g1274_n_spl_;
  wire g1273_n_spl_;
  wire g1274_p_spl_;
  wire g1274_p_spl_0;
  wire g1273_p_spl_;
  wire g1273_p_spl_0;
  wire g1273_p_spl_1;
  wire g1270_n_spl_;
  wire g1275_p_spl_;
  wire g1270_p_spl_;
  wire n2097_lo_buf_o2_p_spl_;
  wire n2097_lo_buf_o2_p_spl_0;
  wire n5326_o2_n_spl_;
  wire n2097_lo_buf_o2_n_spl_;
  wire n5326_o2_p_spl_;
  wire n5326_o2_p_spl_0;
  wire n2133_lo_buf_o2_n_spl_;
  wire n5327_o2_p_spl_;
  wire n5327_o2_p_spl_0;
  wire n2133_lo_buf_o2_p_spl_;
  wire n2133_lo_buf_o2_p_spl_0;
  wire n5327_o2_n_spl_;
  wire g1074_n_spl_;
  wire g1074_n_spl_0;
  wire g1045_n_spl_;
  wire g1045_n_spl_0;
  wire g1045_n_spl_00;
  wire g1045_n_spl_01;
  wire g1045_n_spl_1;
  wire g1269_n_spl_;
  wire n1557_inv_n_spl_;
  wire G2393_o2_n_spl_;
  wire n1557_inv_p_spl_;
  wire n1557_inv_p_spl_0;
  wire G2393_o2_p_spl_;
  wire G2393_o2_p_spl_0;
  wire g1289_p_spl_;
  wire g1288_p_spl_;
  wire g1288_p_spl_0;
  wire g1289_n_spl_;
  wire g1288_n_spl_;
  wire g1288_n_spl_0;
  wire g1288_n_spl_1;
  wire G2577_o2_n_spl_;
  wire G2281_o2_n_spl_;
  wire G2577_o2_p_spl_;
  wire G2281_o2_p_spl_;
  wire g1293_p_spl_;
  wire g1293_p_spl_0;
  wire g1293_p_spl_1;
  wire g1293_n_spl_;
  wire g1293_n_spl_0;
  wire g1293_n_spl_00;
  wire g1293_n_spl_01;
  wire g1293_n_spl_1;
  wire g1295_p_spl_;
  wire g1294_n_spl_;
  wire g1294_n_spl_0;
  wire g1295_n_spl_;
  wire g1294_p_spl_;
  wire g1294_p_spl_0;
  wire g1055_p_spl_;
  wire g1055_p_spl_0;
  wire g1055_p_spl_1;
  wire g1055_n_spl_;
  wire g1055_n_spl_0;
  wire g1055_n_spl_00;
  wire g1055_n_spl_1;
  wire g1045_p_spl_;
  wire g1045_p_spl_0;
  wire g1045_p_spl_00;
  wire g1045_p_spl_1;
  wire n4921_o2_p_spl_;
  wire n4920_o2_p_spl_;
  wire n4920_o2_p_spl_0;
  wire g1302_p_spl_;
  wire g1254_p_spl_;
  wire g1254_p_spl_0;
  wire g1256_p_spl_;
  wire g1256_p_spl_0;
  wire G1189_o2_p_spl_;
  wire G1189_o2_n_spl_;
  wire g1305_n_spl_;
  wire g1305_p_spl_;
  wire g1305_p_spl_0;
  wire n1761_lo_buf_o2_p_spl_;
  wire n1761_lo_buf_o2_p_spl_0;
  wire n1761_lo_buf_o2_p_spl_1;
  wire n1749_lo_buf_o2_p_spl_;
  wire n1749_lo_buf_o2_p_spl_0;
  wire n1749_lo_buf_o2_p_spl_00;
  wire n1749_lo_buf_o2_p_spl_01;
  wire n1749_lo_buf_o2_p_spl_1;
  wire n1749_lo_buf_o2_p_spl_10;
  wire n1749_lo_buf_o2_p_spl_11;
  wire n1749_lo_buf_o2_n_spl_;
  wire n1749_lo_buf_o2_n_spl_0;
  wire n1749_lo_buf_o2_n_spl_00;
  wire n1749_lo_buf_o2_n_spl_01;
  wire n1749_lo_buf_o2_n_spl_1;
  wire g1309_p_spl_;
  wire g1309_p_spl_0;
  wire g1309_n_spl_;
  wire g1309_n_spl_0;
  wire n1809_lo_buf_o2_n_spl_;
  wire n1809_lo_buf_o2_p_spl_;
  wire n1809_lo_buf_o2_p_spl_0;
  wire g1310_n_spl_;
  wire g1310_n_spl_0;
  wire g1310_n_spl_00;
  wire g1310_n_spl_000;
  wire g1310_n_spl_01;
  wire g1310_n_spl_1;
  wire g1310_n_spl_10;
  wire g1310_n_spl_11;
  wire n2139_lo_buf_o2_p_spl_;
  wire n2139_lo_buf_o2_p_spl_0;
  wire n2139_lo_buf_o2_p_spl_1;
  wire g1310_p_spl_;
  wire g1310_p_spl_0;
  wire g1310_p_spl_00;
  wire g1310_p_spl_01;
  wire g1310_p_spl_1;
  wire g1310_p_spl_10;
  wire n2139_lo_buf_o2_n_spl_;
  wire n2139_lo_buf_o2_n_spl_0;
  wire g1311_n_spl_;
  wire g1311_p_spl_;
  wire n2187_lo_buf_o2_p_spl_;
  wire n2187_lo_buf_o2_n_spl_;
  wire g1314_p_spl_;
  wire g1314_n_spl_;
  wire n1899_lo_buf_o2_p_spl_;
  wire n1899_lo_buf_o2_p_spl_0;
  wire n1899_lo_buf_o2_p_spl_00;
  wire n1899_lo_buf_o2_p_spl_01;
  wire n1899_lo_buf_o2_p_spl_1;
  wire G831_o2_n_spl_;
  wire G831_o2_n_spl_0;
  wire G831_o2_n_spl_00;
  wire G831_o2_n_spl_01;
  wire G831_o2_n_spl_1;
  wire G831_o2_n_spl_10;
  wire G831_o2_n_spl_11;
  wire n1899_lo_buf_o2_n_spl_;
  wire n1899_lo_buf_o2_n_spl_0;
  wire n1899_lo_buf_o2_n_spl_00;
  wire n1899_lo_buf_o2_n_spl_1;
  wire G831_o2_p_spl_;
  wire G831_o2_p_spl_0;
  wire G831_o2_p_spl_00;
  wire G831_o2_p_spl_01;
  wire G831_o2_p_spl_1;
  wire n2121_lo_buf_o2_p_spl_;
  wire n2121_lo_buf_o2_p_spl_0;
  wire n2121_lo_buf_o2_p_spl_1;
  wire G594_o2_n_spl_;
  wire G594_o2_n_spl_0;
  wire G594_o2_n_spl_00;
  wire G594_o2_n_spl_01;
  wire G594_o2_n_spl_1;
  wire G594_o2_n_spl_10;
  wire G594_o2_n_spl_11;
  wire n2121_lo_buf_o2_n_spl_;
  wire n2121_lo_buf_o2_n_spl_0;
  wire G594_o2_p_spl_;
  wire G594_o2_p_spl_0;
  wire G594_o2_p_spl_00;
  wire G594_o2_p_spl_01;
  wire G594_o2_p_spl_1;
  wire g1318_p_spl_;
  wire g1318_p_spl_0;
  wire g1318_p_spl_00;
  wire g1318_p_spl_01;
  wire g1318_p_spl_1;
  wire g1318_p_spl_10;
  wire n2127_lo_buf_o2_p_spl_;
  wire n2127_lo_buf_o2_p_spl_0;
  wire n2127_lo_buf_o2_p_spl_1;
  wire g1318_n_spl_;
  wire g1318_n_spl_0;
  wire g1318_n_spl_00;
  wire g1318_n_spl_1;
  wire n2127_lo_buf_o2_n_spl_;
  wire n2127_lo_buf_o2_n_spl_0;
  wire G477_o2_n_spl_;
  wire G477_o2_p_spl_;
  wire n1797_lo_buf_o2_p_spl_;
  wire n2151_lo_buf_o2_p_spl_;
  wire n2151_lo_buf_o2_p_spl_0;
  wire n2151_lo_buf_o2_p_spl_1;
  wire n2151_lo_buf_o2_n_spl_;
  wire g1326_n_spl_;
  wire g1326_n_spl_0;
  wire g1326_n_spl_1;
  wire g1326_p_spl_;
  wire g1326_p_spl_0;
  wire n2199_lo_buf_o2_p_spl_;
  wire n2199_lo_buf_o2_p_spl_0;
  wire n2199_lo_buf_o2_n_spl_;
  wire g1329_n_spl_;
  wire g1329_p_spl_;
  wire g1329_p_spl_0;
  wire n2163_lo_p_spl_;
  wire n2163_lo_p_spl_0;
  wire n2211_lo_buf_o2_p_spl_;
  wire G501_o2_p_spl_;
  wire G501_o2_p_spl_0;
  wire G501_o2_p_spl_00;
  wire G501_o2_p_spl_000;
  wire G501_o2_p_spl_01;
  wire G501_o2_p_spl_1;
  wire G501_o2_p_spl_10;
  wire G501_o2_p_spl_11;
  wire n1854_lo_buf_o2_p_spl_;
  wire n1854_lo_buf_o2_p_spl_0;
  wire n1854_lo_buf_o2_p_spl_00;
  wire n1854_lo_buf_o2_p_spl_01;
  wire n1854_lo_buf_o2_p_spl_1;
  wire n1854_lo_buf_o2_p_spl_10;
  wire G501_o2_n_spl_;
  wire G501_o2_n_spl_0;
  wire G501_o2_n_spl_00;
  wire G501_o2_n_spl_01;
  wire G501_o2_n_spl_1;
  wire G501_o2_n_spl_10;
  wire G501_o2_n_spl_11;
  wire n1854_lo_buf_o2_n_spl_;
  wire n1854_lo_buf_o2_n_spl_0;
  wire n1854_lo_buf_o2_n_spl_00;
  wire n1854_lo_buf_o2_n_spl_1;
  wire n1869_lo_buf_o2_n_spl_;
  wire n1869_lo_buf_o2_n_spl_0;
  wire n1869_lo_buf_o2_n_spl_00;
  wire n1869_lo_buf_o2_n_spl_01;
  wire n1869_lo_buf_o2_n_spl_1;
  wire G667_o2_p_spl_;
  wire G667_o2_p_spl_0;
  wire G667_o2_p_spl_00;
  wire G667_o2_p_spl_000;
  wire G667_o2_p_spl_01;
  wire G667_o2_p_spl_1;
  wire G667_o2_p_spl_10;
  wire G667_o2_p_spl_11;
  wire n1869_lo_buf_o2_p_spl_;
  wire n1869_lo_buf_o2_p_spl_0;
  wire n1869_lo_buf_o2_p_spl_00;
  wire n1869_lo_buf_o2_p_spl_01;
  wire n1869_lo_buf_o2_p_spl_1;
  wire n1869_lo_buf_o2_p_spl_10;
  wire n1869_lo_buf_o2_p_spl_11;
  wire G667_o2_n_spl_;
  wire G667_o2_n_spl_0;
  wire G667_o2_n_spl_00;
  wire G667_o2_n_spl_01;
  wire G667_o2_n_spl_1;
  wire G667_o2_n_spl_10;
  wire G667_o2_n_spl_11;
  wire g1350_p_spl_;
  wire g1350_p_spl_0;
  wire g1350_p_spl_00;
  wire g1350_p_spl_01;
  wire g1350_p_spl_1;
  wire g1350_p_spl_10;
  wire g1350_p_spl_11;
  wire n1833_lo_buf_o2_n_spl_;
  wire n1833_lo_buf_o2_n_spl_0;
  wire n1833_lo_buf_o2_n_spl_1;
  wire g1350_n_spl_;
  wire g1350_n_spl_0;
  wire g1350_n_spl_00;
  wire g1350_n_spl_01;
  wire g1350_n_spl_1;
  wire g1350_n_spl_10;
  wire n1833_lo_buf_o2_p_spl_;
  wire n1833_lo_buf_o2_p_spl_0;
  wire n1833_lo_buf_o2_p_spl_00;
  wire n1833_lo_buf_o2_p_spl_01;
  wire n1833_lo_buf_o2_p_spl_1;
  wire n1773_lo_buf_o2_p_spl_;
  wire n1773_lo_buf_o2_p_spl_0;
  wire n1773_lo_buf_o2_p_spl_00;
  wire n1773_lo_buf_o2_p_spl_1;
  wire n1773_lo_buf_o2_n_spl_;
  wire n1785_lo_buf_o2_p_spl_;
  wire n1785_lo_buf_o2_p_spl_0;
  wire n1785_lo_buf_o2_n_spl_;
  wire g1356_n_spl_;
  wire g1356_n_spl_0;
  wire g1356_n_spl_00;
  wire g1356_n_spl_000;
  wire g1356_n_spl_01;
  wire g1356_n_spl_1;
  wire g1356_n_spl_10;
  wire g1356_n_spl_11;
  wire g1356_p_spl_;
  wire g1356_p_spl_0;
  wire g1356_p_spl_00;
  wire g1356_p_spl_01;
  wire g1356_p_spl_1;
  wire g1356_p_spl_10;
  wire g1356_p_spl_11;
  wire g1358_p_spl_;
  wire g1358_p_spl_0;
  wire g1358_p_spl_00;
  wire g1358_p_spl_000;
  wire g1358_p_spl_01;
  wire g1358_p_spl_1;
  wire g1358_p_spl_10;
  wire g1358_p_spl_11;
  wire g1358_n_spl_;
  wire g1358_n_spl_0;
  wire g1358_n_spl_00;
  wire g1358_n_spl_01;
  wire g1358_n_spl_1;
  wire g1358_n_spl_10;
  wire g1358_n_spl_11;
  wire g1360_n_spl_;
  wire g1360_n_spl_0;
  wire g1360_n_spl_1;
  wire g1360_p_spl_;
  wire g1360_p_spl_0;
  wire g1361_p_spl_;
  wire g1361_p_spl_0;
  wire g1361_p_spl_00;
  wire g1361_p_spl_01;
  wire g1361_p_spl_1;
  wire g1361_p_spl_10;
  wire g1361_p_spl_11;
  wire g1361_n_spl_;
  wire g1361_n_spl_0;
  wire g1361_n_spl_00;
  wire g1361_n_spl_01;
  wire g1361_n_spl_1;
  wire g1361_n_spl_10;
  wire g1366_n_spl_;
  wire g1366_n_spl_0;
  wire g1366_n_spl_00;
  wire g1366_n_spl_000;
  wire g1366_n_spl_01;
  wire g1366_n_spl_1;
  wire g1366_n_spl_10;
  wire g1366_n_spl_11;
  wire g1366_p_spl_;
  wire g1366_p_spl_0;
  wire g1366_p_spl_00;
  wire g1366_p_spl_01;
  wire g1366_p_spl_1;
  wire g1366_p_spl_10;
  wire g1367_n_spl_;
  wire g1367_n_spl_0;
  wire g1367_n_spl_00;
  wire g1367_n_spl_1;
  wire g1367_p_spl_;
  wire g1367_p_spl_0;
  wire g1367_p_spl_1;
  wire n1893_lo_buf_o2_p_spl_;
  wire n1893_lo_buf_o2_p_spl_0;
  wire n1893_lo_buf_o2_p_spl_00;
  wire n1893_lo_buf_o2_p_spl_01;
  wire n1893_lo_buf_o2_p_spl_1;
  wire n1893_lo_buf_o2_p_spl_10;
  wire n1893_lo_buf_o2_p_spl_11;
  wire n1893_lo_buf_o2_n_spl_;
  wire n1893_lo_buf_o2_n_spl_0;
  wire n1893_lo_buf_o2_n_spl_00;
  wire n1893_lo_buf_o2_n_spl_01;
  wire n1893_lo_buf_o2_n_spl_1;
  wire n2109_lo_buf_o2_p_spl_;
  wire n2109_lo_buf_o2_p_spl_0;
  wire n2109_lo_buf_o2_p_spl_1;
  wire n2109_lo_buf_o2_n_spl_;
  wire n2109_lo_buf_o2_n_spl_0;
  wire g1371_n_spl_;
  wire g1371_n_spl_0;
  wire g1371_p_spl_;
  wire g1371_p_spl_0;
  wire g1371_p_spl_1;
  wire g1365_p_spl_;
  wire g1365_p_spl_0;
  wire g1365_p_spl_00;
  wire g1365_p_spl_1;
  wire n2007_lo_n_spl_;
  wire n2007_lo_n_spl_0;
  wire n2007_lo_n_spl_00;
  wire n2007_lo_n_spl_01;
  wire n2007_lo_n_spl_1;
  wire g1379_n_spl_;
  wire n2019_lo_n_spl_;
  wire n2019_lo_n_spl_0;
  wire n2019_lo_n_spl_00;
  wire n2019_lo_n_spl_01;
  wire n2019_lo_n_spl_1;
  wire g1252_p_spl_;
  wire g1252_p_spl_0;
  wire n1845_lo_buf_o2_n_spl_;
  wire n1845_lo_buf_o2_n_spl_0;
  wire n1845_lo_buf_o2_n_spl_00;
  wire n1845_lo_buf_o2_n_spl_1;
  wire n1845_lo_buf_o2_p_spl_;
  wire n1845_lo_buf_o2_p_spl_0;
  wire n1845_lo_buf_o2_p_spl_00;
  wire n1845_lo_buf_o2_p_spl_01;
  wire n1845_lo_buf_o2_p_spl_1;
  wire n1845_lo_buf_o2_p_spl_10;
  wire n1845_lo_buf_o2_p_spl_11;
  wire n1815_lo_buf_o2_p_spl_;
  wire n1815_lo_buf_o2_p_spl_0;
  wire n1815_lo_buf_o2_p_spl_00;
  wire n1815_lo_buf_o2_p_spl_1;
  wire n1815_lo_buf_o2_n_spl_;
  wire n1881_lo_buf_o2_p_spl_;
  wire n1881_lo_buf_o2_p_spl_0;
  wire n1881_lo_buf_o2_p_spl_00;
  wire n1881_lo_buf_o2_p_spl_01;
  wire n1881_lo_buf_o2_p_spl_1;
  wire n1881_lo_buf_o2_p_spl_10;
  wire n1881_lo_buf_o2_p_spl_11;
  wire n1881_lo_buf_o2_n_spl_;
  wire n1881_lo_buf_o2_n_spl_0;
  wire n1881_lo_buf_o2_n_spl_00;
  wire n1881_lo_buf_o2_n_spl_01;
  wire n1881_lo_buf_o2_n_spl_1;
  wire n2094_lo_buf_o2_p_spl_;
  wire n2094_lo_buf_o2_p_spl_0;
  wire n2094_lo_buf_o2_p_spl_1;
  wire n2094_lo_buf_o2_n_spl_;
  wire g1400_p_spl_;
  wire g1400_p_spl_0;
  wire g1400_p_spl_00;
  wire g1400_p_spl_1;
  wire g1410_n_spl_;
  wire g1425_n_spl_;
  wire g1425_n_spl_0;
  wire g1425_n_spl_1;
  wire g1425_p_spl_;
  wire g1425_p_spl_0;
  wire g1425_p_spl_1;
  wire n2175_lo_p_spl_;
  wire n2223_lo_p_spl_;
  wire n1995_lo_p_spl_;
  wire n2079_lo_buf_o2_p_spl_;
  wire g1466_p_spl_;
  wire g1466_p_spl_0;
  wire g1466_p_spl_00;
  wire g1466_p_spl_1;
  wire g1476_n_spl_;
  wire g1389_n_spl_;
  wire g1481_n_spl_;
  wire g1481_n_spl_0;
  wire g1383_n_spl_;
  wire g1381_n_spl_;
  wire n2031_lo_p_spl_;
  wire n2031_lo_p_spl_0;
  wire n2031_lo_p_spl_1;
  wire g1379_p_spl_;
  wire n2043_lo_p_spl_;
  wire n2043_lo_p_spl_0;
  wire n2043_lo_p_spl_1;
  wire g1252_n_spl_;
  wire n2298_lo_n_spl_;
  wire n2298_lo_n_spl_0;
  wire n2298_lo_n_spl_00;
  wire n2298_lo_n_spl_01;
  wire n2298_lo_n_spl_1;
  wire n2298_lo_n_spl_10;
  wire g1385_n_spl_;
  wire n1905_lo_buf_o2_p_spl_;
  wire n1905_lo_buf_o2_p_spl_0;
  wire n1905_lo_buf_o2_p_spl_1;
  wire g1087_p_spl_;
  wire g1087_p_spl_0;
  wire g1081_n_spl_;
  wire g1081_n_spl_0;
  wire g1240_n_spl_;
  wire g1240_n_spl_0;
  wire g1083_p_spl_;
  wire g1083_p_spl_0;
  wire g1512_n_spl_;
  wire g1512_p_spl_;
  wire g1512_p_spl_0;
  wire g1515_p_spl_;
  wire g1515_p_spl_0;
  wire g1515_p_spl_1;
  wire g1386_n_spl_;
  wire g1386_n_spl_0;
  wire g1493_p_spl_;
  wire g1452_n_spl_;
  wire g1452_n_spl_0;
  wire g1452_n_spl_00;
  wire g1452_n_spl_1;
  wire g1482_n_spl_;
  wire g1482_n_spl_0;
  wire g1482_n_spl_00;
  wire g1482_n_spl_1;
  wire g1308_p_spl_;
  wire n2145_lo_buf_o2_p_spl_;
  wire n2157_lo_buf_o2_p_spl_;
  wire n2169_lo_buf_o2_p_spl_;
  wire n2181_lo_buf_o2_p_spl_;
  wire g1515_n_spl_;
  wire g1515_n_spl_0;
  wire g1276_p_spl_;
  wire n5101_o2_p_spl_;
  wire n5101_o2_p_spl_0;
  wire n5267_o2_p_spl_;
  wire n5267_o2_p_spl_0;
  wire n5267_o2_p_spl_1;
  wire n5325_o2_p_spl_;
  wire n5325_o2_p_spl_0;
  wire n5325_o2_p_spl_1;
  wire g1542_n_spl_;
  wire g1542_p_spl_;
  wire g1542_p_spl_0;
  wire n5294_o2_p_spl_;
  wire n5294_o2_p_spl_0;
  wire n5294_o2_p_spl_00;
  wire n5294_o2_p_spl_1;
  wire n5294_o2_n_spl_;
  wire n5294_o2_n_spl_0;
  wire g1556_p_spl_;
  wire g1556_p_spl_0;
  wire g1557_n_spl_;
  wire g1555_n_spl_;
  wire g1555_n_spl_0;
  wire g1555_n_spl_1;
  wire g1555_p_spl_;
  wire g1555_p_spl_0;
  wire g1555_p_spl_1;
  wire g1560_n_spl_;
  wire g1561_p_spl_;
  wire g1563_n_spl_;
  wire g1565_n_spl_;
  wire g1414_n_spl_;
  wire g1412_n_spl_;
  wire g1410_p_spl_;
  wire n1857_lo_buf_o2_n_spl_;
  wire n1857_lo_buf_o2_n_spl_0;
  wire n5100_o2_n_spl_;
  wire n5100_o2_n_spl_0;
  wire g1507_n_spl_;
  wire n1821_lo_buf_o2_p_spl_;
  wire n1821_lo_buf_o2_p_spl_0;
  wire n1821_lo_buf_o2_p_spl_00;
  wire n1821_lo_buf_o2_p_spl_1;
  wire n5266_o2_n_spl_;
  wire n5266_o2_n_spl_0;
  wire g1582_n_spl_;
  wire g1504_n_spl_;
  wire g1526_n_spl_;
  wire g1526_n_spl_0;
  wire g1526_n_spl_1;
  wire g1524_n_spl_;
  wire g1524_n_spl_0;
  wire g1524_n_spl_1;
  wire g1591_n_spl_;
  wire g1591_n_spl_0;
  wire g1586_n_spl_;
  wire g1586_n_spl_0;
  wire g1607_n_spl_;
  wire g1607_n_spl_0;
  wire g1607_n_spl_1;
  wire n2007_lo_p_spl_;
  wire n2007_lo_p_spl_0;
  wire n2007_lo_p_spl_1;
  wire g1607_p_spl_;
  wire g1607_p_spl_0;
  wire g1607_p_spl_1;
  wire g1347_p_spl_;
  wire g1347_n_spl_;
  wire g1347_n_spl_0;
  wire g1347_n_spl_00;
  wire g1347_n_spl_1;
  wire n2019_lo_p_spl_;
  wire n2019_lo_p_spl_0;
  wire n2019_lo_p_spl_00;
  wire n2019_lo_p_spl_1;
  wire g1429_n_spl_;
  wire g1429_n_spl_0;
  wire g1429_n_spl_00;
  wire g1429_n_spl_1;
  wire g1429_p_spl_;
  wire g1429_p_spl_0;
  wire g1337_p_spl_;
  wire g1337_n_spl_;
  wire g1337_n_spl_0;
  wire g1337_n_spl_00;
  wire g1337_n_spl_1;
  wire n5293_o2_p_spl_;
  wire n5292_o2_p_spl_;
  wire n5292_o2_p_spl_0;
  wire n5266_o2_p_spl_;
  wire n5266_o2_p_spl_0;
  wire n5266_o2_p_spl_00;
  wire n5266_o2_p_spl_01;
  wire n5266_o2_p_spl_1;
  wire n5100_o2_p_spl_;
  wire n5100_o2_p_spl_0;
  wire n5100_o2_p_spl_00;
  wire n5100_o2_p_spl_01;
  wire n5100_o2_p_spl_1;
  wire n1821_lo_buf_o2_n_spl_;
  wire n1821_lo_buf_o2_n_spl_0;
  wire g1506_n_spl_;
  wire g1387_p_spl_;
  wire n2298_lo_p_spl_;
  wire g1284_n_spl_;
  wire g1522_n_spl_;
  wire g1520_n_spl_;
  wire n1857_lo_buf_o2_p_spl_;
  wire n1857_lo_buf_o2_p_spl_0;
  wire n1857_lo_buf_o2_p_spl_00;
  wire n1857_lo_buf_o2_p_spl_1;
  wire g1079_n_spl_;
  wire g1079_p_spl_;
  wire g1079_p_spl_0;
  wire g1301_n_spl_;
  wire g1279_n_spl_;
  wire g1282_n_spl_;
  wire g1442_n_spl_;
  wire g1442_n_spl_0;
  wire g1442_n_spl_00;
  wire g1442_n_spl_1;
  wire g1324_p_spl_;
  wire n2031_lo_n_spl_;
  wire n2031_lo_n_spl_0;
  wire n2031_lo_n_spl_1;
  wire g1324_n_spl_;
  wire g1324_n_spl_0;
  wire n2043_lo_n_spl_;
  wire n2043_lo_n_spl_0;
  wire n2043_lo_n_spl_1;
  wire g1656_n_spl_;
  wire g1612_n_spl_;
  wire g1480_n_spl_;
  wire g1478_n_spl_;
  wire g1476_p_spl_;
  wire g1617_n_spl_;
  wire g1493_n_spl_;
  wire g1493_n_spl_0;
  wire g1493_n_spl_1;
  wire G5_p_spl_;
  wire G5_p_spl_0;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_00;
  wire G4_p_spl_01;
  wire G4_p_spl_1;
  wire G4_p_spl_10;
  wire G4_p_spl_11;
  wire n1983_lo_p_spl_;
  wire g1685_n_spl_;
  wire g1685_n_spl_0;
  wire g1663_n_spl_;
  wire g1663_n_spl_0;
  wire g1663_n_spl_1;
  wire g1625_p_spl_;
  wire g1670_n_spl_;
  wire g1670_n_spl_0;
  wire G6_p_spl_;
  wire g1693_n_spl_;
  wire g1693_n_spl_0;
  wire G3_p_spl_;
  wire G3_p_spl_0;
  wire G2_p_spl_;
  wire n5295_o2_p_spl_;
  wire n5295_o2_p_spl_0;
  wire n5295_o2_p_spl_00;
  wire n5295_o2_p_spl_1;
  wire g1085_p_spl_;
  wire g1085_p_spl_0;
  wire g1085_p_spl_1;
  wire g1258_p_spl_;
  wire g1258_p_spl_0;
  wire g1258_p_spl_1;
  wire g1303_n_spl_;
  wire g1304_n_spl_;
  wire g1501_p_spl_;
  wire g1501_p_spl_0;
  wire g1501_p_spl_1;
  wire g1517_n_spl_;
  wire g1518_n_spl_;
  wire g1523_n_spl_;
  wire g1523_n_spl_0;
  wire g1529_n_spl_;
  wire g1532_n_spl_;
  wire g1535_n_spl_;
  wire g1538_n_spl_;
  wire g1541_n_spl_;
  wire g1554_n_spl_;
  wire g1558_n_spl_;
  wire g1558_n_spl_0;
  wire g1558_n_spl_00;
  wire g1558_n_spl_000;
  wire g1558_n_spl_001;
  wire g1558_n_spl_01;
  wire g1558_n_spl_010;
  wire g1558_n_spl_011;
  wire g1558_n_spl_1;
  wire g1558_n_spl_10;
  wire g1558_n_spl_11;
  wire g1559_n_spl_;
  wire g1559_n_spl_0;
  wire g1559_n_spl_00;
  wire g1559_n_spl_000;
  wire g1559_n_spl_001;
  wire g1559_n_spl_01;
  wire g1559_n_spl_010;
  wire g1559_n_spl_011;
  wire g1559_n_spl_1;
  wire g1559_n_spl_10;
  wire g1559_n_spl_11;
  wire g1562_p_spl_;
  wire g1562_p_spl_0;
  wire g1562_p_spl_00;
  wire g1562_p_spl_000;
  wire g1562_p_spl_001;
  wire g1562_p_spl_01;
  wire g1562_p_spl_010;
  wire g1562_p_spl_011;
  wire g1562_p_spl_1;
  wire g1562_p_spl_10;
  wire g1562_p_spl_11;
  wire g1564_n_spl_;
  wire g1564_n_spl_0;
  wire g1564_n_spl_00;
  wire g1564_n_spl_000;
  wire g1564_n_spl_001;
  wire g1564_n_spl_01;
  wire g1564_n_spl_010;
  wire g1564_n_spl_011;
  wire g1564_n_spl_1;
  wire g1564_n_spl_10;
  wire g1564_n_spl_11;
  wire g1566_n_spl_;
  wire g1566_n_spl_0;
  wire g1566_n_spl_00;
  wire g1566_n_spl_000;
  wire g1566_n_spl_001;
  wire g1566_n_spl_01;
  wire g1566_n_spl_010;
  wire g1566_n_spl_011;
  wire g1566_n_spl_1;
  wire g1566_n_spl_10;
  wire g1566_n_spl_11;
  wire g1567_p_spl_;
  wire g1567_p_spl_0;
  wire g1567_p_spl_00;
  wire g1567_p_spl_000;
  wire g1567_p_spl_001;
  wire g1567_p_spl_01;
  wire g1567_p_spl_010;
  wire g1567_p_spl_011;
  wire g1567_p_spl_1;
  wire g1567_p_spl_10;
  wire g1567_p_spl_11;
  wire g1568_n_spl_;
  wire g1568_n_spl_0;
  wire g1568_n_spl_00;
  wire g1568_n_spl_000;
  wire g1568_n_spl_001;
  wire g1568_n_spl_01;
  wire g1568_n_spl_010;
  wire g1568_n_spl_011;
  wire g1568_n_spl_1;
  wire g1568_n_spl_10;
  wire g1568_n_spl_11;
  wire g1569_n_spl_;
  wire g1569_n_spl_0;
  wire g1569_n_spl_00;
  wire g1569_n_spl_000;
  wire g1569_n_spl_001;
  wire g1569_n_spl_01;
  wire g1569_n_spl_010;
  wire g1569_n_spl_011;
  wire g1569_n_spl_1;
  wire g1569_n_spl_10;
  wire g1569_n_spl_11;
  wire g1577_p_spl_;
  wire g1577_p_spl_0;
  wire G9_p_spl_;
  wire G9_p_spl_0;
  wire G9_p_spl_1;
  wire G13_p_spl_;
  wire G13_p_spl_0;
  wire G13_p_spl_1;
  wire g1592_n_spl_;
  wire g1678_p_spl_;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire g1692_p_spl_;
  wire g1706_n_spl_;
  wire G1_p_spl_;
  wire g1719_n_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  buf

  (
    G42_p,
    G42
  );


  not

  (
    G42_n,
    G42
  );


  buf

  (
    G43_p,
    G43
  );


  not

  (
    G43_n,
    G43
  );


  buf

  (
    G44_p,
    G44
  );


  not

  (
    G44_n,
    G44
  );


  buf

  (
    G45_p,
    G45
  );


  not

  (
    G45_n,
    G45
  );


  buf

  (
    G46_p,
    G46
  );


  not

  (
    G46_n,
    G46
  );


  buf

  (
    G47_p,
    G47
  );


  not

  (
    G47_n,
    G47
  );


  buf

  (
    G48_p,
    G48
  );


  not

  (
    G48_n,
    G48
  );


  buf

  (
    G49_p,
    G49
  );


  not

  (
    G49_n,
    G49
  );


  buf

  (
    G50_p,
    G50
  );


  not

  (
    G50_n,
    G50
  );


  buf

  (
    n1836_lo_p,
    n1836_lo
  );


  not

  (
    n1836_lo_n,
    n1836_lo
  );


  buf

  (
    n1872_lo_p,
    n1872_lo
  );


  not

  (
    n1872_lo_n,
    n1872_lo
  );


  buf

  (
    n1884_lo_p,
    n1884_lo
  );


  not

  (
    n1884_lo_n,
    n1884_lo
  );


  buf

  (
    n1911_lo_p,
    n1911_lo
  );


  not

  (
    n1911_lo_n,
    n1911_lo
  );


  buf

  (
    n1914_lo_p,
    n1914_lo
  );


  not

  (
    n1914_lo_n,
    n1914_lo
  );


  buf

  (
    n1917_lo_p,
    n1917_lo
  );


  not

  (
    n1917_lo_n,
    n1917_lo
  );


  buf

  (
    n1923_lo_p,
    n1923_lo
  );


  not

  (
    n1923_lo_n,
    n1923_lo
  );


  buf

  (
    n1926_lo_p,
    n1926_lo
  );


  not

  (
    n1926_lo_n,
    n1926_lo
  );


  buf

  (
    n1929_lo_p,
    n1929_lo
  );


  not

  (
    n1929_lo_n,
    n1929_lo
  );


  buf

  (
    n1935_lo_p,
    n1935_lo
  );


  not

  (
    n1935_lo_n,
    n1935_lo
  );


  buf

  (
    n1938_lo_p,
    n1938_lo
  );


  not

  (
    n1938_lo_n,
    n1938_lo
  );


  buf

  (
    n1947_lo_p,
    n1947_lo
  );


  not

  (
    n1947_lo_n,
    n1947_lo
  );


  buf

  (
    n1950_lo_p,
    n1950_lo
  );


  not

  (
    n1950_lo_n,
    n1950_lo
  );


  buf

  (
    n1959_lo_p,
    n1959_lo
  );


  not

  (
    n1959_lo_n,
    n1959_lo
  );


  buf

  (
    n1962_lo_p,
    n1962_lo
  );


  not

  (
    n1962_lo_n,
    n1962_lo
  );


  buf

  (
    n1971_lo_p,
    n1971_lo
  );


  not

  (
    n1971_lo_n,
    n1971_lo
  );


  buf

  (
    n1974_lo_p,
    n1974_lo
  );


  not

  (
    n1974_lo_n,
    n1974_lo
  );


  buf

  (
    n1983_lo_p,
    n1983_lo
  );


  not

  (
    n1983_lo_n,
    n1983_lo
  );


  buf

  (
    n1995_lo_p,
    n1995_lo
  );


  not

  (
    n1995_lo_n,
    n1995_lo
  );


  buf

  (
    n2007_lo_p,
    n2007_lo
  );


  not

  (
    n2007_lo_n,
    n2007_lo
  );


  buf

  (
    n2019_lo_p,
    n2019_lo
  );


  not

  (
    n2019_lo_n,
    n2019_lo
  );


  buf

  (
    n2031_lo_p,
    n2031_lo
  );


  not

  (
    n2031_lo_n,
    n2031_lo
  );


  buf

  (
    n2043_lo_p,
    n2043_lo
  );


  not

  (
    n2043_lo_n,
    n2043_lo
  );


  buf

  (
    n2055_lo_p,
    n2055_lo
  );


  not

  (
    n2055_lo_n,
    n2055_lo
  );


  buf

  (
    n2064_lo_p,
    n2064_lo
  );


  not

  (
    n2064_lo_n,
    n2064_lo
  );


  buf

  (
    n2067_lo_p,
    n2067_lo
  );


  not

  (
    n2067_lo_n,
    n2067_lo
  );


  buf

  (
    n2100_lo_p,
    n2100_lo
  );


  not

  (
    n2100_lo_n,
    n2100_lo
  );


  buf

  (
    n2112_lo_p,
    n2112_lo
  );


  not

  (
    n2112_lo_n,
    n2112_lo
  );


  buf

  (
    n2124_lo_p,
    n2124_lo
  );


  not

  (
    n2124_lo_n,
    n2124_lo
  );


  buf

  (
    n2136_lo_p,
    n2136_lo
  );


  not

  (
    n2136_lo_n,
    n2136_lo
  );


  buf

  (
    n2148_lo_p,
    n2148_lo
  );


  not

  (
    n2148_lo_n,
    n2148_lo
  );


  buf

  (
    n2160_lo_p,
    n2160_lo
  );


  not

  (
    n2160_lo_n,
    n2160_lo
  );


  buf

  (
    n2163_lo_p,
    n2163_lo
  );


  not

  (
    n2163_lo_n,
    n2163_lo
  );


  buf

  (
    n2172_lo_p,
    n2172_lo
  );


  not

  (
    n2172_lo_n,
    n2172_lo
  );


  buf

  (
    n2175_lo_p,
    n2175_lo
  );


  not

  (
    n2175_lo_n,
    n2175_lo
  );


  buf

  (
    n2184_lo_p,
    n2184_lo
  );


  not

  (
    n2184_lo_n,
    n2184_lo
  );


  buf

  (
    n2223_lo_p,
    n2223_lo
  );


  not

  (
    n2223_lo_n,
    n2223_lo
  );


  buf

  (
    n2235_lo_p,
    n2235_lo
  );


  not

  (
    n2235_lo_n,
    n2235_lo
  );


  buf

  (
    n2238_lo_p,
    n2238_lo
  );


  not

  (
    n2238_lo_n,
    n2238_lo
  );


  buf

  (
    n2247_lo_p,
    n2247_lo
  );


  not

  (
    n2247_lo_n,
    n2247_lo
  );


  buf

  (
    n2250_lo_p,
    n2250_lo
  );


  not

  (
    n2250_lo_n,
    n2250_lo
  );


  buf

  (
    n2259_lo_p,
    n2259_lo
  );


  not

  (
    n2259_lo_n,
    n2259_lo
  );


  buf

  (
    n2262_lo_p,
    n2262_lo
  );


  not

  (
    n2262_lo_n,
    n2262_lo
  );


  buf

  (
    n2271_lo_p,
    n2271_lo
  );


  not

  (
    n2271_lo_n,
    n2271_lo
  );


  buf

  (
    n2274_lo_p,
    n2274_lo
  );


  not

  (
    n2274_lo_n,
    n2274_lo
  );


  buf

  (
    n2283_lo_p,
    n2283_lo
  );


  not

  (
    n2283_lo_n,
    n2283_lo
  );


  buf

  (
    n2286_lo_p,
    n2286_lo
  );


  not

  (
    n2286_lo_n,
    n2286_lo
  );


  buf

  (
    n2295_lo_p,
    n2295_lo
  );


  not

  (
    n2295_lo_n,
    n2295_lo
  );


  buf

  (
    n2298_lo_p,
    n2298_lo
  );


  not

  (
    n2298_lo_n,
    n2298_lo
  );


  buf

  (
    n2304_lo_p,
    n2304_lo
  );


  not

  (
    n2304_lo_n,
    n2304_lo
  );


  buf

  (
    n2307_lo_p,
    n2307_lo
  );


  not

  (
    n2307_lo_n,
    n2307_lo
  );


  buf

  (
    n2331_lo_p,
    n2331_lo
  );


  not

  (
    n2331_lo_n,
    n2331_lo
  );


  buf

  (
    n2334_lo_p,
    n2334_lo
  );


  not

  (
    n2334_lo_n,
    n2334_lo
  );


  buf

  (
    n2337_lo_p,
    n2337_lo
  );


  not

  (
    n2337_lo_n,
    n2337_lo
  );


  buf

  (
    n2340_lo_p,
    n2340_lo
  );


  not

  (
    n2340_lo_n,
    n2340_lo
  );


  buf

  (
    n3241_o2_p,
    n3241_o2
  );


  not

  (
    n3241_o2_n,
    n3241_o2
  );


  buf

  (
    n3242_o2_p,
    n3242_o2
  );


  not

  (
    n3242_o2_n,
    n3242_o2
  );


  buf

  (
    n3610_o2_p,
    n3610_o2
  );


  not

  (
    n3610_o2_n,
    n3610_o2
  );


  buf

  (
    n3980_o2_p,
    n3980_o2
  );


  not

  (
    n3980_o2_n,
    n3980_o2
  );


  buf

  (
    n3968_o2_p,
    n3968_o2
  );


  not

  (
    n3968_o2_n,
    n3968_o2
  );


  buf

  (
    n4298_o2_p,
    n4298_o2
  );


  not

  (
    n4298_o2_n,
    n4298_o2
  );


  buf

  (
    n4371_o2_p,
    n4371_o2
  );


  not

  (
    n4371_o2_n,
    n4371_o2
  );


  buf

  (
    n4413_o2_p,
    n4413_o2
  );


  not

  (
    n4413_o2_n,
    n4413_o2
  );


  buf

  (
    n4418_o2_p,
    n4418_o2
  );


  not

  (
    n4418_o2_n,
    n4418_o2
  );


  buf

  (
    n4628_o2_p,
    n4628_o2
  );


  not

  (
    n4628_o2_n,
    n4628_o2
  );


  buf

  (
    n4629_o2_p,
    n4629_o2
  );


  not

  (
    n4629_o2_n,
    n4629_o2
  );


  buf

  (
    n4633_o2_p,
    n4633_o2
  );


  not

  (
    n4633_o2_n,
    n4633_o2
  );


  buf

  (
    n4634_o2_p,
    n4634_o2
  );


  not

  (
    n4634_o2_n,
    n4634_o2
  );


  buf

  (
    n4732_o2_p,
    n4732_o2
  );


  not

  (
    n4732_o2_n,
    n4732_o2
  );


  buf

  (
    n4733_o2_p,
    n4733_o2
  );


  not

  (
    n4733_o2_n,
    n4733_o2
  );


  buf

  (
    n4884_o2_p,
    n4884_o2
  );


  not

  (
    n4884_o2_n,
    n4884_o2
  );


  buf

  (
    n4886_o2_p,
    n4886_o2
  );


  not

  (
    n4886_o2_n,
    n4886_o2
  );


  buf

  (
    n4890_o2_p,
    n4890_o2
  );


  not

  (
    n4890_o2_n,
    n4890_o2
  );


  buf

  (
    n5011_o2_p,
    n5011_o2
  );


  not

  (
    n5011_o2_n,
    n5011_o2
  );


  buf

  (
    n5012_o2_p,
    n5012_o2
  );


  not

  (
    n5012_o2_n,
    n5012_o2
  );


  buf

  (
    n5013_o2_p,
    n5013_o2
  );


  not

  (
    n5013_o2_n,
    n5013_o2
  );


  buf

  (
    n5014_o2_p,
    n5014_o2
  );


  not

  (
    n5014_o2_n,
    n5014_o2
  );


  buf

  (
    n5015_o2_p,
    n5015_o2
  );


  not

  (
    n5015_o2_n,
    n5015_o2
  );


  buf

  (
    n5021_o2_p,
    n5021_o2
  );


  not

  (
    n5021_o2_n,
    n5021_o2
  );


  buf

  (
    n5016_o2_p,
    n5016_o2
  );


  not

  (
    n5016_o2_n,
    n5016_o2
  );


  buf

  (
    n5026_o2_p,
    n5026_o2
  );


  not

  (
    n5026_o2_n,
    n5026_o2
  );


  buf

  (
    n4377_o2_p,
    n4377_o2
  );


  not

  (
    n4377_o2_n,
    n4377_o2
  );


  buf

  (
    n4378_o2_p,
    n4378_o2
  );


  not

  (
    n4378_o2_n,
    n4378_o2
  );


  buf

  (
    n4389_o2_p,
    n4389_o2
  );


  not

  (
    n4389_o2_n,
    n4389_o2
  );


  buf

  (
    n327_inv_p,
    n327_inv
  );


  not

  (
    n327_inv_n,
    n327_inv
  );


  buf

  (
    n330_inv_p,
    n330_inv
  );


  not

  (
    n330_inv_n,
    n330_inv
  );


  buf

  (
    n4398_o2_p,
    n4398_o2
  );


  not

  (
    n4398_o2_n,
    n4398_o2
  );


  buf

  (
    n4401_o2_p,
    n4401_o2
  );


  not

  (
    n4401_o2_n,
    n4401_o2
  );


  buf

  (
    n5117_o2_p,
    n5117_o2
  );


  not

  (
    n5117_o2_n,
    n5117_o2
  );


  buf

  (
    n5115_o2_p,
    n5115_o2
  );


  not

  (
    n5115_o2_n,
    n5115_o2
  );


  buf

  (
    n5122_o2_p,
    n5122_o2
  );


  not

  (
    n5122_o2_n,
    n5122_o2
  );


  buf

  (
    n5121_o2_p,
    n5121_o2
  );


  not

  (
    n5121_o2_n,
    n5121_o2
  );


  buf

  (
    n5119_o2_p,
    n5119_o2
  );


  not

  (
    n5119_o2_n,
    n5119_o2
  );


  buf

  (
    n5116_o2_p,
    n5116_o2
  );


  not

  (
    n5116_o2_n,
    n5116_o2
  );


  buf

  (
    n5123_o2_p,
    n5123_o2
  );


  not

  (
    n5123_o2_n,
    n5123_o2
  );


  buf

  (
    n5156_o2_p,
    n5156_o2
  );


  not

  (
    n5156_o2_n,
    n5156_o2
  );


  buf

  (
    n5167_o2_p,
    n5167_o2
  );


  not

  (
    n5167_o2_n,
    n5167_o2
  );


  buf

  (
    n4454_o2_p,
    n4454_o2
  );


  not

  (
    n4454_o2_n,
    n4454_o2
  );


  buf

  (
    n4455_o2_p,
    n4455_o2
  );


  not

  (
    n4455_o2_n,
    n4455_o2
  );


  buf

  (
    n4456_o2_p,
    n4456_o2
  );


  not

  (
    n4456_o2_n,
    n4456_o2
  );


  buf

  (
    n4505_o2_p,
    n4505_o2
  );


  not

  (
    n4505_o2_n,
    n4505_o2
  );


  buf

  (
    G742_o2_p,
    G742_o2
  );


  not

  (
    G742_o2_n,
    G742_o2
  );


  buf

  (
    G727_o2_p,
    G727_o2
  );


  not

  (
    G727_o2_n,
    G727_o2
  );


  buf

  (
    n4567_o2_p,
    n4567_o2
  );


  not

  (
    n4567_o2_n,
    n4567_o2
  );


  buf

  (
    n4568_o2_p,
    n4568_o2
  );


  not

  (
    n4568_o2_n,
    n4568_o2
  );


  buf

  (
    n4569_o2_p,
    n4569_o2
  );


  not

  (
    n4569_o2_n,
    n4569_o2
  );


  buf

  (
    n4571_o2_p,
    n4571_o2
  );


  not

  (
    n4571_o2_n,
    n4571_o2
  );


  buf

  (
    n4572_o2_p,
    n4572_o2
  );


  not

  (
    n4572_o2_n,
    n4572_o2
  );


  buf

  (
    n399_inv_p,
    n399_inv
  );


  not

  (
    n399_inv_n,
    n399_inv
  );


  buf

  (
    n4539_o2_p,
    n4539_o2
  );


  not

  (
    n4539_o2_n,
    n4539_o2
  );


  buf

  (
    n4651_o2_p,
    n4651_o2
  );


  not

  (
    n4651_o2_n,
    n4651_o2
  );


  buf

  (
    n4652_o2_p,
    n4652_o2
  );


  not

  (
    n4652_o2_n,
    n4652_o2
  );


  buf

  (
    n4653_o2_p,
    n4653_o2
  );


  not

  (
    n4653_o2_n,
    n4653_o2
  );


  buf

  (
    G1514_o2_p,
    G1514_o2
  );


  not

  (
    G1514_o2_n,
    G1514_o2
  );


  buf

  (
    G1823_o2_p,
    G1823_o2
  );


  not

  (
    G1823_o2_n,
    G1823_o2
  );


  buf

  (
    n4783_o2_p,
    n4783_o2
  );


  not

  (
    n4783_o2_n,
    n4783_o2
  );


  buf

  (
    n4787_o2_p,
    n4787_o2
  );


  not

  (
    n4787_o2_n,
    n4787_o2
  );


  buf

  (
    n426_inv_p,
    n426_inv
  );


  not

  (
    n426_inv_n,
    n426_inv
  );


  buf

  (
    n429_inv_p,
    n429_inv
  );


  not

  (
    n429_inv_n,
    n429_inv
  );


  buf

  (
    n4816_o2_p,
    n4816_o2
  );


  not

  (
    n4816_o2_n,
    n4816_o2
  );


  buf

  (
    n435_inv_p,
    n435_inv
  );


  not

  (
    n435_inv_n,
    n435_inv
  );


  buf

  (
    G572_o2_p,
    G572_o2
  );


  not

  (
    G572_o2_n,
    G572_o2
  );


  buf

  (
    n4919_o2_p,
    n4919_o2
  );


  not

  (
    n4919_o2_n,
    n4919_o2
  );


  buf

  (
    n4920_o2_p,
    n4920_o2
  );


  not

  (
    n4920_o2_n,
    n4920_o2
  );


  buf

  (
    n4921_o2_p,
    n4921_o2
  );


  not

  (
    n4921_o2_n,
    n4921_o2
  );


  buf

  (
    G1048_o2_p,
    G1048_o2
  );


  not

  (
    G1048_o2_n,
    G1048_o2
  );


  buf

  (
    n5041_o2_p,
    n5041_o2
  );


  not

  (
    n5041_o2_n,
    n5041_o2
  );


  buf

  (
    n5094_o2_p,
    n5094_o2
  );


  not

  (
    n5094_o2_n,
    n5094_o2
  );


  buf

  (
    n5278_o2_p,
    n5278_o2
  );


  not

  (
    n5278_o2_n,
    n5278_o2
  );


  buf

  (
    n5301_o2_p,
    n5301_o2
  );


  not

  (
    n5301_o2_n,
    n5301_o2
  );


  buf

  (
    G2610_o2_p,
    G2610_o2
  );


  not

  (
    G2610_o2_n,
    G2610_o2
  );


  buf

  (
    G3174_o2_p,
    G3174_o2
  );


  not

  (
    G3174_o2_n,
    G3174_o2
  );


  buf

  (
    G3146_o2_p,
    G3146_o2
  );


  not

  (
    G3146_o2_n,
    G3146_o2
  );


  buf

  (
    G3217_o2_p,
    G3217_o2
  );


  not

  (
    G3217_o2_n,
    G3217_o2
  );


  buf

  (
    G3220_o2_p,
    G3220_o2
  );


  not

  (
    G3220_o2_n,
    G3220_o2
  );


  buf

  (
    G2839_o2_p,
    G2839_o2
  );


  not

  (
    G2839_o2_n,
    G2839_o2
  );


  buf

  (
    G3251_o2_p,
    G3251_o2
  );


  not

  (
    G3251_o2_n,
    G3251_o2
  );


  buf

  (
    G3042_o2_p,
    G3042_o2
  );


  not

  (
    G3042_o2_n,
    G3042_o2
  );


  buf

  (
    G3045_o2_p,
    G3045_o2
  );


  not

  (
    G3045_o2_n,
    G3045_o2
  );


  buf

  (
    G3262_o2_p,
    G3262_o2
  );


  not

  (
    G3262_o2_n,
    G3262_o2
  );


  buf

  (
    G2845_o2_p,
    G2845_o2
  );


  not

  (
    G2845_o2_n,
    G2845_o2
  );


  buf

  (
    G2929_o2_p,
    G2929_o2
  );


  not

  (
    G2929_o2_n,
    G2929_o2
  );


  buf

  (
    G2848_o2_p,
    G2848_o2
  );


  not

  (
    G2848_o2_n,
    G2848_o2
  );


  buf

  (
    G2851_o2_p,
    G2851_o2
  );


  not

  (
    G2851_o2_n,
    G2851_o2
  );


  buf

  (
    G3291_o2_p,
    G3291_o2
  );


  not

  (
    G3291_o2_n,
    G3291_o2
  );


  buf

  (
    G3254_o2_p,
    G3254_o2
  );


  not

  (
    G3254_o2_n,
    G3254_o2
  );


  buf

  (
    G2666_o2_p,
    G2666_o2
  );


  not

  (
    G2666_o2_n,
    G2666_o2
  );


  buf

  (
    n5099_o2_p,
    n5099_o2
  );


  not

  (
    n5099_o2_n,
    n5099_o2
  );


  buf

  (
    n5100_o2_p,
    n5100_o2
  );


  not

  (
    n5100_o2_n,
    n5100_o2
  );


  buf

  (
    n5101_o2_p,
    n5101_o2
  );


  not

  (
    n5101_o2_n,
    n5101_o2
  );


  buf

  (
    G2558_o2_p,
    G2558_o2
  );


  not

  (
    G2558_o2_n,
    G2558_o2
  );


  buf

  (
    n5266_o2_p,
    n5266_o2
  );


  not

  (
    n5266_o2_n,
    n5266_o2
  );


  buf

  (
    n5267_o2_p,
    n5267_o2
  );


  not

  (
    n5267_o2_n,
    n5267_o2
  );


  buf

  (
    G2759_o2_p,
    G2759_o2
  );


  not

  (
    G2759_o2_n,
    G2759_o2
  );


  buf

  (
    n537_inv_p,
    n537_inv
  );


  not

  (
    n537_inv_n,
    n537_inv
  );


  buf

  (
    n540_inv_p,
    n540_inv
  );


  not

  (
    n540_inv_n,
    n540_inv
  );


  buf

  (
    n543_inv_p,
    n543_inv
  );


  not

  (
    n543_inv_n,
    n543_inv
  );


  buf

  (
    n5292_o2_p,
    n5292_o2
  );


  not

  (
    n5292_o2_n,
    n5292_o2
  );


  buf

  (
    n5293_o2_p,
    n5293_o2
  );


  not

  (
    n5293_o2_n,
    n5293_o2
  );


  buf

  (
    n5294_o2_p,
    n5294_o2
  );


  not

  (
    n5294_o2_n,
    n5294_o2
  );


  buf

  (
    n5295_o2_p,
    n5295_o2
  );


  not

  (
    n5295_o2_n,
    n5295_o2
  );


  buf

  (
    G618_o2_p,
    G618_o2
  );


  not

  (
    G618_o2_n,
    G618_o2
  );


  buf

  (
    G621_o2_p,
    G621_o2
  );


  not

  (
    G621_o2_n,
    G621_o2
  );


  buf

  (
    G384_o2_p,
    G384_o2
  );


  not

  (
    G384_o2_n,
    G384_o2
  );


  buf

  (
    G377_o2_p,
    G377_o2
  );


  not

  (
    G377_o2_n,
    G377_o2
  );


  buf

  (
    n570_inv_p,
    n570_inv
  );


  not

  (
    n570_inv_n,
    n570_inv
  );


  buf

  (
    G3171_o2_p,
    G3171_o2
  );


  not

  (
    G3171_o2_n,
    G3171_o2
  );


  buf

  (
    G2552_o2_p,
    G2552_o2
  );


  not

  (
    G2552_o2_n,
    G2552_o2
  );


  buf

  (
    G3272_o2_p,
    G3272_o2
  );


  not

  (
    G3272_o2_n,
    G3272_o2
  );


  buf

  (
    G2015_o2_p,
    G2015_o2
  );


  not

  (
    G2015_o2_n,
    G2015_o2
  );


  buf

  (
    G3294_o2_p,
    G3294_o2
  );


  not

  (
    G3294_o2_n,
    G3294_o2
  );


  buf

  (
    G3281_o2_p,
    G3281_o2
  );


  not

  (
    G3281_o2_n,
    G3281_o2
  );


  buf

  (
    G3320_o2_p,
    G3320_o2
  );


  not

  (
    G3320_o2_n,
    G3320_o2
  );


  buf

  (
    G3275_o2_p,
    G3275_o2
  );


  not

  (
    G3275_o2_n,
    G3275_o2
  );


  buf

  (
    G3140_o2_p,
    G3140_o2
  );


  not

  (
    G3140_o2_n,
    G3140_o2
  );


  buf

  (
    G2836_o2_p,
    G2836_o2
  );


  not

  (
    G2836_o2_n,
    G2836_o2
  );


  buf

  (
    G2926_o2_p,
    G2926_o2
  );


  not

  (
    G2926_o2_n,
    G2926_o2
  );


  buf

  (
    G2842_o2_p,
    G2842_o2
  );


  not

  (
    G2842_o2_n,
    G2842_o2
  );


  buf

  (
    G3302_o2_p,
    G3302_o2
  );


  not

  (
    G3302_o2_n,
    G3302_o2
  );


  buf

  (
    G3288_o2_p,
    G3288_o2
  );


  not

  (
    G3288_o2_n,
    G3288_o2
  );


  buf

  (
    G3143_o2_p,
    G3143_o2
  );


  not

  (
    G3143_o2_n,
    G3143_o2
  );


  buf

  (
    G3100_o2_p,
    G3100_o2
  );


  not

  (
    G3100_o2_n,
    G3100_o2
  );


  buf

  (
    G2512_o2_p,
    G2512_o2
  );


  not

  (
    G2512_o2_n,
    G2512_o2
  );


  buf

  (
    n5325_o2_p,
    n5325_o2
  );


  not

  (
    n5325_o2_n,
    n5325_o2
  );


  buf

  (
    n5326_o2_p,
    n5326_o2
  );


  not

  (
    n5326_o2_n,
    n5326_o2
  );


  buf

  (
    n5327_o2_p,
    n5327_o2
  );


  not

  (
    n5327_o2_n,
    n5327_o2
  );


  buf

  (
    n1857_lo_buf_o2_p,
    n1857_lo_buf_o2
  );


  not

  (
    n1857_lo_buf_o2_n,
    n1857_lo_buf_o2
  );


  buf

  (
    n2097_lo_buf_o2_p,
    n2097_lo_buf_o2
  );


  not

  (
    n2097_lo_buf_o2_n,
    n2097_lo_buf_o2
  );


  buf

  (
    G2669_o2_p,
    G2669_o2
  );


  not

  (
    G2669_o2_n,
    G2669_o2
  );


  buf

  (
    n642_inv_p,
    n642_inv
  );


  not

  (
    n642_inv_n,
    n642_inv
  );


  buf

  (
    G568_o2_p,
    G568_o2
  );


  not

  (
    G568_o2_n,
    G568_o2
  );


  buf

  (
    n648_inv_p,
    n648_inv
  );


  not

  (
    n648_inv_n,
    n648_inv
  );


  buf

  (
    G565_o2_p,
    G565_o2
  );


  not

  (
    G565_o2_n,
    G565_o2
  );


  buf

  (
    G559_o2_p,
    G559_o2
  );


  not

  (
    G559_o2_n,
    G559_o2
  );


  buf

  (
    n1821_lo_buf_o2_p,
    n1821_lo_buf_o2
  );


  not

  (
    n1821_lo_buf_o2_n,
    n1821_lo_buf_o2
  );


  buf

  (
    n1905_lo_buf_o2_p,
    n1905_lo_buf_o2
  );


  not

  (
    n1905_lo_buf_o2_n,
    n1905_lo_buf_o2
  );


  buf

  (
    n2133_lo_buf_o2_p,
    n2133_lo_buf_o2
  );


  not

  (
    n2133_lo_buf_o2_n,
    n2133_lo_buf_o2
  );


  buf

  (
    n2145_lo_buf_o2_p,
    n2145_lo_buf_o2
  );


  not

  (
    n2145_lo_buf_o2_n,
    n2145_lo_buf_o2
  );


  buf

  (
    n2157_lo_buf_o2_p,
    n2157_lo_buf_o2
  );


  not

  (
    n2157_lo_buf_o2_n,
    n2157_lo_buf_o2
  );


  buf

  (
    n2205_lo_buf_o2_p,
    n2205_lo_buf_o2
  );


  not

  (
    n2205_lo_buf_o2_n,
    n2205_lo_buf_o2
  );


  buf

  (
    n2217_lo_buf_o2_p,
    n2217_lo_buf_o2
  );


  not

  (
    n2217_lo_buf_o2_n,
    n2217_lo_buf_o2
  );


  buf

  (
    G447_o2_p,
    G447_o2
  );


  not

  (
    G447_o2_n,
    G447_o2
  );


  buf

  (
    G434_o2_p,
    G434_o2
  );


  not

  (
    G434_o2_n,
    G434_o2
  );


  buf

  (
    G422_o2_p,
    G422_o2
  );


  not

  (
    G422_o2_n,
    G422_o2
  );


  buf

  (
    G461_o2_p,
    G461_o2
  );


  not

  (
    G461_o2_n,
    G461_o2
  );


  buf

  (
    G3312_o2_p,
    G3312_o2
  );


  not

  (
    G3312_o2_n,
    G3312_o2
  );


  buf

  (
    G3332_o2_p,
    G3332_o2
  );


  not

  (
    G3332_o2_n,
    G3332_o2
  );


  buf

  (
    G3195_o2_p,
    G3195_o2
  );


  not

  (
    G3195_o2_n,
    G3195_o2
  );


  buf

  (
    G2607_o2_p,
    G2607_o2
  );


  not

  (
    G2607_o2_n,
    G2607_o2
  );


  buf

  (
    n702_inv_p,
    n702_inv
  );


  not

  (
    n702_inv_n,
    n702_inv
  );


  buf

  (
    G1005_o2_p,
    G1005_o2
  );


  not

  (
    G1005_o2_n,
    G1005_o2
  );


  buf

  (
    G1008_o2_p,
    G1008_o2
  );


  not

  (
    G1008_o2_n,
    G1008_o2
  );


  buf

  (
    n2001_lo_buf_o2_p,
    n2001_lo_buf_o2
  );


  not

  (
    n2001_lo_buf_o2_n,
    n2001_lo_buf_o2
  );


  buf

  (
    n2169_lo_buf_o2_p,
    n2169_lo_buf_o2
  );


  not

  (
    n2169_lo_buf_o2_n,
    n2169_lo_buf_o2
  );


  buf

  (
    n2229_lo_buf_o2_p,
    n2229_lo_buf_o2
  );


  not

  (
    n2229_lo_buf_o2_n,
    n2229_lo_buf_o2
  );


  buf

  (
    n2301_lo_buf_o2_p,
    n2301_lo_buf_o2
  );


  not

  (
    n2301_lo_buf_o2_n,
    n2301_lo_buf_o2
  );


  buf

  (
    n723_inv_p,
    n723_inv
  );


  not

  (
    n723_inv_n,
    n723_inv
  );


  buf

  (
    G2947_o2_p,
    G2947_o2
  );


  not

  (
    G2947_o2_n,
    G2947_o2
  );


  buf

  (
    n2013_lo_buf_o2_p,
    n2013_lo_buf_o2
  );


  not

  (
    n2013_lo_buf_o2_n,
    n2013_lo_buf_o2
  );


  buf

  (
    n2025_lo_buf_o2_p,
    n2025_lo_buf_o2
  );


  not

  (
    n2025_lo_buf_o2_n,
    n2025_lo_buf_o2
  );


  buf

  (
    n2037_lo_buf_o2_p,
    n2037_lo_buf_o2
  );


  not

  (
    n2037_lo_buf_o2_n,
    n2037_lo_buf_o2
  );


  buf

  (
    n2049_lo_buf_o2_p,
    n2049_lo_buf_o2
  );


  not

  (
    n2049_lo_buf_o2_n,
    n2049_lo_buf_o2
  );


  buf

  (
    n2181_lo_buf_o2_p,
    n2181_lo_buf_o2
  );


  not

  (
    n2181_lo_buf_o2_n,
    n2181_lo_buf_o2
  );


  buf

  (
    n744_inv_p,
    n744_inv
  );


  not

  (
    n744_inv_n,
    n744_inv
  );


  buf

  (
    n747_inv_p,
    n747_inv
  );


  not

  (
    n747_inv_n,
    n747_inv
  );


  buf

  (
    n750_inv_p,
    n750_inv
  );


  not

  (
    n750_inv_n,
    n750_inv
  );


  buf

  (
    n753_inv_p,
    n753_inv
  );


  not

  (
    n753_inv_n,
    n753_inv
  );


  buf

  (
    G3350_o2_p,
    G3350_o2
  );


  not

  (
    G3350_o2_n,
    G3350_o2
  );


  buf

  (
    G3360_o2_p,
    G3360_o2
  );


  not

  (
    G3360_o2_n,
    G3360_o2
  );


  buf

  (
    G3373_o2_p,
    G3373_o2
  );


  not

  (
    G3373_o2_n,
    G3373_o2
  );


  buf

  (
    G3237_o2_p,
    G3237_o2
  );


  not

  (
    G3237_o2_n,
    G3237_o2
  );


  buf

  (
    G2773_o2_p,
    G2773_o2
  );


  not

  (
    G2773_o2_n,
    G2773_o2
  );


  buf

  (
    G1733_o2_p,
    G1733_o2
  );


  not

  (
    G1733_o2_n,
    G1733_o2
  );


  buf

  (
    G1738_o2_p,
    G1738_o2
  );


  not

  (
    G1738_o2_n,
    G1738_o2
  );


  buf

  (
    G1751_o2_p,
    G1751_o2
  );


  not

  (
    G1751_o2_n,
    G1751_o2
  );


  buf

  (
    G2216_o2_p,
    G2216_o2
  );


  not

  (
    G2216_o2_n,
    G2216_o2
  );


  buf

  (
    G2219_o2_p,
    G2219_o2
  );


  not

  (
    G2219_o2_n,
    G2219_o2
  );


  buf

  (
    n786_inv_p,
    n786_inv
  );


  not

  (
    n786_inv_n,
    n786_inv
  );


  buf

  (
    n789_inv_p,
    n789_inv
  );


  not

  (
    n789_inv_n,
    n789_inv
  );


  buf

  (
    G787_o2_p,
    G787_o2
  );


  not

  (
    G787_o2_n,
    G787_o2
  );


  buf

  (
    G2823_o2_p,
    G2823_o2
  );


  not

  (
    G2823_o2_n,
    G2823_o2
  );


  buf

  (
    G2796_o2_p,
    G2796_o2
  );


  not

  (
    G2796_o2_n,
    G2796_o2
  );


  buf

  (
    G875_o2_p,
    G875_o2
  );


  not

  (
    G875_o2_n,
    G875_o2
  );


  buf

  (
    G2208_o2_p,
    G2208_o2
  );


  not

  (
    G2208_o2_n,
    G2208_o2
  );


  buf

  (
    G2211_o2_p,
    G2211_o2
  );


  not

  (
    G2211_o2_n,
    G2211_o2
  );


  buf

  (
    n1989_lo_buf_o2_p,
    n1989_lo_buf_o2
  );


  not

  (
    n1989_lo_buf_o2_n,
    n1989_lo_buf_o2
  );


  buf

  (
    n2061_lo_buf_o2_p,
    n2061_lo_buf_o2
  );


  not

  (
    n2061_lo_buf_o2_n,
    n2061_lo_buf_o2
  );


  buf

  (
    n2313_lo_buf_o2_p,
    n2313_lo_buf_o2
  );


  not

  (
    n2313_lo_buf_o2_n,
    n2313_lo_buf_o2
  );


  buf

  (
    G2232_o2_p,
    G2232_o2
  );


  not

  (
    G2232_o2_n,
    G2232_o2
  );


  buf

  (
    G1725_o2_p,
    G1725_o2
  );


  not

  (
    G1725_o2_n,
    G1725_o2
  );


  buf

  (
    G1764_o2_p,
    G1764_o2
  );


  not

  (
    G1764_o2_n,
    G1764_o2
  );


  buf

  (
    G2356_o2_p,
    G2356_o2
  );


  not

  (
    G2356_o2_n,
    G2356_o2
  );


  buf

  (
    G2359_o2_p,
    G2359_o2
  );


  not

  (
    G2359_o2_n,
    G2359_o2
  );


  buf

  (
    G1180_o2_p,
    G1180_o2
  );


  not

  (
    G1180_o2_n,
    G1180_o2
  );


  buf

  (
    G1756_o2_p,
    G1756_o2
  );


  not

  (
    G1756_o2_n,
    G1756_o2
  );


  buf

  (
    G2441_o2_p,
    G2441_o2
  );


  not

  (
    G2441_o2_n,
    G2441_o2
  );


  buf

  (
    G2887_o2_p,
    G2887_o2
  );


  not

  (
    G2887_o2_n,
    G2887_o2
  );


  buf

  (
    G2991_o2_p,
    G2991_o2
  );


  not

  (
    G2991_o2_n,
    G2991_o2
  );


  buf

  (
    n849_inv_p,
    n849_inv
  );


  not

  (
    n849_inv_n,
    n849_inv
  );


  buf

  (
    n852_inv_p,
    n852_inv
  );


  not

  (
    n852_inv_n,
    n852_inv
  );


  buf

  (
    n855_inv_p,
    n855_inv
  );


  not

  (
    n855_inv_n,
    n855_inv
  );


  buf

  (
    n858_inv_p,
    n858_inv
  );


  not

  (
    n858_inv_n,
    n858_inv
  );


  buf

  (
    n861_inv_p,
    n861_inv
  );


  not

  (
    n861_inv_n,
    n861_inv
  );


  buf

  (
    G2805_o2_p,
    G2805_o2
  );


  not

  (
    G2805_o2_n,
    G2805_o2
  );


  buf

  (
    G2906_o2_p,
    G2906_o2
  );


  not

  (
    G2906_o2_n,
    G2906_o2
  );


  buf

  (
    G2833_o2_p,
    G2833_o2
  );


  not

  (
    G2833_o2_n,
    G2833_o2
  );


  buf

  (
    n873_inv_p,
    n873_inv
  );


  not

  (
    n873_inv_n,
    n873_inv
  );


  buf

  (
    G3353_o2_p,
    G3353_o2
  );


  not

  (
    G3353_o2_n,
    G3353_o2
  );


  buf

  (
    G3367_o2_p,
    G3367_o2
  );


  not

  (
    G3367_o2_n,
    G3367_o2
  );


  buf

  (
    G3346_o2_p,
    G3346_o2
  );


  not

  (
    G3346_o2_n,
    G3346_o2
  );


  buf

  (
    G3340_o2_p,
    G3340_o2
  );


  not

  (
    G3340_o2_n,
    G3340_o2
  );


  buf

  (
    G3376_o2_p,
    G3376_o2
  );


  not

  (
    G3376_o2_n,
    G3376_o2
  );


  buf

  (
    G3359_o2_p,
    G3359_o2
  );


  not

  (
    G3359_o2_n,
    G3359_o2
  );


  buf

  (
    G3240_o2_p,
    G3240_o2
  );


  not

  (
    G3240_o2_n,
    G3240_o2
  );


  buf

  (
    G3344_o2_p,
    G3344_o2
  );


  not

  (
    G3344_o2_n,
    G3344_o2
  );


  buf

  (
    G2880_o2_p,
    G2880_o2
  );


  not

  (
    G2880_o2_n,
    G2880_o2
  );


  buf

  (
    G2939_o2_p,
    G2939_o2
  );


  not

  (
    G2939_o2_n,
    G2939_o2
  );


  buf

  (
    G2248_o2_p,
    G2248_o2
  );


  not

  (
    G2248_o2_n,
    G2248_o2
  );


  buf

  (
    G2251_o2_p,
    G2251_o2
  );


  not

  (
    G2251_o2_n,
    G2251_o2
  );


  buf

  (
    G2021_o2_p,
    G2021_o2
  );


  not

  (
    G2021_o2_n,
    G2021_o2
  );


  buf

  (
    G3383_o2_p,
    G3383_o2
  );


  not

  (
    G3383_o2_n,
    G3383_o2
  );


  buf

  (
    G3399_o2_p,
    G3399_o2
  );


  not

  (
    G3399_o2_n,
    G3399_o2
  );


  buf

  (
    G3404_o2_p,
    G3404_o2
  );


  not

  (
    G3404_o2_n,
    G3404_o2
  );


  buf

  (
    G3265_o2_p,
    G3265_o2
  );


  not

  (
    G3265_o2_n,
    G3265_o2
  );


  buf

  (
    G2866_o2_p,
    G2866_o2
  );


  not

  (
    G2866_o2_n,
    G2866_o2
  );


  buf

  (
    G2999_o2_p,
    G2999_o2
  );


  not

  (
    G2999_o2_n,
    G2999_o2
  );


  buf

  (
    G736_o2_p,
    G736_o2
  );


  not

  (
    G736_o2_n,
    G736_o2
  );


  buf

  (
    G739_o2_p,
    G739_o2
  );


  not

  (
    G739_o2_n,
    G739_o2
  );


  buf

  (
    G1200_o2_p,
    G1200_o2
  );


  not

  (
    G1200_o2_n,
    G1200_o2
  );


  buf

  (
    G1203_o2_p,
    G1203_o2
  );


  not

  (
    G1203_o2_n,
    G1203_o2
  );


  buf

  (
    G3027_o2_p,
    G3027_o2
  );


  not

  (
    G3027_o2_n,
    G3027_o2
  );


  buf

  (
    G1463_o2_p,
    G1463_o2
  );


  not

  (
    G1463_o2_n,
    G1463_o2
  );


  buf

  (
    G1460_o2_p,
    G1460_o2
  );


  not

  (
    G1460_o2_n,
    G1460_o2
  );


  buf

  (
    G3012_o2_p,
    G3012_o2
  );


  not

  (
    G3012_o2_n,
    G3012_o2
  );


  buf

  (
    G1574_o2_p,
    G1574_o2
  );


  not

  (
    G1574_o2_n,
    G1574_o2
  );


  buf

  (
    G1646_o2_p,
    G1646_o2
  );


  not

  (
    G1646_o2_n,
    G1646_o2
  );


  buf

  (
    G1592_o2_p,
    G1592_o2
  );


  not

  (
    G1592_o2_n,
    G1592_o2
  );


  buf

  (
    G1664_o2_p,
    G1664_o2
  );


  not

  (
    G1664_o2_n,
    G1664_o2
  );


  buf

  (
    G1547_o2_p,
    G1547_o2
  );


  not

  (
    G1547_o2_n,
    G1547_o2
  );


  buf

  (
    G1619_o2_p,
    G1619_o2
  );


  not

  (
    G1619_o2_n,
    G1619_o2
  );


  buf

  (
    G1556_o2_p,
    G1556_o2
  );


  not

  (
    G1556_o2_n,
    G1556_o2
  );


  buf

  (
    G1628_o2_p,
    G1628_o2
  );


  not

  (
    G1628_o2_n,
    G1628_o2
  );


  buf

  (
    G1583_o2_p,
    G1583_o2
  );


  not

  (
    G1583_o2_n,
    G1583_o2
  );


  buf

  (
    G1655_o2_p,
    G1655_o2
  );


  not

  (
    G1655_o2_n,
    G1655_o2
  );


  buf

  (
    G1529_o2_p,
    G1529_o2
  );


  not

  (
    G1529_o2_n,
    G1529_o2
  );


  buf

  (
    G1601_o2_p,
    G1601_o2
  );


  not

  (
    G1601_o2_n,
    G1601_o2
  );


  buf

  (
    G1538_o2_p,
    G1538_o2
  );


  not

  (
    G1538_o2_n,
    G1538_o2
  );


  buf

  (
    G1610_o2_p,
    G1610_o2
  );


  not

  (
    G1610_o2_n,
    G1610_o2
  );


  buf

  (
    G1565_o2_p,
    G1565_o2
  );


  not

  (
    G1565_o2_n,
    G1565_o2
  );


  buf

  (
    G1637_o2_p,
    G1637_o2
  );


  not

  (
    G1637_o2_n,
    G1637_o2
  );


  buf

  (
    G2437_o2_p,
    G2437_o2
  );


  not

  (
    G2437_o2_n,
    G2437_o2
  );


  buf

  (
    n1008_inv_p,
    n1008_inv
  );


  not

  (
    n1008_inv_n,
    n1008_inv
  );


  buf

  (
    n1785_lo_buf_o2_p,
    n1785_lo_buf_o2
  );


  not

  (
    n1785_lo_buf_o2_n,
    n1785_lo_buf_o2
  );


  buf

  (
    n1845_lo_buf_o2_p,
    n1845_lo_buf_o2
  );


  not

  (
    n1845_lo_buf_o2_n,
    n1845_lo_buf_o2
  );


  buf

  (
    n1893_lo_buf_o2_p,
    n1893_lo_buf_o2
  );


  not

  (
    n1893_lo_buf_o2_n,
    n1893_lo_buf_o2
  );


  buf

  (
    n1941_lo_buf_o2_p,
    n1941_lo_buf_o2
  );


  not

  (
    n1941_lo_buf_o2_n,
    n1941_lo_buf_o2
  );


  buf

  (
    n1953_lo_buf_o2_p,
    n1953_lo_buf_o2
  );


  not

  (
    n1953_lo_buf_o2_n,
    n1953_lo_buf_o2
  );


  buf

  (
    n1965_lo_buf_o2_p,
    n1965_lo_buf_o2
  );


  not

  (
    n1965_lo_buf_o2_n,
    n1965_lo_buf_o2
  );


  buf

  (
    n1977_lo_buf_o2_p,
    n1977_lo_buf_o2
  );


  not

  (
    n1977_lo_buf_o2_n,
    n1977_lo_buf_o2
  );


  buf

  (
    n2241_lo_buf_o2_p,
    n2241_lo_buf_o2
  );


  not

  (
    n2241_lo_buf_o2_n,
    n2241_lo_buf_o2
  );


  buf

  (
    n2253_lo_buf_o2_p,
    n2253_lo_buf_o2
  );


  not

  (
    n2253_lo_buf_o2_n,
    n2253_lo_buf_o2
  );


  buf

  (
    n2265_lo_buf_o2_p,
    n2265_lo_buf_o2
  );


  not

  (
    n2265_lo_buf_o2_n,
    n2265_lo_buf_o2
  );


  buf

  (
    n2277_lo_buf_o2_p,
    n2277_lo_buf_o2
  );


  not

  (
    n2277_lo_buf_o2_n,
    n2277_lo_buf_o2
  );


  buf

  (
    n2289_lo_buf_o2_p,
    n2289_lo_buf_o2
  );


  not

  (
    n2289_lo_buf_o2_n,
    n2289_lo_buf_o2
  );


  buf

  (
    G519_o2_p,
    G519_o2
  );


  not

  (
    G519_o2_n,
    G519_o2
  );


  buf

  (
    n1050_inv_p,
    n1050_inv
  );


  not

  (
    n1050_inv_n,
    n1050_inv
  );


  buf

  (
    n1053_inv_p,
    n1053_inv
  );


  not

  (
    n1053_inv_n,
    n1053_inv
  );


  buf

  (
    n1056_inv_p,
    n1056_inv
  );


  not

  (
    n1056_inv_n,
    n1056_inv
  );


  buf

  (
    G1318_o2_p,
    G1318_o2
  );


  not

  (
    G1318_o2_n,
    G1318_o2
  );


  buf

  (
    n1062_inv_p,
    n1062_inv
  );


  not

  (
    n1062_inv_n,
    n1062_inv
  );


  buf

  (
    G593_o2_p,
    G593_o2
  );


  not

  (
    G593_o2_n,
    G593_o2
  );


  buf

  (
    n1068_inv_p,
    n1068_inv
  );


  not

  (
    n1068_inv_n,
    n1068_inv
  );


  buf

  (
    n1071_inv_p,
    n1071_inv
  );


  not

  (
    n1071_inv_n,
    n1071_inv
  );


  buf

  (
    n1074_inv_p,
    n1074_inv
  );


  not

  (
    n1074_inv_n,
    n1074_inv
  );


  buf

  (
    G2284_o2_p,
    G2284_o2
  );


  not

  (
    G2284_o2_n,
    G2284_o2
  );


  buf

  (
    G2580_o2_p,
    G2580_o2
  );


  not

  (
    G2580_o2_n,
    G2580_o2
  );


  buf

  (
    G2302_o2_p,
    G2302_o2
  );


  not

  (
    G2302_o2_n,
    G2302_o2
  );


  buf

  (
    G2598_o2_p,
    G2598_o2
  );


  not

  (
    G2598_o2_n,
    G2598_o2
  );


  buf

  (
    G2497_o2_p,
    G2497_o2
  );


  not

  (
    G2497_o2_n,
    G2497_o2
  );


  buf

  (
    G2651_o2_p,
    G2651_o2
  );


  not

  (
    G2651_o2_n,
    G2651_o2
  );


  buf

  (
    G2296_o2_p,
    G2296_o2
  );


  not

  (
    G2296_o2_n,
    G2296_o2
  );


  buf

  (
    G2308_o2_p,
    G2308_o2
  );


  not

  (
    G2308_o2_n,
    G2308_o2
  );


  buf

  (
    G2592_o2_p,
    G2592_o2
  );


  not

  (
    G2592_o2_n,
    G2592_o2
  );


  buf

  (
    G2604_o2_p,
    G2604_o2
  );


  not

  (
    G2604_o2_n,
    G2604_o2
  );


  buf

  (
    G2902_o2_p,
    G2902_o2
  );


  not

  (
    G2902_o2_n,
    G2902_o2
  );


  buf

  (
    G2975_o2_p,
    G2975_o2
  );


  not

  (
    G2975_o2_n,
    G2975_o2
  );


  buf

  (
    G2962_o2_p,
    G2962_o2
  );


  not

  (
    G2962_o2_n,
    G2962_o2
  );


  buf

  (
    G3069_o2_p,
    G3069_o2
  );


  not

  (
    G3069_o2_n,
    G3069_o2
  );


  buf

  (
    G2018_o2_p,
    G2018_o2
  );


  not

  (
    G2018_o2_n,
    G2018_o2
  );


  buf

  (
    G1176_o2_p,
    G1176_o2
  );


  not

  (
    G1176_o2_n,
    G1176_o2
  );


  buf

  (
    G1189_o2_p,
    G1189_o2
  );


  not

  (
    G1189_o2_n,
    G1189_o2
  );


  buf

  (
    G3066_o2_p,
    G3066_o2
  );


  not

  (
    G3066_o2_n,
    G3066_o2
  );


  buf

  (
    G3137_o2_p,
    G3137_o2
  );


  not

  (
    G3137_o2_n,
    G3137_o2
  );


  buf

  (
    G3038_o2_p,
    G3038_o2
  );


  not

  (
    G3038_o2_n,
    G3038_o2
  );


  buf

  (
    G3117_o2_p,
    G3117_o2
  );


  not

  (
    G3117_o2_n,
    G3117_o2
  );


  buf

  (
    G2384_o2_p,
    G2384_o2
  );


  not

  (
    G2384_o2_n,
    G2384_o2
  );


  buf

  (
    G2472_o2_p,
    G2472_o2
  );


  not

  (
    G2472_o2_n,
    G2472_o2
  );


  buf

  (
    G772_o2_p,
    G772_o2
  );


  not

  (
    G772_o2_n,
    G772_o2
  );


  buf

  (
    G935_o2_p,
    G935_o2
  );


  not

  (
    G935_o2_n,
    G935_o2
  );


  buf

  (
    G2923_o2_p,
    G2923_o2
  );


  not

  (
    G2923_o2_n,
    G2923_o2
  );


  buf

  (
    G2971_o2_p,
    G2971_o2
  );


  not

  (
    G2971_o2_n,
    G2971_o2
  );


  buf

  (
    G2980_o2_p,
    G2980_o2
  );


  not

  (
    G2980_o2_n,
    G2980_o2
  );


  buf

  (
    G3039_o2_p,
    G3039_o2
  );


  not

  (
    G3039_o2_n,
    G3039_o2
  );


  buf

  (
    G2388_o2_p,
    G2388_o2
  );


  not

  (
    G2388_o2_n,
    G2388_o2
  );


  buf

  (
    G2287_o2_p,
    G2287_o2
  );


  not

  (
    G2287_o2_n,
    G2287_o2
  );


  buf

  (
    G3024_o2_p,
    G3024_o2
  );


  not

  (
    G3024_o2_n,
    G3024_o2
  );


  buf

  (
    G2916_o2_p,
    G2916_o2
  );


  not

  (
    G2916_o2_n,
    G2916_o2
  );


  buf

  (
    n1176_inv_p,
    n1176_inv
  );


  not

  (
    n1176_inv_n,
    n1176_inv
  );


  buf

  (
    G3035_o2_p,
    G3035_o2
  );


  not

  (
    G3035_o2_n,
    G3035_o2
  );


  buf

  (
    G3107_o2_p,
    G3107_o2
  );


  not

  (
    G3107_o2_n,
    G3107_o2
  );


  buf

  (
    G1023_o2_p,
    G1023_o2
  );


  not

  (
    G1023_o2_n,
    G1023_o2
  );


  buf

  (
    G1024_o2_p,
    G1024_o2
  );


  not

  (
    G1024_o2_n,
    G1024_o2
  );


  buf

  (
    G1311_o2_p,
    G1311_o2
  );


  not

  (
    G1311_o2_n,
    G1311_o2
  );


  buf

  (
    G1312_o2_p,
    G1312_o2
  );


  not

  (
    G1312_o2_n,
    G1312_o2
  );


  buf

  (
    G3063_o2_p,
    G3063_o2
  );


  not

  (
    G3063_o2_n,
    G3063_o2
  );


  buf

  (
    G1520_o2_p,
    G1520_o2
  );


  not

  (
    G1520_o2_n,
    G1520_o2
  );


  buf

  (
    G1519_o2_p,
    G1519_o2
  );


  not

  (
    G1519_o2_n,
    G1519_o2
  );


  buf

  (
    G3078_o2_p,
    G3078_o2
  );


  not

  (
    G3078_o2_n,
    G3078_o2
  );


  buf

  (
    G2038_o2_p,
    G2038_o2
  );


  not

  (
    G2038_o2_n,
    G2038_o2
  );


  buf

  (
    G1848_o2_p,
    G1848_o2
  );


  not

  (
    G1848_o2_n,
    G1848_o2
  );


  buf

  (
    G1864_o2_p,
    G1864_o2
  );


  not

  (
    G1864_o2_n,
    G1864_o2
  );


  buf

  (
    G1872_o2_p,
    G1872_o2
  );


  not

  (
    G1872_o2_n,
    G1872_o2
  );


  buf

  (
    G1880_o2_p,
    G1880_o2
  );


  not

  (
    G1880_o2_n,
    G1880_o2
  );


  buf

  (
    G1888_o2_p,
    G1888_o2
  );


  not

  (
    G1888_o2_n,
    G1888_o2
  );


  buf

  (
    G1912_o2_p,
    G1912_o2
  );


  not

  (
    G1912_o2_n,
    G1912_o2
  );


  buf

  (
    G1928_o2_p,
    G1928_o2
  );


  not

  (
    G1928_o2_n,
    G1928_o2
  );


  buf

  (
    G1936_o2_p,
    G1936_o2
  );


  not

  (
    G1936_o2_n,
    G1936_o2
  );


  buf

  (
    G1944_o2_p,
    G1944_o2
  );


  not

  (
    G1944_o2_n,
    G1944_o2
  );


  buf

  (
    G1952_o2_p,
    G1952_o2
  );


  not

  (
    G1952_o2_n,
    G1952_o2
  );


  buf

  (
    G1850_o2_p,
    G1850_o2
  );


  not

  (
    G1850_o2_n,
    G1850_o2
  );


  buf

  (
    G1866_o2_p,
    G1866_o2
  );


  not

  (
    G1866_o2_n,
    G1866_o2
  );


  buf

  (
    G1874_o2_p,
    G1874_o2
  );


  not

  (
    G1874_o2_n,
    G1874_o2
  );


  buf

  (
    G1882_o2_p,
    G1882_o2
  );


  not

  (
    G1882_o2_n,
    G1882_o2
  );


  buf

  (
    G1890_o2_p,
    G1890_o2
  );


  not

  (
    G1890_o2_n,
    G1890_o2
  );


  buf

  (
    G1914_o2_p,
    G1914_o2
  );


  not

  (
    G1914_o2_n,
    G1914_o2
  );


  buf

  (
    G1930_o2_p,
    G1930_o2
  );


  not

  (
    G1930_o2_n,
    G1930_o2
  );


  buf

  (
    G1938_o2_p,
    G1938_o2
  );


  not

  (
    G1938_o2_n,
    G1938_o2
  );


  buf

  (
    G1946_o2_p,
    G1946_o2
  );


  not

  (
    G1946_o2_n,
    G1946_o2
  );


  buf

  (
    G1954_o2_p,
    G1954_o2
  );


  not

  (
    G1954_o2_n,
    G1954_o2
  );


  buf

  (
    G1845_o2_p,
    G1845_o2
  );


  not

  (
    G1845_o2_n,
    G1845_o2
  );


  buf

  (
    G1861_o2_p,
    G1861_o2
  );


  not

  (
    G1861_o2_n,
    G1861_o2
  );


  buf

  (
    G1869_o2_p,
    G1869_o2
  );


  not

  (
    G1869_o2_n,
    G1869_o2
  );


  buf

  (
    G1877_o2_p,
    G1877_o2
  );


  not

  (
    G1877_o2_n,
    G1877_o2
  );


  buf

  (
    G1885_o2_p,
    G1885_o2
  );


  not

  (
    G1885_o2_n,
    G1885_o2
  );


  buf

  (
    G1909_o2_p,
    G1909_o2
  );


  not

  (
    G1909_o2_n,
    G1909_o2
  );


  buf

  (
    G1925_o2_p,
    G1925_o2
  );


  not

  (
    G1925_o2_n,
    G1925_o2
  );


  buf

  (
    G1933_o2_p,
    G1933_o2
  );


  not

  (
    G1933_o2_n,
    G1933_o2
  );


  buf

  (
    G1941_o2_p,
    G1941_o2
  );


  not

  (
    G1941_o2_n,
    G1941_o2
  );


  buf

  (
    G1949_o2_p,
    G1949_o2
  );


  not

  (
    G1949_o2_n,
    G1949_o2
  );


  buf

  (
    G1846_o2_p,
    G1846_o2
  );


  not

  (
    G1846_o2_n,
    G1846_o2
  );


  buf

  (
    G1862_o2_p,
    G1862_o2
  );


  not

  (
    G1862_o2_n,
    G1862_o2
  );


  buf

  (
    G1870_o2_p,
    G1870_o2
  );


  not

  (
    G1870_o2_n,
    G1870_o2
  );


  buf

  (
    G1878_o2_p,
    G1878_o2
  );


  not

  (
    G1878_o2_n,
    G1878_o2
  );


  buf

  (
    G1886_o2_p,
    G1886_o2
  );


  not

  (
    G1886_o2_n,
    G1886_o2
  );


  buf

  (
    G1910_o2_p,
    G1910_o2
  );


  not

  (
    G1910_o2_n,
    G1910_o2
  );


  buf

  (
    G1926_o2_p,
    G1926_o2
  );


  not

  (
    G1926_o2_n,
    G1926_o2
  );


  buf

  (
    G1934_o2_p,
    G1934_o2
  );


  not

  (
    G1934_o2_n,
    G1934_o2
  );


  buf

  (
    G1942_o2_p,
    G1942_o2
  );


  not

  (
    G1942_o2_n,
    G1942_o2
  );


  buf

  (
    G1950_o2_p,
    G1950_o2
  );


  not

  (
    G1950_o2_n,
    G1950_o2
  );


  buf

  (
    G1849_o2_p,
    G1849_o2
  );


  not

  (
    G1849_o2_n,
    G1849_o2
  );


  buf

  (
    G1865_o2_p,
    G1865_o2
  );


  not

  (
    G1865_o2_n,
    G1865_o2
  );


  buf

  (
    G1873_o2_p,
    G1873_o2
  );


  not

  (
    G1873_o2_n,
    G1873_o2
  );


  buf

  (
    G1881_o2_p,
    G1881_o2
  );


  not

  (
    G1881_o2_n,
    G1881_o2
  );


  buf

  (
    G1889_o2_p,
    G1889_o2
  );


  not

  (
    G1889_o2_n,
    G1889_o2
  );


  buf

  (
    G1913_o2_p,
    G1913_o2
  );


  not

  (
    G1913_o2_n,
    G1913_o2
  );


  buf

  (
    G1929_o2_p,
    G1929_o2
  );


  not

  (
    G1929_o2_n,
    G1929_o2
  );


  buf

  (
    G1937_o2_p,
    G1937_o2
  );


  not

  (
    G1937_o2_n,
    G1937_o2
  );


  buf

  (
    G1945_o2_p,
    G1945_o2
  );


  not

  (
    G1945_o2_n,
    G1945_o2
  );


  buf

  (
    G1953_o2_p,
    G1953_o2
  );


  not

  (
    G1953_o2_n,
    G1953_o2
  );


  buf

  (
    G1843_o2_p,
    G1843_o2
  );


  not

  (
    G1843_o2_n,
    G1843_o2
  );


  buf

  (
    G1859_o2_p,
    G1859_o2
  );


  not

  (
    G1859_o2_n,
    G1859_o2
  );


  buf

  (
    G1867_o2_p,
    G1867_o2
  );


  not

  (
    G1867_o2_n,
    G1867_o2
  );


  buf

  (
    G1875_o2_p,
    G1875_o2
  );


  not

  (
    G1875_o2_n,
    G1875_o2
  );


  buf

  (
    G1883_o2_p,
    G1883_o2
  );


  not

  (
    G1883_o2_n,
    G1883_o2
  );


  buf

  (
    G1907_o2_p,
    G1907_o2
  );


  not

  (
    G1907_o2_n,
    G1907_o2
  );


  buf

  (
    G1923_o2_p,
    G1923_o2
  );


  not

  (
    G1923_o2_n,
    G1923_o2
  );


  buf

  (
    G1931_o2_p,
    G1931_o2
  );


  not

  (
    G1931_o2_n,
    G1931_o2
  );


  buf

  (
    G1939_o2_p,
    G1939_o2
  );


  not

  (
    G1939_o2_n,
    G1939_o2
  );


  buf

  (
    G1947_o2_p,
    G1947_o2
  );


  not

  (
    G1947_o2_n,
    G1947_o2
  );


  buf

  (
    G1844_o2_p,
    G1844_o2
  );


  not

  (
    G1844_o2_n,
    G1844_o2
  );


  buf

  (
    G1860_o2_p,
    G1860_o2
  );


  not

  (
    G1860_o2_n,
    G1860_o2
  );


  buf

  (
    G1868_o2_p,
    G1868_o2
  );


  not

  (
    G1868_o2_n,
    G1868_o2
  );


  buf

  (
    G1876_o2_p,
    G1876_o2
  );


  not

  (
    G1876_o2_n,
    G1876_o2
  );


  buf

  (
    G1884_o2_p,
    G1884_o2
  );


  not

  (
    G1884_o2_n,
    G1884_o2
  );


  buf

  (
    G1908_o2_p,
    G1908_o2
  );


  not

  (
    G1908_o2_n,
    G1908_o2
  );


  buf

  (
    G1924_o2_p,
    G1924_o2
  );


  not

  (
    G1924_o2_n,
    G1924_o2
  );


  buf

  (
    G1932_o2_p,
    G1932_o2
  );


  not

  (
    G1932_o2_n,
    G1932_o2
  );


  buf

  (
    G1940_o2_p,
    G1940_o2
  );


  not

  (
    G1940_o2_n,
    G1940_o2
  );


  buf

  (
    G1948_o2_p,
    G1948_o2
  );


  not

  (
    G1948_o2_n,
    G1948_o2
  );


  buf

  (
    G1847_o2_p,
    G1847_o2
  );


  not

  (
    G1847_o2_n,
    G1847_o2
  );


  buf

  (
    G1863_o2_p,
    G1863_o2
  );


  not

  (
    G1863_o2_n,
    G1863_o2
  );


  buf

  (
    G1871_o2_p,
    G1871_o2
  );


  not

  (
    G1871_o2_n,
    G1871_o2
  );


  buf

  (
    G1879_o2_p,
    G1879_o2
  );


  not

  (
    G1879_o2_n,
    G1879_o2
  );


  buf

  (
    G1887_o2_p,
    G1887_o2
  );


  not

  (
    G1887_o2_n,
    G1887_o2
  );


  buf

  (
    G1911_o2_p,
    G1911_o2
  );


  not

  (
    G1911_o2_n,
    G1911_o2
  );


  buf

  (
    G1927_o2_p,
    G1927_o2
  );


  not

  (
    G1927_o2_n,
    G1927_o2
  );


  buf

  (
    G1935_o2_p,
    G1935_o2
  );


  not

  (
    G1935_o2_n,
    G1935_o2
  );


  buf

  (
    G1943_o2_p,
    G1943_o2
  );


  not

  (
    G1943_o2_n,
    G1943_o2
  );


  buf

  (
    G1951_o2_p,
    G1951_o2
  );


  not

  (
    G1951_o2_n,
    G1951_o2
  );


  buf

  (
    G2444_o2_p,
    G2444_o2
  );


  not

  (
    G2444_o2_n,
    G2444_o2
  );


  buf

  (
    G2451_o2_p,
    G2451_o2
  );


  not

  (
    G2451_o2_n,
    G2451_o2
  );


  buf

  (
    G2502_o2_p,
    G2502_o2
  );


  not

  (
    G2502_o2_n,
    G2502_o2
  );


  buf

  (
    G2507_o2_p,
    G2507_o2
  );


  not

  (
    G2507_o2_n,
    G2507_o2
  );


  buf

  (
    n1464_inv_p,
    n1464_inv
  );


  not

  (
    n1464_inv_n,
    n1464_inv
  );


  buf

  (
    G2583_o2_p,
    G2583_o2
  );


  not

  (
    G2583_o2_n,
    G2583_o2
  );


  buf

  (
    n1797_lo_buf_o2_p,
    n1797_lo_buf_o2
  );


  not

  (
    n1797_lo_buf_o2_n,
    n1797_lo_buf_o2
  );


  buf

  (
    n1833_lo_buf_o2_p,
    n1833_lo_buf_o2
  );


  not

  (
    n1833_lo_buf_o2_n,
    n1833_lo_buf_o2
  );


  buf

  (
    n1881_lo_buf_o2_p,
    n1881_lo_buf_o2
  );


  not

  (
    n1881_lo_buf_o2_n,
    n1881_lo_buf_o2
  );


  buf

  (
    n1479_inv_p,
    n1479_inv
  );


  not

  (
    n1479_inv_n,
    n1479_inv
  );


  buf

  (
    n1482_inv_p,
    n1482_inv
  );


  not

  (
    n1482_inv_n,
    n1482_inv
  );


  buf

  (
    n1485_inv_p,
    n1485_inv
  );


  not

  (
    n1485_inv_n,
    n1485_inv
  );


  buf

  (
    G615_o2_p,
    G615_o2
  );


  not

  (
    G615_o2_n,
    G615_o2
  );


  buf

  (
    G2254_o2_p,
    G2254_o2
  );


  not

  (
    G2254_o2_n,
    G2254_o2
  );


  buf

  (
    G2255_o2_p,
    G2255_o2
  );


  not

  (
    G2255_o2_n,
    G2255_o2
  );


  buf

  (
    G2027_o2_p,
    G2027_o2
  );


  not

  (
    G2027_o2_n,
    G2027_o2
  );


  buf

  (
    G2393_o2_p,
    G2393_o2
  );


  not

  (
    G2393_o2_n,
    G2393_o2
  );


  buf

  (
    G527_o2_p,
    G527_o2
  );


  not

  (
    G527_o2_n,
    G527_o2
  );


  buf

  (
    G594_o2_p,
    G594_o2
  );


  not

  (
    G594_o2_n,
    G594_o2
  );


  buf

  (
    G1689_o2_p,
    G1689_o2
  );


  not

  (
    G1689_o2_n,
    G1689_o2
  );


  buf

  (
    G1693_o2_p,
    G1693_o2
  );


  not

  (
    G1693_o2_n,
    G1693_o2
  );


  buf

  (
    G2281_o2_p,
    G2281_o2
  );


  not

  (
    G2281_o2_n,
    G2281_o2
  );


  buf

  (
    G2014_o2_p,
    G2014_o2
  );


  not

  (
    G2014_o2_n,
    G2014_o2
  );


  buf

  (
    G2459_o2_p,
    G2459_o2
  );


  not

  (
    G2459_o2_n,
    G2459_o2
  );


  buf

  (
    G2561_o2_p,
    G2561_o2
  );


  not

  (
    G2561_o2_n,
    G2561_o2
  );


  buf

  (
    G2533_o2_p,
    G2533_o2
  );


  not

  (
    G2533_o2_n,
    G2533_o2
  );


  buf

  (
    n1749_lo_buf_o2_p,
    n1749_lo_buf_o2
  );


  not

  (
    n1749_lo_buf_o2_n,
    n1749_lo_buf_o2
  );


  buf

  (
    n1761_lo_buf_o2_p,
    n1761_lo_buf_o2
  );


  not

  (
    n1761_lo_buf_o2_n,
    n1761_lo_buf_o2
  );


  buf

  (
    n1773_lo_buf_o2_p,
    n1773_lo_buf_o2
  );


  not

  (
    n1773_lo_buf_o2_n,
    n1773_lo_buf_o2
  );


  buf

  (
    n1809_lo_buf_o2_p,
    n1809_lo_buf_o2
  );


  not

  (
    n1809_lo_buf_o2_n,
    n1809_lo_buf_o2
  );


  buf

  (
    G1955_o2_p,
    G1955_o2
  );


  not

  (
    G1955_o2_n,
    G1955_o2
  );


  buf

  (
    G1958_o2_p,
    G1958_o2
  );


  not

  (
    G1958_o2_n,
    G1958_o2
  );


  buf

  (
    G2562_o2_p,
    G2562_o2
  );


  not

  (
    G2562_o2_n,
    G2562_o2
  );


  buf

  (
    G2398_o2_p,
    G2398_o2
  );


  not

  (
    G2398_o2_n,
    G2398_o2
  );


  buf

  (
    n1554_inv_p,
    n1554_inv
  );


  not

  (
    n1554_inv_n,
    n1554_inv
  );


  buf

  (
    n1557_inv_p,
    n1557_inv
  );


  not

  (
    n1557_inv_n,
    n1557_inv
  );


  buf

  (
    G2577_o2_p,
    G2577_o2
  );


  not

  (
    G2577_o2_n,
    G2577_o2
  );


  buf

  (
    G2627_o2_p,
    G2627_o2
  );


  not

  (
    G2627_o2_n,
    G2627_o2
  );


  buf

  (
    G654_o2_p,
    G654_o2
  );


  not

  (
    G654_o2_n,
    G654_o2
  );


  buf

  (
    G660_o2_p,
    G660_o2
  );


  not

  (
    G660_o2_n,
    G660_o2
  );


  buf

  (
    G831_o2_p,
    G831_o2
  );


  not

  (
    G831_o2_n,
    G831_o2
  );


  buf

  (
    G919_o2_p,
    G919_o2
  );


  not

  (
    G919_o2_n,
    G919_o2
  );


  buf

  (
    G925_o2_p,
    G925_o2
  );


  not

  (
    G925_o2_n,
    G925_o2
  );


  buf

  (
    n1815_lo_buf_o2_p,
    n1815_lo_buf_o2
  );


  not

  (
    n1815_lo_buf_o2_n,
    n1815_lo_buf_o2
  );


  buf

  (
    n1899_lo_buf_o2_p,
    n1899_lo_buf_o2
  );


  not

  (
    n1899_lo_buf_o2_n,
    n1899_lo_buf_o2
  );


  buf

  (
    n2079_lo_buf_o2_p,
    n2079_lo_buf_o2
  );


  not

  (
    n2079_lo_buf_o2_n,
    n2079_lo_buf_o2
  );


  buf

  (
    n2127_lo_buf_o2_p,
    n2127_lo_buf_o2
  );


  not

  (
    n2127_lo_buf_o2_n,
    n2127_lo_buf_o2
  );


  buf

  (
    n2139_lo_buf_o2_p,
    n2139_lo_buf_o2
  );


  not

  (
    n2139_lo_buf_o2_n,
    n2139_lo_buf_o2
  );


  buf

  (
    n2151_lo_buf_o2_p,
    n2151_lo_buf_o2
  );


  not

  (
    n2151_lo_buf_o2_n,
    n2151_lo_buf_o2
  );


  buf

  (
    n2187_lo_buf_o2_p,
    n2187_lo_buf_o2
  );


  not

  (
    n2187_lo_buf_o2_n,
    n2187_lo_buf_o2
  );


  buf

  (
    n2199_lo_buf_o2_p,
    n2199_lo_buf_o2
  );


  not

  (
    n2199_lo_buf_o2_n,
    n2199_lo_buf_o2
  );


  buf

  (
    n2211_lo_buf_o2_p,
    n2211_lo_buf_o2
  );


  not

  (
    n2211_lo_buf_o2_n,
    n2211_lo_buf_o2
  );


  buf

  (
    G533_o2_p,
    G533_o2
  );


  not

  (
    G533_o2_n,
    G533_o2
  );


  buf

  (
    n1854_lo_buf_o2_p,
    n1854_lo_buf_o2
  );


  not

  (
    n1854_lo_buf_o2_n,
    n1854_lo_buf_o2
  );


  buf

  (
    n2094_lo_buf_o2_p,
    n2094_lo_buf_o2
  );


  not

  (
    n2094_lo_buf_o2_n,
    n2094_lo_buf_o2
  );


  buf

  (
    G667_o2_p,
    G667_o2
  );


  not

  (
    G667_o2_n,
    G667_o2
  );


  buf

  (
    G874_o2_p,
    G874_o2
  );


  not

  (
    G874_o2_n,
    G874_o2
  );


  buf

  (
    G851_o2_p,
    G851_o2
  );


  not

  (
    G851_o2_n,
    G851_o2
  );


  buf

  (
    G1127_o2_p,
    G1127_o2
  );


  not

  (
    G1127_o2_n,
    G1127_o2
  );


  buf

  (
    n1869_lo_buf_o2_p,
    n1869_lo_buf_o2
  );


  not

  (
    n1869_lo_buf_o2_n,
    n1869_lo_buf_o2
  );


  buf

  (
    n2109_lo_buf_o2_p,
    n2109_lo_buf_o2
  );


  not

  (
    n2109_lo_buf_o2_n,
    n2109_lo_buf_o2
  );


  buf

  (
    n2121_lo_buf_o2_p,
    n2121_lo_buf_o2
  );


  not

  (
    n2121_lo_buf_o2_n,
    n2121_lo_buf_o2
  );


  buf

  (
    G477_o2_p,
    G477_o2
  );


  not

  (
    G477_o2_n,
    G477_o2
  );


  buf

  (
    G491_o2_p,
    G491_o2
  );


  not

  (
    G491_o2_n,
    G491_o2
  );


  buf

  (
    G501_o2_p,
    G501_o2
  );


  not

  (
    G501_o2_n,
    G501_o2
  );


  buf

  (
    G786_o2_p,
    G786_o2
  );


  not

  (
    G786_o2_n,
    G786_o2
  );


  buf

  (
    G791_o2_p,
    G791_o2
  );


  not

  (
    G791_o2_n,
    G791_o2
  );


  buf

  (
    G1126_o2_p,
    G1126_o2
  );


  not

  (
    G1126_o2_n,
    G1126_o2
  );


  buf

  (
    G1052_o2_p,
    G1052_o2
  );


  not

  (
    G1052_o2_n,
    G1052_o2
  );


  buf

  (
    G1054_o2_p,
    G1054_o2
  );


  not

  (
    G1054_o2_n,
    G1054_o2
  );


  and

  (
    g580_p,
    n3968_o2_n,
    n3980_o2_n
  );


  and

  (
    g581_p,
    g580_p,
    n3610_o2_n
  );


  and

  (
    g582_p,
    g581_p,
    n4413_o2_n
  );


  or

  (
    g583_n,
    G727_o2_n,
    n1872_lo_n
  );


  and

  (
    g584_p,
    G742_o2_p,
    n5011_o2_n_spl_
  );


  or

  (
    g584_n,
    G742_o2_n,
    n5011_o2_p_spl_
  );


  and

  (
    g585_p,
    g584_p,
    n5013_o2_n_spl_
  );


  or

  (
    g585_n,
    g584_n,
    n5013_o2_p_spl_
  );


  or

  (
    g586_n,
    g585_n_spl_,
    n5156_o2_n
  );


  and

  (
    g587_p,
    n2172_lo_n_spl_,
    n2160_lo_n_spl_
  );


  or

  (
    g588_n,
    g587_p,
    n2148_lo_n_spl_
  );


  and

  (
    g589_p,
    n5012_o2_n,
    n5011_o2_n_spl_
  );


  or

  (
    g589_n,
    n5012_o2_p,
    n5011_o2_p_spl_
  );


  and

  (
    g590_p,
    g589_p_spl_,
    n5013_o2_n_spl_
  );


  or

  (
    g590_n,
    g589_n_spl_,
    n5013_o2_p_spl_
  );


  or

  (
    g591_n,
    g590_n,
    g588_n
  );


  or

  (
    g592_n,
    n5014_o2_p,
    n2100_lo_n
  );


  or

  (
    g593_n,
    n5117_o2_p,
    n2112_lo_n
  );


  or

  (
    g594_n,
    n5115_o2_p,
    n2124_lo_n
  );


  or

  (
    g595_n,
    n5122_o2_p,
    n2136_lo_n
  );


  and

  (
    g596_p,
    g593_n,
    g592_n
  );


  and

  (
    g597_p,
    g596_p,
    g594_n
  );


  and

  (
    g598_p,
    g597_p,
    g595_n
  );


  or

  (
    g599_n,
    n5121_o2_p,
    n2148_lo_n_spl_
  );


  or

  (
    g600_n,
    n5119_o2_p,
    n2160_lo_n_spl_
  );


  or

  (
    g601_n,
    n5116_o2_p,
    n2172_lo_n_spl_
  );


  or

  (
    g602_n,
    n5123_o2_p,
    n2184_lo_n
  );


  and

  (
    g603_p,
    g600_n,
    g599_n
  );


  and

  (
    g604_p,
    g603_p,
    g601_n
  );


  and

  (
    g605_p,
    g604_p,
    g602_n
  );


  and

  (
    g606_p,
    g605_p,
    g598_p
  );


  or

  (
    g607_n,
    g590_p,
    g585_p_spl_
  );


  or

  (
    g608_n,
    g607_n,
    g606_p
  );


  and

  (
    g609_p,
    g591_n,
    g586_n
  );


  and

  (
    g610_p,
    g609_p,
    g608_n
  );


  and

  (
    g611_p,
    n4634_o2_n_spl_,
    n4633_o2_p_spl_
  );


  or

  (
    g611_n,
    n4634_o2_p_spl_,
    n4633_o2_n_spl_
  );


  and

  (
    g612_p,
    n4634_o2_p_spl_,
    n4633_o2_n_spl_
  );


  or

  (
    g612_n,
    n4634_o2_n_spl_,
    n4633_o2_p_spl_
  );


  and

  (
    g613_p,
    g612_n,
    g611_n
  );


  or

  (
    g613_n,
    g612_p,
    g611_p
  );


  or

  (
    g614_n,
    g613_p,
    G1514_o2_n
  );


  or

  (
    g615_n,
    g613_n,
    G1514_o2_p
  );


  and

  (
    g616_p,
    g615_n,
    g614_n
  );


  and

  (
    g617_p,
    G1823_o2_p,
    n5167_o2_n
  );


  and

  (
    g618_p,
    G1823_o2_n,
    n5167_o2_p
  );


  or

  (
    g619_n,
    g618_p,
    g617_p
  );


  and

  (
    g620_p,
    n4418_o2_p_spl_,
    n4371_o2_p
  );


  and

  (
    g621_p,
    n4418_o2_p_spl_,
    n4298_o2_p
  );


  or

  (
    g622_n,
    g621_p,
    n4628_o2_p
  );


  and

  (
    g623_p,
    n4890_o2_p,
    n2304_lo_p_spl_
  );


  and

  (
    g624_p,
    g623_p,
    n4629_o2_n
  );


  and

  (
    g625_p,
    G1048_o2_n,
    n5156_o2_p
  );


  or

  (
    g626_n,
    n5016_o2_p,
    n5021_o2_p
  );


  and

  (
    g627_p,
    g626_n,
    G572_o2_n
  );


  and

  (
    g628_p,
    G1048_o2_p,
    G572_o2_p
  );


  and

  (
    g629_p,
    g628_p,
    n5026_o2_n
  );


  or

  (
    g630_n,
    g627_p,
    g625_p
  );


  or

  (
    g631_n,
    g630_n,
    g629_p
  );


  or

  (
    g632_n,
    G3045_o2_n,
    G3042_o2_p
  );


  or

  (
    g633_n,
    g632_n,
    G2851_o2_p
  );


  and

  (
    g634_p,
    g633_n_spl_,
    G3100_o2_n
  );


  or

  (
    g635_n,
    G3143_o2_p,
    G3140_o2_p
  );


  or

  (
    g636_n,
    g635_n,
    G2842_o2_p
  );


  and

  (
    g637_p,
    g636_n_spl_,
    G3195_o2_p
  );


  and

  (
    g638_p,
    n3241_o2_p,
    n1836_lo_p
  );


  and

  (
    g639_p,
    n3241_o2_n,
    n1836_lo_n
  );


  or

  (
    g640_n,
    g639_p,
    g638_p
  );


  and

  (
    g641_p,
    g640_n,
    n4886_o2_n
  );


  and

  (
    g642_p,
    g641_p,
    n5015_o2_n
  );


  and

  (
    g643_p,
    n5015_o2_p,
    n4884_o2_n
  );


  or

  (
    g644_n,
    g643_p,
    g642_p
  );


  and

  (
    g645_p,
    g644_n,
    g589_p_spl_
  );


  and

  (
    g646_p,
    n3242_o2_p,
    n1884_lo_p
  );


  and

  (
    g647_p,
    n3242_o2_n,
    n1884_lo_n
  );


  or

  (
    g648_n,
    g647_p,
    g646_p
  );


  and

  (
    g649_p,
    g648_n,
    n5123_o2_n
  );


  and

  (
    g650_p,
    g649_p,
    g585_p_spl_
  );


  and

  (
    g651_p,
    G2991_o2_n_spl_,
    G2887_o2_p_spl_
  );


  or

  (
    g651_n,
    G2991_o2_p_spl_,
    G2887_o2_n_spl_
  );


  and

  (
    g652_p,
    G2991_o2_p_spl_,
    G2887_o2_n_spl_
  );


  or

  (
    g652_n,
    G2991_o2_n_spl_,
    G2887_o2_p_spl_
  );


  and

  (
    g653_p,
    g652_n,
    g651_n
  );


  or

  (
    g653_n,
    g652_p,
    g651_p
  );


  and

  (
    g654_p,
    g653_n,
    n2304_lo_p_spl_
  );


  or

  (
    g654_n,
    g653_p,
    n2304_lo_n
  );


  and

  (
    g655_p,
    n4733_o2_p_spl_,
    n4732_o2_p_spl_
  );


  or

  (
    g655_n,
    n4733_o2_n_spl_,
    n4732_o2_n_spl_
  );


  and

  (
    g656_p,
    n4733_o2_n_spl_,
    n4732_o2_n_spl_
  );


  or

  (
    g656_n,
    n4733_o2_p_spl_,
    n4732_o2_p_spl_
  );


  and

  (
    g657_p,
    g656_n,
    g655_n
  );


  or

  (
    g657_n,
    g656_p,
    g655_p
  );


  and

  (
    g658_p,
    g657_p,
    g654_p
  );


  and

  (
    g659_p,
    g657_n,
    g654_n
  );


  or

  (
    g660_n,
    g659_p,
    g658_p
  );


  and

  (
    g661_p,
    g589_n_spl_,
    g585_n_spl_
  );


  and

  (
    g662_p,
    g661_p,
    g660_n
  );


  or

  (
    g663_n,
    g650_p,
    g645_p
  );


  or

  (
    g664_n,
    g663_n,
    g662_p
  );


  or

  (
    g665_n,
    G3251_o2_p,
    G3220_o2_p
  );


  or

  (
    g666_n,
    g665_n,
    G2845_o2_p
  );


  and

  (
    g667_p,
    g666_n_spl_,
    G3275_o2_p
  );


  or

  (
    g668_n,
    G3254_o2_p,
    G3146_o2_p
  );


  or

  (
    g669_n,
    g668_n,
    G2848_o2_p
  );


  and

  (
    g670_p,
    g669_n_spl_,
    G3281_o2_p
  );


  or

  (
    g671_n,
    G3262_o2_p,
    G3174_o2_p
  );


  or

  (
    g672_n,
    g671_n,
    G2929_o2_p
  );


  and

  (
    g673_p,
    g672_n_spl_,
    G3294_o2_p
  );


  or

  (
    g674_n,
    G3291_o2_p,
    G3217_o2_p
  );


  or

  (
    g675_n,
    g674_n,
    G2839_o2_p
  );


  and

  (
    g676_p,
    g675_n_spl_,
    G3320_o2_p
  );


  or

  (
    g677_n,
    g669_n_spl_,
    g633_n_spl_
  );


  or

  (
    g678_n,
    g677_n,
    g672_n_spl_
  );


  or

  (
    g679_n,
    g678_n,
    g666_n_spl_
  );


  or

  (
    g680_n,
    G3288_o2_p,
    G3171_o2_p
  );


  or

  (
    g681_n,
    g680_n,
    G2926_o2_p
  );


  or

  (
    g682_n,
    G3302_o2_p,
    G3272_o2_p
  );


  or

  (
    g683_n,
    g682_n,
    G2836_o2_p
  );


  or

  (
    g684_n,
    g675_n_spl_,
    g636_n_spl_
  );


  or

  (
    g685_n,
    g684_n,
    g681_n_spl_
  );


  or

  (
    g686_n,
    g685_n,
    g683_n_spl_
  );


  or

  (
    g687_n,
    g686_n,
    g679_n
  );


  and

  (
    g688_p,
    G621_o2_p,
    G618_o2_p
  );


  or

  (
    g688_n,
    G621_o2_n,
    G618_o2_n
  );


  or

  (
    g689_n,
    g683_n_spl_,
    g681_n_spl_
  );


  or

  (
    g690_n,
    g689_n,
    g688_n_spl_
  );


  and

  (
    g691_p,
    g690_n,
    g687_n_spl_
  );


  and

  (
    g692_p,
    g691_p,
    n2064_lo_p
  );


  and

  (
    g693_p,
    G3359_o2_n,
    G3346_o2_n
  );


  or

  (
    g693_n,
    G3359_o2_p,
    G3346_o2_p
  );


  and

  (
    g694_p,
    G3344_o2_n,
    G3340_o2_p
  );


  or

  (
    g694_n,
    G3344_o2_p,
    G3340_o2_n
  );


  and

  (
    g695_p,
    g694_n_spl_,
    g693_p_spl_
  );


  or

  (
    g695_n,
    g694_p_spl_,
    g693_n_spl_
  );


  and

  (
    g696_p,
    g694_p_spl_,
    g693_n_spl_
  );


  or

  (
    g696_n,
    g694_n_spl_,
    g693_p_spl_
  );


  and

  (
    g697_p,
    g696_n,
    g695_n
  );


  or

  (
    g697_n,
    g696_p,
    g695_p
  );


  and

  (
    g698_p,
    G3265_o2_p,
    G3373_o2_p
  );


  or

  (
    g698_n,
    G3265_o2_n,
    G3373_o2_n
  );


  and

  (
    g699_p,
    G3404_o2_n,
    G3237_o2_n
  );


  or

  (
    g699_n,
    G3404_o2_p,
    G3237_o2_p
  );


  and

  (
    g700_p,
    g699_n,
    g698_n
  );


  or

  (
    g700_n,
    g699_p,
    g698_p
  );


  and

  (
    g701_p,
    G3360_o2_p_spl_,
    G3350_o2_n_spl_
  );


  or

  (
    g701_n,
    G3360_o2_n_spl_,
    G3350_o2_p_spl_
  );


  and

  (
    g702_p,
    G3360_o2_n_spl_,
    G3350_o2_p_spl_
  );


  or

  (
    g702_n,
    G3360_o2_p_spl_,
    G3350_o2_n_spl_
  );


  and

  (
    g703_p,
    g702_n,
    g701_n
  );


  or

  (
    g703_n,
    g702_p,
    g701_p
  );


  and

  (
    g704_p,
    g688_n_spl_,
    n2340_lo_p
  );


  or

  (
    g704_n,
    g688_p,
    n2340_lo_n
  );


  and

  (
    g705_p,
    g703_n_spl_,
    g700_n_spl_0
  );


  or

  (
    g705_n,
    g703_p_spl_,
    g700_p_spl_0
  );


  and

  (
    g706_p,
    g705_p,
    g704_p_spl_0
  );


  or

  (
    g706_n,
    g705_n,
    g704_n_spl_0
  );


  and

  (
    g707_p,
    G3399_o2_p_spl_,
    G3383_o2_n_spl_
  );


  or

  (
    g707_n,
    G3399_o2_n_spl_,
    G3383_o2_p_spl_
  );


  and

  (
    g708_p,
    G3399_o2_n_spl_,
    G3383_o2_p_spl_
  );


  or

  (
    g708_n,
    G3399_o2_p_spl_,
    G3383_o2_n_spl_
  );


  and

  (
    g709_p,
    g708_n,
    g707_n
  );


  or

  (
    g709_n,
    g708_p,
    g707_p
  );


  and

  (
    g710_p,
    g709_p_spl_,
    g700_n_spl_0
  );


  or

  (
    g710_n,
    g709_n_spl_,
    g700_p_spl_0
  );


  and

  (
    g711_p,
    g710_p,
    g704_n_spl_0
  );


  or

  (
    g711_n,
    g710_n,
    g704_p_spl_0
  );


  and

  (
    g712_p,
    G3240_o2_p_spl_,
    G3376_o2_p_spl_
  );


  or

  (
    g712_n,
    G3240_o2_n_spl_,
    G3376_o2_n_spl_
  );


  and

  (
    g713_p,
    G3240_o2_n_spl_,
    G3376_o2_n_spl_
  );


  or

  (
    g713_n,
    G3240_o2_p_spl_,
    G3376_o2_p_spl_
  );


  and

  (
    g714_p,
    g713_n,
    g712_n
  );


  or

  (
    g714_n,
    g713_p,
    g712_p
  );


  and

  (
    g715_p,
    g714_p_spl_,
    g703_n_spl_
  );


  or

  (
    g715_n,
    g714_n_spl_,
    g703_p_spl_
  );


  and

  (
    g716_p,
    g715_p,
    g704_n_spl_1
  );


  or

  (
    g716_n,
    g715_n,
    g704_p_spl_1
  );


  and

  (
    g717_p,
    g714_p_spl_,
    g709_p_spl_
  );


  or

  (
    g717_n,
    g714_n_spl_,
    g709_n_spl_
  );


  and

  (
    g718_p,
    g717_p,
    g704_p_spl_1
  );


  or

  (
    g718_n,
    g717_n,
    g704_n_spl_1
  );


  and

  (
    g719_p,
    g711_n,
    g706_n
  );


  or

  (
    g719_n,
    g711_p,
    g706_p
  );


  and

  (
    g720_p,
    g719_p,
    g716_n
  );


  or

  (
    g720_n,
    g719_n,
    g716_p
  );


  and

  (
    g721_p,
    g720_p,
    g718_n
  );


  or

  (
    g721_n,
    g720_n,
    g718_p
  );


  and

  (
    g722_p,
    g721_n,
    g697_n_spl_
  );


  and

  (
    g723_p,
    g721_p,
    g697_p_spl_
  );


  or

  (
    g724_n,
    g723_p,
    g722_p
  );


  and

  (
    g725_p,
    G3367_o2_n_spl_,
    G3353_o2_p_spl_
  );


  or

  (
    g725_n,
    G3367_o2_p_spl_,
    G3353_o2_n_spl_
  );


  and

  (
    g726_p,
    G3367_o2_p_spl_,
    G3353_o2_n_spl_
  );


  or

  (
    g726_n,
    G3367_o2_n_spl_,
    G3353_o2_p_spl_
  );


  and

  (
    g727_p,
    g726_n,
    g725_n
  );


  or

  (
    g727_n,
    g726_p,
    g725_p
  );


  and

  (
    g728_p,
    g727_n_spl_,
    g700_n_spl_1
  );


  or

  (
    g728_n,
    g727_p_spl_,
    g700_p_spl_1
  );


  and

  (
    g729_p,
    g727_p_spl_,
    g700_p_spl_1
  );


  or

  (
    g729_n,
    g727_n_spl_,
    g700_n_spl_1
  );


  and

  (
    g730_p,
    g729_n,
    g728_n
  );


  or

  (
    g730_n,
    g729_p,
    g728_p
  );


  or

  (
    g731_n,
    g730_n,
    g697_p_spl_
  );


  or

  (
    g732_n,
    g730_p,
    g697_n_spl_
  );


  and

  (
    g733_p,
    g732_n,
    g731_n
  );


  or

  (
    g734_n,
    G434_o2_p_spl_,
    G447_o2_p
  );


  and

  (
    g735_p,
    G1311_o2_n,
    G1203_o2_p
  );


  and

  (
    g736_p,
    G1312_o2_n,
    G1200_o2_p
  );


  or

  (
    g737_n,
    g736_p,
    g735_p
  );


  or

  (
    g738_n,
    G1519_o2_p,
    G1463_o2_n
  );


  or

  (
    g739_n,
    G1520_o2_p,
    G1460_o2_n
  );


  and

  (
    g740_p,
    g739_n,
    g738_n
  );


  and

  (
    g741_p,
    n852_inv_n_spl_0,
    n849_inv_n_spl_
  );


  or

  (
    g741_n,
    n852_inv_p_spl_0,
    n849_inv_p_spl_0
  );


  and

  (
    g742_p,
    g741_p,
    n855_inv_n
  );


  or

  (
    g742_n,
    g741_n,
    n855_inv_p_spl_
  );


  and

  (
    g743_p,
    g742_p,
    n4539_o2_p_spl_0
  );


  or

  (
    g743_n,
    g742_n,
    n4539_o2_n_spl_0
  );


  and

  (
    g744_p,
    G2533_o2_n,
    G2459_o2_n
  );


  or

  (
    g744_n,
    G2533_o2_p,
    G2459_o2_p
  );


  and

  (
    g745_p,
    g744_p,
    G2561_o2_n
  );


  or

  (
    g745_n,
    g744_n,
    G2561_o2_p
  );


  and

  (
    g746_p,
    g745_p,
    G2562_o2_n
  );


  or

  (
    g746_n,
    g745_n,
    G2562_o2_p
  );


  and

  (
    g747_p,
    G3063_o2_n,
    G2939_o2_p
  );


  or

  (
    g747_n,
    G3063_o2_p,
    G2939_o2_n
  );


  and

  (
    g748_p,
    G2980_o2_n,
    G3027_o2_p
  );


  or

  (
    g748_n,
    G2980_o2_p,
    G3027_o2_n
  );


  and

  (
    g749_p,
    g748_n,
    g747_n
  );


  or

  (
    g749_n,
    g748_p,
    g747_p
  );


  and

  (
    g750_p,
    n4816_o2_n_spl_,
    n429_inv_n_spl_
  );


  or

  (
    g750_n,
    n4816_o2_p_spl_,
    n429_inv_p_spl_0
  );


  and

  (
    g751_p,
    g750_p,
    n4401_o2_p
  );


  or

  (
    g751_n,
    g750_n,
    n4401_o2_n
  );


  and

  (
    g752_p,
    g751_n,
    n4398_o2_n
  );


  or

  (
    g752_n,
    g751_p,
    n4398_o2_p_spl_
  );


  and

  (
    g753_p,
    g752_n_spl_0,
    g749_n_spl_
  );


  and

  (
    g754_p,
    G3035_o2_n,
    G2866_o2_n
  );


  or

  (
    g754_n,
    G3035_o2_p,
    G2866_o2_p
  );


  and

  (
    g755_p,
    G2916_o2_p,
    G2999_o2_p
  );


  or

  (
    g755_n,
    G2916_o2_n,
    G2999_o2_n
  );


  and

  (
    g756_p,
    g755_n,
    g754_n
  );


  or

  (
    g756_n,
    g755_p,
    g754_p
  );


  or

  (
    g757_n,
    g756_p_spl_0,
    g752_p_spl_00
  );


  and

  (
    g758_p,
    G3069_o2_n_spl_,
    G2962_o2_n_spl_
  );


  or

  (
    g758_n,
    G3069_o2_p_spl_,
    G2962_o2_p_spl_
  );


  and

  (
    g759_p,
    G3069_o2_p_spl_,
    G2962_o2_p_spl_
  );


  or

  (
    g759_n,
    G3069_o2_n_spl_,
    G2962_o2_n_spl_
  );


  and

  (
    g760_p,
    g759_n,
    g758_n
  );


  or

  (
    g760_n,
    g759_p,
    g758_p
  );


  or

  (
    g761_n,
    g760_p_spl_0,
    g752_p_spl_00
  );


  or

  (
    g762_n,
    G3012_o2_n,
    G2880_o2_p
  );


  or

  (
    g763_n,
    G3012_o2_p,
    G2880_o2_n
  );


  and

  (
    g764_p,
    g763_n,
    g762_n
  );


  or

  (
    g765_n,
    g764_p_spl_,
    g752_p_spl_01
  );


  or

  (
    g766_n,
    G1843_o2_p,
    n1941_lo_buf_o2_n_spl_0
  );


  or

  (
    g767_n,
    G1844_o2_p,
    n1056_inv_p_spl_00
  );


  or

  (
    g768_n,
    G1845_o2_n,
    n858_inv_p_spl_00
  );


  or

  (
    g769_n,
    G1846_o2_p,
    n4651_o2_n_spl_00
  );


  or

  (
    g770_n,
    G1847_o2_p,
    n4919_o2_n_spl_00
  );


  or

  (
    g771_n,
    G1848_o2_p,
    n1977_lo_buf_o2_n_spl_00
  );


  or

  (
    g772_n,
    G1849_o2_n,
    n1965_lo_buf_o2_n_spl_00
  );


  or

  (
    g773_n,
    G1850_o2_p,
    n1953_lo_buf_o2_n_spl_0
  );


  and

  (
    g774_p,
    g767_n,
    g766_n
  );


  and

  (
    g775_p,
    g774_p,
    g768_n
  );


  and

  (
    g776_p,
    g775_p,
    g769_n
  );


  and

  (
    g777_p,
    g776_p,
    g770_n
  );


  and

  (
    g778_p,
    g777_p,
    g771_n
  );


  and

  (
    g779_p,
    g778_p,
    g772_n
  );


  and

  (
    g780_p,
    g779_p,
    g773_n
  );


  and

  (
    g781_p,
    g780_p,
    G519_o2_n_spl_000
  );


  or

  (
    g782_n,
    G1907_o2_p,
    n4653_o2_n_spl_0
  );


  or

  (
    g783_n,
    G1908_o2_p,
    n1071_inv_p_spl_00
  );


  or

  (
    g784_n,
    G1909_o2_n,
    n1068_inv_p_spl_00
  );


  or

  (
    g785_n,
    G1910_o2_p,
    n1062_inv_p_spl_00
  );


  or

  (
    g786_n,
    G1911_o2_p,
    n1053_inv_p_spl_00
  );


  or

  (
    g787_n,
    G1912_o2_p,
    n1074_inv_p_spl_00
  );


  or

  (
    g788_n,
    G1913_o2_n,
    n4571_o2_n_spl_00
  );


  or

  (
    g789_n,
    G1914_o2_p,
    n4572_o2_n_spl_00
  );


  and

  (
    g790_p,
    g783_n,
    g782_n
  );


  and

  (
    g791_p,
    g790_p,
    g784_n
  );


  and

  (
    g792_p,
    g791_p,
    g785_n
  );


  and

  (
    g793_p,
    g792_p,
    g786_n
  );


  and

  (
    g794_p,
    g793_p,
    g787_n
  );


  and

  (
    g795_p,
    g794_p,
    g788_n
  );


  and

  (
    g796_p,
    g795_p,
    g789_n
  );


  and

  (
    g797_p,
    g796_p,
    G519_o2_p_spl_000
  );


  or

  (
    g798_n,
    g797_p,
    g781_p
  );


  and

  (
    g799_p,
    G593_o2_p,
    n4783_o2_n
  );


  or

  (
    g799_n,
    G593_o2_n,
    n4783_o2_p
  );


  and

  (
    g800_p,
    n849_inv_n_spl_,
    n429_inv_p_spl_0
  );


  or

  (
    g800_n,
    n849_inv_p_spl_0,
    n429_inv_n_spl_
  );


  and

  (
    g801_p,
    g800_p,
    g799_n
  );


  or

  (
    g801_n,
    g800_n,
    g799_p
  );


  and

  (
    g802_p,
    g801_n_spl_00,
    g798_n
  );


  or

  (
    g803_n,
    G2580_o2_p,
    G2284_o2_p
  );


  or

  (
    g804_n,
    G2580_o2_n,
    G2284_o2_n
  );


  and

  (
    g805_p,
    g804_n,
    g803_n
  );


  and

  (
    g806_p,
    n852_inv_n_spl_0,
    n4389_o2_p_spl_0
  );


  or

  (
    g806_n,
    n852_inv_p_spl_0,
    n4389_o2_n_spl_0
  );


  and

  (
    g807_p,
    g806_p_spl_0,
    g805_p
  );


  and

  (
    g808_p,
    g806_n,
    g801_p_spl_0
  );


  and

  (
    g809_p,
    g808_p_spl_0,
    G384_o2_n
  );


  or

  (
    g810_n,
    g807_p,
    g802_p
  );


  or

  (
    g811_n,
    g810_n,
    g809_p
  );


  and

  (
    g812_p,
    g752_p_spl_01,
    g743_p_spl_00
  );


  or

  (
    g812_n,
    g752_n_spl_0,
    g743_n_spl_0
  );


  or

  (
    g813_n,
    g812_n_spl_00,
    g811_n
  );


  or

  (
    g814_n,
    G3078_o2_n,
    G2971_o2_p
  );


  or

  (
    g815_n,
    G3078_o2_p,
    G2971_o2_n
  );


  and

  (
    g816_p,
    g815_n,
    g814_n
  );


  or

  (
    g817_n,
    g816_p,
    G2923_o2_p_spl_0
  );


  or

  (
    g818_n,
    g756_p_spl_0,
    g749_p_spl_
  );


  or

  (
    g819_n,
    g818_n,
    g764_p_spl_
  );


  or

  (
    g820_n,
    g819_n,
    G2923_o2_n_spl_0
  );


  and

  (
    g821_p,
    g820_n,
    g817_n
  );


  or

  (
    g822_n,
    g821_p,
    g743_p_spl_00
  );


  and

  (
    g823_p,
    G2773_o2_p,
    n2301_lo_buf_o2_p_spl_0
  );


  and

  (
    g824_p,
    G2773_o2_n,
    n2301_lo_buf_o2_n_spl_
  );


  or

  (
    g825_n,
    g824_p,
    g823_p
  );


  and

  (
    g826_p,
    g825_n_spl_,
    g752_n_spl_
  );


  and

  (
    g827_p,
    g825_n_spl_,
    g743_n_spl_0
  );


  and

  (
    g828_p,
    g756_n,
    G2923_o2_n_spl_0
  );


  or

  (
    g828_n,
    g756_p_spl_,
    G2923_o2_p_spl_0
  );


  and

  (
    g829_p,
    g828_p,
    g749_n_spl_
  );


  and

  (
    g830_p,
    g828_n,
    g749_p_spl_
  );


  or

  (
    g831_n,
    g830_p,
    g829_p
  );


  and

  (
    g832_p,
    g831_n,
    g743_n_spl_
  );


  or

  (
    g833_n,
    G1859_o2_p,
    n1965_lo_buf_o2_n_spl_00
  );


  or

  (
    g834_n,
    G1860_o2_p,
    n1071_inv_p_spl_00
  );


  or

  (
    g835_n,
    G1861_o2_n,
    n1050_inv_p_spl_00
  );


  or

  (
    g836_n,
    G1862_o2_p,
    n1056_inv_p_spl_00
  );


  or

  (
    g837_n,
    G1863_o2_p,
    n858_inv_p_spl_00
  );


  or

  (
    g838_n,
    G1864_o2_p,
    n4651_o2_n_spl_00
  );


  or

  (
    g839_n,
    G1865_o2_n,
    n4919_o2_n_spl_00
  );


  or

  (
    g840_n,
    G1866_o2_p,
    n1977_lo_buf_o2_n_spl_00
  );


  and

  (
    g841_p,
    g834_n,
    g833_n
  );


  and

  (
    g842_p,
    g841_p,
    g835_n
  );


  and

  (
    g843_p,
    g842_p,
    g836_n
  );


  and

  (
    g844_p,
    g843_p,
    g837_n
  );


  and

  (
    g845_p,
    g844_p,
    g838_n
  );


  and

  (
    g846_p,
    g845_p,
    g839_n
  );


  and

  (
    g847_p,
    g846_p,
    g840_n
  );


  and

  (
    g848_p,
    g847_p,
    G519_o2_n_spl_000
  );


  or

  (
    g849_n,
    G1923_o2_p,
    n2253_lo_buf_o2_n_spl_
  );


  or

  (
    g850_n,
    G1924_o2_p,
    n1062_inv_p_spl_00
  );


  or

  (
    g851_n,
    G1925_o2_n,
    n1053_inv_p_spl_00
  );


  or

  (
    g852_n,
    G1926_o2_p,
    n1074_inv_p_spl_00
  );


  or

  (
    g853_n,
    G1927_o2_p,
    n4571_o2_n_spl_00
  );


  or

  (
    g854_n,
    G1928_o2_p,
    n4572_o2_n_spl_00
  );


  or

  (
    g855_n,
    G1929_o2_n,
    n4653_o2_n_spl_0
  );


  or

  (
    g856_n,
    G1930_o2_p,
    n2241_lo_buf_o2_n_spl_0
  );


  and

  (
    g857_p,
    g850_n,
    g849_n
  );


  and

  (
    g858_p,
    g857_p,
    g851_n
  );


  and

  (
    g859_p,
    g858_p,
    g852_n
  );


  and

  (
    g860_p,
    g859_p,
    g853_n
  );


  and

  (
    g861_p,
    g860_p,
    g854_n
  );


  and

  (
    g862_p,
    g861_p,
    g855_n
  );


  and

  (
    g863_p,
    g862_p,
    g856_n
  );


  and

  (
    g864_p,
    g863_p,
    G519_o2_p_spl_000
  );


  or

  (
    g865_n,
    g864_p,
    g848_p
  );


  and

  (
    g866_p,
    g865_n,
    g801_n_spl_00
  );


  or

  (
    g867_n,
    G2592_o2_p,
    G2296_o2_p
  );


  or

  (
    g868_n,
    G2592_o2_n,
    G2296_o2_n
  );


  and

  (
    g869_p,
    g868_n,
    g867_n
  );


  and

  (
    g870_p,
    n852_inv_n_spl_,
    n4816_o2_n_spl_
  );


  or

  (
    g870_n,
    n852_inv_p_spl_1,
    n4816_o2_p_spl_
  );


  and

  (
    g871_p,
    g870_p,
    n4389_o2_p_spl_0
  );


  or

  (
    g871_n,
    g870_n,
    n4389_o2_n_spl_0
  );


  and

  (
    g872_p,
    g871_p_spl_0,
    g869_p
  );


  and

  (
    g873_p,
    G772_o2_n_spl_,
    G519_o2_n_spl_00
  );


  or

  (
    g873_n,
    G772_o2_p_spl_,
    G519_o2_p_spl_00
  );


  and

  (
    g874_p,
    g873_p_spl_0,
    g737_n_spl_
  );


  and

  (
    g875_p,
    G772_o2_n_spl_,
    n4389_o2_n_spl_1
  );


  or

  (
    g875_n,
    G772_o2_p_spl_,
    n4389_o2_p_spl_1
  );


  and

  (
    g876_p,
    g875_n_spl_0,
    g873_n_spl_0
  );


  or

  (
    g876_n,
    g875_p_spl_0,
    g873_p_spl_0
  );


  and

  (
    g877_p,
    g876_p_spl_,
    G422_o2_n
  );


  or

  (
    g878_n,
    g875_p_spl_0,
    g874_p
  );


  or

  (
    g879_n,
    g878_n,
    g877_p
  );


  and

  (
    g880_p,
    g871_n_spl_0,
    g801_p_spl_0
  );


  or

  (
    g880_n,
    g871_p_spl_0,
    g801_n_spl_01
  );


  and

  (
    g881_p,
    g880_p_spl_,
    g879_n
  );


  or

  (
    g882_n,
    g872_p,
    g866_p
  );


  or

  (
    g883_n,
    g882_n,
    g881_p
  );


  or

  (
    g884_n,
    g883_n,
    g812_n_spl_00
  );


  and

  (
    g885_p,
    G1867_o2_n,
    n1977_lo_buf_o2_p
  );


  and

  (
    g886_p,
    G1868_o2_n,
    n1068_inv_n_spl_
  );


  and

  (
    g887_p,
    G1869_o2_p,
    n1071_inv_n_spl_
  );


  and

  (
    g888_p,
    G1870_o2_n,
    n1050_inv_n_spl_
  );


  and

  (
    g889_p,
    G1871_o2_n,
    n1056_inv_n_spl_
  );


  and

  (
    g890_p,
    G1872_o2_n,
    n858_inv_n_spl_
  );


  and

  (
    g891_p,
    G1873_o2_p,
    n4651_o2_p_spl_
  );


  and

  (
    g892_p,
    G1874_o2_n,
    n4919_o2_p
  );


  or

  (
    g893_n,
    g886_p,
    g885_p
  );


  or

  (
    g894_n,
    g893_n,
    g887_p
  );


  or

  (
    g895_n,
    g894_n,
    g888_p
  );


  or

  (
    g896_n,
    g895_n,
    g889_p
  );


  or

  (
    g897_n,
    g896_n,
    g890_p
  );


  or

  (
    g898_n,
    g897_n,
    g891_p
  );


  or

  (
    g899_n,
    g898_n,
    g892_p
  );


  or

  (
    g900_n,
    g899_n,
    G519_o2_p_spl_01
  );


  and

  (
    g901_p,
    G1931_o2_n,
    n2265_lo_buf_o2_p_spl_
  );


  and

  (
    g902_p,
    G1932_o2_n,
    n1053_inv_n_spl_
  );


  and

  (
    g903_p,
    G1933_o2_p,
    n1074_inv_n
  );


  and

  (
    g904_p,
    G1934_o2_n,
    n4571_o2_p_spl_
  );


  and

  (
    g905_p,
    G1935_o2_n,
    n4572_o2_p_spl_
  );


  and

  (
    g906_p,
    G1936_o2_n,
    n4653_o2_p_spl_
  );


  and

  (
    g907_p,
    G1937_o2_p,
    n2241_lo_buf_o2_p_spl_
  );


  and

  (
    g908_p,
    G1938_o2_n,
    n2253_lo_buf_o2_p_spl_
  );


  or

  (
    g909_n,
    g902_p,
    g901_p
  );


  or

  (
    g910_n,
    g909_n,
    g903_p
  );


  or

  (
    g911_n,
    g910_n,
    g904_p
  );


  or

  (
    g912_n,
    g911_n,
    g905_p
  );


  or

  (
    g913_n,
    g912_n,
    g906_p
  );


  or

  (
    g914_n,
    g913_n,
    g907_p
  );


  or

  (
    g915_n,
    g914_n,
    g908_p
  );


  or

  (
    g916_n,
    g915_n,
    G519_o2_n_spl_01
  );


  and

  (
    g917_p,
    g916_n,
    g900_n
  );


  or

  (
    g918_n,
    g917_p,
    g801_p_spl_1
  );


  and

  (
    g919_p,
    G2651_o2_n,
    G2497_o2_n
  );


  and

  (
    g920_p,
    G2651_o2_p,
    G2497_o2_p
  );


  or

  (
    g921_n,
    g920_p,
    g919_p
  );


  or

  (
    g922_n,
    g921_n,
    g871_n_spl_0
  );


  or

  (
    g923_n,
    g873_n_spl_0,
    g740_p_spl_
  );


  or

  (
    g924_n,
    g876_n_spl_,
    G434_o2_p_spl_
  );


  and

  (
    g925_p,
    g923_n,
    g875_n_spl_0
  );


  and

  (
    g926_p,
    g925_p,
    g924_n
  );


  or

  (
    g927_n,
    g926_p,
    g880_n_spl_
  );


  and

  (
    g928_p,
    g922_n,
    g918_n
  );


  and

  (
    g929_p,
    g928_p,
    g927_n
  );


  and

  (
    g930_p,
    g929_p,
    g812_p_spl_
  );


  or

  (
    g931_n,
    G1875_o2_p,
    n4919_o2_n_spl_01
  );


  or

  (
    g932_n,
    G1876_o2_p,
    n1062_inv_p_spl_01
  );


  or

  (
    g933_n,
    G1877_o2_n,
    n1068_inv_p_spl_00
  );


  or

  (
    g934_n,
    G1878_o2_p,
    n1071_inv_p_spl_01
  );


  or

  (
    g935_n,
    G1879_o2_p,
    n1050_inv_p_spl_00
  );


  or

  (
    g936_n,
    G1880_o2_p,
    n1056_inv_p_spl_01
  );


  or

  (
    g937_n,
    G1881_o2_n,
    n858_inv_p_spl_01
  );


  or

  (
    g938_n,
    G1882_o2_p,
    n4651_o2_n_spl_01
  );


  and

  (
    g939_p,
    g932_n,
    g931_n
  );


  and

  (
    g940_p,
    g939_p,
    g933_n
  );


  and

  (
    g941_p,
    g940_p,
    g934_n
  );


  and

  (
    g942_p,
    g941_p,
    g935_n
  );


  and

  (
    g943_p,
    g942_p,
    g936_n
  );


  and

  (
    g944_p,
    g943_p,
    g937_n
  );


  and

  (
    g945_p,
    g944_p,
    g938_n
  );


  and

  (
    g946_p,
    g945_p,
    G519_o2_n_spl_01
  );


  or

  (
    g947_n,
    G1939_o2_p,
    n2277_lo_buf_o2_n
  );


  or

  (
    g948_n,
    G1940_o2_p,
    n1074_inv_p_spl_01
  );


  or

  (
    g949_n,
    G1941_o2_n,
    n4571_o2_n_spl_01
  );


  or

  (
    g950_n,
    G1942_o2_p,
    n4572_o2_n_spl_0
  );


  or

  (
    g951_n,
    G1943_o2_p,
    n4653_o2_n_spl_1
  );


  or

  (
    g952_n,
    G1944_o2_p,
    n2241_lo_buf_o2_n_spl_0
  );


  or

  (
    g953_n,
    G1945_o2_n,
    n2253_lo_buf_o2_n_spl_
  );


  or

  (
    g954_n,
    G1946_o2_p,
    n2265_lo_buf_o2_n
  );


  and

  (
    g955_p,
    g948_n,
    g947_n
  );


  and

  (
    g956_p,
    g955_p,
    g949_n
  );


  and

  (
    g957_p,
    g956_p,
    g950_n
  );


  and

  (
    g958_p,
    g957_p,
    g951_n
  );


  and

  (
    g959_p,
    g958_p,
    g952_n
  );


  and

  (
    g960_p,
    g959_p,
    g953_n
  );


  and

  (
    g961_p,
    g960_p,
    g954_n
  );


  and

  (
    g962_p,
    g961_p,
    G519_o2_p_spl_01
  );


  or

  (
    g963_n,
    g962_p,
    g946_p
  );


  and

  (
    g964_p,
    g963_n,
    g801_n_spl_01
  );


  or

  (
    g965_n,
    G2598_o2_p,
    G2302_o2_p
  );


  or

  (
    g966_n,
    G2598_o2_n,
    G2302_o2_n
  );


  and

  (
    g967_p,
    g966_n,
    g965_n
  );


  and

  (
    g968_p,
    g967_p,
    g871_p_spl_
  );


  or

  (
    g969_n,
    G2038_o2_p,
    G1023_o2_p
  );


  or

  (
    g970_n,
    G1318_o2_n,
    G736_o2_n
  );


  and

  (
    g971_p,
    g970_n,
    g969_n
  );


  and

  (
    g972_p,
    g971_p,
    g873_p_spl_
  );


  or

  (
    g973_n,
    G787_o2_p,
    G461_o2_p_spl_
  );


  and

  (
    g974_p,
    g973_n,
    g875_p_spl_
  );


  and

  (
    g975_p,
    g876_p_spl_,
    G447_o2_n
  );


  or

  (
    g976_n,
    g974_p,
    g972_p
  );


  or

  (
    g977_n,
    g976_n,
    g975_p
  );


  and

  (
    g978_p,
    g977_n,
    g880_p_spl_
  );


  or

  (
    g979_n,
    g968_p,
    g964_p
  );


  or

  (
    g980_n,
    g979_n,
    g978_p
  );


  or

  (
    g981_n,
    g980_n,
    g812_n_spl_01
  );


  and

  (
    g982_p,
    G1883_o2_n,
    n4651_o2_p_spl_
  );


  and

  (
    g983_p,
    G1884_o2_n,
    n1053_inv_n_spl_
  );


  and

  (
    g984_p,
    G1885_o2_p,
    n1062_inv_n
  );


  and

  (
    g985_p,
    G1886_o2_n,
    n1068_inv_n_spl_
  );


  and

  (
    g986_p,
    G1887_o2_n,
    n1071_inv_n_spl_
  );


  and

  (
    g987_p,
    G1888_o2_n,
    n1050_inv_n_spl_
  );


  and

  (
    g988_p,
    G1889_o2_p,
    n1056_inv_n_spl_
  );


  and

  (
    g989_p,
    G1890_o2_n,
    n858_inv_n_spl_
  );


  or

  (
    g990_n,
    g983_p,
    g982_p
  );


  or

  (
    g991_n,
    g990_n,
    g984_p
  );


  or

  (
    g992_n,
    g991_n,
    g985_p
  );


  or

  (
    g993_n,
    g992_n,
    g986_p
  );


  or

  (
    g994_n,
    g993_n,
    g987_p
  );


  or

  (
    g995_n,
    g994_n,
    g988_p
  );


  or

  (
    g996_n,
    g995_n,
    g989_p
  );


  or

  (
    g997_n,
    g996_n,
    G519_o2_p_spl_10
  );


  and

  (
    g998_p,
    G1947_o2_n,
    n2289_lo_buf_o2_p
  );


  and

  (
    g999_p,
    G1948_o2_n,
    n4571_o2_p_spl_
  );


  and

  (
    g1000_p,
    G1949_o2_p,
    n4572_o2_p_spl_
  );


  and

  (
    g1001_p,
    G1950_o2_n,
    n4653_o2_p_spl_
  );


  and

  (
    g1002_p,
    G1951_o2_n,
    n2241_lo_buf_o2_p_spl_
  );


  and

  (
    g1003_p,
    G1952_o2_n,
    n2253_lo_buf_o2_p_spl_
  );


  and

  (
    g1004_p,
    G1953_o2_p,
    n2265_lo_buf_o2_p_spl_
  );


  and

  (
    g1005_p,
    G1954_o2_n,
    n2277_lo_buf_o2_p
  );


  or

  (
    g1006_n,
    g999_p,
    g998_p
  );


  or

  (
    g1007_n,
    g1006_n,
    g1000_p
  );


  or

  (
    g1008_n,
    g1007_n,
    g1001_p
  );


  or

  (
    g1009_n,
    g1008_n,
    g1002_p
  );


  or

  (
    g1010_n,
    g1009_n,
    g1003_p
  );


  or

  (
    g1011_n,
    g1010_n,
    g1004_p
  );


  or

  (
    g1012_n,
    g1011_n,
    g1005_p
  );


  or

  (
    g1013_n,
    g1012_n,
    G519_o2_n_spl_10
  );


  and

  (
    g1014_p,
    g1013_n,
    g997_n
  );


  or

  (
    g1015_n,
    g1014_p,
    g801_p_spl_1
  );


  and

  (
    g1016_p,
    G2604_o2_n,
    G2308_o2_n
  );


  and

  (
    g1017_p,
    G2604_o2_p,
    G2308_o2_p
  );


  or

  (
    g1018_n,
    g1017_p,
    g1016_p
  );


  or

  (
    g1019_n,
    g1018_n,
    g871_n_spl_
  );


  and

  (
    g1020_p,
    G1024_o2_n,
    n1176_inv_n
  );


  and

  (
    g1021_p,
    G935_o2_p_spl_,
    G739_o2_p
  );


  or

  (
    g1022_n,
    g1021_p,
    g1020_p
  );


  or

  (
    g1023_n,
    g1022_n,
    g873_n_spl_
  );


  and

  (
    g1024_p,
    g734_n_spl_,
    n4454_o2_p_spl_
  );


  or

  (
    g1025_n,
    g1024_p,
    g875_n_spl_
  );


  or

  (
    g1026_n,
    g876_n_spl_,
    G461_o2_p_spl_
  );


  and

  (
    g1027_p,
    g1025_n,
    g1023_n
  );


  and

  (
    g1028_p,
    g1027_p,
    g1026_n
  );


  or

  (
    g1029_n,
    g1028_p,
    g880_n_spl_
  );


  and

  (
    g1030_p,
    g1019_n,
    g1015_n
  );


  and

  (
    g1031_p,
    g1030_p,
    g1029_n
  );


  and

  (
    g1032_p,
    g1031_p,
    g812_p_spl_
  );


  and

  (
    g1033_p,
    G3117_o2_n,
    G3137_o2_p
  );


  or

  (
    g1033_n,
    G3117_o2_p,
    G3137_o2_n
  );


  and

  (
    g1034_p,
    g1033_n,
    G3039_o2_n_spl_0
  );


  and

  (
    g1035_p,
    g1033_p,
    G3039_o2_p_spl_0
  );


  or

  (
    g1036_n,
    g1035_p,
    g1034_p
  );


  or

  (
    g1037_n,
    g1036_n,
    g743_p_spl_01
  );


  and

  (
    g1038_p,
    G3038_o2_n,
    G3066_o2_p
  );


  or

  (
    g1038_n,
    G3038_o2_p,
    G3066_o2_n
  );


  and

  (
    g1039_p,
    g1038_n,
    G2923_o2_n_spl_
  );


  and

  (
    g1040_p,
    g1038_p,
    G2923_o2_p_spl_
  );


  or

  (
    g1041_n,
    g1040_p,
    g1039_p
  );


  or

  (
    g1042_n,
    g1041_n,
    g743_p_spl_01
  );


  and

  (
    g1043_p,
    n2061_lo_buf_o2_p_spl_,
    G875_o2_n
  );


  or

  (
    g1043_n,
    n2061_lo_buf_o2_n,
    G875_o2_p
  );


  and

  (
    g1044_p,
    g1043_p_spl_,
    n2313_lo_buf_o2_p_spl_
  );


  or

  (
    g1044_n,
    g1043_n_spl_,
    n2313_lo_buf_o2_n
  );


  and

  (
    g1045_p,
    g1044_n_spl_00,
    g746_n_spl_
  );


  or

  (
    g1045_n,
    g1044_p_spl_00,
    g746_p
  );


  and

  (
    g1046_p,
    G2251_o2_n,
    G2248_o2_n
  );


  or

  (
    g1046_n,
    G2251_o2_p,
    G2248_o2_p
  );


  and

  (
    g1047_p,
    G2255_o2_n,
    G2254_o2_n
  );


  or

  (
    g1047_n,
    G2255_o2_p,
    G2254_o2_p
  );


  and

  (
    g1048_p,
    g1047_p,
    G2014_o2_n
  );


  or

  (
    g1048_n,
    g1047_n,
    G2014_o2_p
  );


  and

  (
    g1049_p,
    g1048_n,
    g1046_p
  );


  or

  (
    g1049_n,
    g1048_p,
    g1046_n
  );


  and

  (
    g1050_p,
    G2507_o2_p_spl_0,
    G2444_o2_p_spl_0
  );


  or

  (
    g1050_n,
    G2507_o2_n_spl_0,
    G2444_o2_n_spl_0
  );


  and

  (
    g1051_p,
    g1050_p,
    G2451_o2_p
  );


  or

  (
    g1051_n,
    g1050_n,
    G2451_o2_n
  );


  and

  (
    g1052_p,
    g1051_p,
    g1049_p_spl_0
  );


  or

  (
    g1052_n,
    g1051_n,
    g1049_n_spl_0
  );


  and

  (
    g1053_p,
    G2627_o2_n,
    G2287_o2_n
  );


  or

  (
    g1053_n,
    G2627_o2_p,
    G2287_o2_p
  );


  and

  (
    g1054_p,
    G2398_o2_p,
    G2583_o2_p
  );


  or

  (
    g1054_n,
    G2398_o2_n,
    G2583_o2_n
  );


  and

  (
    g1055_p,
    g1054_n,
    g1053_n
  );


  or

  (
    g1055_n,
    g1054_p,
    g1053_p
  );


  and

  (
    g1056_p,
    G3024_o2_n_spl_,
    G2902_o2_p_spl_
  );


  or

  (
    g1056_n,
    G3024_o2_p_spl_,
    G2902_o2_n_spl_
  );


  and

  (
    g1057_p,
    G3024_o2_p_spl_,
    G2902_o2_n_spl_
  );


  or

  (
    g1057_n,
    G3024_o2_n_spl_,
    G2902_o2_p_spl_
  );


  and

  (
    g1058_p,
    g1057_n,
    g1056_n
  );


  or

  (
    g1058_n,
    g1057_p,
    g1056_p
  );


  or

  (
    g1059_n,
    g1058_p_spl_0,
    g752_p_spl_10
  );


  and

  (
    g1060_p,
    G1689_o2_p_spl_0,
    n2013_lo_buf_o2_p_spl_
  );


  or

  (
    g1060_n,
    G1689_o2_n_spl_0,
    n2013_lo_buf_o2_n
  );


  and

  (
    g1061_p,
    g1060_p,
    G1955_o2_n_spl_
  );


  or

  (
    g1061_n,
    g1060_n,
    G1955_o2_p_spl_
  );


  and

  (
    g1062_p,
    G1689_o2_p_spl_0,
    n2025_lo_buf_o2_p_spl_
  );


  or

  (
    g1062_n,
    G1689_o2_n_spl_0,
    n2025_lo_buf_o2_n_spl_
  );


  and

  (
    g1063_p,
    g1062_p,
    G1958_o2_n_spl_
  );


  or

  (
    g1063_n,
    g1062_n,
    G1958_o2_p_spl_
  );


  and

  (
    g1064_p,
    g1063_n,
    g1061_n
  );


  or

  (
    g1064_n,
    g1063_p,
    g1061_p
  );


  and

  (
    g1065_p,
    G1693_o2_n_spl_0,
    n2037_lo_buf_o2_p_spl_
  );


  or

  (
    g1065_n,
    G1693_o2_p_spl_0,
    n2037_lo_buf_o2_n_spl_
  );


  and

  (
    g1066_p,
    g1065_p,
    G1958_o2_n_spl_
  );


  or

  (
    g1066_n,
    g1065_n,
    G1958_o2_p_spl_
  );


  and

  (
    g1067_p,
    G1693_o2_n_spl_0,
    n2049_lo_buf_o2_p_spl_
  );


  or

  (
    g1067_n,
    G1693_o2_p_spl_0,
    n2049_lo_buf_o2_n_spl_0
  );


  and

  (
    g1068_p,
    g1067_p,
    G1955_o2_n_spl_
  );


  or

  (
    g1068_n,
    g1067_n,
    G1955_o2_p_spl_
  );


  and

  (
    g1069_p,
    g1068_n,
    g1066_n
  );


  or

  (
    g1069_n,
    g1068_p,
    g1066_p
  );


  and

  (
    g1070_p,
    g1069_p,
    G1693_o2_n_spl_
  );


  or

  (
    g1070_n,
    g1069_n,
    G1693_o2_p_spl_
  );


  and

  (
    g1071_p,
    g1070_n,
    g1064_p
  );


  or

  (
    g1071_n,
    g1070_p,
    g1064_n_spl_
  );


  and

  (
    g1072_p,
    g1071_p_spl_00,
    G2502_o2_p_spl_
  );


  or

  (
    g1072_n,
    g1071_n_spl_0,
    G2502_o2_n
  );


  or

  (
    g1073_n,
    g1072_n,
    G2437_o2_n
  );


  or

  (
    g1074_n,
    g1073_n,
    G2441_o2_n
  );


  or

  (
    g1075_n,
    G3107_o2_n,
    G2975_o2_p
  );


  or

  (
    g1076_n,
    G3107_o2_p,
    G2975_o2_n
  );


  and

  (
    g1077_p,
    g1076_n,
    g1075_n
  );


  or

  (
    g1078_n,
    g1077_p_spl_0,
    g752_p_spl_10
  );


  and

  (
    g1079_p,
    G1689_o2_p_spl_,
    G1176_o2_p
  );


  or

  (
    g1079_n,
    G1689_o2_n_spl_,
    G1176_o2_n
  );


  or

  (
    g1080_n,
    g832_p_spl_,
    g753_p_spl_
  );


  or

  (
    g1081_n,
    g1080_n,
    g930_p_spl_
  );


  and

  (
    g1082_p,
    g1042_n_spl_,
    g757_n_spl_
  );


  and

  (
    g1083_p,
    g1082_p,
    g981_n_spl_
  );


  and

  (
    g1084_p,
    g1037_n_spl_,
    g761_n_spl_
  );


  and

  (
    g1085_p,
    g1084_p,
    g813_n_spl_
  );


  and

  (
    g1086_p,
    g822_n_spl_,
    g765_n_spl_
  );


  and

  (
    g1087_p,
    g1086_p,
    g884_n_spl_
  );


  and

  (
    g1088_p,
    n2301_lo_buf_o2_p_spl_0,
    G2669_o2_n
  );


  or

  (
    g1088_n,
    n2301_lo_buf_o2_n_spl_,
    G2669_o2_p
  );


  and

  (
    g1089_p,
    G2759_o2_n_spl_,
    G2666_o2_p_spl_
  );


  or

  (
    g1089_n,
    G2759_o2_p_spl_,
    G2666_o2_n_spl_
  );


  and

  (
    g1090_p,
    G2759_o2_p_spl_,
    G2666_o2_n_spl_
  );


  or

  (
    g1090_n,
    G2759_o2_n_spl_,
    G2666_o2_p_spl_
  );


  and

  (
    g1091_p,
    g1090_n,
    g1089_n
  );


  or

  (
    g1091_n,
    g1090_p,
    g1089_p
  );


  or

  (
    g1092_n,
    g1091_n,
    g1088_n
  );


  or

  (
    g1093_n,
    g1091_p,
    g1088_p
  );


  and

  (
    g1094_p,
    g1093_n,
    g1092_n
  );


  or

  (
    g1095_n,
    g1094_p_spl_,
    g752_p_spl_1
  );


  or

  (
    g1096_n,
    G1529_o2_p_spl_0,
    n1917_lo_n
  );


  or

  (
    g1097_n,
    G1538_o2_p_spl_0,
    n4651_o2_n_spl_01
  );


  or

  (
    g1098_n,
    G1547_o2_n_spl_0,
    n4919_o2_n_spl_01
  );


  or

  (
    g1099_n,
    n1977_lo_buf_o2_n_spl_0,
    G1556_o2_p_spl_0
  );


  or

  (
    g1100_n,
    n1965_lo_buf_o2_n_spl_0,
    G1565_o2_p_spl_0
  );


  or

  (
    g1101_n,
    n1953_lo_buf_o2_n_spl_0,
    G1574_o2_p_spl_0
  );


  or

  (
    g1102_n,
    n1941_lo_buf_o2_n_spl_0,
    G1583_o2_n_spl_0
  );


  or

  (
    g1103_n,
    G1592_o2_p_spl_0,
    n1929_lo_n_spl_
  );


  and

  (
    g1104_p,
    g1097_n,
    g1096_n
  );


  and

  (
    g1105_p,
    g1104_p,
    g1098_n
  );


  and

  (
    g1106_p,
    g1105_p,
    g1099_n
  );


  and

  (
    g1107_p,
    g1106_p,
    g1100_n
  );


  and

  (
    g1108_p,
    g1107_p,
    g1101_n
  );


  and

  (
    g1109_p,
    g1108_p,
    g1102_n
  );


  and

  (
    g1110_p,
    g1109_p,
    g1103_n
  );


  and

  (
    g1111_p,
    n4539_o2_p_spl_0,
    n4389_o2_p_spl_1
  );


  or

  (
    g1111_n,
    n4539_o2_n_spl_0,
    n4389_o2_n_spl_1
  );


  and

  (
    g1112_p,
    g1111_p,
    g1110_p
  );


  or

  (
    g1113_n,
    G1601_o2_p_spl_0,
    n4571_o2_n_spl_01
  );


  or

  (
    g1114_n,
    n1056_inv_p_spl_01,
    G1610_o2_p_spl_0
  );


  or

  (
    g1115_n,
    n1050_inv_p_spl_01,
    G1619_o2_n_spl_0
  );


  or

  (
    g1116_n,
    n1071_inv_p_spl_01,
    G1628_o2_p_spl_0
  );


  or

  (
    g1117_n,
    n1068_inv_p_spl_01,
    G1637_o2_p_spl_0
  );


  or

  (
    g1118_n,
    n1062_inv_p_spl_01,
    G1646_o2_p_spl_0
  );


  or

  (
    g1119_n,
    n1053_inv_p_spl_01,
    G1655_o2_n_spl_0
  );


  or

  (
    g1120_n,
    n1074_inv_p_spl_01,
    G1664_o2_p_spl_0
  );


  and

  (
    g1121_p,
    g1114_n,
    g1113_n
  );


  and

  (
    g1122_p,
    g1121_p,
    g1115_n
  );


  and

  (
    g1123_p,
    g1122_p,
    g1116_n
  );


  and

  (
    g1124_p,
    g1123_p,
    g1117_n
  );


  and

  (
    g1125_p,
    g1124_p,
    g1118_n
  );


  and

  (
    g1126_p,
    g1125_p,
    g1119_n
  );


  and

  (
    g1127_p,
    g1126_p,
    g1120_n
  );


  and

  (
    g1128_p,
    G519_o2_n_spl_10,
    n4539_o2_p_spl_
  );


  or

  (
    g1128_n,
    G519_o2_p_spl_10,
    n4539_o2_n_spl_
  );


  and

  (
    g1129_p,
    g1128_p,
    g1127_p
  );


  and

  (
    g1130_p,
    g1128_n,
    g1111_n
  );


  and

  (
    g1131_p,
    g1130_p,
    n861_inv_n_spl_
  );


  or

  (
    g1132_n,
    g1129_p,
    g1112_p
  );


  or

  (
    g1133_n,
    g1132_n,
    g1131_p
  );


  and

  (
    g1134_p,
    g1133_n,
    g801_n_spl_10
  );


  or

  (
    g1135_n,
    G2512_o2_p,
    G2015_o2_p
  );


  or

  (
    g1136_n,
    G2512_o2_n,
    G2015_o2_n
  );


  and

  (
    g1137_p,
    g1136_n,
    g1135_n
  );


  and

  (
    g1138_p,
    g1137_p,
    g806_p_spl_0
  );


  and

  (
    g1139_p,
    g808_p_spl_0,
    n861_inv_n_spl_
  );


  or

  (
    g1140_n,
    g1138_p,
    g1134_p
  );


  or

  (
    g1141_n,
    g1140_n,
    g1139_p
  );


  or

  (
    g1142_n,
    g1141_n,
    g812_n_spl_01
  );


  or

  (
    g1143_n,
    G1529_o2_p_spl_0,
    n1929_lo_n_spl_
  );


  or

  (
    g1144_n,
    G1538_o2_p_spl_0,
    n858_inv_p_spl_01
  );


  or

  (
    g1145_n,
    G1547_o2_n_spl_0,
    n4651_o2_n_spl_1
  );


  or

  (
    g1146_n,
    G1556_o2_p_spl_0,
    n4919_o2_n_spl_1
  );


  or

  (
    g1147_n,
    n1977_lo_buf_o2_n_spl_1,
    G1565_o2_p_spl_0
  );


  or

  (
    g1148_n,
    n1965_lo_buf_o2_n_spl_1,
    G1574_o2_p_spl_0
  );


  or

  (
    g1149_n,
    n1953_lo_buf_o2_n_spl_1,
    G1583_o2_n_spl_0
  );


  or

  (
    g1150_n,
    n1941_lo_buf_o2_n_spl_,
    G1592_o2_p_spl_0
  );


  and

  (
    g1151_p,
    g1144_n,
    g1143_n
  );


  and

  (
    g1152_p,
    g1151_p,
    g1145_n
  );


  and

  (
    g1153_p,
    g1152_p,
    g1146_n
  );


  and

  (
    g1154_p,
    g1153_p,
    g1147_n
  );


  and

  (
    g1155_p,
    g1154_p,
    g1148_n
  );


  and

  (
    g1156_p,
    g1155_p,
    g1149_n
  );


  and

  (
    g1157_p,
    g1156_p,
    g1150_n
  );


  and

  (
    g1158_p,
    g1157_p,
    G519_o2_n_spl_11
  );


  or

  (
    g1159_n,
    G1601_o2_p_spl_0,
    n4572_o2_n_spl_1
  );


  or

  (
    g1160_n,
    n1050_inv_p_spl_01,
    G1610_o2_p_spl_0
  );


  or

  (
    g1161_n,
    n1071_inv_p_spl_1,
    G1619_o2_n_spl_0
  );


  or

  (
    g1162_n,
    n1068_inv_p_spl_01,
    G1628_o2_p_spl_0
  );


  or

  (
    g1163_n,
    n1062_inv_p_spl_10,
    G1637_o2_p_spl_0
  );


  or

  (
    g1164_n,
    n1053_inv_p_spl_01,
    G1646_o2_p_spl_0
  );


  or

  (
    g1165_n,
    n1074_inv_p_spl_10,
    G1655_o2_n_spl_0
  );


  or

  (
    g1166_n,
    G1664_o2_p_spl_0,
    n4571_o2_n_spl_1
  );


  and

  (
    g1167_p,
    g1160_n,
    g1159_n
  );


  and

  (
    g1168_p,
    g1167_p,
    g1161_n
  );


  and

  (
    g1169_p,
    g1168_p,
    g1162_n
  );


  and

  (
    g1170_p,
    g1169_p,
    g1163_n
  );


  and

  (
    g1171_p,
    g1170_p,
    g1164_n
  );


  and

  (
    g1172_p,
    g1171_p,
    g1165_n
  );


  and

  (
    g1173_p,
    g1172_p,
    g1166_n
  );


  and

  (
    g1174_p,
    g1173_p,
    G519_o2_p_spl_11
  );


  or

  (
    g1175_n,
    g1174_p,
    g1158_p
  );


  and

  (
    g1176_p,
    g1175_n,
    g801_n_spl_10
  );


  or

  (
    g1177_n,
    n5301_o2_p,
    n5278_o2_p
  );


  or

  (
    g1178_n,
    n5301_o2_n,
    n5278_o2_n
  );


  and

  (
    g1179_p,
    g1178_n,
    g1177_n
  );


  and

  (
    g1180_p,
    g1179_p,
    g806_p_spl_1
  );


  and

  (
    g1181_p,
    g808_p_spl_1,
    G377_o2_n
  );


  or

  (
    g1182_n,
    g1180_p,
    g1176_p
  );


  or

  (
    g1183_n,
    g1182_n,
    g1181_p
  );


  or

  (
    g1184_n,
    g1183_n,
    g812_n_spl_1
  );


  or

  (
    g1185_n,
    n1953_lo_buf_o2_n_spl_1,
    G1529_o2_p_spl_
  );


  or

  (
    g1186_n,
    n1050_inv_p_spl_1,
    G1538_o2_p_spl_
  );


  or

  (
    g1187_n,
    n1056_inv_p_spl_1,
    G1547_o2_n_spl_
  );


  or

  (
    g1188_n,
    G1556_o2_p_spl_,
    n858_inv_p_spl_1
  );


  or

  (
    g1189_n,
    G1565_o2_p_spl_,
    n4651_o2_n_spl_1
  );


  or

  (
    g1190_n,
    G1574_o2_p_spl_,
    n4919_o2_n_spl_1
  );


  or

  (
    g1191_n,
    n1977_lo_buf_o2_n_spl_1,
    G1583_o2_n_spl_
  );


  or

  (
    g1192_n,
    n1965_lo_buf_o2_n_spl_1,
    G1592_o2_p_spl_
  );


  and

  (
    g1193_p,
    g1186_n,
    g1185_n
  );


  and

  (
    g1194_p,
    g1193_p,
    g1187_n
  );


  and

  (
    g1195_p,
    g1194_p,
    g1188_n
  );


  and

  (
    g1196_p,
    g1195_p,
    g1189_n
  );


  and

  (
    g1197_p,
    g1196_p,
    g1190_n
  );


  and

  (
    g1198_p,
    g1197_p,
    g1191_n
  );


  and

  (
    g1199_p,
    g1198_p,
    g1192_n
  );


  and

  (
    g1200_p,
    g1199_p,
    G519_o2_n_spl_11
  );


  or

  (
    g1201_n,
    n2241_lo_buf_o2_n_spl_,
    G1601_o2_p_spl_
  );


  or

  (
    g1202_n,
    n1068_inv_p_spl_1,
    G1610_o2_p_spl_
  );


  or

  (
    g1203_n,
    n1062_inv_p_spl_10,
    G1619_o2_n_spl_
  );


  or

  (
    g1204_n,
    n1053_inv_p_spl_1,
    G1628_o2_p_spl_
  );


  or

  (
    g1205_n,
    n1074_inv_p_spl_10,
    G1637_o2_p_spl_
  );


  or

  (
    g1206_n,
    G1646_o2_p_spl_,
    n4571_o2_n_spl_1
  );


  or

  (
    g1207_n,
    G1655_o2_n_spl_,
    n4572_o2_n_spl_1
  );


  or

  (
    g1208_n,
    G1664_o2_p_spl_,
    n4653_o2_n_spl_1
  );


  and

  (
    g1209_p,
    g1202_n,
    g1201_n
  );


  and

  (
    g1210_p,
    g1209_p,
    g1203_n
  );


  and

  (
    g1211_p,
    g1210_p,
    g1204_n
  );


  and

  (
    g1212_p,
    g1211_p,
    g1205_n
  );


  and

  (
    g1213_p,
    g1212_p,
    g1206_n
  );


  and

  (
    g1214_p,
    g1213_p,
    g1207_n
  );


  and

  (
    g1215_p,
    g1214_p,
    g1208_n
  );


  and

  (
    g1216_p,
    g1215_p,
    G519_o2_p_spl_11
  );


  or

  (
    g1217_n,
    g1216_p,
    g1200_p
  );


  and

  (
    g1218_p,
    g1217_n,
    g801_n_spl_1
  );


  or

  (
    g1219_n,
    n5094_o2_p,
    n5041_o2_p
  );


  or

  (
    g1220_n,
    n5094_o2_n,
    n5041_o2_n
  );


  and

  (
    g1221_p,
    g1220_n,
    g1219_n
  );


  and

  (
    g1222_p,
    g1221_p,
    g806_p_spl_1
  );


  and

  (
    g1223_p,
    g808_p_spl_1,
    n570_inv_n
  );


  or

  (
    g1224_n,
    g1222_p,
    g1218_p
  );


  or

  (
    g1225_n,
    g1224_n,
    g1223_p
  );


  or

  (
    g1226_n,
    g1225_n,
    g812_n_spl_1
  );


  or

  (
    g1227_n,
    g1077_p_spl_0,
    G3039_o2_p_spl_0
  );


  or

  (
    g1228_n,
    g1058_p_spl_0,
    g760_p_spl_0
  );


  or

  (
    g1229_n,
    g1228_n,
    g1077_p_spl_
  );


  or

  (
    g1230_n,
    g1229_n,
    G3039_o2_n_spl_0
  );


  and

  (
    g1231_p,
    g1230_n,
    g1227_n
  );


  or

  (
    g1232_n,
    g1231_p,
    g743_p_spl_10
  );


  and

  (
    g1233_p,
    g760_n,
    G3039_o2_n_spl_
  );


  or

  (
    g1233_n,
    g760_p_spl_,
    G3039_o2_p_spl_
  );


  or

  (
    g1234_n,
    g1233_n,
    g1058_p_spl_
  );


  or

  (
    g1235_n,
    g1233_p,
    g1058_n
  );


  and

  (
    g1236_p,
    g1235_n,
    g1234_n
  );


  or

  (
    g1237_n,
    g1236_p,
    g743_p_spl_10
  );


  or

  (
    g1238_n,
    g1094_p_spl_,
    g743_p_spl_11
  );


  or

  (
    g1239_n,
    g827_p_spl_,
    g826_p_spl_
  );


  or

  (
    g1240_n,
    g1239_n,
    g1032_p_spl_
  );


  and

  (
    g1241_p,
    G1738_o2_p_spl_,
    G1733_o2_p_spl_
  );


  or

  (
    g1241_n,
    G1738_o2_n_spl_,
    G1733_o2_n_spl_
  );


  and

  (
    g1242_p,
    g1241_p,
    G1751_o2_p_spl_
  );


  or

  (
    g1242_n,
    g1241_n,
    G1751_o2_n_spl_
  );


  and

  (
    g1243_p,
    g1242_p,
    G1764_o2_p_spl_
  );


  or

  (
    g1243_n,
    g1242_n,
    G1764_o2_n_spl_
  );


  and

  (
    g1244_p,
    g1243_p,
    G615_o2_p_spl_
  );


  or

  (
    g1244_n,
    g1243_n,
    G615_o2_n_spl_
  );


  and

  (
    g1245_p,
    G1738_o2_n_spl_,
    G1733_o2_n_spl_
  );


  or

  (
    g1245_n,
    G1738_o2_p_spl_,
    G1733_o2_p_spl_
  );


  and

  (
    g1246_p,
    g1245_p,
    G1751_o2_n_spl_
  );


  or

  (
    g1246_n,
    g1245_n,
    G1751_o2_p_spl_
  );


  and

  (
    g1247_p,
    g1246_p,
    G1764_o2_n_spl_
  );


  or

  (
    g1247_n,
    g1246_n,
    G1764_o2_p_spl_
  );


  and

  (
    g1248_p,
    g1247_p,
    G615_o2_n_spl_
  );


  or

  (
    g1248_n,
    g1247_n,
    G615_o2_p_spl_
  );


  and

  (
    g1249_p,
    g1248_n,
    g1244_n
  );


  or

  (
    g1249_n,
    g1248_p,
    g1244_p
  );


  and

  (
    g1250_p,
    g1249_n,
    g1044_n_spl_00
  );


  or

  (
    g1250_n,
    g1249_p,
    g1044_p_spl_00
  );


  and

  (
    g1251_p,
    g1052_p_spl_,
    g1044_p_spl_01
  );


  or

  (
    g1251_n,
    g1052_n,
    g1044_n_spl_01
  );


  and

  (
    g1252_p,
    g1251_n,
    g1250_n
  );


  or

  (
    g1252_n,
    g1251_p,
    g1250_p
  );


  and

  (
    g1253_p,
    g1237_n_spl_,
    g1059_n_spl_
  );


  and

  (
    g1254_p,
    g1253_p,
    g1184_n_spl_
  );


  and

  (
    g1255_p,
    g1232_n_spl_,
    g1078_n_spl_
  );


  and

  (
    g1256_p,
    g1255_p,
    g1142_n_spl_
  );


  and

  (
    g1257_p,
    g1238_n_spl_,
    g1095_n_spl_
  );


  and

  (
    g1258_p,
    g1257_p,
    g1226_n_spl_
  );


  and

  (
    g1259_p,
    G2359_o2_n,
    G2356_o2_n
  );


  or

  (
    g1259_n,
    G2359_o2_p,
    G2356_o2_p
  );


  and

  (
    g1260_p,
    g1259_n_spl_,
    g1071_p_spl_00
  );


  and

  (
    g1261_p,
    G2211_o2_n,
    G2208_o2_n
  );


  or

  (
    g1261_n,
    G2211_o2_p,
    G2208_o2_p
  );


  and

  (
    g1262_p,
    g1261_n_spl_,
    g1072_p
  );


  and

  (
    g1263_p,
    G2219_o2_n,
    G2216_o2_n
  );


  or

  (
    g1263_n,
    G2219_o2_p,
    G2216_o2_p
  );


  and

  (
    g1264_p,
    g1263_n_spl_,
    G2502_o2_p_spl_
  );


  and

  (
    g1265_p,
    g1264_p,
    G2437_o2_p
  );


  and

  (
    g1266_p,
    g1265_p,
    g1071_p_spl_01
  );


  or

  (
    g1267_n,
    g1260_p,
    g1064_n_spl_
  );


  or

  (
    g1268_n,
    g1267_n,
    g1262_p
  );


  or

  (
    g1269_n,
    g1268_n,
    g1266_p
  );


  and

  (
    g1270_p,
    g1044_n_spl_01,
    G2384_o2_p
  );


  or

  (
    g1270_n,
    g1044_p_spl_01,
    G2384_o2_n
  );


  and

  (
    g1271_p,
    n1554_inv_n_spl_,
    G2027_o2_n_spl_
  );


  or

  (
    g1271_n,
    n1554_inv_p_spl_0,
    G2027_o2_p_spl_0
  );


  and

  (
    g1272_p,
    n1554_inv_p_spl_0,
    G2027_o2_p_spl_0
  );


  or

  (
    g1272_n,
    n1554_inv_n_spl_,
    G2027_o2_n_spl_
  );


  and

  (
    g1273_p,
    g1272_n,
    g1271_n
  );


  or

  (
    g1273_n,
    g1272_p,
    g1271_p
  );


  and

  (
    g1274_p,
    g1044_n_spl_10,
    G2388_o2_p
  );


  or

  (
    g1274_n,
    g1044_p_spl_10,
    G2388_o2_n
  );


  and

  (
    g1275_p,
    g1274_n_spl_,
    g1273_n_spl_
  );


  or

  (
    g1275_n,
    g1274_p_spl_0,
    g1273_p_spl_0
  );


  and

  (
    g1276_p,
    g1275_n,
    g1270_n_spl_
  );


  or

  (
    g1276_n,
    g1275_p_spl_,
    g1270_p_spl_
  );


  and

  (
    g1277_p,
    n2097_lo_buf_o2_p_spl_0,
    n5326_o2_n_spl_
  );


  or

  (
    g1277_n,
    n2097_lo_buf_o2_n_spl_,
    n5326_o2_p_spl_0
  );


  and

  (
    g1278_p,
    n2097_lo_buf_o2_n_spl_,
    n5326_o2_p_spl_0
  );


  or

  (
    g1278_n,
    n2097_lo_buf_o2_p_spl_0,
    n5326_o2_n_spl_
  );


  and

  (
    g1279_p,
    g1278_n,
    g1277_n
  );


  or

  (
    g1279_n,
    g1278_p,
    g1277_p
  );


  and

  (
    g1280_p,
    n2133_lo_buf_o2_n_spl_,
    n5327_o2_p_spl_0
  );


  or

  (
    g1280_n,
    n2133_lo_buf_o2_p_spl_0,
    n5327_o2_n_spl_
  );


  and

  (
    g1281_p,
    n2133_lo_buf_o2_p_spl_0,
    n5327_o2_n_spl_
  );


  or

  (
    g1281_n,
    n2133_lo_buf_o2_n_spl_,
    n5327_o2_p_spl_0
  );


  and

  (
    g1282_p,
    g1281_n,
    g1280_n
  );


  or

  (
    g1282_n,
    g1281_p,
    g1280_p
  );


  and

  (
    g1283_p,
    g1074_n_spl_0,
    g1045_n_spl_00
  );


  or

  (
    g1284_n,
    g1283_p,
    g1269_n_spl_
  );


  and

  (
    g1285_p,
    g1259_n_spl_,
    g1043_n_spl_
  );


  or

  (
    g1285_n,
    g1259_p,
    g1043_p_spl_
  );


  and

  (
    g1286_p,
    n1557_inv_n_spl_,
    G2393_o2_n_spl_
  );


  or

  (
    g1286_n,
    n1557_inv_p_spl_0,
    G2393_o2_p_spl_0
  );


  and

  (
    g1287_p,
    n1557_inv_p_spl_0,
    G2393_o2_p_spl_0
  );


  or

  (
    g1287_n,
    n1557_inv_n_spl_,
    G2393_o2_n_spl_
  );


  and

  (
    g1288_p,
    g1287_n,
    g1286_n
  );


  or

  (
    g1288_n,
    g1287_p,
    g1286_p
  );


  and

  (
    g1289_p,
    g1261_n_spl_,
    g1044_n_spl_10
  );


  or

  (
    g1289_n,
    g1261_p,
    g1044_p_spl_10
  );


  and

  (
    g1290_p,
    g1289_p_spl_,
    g1288_p_spl_0
  );


  or

  (
    g1290_n,
    g1289_n_spl_,
    g1288_n_spl_0
  );


  and

  (
    g1291_p,
    G2577_o2_n_spl_,
    G2281_o2_n_spl_
  );


  or

  (
    g1291_n,
    G2577_o2_p_spl_,
    G2281_o2_p_spl_
  );


  and

  (
    g1292_p,
    G2577_o2_p_spl_,
    G2281_o2_p_spl_
  );


  or

  (
    g1292_n,
    G2577_o2_n_spl_,
    G2281_o2_n_spl_
  );


  and

  (
    g1293_p,
    g1292_n,
    g1291_n
  );


  or

  (
    g1293_n,
    g1292_p,
    g1291_p
  );


  and

  (
    g1294_p,
    g1263_n_spl_,
    g1044_n_spl_11
  );


  or

  (
    g1294_n,
    g1263_p,
    g1044_p_spl_11
  );


  and

  (
    g1295_p,
    g1293_p_spl_0,
    g1288_p_spl_0
  );


  or

  (
    g1295_n,
    g1293_n_spl_00,
    g1288_n_spl_0
  );


  and

  (
    g1296_p,
    g1295_p_spl_,
    g1294_n_spl_0
  );


  or

  (
    g1296_n,
    g1295_n_spl_,
    g1294_p_spl_0
  );


  and

  (
    g1297_p,
    g1295_p_spl_,
    g1055_p_spl_0
  );


  or

  (
    g1297_n,
    g1295_n_spl_,
    g1055_n_spl_00
  );


  and

  (
    g1298_p,
    g1297_p,
    g1045_n_spl_00
  );


  or

  (
    g1298_n,
    g1297_n,
    g1045_p_spl_00
  );


  and

  (
    g1299_p,
    g1290_n,
    g1285_n
  );


  or

  (
    g1299_n,
    g1290_p,
    g1285_p
  );


  and

  (
    g1300_p,
    g1299_p,
    g1296_n
  );


  or

  (
    g1300_n,
    g1299_n,
    g1296_p
  );


  and

  (
    g1301_p,
    g1300_p,
    g1298_n
  );


  or

  (
    g1301_n,
    g1300_n,
    g1298_p
  );


  and

  (
    g1302_p,
    n4921_o2_p_spl_,
    n4920_o2_p_spl_0
  );


  or

  (
    g1303_n,
    g1302_p_spl_,
    g1254_p_spl_0
  );


  or

  (
    g1304_n,
    g1302_p_spl_,
    g1256_p_spl_0
  );


  and

  (
    g1305_p,
    G1189_o2_p_spl_,
    G1756_o2_p
  );


  or

  (
    g1305_n,
    G1189_o2_n_spl_,
    G1756_o2_n
  );


  and

  (
    g1306_p,
    g1305_n_spl_,
    g1049_n_spl_0
  );


  or

  (
    g1306_n,
    g1305_p_spl_0,
    g1049_p_spl_0
  );


  and

  (
    g1307_p,
    g1305_p_spl_0,
    g1049_p_spl_1
  );


  or

  (
    g1307_n,
    g1305_n_spl_,
    g1049_n_spl_
  );


  and

  (
    g1308_p,
    g1307_n,
    g1306_n
  );


  or

  (
    g1308_n,
    g1307_p,
    g1306_p
  );


  and

  (
    g1309_p,
    n1761_lo_buf_o2_p_spl_0,
    n1749_lo_buf_o2_p_spl_00
  );


  or

  (
    g1309_n,
    n1761_lo_buf_o2_n,
    n1749_lo_buf_o2_n_spl_00
  );


  and

  (
    g1310_p,
    g1309_p_spl_0,
    G527_o2_n
  );


  or

  (
    g1310_n,
    g1309_n_spl_0,
    G527_o2_p
  );


  and

  (
    g1311_p,
    n1809_lo_buf_o2_n_spl_,
    n1749_lo_buf_o2_n_spl_00
  );


  or

  (
    g1311_n,
    n1809_lo_buf_o2_p_spl_0,
    n1749_lo_buf_o2_p_spl_00
  );


  and

  (
    g1312_p,
    g1310_n_spl_000,
    n2139_lo_buf_o2_p_spl_0
  );


  or

  (
    g1312_n,
    g1310_p_spl_00,
    n2139_lo_buf_o2_n_spl_0
  );


  and

  (
    g1313_p,
    g1312_p,
    g1311_n_spl_
  );


  or

  (
    g1313_n,
    g1312_n,
    g1311_p_spl_
  );


  and

  (
    g1314_p,
    g1310_n_spl_000,
    n2187_lo_buf_o2_p_spl_
  );


  or

  (
    g1314_n,
    g1310_p_spl_00,
    n2187_lo_buf_o2_n_spl_
  );


  and

  (
    g1315_p,
    g1314_p_spl_,
    g1311_p_spl_
  );


  or

  (
    g1315_n,
    g1314_n_spl_,
    g1311_n_spl_
  );


  and

  (
    g1316_p,
    n1899_lo_buf_o2_p_spl_00,
    G831_o2_n_spl_00
  );


  or

  (
    g1316_n,
    n1899_lo_buf_o2_n_spl_00,
    G831_o2_p_spl_00
  );


  and

  (
    g1317_p,
    n2121_lo_buf_o2_p_spl_0,
    G594_o2_n_spl_00
  );


  or

  (
    g1317_n,
    n2121_lo_buf_o2_n_spl_0,
    G594_o2_p_spl_00
  );


  and

  (
    g1318_p,
    G831_o2_p_spl_00,
    G594_o2_p_spl_00
  );


  or

  (
    g1318_n,
    G831_o2_n_spl_00,
    G594_o2_n_spl_00
  );


  and

  (
    g1319_p,
    g1318_p_spl_00,
    n2127_lo_buf_o2_p_spl_0
  );


  or

  (
    g1319_n,
    g1318_n_spl_00,
    n2127_lo_buf_o2_n_spl_0
  );


  and

  (
    g1320_p,
    g1317_n,
    g1316_n
  );


  or

  (
    g1320_n,
    g1317_p,
    g1316_p
  );


  and

  (
    g1321_p,
    g1320_p,
    g1319_n
  );


  or

  (
    g1321_n,
    g1320_n,
    g1319_p
  );


  and

  (
    g1322_p,
    g1321_n,
    g1310_n_spl_00
  );


  or

  (
    g1322_n,
    g1321_p,
    g1310_p_spl_01
  );


  and

  (
    g1323_p,
    g1315_n,
    g1313_n
  );


  or

  (
    g1323_n,
    g1315_p,
    g1313_p
  );


  and

  (
    g1324_p,
    g1323_p,
    g1322_n
  );


  or

  (
    g1324_n,
    g1323_n,
    g1322_p
  );


  and

  (
    g1325_p,
    G477_o2_n_spl_,
    n1809_lo_buf_o2_n_spl_
  );


  or

  (
    g1325_n,
    G477_o2_p_spl_,
    n1809_lo_buf_o2_p_spl_0
  );


  and

  (
    g1326_p,
    g1325_p,
    n1797_lo_buf_o2_n
  );


  or

  (
    g1326_n,
    g1325_n,
    n1797_lo_buf_o2_p_spl_
  );


  and

  (
    g1327_p,
    g1310_n_spl_01,
    n2151_lo_buf_o2_p_spl_0
  );


  or

  (
    g1327_n,
    g1310_p_spl_01,
    n2151_lo_buf_o2_n_spl_
  );


  and

  (
    g1328_p,
    g1327_p,
    g1326_n_spl_0
  );


  or

  (
    g1328_n,
    g1327_n,
    g1326_p_spl_0
  );


  and

  (
    g1329_p,
    g1326_p_spl_0,
    g1314_p_spl_
  );


  or

  (
    g1329_n,
    g1326_n_spl_0,
    g1314_n_spl_
  );


  and

  (
    g1330_p,
    n2199_lo_buf_o2_p_spl_0,
    G831_o2_n_spl_01
  );


  or

  (
    g1330_n,
    n2199_lo_buf_o2_n_spl_,
    G831_o2_p_spl_01
  );


  and

  (
    g1331_p,
    n2127_lo_buf_o2_p_spl_0,
    G594_o2_n_spl_01
  );


  or

  (
    g1331_n,
    n2127_lo_buf_o2_n_spl_0,
    G594_o2_p_spl_01
  );


  and

  (
    g1332_p,
    g1318_p_spl_00,
    n2139_lo_buf_o2_p_spl_0
  );


  or

  (
    g1332_n,
    g1318_n_spl_00,
    n2139_lo_buf_o2_n_spl_0
  );


  and

  (
    g1333_p,
    g1331_n,
    g1330_n
  );


  or

  (
    g1333_n,
    g1331_p,
    g1330_p
  );


  and

  (
    g1334_p,
    g1333_p,
    g1332_n
  );


  or

  (
    g1334_n,
    g1333_n,
    g1332_p
  );


  and

  (
    g1335_p,
    g1334_n,
    g1310_n_spl_01
  );


  or

  (
    g1335_n,
    g1334_p,
    g1310_p_spl_10
  );


  and

  (
    g1336_p,
    g1329_n_spl_,
    g1328_n
  );


  or

  (
    g1336_n,
    g1329_p_spl_0,
    g1328_p
  );


  and

  (
    g1337_p,
    g1336_p,
    g1335_n
  );


  or

  (
    g1337_n,
    g1336_n,
    g1335_p
  );


  and

  (
    g1338_p,
    g1310_n_spl_10,
    n2163_lo_p_spl_0
  );


  or

  (
    g1338_n,
    g1310_p_spl_10,
    n2163_lo_n
  );


  and

  (
    g1339_p,
    g1338_p,
    g1326_n_spl_1
  );


  or

  (
    g1339_n,
    g1338_n,
    g1326_p_spl_
  );


  and

  (
    g1340_p,
    n2211_lo_buf_o2_p_spl_,
    G831_o2_n_spl_01
  );


  or

  (
    g1340_n,
    n2211_lo_buf_o2_n,
    G831_o2_p_spl_01
  );


  and

  (
    g1341_p,
    n2139_lo_buf_o2_p_spl_1,
    G594_o2_n_spl_01
  );


  or

  (
    g1341_n,
    n2139_lo_buf_o2_n_spl_,
    G594_o2_p_spl_01
  );


  and

  (
    g1342_p,
    g1318_p_spl_01,
    n2151_lo_buf_o2_p_spl_0
  );


  or

  (
    g1342_n,
    g1318_n_spl_0,
    n2151_lo_buf_o2_n_spl_
  );


  and

  (
    g1343_p,
    g1341_n,
    g1340_n
  );


  or

  (
    g1343_n,
    g1341_p,
    g1340_p
  );


  and

  (
    g1344_p,
    g1343_p,
    g1342_n
  );


  or

  (
    g1344_n,
    g1343_n,
    g1342_p
  );


  and

  (
    g1345_p,
    g1344_n,
    g1310_n_spl_10
  );


  or

  (
    g1345_n,
    g1344_p,
    g1310_p_spl_1
  );


  and

  (
    g1346_p,
    g1339_n,
    g1329_n_spl_
  );


  or

  (
    g1346_n,
    g1339_p,
    g1329_p_spl_0
  );


  and

  (
    g1347_p,
    g1346_p,
    g1345_n
  );


  or

  (
    g1347_n,
    g1346_n,
    g1345_p
  );


  and

  (
    g1348_p,
    G501_o2_p_spl_000,
    n1854_lo_buf_o2_p_spl_00
  );


  or

  (
    g1348_n,
    G501_o2_n_spl_00,
    n1854_lo_buf_o2_n_spl_00
  );


  and

  (
    g1349_p,
    n1869_lo_buf_o2_n_spl_00,
    G667_o2_p_spl_000
  );


  or

  (
    g1349_n,
    n1869_lo_buf_o2_p_spl_00,
    G667_o2_n_spl_00
  );


  and

  (
    g1350_p,
    G501_o2_n_spl_00,
    G667_o2_n_spl_00
  );


  or

  (
    g1350_n,
    G501_o2_p_spl_000,
    G667_o2_p_spl_000
  );


  and

  (
    g1351_p,
    g1350_p_spl_00,
    n1833_lo_buf_o2_n_spl_0
  );


  or

  (
    g1351_n,
    g1350_n_spl_00,
    n1833_lo_buf_o2_p_spl_00
  );


  and

  (
    g1352_p,
    g1349_n,
    g1348_n
  );


  or

  (
    g1352_n,
    g1349_p,
    g1348_p
  );


  and

  (
    g1353_p,
    g1352_p,
    g1351_n
  );


  or

  (
    g1353_n,
    g1352_n,
    g1351_p
  );


  and

  (
    g1354_p,
    n1773_lo_buf_o2_p_spl_00,
    n1749_lo_buf_o2_p_spl_01
  );


  or

  (
    g1354_n,
    n1773_lo_buf_o2_n_spl_,
    n1749_lo_buf_o2_n_spl_01
  );


  and

  (
    g1355_p,
    g1354_p,
    n1785_lo_buf_o2_p_spl_0
  );


  or

  (
    g1355_n,
    g1354_n,
    n1785_lo_buf_o2_n_spl_
  );


  and

  (
    g1356_p,
    g1355_n,
    g1309_n_spl_0
  );


  or

  (
    g1356_n,
    g1355_p,
    g1309_p_spl_0
  );


  and

  (
    g1357_p,
    g1356_n_spl_000,
    g1353_n
  );


  or

  (
    g1357_n,
    g1356_p_spl_00,
    g1353_p
  );


  and

  (
    g1358_p,
    G491_o2_p,
    n1749_lo_buf_o2_n_spl_01
  );


  or

  (
    g1358_n,
    G491_o2_n,
    n1749_lo_buf_o2_p_spl_01
  );


  and

  (
    g1359_p,
    g1358_p_spl_000,
    n1854_lo_buf_o2_n_spl_00
  );


  or

  (
    g1359_n,
    g1358_n_spl_00,
    n1854_lo_buf_o2_p_spl_00
  );


  and

  (
    g1360_p,
    n1773_lo_buf_o2_p_spl_00,
    n1749_lo_buf_o2_n_spl_1
  );


  or

  (
    g1360_n,
    n1773_lo_buf_o2_n_spl_,
    n1749_lo_buf_o2_p_spl_10
  );


  and

  (
    g1361_p,
    g1358_n_spl_00,
    g1356_p_spl_00
  );


  or

  (
    g1361_n,
    g1358_p_spl_000,
    g1356_n_spl_000
  );


  and

  (
    g1362_p,
    g1360_n_spl_0,
    n1854_lo_buf_o2_p_spl_01
  );


  or

  (
    g1362_n,
    g1360_p_spl_0,
    n1854_lo_buf_o2_n_spl_0
  );


  and

  (
    g1363_p,
    g1362_p,
    g1361_p_spl_00
  );


  or

  (
    g1363_n,
    g1362_n,
    g1361_n_spl_00
  );


  and

  (
    g1364_p,
    g1359_n,
    g1357_n
  );


  or

  (
    g1364_n,
    g1359_p,
    g1357_p
  );


  and

  (
    g1365_p,
    g1364_p,
    g1363_n
  );


  or

  (
    g1365_n,
    g1364_n,
    g1363_p
  );


  and

  (
    g1366_p,
    g1309_p_spl_,
    G874_o2_n
  );


  or

  (
    g1366_n,
    g1309_n_spl_,
    G874_o2_p
  );


  and

  (
    g1367_p,
    G477_o2_n_spl_,
    G533_o2_p
  );


  or

  (
    g1367_n,
    G477_o2_p_spl_,
    G533_o2_n
  );


  and

  (
    g1368_p,
    g1366_n_spl_000,
    n2127_lo_buf_o2_p_spl_1
  );


  or

  (
    g1368_n,
    g1366_p_spl_00,
    n2127_lo_buf_o2_n_spl_
  );


  and

  (
    g1369_p,
    g1368_p,
    g1367_n_spl_00
  );


  or

  (
    g1369_n,
    g1368_n,
    g1367_p_spl_0
  );


  and

  (
    g1370_p,
    g1366_n_spl_000,
    n2187_lo_buf_o2_p_spl_
  );


  or

  (
    g1370_n,
    g1366_p_spl_00,
    n2187_lo_buf_o2_n_spl_
  );


  and

  (
    g1371_p,
    g1370_p,
    g1367_p_spl_0
  );


  or

  (
    g1371_n,
    g1370_n,
    g1367_n_spl_00
  );


  and

  (
    g1372_p,
    G1126_o2_n,
    n1893_lo_buf_o2_p_spl_00
  );


  or

  (
    g1372_n,
    G1126_o2_p,
    n1893_lo_buf_o2_n_spl_00
  );


  and

  (
    g1373_p,
    n2109_lo_buf_o2_p_spl_0,
    G851_o2_n
  );


  or

  (
    g1373_n,
    n2109_lo_buf_o2_n_spl_0,
    G851_o2_p
  );


  and

  (
    g1374_p,
    n2121_lo_buf_o2_p_spl_0,
    G1127_o2_p
  );


  or

  (
    g1374_n,
    n2121_lo_buf_o2_n_spl_0,
    G1127_o2_n
  );


  and

  (
    g1375_p,
    g1373_n,
    g1372_n
  );


  or

  (
    g1375_n,
    g1373_p,
    g1372_p
  );


  and

  (
    g1376_p,
    g1375_p,
    g1374_n
  );


  or

  (
    g1376_n,
    g1375_n,
    g1374_p
  );


  and

  (
    g1377_p,
    g1376_n,
    g1366_n_spl_00
  );


  or

  (
    g1377_n,
    g1376_p,
    g1366_p_spl_01
  );


  and

  (
    g1378_p,
    g1371_n_spl_0,
    g1369_n
  );


  or

  (
    g1378_n,
    g1371_p_spl_0,
    g1369_p
  );


  and

  (
    g1379_p,
    g1378_p,
    g1377_n
  );


  or

  (
    g1379_n,
    g1378_n,
    g1377_p
  );


  or

  (
    g1380_n,
    g1365_p_spl_00,
    n2007_lo_n_spl_00
  );


  or

  (
    g1381_n,
    g1380_n,
    g1379_n_spl_
  );


  or

  (
    g1382_n,
    g1365_p_spl_00,
    n2019_lo_n_spl_00
  );


  or

  (
    g1383_n,
    g1382_n,
    g1379_n_spl_
  );


  or

  (
    g1384_n,
    G559_o2_p,
    G565_o2_p
  );


  or

  (
    g1385_n,
    g1384_n,
    G568_o2_p
  );


  or

  (
    g1386_n,
    g1308_n,
    g1273_p_spl_0
  );


  and

  (
    g1387_p,
    g1252_p_spl_0,
    g1074_n_spl_0
  );


  or

  (
    g1388_n,
    n1761_lo_buf_o2_p_spl_0,
    n1749_lo_buf_o2_p_spl_10
  );


  or

  (
    g1389_n,
    g1388_n,
    n1773_lo_buf_o2_p_spl_0
  );


  and

  (
    g1390_p,
    G501_o2_p_spl_00,
    n1845_lo_buf_o2_n_spl_00
  );


  or

  (
    g1390_n,
    G501_o2_n_spl_01,
    n1845_lo_buf_o2_p_spl_00
  );


  and

  (
    g1391_p,
    G667_o2_p_spl_00,
    n1854_lo_buf_o2_p_spl_01
  );


  or

  (
    g1391_n,
    G667_o2_n_spl_01,
    n1854_lo_buf_o2_n_spl_1
  );


  and

  (
    g1392_p,
    g1350_p_spl_00,
    n1815_lo_buf_o2_p_spl_00
  );


  or

  (
    g1392_n,
    g1350_n_spl_00,
    n1815_lo_buf_o2_n_spl_
  );


  and

  (
    g1393_p,
    g1391_n,
    g1390_n
  );


  or

  (
    g1393_n,
    g1391_p,
    g1390_p
  );


  and

  (
    g1394_p,
    g1393_p,
    g1392_n
  );


  or

  (
    g1394_n,
    g1393_n,
    g1392_p
  );


  and

  (
    g1395_p,
    g1394_n,
    g1356_n_spl_00
  );


  or

  (
    g1395_n,
    g1394_p,
    g1356_p_spl_01
  );


  and

  (
    g1396_p,
    g1358_p_spl_00,
    n1845_lo_buf_o2_n_spl_00
  );


  or

  (
    g1396_n,
    g1358_n_spl_01,
    n1845_lo_buf_o2_p_spl_00
  );


  and

  (
    g1397_p,
    g1360_n_spl_0,
    n1845_lo_buf_o2_p_spl_01
  );


  or

  (
    g1397_n,
    g1360_p_spl_0,
    n1845_lo_buf_o2_n_spl_0
  );


  and

  (
    g1398_p,
    g1397_p,
    g1361_p_spl_00
  );


  or

  (
    g1398_n,
    g1397_n,
    g1361_n_spl_00
  );


  and

  (
    g1399_p,
    g1396_n,
    g1395_n
  );


  or

  (
    g1399_n,
    g1396_p,
    g1395_p
  );


  and

  (
    g1400_p,
    g1399_p,
    g1398_n
  );


  or

  (
    g1400_n,
    g1399_n,
    g1398_p
  );


  and

  (
    g1401_p,
    g1366_n_spl_01,
    n2121_lo_buf_o2_p_spl_1
  );


  or

  (
    g1401_n,
    g1366_p_spl_01,
    n2121_lo_buf_o2_n_spl_
  );


  and

  (
    g1402_p,
    g1401_p,
    g1367_n_spl_0
  );


  or

  (
    g1402_n,
    g1401_n,
    g1367_p_spl_1
  );


  and

  (
    g1403_p,
    G831_o2_n_spl_10,
    n1881_lo_buf_o2_p_spl_00
  );


  or

  (
    g1403_n,
    G831_o2_p_spl_1,
    n1881_lo_buf_o2_n_spl_00
  );


  and

  (
    g1404_p,
    n2094_lo_buf_o2_p_spl_0,
    G594_o2_n_spl_10
  );


  or

  (
    g1404_n,
    n2094_lo_buf_o2_n_spl_,
    G594_o2_p_spl_1
  );


  and

  (
    g1405_p,
    g1318_p_spl_01,
    n2109_lo_buf_o2_p_spl_0
  );


  or

  (
    g1405_n,
    g1318_n_spl_1,
    n2109_lo_buf_o2_n_spl_0
  );


  and

  (
    g1406_p,
    g1404_n,
    g1403_n
  );


  or

  (
    g1406_n,
    g1404_p,
    g1403_p
  );


  and

  (
    g1407_p,
    g1406_p,
    g1405_n
  );


  or

  (
    g1407_n,
    g1406_n,
    g1405_p
  );


  and

  (
    g1408_p,
    g1407_n,
    g1366_n_spl_01
  );


  or

  (
    g1408_n,
    g1407_p,
    g1366_p_spl_10
  );


  and

  (
    g1409_p,
    g1402_n,
    g1371_n_spl_0
  );


  or

  (
    g1409_n,
    g1402_p,
    g1371_p_spl_0
  );


  and

  (
    g1410_p,
    g1409_p,
    g1408_n
  );


  or

  (
    g1410_n,
    g1409_n,
    g1408_p
  );


  or

  (
    g1411_n,
    g1400_p_spl_00,
    n2007_lo_n_spl_00
  );


  or

  (
    g1412_n,
    g1411_n,
    g1410_n_spl_
  );


  or

  (
    g1413_n,
    g1400_p_spl_00,
    n2019_lo_n_spl_00
  );


  or

  (
    g1414_n,
    g1413_n,
    g1410_n_spl_
  );


  and

  (
    g1415_p,
    G791_o2_p,
    G925_o2_p
  );


  or

  (
    g1415_n,
    G791_o2_n,
    G925_o2_n
  );


  and

  (
    g1416_p,
    G1054_o2_n,
    G660_o2_n
  );


  or

  (
    g1416_n,
    G1054_o2_p,
    G660_o2_p
  );


  and

  (
    g1417_p,
    g1416_n,
    g1415_n
  );


  or

  (
    g1417_n,
    g1416_p,
    g1415_p
  );


  and

  (
    g1418_p,
    g1417_p,
    G501_o2_p_spl_01
  );


  or

  (
    g1418_n,
    g1417_n,
    G501_o2_n_spl_01
  );


  and

  (
    g1419_p,
    G667_o2_p_spl_01,
    n1893_lo_buf_o2_p_spl_00
  );


  or

  (
    g1419_n,
    G667_o2_n_spl_01,
    n1893_lo_buf_o2_n_spl_00
  );


  and

  (
    g1420_p,
    g1350_p_spl_01,
    n1854_lo_buf_o2_p_spl_10
  );


  or

  (
    g1420_n,
    g1350_n_spl_01,
    n1854_lo_buf_o2_n_spl_1
  );


  and

  (
    g1421_p,
    g1419_n,
    g1418_n
  );


  or

  (
    g1421_n,
    g1419_p,
    g1418_p
  );


  and

  (
    g1422_p,
    g1421_p,
    g1420_n
  );


  or

  (
    g1422_n,
    g1421_n,
    g1420_p
  );


  and

  (
    g1423_p,
    g1422_n,
    g1356_n_spl_01
  );


  or

  (
    g1423_n,
    g1422_p,
    g1356_p_spl_01
  );


  and

  (
    g1424_p,
    g1358_p_spl_01,
    n1881_lo_buf_o2_n_spl_00
  );


  or

  (
    g1424_n,
    g1358_n_spl_01,
    n1881_lo_buf_o2_p_spl_00
  );


  and

  (
    g1425_p,
    n1749_lo_buf_o2_n_spl_1,
    n1785_lo_buf_o2_p_spl_0
  );


  or

  (
    g1425_n,
    n1749_lo_buf_o2_p_spl_11,
    n1785_lo_buf_o2_n_spl_
  );


  and

  (
    g1426_p,
    g1425_n_spl_0,
    n1881_lo_buf_o2_p_spl_01
  );


  or

  (
    g1426_n,
    g1425_p_spl_0,
    n1881_lo_buf_o2_n_spl_01
  );


  and

  (
    g1427_p,
    g1426_p,
    g1361_p_spl_01
  );


  or

  (
    g1427_n,
    g1426_n,
    g1361_n_spl_01
  );


  and

  (
    g1428_p,
    g1424_n,
    g1423_n
  );


  or

  (
    g1428_n,
    g1424_p,
    g1423_p
  );


  and

  (
    g1429_p,
    g1428_p,
    g1427_n
  );


  or

  (
    g1429_n,
    g1428_n,
    g1427_p
  );


  and

  (
    g1430_p,
    n1869_lo_buf_o2_n_spl_00,
    n1881_lo_buf_o2_n_spl_01
  );


  or

  (
    g1430_n,
    n1869_lo_buf_o2_p_spl_00,
    n1881_lo_buf_o2_p_spl_01
  );


  and

  (
    g1431_p,
    g1430_p,
    n1893_lo_buf_o2_n_spl_01
  );


  or

  (
    g1431_n,
    g1430_n,
    n1893_lo_buf_o2_p_spl_01
  );


  and

  (
    g1432_p,
    g1431_n,
    G501_o2_p_spl_01
  );


  or

  (
    g1432_n,
    g1431_p,
    G501_o2_n_spl_10
  );


  and

  (
    g1433_p,
    G667_o2_p_spl_01,
    n1881_lo_buf_o2_n_spl_1
  );


  or

  (
    g1433_n,
    G667_o2_n_spl_10,
    n1881_lo_buf_o2_p_spl_10
  );


  and

  (
    g1434_p,
    g1350_p_spl_01,
    n1845_lo_buf_o2_n_spl_1
  );


  or

  (
    g1434_n,
    g1350_n_spl_01,
    n1845_lo_buf_o2_p_spl_01
  );


  and

  (
    g1435_p,
    g1433_n,
    g1432_n
  );


  or

  (
    g1435_n,
    g1433_p,
    g1432_p
  );


  and

  (
    g1436_p,
    g1435_p,
    g1434_n
  );


  or

  (
    g1436_n,
    g1435_n,
    g1434_p
  );


  and

  (
    g1437_p,
    g1436_n,
    g1356_n_spl_01
  );


  or

  (
    g1437_n,
    g1436_p,
    g1356_p_spl_10
  );


  and

  (
    g1438_p,
    g1358_p_spl_01,
    n1869_lo_buf_o2_n_spl_01
  );


  or

  (
    g1438_n,
    g1358_n_spl_10,
    n1869_lo_buf_o2_p_spl_01
  );


  and

  (
    g1439_p,
    g1425_n_spl_0,
    n1869_lo_buf_o2_p_spl_01
  );


  or

  (
    g1439_n,
    g1425_p_spl_0,
    n1869_lo_buf_o2_n_spl_01
  );


  and

  (
    g1440_p,
    g1439_p,
    g1361_p_spl_01
  );


  or

  (
    g1440_n,
    g1439_n,
    g1361_n_spl_01
  );


  and

  (
    g1441_p,
    g1438_n,
    g1437_n
  );


  or

  (
    g1441_n,
    g1438_p,
    g1437_p
  );


  and

  (
    g1442_p,
    g1441_p,
    g1440_n
  );


  or

  (
    g1442_n,
    g1441_n,
    g1440_p
  );


  and

  (
    g1443_p,
    g1310_n_spl_11,
    n2175_lo_p_spl_
  );


  and

  (
    g1444_p,
    g1443_p,
    g1326_n_spl_1
  );


  and

  (
    g1445_p,
    G831_o2_n_spl_10,
    n2223_lo_p_spl_
  );


  and

  (
    g1446_p,
    n2151_lo_buf_o2_p_spl_1,
    G594_o2_n_spl_10
  );


  and

  (
    g1447_p,
    g1318_p_spl_10,
    n2163_lo_p_spl_0
  );


  or

  (
    g1448_n,
    g1446_p,
    g1445_p
  );


  or

  (
    g1449_n,
    g1448_n,
    g1447_p
  );


  and

  (
    g1450_p,
    g1449_n,
    g1310_n_spl_11
  );


  or

  (
    g1451_n,
    g1444_p,
    g1329_p_spl_
  );


  or

  (
    g1452_n,
    g1451_n,
    g1450_p
  );


  and

  (
    g1453_p,
    G786_o2_p,
    G919_o2_p
  );


  or

  (
    g1453_n,
    G786_o2_n,
    G919_o2_n
  );


  and

  (
    g1454_p,
    G1052_o2_n,
    G654_o2_n
  );


  or

  (
    g1454_n,
    G1052_o2_p,
    G654_o2_p
  );


  and

  (
    g1455_p,
    g1454_n,
    g1453_n
  );


  or

  (
    g1455_n,
    g1454_p,
    g1453_p
  );


  and

  (
    g1456_p,
    g1455_p,
    G501_o2_p_spl_10
  );


  or

  (
    g1456_n,
    g1455_n,
    G501_o2_n_spl_10
  );


  and

  (
    g1457_p,
    G667_o2_p_spl_10,
    n1845_lo_buf_o2_n_spl_1
  );


  or

  (
    g1457_n,
    G667_o2_n_spl_10,
    n1845_lo_buf_o2_p_spl_10
  );


  and

  (
    g1458_p,
    g1350_p_spl_10,
    n1995_lo_p_spl_
  );


  or

  (
    g1458_n,
    g1350_n_spl_10,
    n1995_lo_n
  );


  and

  (
    g1459_p,
    g1457_n,
    g1456_n
  );


  or

  (
    g1459_n,
    g1457_p,
    g1456_p
  );


  and

  (
    g1460_p,
    g1459_p,
    g1458_n
  );


  or

  (
    g1460_n,
    g1459_n,
    g1458_p
  );


  and

  (
    g1461_p,
    g1460_n,
    g1356_n_spl_10
  );


  or

  (
    g1461_n,
    g1460_p,
    g1356_p_spl_10
  );


  and

  (
    g1462_p,
    g1358_p_spl_10,
    n1833_lo_buf_o2_n_spl_0
  );


  or

  (
    g1462_n,
    g1358_n_spl_10,
    n1833_lo_buf_o2_p_spl_00
  );


  and

  (
    g1463_p,
    g1360_n_spl_1,
    n1833_lo_buf_o2_p_spl_01
  );


  or

  (
    g1463_n,
    g1360_p_spl_,
    n1833_lo_buf_o2_n_spl_1
  );


  and

  (
    g1464_p,
    g1463_p,
    g1361_p_spl_10
  );


  or

  (
    g1464_n,
    g1463_n,
    g1361_n_spl_10
  );


  and

  (
    g1465_p,
    g1462_n,
    g1461_n
  );


  or

  (
    g1465_n,
    g1462_p,
    g1461_p
  );


  and

  (
    g1466_p,
    g1465_p,
    g1464_n
  );


  or

  (
    g1466_n,
    g1465_n,
    g1464_p
  );


  and

  (
    g1467_p,
    g1366_n_spl_10,
    n2109_lo_buf_o2_p_spl_1
  );


  or

  (
    g1467_n,
    g1366_p_spl_10,
    n2109_lo_buf_o2_n_spl_
  );


  and

  (
    g1468_p,
    g1467_p,
    g1367_n_spl_1
  );


  or

  (
    g1468_n,
    g1467_n,
    g1367_p_spl_1
  );


  and

  (
    g1469_p,
    n1869_lo_buf_o2_p_spl_10,
    G831_o2_n_spl_11
  );


  or

  (
    g1469_n,
    n1869_lo_buf_o2_n_spl_1,
    G831_o2_p_spl_1
  );


  and

  (
    g1470_p,
    n2079_lo_buf_o2_p_spl_,
    G594_o2_n_spl_11
  );


  or

  (
    g1470_n,
    n2079_lo_buf_o2_n,
    G594_o2_p_spl_1
  );


  and

  (
    g1471_p,
    g1318_p_spl_10,
    n2094_lo_buf_o2_p_spl_0
  );


  or

  (
    g1471_n,
    g1318_n_spl_1,
    n2094_lo_buf_o2_n_spl_
  );


  and

  (
    g1472_p,
    g1470_n,
    g1469_n
  );


  or

  (
    g1472_n,
    g1470_p,
    g1469_p
  );


  and

  (
    g1473_p,
    g1472_p,
    g1471_n
  );


  or

  (
    g1473_n,
    g1472_n,
    g1471_p
  );


  and

  (
    g1474_p,
    g1473_n,
    g1366_n_spl_10
  );


  or

  (
    g1474_n,
    g1473_p,
    g1366_p_spl_1
  );


  and

  (
    g1475_p,
    g1468_n,
    g1371_n_spl_
  );


  or

  (
    g1475_n,
    g1468_p,
    g1371_p_spl_1
  );


  and

  (
    g1476_p,
    g1475_p,
    g1474_n
  );


  or

  (
    g1476_n,
    g1475_n,
    g1474_p
  );


  or

  (
    g1477_n,
    g1466_p_spl_00,
    n2007_lo_n_spl_01
  );


  or

  (
    g1478_n,
    g1477_n,
    g1476_n_spl_
  );


  or

  (
    g1479_n,
    g1466_p_spl_00,
    n2019_lo_n_spl_01
  );


  or

  (
    g1480_n,
    g1479_n,
    g1476_n_spl_
  );


  or

  (
    g1481_n,
    g1389_n_spl_,
    n2055_lo_n
  );


  or

  (
    g1482_n,
    g1481_n_spl_0,
    n2307_lo_n
  );


  and

  (
    g1483_p,
    G501_o2_p_spl_10,
    n1899_lo_buf_o2_p_spl_00
  );


  or

  (
    g1483_n,
    G501_o2_n_spl_11,
    n1899_lo_buf_o2_n_spl_00
  );


  and

  (
    g1484_p,
    G667_o2_p_spl_10,
    n2199_lo_buf_o2_p_spl_0
  );


  or

  (
    g1484_n,
    G667_o2_n_spl_11,
    n2199_lo_buf_o2_n_spl_
  );


  and

  (
    g1485_p,
    g1350_p_spl_10,
    n1881_lo_buf_o2_n_spl_1
  );


  or

  (
    g1485_n,
    g1350_n_spl_10,
    n1881_lo_buf_o2_p_spl_10
  );


  and

  (
    g1486_p,
    g1484_n,
    g1483_n
  );


  or

  (
    g1486_n,
    g1484_p,
    g1483_p
  );


  and

  (
    g1487_p,
    g1486_p,
    g1485_n
  );


  or

  (
    g1487_n,
    g1486_n,
    g1485_p
  );


  and

  (
    g1488_p,
    g1487_n,
    g1356_n_spl_10
  );


  or

  (
    g1488_n,
    g1487_p,
    g1356_p_spl_11
  );


  and

  (
    g1489_p,
    g1358_p_spl_10,
    n1899_lo_buf_o2_n_spl_0
  );


  or

  (
    g1489_n,
    g1358_n_spl_11,
    n1899_lo_buf_o2_p_spl_01
  );


  and

  (
    g1490_p,
    g1425_n_spl_1,
    n1899_lo_buf_o2_p_spl_01
  );


  or

  (
    g1490_n,
    g1425_p_spl_1,
    n1899_lo_buf_o2_n_spl_1
  );


  and

  (
    g1491_p,
    g1490_p,
    g1361_p_spl_10
  );


  or

  (
    g1491_n,
    g1490_n,
    g1361_n_spl_10
  );


  and

  (
    g1492_p,
    g1489_n,
    g1488_n
  );


  or

  (
    g1492_n,
    g1489_p,
    g1488_p
  );


  and

  (
    g1493_p,
    g1492_p,
    g1491_n
  );


  or

  (
    g1493_n,
    g1492_n,
    g1491_p
  );


  and

  (
    g1494_p,
    g1383_n_spl_,
    g1381_n_spl_
  );


  and

  (
    g1495_p,
    g1365_p_spl_0,
    n2031_lo_p_spl_0
  );


  and

  (
    g1496_p,
    g1495_p,
    g1379_p_spl_
  );


  and

  (
    g1497_p,
    g1365_p_spl_1,
    n2043_lo_p_spl_0
  );


  and

  (
    g1498_p,
    g1497_p,
    g1379_p_spl_
  );


  or

  (
    g1499_n,
    g1498_p,
    g1496_p
  );


  or

  (
    g1500_n,
    g1499_n,
    g1365_n
  );


  and

  (
    g1501_p,
    g1500_n,
    g1494_p
  );


  or

  (
    g1502_n,
    g1288_n_spl_1,
    g1252_n_spl_
  );


  or

  (
    g1503_n,
    g1502_n,
    g1293_n_spl_00
  );


  or

  (
    g1504_n,
    g1503_n,
    g1055_n_spl_00
  );


  or

  (
    g1505_n,
    g1252_p_spl_0,
    n2298_lo_n_spl_00
  );


  or

  (
    g1506_n,
    g1505_n,
    g1045_n_spl_01
  );


  or

  (
    g1507_n,
    g1385_n_spl_,
    n1905_lo_buf_o2_p_spl_0
  );


  or

  (
    g1508_n,
    g1087_p_spl_0,
    g1081_n_spl_0
  );


  and

  (
    g1509_p,
    g1240_n_spl_0,
    g1083_p_spl_0
  );


  and

  (
    g1510_p,
    g1087_p_spl_0,
    g1081_n_spl_0
  );


  or

  (
    g1511_n,
    g1240_n_spl_0,
    g1083_p_spl_0
  );


  and

  (
    g1512_p,
    G1189_o2_p_spl_,
    G2232_o2_p
  );


  or

  (
    g1512_n,
    G1189_o2_n_spl_,
    G2232_o2_n
  );


  and

  (
    g1513_p,
    g1512_n_spl_,
    G2507_o2_n_spl_0
  );


  or

  (
    g1513_n,
    g1512_p_spl_0,
    G2507_o2_p_spl_0
  );


  and

  (
    g1514_p,
    g1512_p_spl_0,
    G2507_o2_p_spl_1
  );


  or

  (
    g1514_n,
    g1512_n_spl_,
    G2507_o2_n_spl_
  );


  and

  (
    g1515_p,
    g1514_n,
    g1513_n
  );


  or

  (
    g1515_n,
    g1514_p,
    g1513_p
  );


  or

  (
    g1516_n,
    g1515_p_spl_0,
    g1386_n_spl_0
  );


  or

  (
    g1517_n,
    g1516_n,
    n2298_lo_n_spl_00
  );


  or

  (
    g1518_n,
    g1386_n_spl_0,
    n2298_lo_n_spl_01
  );


  or

  (
    g1519_n,
    g1493_p_spl_,
    n2007_lo_n_spl_01
  );


  or

  (
    g1520_n,
    g1519_n,
    g1452_n_spl_00
  );


  or

  (
    g1521_n,
    g1493_p_spl_,
    n2019_lo_n_spl_01
  );


  or

  (
    g1522_n,
    g1521_n,
    g1452_n_spl_00
  );


  or

  (
    g1523_n,
    g1482_n_spl_00,
    g1365_p_spl_1
  );


  or

  (
    g1524_n,
    g1308_p_spl_,
    n2298_lo_n_spl_01
  );


  and

  (
    g1525_p,
    g1274_p_spl_0,
    g1273_p_spl_1
  );


  or

  (
    g1526_n,
    g1525_p,
    g1275_p_spl_
  );


  and

  (
    g1527_p,
    n2157_lo_buf_o2_n,
    n2145_lo_buf_o2_p_spl_
  );


  and

  (
    g1528_p,
    n2157_lo_buf_o2_p_spl_,
    n2145_lo_buf_o2_n
  );


  or

  (
    g1529_n,
    g1528_p,
    g1527_p
  );


  and

  (
    g1530_p,
    n2181_lo_buf_o2_n,
    n2169_lo_buf_o2_p_spl_
  );


  and

  (
    g1531_p,
    n2181_lo_buf_o2_p_spl_,
    n2169_lo_buf_o2_n
  );


  or

  (
    g1532_n,
    g1531_p,
    g1530_p
  );


  and

  (
    g1533_p,
    g1515_p_spl_0,
    g1276_n
  );


  and

  (
    g1534_p,
    g1515_n_spl_0,
    g1276_p_spl_
  );


  or

  (
    g1535_n,
    g1534_p,
    g1533_p
  );


  and

  (
    g1536_p,
    n1905_lo_buf_o2_p_spl_0,
    n5101_o2_n
  );


  and

  (
    g1537_p,
    n1905_lo_buf_o2_n,
    n5101_o2_p_spl_0
  );


  or

  (
    g1538_n,
    g1537_p,
    g1536_p
  );


  and

  (
    g1539_p,
    n5325_o2_n,
    n5267_o2_p_spl_0
  );


  and

  (
    g1540_p,
    n5325_o2_p_spl_0,
    n5267_o2_n
  );


  or

  (
    g1541_n,
    g1540_p,
    g1539_p
  );


  and

  (
    g1542_p,
    G1180_o2_p,
    G1725_o2_p
  );


  or

  (
    g1542_n,
    G1180_o2_n,
    G1725_o2_n
  );


  and

  (
    g1543_p,
    g1542_n_spl_,
    G2444_o2_n_spl_0
  );


  or

  (
    g1543_n,
    g1542_p_spl_0,
    G2444_o2_p_spl_0
  );


  and

  (
    g1544_p,
    g1542_p_spl_0,
    G2444_o2_p_spl_1
  );


  or

  (
    g1544_n,
    g1542_n_spl_,
    G2444_o2_n_spl_
  );


  and

  (
    g1545_p,
    g1544_n,
    g1543_n
  );


  or

  (
    g1545_n,
    g1544_p,
    g1543_p
  );


  and

  (
    g1546_p,
    g1044_n_spl_11,
    G2472_o2_p
  );


  or

  (
    g1546_n,
    g1044_p_spl_11,
    G2472_o2_n
  );


  and

  (
    g1547_p,
    g1515_n_spl_0,
    g1270_p_spl_
  );


  or

  (
    g1547_n,
    g1515_p_spl_1,
    g1270_n_spl_
  );


  and

  (
    g1548_p,
    g1515_n_spl_,
    g1273_n_spl_
  );


  or

  (
    g1548_n,
    g1515_p_spl_1,
    g1273_p_spl_1
  );


  and

  (
    g1549_p,
    g1548_p,
    g1274_n_spl_
  );


  or

  (
    g1549_n,
    g1548_n,
    g1274_p_spl_
  );


  and

  (
    g1550_p,
    g1547_n,
    g1546_n
  );


  or

  (
    g1550_n,
    g1547_p,
    g1546_p
  );


  and

  (
    g1551_p,
    g1550_p,
    g1549_n
  );


  or

  (
    g1551_n,
    g1550_n,
    g1549_p
  );


  and

  (
    g1552_p,
    g1551_p,
    g1545_n
  );


  and

  (
    g1553_p,
    g1551_n,
    g1545_p
  );


  or

  (
    g1554_n,
    g1553_p,
    g1552_p
  );


  and

  (
    g1555_p,
    n2037_lo_buf_o2_p_spl_,
    n5294_o2_p_spl_00
  );


  or

  (
    g1555_n,
    n2037_lo_buf_o2_n_spl_,
    n5294_o2_n_spl_0
  );


  and

  (
    g1556_p,
    n2025_lo_buf_o2_p_spl_,
    n5294_o2_p_spl_00
  );


  or

  (
    g1556_n,
    n2025_lo_buf_o2_n_spl_,
    n5294_o2_n_spl_0
  );


  or

  (
    g1557_n,
    g1556_p_spl_0,
    n2049_lo_buf_o2_n_spl_0
  );


  or

  (
    g1558_n,
    g1557_n_spl_,
    g1555_n_spl_0
  );


  or

  (
    g1559_n,
    g1557_n_spl_,
    g1555_p_spl_0
  );


  or

  (
    g1560_n,
    n2049_lo_buf_o2_n_spl_,
    n5294_o2_n_spl_
  );


  and

  (
    g1561_p,
    g1560_n_spl_,
    g1556_n
  );


  and

  (
    g1562_p,
    g1561_p_spl_,
    g1555_n_spl_0
  );


  or

  (
    g1563_n,
    g1560_n_spl_,
    g1556_p_spl_0
  );


  or

  (
    g1564_n,
    g1563_n_spl_,
    g1555_p_spl_0
  );


  or

  (
    g1565_n,
    g1556_p_spl_,
    n2049_lo_buf_o2_p_spl_
  );


  or

  (
    g1566_n,
    g1565_n_spl_,
    g1555_p_spl_1
  );


  and

  (
    g1567_p,
    g1561_p_spl_,
    g1555_p_spl_1
  );


  or

  (
    g1568_n,
    g1563_n_spl_,
    g1555_n_spl_1
  );


  or

  (
    g1569_n,
    g1565_n_spl_,
    g1555_n_spl_1
  );


  and

  (
    g1570_p,
    g1414_n_spl_,
    g1412_n_spl_
  );


  and

  (
    g1571_p,
    g1400_p_spl_0,
    n2031_lo_p_spl_0
  );


  and

  (
    g1572_p,
    g1571_p,
    g1410_p_spl_
  );


  and

  (
    g1573_p,
    g1400_p_spl_1,
    n2043_lo_p_spl_0
  );


  and

  (
    g1574_p,
    g1573_p,
    g1410_p_spl_
  );


  or

  (
    g1575_n,
    g1574_p,
    g1572_p
  );


  or

  (
    g1576_n,
    g1575_n,
    g1400_n
  );


  and

  (
    g1577_p,
    g1576_n,
    g1570_p
  );


  and

  (
    g1578_p,
    n1857_lo_buf_o2_n_spl_0,
    n5100_o2_n_spl_0
  );


  or

  (
    g1579_n,
    g1578_p,
    g1507_n_spl_
  );


  or

  (
    g1580_n,
    g1579_n,
    n1821_lo_buf_o2_p_spl_00
  );


  or

  (
    g1581_n,
    g1580_n,
    n5266_o2_n_spl_0
  );


  or

  (
    g1582_n,
    g1252_n_spl_,
    g1055_n_spl_0
  );


  or

  (
    g1583_n,
    g1582_n_spl_,
    g1293_n_spl_01
  );


  or

  (
    g1584_n,
    g1583_n,
    n2298_lo_n_spl_10
  );


  or

  (
    g1585_n,
    g1504_n_spl_,
    n2298_lo_n_spl_10
  );


  or

  (
    g1586_n,
    g1582_n_spl_,
    n2298_lo_n_spl_1
  );


  and

  (
    g1587_p,
    g1055_p_spl_0,
    g1045_n_spl_01
  );


  or

  (
    g1587_n,
    g1055_n_spl_1,
    g1045_p_spl_00
  );


  and

  (
    g1588_p,
    g1587_n,
    g1294_n_spl_0
  );


  or

  (
    g1588_n,
    g1587_p,
    g1294_p_spl_0
  );


  and

  (
    g1589_p,
    g1588_p,
    g1293_n_spl_01
  );


  and

  (
    g1590_p,
    g1588_n,
    g1293_p_spl_0
  );


  or

  (
    g1591_n,
    g1590_p,
    g1589_p
  );


  or

  (
    g1592_n,
    g1482_n_spl_00,
    g1400_p_spl_1
  );


  and

  (
    g1593_p,
    g1526_n_spl_0,
    g1524_n_spl_0
  );


  and

  (
    g1594_p,
    g1591_n_spl_0,
    g1586_n_spl_0
  );


  or

  (
    g1595_n,
    g1526_n_spl_0,
    g1524_n_spl_0
  );


  or

  (
    g1596_n,
    g1591_n_spl_0,
    g1586_n_spl_0
  );


  and

  (
    g1597_p,
    G501_o2_p_spl_11,
    n1893_lo_buf_o2_n_spl_01
  );


  or

  (
    g1597_n,
    G501_o2_n_spl_11,
    n1893_lo_buf_o2_p_spl_01
  );


  and

  (
    g1598_p,
    G667_o2_p_spl_11,
    n1899_lo_buf_o2_p_spl_1
  );


  or

  (
    g1598_n,
    G667_o2_n_spl_11,
    n1899_lo_buf_o2_n_spl_1
  );


  and

  (
    g1599_p,
    g1350_p_spl_11,
    n1869_lo_buf_o2_n_spl_1
  );


  or

  (
    g1599_n,
    g1350_n_spl_1,
    n1869_lo_buf_o2_p_spl_10
  );


  and

  (
    g1600_p,
    g1598_n,
    g1597_n
  );


  or

  (
    g1600_n,
    g1598_p,
    g1597_p
  );


  and

  (
    g1601_p,
    g1600_p,
    g1599_n
  );


  or

  (
    g1601_n,
    g1600_n,
    g1599_p
  );


  and

  (
    g1602_p,
    g1601_n,
    g1356_n_spl_11
  );


  or

  (
    g1602_n,
    g1601_p,
    g1356_p_spl_11
  );


  and

  (
    g1603_p,
    g1358_p_spl_11,
    n1893_lo_buf_o2_n_spl_1
  );


  or

  (
    g1603_n,
    g1358_n_spl_11,
    n1893_lo_buf_o2_p_spl_10
  );


  and

  (
    g1604_p,
    g1425_n_spl_1,
    n1893_lo_buf_o2_p_spl_10
  );


  or

  (
    g1604_n,
    g1425_p_spl_1,
    n1893_lo_buf_o2_n_spl_1
  );


  and

  (
    g1605_p,
    g1604_p,
    g1361_p_spl_11
  );


  or

  (
    g1605_n,
    g1604_n,
    g1361_n_spl_1
  );


  and

  (
    g1606_p,
    g1603_n,
    g1602_n
  );


  or

  (
    g1606_n,
    g1603_p,
    g1602_p
  );


  and

  (
    g1607_p,
    g1606_p,
    g1605_n
  );


  or

  (
    g1607_n,
    g1606_n,
    g1605_p
  );


  and

  (
    g1608_p,
    g1607_n_spl_0,
    n2007_lo_p_spl_0
  );


  or

  (
    g1608_n,
    g1607_p_spl_0,
    n2007_lo_n_spl_1
  );


  and

  (
    g1609_p,
    g1608_p,
    g1347_p_spl_
  );


  or

  (
    g1609_n,
    g1608_n,
    g1347_n_spl_00
  );


  and

  (
    g1610_p,
    g1607_n_spl_0,
    n2019_lo_p_spl_00
  );


  or

  (
    g1610_n,
    g1607_p_spl_0,
    n2019_lo_n_spl_1
  );


  and

  (
    g1611_p,
    g1610_p,
    g1347_p_spl_
  );


  or

  (
    g1611_n,
    g1610_n,
    g1347_n_spl_00
  );


  and

  (
    g1612_p,
    g1611_n,
    g1609_n
  );


  or

  (
    g1612_n,
    g1611_p,
    g1609_p
  );


  and

  (
    g1613_p,
    g1429_n_spl_00,
    n2007_lo_p_spl_0
  );


  or

  (
    g1613_n,
    g1429_p_spl_0,
    n2007_lo_n_spl_1
  );


  and

  (
    g1614_p,
    g1613_p,
    g1337_p_spl_
  );


  or

  (
    g1614_n,
    g1613_n,
    g1337_n_spl_00
  );


  and

  (
    g1615_p,
    g1429_n_spl_00,
    n2019_lo_p_spl_00
  );


  or

  (
    g1615_n,
    g1429_p_spl_0,
    n2019_lo_n_spl_1
  );


  and

  (
    g1616_p,
    g1615_p,
    g1337_p_spl_
  );


  or

  (
    g1616_n,
    g1615_n,
    g1337_n_spl_00
  );


  and

  (
    g1617_p,
    g1616_n,
    g1614_n
  );


  or

  (
    g1617_n,
    g1616_p,
    g1614_p
  );


  or

  (
    g1618_n,
    n5293_o2_p_spl_,
    n5292_o2_p_spl_0
  );


  or

  (
    g1619_n,
    g1618_n,
    n5294_o2_p_spl_0
  );


  or

  (
    g1620_n,
    n5266_o2_p_spl_00,
    n5100_o2_p_spl_00
  );


  and

  (
    g1621_p,
    g1620_n,
    n1821_lo_buf_o2_n_spl_0
  );


  and

  (
    g1622_p,
    g1506_n_spl_,
    g1045_n_spl_1
  );


  and

  (
    g1623_p,
    g1387_p_spl_,
    n2298_lo_p_spl_
  );


  and

  (
    g1624_p,
    g1623_p,
    g1284_n_spl_
  );


  and

  (
    g1625_p,
    g1522_n_spl_,
    g1520_n_spl_
  );


  and

  (
    g1626_p,
    g1294_n_spl_,
    g1293_p_spl_1
  );


  or

  (
    g1626_n,
    g1294_p_spl_,
    g1293_n_spl_1
  );


  and

  (
    g1627_p,
    g1293_p_spl_1,
    g1055_p_spl_1
  );


  or

  (
    g1627_n,
    g1293_n_spl_1,
    g1055_n_spl_1
  );


  and

  (
    g1628_p,
    g1627_p,
    g1045_n_spl_1
  );


  or

  (
    g1628_n,
    g1627_n,
    g1045_p_spl_0
  );


  and

  (
    g1629_p,
    g1626_n,
    g1289_n_spl_
  );


  or

  (
    g1629_n,
    g1626_p,
    g1289_p_spl_
  );


  and

  (
    g1630_p,
    g1629_p,
    g1628_n
  );


  or

  (
    g1630_n,
    g1629_n,
    g1628_p
  );


  and

  (
    g1631_p,
    g1630_p,
    g1288_p_spl_
  );


  and

  (
    g1632_p,
    g1630_n,
    g1288_n_spl_1
  );


  or

  (
    g1633_n,
    g1632_p,
    g1631_p
  );


  and

  (
    g1634_p,
    n1857_lo_buf_o2_p_spl_00,
    n5100_o2_n_spl_0
  );


  or

  (
    g1634_n,
    n1857_lo_buf_o2_n_spl_0,
    n5100_o2_p_spl_00
  );


  and

  (
    g1635_p,
    n1857_lo_buf_o2_n_spl_,
    n5100_o2_p_spl_01
  );


  or

  (
    g1635_n,
    n1857_lo_buf_o2_p_spl_00,
    n5100_o2_n_spl_
  );


  and

  (
    g1636_p,
    g1635_n,
    g1634_n
  );


  or

  (
    g1636_n,
    g1635_p,
    g1634_p
  );


  and

  (
    g1637_p,
    n1821_lo_buf_o2_p_spl_00,
    n5266_o2_p_spl_00
  );


  or

  (
    g1637_n,
    n1821_lo_buf_o2_n_spl_0,
    n5266_o2_n_spl_0
  );


  and

  (
    g1638_p,
    n1821_lo_buf_o2_n_spl_,
    n5266_o2_n_spl_
  );


  or

  (
    g1638_n,
    n1821_lo_buf_o2_p_spl_0,
    n5266_o2_p_spl_01
  );


  and

  (
    g1639_p,
    g1638_n,
    g1637_n
  );


  or

  (
    g1639_n,
    g1638_p,
    g1637_p
  );


  or

  (
    g1640_n,
    g1639_n,
    g1636_p
  );


  or

  (
    g1641_n,
    g1639_p,
    g1636_n
  );


  and

  (
    g1642_p,
    g1641_n,
    g1640_n
  );


  and

  (
    g1643_p,
    g1079_n_spl_,
    g1071_n_spl_0
  );


  or

  (
    g1643_n,
    g1079_p_spl_0,
    g1071_p_spl_01
  );


  and

  (
    g1644_p,
    g1079_p_spl_0,
    g1071_p_spl_1
  );


  or

  (
    g1644_n,
    g1079_n_spl_,
    g1071_n_spl_
  );


  and

  (
    g1645_p,
    g1644_n,
    g1643_n
  );


  or

  (
    g1645_n,
    g1644_p,
    g1643_p
  );


  and

  (
    g1646_p,
    g1645_n,
    g1301_n_spl_
  );


  and

  (
    g1647_p,
    g1645_p,
    g1301_p
  );


  or

  (
    g1648_n,
    g1647_p,
    g1646_p
  );


  and

  (
    g1649_p,
    g1282_p,
    g1279_n_spl_
  );


  and

  (
    g1650_p,
    g1282_n_spl_,
    g1279_p
  );


  or

  (
    g1651_n,
    g1650_p,
    g1649_p
  );


  and

  (
    g1652_p,
    g1442_n_spl_00,
    n2007_lo_p_spl_1
  );


  and

  (
    g1653_p,
    g1652_p,
    g1324_p_spl_
  );


  and

  (
    g1654_p,
    g1442_n_spl_00,
    n2019_lo_p_spl_0
  );


  and

  (
    g1655_p,
    g1654_p,
    g1324_p_spl_
  );


  or

  (
    g1656_n,
    g1655_p,
    g1653_p
  );


  or

  (
    g1657_n,
    g1442_n_spl_0,
    n2031_lo_n_spl_0
  );


  or

  (
    g1658_n,
    g1657_n,
    g1324_n_spl_0
  );


  or

  (
    g1659_n,
    g1442_n_spl_1,
    n2043_lo_n_spl_0
  );


  or

  (
    g1660_n,
    g1659_n,
    g1324_n_spl_0
  );


  and

  (
    g1661_p,
    g1660_n,
    g1658_n
  );


  and

  (
    g1662_p,
    g1661_p,
    g1442_p
  );


  or

  (
    g1663_n,
    g1662_p,
    g1656_n_spl_
  );


  or

  (
    g1664_n,
    g1607_n_spl_1,
    n2031_lo_n_spl_0
  );


  or

  (
    g1665_n,
    g1664_n,
    g1347_n_spl_0
  );


  or

  (
    g1666_n,
    g1607_n_spl_1,
    n2043_lo_n_spl_0
  );


  or

  (
    g1667_n,
    g1666_n,
    g1347_n_spl_1
  );


  and

  (
    g1668_p,
    g1667_n,
    g1665_n
  );


  and

  (
    g1669_p,
    g1668_p,
    g1607_p_spl_1
  );


  or

  (
    g1670_n,
    g1669_p,
    g1612_n_spl_
  );


  and

  (
    g1671_p,
    g1480_n_spl_,
    g1478_n_spl_
  );


  and

  (
    g1672_p,
    g1466_p_spl_0,
    n2031_lo_p_spl_1
  );


  and

  (
    g1673_p,
    g1672_p,
    g1476_p_spl_
  );


  and

  (
    g1674_p,
    g1466_p_spl_1,
    n2043_lo_p_spl_1
  );


  and

  (
    g1675_p,
    g1674_p,
    g1476_p_spl_
  );


  or

  (
    g1676_n,
    g1675_p,
    g1673_p
  );


  or

  (
    g1677_n,
    g1676_n,
    g1466_n
  );


  and

  (
    g1678_p,
    g1677_n,
    g1671_p
  );


  or

  (
    g1679_n,
    g1429_n_spl_0,
    n2031_lo_n_spl_1
  );


  or

  (
    g1680_n,
    g1679_n,
    g1337_n_spl_0
  );


  or

  (
    g1681_n,
    g1429_n_spl_1,
    n2043_lo_n_spl_1
  );


  or

  (
    g1682_n,
    g1681_n,
    g1337_n_spl_1
  );


  and

  (
    g1683_p,
    g1682_n,
    g1680_n
  );


  and

  (
    g1684_p,
    g1683_p,
    g1429_p_spl_
  );


  or

  (
    g1685_n,
    g1684_p,
    g1617_n_spl_
  );


  or

  (
    g1686_n,
    g1493_n_spl_0,
    n2031_lo_n_spl_1
  );


  or

  (
    g1687_n,
    g1686_n,
    g1452_n_spl_0
  );


  or

  (
    g1688_n,
    g1493_n_spl_0,
    n2043_lo_n_spl_1
  );


  or

  (
    g1689_n,
    g1688_n,
    g1452_n_spl_1
  );


  or

  (
    g1690_n,
    g1607_p_spl_1,
    g1482_n_spl_0
  );


  or

  (
    g1691_n,
    g1481_n_spl_0,
    g1466_p_spl_1
  );


  and

  (
    g1692_p,
    G5_p_spl_0,
    G4_p_spl_00
  );


  or

  (
    g1693_n,
    G49_p,
    G4_p_spl_00
  );


  or

  (
    g1694_n,
    n1815_lo_buf_o2_p_spl_00,
    n1833_lo_buf_o2_p_spl_01
  );


  or

  (
    g1695_n,
    g1694_n,
    n1845_lo_buf_o2_p_spl_10
  );


  and

  (
    g1696_p,
    g1695_n,
    G501_o2_p_spl_11
  );


  and

  (
    g1697_p,
    G667_o2_p_spl_11,
    n1833_lo_buf_o2_n_spl_1
  );


  and

  (
    g1698_p,
    g1350_p_spl_11,
    n1983_lo_p_spl_
  );


  or

  (
    g1699_n,
    g1697_p,
    g1696_p
  );


  or

  (
    g1700_n,
    g1699_n,
    g1698_p
  );


  and

  (
    g1701_p,
    g1700_n,
    g1356_n_spl_11
  );


  and

  (
    g1702_p,
    g1358_p_spl_11,
    n1815_lo_buf_o2_n_spl_
  );


  and

  (
    g1703_p,
    g1360_n_spl_1,
    n1815_lo_buf_o2_p_spl_0
  );


  and

  (
    g1704_p,
    g1703_p,
    g1361_p_spl_11
  );


  or

  (
    g1705_n,
    g1702_p,
    g1701_p
  );


  or

  (
    g1706_n,
    g1705_n,
    g1704_p
  );


  or

  (
    g1707_n,
    g1685_n_spl_0,
    g1663_n_spl_0
  );


  or

  (
    g1708_n,
    g1707_n,
    g1612_p
  );


  or

  (
    g1709_n,
    g1663_n_spl_0,
    g1617_p
  );


  and

  (
    g1710_p,
    g1366_n_spl_11,
    n2094_lo_buf_o2_p_spl_1
  );


  and

  (
    g1711_p,
    g1710_p,
    g1367_n_spl_1
  );


  and

  (
    g1712_p,
    n1854_lo_buf_o2_p_spl_10,
    G831_o2_n_spl_11
  );


  and

  (
    g1713_p,
    G594_o2_n_spl_11,
    n2067_lo_p
  );


  and

  (
    g1714_p,
    g1318_p_spl_1,
    n2079_lo_buf_o2_p_spl_
  );


  or

  (
    g1715_n,
    g1713_p,
    g1712_p
  );


  or

  (
    g1716_n,
    g1715_n,
    g1714_p
  );


  and

  (
    g1717_p,
    g1716_n,
    g1366_n_spl_11
  );


  or

  (
    g1718_n,
    g1711_p,
    g1371_p_spl_1
  );


  or

  (
    g1719_n,
    g1718_n,
    g1717_p
  );


  or

  (
    g1720_n,
    g1685_n_spl_0,
    g1625_p_spl_
  );


  or

  (
    g1721_n,
    g1720_n,
    g1670_n_spl_0
  );


  or

  (
    g1722_n,
    g1721_n,
    g1663_n_spl_1
  );


  or

  (
    g1723_n,
    G6_p_spl_,
    G5_p_spl_0
  );


  and

  (
    g1724_p,
    G4_p_spl_01,
    G3_n
  );


  and

  (
    g1725_p,
    g1693_n_spl_0,
    G4_p_spl_01
  );


  and

  (
    g1726_p,
    G3_p_spl_0,
    G2_p_spl_
  );


  buf

  (
    G3519,
    g582_p
  );


  buf

  (
    G3520,
    g583_n
  );


  buf

  (
    G3521,
    g610_p
  );


  buf

  (
    G3522,
    g616_p
  );


  buf

  (
    G3523,
    g619_n
  );


  buf

  (
    G3524,
    g620_p
  );


  buf

  (
    G3525,
    g622_n
  );


  buf

  (
    G3526,
    g624_p
  );


  buf

  (
    G3527,
    g631_n
  );


  buf

  (
    G3528,
    g634_p
  );


  buf

  (
    G3529,
    g637_p
  );


  buf

  (
    G3530,
    g664_n
  );


  buf

  (
    G3531,
    g667_p
  );


  buf

  (
    G3532,
    g670_p
  );


  buf

  (
    G3533,
    g673_p
  );


  buf

  (
    G3534,
    G3312_o2_p
  );


  buf

  (
    G3535,
    G3332_o2_p
  );


  buf

  (
    G3536,
    g676_p
  );


  buf

  (
    G3537,
    g687_n_spl_
  );


  not

  (
    G3538,
    g692_p
  );


  buf

  (
    G3539,
    g724_n
  );


  buf

  (
    G3540,
    g733_p
  );


  buf

  (
    n1836_li,
    n4377_o2_p
  );


  buf

  (
    n1872_li,
    n4454_o2_p_spl_
  );


  buf

  (
    n1884_li,
    n4378_o2_p
  );


  buf

  (
    n1911_li,
    G15_p
  );


  buf

  (
    n1914_li,
    n1911_lo_p
  );


  buf

  (
    n1917_li,
    n1914_lo_p
  );


  buf

  (
    n1923_li,
    G16_p
  );


  buf

  (
    n1926_li,
    n1923_lo_p
  );


  buf

  (
    n1929_li,
    n1926_lo_p
  );


  buf

  (
    n1935_li,
    G17_p
  );


  buf

  (
    n1938_li,
    n1935_lo_p
  );


  buf

  (
    n1947_li,
    G18_p
  );


  buf

  (
    n1950_li,
    n1947_lo_p
  );


  buf

  (
    n1959_li,
    G19_p
  );


  buf

  (
    n1962_li,
    n1959_lo_p
  );


  buf

  (
    n1971_li,
    G20_p
  );


  buf

  (
    n1974_li,
    n1971_lo_p
  );


  buf

  (
    n1983_li,
    G21_p
  );


  buf

  (
    n1995_li,
    G22_p
  );


  buf

  (
    n2007_li,
    G23_p
  );


  buf

  (
    n2019_li,
    G24_p
  );


  buf

  (
    n2031_li,
    G25_p
  );


  buf

  (
    n2043_li,
    G26_p
  );


  buf

  (
    n2055_li,
    G27_p
  );


  buf

  (
    n2064_li,
    n4920_o2_p_spl_0
  );


  buf

  (
    n2067_li,
    G28_p
  );


  buf

  (
    n2100_li,
    n4505_o2_p
  );


  buf

  (
    n2112_li,
    n4455_o2_p
  );


  buf

  (
    n2124_li,
    n4456_o2_p
  );


  buf

  (
    n2136_li,
    n4567_o2_p
  );


  buf

  (
    n2148_li,
    n4568_o2_p
  );


  buf

  (
    n2160_li,
    n4569_o2_p
  );


  buf

  (
    n2163_li,
    G36_p
  );


  buf

  (
    n2172_li,
    n4652_o2_p
  );


  buf

  (
    n2175_li,
    G37_p
  );


  buf

  (
    n2184_li,
    n4787_o2_p
  );


  buf

  (
    n2223_li,
    G41_p
  );


  buf

  (
    n2235_li,
    G42_p
  );


  buf

  (
    n2238_li,
    n2235_lo_p
  );


  buf

  (
    n2247_li,
    G43_p
  );


  buf

  (
    n2250_li,
    n2247_lo_p
  );


  buf

  (
    n2259_li,
    G44_p
  );


  buf

  (
    n2262_li,
    n2259_lo_p
  );


  buf

  (
    n2271_li,
    G45_p
  );


  buf

  (
    n2274_li,
    n2271_lo_p
  );


  buf

  (
    n2283_li,
    G46_p
  );


  buf

  (
    n2286_li,
    n2283_lo_p
  );


  buf

  (
    n2295_li,
    G47_p
  );


  buf

  (
    n2298_li,
    n2295_lo_p
  );


  buf

  (
    n2304_li,
    n2301_lo_buf_o2_p_spl_
  );


  buf

  (
    n2307_li,
    G48_p
  );


  buf

  (
    n2331_li,
    G50_p
  );


  buf

  (
    n2334_li,
    n2331_lo_p
  );


  buf

  (
    n2337_li,
    n2334_lo_p
  );


  buf

  (
    n2340_li,
    n2337_lo_p
  );


  buf

  (
    n3241_i2,
    n327_inv_p
  );


  buf

  (
    n3242_i2,
    n330_inv_p
  );


  buf

  (
    n3610_i2,
    n399_inv_p
  );


  buf

  (
    n3980_i2,
    n435_inv_p
  );


  buf

  (
    n3968_i2,
    n426_inv_p
  );


  buf

  (
    n4298_i2,
    G2610_o2_p
  );


  buf

  (
    n4371_i2,
    G2558_o2_p
  );


  buf

  (
    n4413_i2,
    n570_inv_p
  );


  buf

  (
    n4418_i2,
    G2552_o2_p
  );


  buf

  (
    n4628_i2,
    G2607_o2_p
  );


  buf

  (
    n4629_i2,
    n702_inv_p
  );


  buf

  (
    n4633_i2,
    G1005_o2_p
  );


  buf

  (
    n4634_i2,
    G1008_o2_p
  );


  buf

  (
    n4732_i2,
    n723_inv_p
  );


  buf

  (
    n4733_i2,
    G2947_o2_p
  );


  buf

  (
    n4884_i2,
    n786_inv_p
  );


  buf

  (
    n4886_i2,
    n789_inv_p
  );


  buf

  (
    n4890_i2,
    G2823_o2_p
  );


  buf

  (
    n5011_i2,
    n849_inv_p_spl_
  );


  buf

  (
    n5012_i2,
    n852_inv_p_spl_1
  );


  buf

  (
    n5013_i2,
    n855_inv_p_spl_
  );


  buf

  (
    n5014_i2,
    n858_inv_p_spl_1
  );


  buf

  (
    n5015_i2,
    n861_inv_p
  );


  buf

  (
    n5021_i2,
    G2833_o2_p
  );


  buf

  (
    n5016_i2,
    G2805_o2_p
  );


  buf

  (
    n5026_i2,
    n873_inv_p
  );


  buf

  (
    n4377_i2,
    n5266_o2_p_spl_01
  );


  buf

  (
    n4378_i2,
    n5267_o2_p_spl_0
  );


  buf

  (
    n4389_i2,
    n537_inv_p
  );


  buf

  (
    n4390_i2,
    n540_inv_p
  );


  buf

  (
    n4391_i2,
    n543_inv_p
  );


  buf

  (
    n4398_i2,
    n5292_o2_p_spl_0
  );


  buf

  (
    n4401_i2,
    n5295_o2_p_spl_00
  );


  buf

  (
    n5117_i2,
    n1056_inv_p_spl_1
  );


  buf

  (
    n5115_i2,
    n1050_inv_p_spl_1
  );


  buf

  (
    n5122_i2,
    n1071_inv_p_spl_1
  );


  buf

  (
    n5121_i2,
    n1068_inv_p_spl_1
  );


  buf

  (
    n5119_i2,
    n1062_inv_p_spl_1
  );


  buf

  (
    n5116_i2,
    n1053_inv_p_spl_1
  );


  buf

  (
    n5123_i2,
    n1074_inv_p_spl_1
  );


  buf

  (
    n5156_i2,
    G935_o2_p_spl_
  );


  buf

  (
    n5167_i2,
    n1176_inv_p
  );


  buf

  (
    n4454_i2,
    n5325_o2_p_spl_0
  );


  buf

  (
    n4455_i2,
    n5326_o2_p_spl_
  );


  buf

  (
    n4456_i2,
    n5327_o2_p_spl_
  );


  buf

  (
    n4505_i2,
    n2097_lo_buf_o2_p_spl_
  );


  buf

  (
    G742_i2,
    n429_inv_p_spl_
  );


  buf

  (
    G727_i2,
    g734_n_spl_
  );


  buf

  (
    n4567_i2,
    n2133_lo_buf_o2_p_spl_
  );


  buf

  (
    n4568_i2,
    n2145_lo_buf_o2_p_spl_
  );


  buf

  (
    n4569_i2,
    n2157_lo_buf_o2_p_spl_
  );


  buf

  (
    n4571_i2,
    n2205_lo_buf_o2_p
  );


  buf

  (
    n4572_i2,
    n2217_lo_buf_o2_p
  );


  buf

  (
    n4537_i2,
    n642_inv_p
  );


  buf

  (
    n4539_i2,
    n648_inv_p
  );


  buf

  (
    n4651_i2,
    n2001_lo_buf_o2_p
  );


  buf

  (
    n4652_i2,
    n2169_lo_buf_o2_p_spl_
  );


  buf

  (
    n4653_i2,
    n2229_lo_buf_o2_p
  );


  buf

  (
    G1514_i2,
    g737_n_spl_
  );


  not

  (
    G1823_i2,
    g740_p_spl_
  );


  buf

  (
    n4783_i2,
    n2013_lo_buf_o2_p_spl_
  );


  buf

  (
    n4787_i2,
    n2181_lo_buf_o2_p_spl_
  );


  buf

  (
    n4808_i2,
    n744_inv_p
  );


  buf

  (
    n4815_i2,
    n747_inv_p
  );


  buf

  (
    n4816_i2,
    n750_inv_p
  );


  buf

  (
    n4822_i2,
    n753_inv_p
  );


  buf

  (
    G572_i2,
    n4398_o2_p_spl_
  );


  buf

  (
    n4919_i2,
    n1989_lo_buf_o2_p
  );


  buf

  (
    n4920_i2,
    n2061_lo_buf_o2_p_spl_
  );


  buf

  (
    n4921_i2,
    n2313_lo_buf_o2_p_spl_
  );


  buf

  (
    G1048_i2,
    g743_p_spl_11
  );


  buf

  (
    n5041_i2,
    G2021_o2_p
  );


  buf

  (
    n5094_i2,
    n1008_inv_p
  );


  buf

  (
    n5278_i2,
    G2393_o2_p_spl_
  );


  buf

  (
    n5301_i2,
    n1557_inv_p_spl_
  );


  buf

  (
    G2610_i2,
    g746_n_spl_
  );


  buf

  (
    G3174_i2,
    g753_p_spl_
  );


  not

  (
    G3146_i2,
    g757_n_spl_
  );


  not

  (
    G3217_i2,
    g761_n_spl_
  );


  not

  (
    G3220_i2,
    g765_n_spl_
  );


  not

  (
    G2839_i2,
    g813_n_spl_
  );


  not

  (
    G3251_i2,
    g822_n_spl_
  );


  buf

  (
    G3042_i2,
    g826_p_spl_
  );


  not

  (
    G3045_i2,
    g827_p_spl_
  );


  buf

  (
    G3262_i2,
    g832_p_spl_
  );


  not

  (
    G2845_i2,
    g884_n_spl_
  );


  buf

  (
    G2929_i2,
    g930_p_spl_
  );


  not

  (
    G2848_i2,
    g981_n_spl_
  );


  buf

  (
    G2851_i2,
    g1032_p_spl_
  );


  not

  (
    G3291_i2,
    g1037_n_spl_
  );


  not

  (
    G3254_i2,
    g1042_n_spl_
  );


  buf

  (
    G2666_i2,
    g1045_p_spl_1
  );


  buf

  (
    n5099_i2,
    n1785_lo_buf_o2_p_spl_
  );


  buf

  (
    n5100_i2,
    n1845_lo_buf_o2_p_spl_11
  );


  buf

  (
    n5101_i2,
    n1893_lo_buf_o2_p_spl_11
  );


  buf

  (
    G2558_i2,
    g1052_p_spl_
  );


  buf

  (
    n5266_i2,
    n1833_lo_buf_o2_p_spl_1
  );


  buf

  (
    n5267_i2,
    n1881_lo_buf_o2_p_spl_11
  );


  buf

  (
    G2759_i2,
    g1055_p_spl_1
  );


  buf

  (
    n5269_i2,
    n1479_inv_p
  );


  buf

  (
    n5270_i2,
    n1482_inv_p
  );


  buf

  (
    n5271_i2,
    n1485_inv_p
  );


  buf

  (
    n5292_i2,
    n1749_lo_buf_o2_p_spl_11
  );


  buf

  (
    n5293_i2,
    n1761_lo_buf_o2_p_spl_1
  );


  buf

  (
    n5294_i2,
    n1773_lo_buf_o2_p_spl_1
  );


  buf

  (
    n5295_i2,
    n1809_lo_buf_o2_p_spl_
  );


  buf

  (
    G618_i2,
    n4920_o2_p_spl_
  );


  buf

  (
    G621_i2,
    n4921_o2_p_spl_
  );


  buf

  (
    G384_i2,
    n5100_o2_p_spl_01
  );


  buf

  (
    G377_i2,
    n5266_o2_p_spl_1
  );


  buf

  (
    G400_i2,
    n1857_lo_buf_o2_p_spl_0
  );


  not

  (
    G3171_i2,
    g1059_n_spl_
  );


  not

  (
    G2552_i2,
    g1074_n_spl_
  );


  not

  (
    G3272_i2,
    g1078_n_spl_
  );


  buf

  (
    G2015_i2,
    g1079_p_spl_
  );


  buf

  (
    G3294_i2,
    g1081_n_spl_
  );


  not

  (
    G3281_i2,
    g1083_p_spl_
  );


  not

  (
    G3320_i2,
    g1085_p_spl_0
  );


  not

  (
    G3275_i2,
    g1087_p_spl_
  );


  not

  (
    G3140_i2,
    g1095_n_spl_
  );


  not

  (
    G2836_i2,
    g1142_n_spl_
  );


  not

  (
    G2926_i2,
    g1184_n_spl_
  );


  not

  (
    G2842_i2,
    g1226_n_spl_
  );


  not

  (
    G3302_i2,
    g1232_n_spl_
  );


  not

  (
    G3288_i2,
    g1237_n_spl_
  );


  not

  (
    G3143_i2,
    g1238_n_spl_
  );


  not

  (
    G3100_i2,
    g1240_n_spl_
  );


  buf

  (
    G2512_i2,
    g1071_p_spl_1
  );


  buf

  (
    n5325_i2,
    n1869_lo_buf_o2_p_spl_11
  );


  buf

  (
    n5326_i2,
    n2109_lo_buf_o2_p_spl_1
  );


  buf

  (
    n5327_i2,
    n2121_lo_buf_o2_p_spl_1
  );


  buf

  (
    n1857_lo_buf_i2,
    n1854_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2097_lo_buf_i2,
    n2094_lo_buf_o2_p_spl_1
  );


  buf

  (
    G2669_i2,
    g1252_p_spl_
  );


  buf

  (
    G552_i2,
    n1845_lo_buf_o2_p_spl_11
  );


  buf

  (
    G568_i2,
    n1893_lo_buf_o2_p_spl_11
  );


  buf

  (
    G530_i2,
    n1797_lo_buf_o2_p_spl_
  );


  buf

  (
    G565_i2,
    n1881_lo_buf_o2_p_spl_11
  );


  buf

  (
    G559_i2,
    n1869_lo_buf_o2_p_spl_11
  );


  buf

  (
    n1821_lo_buf_i2,
    n1815_lo_buf_o2_p_spl_1
  );


  buf

  (
    n1905_lo_buf_i2,
    n1899_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2133_lo_buf_i2,
    n2127_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2145_lo_buf_i2,
    n2139_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2157_lo_buf_i2,
    n2151_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2205_lo_buf_i2,
    n2199_lo_buf_o2_p_spl_
  );


  buf

  (
    n2217_lo_buf_i2,
    n2211_lo_buf_o2_p_spl_
  );


  buf

  (
    G447_i2,
    n5101_o2_p_spl_0
  );


  buf

  (
    G434_i2,
    n5267_o2_p_spl_1
  );


  buf

  (
    G422_i2,
    n5325_o2_p_spl_1
  );


  buf

  (
    G461_i2,
    n1905_lo_buf_o2_p_spl_1
  );


  not

  (
    G3312_i2,
    g1254_p_spl_0
  );


  not

  (
    G3332_i2,
    g1256_p_spl_0
  );


  not

  (
    G3195_i2,
    g1258_p_spl_0
  );


  buf

  (
    G2607_i2,
    g1269_n_spl_
  );


  buf

  (
    G2799_i2,
    g1276_p_spl_
  );


  buf

  (
    G1005_i2,
    g1279_n_spl_
  );


  buf

  (
    G1008_i2,
    g1282_n_spl_
  );


  buf

  (
    n2001_lo_buf_i2,
    n1995_lo_p_spl_
  );


  buf

  (
    n2169_lo_buf_i2,
    n2163_lo_p_spl_
  );


  buf

  (
    n2229_lo_buf_i2,
    n2223_lo_p_spl_
  );


  buf

  (
    n2301_lo_buf_i2,
    n2298_lo_p_spl_
  );


  not

  (
    G2816_i2,
    g1284_n_spl_
  );


  buf

  (
    G2947_i2,
    g1301_n_spl_
  );


  buf

  (
    n2013_lo_buf_i2,
    n2007_lo_p_spl_1
  );


  buf

  (
    n2025_lo_buf_i2,
    n2019_lo_p_spl_1
  );


  buf

  (
    n2037_lo_buf_i2,
    n2031_lo_p_spl_1
  );


  buf

  (
    n2049_lo_buf_i2,
    n2043_lo_p_spl_1
  );


  buf

  (
    n2181_lo_buf_i2,
    n2175_lo_p_spl_
  );


  buf

  (
    G546_i2,
    n1833_lo_buf_o2_p_spl_1
  );


  buf

  (
    G480_i2,
    n1761_lo_buf_o2_p_spl_1
  );


  buf

  (
    G492_i2,
    n1773_lo_buf_o2_p_spl_1
  );


  buf

  (
    G540_i2,
    n1815_lo_buf_o2_p_spl_1
  );


  not

  (
    G3350_i2,
    g1303_n_spl_
  );


  not

  (
    G3360_i2,
    g1304_n_spl_
  );


  not

  (
    G3373_i2,
    g1085_p_spl_0
  );


  not

  (
    G3237_i2,
    g1258_p_spl_0
  );


  buf

  (
    G2773_i2,
    g1308_p_spl_
  );


  buf

  (
    G1733_i2,
    g1324_n_spl_
  );


  buf

  (
    G1738_i2,
    g1337_n_spl_1
  );


  buf

  (
    G1751_i2,
    g1347_n_spl_1
  );


  not

  (
    G2216_i2,
    g1381_n_spl_
  );


  not

  (
    G2219_i2,
    g1383_n_spl_
  );


  buf

  (
    G381_i2,
    n5100_o2_p_spl_1
  );


  buf

  (
    G397_i2,
    n1857_lo_buf_o2_p_spl_1
  );


  buf

  (
    G787_i2,
    g1385_n_spl_
  );


  not

  (
    G2823_i2,
    g1386_n_spl_
  );


  buf

  (
    G2796_i2,
    g1387_p_spl_
  );


  buf

  (
    G875_i2,
    g1389_n_spl_
  );


  not

  (
    G2208_i2,
    g1412_n_spl_
  );


  not

  (
    G2211_i2,
    g1414_n_spl_
  );


  buf

  (
    n1989_lo_buf_i2,
    n1983_lo_p_spl_
  );


  buf

  (
    n2061_lo_buf_i2,
    n2055_lo_p
  );


  buf

  (
    n2313_lo_buf_i2,
    n2307_lo_p
  );


  buf

  (
    G2232_i2,
    g1429_n_spl_1
  );


  buf

  (
    G1725_i2,
    g1442_n_spl_1
  );


  buf

  (
    G1764_i2,
    g1452_n_spl_1
  );


  not

  (
    G2356_i2,
    g1478_n_spl_
  );


  not

  (
    G2359_i2,
    g1480_n_spl_
  );


  not

  (
    G1180_i2,
    g1482_n_spl_1
  );


  buf

  (
    G1756_i2,
    g1493_n_spl_1
  );


  buf

  (
    G2441_i2,
    g1501_p_spl_0
  );


  buf

  (
    G2887_i2,
    G2796_o2_p
  );


  buf

  (
    G2991_i2,
    G2906_o2_p
  );


  buf

  (
    G470_i2,
    n5292_o2_p_spl_
  );


  buf

  (
    G484_i2,
    n5293_o2_p_spl_
  );


  buf

  (
    G496_i2,
    n5294_o2_p_spl_1
  );


  buf

  (
    G353_i2,
    n1821_lo_buf_o2_p_spl_1
  );


  buf

  (
    G363_i2,
    n1821_lo_buf_o2_p_spl_1
  );


  buf

  (
    G2805_i2,
    g1045_p_spl_1
  );


  not

  (
    G2906_i2,
    g1504_n_spl_
  );


  not

  (
    G2833_i2,
    g1506_n_spl_
  );


  buf

  (
    G1012_i2,
    g1507_n_spl_
  );


  not

  (
    G3353_i2,
    g1254_p_spl_
  );


  not

  (
    G3367_i2,
    g1256_p_spl_
  );


  not

  (
    G3346_i2,
    g1508_n
  );


  not

  (
    G3340_i2,
    g1509_p
  );


  not

  (
    G3376_i2,
    g1085_p_spl_1
  );


  buf

  (
    G3359_i2,
    g1510_p
  );


  not

  (
    G3240_i2,
    g1258_p_spl_1
  );


  not

  (
    G3344_i2,
    g1511_n
  );


  not

  (
    G2880_i2,
    g1517_n_spl_
  );


  not

  (
    G2939_i2,
    g1518_n_spl_
  );


  not

  (
    G2248_i2,
    g1520_n_spl_
  );


  not

  (
    G2251_i2,
    g1522_n_spl_
  );


  not

  (
    G2021_i2,
    g1523_n_spl_0
  );


  not

  (
    G3383_i2,
    g1303_n_spl_
  );


  not

  (
    G3399_i2,
    g1304_n_spl_
  );


  not

  (
    G3404_i2,
    g1085_p_spl_1
  );


  not

  (
    G3265_i2,
    g1258_p_spl_1
  );


  not

  (
    G2866_i2,
    g1524_n_spl_1
  );


  not

  (
    G2999_i2,
    g1526_n_spl_1
  );


  buf

  (
    G736_i2,
    n5295_o2_p_spl_00
  );


  buf

  (
    G739_i2,
    n5295_o2_p_spl_0
  );


  buf

  (
    G1200_i2,
    g1529_n_spl_
  );


  buf

  (
    G1203_i2,
    g1532_n_spl_
  );


  buf

  (
    G3027_i2,
    g1535_n_spl_
  );


  buf

  (
    G1463_i2,
    g1538_n_spl_
  );


  buf

  (
    G1460_i2,
    g1541_n_spl_
  );


  buf

  (
    G3012_i2,
    g1554_n_spl_
  );


  not

  (
    G1574_i2,
    g1558_n_spl_000
  );


  not

  (
    G1646_i2,
    g1558_n_spl_000
  );


  not

  (
    G1592_i2,
    g1559_n_spl_000
  );


  not

  (
    G1664_i2,
    g1559_n_spl_000
  );


  not

  (
    G1547_i2,
    g1562_p_spl_000
  );


  not

  (
    G1619_i2,
    g1562_p_spl_000
  );


  not

  (
    G1556_i2,
    g1564_n_spl_000
  );


  not

  (
    G1628_i2,
    g1564_n_spl_000
  );


  buf

  (
    G1583_i2,
    g1566_n_spl_000
  );


  buf

  (
    G1655_i2,
    g1566_n_spl_000
  );


  buf

  (
    G1529_i2,
    g1567_p_spl_000
  );


  buf

  (
    G1601_i2,
    g1567_p_spl_000
  );


  not

  (
    G1538_i2,
    g1568_n_spl_000
  );


  not

  (
    G1610_i2,
    g1568_n_spl_000
  );


  not

  (
    G1565_i2,
    g1569_n_spl_000
  );


  not

  (
    G1637_i2,
    g1569_n_spl_000
  );


  buf

  (
    G2437_i2,
    g1577_p_spl_0
  );


  buf

  (
    G2518_i2,
    g1501_p_spl_0
  );


  buf

  (
    n1785_lo_buf_i2,
    G4_p_spl_10
  );


  buf

  (
    n1845_lo_buf_i2,
    G9_p_spl_0
  );


  buf

  (
    n1893_lo_buf_i2,
    G13_p_spl_0
  );


  buf

  (
    n1941_lo_buf_i2,
    n1938_lo_p
  );


  buf

  (
    n1953_lo_buf_i2,
    n1950_lo_p
  );


  buf

  (
    n1965_lo_buf_i2,
    n1962_lo_p
  );


  buf

  (
    n1977_lo_buf_i2,
    n1974_lo_p
  );


  buf

  (
    n2241_lo_buf_i2,
    n2238_lo_p
  );


  buf

  (
    n2253_lo_buf_i2,
    n2250_lo_p
  );


  buf

  (
    n2265_lo_buf_i2,
    n2262_lo_p
  );


  buf

  (
    n2277_lo_buf_i2,
    n2274_lo_p
  );


  buf

  (
    n2289_lo_buf_i2,
    n2286_lo_p
  );


  buf

  (
    G519_i2,
    n5099_o2_p
  );


  buf

  (
    G388_i2,
    n5100_o2_p_spl_1
  );


  buf

  (
    G438_i2,
    n5101_o2_p_spl_
  );


  buf

  (
    G368_i2,
    n5266_o2_p_spl_1
  );


  not

  (
    G1318_i2,
    g1581_n
  );


  buf

  (
    G425_i2,
    n5267_o2_p_spl_1
  );


  buf

  (
    G593_i2,
    n5294_o2_p_spl_1
  );


  buf

  (
    G413_i2,
    n5325_o2_p_spl_1
  );


  buf

  (
    G404_i2,
    n1857_lo_buf_o2_p_spl_1
  );


  buf

  (
    G451_i2,
    n1905_lo_buf_o2_p_spl_1
  );


  buf

  (
    G2284_i2,
    G2018_o2_p
  );


  buf

  (
    G2580_i2,
    n1464_inv_p
  );


  buf

  (
    G2302_i2,
    G2027_o2_p_spl_
  );


  buf

  (
    G2598_i2,
    n1554_inv_p_spl_
  );


  buf

  (
    G2497_i2,
    g1512_p_spl_
  );


  buf

  (
    G2651_i2,
    G2507_o2_p_spl_1
  );


  buf

  (
    G2296_i2,
    g1542_p_spl_
  );


  buf

  (
    G2308_i2,
    g1305_p_spl_
  );


  buf

  (
    G2592_i2,
    G2444_o2_p_spl_1
  );


  buf

  (
    G2604_i2,
    g1049_p_spl_1
  );


  not

  (
    G2902_i2,
    g1584_n
  );


  not

  (
    G2975_i2,
    g1585_n
  );


  not

  (
    G2962_i2,
    g1586_n_spl_
  );


  not

  (
    G3069_i2,
    g1591_n_spl_
  );


  not

  (
    G2018_i2,
    g1592_n_spl_
  );


  not

  (
    G1176_i2,
    g1481_n_spl_
  );


  not

  (
    G1189_i2,
    g1482_n_spl_1
  );


  not

  (
    G3066_i2,
    g1593_p
  );


  not

  (
    G3137_i2,
    g1594_p
  );


  not

  (
    G3038_i2,
    g1595_n
  );


  not

  (
    G3117_i2,
    g1596_n
  );


  buf

  (
    G2384_i2,
    g1612_n_spl_
  );


  buf

  (
    G2472_i2,
    g1617_n_spl_
  );


  buf

  (
    G772_i2,
    g1619_n
  );


  buf

  (
    G935_i2,
    g1621_p
  );


  not

  (
    G2923_i2,
    g1622_p
  );


  not

  (
    G2971_i2,
    g1517_n_spl_
  );


  not

  (
    G2980_i2,
    g1518_n_spl_
  );


  buf

  (
    G3039_i2,
    g1624_p
  );


  not

  (
    G2388_i2,
    g1625_p_spl_
  );


  not

  (
    G2287_i2,
    g1523_n_spl_0
  );


  buf

  (
    G3024_i2,
    g1633_n
  );


  not

  (
    G2916_i2,
    g1524_n_spl_1
  );


  buf

  (
    G1819_i2,
    g1642_p
  );


  not

  (
    G3035_i2,
    g1526_n_spl_1
  );


  buf

  (
    G3107_i2,
    g1648_n
  );


  buf

  (
    G1023_i2,
    n5295_o2_p_spl_1
  );


  buf

  (
    G1024_i2,
    n5295_o2_p_spl_1
  );


  buf

  (
    G1311_i2,
    g1529_n_spl_
  );


  buf

  (
    G1312_i2,
    g1532_n_spl_
  );


  buf

  (
    G3063_i2,
    g1535_n_spl_
  );


  buf

  (
    G1520_i2,
    g1538_n_spl_
  );


  buf

  (
    G1519_i2,
    g1541_n_spl_
  );


  buf

  (
    G3078_i2,
    g1554_n_spl_
  );


  buf

  (
    G2038_i2,
    g1651_n
  );


  not

  (
    G1848_i2,
    g1558_n_spl_001
  );


  not

  (
    G1864_i2,
    g1558_n_spl_001
  );


  not

  (
    G1872_i2,
    g1558_n_spl_010
  );


  not

  (
    G1880_i2,
    g1558_n_spl_010
  );


  not

  (
    G1888_i2,
    g1558_n_spl_011
  );


  not

  (
    G1912_i2,
    g1558_n_spl_011
  );


  not

  (
    G1928_i2,
    g1558_n_spl_10
  );


  not

  (
    G1936_i2,
    g1558_n_spl_10
  );


  not

  (
    G1944_i2,
    g1558_n_spl_11
  );


  not

  (
    G1952_i2,
    g1558_n_spl_11
  );


  not

  (
    G1850_i2,
    g1559_n_spl_001
  );


  not

  (
    G1866_i2,
    g1559_n_spl_001
  );


  not

  (
    G1874_i2,
    g1559_n_spl_010
  );


  not

  (
    G1882_i2,
    g1559_n_spl_010
  );


  not

  (
    G1890_i2,
    g1559_n_spl_011
  );


  not

  (
    G1914_i2,
    g1559_n_spl_011
  );


  not

  (
    G1930_i2,
    g1559_n_spl_10
  );


  not

  (
    G1938_i2,
    g1559_n_spl_10
  );


  not

  (
    G1946_i2,
    g1559_n_spl_11
  );


  not

  (
    G1954_i2,
    g1559_n_spl_11
  );


  not

  (
    G1845_i2,
    g1562_p_spl_001
  );


  not

  (
    G1861_i2,
    g1562_p_spl_001
  );


  not

  (
    G1869_i2,
    g1562_p_spl_010
  );


  not

  (
    G1877_i2,
    g1562_p_spl_010
  );


  not

  (
    G1885_i2,
    g1562_p_spl_011
  );


  not

  (
    G1909_i2,
    g1562_p_spl_011
  );


  not

  (
    G1925_i2,
    g1562_p_spl_10
  );


  not

  (
    G1933_i2,
    g1562_p_spl_10
  );


  not

  (
    G1941_i2,
    g1562_p_spl_11
  );


  not

  (
    G1949_i2,
    g1562_p_spl_11
  );


  not

  (
    G1846_i2,
    g1564_n_spl_001
  );


  not

  (
    G1862_i2,
    g1564_n_spl_001
  );


  not

  (
    G1870_i2,
    g1564_n_spl_010
  );


  not

  (
    G1878_i2,
    g1564_n_spl_010
  );


  not

  (
    G1886_i2,
    g1564_n_spl_011
  );


  not

  (
    G1910_i2,
    g1564_n_spl_011
  );


  not

  (
    G1926_i2,
    g1564_n_spl_10
  );


  not

  (
    G1934_i2,
    g1564_n_spl_10
  );


  not

  (
    G1942_i2,
    g1564_n_spl_11
  );


  not

  (
    G1950_i2,
    g1564_n_spl_11
  );


  buf

  (
    G1849_i2,
    g1566_n_spl_001
  );


  buf

  (
    G1865_i2,
    g1566_n_spl_001
  );


  buf

  (
    G1873_i2,
    g1566_n_spl_010
  );


  buf

  (
    G1881_i2,
    g1566_n_spl_010
  );


  buf

  (
    G1889_i2,
    g1566_n_spl_011
  );


  buf

  (
    G1913_i2,
    g1566_n_spl_011
  );


  buf

  (
    G1929_i2,
    g1566_n_spl_10
  );


  buf

  (
    G1937_i2,
    g1566_n_spl_10
  );


  buf

  (
    G1945_i2,
    g1566_n_spl_11
  );


  buf

  (
    G1953_i2,
    g1566_n_spl_11
  );


  buf

  (
    G1843_i2,
    g1567_p_spl_001
  );


  buf

  (
    G1859_i2,
    g1567_p_spl_001
  );


  buf

  (
    G1867_i2,
    g1567_p_spl_010
  );


  buf

  (
    G1875_i2,
    g1567_p_spl_010
  );


  buf

  (
    G1883_i2,
    g1567_p_spl_011
  );


  buf

  (
    G1907_i2,
    g1567_p_spl_011
  );


  buf

  (
    G1923_i2,
    g1567_p_spl_10
  );


  buf

  (
    G1931_i2,
    g1567_p_spl_10
  );


  buf

  (
    G1939_i2,
    g1567_p_spl_11
  );


  buf

  (
    G1947_i2,
    g1567_p_spl_11
  );


  not

  (
    G1844_i2,
    g1568_n_spl_001
  );


  not

  (
    G1860_i2,
    g1568_n_spl_001
  );


  not

  (
    G1868_i2,
    g1568_n_spl_010
  );


  not

  (
    G1876_i2,
    g1568_n_spl_010
  );


  not

  (
    G1884_i2,
    g1568_n_spl_011
  );


  not

  (
    G1908_i2,
    g1568_n_spl_011
  );


  not

  (
    G1924_i2,
    g1568_n_spl_10
  );


  not

  (
    G1932_i2,
    g1568_n_spl_10
  );


  not

  (
    G1940_i2,
    g1568_n_spl_11
  );


  not

  (
    G1948_i2,
    g1568_n_spl_11
  );


  not

  (
    G1847_i2,
    g1569_n_spl_001
  );


  not

  (
    G1863_i2,
    g1569_n_spl_001
  );


  not

  (
    G1871_i2,
    g1569_n_spl_010
  );


  not

  (
    G1879_i2,
    g1569_n_spl_010
  );


  not

  (
    G1887_i2,
    g1569_n_spl_011
  );


  not

  (
    G1911_i2,
    g1569_n_spl_011
  );


  not

  (
    G1927_i2,
    g1569_n_spl_10
  );


  not

  (
    G1935_i2,
    g1569_n_spl_10
  );


  not

  (
    G1943_i2,
    g1569_n_spl_11
  );


  not

  (
    G1951_i2,
    g1569_n_spl_11
  );


  not

  (
    G2444_i2,
    g1663_n_spl_1
  );


  not

  (
    G2451_i2,
    g1670_n_spl_0
  );


  buf

  (
    G2502_i2,
    g1678_p_spl_
  );


  not

  (
    G2507_i2,
    g1685_n_spl_
  );


  buf

  (
    G2515_i2,
    g1577_p_spl_0
  );


  buf

  (
    G2583_i2,
    g1501_p_spl_1
  );


  buf

  (
    n1797_lo_buf_i2,
    G5_p_spl_
  );


  buf

  (
    n1833_lo_buf_i2,
    G8_p_spl_0
  );


  buf

  (
    n1881_lo_buf_i2,
    G12_p_spl_0
  );


  buf

  (
    G523_i2,
    G4_p_spl_10
  );


  buf

  (
    G575_i2,
    G9_p_spl_0
  );


  buf

  (
    G578_i2,
    G13_p_spl_0
  );


  buf

  (
    G615_i2,
    n2019_lo_p_spl_1
  );


  not

  (
    G2254_i2,
    g1687_n
  );


  not

  (
    G2255_i2,
    g1689_n
  );


  not

  (
    G2027_i2,
    g1690_n
  );


  not

  (
    G2393_i2,
    g1691_n
  );


  buf

  (
    G527_i2,
    g1692_p_spl_
  );


  buf

  (
    G594_i2,
    g1693_n_spl_0
  );


  buf

  (
    G1689_i2,
    g1706_n_spl_
  );


  buf

  (
    G1693_i2,
    g1706_n_spl_
  );


  not

  (
    G2281_i2,
    g1592_n_spl_
  );


  buf

  (
    G2014_i2,
    g1493_n_spl_1
  );


  buf

  (
    G2459_i2,
    g1656_n_spl_
  );


  not

  (
    G2561_i2,
    g1708_n
  );


  not

  (
    G2533_i2,
    g1709_n
  );


  buf

  (
    n1749_lo_buf_i2,
    G1_p_spl_
  );


  buf

  (
    n1761_lo_buf_i2,
    G2_p_spl_
  );


  buf

  (
    n1773_lo_buf_i2,
    G3_p_spl_0
  );


  buf

  (
    n1809_lo_buf_i2,
    G6_p_spl_
  );


  buf

  (
    G1955_i2,
    g1719_n_spl_
  );


  buf

  (
    G1958_i2,
    g1719_n_spl_
  );


  not

  (
    G2562_i2,
    g1722_n
  );


  not

  (
    G2398_i2,
    g1523_n_spl_
  );


  not

  (
    G2524_i2,
    g1670_n_spl_
  );


  buf

  (
    G2563_i2,
    g1678_p_spl_
  );


  buf

  (
    G2577_i2,
    g1577_p_spl_
  );


  buf

  (
    G2627_i2,
    g1501_p_spl_1
  );


  buf

  (
    G654_i2,
    G8_p_spl_0
  );


  buf

  (
    G660_i2,
    G12_p_spl_0
  );


  buf

  (
    G831_i2,
    G4_p_spl_11
  );


  buf

  (
    G919_i2,
    G9_p_spl_1
  );


  buf

  (
    G925_i2,
    G13_p_spl_1
  );


  buf

  (
    n1815_lo_buf_i2,
    G7_p
  );


  buf

  (
    n1899_lo_buf_i2,
    G14_p
  );


  buf

  (
    n2079_lo_buf_i2,
    G29_p
  );


  buf

  (
    n2127_lo_buf_i2,
    G33_p
  );


  buf

  (
    n2139_lo_buf_i2,
    G34_p
  );


  buf

  (
    n2151_lo_buf_i2,
    G35_p
  );


  buf

  (
    n2187_lo_buf_i2,
    G38_p
  );


  buf

  (
    n2199_lo_buf_i2,
    G39_p
  );


  buf

  (
    n2211_lo_buf_i2,
    G40_p
  );


  buf

  (
    G533_i2,
    g1723_n
  );


  buf

  (
    n1854_lo_buf_i2,
    G10_p
  );


  buf

  (
    n2094_lo_buf_i2,
    G30_p
  );


  buf

  (
    G667_i2,
    g1724_p
  );


  buf

  (
    G874_i2,
    g1692_p_spl_
  );


  buf

  (
    G851_i2,
    g1693_n_spl_
  );


  buf

  (
    G1127_i2,
    g1725_p
  );


  buf

  (
    n1869_lo_buf_i2,
    G11_p
  );


  buf

  (
    n2109_lo_buf_i2,
    G31_p
  );


  buf

  (
    n2121_lo_buf_i2,
    G32_p
  );


  buf

  (
    G477_i2,
    G1_p_spl_
  );


  buf

  (
    G491_i2,
    g1726_p
  );


  buf

  (
    G501_i2,
    G3_p_spl_
  );


  buf

  (
    G786_i2,
    G8_p_spl_
  );


  buf

  (
    G791_i2,
    G12_p_spl_
  );


  buf

  (
    G1126_i2,
    G4_p_spl_11
  );


  buf

  (
    G1052_i2,
    G9_p_spl_1
  );


  buf

  (
    G1054_i2,
    G13_p_spl_1
  );


  buf

  (
    n5011_o2_n_spl_,
    n5011_o2_n
  );


  buf

  (
    n5011_o2_p_spl_,
    n5011_o2_p
  );


  buf

  (
    n5013_o2_n_spl_,
    n5013_o2_n
  );


  buf

  (
    n5013_o2_p_spl_,
    n5013_o2_p
  );


  buf

  (
    g585_n_spl_,
    g585_n
  );


  buf

  (
    n2172_lo_n_spl_,
    n2172_lo_n
  );


  buf

  (
    n2160_lo_n_spl_,
    n2160_lo_n
  );


  buf

  (
    n2148_lo_n_spl_,
    n2148_lo_n
  );


  buf

  (
    g589_p_spl_,
    g589_p
  );


  buf

  (
    g589_n_spl_,
    g589_n
  );


  buf

  (
    g585_p_spl_,
    g585_p
  );


  buf

  (
    n4634_o2_n_spl_,
    n4634_o2_n
  );


  buf

  (
    n4633_o2_p_spl_,
    n4633_o2_p
  );


  buf

  (
    n4634_o2_p_spl_,
    n4634_o2_p
  );


  buf

  (
    n4633_o2_n_spl_,
    n4633_o2_n
  );


  buf

  (
    n4418_o2_p_spl_,
    n4418_o2_p
  );


  buf

  (
    n2304_lo_p_spl_,
    n2304_lo_p
  );


  buf

  (
    g633_n_spl_,
    g633_n
  );


  buf

  (
    g636_n_spl_,
    g636_n
  );


  buf

  (
    G2991_o2_n_spl_,
    G2991_o2_n
  );


  buf

  (
    G2887_o2_p_spl_,
    G2887_o2_p
  );


  buf

  (
    G2991_o2_p_spl_,
    G2991_o2_p
  );


  buf

  (
    G2887_o2_n_spl_,
    G2887_o2_n
  );


  buf

  (
    n4733_o2_p_spl_,
    n4733_o2_p
  );


  buf

  (
    n4732_o2_p_spl_,
    n4732_o2_p
  );


  buf

  (
    n4733_o2_n_spl_,
    n4733_o2_n
  );


  buf

  (
    n4732_o2_n_spl_,
    n4732_o2_n
  );


  buf

  (
    g666_n_spl_,
    g666_n
  );


  buf

  (
    g669_n_spl_,
    g669_n
  );


  buf

  (
    g672_n_spl_,
    g672_n
  );


  buf

  (
    g675_n_spl_,
    g675_n
  );


  buf

  (
    g681_n_spl_,
    g681_n
  );


  buf

  (
    g683_n_spl_,
    g683_n
  );


  buf

  (
    g688_n_spl_,
    g688_n
  );


  buf

  (
    g687_n_spl_,
    g687_n
  );


  buf

  (
    g694_n_spl_,
    g694_n
  );


  buf

  (
    g693_p_spl_,
    g693_p
  );


  buf

  (
    g694_p_spl_,
    g694_p
  );


  buf

  (
    g693_n_spl_,
    g693_n
  );


  buf

  (
    G3360_o2_p_spl_,
    G3360_o2_p
  );


  buf

  (
    G3350_o2_n_spl_,
    G3350_o2_n
  );


  buf

  (
    G3360_o2_n_spl_,
    G3360_o2_n
  );


  buf

  (
    G3350_o2_p_spl_,
    G3350_o2_p
  );


  buf

  (
    g703_n_spl_,
    g703_n
  );


  buf

  (
    g700_n_spl_,
    g700_n
  );


  buf

  (
    g700_n_spl_0,
    g700_n_spl_
  );


  buf

  (
    g700_n_spl_1,
    g700_n_spl_
  );


  buf

  (
    g703_p_spl_,
    g703_p
  );


  buf

  (
    g700_p_spl_,
    g700_p
  );


  buf

  (
    g700_p_spl_0,
    g700_p_spl_
  );


  buf

  (
    g700_p_spl_1,
    g700_p_spl_
  );


  buf

  (
    g704_p_spl_,
    g704_p
  );


  buf

  (
    g704_p_spl_0,
    g704_p_spl_
  );


  buf

  (
    g704_p_spl_1,
    g704_p_spl_
  );


  buf

  (
    g704_n_spl_,
    g704_n
  );


  buf

  (
    g704_n_spl_0,
    g704_n_spl_
  );


  buf

  (
    g704_n_spl_1,
    g704_n_spl_
  );


  buf

  (
    G3399_o2_p_spl_,
    G3399_o2_p
  );


  buf

  (
    G3383_o2_n_spl_,
    G3383_o2_n
  );


  buf

  (
    G3399_o2_n_spl_,
    G3399_o2_n
  );


  buf

  (
    G3383_o2_p_spl_,
    G3383_o2_p
  );


  buf

  (
    g709_p_spl_,
    g709_p
  );


  buf

  (
    g709_n_spl_,
    g709_n
  );


  buf

  (
    G3240_o2_p_spl_,
    G3240_o2_p
  );


  buf

  (
    G3376_o2_p_spl_,
    G3376_o2_p
  );


  buf

  (
    G3240_o2_n_spl_,
    G3240_o2_n
  );


  buf

  (
    G3376_o2_n_spl_,
    G3376_o2_n
  );


  buf

  (
    g714_p_spl_,
    g714_p
  );


  buf

  (
    g714_n_spl_,
    g714_n
  );


  buf

  (
    g697_n_spl_,
    g697_n
  );


  buf

  (
    g697_p_spl_,
    g697_p
  );


  buf

  (
    G3367_o2_n_spl_,
    G3367_o2_n
  );


  buf

  (
    G3353_o2_p_spl_,
    G3353_o2_p
  );


  buf

  (
    G3367_o2_p_spl_,
    G3367_o2_p
  );


  buf

  (
    G3353_o2_n_spl_,
    G3353_o2_n
  );


  buf

  (
    g727_n_spl_,
    g727_n
  );


  buf

  (
    g727_p_spl_,
    g727_p
  );


  buf

  (
    G434_o2_p_spl_,
    G434_o2_p
  );


  buf

  (
    n852_inv_n_spl_,
    n852_inv_n
  );


  buf

  (
    n852_inv_n_spl_0,
    n852_inv_n_spl_
  );


  buf

  (
    n849_inv_n_spl_,
    n849_inv_n
  );


  buf

  (
    n852_inv_p_spl_,
    n852_inv_p
  );


  buf

  (
    n852_inv_p_spl_0,
    n852_inv_p_spl_
  );


  buf

  (
    n852_inv_p_spl_1,
    n852_inv_p_spl_
  );


  buf

  (
    n849_inv_p_spl_,
    n849_inv_p
  );


  buf

  (
    n849_inv_p_spl_0,
    n849_inv_p_spl_
  );


  buf

  (
    n855_inv_p_spl_,
    n855_inv_p
  );


  buf

  (
    n4539_o2_p_spl_,
    n4539_o2_p
  );


  buf

  (
    n4539_o2_p_spl_0,
    n4539_o2_p_spl_
  );


  buf

  (
    n4539_o2_n_spl_,
    n4539_o2_n
  );


  buf

  (
    n4539_o2_n_spl_0,
    n4539_o2_n_spl_
  );


  buf

  (
    n4816_o2_n_spl_,
    n4816_o2_n
  );


  buf

  (
    n429_inv_n_spl_,
    n429_inv_n
  );


  buf

  (
    n4816_o2_p_spl_,
    n4816_o2_p
  );


  buf

  (
    n429_inv_p_spl_,
    n429_inv_p
  );


  buf

  (
    n429_inv_p_spl_0,
    n429_inv_p_spl_
  );


  buf

  (
    n4398_o2_p_spl_,
    n4398_o2_p
  );


  buf

  (
    g752_n_spl_,
    g752_n
  );


  buf

  (
    g752_n_spl_0,
    g752_n_spl_
  );


  buf

  (
    g749_n_spl_,
    g749_n
  );


  buf

  (
    g756_p_spl_,
    g756_p
  );


  buf

  (
    g756_p_spl_0,
    g756_p_spl_
  );


  buf

  (
    g752_p_spl_,
    g752_p
  );


  buf

  (
    g752_p_spl_0,
    g752_p_spl_
  );


  buf

  (
    g752_p_spl_00,
    g752_p_spl_0
  );


  buf

  (
    g752_p_spl_01,
    g752_p_spl_0
  );


  buf

  (
    g752_p_spl_1,
    g752_p_spl_
  );


  buf

  (
    g752_p_spl_10,
    g752_p_spl_1
  );


  buf

  (
    G3069_o2_n_spl_,
    G3069_o2_n
  );


  buf

  (
    G2962_o2_n_spl_,
    G2962_o2_n
  );


  buf

  (
    G3069_o2_p_spl_,
    G3069_o2_p
  );


  buf

  (
    G2962_o2_p_spl_,
    G2962_o2_p
  );


  buf

  (
    g760_p_spl_,
    g760_p
  );


  buf

  (
    g760_p_spl_0,
    g760_p_spl_
  );


  buf

  (
    g764_p_spl_,
    g764_p
  );


  buf

  (
    n1941_lo_buf_o2_n_spl_,
    n1941_lo_buf_o2_n
  );


  buf

  (
    n1941_lo_buf_o2_n_spl_0,
    n1941_lo_buf_o2_n_spl_
  );


  buf

  (
    n1056_inv_p_spl_,
    n1056_inv_p
  );


  buf

  (
    n1056_inv_p_spl_0,
    n1056_inv_p_spl_
  );


  buf

  (
    n1056_inv_p_spl_00,
    n1056_inv_p_spl_0
  );


  buf

  (
    n1056_inv_p_spl_01,
    n1056_inv_p_spl_0
  );


  buf

  (
    n1056_inv_p_spl_1,
    n1056_inv_p_spl_
  );


  buf

  (
    n858_inv_p_spl_,
    n858_inv_p
  );


  buf

  (
    n858_inv_p_spl_0,
    n858_inv_p_spl_
  );


  buf

  (
    n858_inv_p_spl_00,
    n858_inv_p_spl_0
  );


  buf

  (
    n858_inv_p_spl_01,
    n858_inv_p_spl_0
  );


  buf

  (
    n858_inv_p_spl_1,
    n858_inv_p_spl_
  );


  buf

  (
    n4651_o2_n_spl_,
    n4651_o2_n
  );


  buf

  (
    n4651_o2_n_spl_0,
    n4651_o2_n_spl_
  );


  buf

  (
    n4651_o2_n_spl_00,
    n4651_o2_n_spl_0
  );


  buf

  (
    n4651_o2_n_spl_01,
    n4651_o2_n_spl_0
  );


  buf

  (
    n4651_o2_n_spl_1,
    n4651_o2_n_spl_
  );


  buf

  (
    n4919_o2_n_spl_,
    n4919_o2_n
  );


  buf

  (
    n4919_o2_n_spl_0,
    n4919_o2_n_spl_
  );


  buf

  (
    n4919_o2_n_spl_00,
    n4919_o2_n_spl_0
  );


  buf

  (
    n4919_o2_n_spl_01,
    n4919_o2_n_spl_0
  );


  buf

  (
    n4919_o2_n_spl_1,
    n4919_o2_n_spl_
  );


  buf

  (
    n1977_lo_buf_o2_n_spl_,
    n1977_lo_buf_o2_n
  );


  buf

  (
    n1977_lo_buf_o2_n_spl_0,
    n1977_lo_buf_o2_n_spl_
  );


  buf

  (
    n1977_lo_buf_o2_n_spl_00,
    n1977_lo_buf_o2_n_spl_0
  );


  buf

  (
    n1977_lo_buf_o2_n_spl_1,
    n1977_lo_buf_o2_n_spl_
  );


  buf

  (
    n1965_lo_buf_o2_n_spl_,
    n1965_lo_buf_o2_n
  );


  buf

  (
    n1965_lo_buf_o2_n_spl_0,
    n1965_lo_buf_o2_n_spl_
  );


  buf

  (
    n1965_lo_buf_o2_n_spl_00,
    n1965_lo_buf_o2_n_spl_0
  );


  buf

  (
    n1965_lo_buf_o2_n_spl_1,
    n1965_lo_buf_o2_n_spl_
  );


  buf

  (
    n1953_lo_buf_o2_n_spl_,
    n1953_lo_buf_o2_n
  );


  buf

  (
    n1953_lo_buf_o2_n_spl_0,
    n1953_lo_buf_o2_n_spl_
  );


  buf

  (
    n1953_lo_buf_o2_n_spl_1,
    n1953_lo_buf_o2_n_spl_
  );


  buf

  (
    G519_o2_n_spl_,
    G519_o2_n
  );


  buf

  (
    G519_o2_n_spl_0,
    G519_o2_n_spl_
  );


  buf

  (
    G519_o2_n_spl_00,
    G519_o2_n_spl_0
  );


  buf

  (
    G519_o2_n_spl_000,
    G519_o2_n_spl_00
  );


  buf

  (
    G519_o2_n_spl_01,
    G519_o2_n_spl_0
  );


  buf

  (
    G519_o2_n_spl_1,
    G519_o2_n_spl_
  );


  buf

  (
    G519_o2_n_spl_10,
    G519_o2_n_spl_1
  );


  buf

  (
    G519_o2_n_spl_11,
    G519_o2_n_spl_1
  );


  buf

  (
    n4653_o2_n_spl_,
    n4653_o2_n
  );


  buf

  (
    n4653_o2_n_spl_0,
    n4653_o2_n_spl_
  );


  buf

  (
    n4653_o2_n_spl_1,
    n4653_o2_n_spl_
  );


  buf

  (
    n1071_inv_p_spl_,
    n1071_inv_p
  );


  buf

  (
    n1071_inv_p_spl_0,
    n1071_inv_p_spl_
  );


  buf

  (
    n1071_inv_p_spl_00,
    n1071_inv_p_spl_0
  );


  buf

  (
    n1071_inv_p_spl_01,
    n1071_inv_p_spl_0
  );


  buf

  (
    n1071_inv_p_spl_1,
    n1071_inv_p_spl_
  );


  buf

  (
    n1068_inv_p_spl_,
    n1068_inv_p
  );


  buf

  (
    n1068_inv_p_spl_0,
    n1068_inv_p_spl_
  );


  buf

  (
    n1068_inv_p_spl_00,
    n1068_inv_p_spl_0
  );


  buf

  (
    n1068_inv_p_spl_01,
    n1068_inv_p_spl_0
  );


  buf

  (
    n1068_inv_p_spl_1,
    n1068_inv_p_spl_
  );


  buf

  (
    n1062_inv_p_spl_,
    n1062_inv_p
  );


  buf

  (
    n1062_inv_p_spl_0,
    n1062_inv_p_spl_
  );


  buf

  (
    n1062_inv_p_spl_00,
    n1062_inv_p_spl_0
  );


  buf

  (
    n1062_inv_p_spl_01,
    n1062_inv_p_spl_0
  );


  buf

  (
    n1062_inv_p_spl_1,
    n1062_inv_p_spl_
  );


  buf

  (
    n1062_inv_p_spl_10,
    n1062_inv_p_spl_1
  );


  buf

  (
    n1053_inv_p_spl_,
    n1053_inv_p
  );


  buf

  (
    n1053_inv_p_spl_0,
    n1053_inv_p_spl_
  );


  buf

  (
    n1053_inv_p_spl_00,
    n1053_inv_p_spl_0
  );


  buf

  (
    n1053_inv_p_spl_01,
    n1053_inv_p_spl_0
  );


  buf

  (
    n1053_inv_p_spl_1,
    n1053_inv_p_spl_
  );


  buf

  (
    n1074_inv_p_spl_,
    n1074_inv_p
  );


  buf

  (
    n1074_inv_p_spl_0,
    n1074_inv_p_spl_
  );


  buf

  (
    n1074_inv_p_spl_00,
    n1074_inv_p_spl_0
  );


  buf

  (
    n1074_inv_p_spl_01,
    n1074_inv_p_spl_0
  );


  buf

  (
    n1074_inv_p_spl_1,
    n1074_inv_p_spl_
  );


  buf

  (
    n1074_inv_p_spl_10,
    n1074_inv_p_spl_1
  );


  buf

  (
    n4571_o2_n_spl_,
    n4571_o2_n
  );


  buf

  (
    n4571_o2_n_spl_0,
    n4571_o2_n_spl_
  );


  buf

  (
    n4571_o2_n_spl_00,
    n4571_o2_n_spl_0
  );


  buf

  (
    n4571_o2_n_spl_01,
    n4571_o2_n_spl_0
  );


  buf

  (
    n4571_o2_n_spl_1,
    n4571_o2_n_spl_
  );


  buf

  (
    n4572_o2_n_spl_,
    n4572_o2_n
  );


  buf

  (
    n4572_o2_n_spl_0,
    n4572_o2_n_spl_
  );


  buf

  (
    n4572_o2_n_spl_00,
    n4572_o2_n_spl_0
  );


  buf

  (
    n4572_o2_n_spl_1,
    n4572_o2_n_spl_
  );


  buf

  (
    G519_o2_p_spl_,
    G519_o2_p
  );


  buf

  (
    G519_o2_p_spl_0,
    G519_o2_p_spl_
  );


  buf

  (
    G519_o2_p_spl_00,
    G519_o2_p_spl_0
  );


  buf

  (
    G519_o2_p_spl_000,
    G519_o2_p_spl_00
  );


  buf

  (
    G519_o2_p_spl_01,
    G519_o2_p_spl_0
  );


  buf

  (
    G519_o2_p_spl_1,
    G519_o2_p_spl_
  );


  buf

  (
    G519_o2_p_spl_10,
    G519_o2_p_spl_1
  );


  buf

  (
    G519_o2_p_spl_11,
    G519_o2_p_spl_1
  );


  buf

  (
    g801_n_spl_,
    g801_n
  );


  buf

  (
    g801_n_spl_0,
    g801_n_spl_
  );


  buf

  (
    g801_n_spl_00,
    g801_n_spl_0
  );


  buf

  (
    g801_n_spl_01,
    g801_n_spl_0
  );


  buf

  (
    g801_n_spl_1,
    g801_n_spl_
  );


  buf

  (
    g801_n_spl_10,
    g801_n_spl_1
  );


  buf

  (
    n4389_o2_p_spl_,
    n4389_o2_p
  );


  buf

  (
    n4389_o2_p_spl_0,
    n4389_o2_p_spl_
  );


  buf

  (
    n4389_o2_p_spl_1,
    n4389_o2_p_spl_
  );


  buf

  (
    n4389_o2_n_spl_,
    n4389_o2_n
  );


  buf

  (
    n4389_o2_n_spl_0,
    n4389_o2_n_spl_
  );


  buf

  (
    n4389_o2_n_spl_1,
    n4389_o2_n_spl_
  );


  buf

  (
    g806_p_spl_,
    g806_p
  );


  buf

  (
    g806_p_spl_0,
    g806_p_spl_
  );


  buf

  (
    g806_p_spl_1,
    g806_p_spl_
  );


  buf

  (
    g801_p_spl_,
    g801_p
  );


  buf

  (
    g801_p_spl_0,
    g801_p_spl_
  );


  buf

  (
    g801_p_spl_1,
    g801_p_spl_
  );


  buf

  (
    g808_p_spl_,
    g808_p
  );


  buf

  (
    g808_p_spl_0,
    g808_p_spl_
  );


  buf

  (
    g808_p_spl_1,
    g808_p_spl_
  );


  buf

  (
    g743_p_spl_,
    g743_p
  );


  buf

  (
    g743_p_spl_0,
    g743_p_spl_
  );


  buf

  (
    g743_p_spl_00,
    g743_p_spl_0
  );


  buf

  (
    g743_p_spl_01,
    g743_p_spl_0
  );


  buf

  (
    g743_p_spl_1,
    g743_p_spl_
  );


  buf

  (
    g743_p_spl_10,
    g743_p_spl_1
  );


  buf

  (
    g743_p_spl_11,
    g743_p_spl_1
  );


  buf

  (
    g743_n_spl_,
    g743_n
  );


  buf

  (
    g743_n_spl_0,
    g743_n_spl_
  );


  buf

  (
    g812_n_spl_,
    g812_n
  );


  buf

  (
    g812_n_spl_0,
    g812_n_spl_
  );


  buf

  (
    g812_n_spl_00,
    g812_n_spl_0
  );


  buf

  (
    g812_n_spl_01,
    g812_n_spl_0
  );


  buf

  (
    g812_n_spl_1,
    g812_n_spl_
  );


  buf

  (
    G2923_o2_p_spl_,
    G2923_o2_p
  );


  buf

  (
    G2923_o2_p_spl_0,
    G2923_o2_p_spl_
  );


  buf

  (
    g749_p_spl_,
    g749_p
  );


  buf

  (
    G2923_o2_n_spl_,
    G2923_o2_n
  );


  buf

  (
    G2923_o2_n_spl_0,
    G2923_o2_n_spl_
  );


  buf

  (
    n2301_lo_buf_o2_p_spl_,
    n2301_lo_buf_o2_p
  );


  buf

  (
    n2301_lo_buf_o2_p_spl_0,
    n2301_lo_buf_o2_p_spl_
  );


  buf

  (
    n2301_lo_buf_o2_n_spl_,
    n2301_lo_buf_o2_n
  );


  buf

  (
    g825_n_spl_,
    g825_n
  );


  buf

  (
    n1050_inv_p_spl_,
    n1050_inv_p
  );


  buf

  (
    n1050_inv_p_spl_0,
    n1050_inv_p_spl_
  );


  buf

  (
    n1050_inv_p_spl_00,
    n1050_inv_p_spl_0
  );


  buf

  (
    n1050_inv_p_spl_01,
    n1050_inv_p_spl_0
  );


  buf

  (
    n1050_inv_p_spl_1,
    n1050_inv_p_spl_
  );


  buf

  (
    n2253_lo_buf_o2_n_spl_,
    n2253_lo_buf_o2_n
  );


  buf

  (
    n2241_lo_buf_o2_n_spl_,
    n2241_lo_buf_o2_n
  );


  buf

  (
    n2241_lo_buf_o2_n_spl_0,
    n2241_lo_buf_o2_n_spl_
  );


  buf

  (
    g871_p_spl_,
    g871_p
  );


  buf

  (
    g871_p_spl_0,
    g871_p_spl_
  );


  buf

  (
    G772_o2_n_spl_,
    G772_o2_n
  );


  buf

  (
    G772_o2_p_spl_,
    G772_o2_p
  );


  buf

  (
    g873_p_spl_,
    g873_p
  );


  buf

  (
    g873_p_spl_0,
    g873_p_spl_
  );


  buf

  (
    g737_n_spl_,
    g737_n
  );


  buf

  (
    g875_n_spl_,
    g875_n
  );


  buf

  (
    g875_n_spl_0,
    g875_n_spl_
  );


  buf

  (
    g873_n_spl_,
    g873_n
  );


  buf

  (
    g873_n_spl_0,
    g873_n_spl_
  );


  buf

  (
    g875_p_spl_,
    g875_p
  );


  buf

  (
    g875_p_spl_0,
    g875_p_spl_
  );


  buf

  (
    g876_p_spl_,
    g876_p
  );


  buf

  (
    g871_n_spl_,
    g871_n
  );


  buf

  (
    g871_n_spl_0,
    g871_n_spl_
  );


  buf

  (
    g880_p_spl_,
    g880_p
  );


  buf

  (
    n1068_inv_n_spl_,
    n1068_inv_n
  );


  buf

  (
    n1071_inv_n_spl_,
    n1071_inv_n
  );


  buf

  (
    n1050_inv_n_spl_,
    n1050_inv_n
  );


  buf

  (
    n1056_inv_n_spl_,
    n1056_inv_n
  );


  buf

  (
    n858_inv_n_spl_,
    n858_inv_n
  );


  buf

  (
    n4651_o2_p_spl_,
    n4651_o2_p
  );


  buf

  (
    n2265_lo_buf_o2_p_spl_,
    n2265_lo_buf_o2_p
  );


  buf

  (
    n1053_inv_n_spl_,
    n1053_inv_n
  );


  buf

  (
    n4571_o2_p_spl_,
    n4571_o2_p
  );


  buf

  (
    n4572_o2_p_spl_,
    n4572_o2_p
  );


  buf

  (
    n4653_o2_p_spl_,
    n4653_o2_p
  );


  buf

  (
    n2241_lo_buf_o2_p_spl_,
    n2241_lo_buf_o2_p
  );


  buf

  (
    n2253_lo_buf_o2_p_spl_,
    n2253_lo_buf_o2_p
  );


  buf

  (
    g740_p_spl_,
    g740_p
  );


  buf

  (
    g876_n_spl_,
    g876_n
  );


  buf

  (
    g880_n_spl_,
    g880_n
  );


  buf

  (
    g812_p_spl_,
    g812_p
  );


  buf

  (
    G461_o2_p_spl_,
    G461_o2_p
  );


  buf

  (
    G935_o2_p_spl_,
    G935_o2_p
  );


  buf

  (
    g734_n_spl_,
    g734_n
  );


  buf

  (
    n4454_o2_p_spl_,
    n4454_o2_p
  );


  buf

  (
    G3039_o2_n_spl_,
    G3039_o2_n
  );


  buf

  (
    G3039_o2_n_spl_0,
    G3039_o2_n_spl_
  );


  buf

  (
    G3039_o2_p_spl_,
    G3039_o2_p
  );


  buf

  (
    G3039_o2_p_spl_0,
    G3039_o2_p_spl_
  );


  buf

  (
    n2061_lo_buf_o2_p_spl_,
    n2061_lo_buf_o2_p
  );


  buf

  (
    g1043_p_spl_,
    g1043_p
  );


  buf

  (
    n2313_lo_buf_o2_p_spl_,
    n2313_lo_buf_o2_p
  );


  buf

  (
    g1043_n_spl_,
    g1043_n
  );


  buf

  (
    g1044_n_spl_,
    g1044_n
  );


  buf

  (
    g1044_n_spl_0,
    g1044_n_spl_
  );


  buf

  (
    g1044_n_spl_00,
    g1044_n_spl_0
  );


  buf

  (
    g1044_n_spl_01,
    g1044_n_spl_0
  );


  buf

  (
    g1044_n_spl_1,
    g1044_n_spl_
  );


  buf

  (
    g1044_n_spl_10,
    g1044_n_spl_1
  );


  buf

  (
    g1044_n_spl_11,
    g1044_n_spl_1
  );


  buf

  (
    g746_n_spl_,
    g746_n
  );


  buf

  (
    g1044_p_spl_,
    g1044_p
  );


  buf

  (
    g1044_p_spl_0,
    g1044_p_spl_
  );


  buf

  (
    g1044_p_spl_00,
    g1044_p_spl_0
  );


  buf

  (
    g1044_p_spl_01,
    g1044_p_spl_0
  );


  buf

  (
    g1044_p_spl_1,
    g1044_p_spl_
  );


  buf

  (
    g1044_p_spl_10,
    g1044_p_spl_1
  );


  buf

  (
    g1044_p_spl_11,
    g1044_p_spl_1
  );


  buf

  (
    G2507_o2_p_spl_,
    G2507_o2_p
  );


  buf

  (
    G2507_o2_p_spl_0,
    G2507_o2_p_spl_
  );


  buf

  (
    G2507_o2_p_spl_1,
    G2507_o2_p_spl_
  );


  buf

  (
    G2444_o2_p_spl_,
    G2444_o2_p
  );


  buf

  (
    G2444_o2_p_spl_0,
    G2444_o2_p_spl_
  );


  buf

  (
    G2444_o2_p_spl_1,
    G2444_o2_p_spl_
  );


  buf

  (
    G2507_o2_n_spl_,
    G2507_o2_n
  );


  buf

  (
    G2507_o2_n_spl_0,
    G2507_o2_n_spl_
  );


  buf

  (
    G2444_o2_n_spl_,
    G2444_o2_n
  );


  buf

  (
    G2444_o2_n_spl_0,
    G2444_o2_n_spl_
  );


  buf

  (
    g1049_p_spl_,
    g1049_p
  );


  buf

  (
    g1049_p_spl_0,
    g1049_p_spl_
  );


  buf

  (
    g1049_p_spl_1,
    g1049_p_spl_
  );


  buf

  (
    g1049_n_spl_,
    g1049_n
  );


  buf

  (
    g1049_n_spl_0,
    g1049_n_spl_
  );


  buf

  (
    G3024_o2_n_spl_,
    G3024_o2_n
  );


  buf

  (
    G2902_o2_p_spl_,
    G2902_o2_p
  );


  buf

  (
    G3024_o2_p_spl_,
    G3024_o2_p
  );


  buf

  (
    G2902_o2_n_spl_,
    G2902_o2_n
  );


  buf

  (
    g1058_p_spl_,
    g1058_p
  );


  buf

  (
    g1058_p_spl_0,
    g1058_p_spl_
  );


  buf

  (
    G1689_o2_p_spl_,
    G1689_o2_p
  );


  buf

  (
    G1689_o2_p_spl_0,
    G1689_o2_p_spl_
  );


  buf

  (
    n2013_lo_buf_o2_p_spl_,
    n2013_lo_buf_o2_p
  );


  buf

  (
    G1689_o2_n_spl_,
    G1689_o2_n
  );


  buf

  (
    G1689_o2_n_spl_0,
    G1689_o2_n_spl_
  );


  buf

  (
    G1955_o2_n_spl_,
    G1955_o2_n
  );


  buf

  (
    G1955_o2_p_spl_,
    G1955_o2_p
  );


  buf

  (
    n2025_lo_buf_o2_p_spl_,
    n2025_lo_buf_o2_p
  );


  buf

  (
    n2025_lo_buf_o2_n_spl_,
    n2025_lo_buf_o2_n
  );


  buf

  (
    G1958_o2_n_spl_,
    G1958_o2_n
  );


  buf

  (
    G1958_o2_p_spl_,
    G1958_o2_p
  );


  buf

  (
    G1693_o2_n_spl_,
    G1693_o2_n
  );


  buf

  (
    G1693_o2_n_spl_0,
    G1693_o2_n_spl_
  );


  buf

  (
    n2037_lo_buf_o2_p_spl_,
    n2037_lo_buf_o2_p
  );


  buf

  (
    G1693_o2_p_spl_,
    G1693_o2_p
  );


  buf

  (
    G1693_o2_p_spl_0,
    G1693_o2_p_spl_
  );


  buf

  (
    n2037_lo_buf_o2_n_spl_,
    n2037_lo_buf_o2_n
  );


  buf

  (
    n2049_lo_buf_o2_p_spl_,
    n2049_lo_buf_o2_p
  );


  buf

  (
    n2049_lo_buf_o2_n_spl_,
    n2049_lo_buf_o2_n
  );


  buf

  (
    n2049_lo_buf_o2_n_spl_0,
    n2049_lo_buf_o2_n_spl_
  );


  buf

  (
    g1064_n_spl_,
    g1064_n
  );


  buf

  (
    g1071_p_spl_,
    g1071_p
  );


  buf

  (
    g1071_p_spl_0,
    g1071_p_spl_
  );


  buf

  (
    g1071_p_spl_00,
    g1071_p_spl_0
  );


  buf

  (
    g1071_p_spl_01,
    g1071_p_spl_0
  );


  buf

  (
    g1071_p_spl_1,
    g1071_p_spl_
  );


  buf

  (
    G2502_o2_p_spl_,
    G2502_o2_p
  );


  buf

  (
    g1071_n_spl_,
    g1071_n
  );


  buf

  (
    g1071_n_spl_0,
    g1071_n_spl_
  );


  buf

  (
    g1077_p_spl_,
    g1077_p
  );


  buf

  (
    g1077_p_spl_0,
    g1077_p_spl_
  );


  buf

  (
    g832_p_spl_,
    g832_p
  );


  buf

  (
    g753_p_spl_,
    g753_p
  );


  buf

  (
    g930_p_spl_,
    g930_p
  );


  buf

  (
    g1042_n_spl_,
    g1042_n
  );


  buf

  (
    g757_n_spl_,
    g757_n
  );


  buf

  (
    g981_n_spl_,
    g981_n
  );


  buf

  (
    g1037_n_spl_,
    g1037_n
  );


  buf

  (
    g761_n_spl_,
    g761_n
  );


  buf

  (
    g813_n_spl_,
    g813_n
  );


  buf

  (
    g822_n_spl_,
    g822_n
  );


  buf

  (
    g765_n_spl_,
    g765_n
  );


  buf

  (
    g884_n_spl_,
    g884_n
  );


  buf

  (
    G2759_o2_n_spl_,
    G2759_o2_n
  );


  buf

  (
    G2666_o2_p_spl_,
    G2666_o2_p
  );


  buf

  (
    G2759_o2_p_spl_,
    G2759_o2_p
  );


  buf

  (
    G2666_o2_n_spl_,
    G2666_o2_n
  );


  buf

  (
    g1094_p_spl_,
    g1094_p
  );


  buf

  (
    G1529_o2_p_spl_,
    G1529_o2_p
  );


  buf

  (
    G1529_o2_p_spl_0,
    G1529_o2_p_spl_
  );


  buf

  (
    G1538_o2_p_spl_,
    G1538_o2_p
  );


  buf

  (
    G1538_o2_p_spl_0,
    G1538_o2_p_spl_
  );


  buf

  (
    G1547_o2_n_spl_,
    G1547_o2_n
  );


  buf

  (
    G1547_o2_n_spl_0,
    G1547_o2_n_spl_
  );


  buf

  (
    G1556_o2_p_spl_,
    G1556_o2_p
  );


  buf

  (
    G1556_o2_p_spl_0,
    G1556_o2_p_spl_
  );


  buf

  (
    G1565_o2_p_spl_,
    G1565_o2_p
  );


  buf

  (
    G1565_o2_p_spl_0,
    G1565_o2_p_spl_
  );


  buf

  (
    G1574_o2_p_spl_,
    G1574_o2_p
  );


  buf

  (
    G1574_o2_p_spl_0,
    G1574_o2_p_spl_
  );


  buf

  (
    G1583_o2_n_spl_,
    G1583_o2_n
  );


  buf

  (
    G1583_o2_n_spl_0,
    G1583_o2_n_spl_
  );


  buf

  (
    G1592_o2_p_spl_,
    G1592_o2_p
  );


  buf

  (
    G1592_o2_p_spl_0,
    G1592_o2_p_spl_
  );


  buf

  (
    n1929_lo_n_spl_,
    n1929_lo_n
  );


  buf

  (
    G1601_o2_p_spl_,
    G1601_o2_p
  );


  buf

  (
    G1601_o2_p_spl_0,
    G1601_o2_p_spl_
  );


  buf

  (
    G1610_o2_p_spl_,
    G1610_o2_p
  );


  buf

  (
    G1610_o2_p_spl_0,
    G1610_o2_p_spl_
  );


  buf

  (
    G1619_o2_n_spl_,
    G1619_o2_n
  );


  buf

  (
    G1619_o2_n_spl_0,
    G1619_o2_n_spl_
  );


  buf

  (
    G1628_o2_p_spl_,
    G1628_o2_p
  );


  buf

  (
    G1628_o2_p_spl_0,
    G1628_o2_p_spl_
  );


  buf

  (
    G1637_o2_p_spl_,
    G1637_o2_p
  );


  buf

  (
    G1637_o2_p_spl_0,
    G1637_o2_p_spl_
  );


  buf

  (
    G1646_o2_p_spl_,
    G1646_o2_p
  );


  buf

  (
    G1646_o2_p_spl_0,
    G1646_o2_p_spl_
  );


  buf

  (
    G1655_o2_n_spl_,
    G1655_o2_n
  );


  buf

  (
    G1655_o2_n_spl_0,
    G1655_o2_n_spl_
  );


  buf

  (
    G1664_o2_p_spl_,
    G1664_o2_p
  );


  buf

  (
    G1664_o2_p_spl_0,
    G1664_o2_p_spl_
  );


  buf

  (
    n861_inv_n_spl_,
    n861_inv_n
  );


  buf

  (
    g827_p_spl_,
    g827_p
  );


  buf

  (
    g826_p_spl_,
    g826_p
  );


  buf

  (
    g1032_p_spl_,
    g1032_p
  );


  buf

  (
    G1738_o2_p_spl_,
    G1738_o2_p
  );


  buf

  (
    G1733_o2_p_spl_,
    G1733_o2_p
  );


  buf

  (
    G1738_o2_n_spl_,
    G1738_o2_n
  );


  buf

  (
    G1733_o2_n_spl_,
    G1733_o2_n
  );


  buf

  (
    G1751_o2_p_spl_,
    G1751_o2_p
  );


  buf

  (
    G1751_o2_n_spl_,
    G1751_o2_n
  );


  buf

  (
    G1764_o2_p_spl_,
    G1764_o2_p
  );


  buf

  (
    G1764_o2_n_spl_,
    G1764_o2_n
  );


  buf

  (
    G615_o2_p_spl_,
    G615_o2_p
  );


  buf

  (
    G615_o2_n_spl_,
    G615_o2_n
  );


  buf

  (
    g1052_p_spl_,
    g1052_p
  );


  buf

  (
    g1237_n_spl_,
    g1237_n
  );


  buf

  (
    g1059_n_spl_,
    g1059_n
  );


  buf

  (
    g1184_n_spl_,
    g1184_n
  );


  buf

  (
    g1232_n_spl_,
    g1232_n
  );


  buf

  (
    g1078_n_spl_,
    g1078_n
  );


  buf

  (
    g1142_n_spl_,
    g1142_n
  );


  buf

  (
    g1238_n_spl_,
    g1238_n
  );


  buf

  (
    g1095_n_spl_,
    g1095_n
  );


  buf

  (
    g1226_n_spl_,
    g1226_n
  );


  buf

  (
    g1259_n_spl_,
    g1259_n
  );


  buf

  (
    g1261_n_spl_,
    g1261_n
  );


  buf

  (
    g1263_n_spl_,
    g1263_n
  );


  buf

  (
    n1554_inv_n_spl_,
    n1554_inv_n
  );


  buf

  (
    G2027_o2_n_spl_,
    G2027_o2_n
  );


  buf

  (
    n1554_inv_p_spl_,
    n1554_inv_p
  );


  buf

  (
    n1554_inv_p_spl_0,
    n1554_inv_p_spl_
  );


  buf

  (
    G2027_o2_p_spl_,
    G2027_o2_p
  );


  buf

  (
    G2027_o2_p_spl_0,
    G2027_o2_p_spl_
  );


  buf

  (
    g1274_n_spl_,
    g1274_n
  );


  buf

  (
    g1273_n_spl_,
    g1273_n
  );


  buf

  (
    g1274_p_spl_,
    g1274_p
  );


  buf

  (
    g1274_p_spl_0,
    g1274_p_spl_
  );


  buf

  (
    g1273_p_spl_,
    g1273_p
  );


  buf

  (
    g1273_p_spl_0,
    g1273_p_spl_
  );


  buf

  (
    g1273_p_spl_1,
    g1273_p_spl_
  );


  buf

  (
    g1270_n_spl_,
    g1270_n
  );


  buf

  (
    g1275_p_spl_,
    g1275_p
  );


  buf

  (
    g1270_p_spl_,
    g1270_p
  );


  buf

  (
    n2097_lo_buf_o2_p_spl_,
    n2097_lo_buf_o2_p
  );


  buf

  (
    n2097_lo_buf_o2_p_spl_0,
    n2097_lo_buf_o2_p_spl_
  );


  buf

  (
    n5326_o2_n_spl_,
    n5326_o2_n
  );


  buf

  (
    n2097_lo_buf_o2_n_spl_,
    n2097_lo_buf_o2_n
  );


  buf

  (
    n5326_o2_p_spl_,
    n5326_o2_p
  );


  buf

  (
    n5326_o2_p_spl_0,
    n5326_o2_p_spl_
  );


  buf

  (
    n2133_lo_buf_o2_n_spl_,
    n2133_lo_buf_o2_n
  );


  buf

  (
    n5327_o2_p_spl_,
    n5327_o2_p
  );


  buf

  (
    n5327_o2_p_spl_0,
    n5327_o2_p_spl_
  );


  buf

  (
    n2133_lo_buf_o2_p_spl_,
    n2133_lo_buf_o2_p
  );


  buf

  (
    n2133_lo_buf_o2_p_spl_0,
    n2133_lo_buf_o2_p_spl_
  );


  buf

  (
    n5327_o2_n_spl_,
    n5327_o2_n
  );


  buf

  (
    g1074_n_spl_,
    g1074_n
  );


  buf

  (
    g1074_n_spl_0,
    g1074_n_spl_
  );


  buf

  (
    g1045_n_spl_,
    g1045_n
  );


  buf

  (
    g1045_n_spl_0,
    g1045_n_spl_
  );


  buf

  (
    g1045_n_spl_00,
    g1045_n_spl_0
  );


  buf

  (
    g1045_n_spl_01,
    g1045_n_spl_0
  );


  buf

  (
    g1045_n_spl_1,
    g1045_n_spl_
  );


  buf

  (
    g1269_n_spl_,
    g1269_n
  );


  buf

  (
    n1557_inv_n_spl_,
    n1557_inv_n
  );


  buf

  (
    G2393_o2_n_spl_,
    G2393_o2_n
  );


  buf

  (
    n1557_inv_p_spl_,
    n1557_inv_p
  );


  buf

  (
    n1557_inv_p_spl_0,
    n1557_inv_p_spl_
  );


  buf

  (
    G2393_o2_p_spl_,
    G2393_o2_p
  );


  buf

  (
    G2393_o2_p_spl_0,
    G2393_o2_p_spl_
  );


  buf

  (
    g1289_p_spl_,
    g1289_p
  );


  buf

  (
    g1288_p_spl_,
    g1288_p
  );


  buf

  (
    g1288_p_spl_0,
    g1288_p_spl_
  );


  buf

  (
    g1289_n_spl_,
    g1289_n
  );


  buf

  (
    g1288_n_spl_,
    g1288_n
  );


  buf

  (
    g1288_n_spl_0,
    g1288_n_spl_
  );


  buf

  (
    g1288_n_spl_1,
    g1288_n_spl_
  );


  buf

  (
    G2577_o2_n_spl_,
    G2577_o2_n
  );


  buf

  (
    G2281_o2_n_spl_,
    G2281_o2_n
  );


  buf

  (
    G2577_o2_p_spl_,
    G2577_o2_p
  );


  buf

  (
    G2281_o2_p_spl_,
    G2281_o2_p
  );


  buf

  (
    g1293_p_spl_,
    g1293_p
  );


  buf

  (
    g1293_p_spl_0,
    g1293_p_spl_
  );


  buf

  (
    g1293_p_spl_1,
    g1293_p_spl_
  );


  buf

  (
    g1293_n_spl_,
    g1293_n
  );


  buf

  (
    g1293_n_spl_0,
    g1293_n_spl_
  );


  buf

  (
    g1293_n_spl_00,
    g1293_n_spl_0
  );


  buf

  (
    g1293_n_spl_01,
    g1293_n_spl_0
  );


  buf

  (
    g1293_n_spl_1,
    g1293_n_spl_
  );


  buf

  (
    g1295_p_spl_,
    g1295_p
  );


  buf

  (
    g1294_n_spl_,
    g1294_n
  );


  buf

  (
    g1294_n_spl_0,
    g1294_n_spl_
  );


  buf

  (
    g1295_n_spl_,
    g1295_n
  );


  buf

  (
    g1294_p_spl_,
    g1294_p
  );


  buf

  (
    g1294_p_spl_0,
    g1294_p_spl_
  );


  buf

  (
    g1055_p_spl_,
    g1055_p
  );


  buf

  (
    g1055_p_spl_0,
    g1055_p_spl_
  );


  buf

  (
    g1055_p_spl_1,
    g1055_p_spl_
  );


  buf

  (
    g1055_n_spl_,
    g1055_n
  );


  buf

  (
    g1055_n_spl_0,
    g1055_n_spl_
  );


  buf

  (
    g1055_n_spl_00,
    g1055_n_spl_0
  );


  buf

  (
    g1055_n_spl_1,
    g1055_n_spl_
  );


  buf

  (
    g1045_p_spl_,
    g1045_p
  );


  buf

  (
    g1045_p_spl_0,
    g1045_p_spl_
  );


  buf

  (
    g1045_p_spl_00,
    g1045_p_spl_0
  );


  buf

  (
    g1045_p_spl_1,
    g1045_p_spl_
  );


  buf

  (
    n4921_o2_p_spl_,
    n4921_o2_p
  );


  buf

  (
    n4920_o2_p_spl_,
    n4920_o2_p
  );


  buf

  (
    n4920_o2_p_spl_0,
    n4920_o2_p_spl_
  );


  buf

  (
    g1302_p_spl_,
    g1302_p
  );


  buf

  (
    g1254_p_spl_,
    g1254_p
  );


  buf

  (
    g1254_p_spl_0,
    g1254_p_spl_
  );


  buf

  (
    g1256_p_spl_,
    g1256_p
  );


  buf

  (
    g1256_p_spl_0,
    g1256_p_spl_
  );


  buf

  (
    G1189_o2_p_spl_,
    G1189_o2_p
  );


  buf

  (
    G1189_o2_n_spl_,
    G1189_o2_n
  );


  buf

  (
    g1305_n_spl_,
    g1305_n
  );


  buf

  (
    g1305_p_spl_,
    g1305_p
  );


  buf

  (
    g1305_p_spl_0,
    g1305_p_spl_
  );


  buf

  (
    n1761_lo_buf_o2_p_spl_,
    n1761_lo_buf_o2_p
  );


  buf

  (
    n1761_lo_buf_o2_p_spl_0,
    n1761_lo_buf_o2_p_spl_
  );


  buf

  (
    n1761_lo_buf_o2_p_spl_1,
    n1761_lo_buf_o2_p_spl_
  );


  buf

  (
    n1749_lo_buf_o2_p_spl_,
    n1749_lo_buf_o2_p
  );


  buf

  (
    n1749_lo_buf_o2_p_spl_0,
    n1749_lo_buf_o2_p_spl_
  );


  buf

  (
    n1749_lo_buf_o2_p_spl_00,
    n1749_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1749_lo_buf_o2_p_spl_01,
    n1749_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1749_lo_buf_o2_p_spl_1,
    n1749_lo_buf_o2_p_spl_
  );


  buf

  (
    n1749_lo_buf_o2_p_spl_10,
    n1749_lo_buf_o2_p_spl_1
  );


  buf

  (
    n1749_lo_buf_o2_p_spl_11,
    n1749_lo_buf_o2_p_spl_1
  );


  buf

  (
    n1749_lo_buf_o2_n_spl_,
    n1749_lo_buf_o2_n
  );


  buf

  (
    n1749_lo_buf_o2_n_spl_0,
    n1749_lo_buf_o2_n_spl_
  );


  buf

  (
    n1749_lo_buf_o2_n_spl_00,
    n1749_lo_buf_o2_n_spl_0
  );


  buf

  (
    n1749_lo_buf_o2_n_spl_01,
    n1749_lo_buf_o2_n_spl_0
  );


  buf

  (
    n1749_lo_buf_o2_n_spl_1,
    n1749_lo_buf_o2_n_spl_
  );


  buf

  (
    g1309_p_spl_,
    g1309_p
  );


  buf

  (
    g1309_p_spl_0,
    g1309_p_spl_
  );


  buf

  (
    g1309_n_spl_,
    g1309_n
  );


  buf

  (
    g1309_n_spl_0,
    g1309_n_spl_
  );


  buf

  (
    n1809_lo_buf_o2_n_spl_,
    n1809_lo_buf_o2_n
  );


  buf

  (
    n1809_lo_buf_o2_p_spl_,
    n1809_lo_buf_o2_p
  );


  buf

  (
    n1809_lo_buf_o2_p_spl_0,
    n1809_lo_buf_o2_p_spl_
  );


  buf

  (
    g1310_n_spl_,
    g1310_n
  );


  buf

  (
    g1310_n_spl_0,
    g1310_n_spl_
  );


  buf

  (
    g1310_n_spl_00,
    g1310_n_spl_0
  );


  buf

  (
    g1310_n_spl_000,
    g1310_n_spl_00
  );


  buf

  (
    g1310_n_spl_01,
    g1310_n_spl_0
  );


  buf

  (
    g1310_n_spl_1,
    g1310_n_spl_
  );


  buf

  (
    g1310_n_spl_10,
    g1310_n_spl_1
  );


  buf

  (
    g1310_n_spl_11,
    g1310_n_spl_1
  );


  buf

  (
    n2139_lo_buf_o2_p_spl_,
    n2139_lo_buf_o2_p
  );


  buf

  (
    n2139_lo_buf_o2_p_spl_0,
    n2139_lo_buf_o2_p_spl_
  );


  buf

  (
    n2139_lo_buf_o2_p_spl_1,
    n2139_lo_buf_o2_p_spl_
  );


  buf

  (
    g1310_p_spl_,
    g1310_p
  );


  buf

  (
    g1310_p_spl_0,
    g1310_p_spl_
  );


  buf

  (
    g1310_p_spl_00,
    g1310_p_spl_0
  );


  buf

  (
    g1310_p_spl_01,
    g1310_p_spl_0
  );


  buf

  (
    g1310_p_spl_1,
    g1310_p_spl_
  );


  buf

  (
    g1310_p_spl_10,
    g1310_p_spl_1
  );


  buf

  (
    n2139_lo_buf_o2_n_spl_,
    n2139_lo_buf_o2_n
  );


  buf

  (
    n2139_lo_buf_o2_n_spl_0,
    n2139_lo_buf_o2_n_spl_
  );


  buf

  (
    g1311_n_spl_,
    g1311_n
  );


  buf

  (
    g1311_p_spl_,
    g1311_p
  );


  buf

  (
    n2187_lo_buf_o2_p_spl_,
    n2187_lo_buf_o2_p
  );


  buf

  (
    n2187_lo_buf_o2_n_spl_,
    n2187_lo_buf_o2_n
  );


  buf

  (
    g1314_p_spl_,
    g1314_p
  );


  buf

  (
    g1314_n_spl_,
    g1314_n
  );


  buf

  (
    n1899_lo_buf_o2_p_spl_,
    n1899_lo_buf_o2_p
  );


  buf

  (
    n1899_lo_buf_o2_p_spl_0,
    n1899_lo_buf_o2_p_spl_
  );


  buf

  (
    n1899_lo_buf_o2_p_spl_00,
    n1899_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1899_lo_buf_o2_p_spl_01,
    n1899_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1899_lo_buf_o2_p_spl_1,
    n1899_lo_buf_o2_p_spl_
  );


  buf

  (
    G831_o2_n_spl_,
    G831_o2_n
  );


  buf

  (
    G831_o2_n_spl_0,
    G831_o2_n_spl_
  );


  buf

  (
    G831_o2_n_spl_00,
    G831_o2_n_spl_0
  );


  buf

  (
    G831_o2_n_spl_01,
    G831_o2_n_spl_0
  );


  buf

  (
    G831_o2_n_spl_1,
    G831_o2_n_spl_
  );


  buf

  (
    G831_o2_n_spl_10,
    G831_o2_n_spl_1
  );


  buf

  (
    G831_o2_n_spl_11,
    G831_o2_n_spl_1
  );


  buf

  (
    n1899_lo_buf_o2_n_spl_,
    n1899_lo_buf_o2_n
  );


  buf

  (
    n1899_lo_buf_o2_n_spl_0,
    n1899_lo_buf_o2_n_spl_
  );


  buf

  (
    n1899_lo_buf_o2_n_spl_00,
    n1899_lo_buf_o2_n_spl_0
  );


  buf

  (
    n1899_lo_buf_o2_n_spl_1,
    n1899_lo_buf_o2_n_spl_
  );


  buf

  (
    G831_o2_p_spl_,
    G831_o2_p
  );


  buf

  (
    G831_o2_p_spl_0,
    G831_o2_p_spl_
  );


  buf

  (
    G831_o2_p_spl_00,
    G831_o2_p_spl_0
  );


  buf

  (
    G831_o2_p_spl_01,
    G831_o2_p_spl_0
  );


  buf

  (
    G831_o2_p_spl_1,
    G831_o2_p_spl_
  );


  buf

  (
    n2121_lo_buf_o2_p_spl_,
    n2121_lo_buf_o2_p
  );


  buf

  (
    n2121_lo_buf_o2_p_spl_0,
    n2121_lo_buf_o2_p_spl_
  );


  buf

  (
    n2121_lo_buf_o2_p_spl_1,
    n2121_lo_buf_o2_p_spl_
  );


  buf

  (
    G594_o2_n_spl_,
    G594_o2_n
  );


  buf

  (
    G594_o2_n_spl_0,
    G594_o2_n_spl_
  );


  buf

  (
    G594_o2_n_spl_00,
    G594_o2_n_spl_0
  );


  buf

  (
    G594_o2_n_spl_01,
    G594_o2_n_spl_0
  );


  buf

  (
    G594_o2_n_spl_1,
    G594_o2_n_spl_
  );


  buf

  (
    G594_o2_n_spl_10,
    G594_o2_n_spl_1
  );


  buf

  (
    G594_o2_n_spl_11,
    G594_o2_n_spl_1
  );


  buf

  (
    n2121_lo_buf_o2_n_spl_,
    n2121_lo_buf_o2_n
  );


  buf

  (
    n2121_lo_buf_o2_n_spl_0,
    n2121_lo_buf_o2_n_spl_
  );


  buf

  (
    G594_o2_p_spl_,
    G594_o2_p
  );


  buf

  (
    G594_o2_p_spl_0,
    G594_o2_p_spl_
  );


  buf

  (
    G594_o2_p_spl_00,
    G594_o2_p_spl_0
  );


  buf

  (
    G594_o2_p_spl_01,
    G594_o2_p_spl_0
  );


  buf

  (
    G594_o2_p_spl_1,
    G594_o2_p_spl_
  );


  buf

  (
    g1318_p_spl_,
    g1318_p
  );


  buf

  (
    g1318_p_spl_0,
    g1318_p_spl_
  );


  buf

  (
    g1318_p_spl_00,
    g1318_p_spl_0
  );


  buf

  (
    g1318_p_spl_01,
    g1318_p_spl_0
  );


  buf

  (
    g1318_p_spl_1,
    g1318_p_spl_
  );


  buf

  (
    g1318_p_spl_10,
    g1318_p_spl_1
  );


  buf

  (
    n2127_lo_buf_o2_p_spl_,
    n2127_lo_buf_o2_p
  );


  buf

  (
    n2127_lo_buf_o2_p_spl_0,
    n2127_lo_buf_o2_p_spl_
  );


  buf

  (
    n2127_lo_buf_o2_p_spl_1,
    n2127_lo_buf_o2_p_spl_
  );


  buf

  (
    g1318_n_spl_,
    g1318_n
  );


  buf

  (
    g1318_n_spl_0,
    g1318_n_spl_
  );


  buf

  (
    g1318_n_spl_00,
    g1318_n_spl_0
  );


  buf

  (
    g1318_n_spl_1,
    g1318_n_spl_
  );


  buf

  (
    n2127_lo_buf_o2_n_spl_,
    n2127_lo_buf_o2_n
  );


  buf

  (
    n2127_lo_buf_o2_n_spl_0,
    n2127_lo_buf_o2_n_spl_
  );


  buf

  (
    G477_o2_n_spl_,
    G477_o2_n
  );


  buf

  (
    G477_o2_p_spl_,
    G477_o2_p
  );


  buf

  (
    n1797_lo_buf_o2_p_spl_,
    n1797_lo_buf_o2_p
  );


  buf

  (
    n2151_lo_buf_o2_p_spl_,
    n2151_lo_buf_o2_p
  );


  buf

  (
    n2151_lo_buf_o2_p_spl_0,
    n2151_lo_buf_o2_p_spl_
  );


  buf

  (
    n2151_lo_buf_o2_p_spl_1,
    n2151_lo_buf_o2_p_spl_
  );


  buf

  (
    n2151_lo_buf_o2_n_spl_,
    n2151_lo_buf_o2_n
  );


  buf

  (
    g1326_n_spl_,
    g1326_n
  );


  buf

  (
    g1326_n_spl_0,
    g1326_n_spl_
  );


  buf

  (
    g1326_n_spl_1,
    g1326_n_spl_
  );


  buf

  (
    g1326_p_spl_,
    g1326_p
  );


  buf

  (
    g1326_p_spl_0,
    g1326_p_spl_
  );


  buf

  (
    n2199_lo_buf_o2_p_spl_,
    n2199_lo_buf_o2_p
  );


  buf

  (
    n2199_lo_buf_o2_p_spl_0,
    n2199_lo_buf_o2_p_spl_
  );


  buf

  (
    n2199_lo_buf_o2_n_spl_,
    n2199_lo_buf_o2_n
  );


  buf

  (
    g1329_n_spl_,
    g1329_n
  );


  buf

  (
    g1329_p_spl_,
    g1329_p
  );


  buf

  (
    g1329_p_spl_0,
    g1329_p_spl_
  );


  buf

  (
    n2163_lo_p_spl_,
    n2163_lo_p
  );


  buf

  (
    n2163_lo_p_spl_0,
    n2163_lo_p_spl_
  );


  buf

  (
    n2211_lo_buf_o2_p_spl_,
    n2211_lo_buf_o2_p
  );


  buf

  (
    G501_o2_p_spl_,
    G501_o2_p
  );


  buf

  (
    G501_o2_p_spl_0,
    G501_o2_p_spl_
  );


  buf

  (
    G501_o2_p_spl_00,
    G501_o2_p_spl_0
  );


  buf

  (
    G501_o2_p_spl_000,
    G501_o2_p_spl_00
  );


  buf

  (
    G501_o2_p_spl_01,
    G501_o2_p_spl_0
  );


  buf

  (
    G501_o2_p_spl_1,
    G501_o2_p_spl_
  );


  buf

  (
    G501_o2_p_spl_10,
    G501_o2_p_spl_1
  );


  buf

  (
    G501_o2_p_spl_11,
    G501_o2_p_spl_1
  );


  buf

  (
    n1854_lo_buf_o2_p_spl_,
    n1854_lo_buf_o2_p
  );


  buf

  (
    n1854_lo_buf_o2_p_spl_0,
    n1854_lo_buf_o2_p_spl_
  );


  buf

  (
    n1854_lo_buf_o2_p_spl_00,
    n1854_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1854_lo_buf_o2_p_spl_01,
    n1854_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1854_lo_buf_o2_p_spl_1,
    n1854_lo_buf_o2_p_spl_
  );


  buf

  (
    n1854_lo_buf_o2_p_spl_10,
    n1854_lo_buf_o2_p_spl_1
  );


  buf

  (
    G501_o2_n_spl_,
    G501_o2_n
  );


  buf

  (
    G501_o2_n_spl_0,
    G501_o2_n_spl_
  );


  buf

  (
    G501_o2_n_spl_00,
    G501_o2_n_spl_0
  );


  buf

  (
    G501_o2_n_spl_01,
    G501_o2_n_spl_0
  );


  buf

  (
    G501_o2_n_spl_1,
    G501_o2_n_spl_
  );


  buf

  (
    G501_o2_n_spl_10,
    G501_o2_n_spl_1
  );


  buf

  (
    G501_o2_n_spl_11,
    G501_o2_n_spl_1
  );


  buf

  (
    n1854_lo_buf_o2_n_spl_,
    n1854_lo_buf_o2_n
  );


  buf

  (
    n1854_lo_buf_o2_n_spl_0,
    n1854_lo_buf_o2_n_spl_
  );


  buf

  (
    n1854_lo_buf_o2_n_spl_00,
    n1854_lo_buf_o2_n_spl_0
  );


  buf

  (
    n1854_lo_buf_o2_n_spl_1,
    n1854_lo_buf_o2_n_spl_
  );


  buf

  (
    n1869_lo_buf_o2_n_spl_,
    n1869_lo_buf_o2_n
  );


  buf

  (
    n1869_lo_buf_o2_n_spl_0,
    n1869_lo_buf_o2_n_spl_
  );


  buf

  (
    n1869_lo_buf_o2_n_spl_00,
    n1869_lo_buf_o2_n_spl_0
  );


  buf

  (
    n1869_lo_buf_o2_n_spl_01,
    n1869_lo_buf_o2_n_spl_0
  );


  buf

  (
    n1869_lo_buf_o2_n_spl_1,
    n1869_lo_buf_o2_n_spl_
  );


  buf

  (
    G667_o2_p_spl_,
    G667_o2_p
  );


  buf

  (
    G667_o2_p_spl_0,
    G667_o2_p_spl_
  );


  buf

  (
    G667_o2_p_spl_00,
    G667_o2_p_spl_0
  );


  buf

  (
    G667_o2_p_spl_000,
    G667_o2_p_spl_00
  );


  buf

  (
    G667_o2_p_spl_01,
    G667_o2_p_spl_0
  );


  buf

  (
    G667_o2_p_spl_1,
    G667_o2_p_spl_
  );


  buf

  (
    G667_o2_p_spl_10,
    G667_o2_p_spl_1
  );


  buf

  (
    G667_o2_p_spl_11,
    G667_o2_p_spl_1
  );


  buf

  (
    n1869_lo_buf_o2_p_spl_,
    n1869_lo_buf_o2_p
  );


  buf

  (
    n1869_lo_buf_o2_p_spl_0,
    n1869_lo_buf_o2_p_spl_
  );


  buf

  (
    n1869_lo_buf_o2_p_spl_00,
    n1869_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1869_lo_buf_o2_p_spl_01,
    n1869_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1869_lo_buf_o2_p_spl_1,
    n1869_lo_buf_o2_p_spl_
  );


  buf

  (
    n1869_lo_buf_o2_p_spl_10,
    n1869_lo_buf_o2_p_spl_1
  );


  buf

  (
    n1869_lo_buf_o2_p_spl_11,
    n1869_lo_buf_o2_p_spl_1
  );


  buf

  (
    G667_o2_n_spl_,
    G667_o2_n
  );


  buf

  (
    G667_o2_n_spl_0,
    G667_o2_n_spl_
  );


  buf

  (
    G667_o2_n_spl_00,
    G667_o2_n_spl_0
  );


  buf

  (
    G667_o2_n_spl_01,
    G667_o2_n_spl_0
  );


  buf

  (
    G667_o2_n_spl_1,
    G667_o2_n_spl_
  );


  buf

  (
    G667_o2_n_spl_10,
    G667_o2_n_spl_1
  );


  buf

  (
    G667_o2_n_spl_11,
    G667_o2_n_spl_1
  );


  buf

  (
    g1350_p_spl_,
    g1350_p
  );


  buf

  (
    g1350_p_spl_0,
    g1350_p_spl_
  );


  buf

  (
    g1350_p_spl_00,
    g1350_p_spl_0
  );


  buf

  (
    g1350_p_spl_01,
    g1350_p_spl_0
  );


  buf

  (
    g1350_p_spl_1,
    g1350_p_spl_
  );


  buf

  (
    g1350_p_spl_10,
    g1350_p_spl_1
  );


  buf

  (
    g1350_p_spl_11,
    g1350_p_spl_1
  );


  buf

  (
    n1833_lo_buf_o2_n_spl_,
    n1833_lo_buf_o2_n
  );


  buf

  (
    n1833_lo_buf_o2_n_spl_0,
    n1833_lo_buf_o2_n_spl_
  );


  buf

  (
    n1833_lo_buf_o2_n_spl_1,
    n1833_lo_buf_o2_n_spl_
  );


  buf

  (
    g1350_n_spl_,
    g1350_n
  );


  buf

  (
    g1350_n_spl_0,
    g1350_n_spl_
  );


  buf

  (
    g1350_n_spl_00,
    g1350_n_spl_0
  );


  buf

  (
    g1350_n_spl_01,
    g1350_n_spl_0
  );


  buf

  (
    g1350_n_spl_1,
    g1350_n_spl_
  );


  buf

  (
    g1350_n_spl_10,
    g1350_n_spl_1
  );


  buf

  (
    n1833_lo_buf_o2_p_spl_,
    n1833_lo_buf_o2_p
  );


  buf

  (
    n1833_lo_buf_o2_p_spl_0,
    n1833_lo_buf_o2_p_spl_
  );


  buf

  (
    n1833_lo_buf_o2_p_spl_00,
    n1833_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1833_lo_buf_o2_p_spl_01,
    n1833_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1833_lo_buf_o2_p_spl_1,
    n1833_lo_buf_o2_p_spl_
  );


  buf

  (
    n1773_lo_buf_o2_p_spl_,
    n1773_lo_buf_o2_p
  );


  buf

  (
    n1773_lo_buf_o2_p_spl_0,
    n1773_lo_buf_o2_p_spl_
  );


  buf

  (
    n1773_lo_buf_o2_p_spl_00,
    n1773_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1773_lo_buf_o2_p_spl_1,
    n1773_lo_buf_o2_p_spl_
  );


  buf

  (
    n1773_lo_buf_o2_n_spl_,
    n1773_lo_buf_o2_n
  );


  buf

  (
    n1785_lo_buf_o2_p_spl_,
    n1785_lo_buf_o2_p
  );


  buf

  (
    n1785_lo_buf_o2_p_spl_0,
    n1785_lo_buf_o2_p_spl_
  );


  buf

  (
    n1785_lo_buf_o2_n_spl_,
    n1785_lo_buf_o2_n
  );


  buf

  (
    g1356_n_spl_,
    g1356_n
  );


  buf

  (
    g1356_n_spl_0,
    g1356_n_spl_
  );


  buf

  (
    g1356_n_spl_00,
    g1356_n_spl_0
  );


  buf

  (
    g1356_n_spl_000,
    g1356_n_spl_00
  );


  buf

  (
    g1356_n_spl_01,
    g1356_n_spl_0
  );


  buf

  (
    g1356_n_spl_1,
    g1356_n_spl_
  );


  buf

  (
    g1356_n_spl_10,
    g1356_n_spl_1
  );


  buf

  (
    g1356_n_spl_11,
    g1356_n_spl_1
  );


  buf

  (
    g1356_p_spl_,
    g1356_p
  );


  buf

  (
    g1356_p_spl_0,
    g1356_p_spl_
  );


  buf

  (
    g1356_p_spl_00,
    g1356_p_spl_0
  );


  buf

  (
    g1356_p_spl_01,
    g1356_p_spl_0
  );


  buf

  (
    g1356_p_spl_1,
    g1356_p_spl_
  );


  buf

  (
    g1356_p_spl_10,
    g1356_p_spl_1
  );


  buf

  (
    g1356_p_spl_11,
    g1356_p_spl_1
  );


  buf

  (
    g1358_p_spl_,
    g1358_p
  );


  buf

  (
    g1358_p_spl_0,
    g1358_p_spl_
  );


  buf

  (
    g1358_p_spl_00,
    g1358_p_spl_0
  );


  buf

  (
    g1358_p_spl_000,
    g1358_p_spl_00
  );


  buf

  (
    g1358_p_spl_01,
    g1358_p_spl_0
  );


  buf

  (
    g1358_p_spl_1,
    g1358_p_spl_
  );


  buf

  (
    g1358_p_spl_10,
    g1358_p_spl_1
  );


  buf

  (
    g1358_p_spl_11,
    g1358_p_spl_1
  );


  buf

  (
    g1358_n_spl_,
    g1358_n
  );


  buf

  (
    g1358_n_spl_0,
    g1358_n_spl_
  );


  buf

  (
    g1358_n_spl_00,
    g1358_n_spl_0
  );


  buf

  (
    g1358_n_spl_01,
    g1358_n_spl_0
  );


  buf

  (
    g1358_n_spl_1,
    g1358_n_spl_
  );


  buf

  (
    g1358_n_spl_10,
    g1358_n_spl_1
  );


  buf

  (
    g1358_n_spl_11,
    g1358_n_spl_1
  );


  buf

  (
    g1360_n_spl_,
    g1360_n
  );


  buf

  (
    g1360_n_spl_0,
    g1360_n_spl_
  );


  buf

  (
    g1360_n_spl_1,
    g1360_n_spl_
  );


  buf

  (
    g1360_p_spl_,
    g1360_p
  );


  buf

  (
    g1360_p_spl_0,
    g1360_p_spl_
  );


  buf

  (
    g1361_p_spl_,
    g1361_p
  );


  buf

  (
    g1361_p_spl_0,
    g1361_p_spl_
  );


  buf

  (
    g1361_p_spl_00,
    g1361_p_spl_0
  );


  buf

  (
    g1361_p_spl_01,
    g1361_p_spl_0
  );


  buf

  (
    g1361_p_spl_1,
    g1361_p_spl_
  );


  buf

  (
    g1361_p_spl_10,
    g1361_p_spl_1
  );


  buf

  (
    g1361_p_spl_11,
    g1361_p_spl_1
  );


  buf

  (
    g1361_n_spl_,
    g1361_n
  );


  buf

  (
    g1361_n_spl_0,
    g1361_n_spl_
  );


  buf

  (
    g1361_n_spl_00,
    g1361_n_spl_0
  );


  buf

  (
    g1361_n_spl_01,
    g1361_n_spl_0
  );


  buf

  (
    g1361_n_spl_1,
    g1361_n_spl_
  );


  buf

  (
    g1361_n_spl_10,
    g1361_n_spl_1
  );


  buf

  (
    g1366_n_spl_,
    g1366_n
  );


  buf

  (
    g1366_n_spl_0,
    g1366_n_spl_
  );


  buf

  (
    g1366_n_spl_00,
    g1366_n_spl_0
  );


  buf

  (
    g1366_n_spl_000,
    g1366_n_spl_00
  );


  buf

  (
    g1366_n_spl_01,
    g1366_n_spl_0
  );


  buf

  (
    g1366_n_spl_1,
    g1366_n_spl_
  );


  buf

  (
    g1366_n_spl_10,
    g1366_n_spl_1
  );


  buf

  (
    g1366_n_spl_11,
    g1366_n_spl_1
  );


  buf

  (
    g1366_p_spl_,
    g1366_p
  );


  buf

  (
    g1366_p_spl_0,
    g1366_p_spl_
  );


  buf

  (
    g1366_p_spl_00,
    g1366_p_spl_0
  );


  buf

  (
    g1366_p_spl_01,
    g1366_p_spl_0
  );


  buf

  (
    g1366_p_spl_1,
    g1366_p_spl_
  );


  buf

  (
    g1366_p_spl_10,
    g1366_p_spl_1
  );


  buf

  (
    g1367_n_spl_,
    g1367_n
  );


  buf

  (
    g1367_n_spl_0,
    g1367_n_spl_
  );


  buf

  (
    g1367_n_spl_00,
    g1367_n_spl_0
  );


  buf

  (
    g1367_n_spl_1,
    g1367_n_spl_
  );


  buf

  (
    g1367_p_spl_,
    g1367_p
  );


  buf

  (
    g1367_p_spl_0,
    g1367_p_spl_
  );


  buf

  (
    g1367_p_spl_1,
    g1367_p_spl_
  );


  buf

  (
    n1893_lo_buf_o2_p_spl_,
    n1893_lo_buf_o2_p
  );


  buf

  (
    n1893_lo_buf_o2_p_spl_0,
    n1893_lo_buf_o2_p_spl_
  );


  buf

  (
    n1893_lo_buf_o2_p_spl_00,
    n1893_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1893_lo_buf_o2_p_spl_01,
    n1893_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1893_lo_buf_o2_p_spl_1,
    n1893_lo_buf_o2_p_spl_
  );


  buf

  (
    n1893_lo_buf_o2_p_spl_10,
    n1893_lo_buf_o2_p_spl_1
  );


  buf

  (
    n1893_lo_buf_o2_p_spl_11,
    n1893_lo_buf_o2_p_spl_1
  );


  buf

  (
    n1893_lo_buf_o2_n_spl_,
    n1893_lo_buf_o2_n
  );


  buf

  (
    n1893_lo_buf_o2_n_spl_0,
    n1893_lo_buf_o2_n_spl_
  );


  buf

  (
    n1893_lo_buf_o2_n_spl_00,
    n1893_lo_buf_o2_n_spl_0
  );


  buf

  (
    n1893_lo_buf_o2_n_spl_01,
    n1893_lo_buf_o2_n_spl_0
  );


  buf

  (
    n1893_lo_buf_o2_n_spl_1,
    n1893_lo_buf_o2_n_spl_
  );


  buf

  (
    n2109_lo_buf_o2_p_spl_,
    n2109_lo_buf_o2_p
  );


  buf

  (
    n2109_lo_buf_o2_p_spl_0,
    n2109_lo_buf_o2_p_spl_
  );


  buf

  (
    n2109_lo_buf_o2_p_spl_1,
    n2109_lo_buf_o2_p_spl_
  );


  buf

  (
    n2109_lo_buf_o2_n_spl_,
    n2109_lo_buf_o2_n
  );


  buf

  (
    n2109_lo_buf_o2_n_spl_0,
    n2109_lo_buf_o2_n_spl_
  );


  buf

  (
    g1371_n_spl_,
    g1371_n
  );


  buf

  (
    g1371_n_spl_0,
    g1371_n_spl_
  );


  buf

  (
    g1371_p_spl_,
    g1371_p
  );


  buf

  (
    g1371_p_spl_0,
    g1371_p_spl_
  );


  buf

  (
    g1371_p_spl_1,
    g1371_p_spl_
  );


  buf

  (
    g1365_p_spl_,
    g1365_p
  );


  buf

  (
    g1365_p_spl_0,
    g1365_p_spl_
  );


  buf

  (
    g1365_p_spl_00,
    g1365_p_spl_0
  );


  buf

  (
    g1365_p_spl_1,
    g1365_p_spl_
  );


  buf

  (
    n2007_lo_n_spl_,
    n2007_lo_n
  );


  buf

  (
    n2007_lo_n_spl_0,
    n2007_lo_n_spl_
  );


  buf

  (
    n2007_lo_n_spl_00,
    n2007_lo_n_spl_0
  );


  buf

  (
    n2007_lo_n_spl_01,
    n2007_lo_n_spl_0
  );


  buf

  (
    n2007_lo_n_spl_1,
    n2007_lo_n_spl_
  );


  buf

  (
    g1379_n_spl_,
    g1379_n
  );


  buf

  (
    n2019_lo_n_spl_,
    n2019_lo_n
  );


  buf

  (
    n2019_lo_n_spl_0,
    n2019_lo_n_spl_
  );


  buf

  (
    n2019_lo_n_spl_00,
    n2019_lo_n_spl_0
  );


  buf

  (
    n2019_lo_n_spl_01,
    n2019_lo_n_spl_0
  );


  buf

  (
    n2019_lo_n_spl_1,
    n2019_lo_n_spl_
  );


  buf

  (
    g1252_p_spl_,
    g1252_p
  );


  buf

  (
    g1252_p_spl_0,
    g1252_p_spl_
  );


  buf

  (
    n1845_lo_buf_o2_n_spl_,
    n1845_lo_buf_o2_n
  );


  buf

  (
    n1845_lo_buf_o2_n_spl_0,
    n1845_lo_buf_o2_n_spl_
  );


  buf

  (
    n1845_lo_buf_o2_n_spl_00,
    n1845_lo_buf_o2_n_spl_0
  );


  buf

  (
    n1845_lo_buf_o2_n_spl_1,
    n1845_lo_buf_o2_n_spl_
  );


  buf

  (
    n1845_lo_buf_o2_p_spl_,
    n1845_lo_buf_o2_p
  );


  buf

  (
    n1845_lo_buf_o2_p_spl_0,
    n1845_lo_buf_o2_p_spl_
  );


  buf

  (
    n1845_lo_buf_o2_p_spl_00,
    n1845_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1845_lo_buf_o2_p_spl_01,
    n1845_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1845_lo_buf_o2_p_spl_1,
    n1845_lo_buf_o2_p_spl_
  );


  buf

  (
    n1845_lo_buf_o2_p_spl_10,
    n1845_lo_buf_o2_p_spl_1
  );


  buf

  (
    n1845_lo_buf_o2_p_spl_11,
    n1845_lo_buf_o2_p_spl_1
  );


  buf

  (
    n1815_lo_buf_o2_p_spl_,
    n1815_lo_buf_o2_p
  );


  buf

  (
    n1815_lo_buf_o2_p_spl_0,
    n1815_lo_buf_o2_p_spl_
  );


  buf

  (
    n1815_lo_buf_o2_p_spl_00,
    n1815_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1815_lo_buf_o2_p_spl_1,
    n1815_lo_buf_o2_p_spl_
  );


  buf

  (
    n1815_lo_buf_o2_n_spl_,
    n1815_lo_buf_o2_n
  );


  buf

  (
    n1881_lo_buf_o2_p_spl_,
    n1881_lo_buf_o2_p
  );


  buf

  (
    n1881_lo_buf_o2_p_spl_0,
    n1881_lo_buf_o2_p_spl_
  );


  buf

  (
    n1881_lo_buf_o2_p_spl_00,
    n1881_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1881_lo_buf_o2_p_spl_01,
    n1881_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1881_lo_buf_o2_p_spl_1,
    n1881_lo_buf_o2_p_spl_
  );


  buf

  (
    n1881_lo_buf_o2_p_spl_10,
    n1881_lo_buf_o2_p_spl_1
  );


  buf

  (
    n1881_lo_buf_o2_p_spl_11,
    n1881_lo_buf_o2_p_spl_1
  );


  buf

  (
    n1881_lo_buf_o2_n_spl_,
    n1881_lo_buf_o2_n
  );


  buf

  (
    n1881_lo_buf_o2_n_spl_0,
    n1881_lo_buf_o2_n_spl_
  );


  buf

  (
    n1881_lo_buf_o2_n_spl_00,
    n1881_lo_buf_o2_n_spl_0
  );


  buf

  (
    n1881_lo_buf_o2_n_spl_01,
    n1881_lo_buf_o2_n_spl_0
  );


  buf

  (
    n1881_lo_buf_o2_n_spl_1,
    n1881_lo_buf_o2_n_spl_
  );


  buf

  (
    n2094_lo_buf_o2_p_spl_,
    n2094_lo_buf_o2_p
  );


  buf

  (
    n2094_lo_buf_o2_p_spl_0,
    n2094_lo_buf_o2_p_spl_
  );


  buf

  (
    n2094_lo_buf_o2_p_spl_1,
    n2094_lo_buf_o2_p_spl_
  );


  buf

  (
    n2094_lo_buf_o2_n_spl_,
    n2094_lo_buf_o2_n
  );


  buf

  (
    g1400_p_spl_,
    g1400_p
  );


  buf

  (
    g1400_p_spl_0,
    g1400_p_spl_
  );


  buf

  (
    g1400_p_spl_00,
    g1400_p_spl_0
  );


  buf

  (
    g1400_p_spl_1,
    g1400_p_spl_
  );


  buf

  (
    g1410_n_spl_,
    g1410_n
  );


  buf

  (
    g1425_n_spl_,
    g1425_n
  );


  buf

  (
    g1425_n_spl_0,
    g1425_n_spl_
  );


  buf

  (
    g1425_n_spl_1,
    g1425_n_spl_
  );


  buf

  (
    g1425_p_spl_,
    g1425_p
  );


  buf

  (
    g1425_p_spl_0,
    g1425_p_spl_
  );


  buf

  (
    g1425_p_spl_1,
    g1425_p_spl_
  );


  buf

  (
    n2175_lo_p_spl_,
    n2175_lo_p
  );


  buf

  (
    n2223_lo_p_spl_,
    n2223_lo_p
  );


  buf

  (
    n1995_lo_p_spl_,
    n1995_lo_p
  );


  buf

  (
    n2079_lo_buf_o2_p_spl_,
    n2079_lo_buf_o2_p
  );


  buf

  (
    g1466_p_spl_,
    g1466_p
  );


  buf

  (
    g1466_p_spl_0,
    g1466_p_spl_
  );


  buf

  (
    g1466_p_spl_00,
    g1466_p_spl_0
  );


  buf

  (
    g1466_p_spl_1,
    g1466_p_spl_
  );


  buf

  (
    g1476_n_spl_,
    g1476_n
  );


  buf

  (
    g1389_n_spl_,
    g1389_n
  );


  buf

  (
    g1481_n_spl_,
    g1481_n
  );


  buf

  (
    g1481_n_spl_0,
    g1481_n_spl_
  );


  buf

  (
    g1383_n_spl_,
    g1383_n
  );


  buf

  (
    g1381_n_spl_,
    g1381_n
  );


  buf

  (
    n2031_lo_p_spl_,
    n2031_lo_p
  );


  buf

  (
    n2031_lo_p_spl_0,
    n2031_lo_p_spl_
  );


  buf

  (
    n2031_lo_p_spl_1,
    n2031_lo_p_spl_
  );


  buf

  (
    g1379_p_spl_,
    g1379_p
  );


  buf

  (
    n2043_lo_p_spl_,
    n2043_lo_p
  );


  buf

  (
    n2043_lo_p_spl_0,
    n2043_lo_p_spl_
  );


  buf

  (
    n2043_lo_p_spl_1,
    n2043_lo_p_spl_
  );


  buf

  (
    g1252_n_spl_,
    g1252_n
  );


  buf

  (
    n2298_lo_n_spl_,
    n2298_lo_n
  );


  buf

  (
    n2298_lo_n_spl_0,
    n2298_lo_n_spl_
  );


  buf

  (
    n2298_lo_n_spl_00,
    n2298_lo_n_spl_0
  );


  buf

  (
    n2298_lo_n_spl_01,
    n2298_lo_n_spl_0
  );


  buf

  (
    n2298_lo_n_spl_1,
    n2298_lo_n_spl_
  );


  buf

  (
    n2298_lo_n_spl_10,
    n2298_lo_n_spl_1
  );


  buf

  (
    g1385_n_spl_,
    g1385_n
  );


  buf

  (
    n1905_lo_buf_o2_p_spl_,
    n1905_lo_buf_o2_p
  );


  buf

  (
    n1905_lo_buf_o2_p_spl_0,
    n1905_lo_buf_o2_p_spl_
  );


  buf

  (
    n1905_lo_buf_o2_p_spl_1,
    n1905_lo_buf_o2_p_spl_
  );


  buf

  (
    g1087_p_spl_,
    g1087_p
  );


  buf

  (
    g1087_p_spl_0,
    g1087_p_spl_
  );


  buf

  (
    g1081_n_spl_,
    g1081_n
  );


  buf

  (
    g1081_n_spl_0,
    g1081_n_spl_
  );


  buf

  (
    g1240_n_spl_,
    g1240_n
  );


  buf

  (
    g1240_n_spl_0,
    g1240_n_spl_
  );


  buf

  (
    g1083_p_spl_,
    g1083_p
  );


  buf

  (
    g1083_p_spl_0,
    g1083_p_spl_
  );


  buf

  (
    g1512_n_spl_,
    g1512_n
  );


  buf

  (
    g1512_p_spl_,
    g1512_p
  );


  buf

  (
    g1512_p_spl_0,
    g1512_p_spl_
  );


  buf

  (
    g1515_p_spl_,
    g1515_p
  );


  buf

  (
    g1515_p_spl_0,
    g1515_p_spl_
  );


  buf

  (
    g1515_p_spl_1,
    g1515_p_spl_
  );


  buf

  (
    g1386_n_spl_,
    g1386_n
  );


  buf

  (
    g1386_n_spl_0,
    g1386_n_spl_
  );


  buf

  (
    g1493_p_spl_,
    g1493_p
  );


  buf

  (
    g1452_n_spl_,
    g1452_n
  );


  buf

  (
    g1452_n_spl_0,
    g1452_n_spl_
  );


  buf

  (
    g1452_n_spl_00,
    g1452_n_spl_0
  );


  buf

  (
    g1452_n_spl_1,
    g1452_n_spl_
  );


  buf

  (
    g1482_n_spl_,
    g1482_n
  );


  buf

  (
    g1482_n_spl_0,
    g1482_n_spl_
  );


  buf

  (
    g1482_n_spl_00,
    g1482_n_spl_0
  );


  buf

  (
    g1482_n_spl_1,
    g1482_n_spl_
  );


  buf

  (
    g1308_p_spl_,
    g1308_p
  );


  buf

  (
    n2145_lo_buf_o2_p_spl_,
    n2145_lo_buf_o2_p
  );


  buf

  (
    n2157_lo_buf_o2_p_spl_,
    n2157_lo_buf_o2_p
  );


  buf

  (
    n2169_lo_buf_o2_p_spl_,
    n2169_lo_buf_o2_p
  );


  buf

  (
    n2181_lo_buf_o2_p_spl_,
    n2181_lo_buf_o2_p
  );


  buf

  (
    g1515_n_spl_,
    g1515_n
  );


  buf

  (
    g1515_n_spl_0,
    g1515_n_spl_
  );


  buf

  (
    g1276_p_spl_,
    g1276_p
  );


  buf

  (
    n5101_o2_p_spl_,
    n5101_o2_p
  );


  buf

  (
    n5101_o2_p_spl_0,
    n5101_o2_p_spl_
  );


  buf

  (
    n5267_o2_p_spl_,
    n5267_o2_p
  );


  buf

  (
    n5267_o2_p_spl_0,
    n5267_o2_p_spl_
  );


  buf

  (
    n5267_o2_p_spl_1,
    n5267_o2_p_spl_
  );


  buf

  (
    n5325_o2_p_spl_,
    n5325_o2_p
  );


  buf

  (
    n5325_o2_p_spl_0,
    n5325_o2_p_spl_
  );


  buf

  (
    n5325_o2_p_spl_1,
    n5325_o2_p_spl_
  );


  buf

  (
    g1542_n_spl_,
    g1542_n
  );


  buf

  (
    g1542_p_spl_,
    g1542_p
  );


  buf

  (
    g1542_p_spl_0,
    g1542_p_spl_
  );


  buf

  (
    n5294_o2_p_spl_,
    n5294_o2_p
  );


  buf

  (
    n5294_o2_p_spl_0,
    n5294_o2_p_spl_
  );


  buf

  (
    n5294_o2_p_spl_00,
    n5294_o2_p_spl_0
  );


  buf

  (
    n5294_o2_p_spl_1,
    n5294_o2_p_spl_
  );


  buf

  (
    n5294_o2_n_spl_,
    n5294_o2_n
  );


  buf

  (
    n5294_o2_n_spl_0,
    n5294_o2_n_spl_
  );


  buf

  (
    g1556_p_spl_,
    g1556_p
  );


  buf

  (
    g1556_p_spl_0,
    g1556_p_spl_
  );


  buf

  (
    g1557_n_spl_,
    g1557_n
  );


  buf

  (
    g1555_n_spl_,
    g1555_n
  );


  buf

  (
    g1555_n_spl_0,
    g1555_n_spl_
  );


  buf

  (
    g1555_n_spl_1,
    g1555_n_spl_
  );


  buf

  (
    g1555_p_spl_,
    g1555_p
  );


  buf

  (
    g1555_p_spl_0,
    g1555_p_spl_
  );


  buf

  (
    g1555_p_spl_1,
    g1555_p_spl_
  );


  buf

  (
    g1560_n_spl_,
    g1560_n
  );


  buf

  (
    g1561_p_spl_,
    g1561_p
  );


  buf

  (
    g1563_n_spl_,
    g1563_n
  );


  buf

  (
    g1565_n_spl_,
    g1565_n
  );


  buf

  (
    g1414_n_spl_,
    g1414_n
  );


  buf

  (
    g1412_n_spl_,
    g1412_n
  );


  buf

  (
    g1410_p_spl_,
    g1410_p
  );


  buf

  (
    n1857_lo_buf_o2_n_spl_,
    n1857_lo_buf_o2_n
  );


  buf

  (
    n1857_lo_buf_o2_n_spl_0,
    n1857_lo_buf_o2_n_spl_
  );


  buf

  (
    n5100_o2_n_spl_,
    n5100_o2_n
  );


  buf

  (
    n5100_o2_n_spl_0,
    n5100_o2_n_spl_
  );


  buf

  (
    g1507_n_spl_,
    g1507_n
  );


  buf

  (
    n1821_lo_buf_o2_p_spl_,
    n1821_lo_buf_o2_p
  );


  buf

  (
    n1821_lo_buf_o2_p_spl_0,
    n1821_lo_buf_o2_p_spl_
  );


  buf

  (
    n1821_lo_buf_o2_p_spl_00,
    n1821_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1821_lo_buf_o2_p_spl_1,
    n1821_lo_buf_o2_p_spl_
  );


  buf

  (
    n5266_o2_n_spl_,
    n5266_o2_n
  );


  buf

  (
    n5266_o2_n_spl_0,
    n5266_o2_n_spl_
  );


  buf

  (
    g1582_n_spl_,
    g1582_n
  );


  buf

  (
    g1504_n_spl_,
    g1504_n
  );


  buf

  (
    g1526_n_spl_,
    g1526_n
  );


  buf

  (
    g1526_n_spl_0,
    g1526_n_spl_
  );


  buf

  (
    g1526_n_spl_1,
    g1526_n_spl_
  );


  buf

  (
    g1524_n_spl_,
    g1524_n
  );


  buf

  (
    g1524_n_spl_0,
    g1524_n_spl_
  );


  buf

  (
    g1524_n_spl_1,
    g1524_n_spl_
  );


  buf

  (
    g1591_n_spl_,
    g1591_n
  );


  buf

  (
    g1591_n_spl_0,
    g1591_n_spl_
  );


  buf

  (
    g1586_n_spl_,
    g1586_n
  );


  buf

  (
    g1586_n_spl_0,
    g1586_n_spl_
  );


  buf

  (
    g1607_n_spl_,
    g1607_n
  );


  buf

  (
    g1607_n_spl_0,
    g1607_n_spl_
  );


  buf

  (
    g1607_n_spl_1,
    g1607_n_spl_
  );


  buf

  (
    n2007_lo_p_spl_,
    n2007_lo_p
  );


  buf

  (
    n2007_lo_p_spl_0,
    n2007_lo_p_spl_
  );


  buf

  (
    n2007_lo_p_spl_1,
    n2007_lo_p_spl_
  );


  buf

  (
    g1607_p_spl_,
    g1607_p
  );


  buf

  (
    g1607_p_spl_0,
    g1607_p_spl_
  );


  buf

  (
    g1607_p_spl_1,
    g1607_p_spl_
  );


  buf

  (
    g1347_p_spl_,
    g1347_p
  );


  buf

  (
    g1347_n_spl_,
    g1347_n
  );


  buf

  (
    g1347_n_spl_0,
    g1347_n_spl_
  );


  buf

  (
    g1347_n_spl_00,
    g1347_n_spl_0
  );


  buf

  (
    g1347_n_spl_1,
    g1347_n_spl_
  );


  buf

  (
    n2019_lo_p_spl_,
    n2019_lo_p
  );


  buf

  (
    n2019_lo_p_spl_0,
    n2019_lo_p_spl_
  );


  buf

  (
    n2019_lo_p_spl_00,
    n2019_lo_p_spl_0
  );


  buf

  (
    n2019_lo_p_spl_1,
    n2019_lo_p_spl_
  );


  buf

  (
    g1429_n_spl_,
    g1429_n
  );


  buf

  (
    g1429_n_spl_0,
    g1429_n_spl_
  );


  buf

  (
    g1429_n_spl_00,
    g1429_n_spl_0
  );


  buf

  (
    g1429_n_spl_1,
    g1429_n_spl_
  );


  buf

  (
    g1429_p_spl_,
    g1429_p
  );


  buf

  (
    g1429_p_spl_0,
    g1429_p_spl_
  );


  buf

  (
    g1337_p_spl_,
    g1337_p
  );


  buf

  (
    g1337_n_spl_,
    g1337_n
  );


  buf

  (
    g1337_n_spl_0,
    g1337_n_spl_
  );


  buf

  (
    g1337_n_spl_00,
    g1337_n_spl_0
  );


  buf

  (
    g1337_n_spl_1,
    g1337_n_spl_
  );


  buf

  (
    n5293_o2_p_spl_,
    n5293_o2_p
  );


  buf

  (
    n5292_o2_p_spl_,
    n5292_o2_p
  );


  buf

  (
    n5292_o2_p_spl_0,
    n5292_o2_p_spl_
  );


  buf

  (
    n5266_o2_p_spl_,
    n5266_o2_p
  );


  buf

  (
    n5266_o2_p_spl_0,
    n5266_o2_p_spl_
  );


  buf

  (
    n5266_o2_p_spl_00,
    n5266_o2_p_spl_0
  );


  buf

  (
    n5266_o2_p_spl_01,
    n5266_o2_p_spl_0
  );


  buf

  (
    n5266_o2_p_spl_1,
    n5266_o2_p_spl_
  );


  buf

  (
    n5100_o2_p_spl_,
    n5100_o2_p
  );


  buf

  (
    n5100_o2_p_spl_0,
    n5100_o2_p_spl_
  );


  buf

  (
    n5100_o2_p_spl_00,
    n5100_o2_p_spl_0
  );


  buf

  (
    n5100_o2_p_spl_01,
    n5100_o2_p_spl_0
  );


  buf

  (
    n5100_o2_p_spl_1,
    n5100_o2_p_spl_
  );


  buf

  (
    n1821_lo_buf_o2_n_spl_,
    n1821_lo_buf_o2_n
  );


  buf

  (
    n1821_lo_buf_o2_n_spl_0,
    n1821_lo_buf_o2_n_spl_
  );


  buf

  (
    g1506_n_spl_,
    g1506_n
  );


  buf

  (
    g1387_p_spl_,
    g1387_p
  );


  buf

  (
    n2298_lo_p_spl_,
    n2298_lo_p
  );


  buf

  (
    g1284_n_spl_,
    g1284_n
  );


  buf

  (
    g1522_n_spl_,
    g1522_n
  );


  buf

  (
    g1520_n_spl_,
    g1520_n
  );


  buf

  (
    n1857_lo_buf_o2_p_spl_,
    n1857_lo_buf_o2_p
  );


  buf

  (
    n1857_lo_buf_o2_p_spl_0,
    n1857_lo_buf_o2_p_spl_
  );


  buf

  (
    n1857_lo_buf_o2_p_spl_00,
    n1857_lo_buf_o2_p_spl_0
  );


  buf

  (
    n1857_lo_buf_o2_p_spl_1,
    n1857_lo_buf_o2_p_spl_
  );


  buf

  (
    g1079_n_spl_,
    g1079_n
  );


  buf

  (
    g1079_p_spl_,
    g1079_p
  );


  buf

  (
    g1079_p_spl_0,
    g1079_p_spl_
  );


  buf

  (
    g1301_n_spl_,
    g1301_n
  );


  buf

  (
    g1279_n_spl_,
    g1279_n
  );


  buf

  (
    g1282_n_spl_,
    g1282_n
  );


  buf

  (
    g1442_n_spl_,
    g1442_n
  );


  buf

  (
    g1442_n_spl_0,
    g1442_n_spl_
  );


  buf

  (
    g1442_n_spl_00,
    g1442_n_spl_0
  );


  buf

  (
    g1442_n_spl_1,
    g1442_n_spl_
  );


  buf

  (
    g1324_p_spl_,
    g1324_p
  );


  buf

  (
    n2031_lo_n_spl_,
    n2031_lo_n
  );


  buf

  (
    n2031_lo_n_spl_0,
    n2031_lo_n_spl_
  );


  buf

  (
    n2031_lo_n_spl_1,
    n2031_lo_n_spl_
  );


  buf

  (
    g1324_n_spl_,
    g1324_n
  );


  buf

  (
    g1324_n_spl_0,
    g1324_n_spl_
  );


  buf

  (
    n2043_lo_n_spl_,
    n2043_lo_n
  );


  buf

  (
    n2043_lo_n_spl_0,
    n2043_lo_n_spl_
  );


  buf

  (
    n2043_lo_n_spl_1,
    n2043_lo_n_spl_
  );


  buf

  (
    g1656_n_spl_,
    g1656_n
  );


  buf

  (
    g1612_n_spl_,
    g1612_n
  );


  buf

  (
    g1480_n_spl_,
    g1480_n
  );


  buf

  (
    g1478_n_spl_,
    g1478_n
  );


  buf

  (
    g1476_p_spl_,
    g1476_p
  );


  buf

  (
    g1617_n_spl_,
    g1617_n
  );


  buf

  (
    g1493_n_spl_,
    g1493_n
  );


  buf

  (
    g1493_n_spl_0,
    g1493_n_spl_
  );


  buf

  (
    g1493_n_spl_1,
    g1493_n_spl_
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G5_p_spl_0,
    G5_p_spl_
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_00,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_01,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_10,
    G4_p_spl_1
  );


  buf

  (
    G4_p_spl_11,
    G4_p_spl_1
  );


  buf

  (
    n1983_lo_p_spl_,
    n1983_lo_p
  );


  buf

  (
    g1685_n_spl_,
    g1685_n
  );


  buf

  (
    g1685_n_spl_0,
    g1685_n_spl_
  );


  buf

  (
    g1663_n_spl_,
    g1663_n
  );


  buf

  (
    g1663_n_spl_0,
    g1663_n_spl_
  );


  buf

  (
    g1663_n_spl_1,
    g1663_n_spl_
  );


  buf

  (
    g1625_p_spl_,
    g1625_p
  );


  buf

  (
    g1670_n_spl_,
    g1670_n
  );


  buf

  (
    g1670_n_spl_0,
    g1670_n_spl_
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    g1693_n_spl_,
    g1693_n
  );


  buf

  (
    g1693_n_spl_0,
    g1693_n_spl_
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G3_p_spl_0,
    G3_p_spl_
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    n5295_o2_p_spl_,
    n5295_o2_p
  );


  buf

  (
    n5295_o2_p_spl_0,
    n5295_o2_p_spl_
  );


  buf

  (
    n5295_o2_p_spl_00,
    n5295_o2_p_spl_0
  );


  buf

  (
    n5295_o2_p_spl_1,
    n5295_o2_p_spl_
  );


  buf

  (
    g1085_p_spl_,
    g1085_p
  );


  buf

  (
    g1085_p_spl_0,
    g1085_p_spl_
  );


  buf

  (
    g1085_p_spl_1,
    g1085_p_spl_
  );


  buf

  (
    g1258_p_spl_,
    g1258_p
  );


  buf

  (
    g1258_p_spl_0,
    g1258_p_spl_
  );


  buf

  (
    g1258_p_spl_1,
    g1258_p_spl_
  );


  buf

  (
    g1303_n_spl_,
    g1303_n
  );


  buf

  (
    g1304_n_spl_,
    g1304_n
  );


  buf

  (
    g1501_p_spl_,
    g1501_p
  );


  buf

  (
    g1501_p_spl_0,
    g1501_p_spl_
  );


  buf

  (
    g1501_p_spl_1,
    g1501_p_spl_
  );


  buf

  (
    g1517_n_spl_,
    g1517_n
  );


  buf

  (
    g1518_n_spl_,
    g1518_n
  );


  buf

  (
    g1523_n_spl_,
    g1523_n
  );


  buf

  (
    g1523_n_spl_0,
    g1523_n_spl_
  );


  buf

  (
    g1529_n_spl_,
    g1529_n
  );


  buf

  (
    g1532_n_spl_,
    g1532_n
  );


  buf

  (
    g1535_n_spl_,
    g1535_n
  );


  buf

  (
    g1538_n_spl_,
    g1538_n
  );


  buf

  (
    g1541_n_spl_,
    g1541_n
  );


  buf

  (
    g1554_n_spl_,
    g1554_n
  );


  buf

  (
    g1558_n_spl_,
    g1558_n
  );


  buf

  (
    g1558_n_spl_0,
    g1558_n_spl_
  );


  buf

  (
    g1558_n_spl_00,
    g1558_n_spl_0
  );


  buf

  (
    g1558_n_spl_000,
    g1558_n_spl_00
  );


  buf

  (
    g1558_n_spl_001,
    g1558_n_spl_00
  );


  buf

  (
    g1558_n_spl_01,
    g1558_n_spl_0
  );


  buf

  (
    g1558_n_spl_010,
    g1558_n_spl_01
  );


  buf

  (
    g1558_n_spl_011,
    g1558_n_spl_01
  );


  buf

  (
    g1558_n_spl_1,
    g1558_n_spl_
  );


  buf

  (
    g1558_n_spl_10,
    g1558_n_spl_1
  );


  buf

  (
    g1558_n_spl_11,
    g1558_n_spl_1
  );


  buf

  (
    g1559_n_spl_,
    g1559_n
  );


  buf

  (
    g1559_n_spl_0,
    g1559_n_spl_
  );


  buf

  (
    g1559_n_spl_00,
    g1559_n_spl_0
  );


  buf

  (
    g1559_n_spl_000,
    g1559_n_spl_00
  );


  buf

  (
    g1559_n_spl_001,
    g1559_n_spl_00
  );


  buf

  (
    g1559_n_spl_01,
    g1559_n_spl_0
  );


  buf

  (
    g1559_n_spl_010,
    g1559_n_spl_01
  );


  buf

  (
    g1559_n_spl_011,
    g1559_n_spl_01
  );


  buf

  (
    g1559_n_spl_1,
    g1559_n_spl_
  );


  buf

  (
    g1559_n_spl_10,
    g1559_n_spl_1
  );


  buf

  (
    g1559_n_spl_11,
    g1559_n_spl_1
  );


  buf

  (
    g1562_p_spl_,
    g1562_p
  );


  buf

  (
    g1562_p_spl_0,
    g1562_p_spl_
  );


  buf

  (
    g1562_p_spl_00,
    g1562_p_spl_0
  );


  buf

  (
    g1562_p_spl_000,
    g1562_p_spl_00
  );


  buf

  (
    g1562_p_spl_001,
    g1562_p_spl_00
  );


  buf

  (
    g1562_p_spl_01,
    g1562_p_spl_0
  );


  buf

  (
    g1562_p_spl_010,
    g1562_p_spl_01
  );


  buf

  (
    g1562_p_spl_011,
    g1562_p_spl_01
  );


  buf

  (
    g1562_p_spl_1,
    g1562_p_spl_
  );


  buf

  (
    g1562_p_spl_10,
    g1562_p_spl_1
  );


  buf

  (
    g1562_p_spl_11,
    g1562_p_spl_1
  );


  buf

  (
    g1564_n_spl_,
    g1564_n
  );


  buf

  (
    g1564_n_spl_0,
    g1564_n_spl_
  );


  buf

  (
    g1564_n_spl_00,
    g1564_n_spl_0
  );


  buf

  (
    g1564_n_spl_000,
    g1564_n_spl_00
  );


  buf

  (
    g1564_n_spl_001,
    g1564_n_spl_00
  );


  buf

  (
    g1564_n_spl_01,
    g1564_n_spl_0
  );


  buf

  (
    g1564_n_spl_010,
    g1564_n_spl_01
  );


  buf

  (
    g1564_n_spl_011,
    g1564_n_spl_01
  );


  buf

  (
    g1564_n_spl_1,
    g1564_n_spl_
  );


  buf

  (
    g1564_n_spl_10,
    g1564_n_spl_1
  );


  buf

  (
    g1564_n_spl_11,
    g1564_n_spl_1
  );


  buf

  (
    g1566_n_spl_,
    g1566_n
  );


  buf

  (
    g1566_n_spl_0,
    g1566_n_spl_
  );


  buf

  (
    g1566_n_spl_00,
    g1566_n_spl_0
  );


  buf

  (
    g1566_n_spl_000,
    g1566_n_spl_00
  );


  buf

  (
    g1566_n_spl_001,
    g1566_n_spl_00
  );


  buf

  (
    g1566_n_spl_01,
    g1566_n_spl_0
  );


  buf

  (
    g1566_n_spl_010,
    g1566_n_spl_01
  );


  buf

  (
    g1566_n_spl_011,
    g1566_n_spl_01
  );


  buf

  (
    g1566_n_spl_1,
    g1566_n_spl_
  );


  buf

  (
    g1566_n_spl_10,
    g1566_n_spl_1
  );


  buf

  (
    g1566_n_spl_11,
    g1566_n_spl_1
  );


  buf

  (
    g1567_p_spl_,
    g1567_p
  );


  buf

  (
    g1567_p_spl_0,
    g1567_p_spl_
  );


  buf

  (
    g1567_p_spl_00,
    g1567_p_spl_0
  );


  buf

  (
    g1567_p_spl_000,
    g1567_p_spl_00
  );


  buf

  (
    g1567_p_spl_001,
    g1567_p_spl_00
  );


  buf

  (
    g1567_p_spl_01,
    g1567_p_spl_0
  );


  buf

  (
    g1567_p_spl_010,
    g1567_p_spl_01
  );


  buf

  (
    g1567_p_spl_011,
    g1567_p_spl_01
  );


  buf

  (
    g1567_p_spl_1,
    g1567_p_spl_
  );


  buf

  (
    g1567_p_spl_10,
    g1567_p_spl_1
  );


  buf

  (
    g1567_p_spl_11,
    g1567_p_spl_1
  );


  buf

  (
    g1568_n_spl_,
    g1568_n
  );


  buf

  (
    g1568_n_spl_0,
    g1568_n_spl_
  );


  buf

  (
    g1568_n_spl_00,
    g1568_n_spl_0
  );


  buf

  (
    g1568_n_spl_000,
    g1568_n_spl_00
  );


  buf

  (
    g1568_n_spl_001,
    g1568_n_spl_00
  );


  buf

  (
    g1568_n_spl_01,
    g1568_n_spl_0
  );


  buf

  (
    g1568_n_spl_010,
    g1568_n_spl_01
  );


  buf

  (
    g1568_n_spl_011,
    g1568_n_spl_01
  );


  buf

  (
    g1568_n_spl_1,
    g1568_n_spl_
  );


  buf

  (
    g1568_n_spl_10,
    g1568_n_spl_1
  );


  buf

  (
    g1568_n_spl_11,
    g1568_n_spl_1
  );


  buf

  (
    g1569_n_spl_,
    g1569_n
  );


  buf

  (
    g1569_n_spl_0,
    g1569_n_spl_
  );


  buf

  (
    g1569_n_spl_00,
    g1569_n_spl_0
  );


  buf

  (
    g1569_n_spl_000,
    g1569_n_spl_00
  );


  buf

  (
    g1569_n_spl_001,
    g1569_n_spl_00
  );


  buf

  (
    g1569_n_spl_01,
    g1569_n_spl_0
  );


  buf

  (
    g1569_n_spl_010,
    g1569_n_spl_01
  );


  buf

  (
    g1569_n_spl_011,
    g1569_n_spl_01
  );


  buf

  (
    g1569_n_spl_1,
    g1569_n_spl_
  );


  buf

  (
    g1569_n_spl_10,
    g1569_n_spl_1
  );


  buf

  (
    g1569_n_spl_11,
    g1569_n_spl_1
  );


  buf

  (
    g1577_p_spl_,
    g1577_p
  );


  buf

  (
    g1577_p_spl_0,
    g1577_p_spl_
  );


  buf

  (
    G9_p_spl_,
    G9_p
  );


  buf

  (
    G9_p_spl_0,
    G9_p_spl_
  );


  buf

  (
    G9_p_spl_1,
    G9_p_spl_
  );


  buf

  (
    G13_p_spl_,
    G13_p
  );


  buf

  (
    G13_p_spl_0,
    G13_p_spl_
  );


  buf

  (
    G13_p_spl_1,
    G13_p_spl_
  );


  buf

  (
    g1592_n_spl_,
    g1592_n
  );


  buf

  (
    g1678_p_spl_,
    g1678_p
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    g1692_p_spl_,
    g1692_p
  );


  buf

  (
    g1706_n_spl_,
    g1706_n
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    g1719_n_spl_,
    g1719_n
  );


endmodule
