
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  G42,
  G43,
  G44,
  G45,
  G46,
  G47,
  G48,
  G49,
  G50,
  G51,
  G52,
  G53,
  G54,
  G55,
  G56,
  G57,
  G58,
  G59,
  G60,
  G61,
  G62,
  G63,
  G64,
  G65,
  G66,
  G67,
  G68,
  G69,
  G70,
  G71,
  G72,
  G73,
  G74,
  G75,
  G76,
  G77,
  G78,
  G79,
  G80,
  G81,
  G82,
  G83,
  G84,
  G85,
  G86,
  G87,
  G88,
  G89,
  G90,
  G91,
  G92,
  G93,
  G94,
  G95,
  G96,
  G97,
  G98,
  G99,
  G100,
  G101,
  G102,
  G103,
  G104,
  G105,
  G106,
  G107,
  G108,
  G109,
  G110,
  G111,
  G112,
  G113,
  G114,
  G115,
  G116,
  G117,
  G118,
  G119,
  G120,
  G121,
  G122,
  G123,
  G124,
  G125,
  G126,
  G127,
  G128,
  G129,
  G130,
  G131,
  G132,
  G133,
  G134,
  G135,
  G136,
  G137,
  G138,
  G139,
  G140,
  G141,
  G142,
  G143,
  G144,
  G145,
  G146,
  G147,
  G148,
  G149,
  G150,
  G151,
  G152,
  G153,
  G154,
  G155,
  G156,
  G157,
  n1416_lo,
  n1419_lo,
  n1422_lo,
  n1425_lo,
  n1428_lo,
  n1431_lo,
  n1434_lo,
  n1437_lo,
  n1440_lo,
  n1443_lo,
  n1446_lo,
  n1449_lo,
  n1452_lo,
  n1455_lo,
  n1458_lo,
  n1464_lo,
  n1467_lo,
  n1470_lo,
  n1476_lo,
  n1479_lo,
  n1482_lo,
  n1488_lo,
  n1491_lo,
  n1494_lo,
  n1497_lo,
  n1500_lo,
  n1512_lo,
  n1515_lo,
  n1518_lo,
  n1521_lo,
  n1524_lo,
  n1527_lo,
  n1530_lo,
  n1533_lo,
  n1536_lo,
  n1539_lo,
  n1542_lo,
  n1545_lo,
  n1548_lo,
  n1551_lo,
  n1554_lo,
  n1560_lo,
  n1563_lo,
  n1566_lo,
  n1572_lo,
  n1575_lo,
  n1578_lo,
  n1584_lo,
  n1587_lo,
  n1590_lo,
  n1596_lo,
  n1599_lo,
  n1602_lo,
  n1608_lo,
  n1611_lo,
  n1614_lo,
  n1620_lo,
  n1623_lo,
  n1626_lo,
  n1632_lo,
  n1635_lo,
  n1638_lo,
  n1644_lo,
  n1647_lo,
  n1650_lo,
  n1656_lo,
  n1659_lo,
  n1662_lo,
  n1668_lo,
  n1671_lo,
  n1674_lo,
  n1677_lo,
  n1680_lo,
  n1683_lo,
  n1686_lo,
  n1692_lo,
  n1695_lo,
  n1698_lo,
  n1704_lo,
  n1707_lo,
  n1710_lo,
  n1716_lo,
  n1719_lo,
  n1722_lo,
  n1728_lo,
  n1731_lo,
  n1734_lo,
  n1740_lo,
  n1743_lo,
  n1746_lo,
  n1749_lo,
  n1752_lo,
  n1755_lo,
  n1758_lo,
  n1761_lo,
  n1764_lo,
  n1776_lo,
  n1779_lo,
  n1788_lo,
  n1791_lo,
  n1794_lo,
  n1797_lo,
  n1800_lo,
  n1812_lo,
  n1824_lo,
  n1836_lo,
  n1848_lo,
  n1860_lo,
  n1872_lo,
  n1884_lo,
  n1896_lo,
  n1899_lo,
  n1908_lo,
  n1911_lo,
  n1920_lo,
  n1923_lo,
  n1926_lo,
  n1929_lo,
  n1932_lo,
  n1944_lo,
  n1956_lo,
  n1968_lo,
  n1980_lo,
  n1992_lo,
  n2004_lo,
  n2016_lo,
  n2019_lo,
  n2028_lo,
  n2031_lo,
  n2040_lo,
  n2043_lo,
  n2046_lo,
  n2049_lo,
  n2052_lo,
  n2064_lo,
  n2076_lo,
  n2088_lo,
  n2100_lo,
  n2112_lo,
  n2124_lo,
  n2136_lo,
  n2148_lo,
  n2151_lo,
  n2160_lo,
  n2163_lo,
  n2172_lo,
  n2175_lo,
  n2178_lo,
  n2181_lo,
  n2184_lo,
  n2196_lo,
  n2208_lo,
  n2220_lo,
  n2232_lo,
  n2244_lo,
  n2256_lo,
  n2268_lo,
  n2280_lo,
  n2283_lo,
  n2292_lo,
  n2295_lo,
  n2298_lo,
  n2301_lo,
  n2304_lo,
  n2316_lo,
  n2319_lo,
  n2322_lo,
  n2325_lo,
  n2328_lo,
  n2331_lo,
  n2340_lo,
  n2343_lo,
  n2376_lo,
  n2379_lo,
  n2388_lo,
  n2400_lo,
  n2412_lo,
  n2415_lo,
  n2424_lo,
  n2436_lo,
  n2439_lo,
  n2442_lo,
  n2445_lo,
  n2448_lo,
  n2451_lo,
  n2460_lo,
  n2463_lo,
  n2496_lo,
  n2499_lo,
  n2508_lo,
  n2520_lo,
  n2532_lo,
  n2535_lo,
  n2544_lo,
  n2556_lo,
  n2559_lo,
  n2562_lo,
  n2565_lo,
  n2568_lo,
  n2571_lo,
  n2580_lo,
  n2583_lo,
  n2616_lo,
  n2619_lo,
  n2628_lo,
  n2640_lo,
  n2652_lo,
  n2655_lo,
  n2664_lo,
  n2676_lo,
  n2679_lo,
  n2682_lo,
  n2685_lo,
  n2688_lo,
  n2691_lo,
  n2700_lo,
  n2703_lo,
  n2736_lo,
  n2739_lo,
  n2748_lo,
  n2760_lo,
  n2772_lo,
  n2775_lo,
  n2784_lo,
  n2787_lo,
  n2790_lo,
  n2793_lo,
  n2796_lo,
  n2799_lo,
  n2802_lo,
  n2805_lo,
  n2808_lo,
  n2820_lo,
  n2823_lo,
  n2826_lo,
  n2832_lo,
  n2835_lo,
  n2838_lo,
  n2841_lo,
  n2844_lo,
  n2856_lo,
  n2859_lo,
  n2862_lo,
  n2865_lo,
  n2868_lo,
  n2871_lo,
  n2874_lo,
  n2877_lo,
  n2880_lo,
  n2883_lo,
  n2886_lo,
  n2889_lo,
  n2892_lo,
  n2895_lo,
  n2898_lo,
  n2901_lo,
  n2904_lo,
  n2907_lo,
  n2916_lo,
  n2928_lo,
  n2940_lo,
  n2952_lo,
  n2955_lo,
  n2964_lo,
  n2976_lo,
  n2988_lo,
  n2991_lo,
  n3000_lo,
  n3003_lo,
  n3012_lo,
  n3015_lo,
  n3024_lo,
  n3027_lo,
  n3036_lo,
  n3039_lo,
  n3048_lo,
  n3051_lo,
  n3054_lo,
  n3057_lo,
  n3060_lo,
  n3072_lo,
  n3081_lo,
  n3084_lo,
  n3087_lo,
  n3093_lo,
  n3096_lo,
  n3105_lo,
  n3108_lo,
  n3117_lo,
  n3120_lo,
  n3123_lo,
  n3126_lo,
  n3129_lo,
  n3132_lo,
  n3135_lo,
  n3138_lo,
  n3141_lo,
  n3168_lo,
  n3171_lo,
  n3174_lo,
  n3177_lo,
  n3180_lo,
  n3183_lo,
  n3192_lo,
  n3195_lo,
  n3204_lo,
  n3207_lo,
  n3216_lo,
  n3219_lo,
  n3228_lo,
  n3231_lo,
  n3240_lo,
  n3243_lo,
  n3252_lo,
  n3255_lo,
  n3258_lo,
  n3264_lo,
  n3267_lo,
  n3270_lo,
  n3276_lo,
  n3279_lo,
  n3282_lo,
  n3288_lo,
  n3291_lo,
  n3294_lo,
  n4537_o2,
  n4538_o2,
  n4710_o2,
  n4711_o2,
  n1211_inv,
  n1214_inv,
  n1217_inv,
  n1220_inv,
  n4927_o2,
  n4928_o2,
  n1229_inv,
  n1232_inv,
  n1235_inv,
  n5178_o2,
  n5179_o2,
  n5477_o2,
  n5478_o2,
  n5479_o2,
  n5222_o2,
  n5223_o2,
  n5553_o2,
  n5554_o2,
  G491_o2,
  n2922_lo_buf_o2,
  n2946_lo_buf_o2,
  n2970_lo_buf_o2,
  n2982_lo_buf_o2,
  n3066_lo_buf_o2,
  n3078_lo_buf_o2,
  n3102_lo_buf_o2,
  n3114_lo_buf_o2,
  G1321_o2,
  G1033_o2,
  G1030_o2,
  G1072_o2,
  n1304_inv,
  n1307_inv,
  n2958_lo_buf_o2,
  n2994_lo_buf_o2,
  n3006_lo_buf_o2,
  n3030_lo_buf_o2,
  n3042_lo_buf_o2,
  n3090_lo_buf_o2,
  n1328_inv,
  n1331_inv,
  n1334_inv,
  n1337_inv,
  n1340_inv,
  n1343_inv,
  n1346_inv,
  n1349_inv,
  G1036_o2,
  G1062_o2,
  G1067_o2,
  G1014_o2,
  n1364_inv,
  n1367_inv,
  n3018_lo_buf_o2,
  G766_o2,
  n1376_inv,
  n1379_inv,
  n1382_inv,
  n1385_inv,
  n1388_inv,
  n1391_inv,
  G1017_o2,
  G1008_o2,
  n1400_inv,
  n1403_inv,
  n2910_lo_buf_o2,
  n1409_inv,
  G2138_o2,
  G2147_o2,
  n1418_inv,
  G1137_o2,
  G1329_o2,
  G374_o2,
  G386_o2,
  G663_o2,
  G674_o2,
  G578_o2,
  G575_o2,
  G2505_o2,
  n1448_inv,
  G987_o2,
  G984_o2,
  G1862_o2,
  G1859_o2,
  G1260_o2,
  G1865_o2,
  G2073_o2,
  G1402_o2,
  G2048_o2,
  G2276_o2,
  n1481_inv,
  G2141_o2,
  G2008_o2,
  G2011_o2,
  G2150_o2,
  G2026_o2,
  G2029_o2,
  G2023_o2,
  G2041_o2,
  G2017_o2,
  G2020_o2,
  G2035_o2,
  G2038_o2,
  G2228_o2,
  G2231_o2,
  G2234_o2,
  G2237_o2,
  G1904_o2,
  G1907_o2,
  G1928_o2,
  G1931_o2,
  G1893_o2,
  G1896_o2,
  G1899_o2,
  G1937_o2,
  G1940_o2,
  G1943_o2,
  G1336_o2,
  G1996_o2,
  G1999_o2,
  G2002_o2,
  G2005_o2,
  G2014_o2,
  G2032_o2,
  G1076_o2,
  G1002_o2,
  G998_o2,
  G1890_o2,
  G1934_o2,
  G1044_o2,
  G1039_o2,
  n1770_lo_buf_o2,
  G342_o2,
  G354_o2,
  G1193_o2,
  n3234_lo_buf_o2,
  n3246_lo_buf_o2,
  G783_o2,
  G786_o2,
  G792_o2,
  G795_o2,
  G815_o2,
  G818_o2,
  G824_o2,
  G827_o2,
  G789_o2,
  G798_o2,
  G801_o2,
  G807_o2,
  G812_o2,
  G821_o2,
  G804_o2,
  G780_o2,
  G1231_o2,
  G1572_o2,
  G1377_o2,
  G1253_o2,
  G1359_o2,
  G1258_o2,
  G1367_o2,
  G1358_o2,
  G1366_o2,
  G2057_o2,
  G2117_o2,
  G2118_o2,
  G1254_o2,
  G1259_o2,
  G2058_o2,
  G405_o2,
  G417_o2,
  G1269_o2,
  G1275_o2,
  G1287_o2,
  G1266_o2,
  G1272_o2,
  G1278_o2,
  G1281_o2,
  G1284_o2,
  G1290_o2,
  G1293_o2,
  G1299_o2,
  G1305_o2,
  G1296_o2,
  G1302_o2,
  G1308_o2,
  G1311_o2,
  G811_o2,
  G810_o2,
  G1728_o2,
  G2512_o2,
  G1114_o2,
  G1113_o2,
  G1992_o2,
  G1991_o2,
  G1426_o2,
  G1966_o2,
  G2211_o2,
  G1509_o2,
  G2153_o2,
  G2329_o2,
  G1540_o2,
  G2167_o2,
  G2191_o2,
  G1234_o2,
  G1132_o2,
  G1129_o2,
  G2088_o2,
  G2106_o2,
  G1314_o2,
  G636_o2,
  G647_o2,
  n3186_lo_buf_o2,
  n3198_lo_buf_o2,
  n3210_lo_buf_o2,
  n3222_lo_buf_o2,
  G1225_o2,
  G1342_o2,
  G1222_o2,
  G1228_o2,
  G1348_o2,
  G1345_o2,
  G1351_o2,
  G2242_o2,
  G2260_o2,
  G1374_o2,
  G1537_o2,
  G301_o2,
  G313_o2,
  G2365_o2,
  G2255_o2,
  G2253_o2,
  G2395_o2,
  G2272_o2,
  G2270_o2,
  G2245_o2,
  G2262_o2,
  G2249_o2,
  G2247_o2,
  G2266_o2,
  G2264_o2,
  G2403_o2,
  G2401_o2,
  G2410_o2,
  G2408_o2,
  G2306_o2,
  G2305_o2,
  G2314_o2,
  G2313_o2,
  G2303_o2,
  G2302_o2,
  G2301_o2,
  G2311_o2,
  G2310_o2,
  G2309_o2,
  G2404_o2,
  G2411_o2,
  G2420_o2,
  G2419_o2,
  G2433_o2,
  G2432_o2,
  G402_o2,
  G403_o2,
  G1053_o2,
  G1049_o2,
  n2003_inv,
  G1364_o2,
  G1079_o2,
  G1478_o2,
  G707_o2,
  G718_o2,
  G2417_o2,
  G2414_o2,
  G2431_o2,
  G2428_o2,
  G1653_o2,
  G2213_o2,
  G2221_o2,
  G2250_o2,
  G2267_o2,
  G1365_o2,
  G1368_o2,
  G1371_o2,
  G2218_o2,
  G2225_o2,
  n1503_lo_buf_o2,
  n1863_lo_buf_o2,
  n1887_lo_buf_o2,
  n1983_lo_buf_o2,
  n2007_lo_buf_o2,
  n2115_lo_buf_o2,
  n2139_lo_buf_o2,
  n2247_lo_buf_o2,
  n2271_lo_buf_o2,
  n2919_lo_buf_o2,
  n2943_lo_buf_o2,
  n2967_lo_buf_o2,
  n2979_lo_buf_o2,
  n3063_lo_buf_o2,
  n3075_lo_buf_o2,
  n3099_lo_buf_o2,
  n3111_lo_buf_o2,
  G878_o2,
  G875_o2,
  G661_o2,
  G660_o2,
  G879_o2,
  G876_o2,
  G1320_o2,
  G941_o2,
  G732_o2,
  G942_o2,
  G1493_o2,
  G1498_o2,
  G877_o2,
  G874_o2,
  n1806_lo_buf_o2,
  n1878_lo_buf_o2,
  n1938_lo_buf_o2,
  n1998_lo_buf_o2,
  n2058_lo_buf_o2,
  n2130_lo_buf_o2,
  n2190_lo_buf_o2,
  n2262_lo_buf_o2,
  n2310_lo_buf_o2,
  n2406_lo_buf_o2,
  n2430_lo_buf_o2,
  n2526_lo_buf_o2,
  n2550_lo_buf_o2,
  n2646_lo_buf_o2,
  n2670_lo_buf_o2,
  n2766_lo_buf_o2,
  G603_o2,
  G614_o2,
  G1026_o2,
  G1021_o2,
  G940_o2,
  G1636_o2,
  G1684_o2,
  n2352_lo_buf_o2,
  n2364_lo_buf_o2,
  n2472_lo_buf_o2,
  n2484_lo_buf_o2,
  n2592_lo_buf_o2,
  n2604_lo_buf_o2,
  n2712_lo_buf_o2,
  n2724_lo_buf_o2,
  n3150_lo_buf_o2,
  n3162_lo_buf_o2,
  G2531,
  G2532,
  G2533,
  G2534,
  G2535,
  G2536,
  G2537,
  G2538,
  G2539,
  G2540,
  G2541,
  G2542,
  G2543,
  G2544,
  G2545,
  G2546,
  G2547,
  G2548,
  G2549,
  G2550,
  G2551,
  G2552,
  G2553,
  G2554,
  G2555,
  G2556,
  G2557,
  G2558,
  G2559,
  G2560,
  G2561,
  G2562,
  G2563,
  G2564,
  G2565,
  G2566,
  G2567,
  G2568,
  G2569,
  G2570,
  G2571,
  G2572,
  G2573,
  G2574,
  G2575,
  G2576,
  G2577,
  G2578,
  G2579,
  G2580,
  G2581,
  G2582,
  G2583,
  G2584,
  G2585,
  G2586,
  G2587,
  G2588,
  G2589,
  G2590,
  G2591,
  G2592,
  G2593,
  G2594,
  n1416_li,
  n1419_li,
  n1422_li,
  n1425_li,
  n1428_li,
  n1431_li,
  n1434_li,
  n1437_li,
  n1440_li,
  n1443_li,
  n1446_li,
  n1449_li,
  n1452_li,
  n1455_li,
  n1458_li,
  n1464_li,
  n1467_li,
  n1470_li,
  n1476_li,
  n1479_li,
  n1482_li,
  n1488_li,
  n1491_li,
  n1494_li,
  n1497_li,
  n1500_li,
  n1512_li,
  n1515_li,
  n1518_li,
  n1521_li,
  n1524_li,
  n1527_li,
  n1530_li,
  n1533_li,
  n1536_li,
  n1539_li,
  n1542_li,
  n1545_li,
  n1548_li,
  n1551_li,
  n1554_li,
  n1560_li,
  n1563_li,
  n1566_li,
  n1572_li,
  n1575_li,
  n1578_li,
  n1584_li,
  n1587_li,
  n1590_li,
  n1596_li,
  n1599_li,
  n1602_li,
  n1608_li,
  n1611_li,
  n1614_li,
  n1620_li,
  n1623_li,
  n1626_li,
  n1632_li,
  n1635_li,
  n1638_li,
  n1644_li,
  n1647_li,
  n1650_li,
  n1656_li,
  n1659_li,
  n1662_li,
  n1668_li,
  n1671_li,
  n1674_li,
  n1677_li,
  n1680_li,
  n1683_li,
  n1686_li,
  n1692_li,
  n1695_li,
  n1698_li,
  n1704_li,
  n1707_li,
  n1710_li,
  n1716_li,
  n1719_li,
  n1722_li,
  n1728_li,
  n1731_li,
  n1734_li,
  n1740_li,
  n1743_li,
  n1746_li,
  n1749_li,
  n1752_li,
  n1755_li,
  n1758_li,
  n1761_li,
  n1764_li,
  n1776_li,
  n1779_li,
  n1788_li,
  n1791_li,
  n1794_li,
  n1797_li,
  n1800_li,
  n1812_li,
  n1824_li,
  n1836_li,
  n1848_li,
  n1860_li,
  n1872_li,
  n1884_li,
  n1896_li,
  n1899_li,
  n1908_li,
  n1911_li,
  n1920_li,
  n1923_li,
  n1926_li,
  n1929_li,
  n1932_li,
  n1944_li,
  n1956_li,
  n1968_li,
  n1980_li,
  n1992_li,
  n2004_li,
  n2016_li,
  n2019_li,
  n2028_li,
  n2031_li,
  n2040_li,
  n2043_li,
  n2046_li,
  n2049_li,
  n2052_li,
  n2064_li,
  n2076_li,
  n2088_li,
  n2100_li,
  n2112_li,
  n2124_li,
  n2136_li,
  n2148_li,
  n2151_li,
  n2160_li,
  n2163_li,
  n2172_li,
  n2175_li,
  n2178_li,
  n2181_li,
  n2184_li,
  n2196_li,
  n2208_li,
  n2220_li,
  n2232_li,
  n2244_li,
  n2256_li,
  n2268_li,
  n2280_li,
  n2283_li,
  n2292_li,
  n2295_li,
  n2298_li,
  n2301_li,
  n2304_li,
  n2316_li,
  n2319_li,
  n2322_li,
  n2325_li,
  n2328_li,
  n2331_li,
  n2340_li,
  n2343_li,
  n2376_li,
  n2379_li,
  n2388_li,
  n2400_li,
  n2412_li,
  n2415_li,
  n2424_li,
  n2436_li,
  n2439_li,
  n2442_li,
  n2445_li,
  n2448_li,
  n2451_li,
  n2460_li,
  n2463_li,
  n2496_li,
  n2499_li,
  n2508_li,
  n2520_li,
  n2532_li,
  n2535_li,
  n2544_li,
  n2556_li,
  n2559_li,
  n2562_li,
  n2565_li,
  n2568_li,
  n2571_li,
  n2580_li,
  n2583_li,
  n2616_li,
  n2619_li,
  n2628_li,
  n2640_li,
  n2652_li,
  n2655_li,
  n2664_li,
  n2676_li,
  n2679_li,
  n2682_li,
  n2685_li,
  n2688_li,
  n2691_li,
  n2700_li,
  n2703_li,
  n2736_li,
  n2739_li,
  n2748_li,
  n2760_li,
  n2772_li,
  n2775_li,
  n2784_li,
  n2787_li,
  n2790_li,
  n2793_li,
  n2796_li,
  n2799_li,
  n2802_li,
  n2805_li,
  n2808_li,
  n2820_li,
  n2823_li,
  n2826_li,
  n2832_li,
  n2835_li,
  n2838_li,
  n2841_li,
  n2844_li,
  n2856_li,
  n2859_li,
  n2862_li,
  n2865_li,
  n2868_li,
  n2871_li,
  n2874_li,
  n2877_li,
  n2880_li,
  n2883_li,
  n2886_li,
  n2889_li,
  n2892_li,
  n2895_li,
  n2898_li,
  n2901_li,
  n2904_li,
  n2907_li,
  n2916_li,
  n2928_li,
  n2940_li,
  n2952_li,
  n2955_li,
  n2964_li,
  n2976_li,
  n2988_li,
  n2991_li,
  n3000_li,
  n3003_li,
  n3012_li,
  n3015_li,
  n3024_li,
  n3027_li,
  n3036_li,
  n3039_li,
  n3048_li,
  n3051_li,
  n3054_li,
  n3057_li,
  n3060_li,
  n3072_li,
  n3081_li,
  n3084_li,
  n3087_li,
  n3093_li,
  n3096_li,
  n3105_li,
  n3108_li,
  n3117_li,
  n3120_li,
  n3123_li,
  n3126_li,
  n3129_li,
  n3132_li,
  n3135_li,
  n3138_li,
  n3141_li,
  n3168_li,
  n3171_li,
  n3174_li,
  n3177_li,
  n3180_li,
  n3183_li,
  n3192_li,
  n3195_li,
  n3204_li,
  n3207_li,
  n3216_li,
  n3219_li,
  n3228_li,
  n3231_li,
  n3240_li,
  n3243_li,
  n3252_li,
  n3255_li,
  n3258_li,
  n3264_li,
  n3267_li,
  n3270_li,
  n3276_li,
  n3279_li,
  n3282_li,
  n3288_li,
  n3291_li,
  n3294_li,
  n4537_i2,
  n4538_i2,
  n4710_i2,
  n4711_i2,
  n4803_i2,
  n4804_i2,
  n4843_i2,
  n4844_i2,
  n4927_i2,
  n4928_i2,
  n4945_i2,
  n4946_i2,
  n5009_i2,
  n5178_i2,
  n5179_i2,
  n5477_i2,
  n5478_i2,
  n5479_i2,
  n5222_i2,
  n5223_i2,
  n5553_i2,
  n5554_i2,
  G491_i2,
  n2922_lo_buf_i2,
  n2946_lo_buf_i2,
  n2970_lo_buf_i2,
  n2982_lo_buf_i2,
  n3066_lo_buf_i2,
  n3078_lo_buf_i2,
  n3102_lo_buf_i2,
  n3114_lo_buf_i2,
  G1321_i2,
  G1033_i2,
  G1030_i2,
  G1072_i2,
  G1159_i2,
  G1152_i2,
  n2958_lo_buf_i2,
  n2994_lo_buf_i2,
  n3006_lo_buf_i2,
  n3030_lo_buf_i2,
  n3042_lo_buf_i2,
  n3090_lo_buf_i2,
  G370_i2,
  G447_i2,
  G455_i2,
  G459_i2,
  G497_i2,
  G503_i2,
  G511_i2,
  G515_i2,
  G1036_i2,
  G1062_i2,
  G1067_i2,
  G1014_i2,
  G1171_i2,
  G1166_i2,
  n3018_lo_buf_i2,
  G766_i2,
  G451_i2,
  G463_i2,
  G467_i2,
  G475_i2,
  G479_i2,
  G507_i2,
  G1017_i2,
  G1008_i2,
  G1176_i2,
  G1144_i2,
  n2910_lo_buf_i2,
  G471_i2,
  G2138_i2,
  G2147_i2,
  G1148_i2,
  G1137_i2,
  G1329_i2,
  G374_i2,
  G386_i2,
  G663_i2,
  G674_i2,
  G578_i2,
  G575_i2,
  G2505_i2,
  G2508_i2,
  G987_i2,
  G984_i2,
  G1862_i2,
  G1859_i2,
  G1260_i2,
  G1865_i2,
  G2073_i2,
  G1402_i2,
  G2048_i2,
  G2276_i2,
  G366_i2,
  G2141_i2,
  G2008_i2,
  G2011_i2,
  G2150_i2,
  G2026_i2,
  G2029_i2,
  G2023_i2,
  G2041_i2,
  G2017_i2,
  G2020_i2,
  G2035_i2,
  G2038_i2,
  G2228_i2,
  G2231_i2,
  G2234_i2,
  G2237_i2,
  G1904_i2,
  G1907_i2,
  G1928_i2,
  G1931_i2,
  G1893_i2,
  G1896_i2,
  G1899_i2,
  G1937_i2,
  G1940_i2,
  G1943_i2,
  G1336_i2,
  G1996_i2,
  G1999_i2,
  G2002_i2,
  G2005_i2,
  G2014_i2,
  G2032_i2,
  G1076_i2,
  G1002_i2,
  G998_i2,
  G1890_i2,
  G1934_i2,
  G1044_i2,
  G1039_i2,
  n1770_lo_buf_i2,
  G342_i2,
  G354_i2,
  G1193_i2,
  n3234_lo_buf_i2,
  n3246_lo_buf_i2,
  G783_i2,
  G786_i2,
  G792_i2,
  G795_i2,
  G815_i2,
  G818_i2,
  G824_i2,
  G827_i2,
  G789_i2,
  G798_i2,
  G801_i2,
  G807_i2,
  G812_i2,
  G821_i2,
  G804_i2,
  G780_i2,
  G1231_i2,
  G1572_i2,
  G1377_i2,
  G1253_i2,
  G1359_i2,
  G1258_i2,
  G1367_i2,
  G1358_i2,
  G1366_i2,
  G2057_i2,
  G2117_i2,
  G2118_i2,
  G1254_i2,
  G1259_i2,
  G2058_i2,
  G405_i2,
  G417_i2,
  G1269_i2,
  G1275_i2,
  G1287_i2,
  G1266_i2,
  G1272_i2,
  G1278_i2,
  G1281_i2,
  G1284_i2,
  G1290_i2,
  G1293_i2,
  G1299_i2,
  G1305_i2,
  G1296_i2,
  G1302_i2,
  G1308_i2,
  G1311_i2,
  G811_i2,
  G810_i2,
  G1728_i2,
  G2512_i2,
  G1114_i2,
  G1113_i2,
  G1992_i2,
  G1991_i2,
  G1426_i2,
  G1966_i2,
  G2211_i2,
  G1509_i2,
  G2153_i2,
  G2329_i2,
  G1540_i2,
  G2167_i2,
  G2191_i2,
  G1234_i2,
  G1132_i2,
  G1129_i2,
  G2088_i2,
  G2106_i2,
  G1314_i2,
  G636_i2,
  G647_i2,
  n3186_lo_buf_i2,
  n3198_lo_buf_i2,
  n3210_lo_buf_i2,
  n3222_lo_buf_i2,
  G1225_i2,
  G1342_i2,
  G1222_i2,
  G1228_i2,
  G1348_i2,
  G1345_i2,
  G1351_i2,
  G2242_i2,
  G2260_i2,
  G1374_i2,
  G1537_i2,
  G301_i2,
  G313_i2,
  G2365_i2,
  G2255_i2,
  G2253_i2,
  G2395_i2,
  G2272_i2,
  G2270_i2,
  G2245_i2,
  G2262_i2,
  G2249_i2,
  G2247_i2,
  G2266_i2,
  G2264_i2,
  G2403_i2,
  G2401_i2,
  G2410_i2,
  G2408_i2,
  G2306_i2,
  G2305_i2,
  G2314_i2,
  G2313_i2,
  G2303_i2,
  G2302_i2,
  G2301_i2,
  G2311_i2,
  G2310_i2,
  G2309_i2,
  G2404_i2,
  G2411_i2,
  G2420_i2,
  G2419_i2,
  G2433_i2,
  G2432_i2,
  G402_i2,
  G403_i2,
  G1053_i2,
  G1049_i2,
  G1058_i2,
  G1364_i2,
  G1079_i2,
  G1478_i2,
  G707_i2,
  G718_i2,
  G2417_i2,
  G2414_i2,
  G2431_i2,
  G2428_i2,
  G1653_i2,
  G2213_i2,
  G2221_i2,
  G2250_i2,
  G2267_i2,
  G1365_i2,
  G1368_i2,
  G1371_i2,
  G2218_i2,
  G2225_i2,
  n1503_lo_buf_i2,
  n1863_lo_buf_i2,
  n1887_lo_buf_i2,
  n1983_lo_buf_i2,
  n2007_lo_buf_i2,
  n2115_lo_buf_i2,
  n2139_lo_buf_i2,
  n2247_lo_buf_i2,
  n2271_lo_buf_i2,
  n2919_lo_buf_i2,
  n2943_lo_buf_i2,
  n2967_lo_buf_i2,
  n2979_lo_buf_i2,
  n3063_lo_buf_i2,
  n3075_lo_buf_i2,
  n3099_lo_buf_i2,
  n3111_lo_buf_i2,
  G878_i2,
  G875_i2,
  G661_i2,
  G660_i2,
  G879_i2,
  G876_i2,
  G1320_i2,
  G941_i2,
  G732_i2,
  G942_i2,
  G1493_i2,
  G1498_i2,
  G877_i2,
  G874_i2,
  n1806_lo_buf_i2,
  n1878_lo_buf_i2,
  n1938_lo_buf_i2,
  n1998_lo_buf_i2,
  n2058_lo_buf_i2,
  n2130_lo_buf_i2,
  n2190_lo_buf_i2,
  n2262_lo_buf_i2,
  n2310_lo_buf_i2,
  n2406_lo_buf_i2,
  n2430_lo_buf_i2,
  n2526_lo_buf_i2,
  n2550_lo_buf_i2,
  n2646_lo_buf_i2,
  n2670_lo_buf_i2,
  n2766_lo_buf_i2,
  G603_i2,
  G614_i2,
  G1026_i2,
  G1021_i2,
  G940_i2,
  G1636_i2,
  G1684_i2,
  n2352_lo_buf_i2,
  n2364_lo_buf_i2,
  n2472_lo_buf_i2,
  n2484_lo_buf_i2,
  n2592_lo_buf_i2,
  n2604_lo_buf_i2,
  n2712_lo_buf_i2,
  n2724_lo_buf_i2,
  n3150_lo_buf_i2,
  n3162_lo_buf_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input G42;input G43;input G44;input G45;input G46;input G47;input G48;input G49;input G50;input G51;input G52;input G53;input G54;input G55;input G56;input G57;input G58;input G59;input G60;input G61;input G62;input G63;input G64;input G65;input G66;input G67;input G68;input G69;input G70;input G71;input G72;input G73;input G74;input G75;input G76;input G77;input G78;input G79;input G80;input G81;input G82;input G83;input G84;input G85;input G86;input G87;input G88;input G89;input G90;input G91;input G92;input G93;input G94;input G95;input G96;input G97;input G98;input G99;input G100;input G101;input G102;input G103;input G104;input G105;input G106;input G107;input G108;input G109;input G110;input G111;input G112;input G113;input G114;input G115;input G116;input G117;input G118;input G119;input G120;input G121;input G122;input G123;input G124;input G125;input G126;input G127;input G128;input G129;input G130;input G131;input G132;input G133;input G134;input G135;input G136;input G137;input G138;input G139;input G140;input G141;input G142;input G143;input G144;input G145;input G146;input G147;input G148;input G149;input G150;input G151;input G152;input G153;input G154;input G155;input G156;input G157;input n1416_lo;input n1419_lo;input n1422_lo;input n1425_lo;input n1428_lo;input n1431_lo;input n1434_lo;input n1437_lo;input n1440_lo;input n1443_lo;input n1446_lo;input n1449_lo;input n1452_lo;input n1455_lo;input n1458_lo;input n1464_lo;input n1467_lo;input n1470_lo;input n1476_lo;input n1479_lo;input n1482_lo;input n1488_lo;input n1491_lo;input n1494_lo;input n1497_lo;input n1500_lo;input n1512_lo;input n1515_lo;input n1518_lo;input n1521_lo;input n1524_lo;input n1527_lo;input n1530_lo;input n1533_lo;input n1536_lo;input n1539_lo;input n1542_lo;input n1545_lo;input n1548_lo;input n1551_lo;input n1554_lo;input n1560_lo;input n1563_lo;input n1566_lo;input n1572_lo;input n1575_lo;input n1578_lo;input n1584_lo;input n1587_lo;input n1590_lo;input n1596_lo;input n1599_lo;input n1602_lo;input n1608_lo;input n1611_lo;input n1614_lo;input n1620_lo;input n1623_lo;input n1626_lo;input n1632_lo;input n1635_lo;input n1638_lo;input n1644_lo;input n1647_lo;input n1650_lo;input n1656_lo;input n1659_lo;input n1662_lo;input n1668_lo;input n1671_lo;input n1674_lo;input n1677_lo;input n1680_lo;input n1683_lo;input n1686_lo;input n1692_lo;input n1695_lo;input n1698_lo;input n1704_lo;input n1707_lo;input n1710_lo;input n1716_lo;input n1719_lo;input n1722_lo;input n1728_lo;input n1731_lo;input n1734_lo;input n1740_lo;input n1743_lo;input n1746_lo;input n1749_lo;input n1752_lo;input n1755_lo;input n1758_lo;input n1761_lo;input n1764_lo;input n1776_lo;input n1779_lo;input n1788_lo;input n1791_lo;input n1794_lo;input n1797_lo;input n1800_lo;input n1812_lo;input n1824_lo;input n1836_lo;input n1848_lo;input n1860_lo;input n1872_lo;input n1884_lo;input n1896_lo;input n1899_lo;input n1908_lo;input n1911_lo;input n1920_lo;input n1923_lo;input n1926_lo;input n1929_lo;input n1932_lo;input n1944_lo;input n1956_lo;input n1968_lo;input n1980_lo;input n1992_lo;input n2004_lo;input n2016_lo;input n2019_lo;input n2028_lo;input n2031_lo;input n2040_lo;input n2043_lo;input n2046_lo;input n2049_lo;input n2052_lo;input n2064_lo;input n2076_lo;input n2088_lo;input n2100_lo;input n2112_lo;input n2124_lo;input n2136_lo;input n2148_lo;input n2151_lo;input n2160_lo;input n2163_lo;input n2172_lo;input n2175_lo;input n2178_lo;input n2181_lo;input n2184_lo;input n2196_lo;input n2208_lo;input n2220_lo;input n2232_lo;input n2244_lo;input n2256_lo;input n2268_lo;input n2280_lo;input n2283_lo;input n2292_lo;input n2295_lo;input n2298_lo;input n2301_lo;input n2304_lo;input n2316_lo;input n2319_lo;input n2322_lo;input n2325_lo;input n2328_lo;input n2331_lo;input n2340_lo;input n2343_lo;input n2376_lo;input n2379_lo;input n2388_lo;input n2400_lo;input n2412_lo;input n2415_lo;input n2424_lo;input n2436_lo;input n2439_lo;input n2442_lo;input n2445_lo;input n2448_lo;input n2451_lo;input n2460_lo;input n2463_lo;input n2496_lo;input n2499_lo;input n2508_lo;input n2520_lo;input n2532_lo;input n2535_lo;input n2544_lo;input n2556_lo;input n2559_lo;input n2562_lo;input n2565_lo;input n2568_lo;input n2571_lo;input n2580_lo;input n2583_lo;input n2616_lo;input n2619_lo;input n2628_lo;input n2640_lo;input n2652_lo;input n2655_lo;input n2664_lo;input n2676_lo;input n2679_lo;input n2682_lo;input n2685_lo;input n2688_lo;input n2691_lo;input n2700_lo;input n2703_lo;input n2736_lo;input n2739_lo;input n2748_lo;input n2760_lo;input n2772_lo;input n2775_lo;input n2784_lo;input n2787_lo;input n2790_lo;input n2793_lo;input n2796_lo;input n2799_lo;input n2802_lo;input n2805_lo;input n2808_lo;input n2820_lo;input n2823_lo;input n2826_lo;input n2832_lo;input n2835_lo;input n2838_lo;input n2841_lo;input n2844_lo;input n2856_lo;input n2859_lo;input n2862_lo;input n2865_lo;input n2868_lo;input n2871_lo;input n2874_lo;input n2877_lo;input n2880_lo;input n2883_lo;input n2886_lo;input n2889_lo;input n2892_lo;input n2895_lo;input n2898_lo;input n2901_lo;input n2904_lo;input n2907_lo;input n2916_lo;input n2928_lo;input n2940_lo;input n2952_lo;input n2955_lo;input n2964_lo;input n2976_lo;input n2988_lo;input n2991_lo;input n3000_lo;input n3003_lo;input n3012_lo;input n3015_lo;input n3024_lo;input n3027_lo;input n3036_lo;input n3039_lo;input n3048_lo;input n3051_lo;input n3054_lo;input n3057_lo;input n3060_lo;input n3072_lo;input n3081_lo;input n3084_lo;input n3087_lo;input n3093_lo;input n3096_lo;input n3105_lo;input n3108_lo;input n3117_lo;input n3120_lo;input n3123_lo;input n3126_lo;input n3129_lo;input n3132_lo;input n3135_lo;input n3138_lo;input n3141_lo;input n3168_lo;input n3171_lo;input n3174_lo;input n3177_lo;input n3180_lo;input n3183_lo;input n3192_lo;input n3195_lo;input n3204_lo;input n3207_lo;input n3216_lo;input n3219_lo;input n3228_lo;input n3231_lo;input n3240_lo;input n3243_lo;input n3252_lo;input n3255_lo;input n3258_lo;input n3264_lo;input n3267_lo;input n3270_lo;input n3276_lo;input n3279_lo;input n3282_lo;input n3288_lo;input n3291_lo;input n3294_lo;input n4537_o2;input n4538_o2;input n4710_o2;input n4711_o2;input n1211_inv;input n1214_inv;input n1217_inv;input n1220_inv;input n4927_o2;input n4928_o2;input n1229_inv;input n1232_inv;input n1235_inv;input n5178_o2;input n5179_o2;input n5477_o2;input n5478_o2;input n5479_o2;input n5222_o2;input n5223_o2;input n5553_o2;input n5554_o2;input G491_o2;input n2922_lo_buf_o2;input n2946_lo_buf_o2;input n2970_lo_buf_o2;input n2982_lo_buf_o2;input n3066_lo_buf_o2;input n3078_lo_buf_o2;input n3102_lo_buf_o2;input n3114_lo_buf_o2;input G1321_o2;input G1033_o2;input G1030_o2;input G1072_o2;input n1304_inv;input n1307_inv;input n2958_lo_buf_o2;input n2994_lo_buf_o2;input n3006_lo_buf_o2;input n3030_lo_buf_o2;input n3042_lo_buf_o2;input n3090_lo_buf_o2;input n1328_inv;input n1331_inv;input n1334_inv;input n1337_inv;input n1340_inv;input n1343_inv;input n1346_inv;input n1349_inv;input G1036_o2;input G1062_o2;input G1067_o2;input G1014_o2;input n1364_inv;input n1367_inv;input n3018_lo_buf_o2;input G766_o2;input n1376_inv;input n1379_inv;input n1382_inv;input n1385_inv;input n1388_inv;input n1391_inv;input G1017_o2;input G1008_o2;input n1400_inv;input n1403_inv;input n2910_lo_buf_o2;input n1409_inv;input G2138_o2;input G2147_o2;input n1418_inv;input G1137_o2;input G1329_o2;input G374_o2;input G386_o2;input G663_o2;input G674_o2;input G578_o2;input G575_o2;input G2505_o2;input n1448_inv;input G987_o2;input G984_o2;input G1862_o2;input G1859_o2;input G1260_o2;input G1865_o2;input G2073_o2;input G1402_o2;input G2048_o2;input G2276_o2;input n1481_inv;input G2141_o2;input G2008_o2;input G2011_o2;input G2150_o2;input G2026_o2;input G2029_o2;input G2023_o2;input G2041_o2;input G2017_o2;input G2020_o2;input G2035_o2;input G2038_o2;input G2228_o2;input G2231_o2;input G2234_o2;input G2237_o2;input G1904_o2;input G1907_o2;input G1928_o2;input G1931_o2;input G1893_o2;input G1896_o2;input G1899_o2;input G1937_o2;input G1940_o2;input G1943_o2;input G1336_o2;input G1996_o2;input G1999_o2;input G2002_o2;input G2005_o2;input G2014_o2;input G2032_o2;input G1076_o2;input G1002_o2;input G998_o2;input G1890_o2;input G1934_o2;input G1044_o2;input G1039_o2;input n1770_lo_buf_o2;input G342_o2;input G354_o2;input G1193_o2;input n3234_lo_buf_o2;input n3246_lo_buf_o2;input G783_o2;input G786_o2;input G792_o2;input G795_o2;input G815_o2;input G818_o2;input G824_o2;input G827_o2;input G789_o2;input G798_o2;input G801_o2;input G807_o2;input G812_o2;input G821_o2;input G804_o2;input G780_o2;input G1231_o2;input G1572_o2;input G1377_o2;input G1253_o2;input G1359_o2;input G1258_o2;input G1367_o2;input G1358_o2;input G1366_o2;input G2057_o2;input G2117_o2;input G2118_o2;input G1254_o2;input G1259_o2;input G2058_o2;input G405_o2;input G417_o2;input G1269_o2;input G1275_o2;input G1287_o2;input G1266_o2;input G1272_o2;input G1278_o2;input G1281_o2;input G1284_o2;input G1290_o2;input G1293_o2;input G1299_o2;input G1305_o2;input G1296_o2;input G1302_o2;input G1308_o2;input G1311_o2;input G811_o2;input G810_o2;input G1728_o2;input G2512_o2;input G1114_o2;input G1113_o2;input G1992_o2;input G1991_o2;input G1426_o2;input G1966_o2;input G2211_o2;input G1509_o2;input G2153_o2;input G2329_o2;input G1540_o2;input G2167_o2;input G2191_o2;input G1234_o2;input G1132_o2;input G1129_o2;input G2088_o2;input G2106_o2;input G1314_o2;input G636_o2;input G647_o2;input n3186_lo_buf_o2;input n3198_lo_buf_o2;input n3210_lo_buf_o2;input n3222_lo_buf_o2;input G1225_o2;input G1342_o2;input G1222_o2;input G1228_o2;input G1348_o2;input G1345_o2;input G1351_o2;input G2242_o2;input G2260_o2;input G1374_o2;input G1537_o2;input G301_o2;input G313_o2;input G2365_o2;input G2255_o2;input G2253_o2;input G2395_o2;input G2272_o2;input G2270_o2;input G2245_o2;input G2262_o2;input G2249_o2;input G2247_o2;input G2266_o2;input G2264_o2;input G2403_o2;input G2401_o2;input G2410_o2;input G2408_o2;input G2306_o2;input G2305_o2;input G2314_o2;input G2313_o2;input G2303_o2;input G2302_o2;input G2301_o2;input G2311_o2;input G2310_o2;input G2309_o2;input G2404_o2;input G2411_o2;input G2420_o2;input G2419_o2;input G2433_o2;input G2432_o2;input G402_o2;input G403_o2;input G1053_o2;input G1049_o2;input n2003_inv;input G1364_o2;input G1079_o2;input G1478_o2;input G707_o2;input G718_o2;input G2417_o2;input G2414_o2;input G2431_o2;input G2428_o2;input G1653_o2;input G2213_o2;input G2221_o2;input G2250_o2;input G2267_o2;input G1365_o2;input G1368_o2;input G1371_o2;input G2218_o2;input G2225_o2;input n1503_lo_buf_o2;input n1863_lo_buf_o2;input n1887_lo_buf_o2;input n1983_lo_buf_o2;input n2007_lo_buf_o2;input n2115_lo_buf_o2;input n2139_lo_buf_o2;input n2247_lo_buf_o2;input n2271_lo_buf_o2;input n2919_lo_buf_o2;input n2943_lo_buf_o2;input n2967_lo_buf_o2;input n2979_lo_buf_o2;input n3063_lo_buf_o2;input n3075_lo_buf_o2;input n3099_lo_buf_o2;input n3111_lo_buf_o2;input G878_o2;input G875_o2;input G661_o2;input G660_o2;input G879_o2;input G876_o2;input G1320_o2;input G941_o2;input G732_o2;input G942_o2;input G1493_o2;input G1498_o2;input G877_o2;input G874_o2;input n1806_lo_buf_o2;input n1878_lo_buf_o2;input n1938_lo_buf_o2;input n1998_lo_buf_o2;input n2058_lo_buf_o2;input n2130_lo_buf_o2;input n2190_lo_buf_o2;input n2262_lo_buf_o2;input n2310_lo_buf_o2;input n2406_lo_buf_o2;input n2430_lo_buf_o2;input n2526_lo_buf_o2;input n2550_lo_buf_o2;input n2646_lo_buf_o2;input n2670_lo_buf_o2;input n2766_lo_buf_o2;input G603_o2;input G614_o2;input G1026_o2;input G1021_o2;input G940_o2;input G1636_o2;input G1684_o2;input n2352_lo_buf_o2;input n2364_lo_buf_o2;input n2472_lo_buf_o2;input n2484_lo_buf_o2;input n2592_lo_buf_o2;input n2604_lo_buf_o2;input n2712_lo_buf_o2;input n2724_lo_buf_o2;input n3150_lo_buf_o2;input n3162_lo_buf_o2;
  output G2531;output G2532;output G2533;output G2534;output G2535;output G2536;output G2537;output G2538;output G2539;output G2540;output G2541;output G2542;output G2543;output G2544;output G2545;output G2546;output G2547;output G2548;output G2549;output G2550;output G2551;output G2552;output G2553;output G2554;output G2555;output G2556;output G2557;output G2558;output G2559;output G2560;output G2561;output G2562;output G2563;output G2564;output G2565;output G2566;output G2567;output G2568;output G2569;output G2570;output G2571;output G2572;output G2573;output G2574;output G2575;output G2576;output G2577;output G2578;output G2579;output G2580;output G2581;output G2582;output G2583;output G2584;output G2585;output G2586;output G2587;output G2588;output G2589;output G2590;output G2591;output G2592;output G2593;output G2594;output n1416_li;output n1419_li;output n1422_li;output n1425_li;output n1428_li;output n1431_li;output n1434_li;output n1437_li;output n1440_li;output n1443_li;output n1446_li;output n1449_li;output n1452_li;output n1455_li;output n1458_li;output n1464_li;output n1467_li;output n1470_li;output n1476_li;output n1479_li;output n1482_li;output n1488_li;output n1491_li;output n1494_li;output n1497_li;output n1500_li;output n1512_li;output n1515_li;output n1518_li;output n1521_li;output n1524_li;output n1527_li;output n1530_li;output n1533_li;output n1536_li;output n1539_li;output n1542_li;output n1545_li;output n1548_li;output n1551_li;output n1554_li;output n1560_li;output n1563_li;output n1566_li;output n1572_li;output n1575_li;output n1578_li;output n1584_li;output n1587_li;output n1590_li;output n1596_li;output n1599_li;output n1602_li;output n1608_li;output n1611_li;output n1614_li;output n1620_li;output n1623_li;output n1626_li;output n1632_li;output n1635_li;output n1638_li;output n1644_li;output n1647_li;output n1650_li;output n1656_li;output n1659_li;output n1662_li;output n1668_li;output n1671_li;output n1674_li;output n1677_li;output n1680_li;output n1683_li;output n1686_li;output n1692_li;output n1695_li;output n1698_li;output n1704_li;output n1707_li;output n1710_li;output n1716_li;output n1719_li;output n1722_li;output n1728_li;output n1731_li;output n1734_li;output n1740_li;output n1743_li;output n1746_li;output n1749_li;output n1752_li;output n1755_li;output n1758_li;output n1761_li;output n1764_li;output n1776_li;output n1779_li;output n1788_li;output n1791_li;output n1794_li;output n1797_li;output n1800_li;output n1812_li;output n1824_li;output n1836_li;output n1848_li;output n1860_li;output n1872_li;output n1884_li;output n1896_li;output n1899_li;output n1908_li;output n1911_li;output n1920_li;output n1923_li;output n1926_li;output n1929_li;output n1932_li;output n1944_li;output n1956_li;output n1968_li;output n1980_li;output n1992_li;output n2004_li;output n2016_li;output n2019_li;output n2028_li;output n2031_li;output n2040_li;output n2043_li;output n2046_li;output n2049_li;output n2052_li;output n2064_li;output n2076_li;output n2088_li;output n2100_li;output n2112_li;output n2124_li;output n2136_li;output n2148_li;output n2151_li;output n2160_li;output n2163_li;output n2172_li;output n2175_li;output n2178_li;output n2181_li;output n2184_li;output n2196_li;output n2208_li;output n2220_li;output n2232_li;output n2244_li;output n2256_li;output n2268_li;output n2280_li;output n2283_li;output n2292_li;output n2295_li;output n2298_li;output n2301_li;output n2304_li;output n2316_li;output n2319_li;output n2322_li;output n2325_li;output n2328_li;output n2331_li;output n2340_li;output n2343_li;output n2376_li;output n2379_li;output n2388_li;output n2400_li;output n2412_li;output n2415_li;output n2424_li;output n2436_li;output n2439_li;output n2442_li;output n2445_li;output n2448_li;output n2451_li;output n2460_li;output n2463_li;output n2496_li;output n2499_li;output n2508_li;output n2520_li;output n2532_li;output n2535_li;output n2544_li;output n2556_li;output n2559_li;output n2562_li;output n2565_li;output n2568_li;output n2571_li;output n2580_li;output n2583_li;output n2616_li;output n2619_li;output n2628_li;output n2640_li;output n2652_li;output n2655_li;output n2664_li;output n2676_li;output n2679_li;output n2682_li;output n2685_li;output n2688_li;output n2691_li;output n2700_li;output n2703_li;output n2736_li;output n2739_li;output n2748_li;output n2760_li;output n2772_li;output n2775_li;output n2784_li;output n2787_li;output n2790_li;output n2793_li;output n2796_li;output n2799_li;output n2802_li;output n2805_li;output n2808_li;output n2820_li;output n2823_li;output n2826_li;output n2832_li;output n2835_li;output n2838_li;output n2841_li;output n2844_li;output n2856_li;output n2859_li;output n2862_li;output n2865_li;output n2868_li;output n2871_li;output n2874_li;output n2877_li;output n2880_li;output n2883_li;output n2886_li;output n2889_li;output n2892_li;output n2895_li;output n2898_li;output n2901_li;output n2904_li;output n2907_li;output n2916_li;output n2928_li;output n2940_li;output n2952_li;output n2955_li;output n2964_li;output n2976_li;output n2988_li;output n2991_li;output n3000_li;output n3003_li;output n3012_li;output n3015_li;output n3024_li;output n3027_li;output n3036_li;output n3039_li;output n3048_li;output n3051_li;output n3054_li;output n3057_li;output n3060_li;output n3072_li;output n3081_li;output n3084_li;output n3087_li;output n3093_li;output n3096_li;output n3105_li;output n3108_li;output n3117_li;output n3120_li;output n3123_li;output n3126_li;output n3129_li;output n3132_li;output n3135_li;output n3138_li;output n3141_li;output n3168_li;output n3171_li;output n3174_li;output n3177_li;output n3180_li;output n3183_li;output n3192_li;output n3195_li;output n3204_li;output n3207_li;output n3216_li;output n3219_li;output n3228_li;output n3231_li;output n3240_li;output n3243_li;output n3252_li;output n3255_li;output n3258_li;output n3264_li;output n3267_li;output n3270_li;output n3276_li;output n3279_li;output n3282_li;output n3288_li;output n3291_li;output n3294_li;output n4537_i2;output n4538_i2;output n4710_i2;output n4711_i2;output n4803_i2;output n4804_i2;output n4843_i2;output n4844_i2;output n4927_i2;output n4928_i2;output n4945_i2;output n4946_i2;output n5009_i2;output n5178_i2;output n5179_i2;output n5477_i2;output n5478_i2;output n5479_i2;output n5222_i2;output n5223_i2;output n5553_i2;output n5554_i2;output G491_i2;output n2922_lo_buf_i2;output n2946_lo_buf_i2;output n2970_lo_buf_i2;output n2982_lo_buf_i2;output n3066_lo_buf_i2;output n3078_lo_buf_i2;output n3102_lo_buf_i2;output n3114_lo_buf_i2;output G1321_i2;output G1033_i2;output G1030_i2;output G1072_i2;output G1159_i2;output G1152_i2;output n2958_lo_buf_i2;output n2994_lo_buf_i2;output n3006_lo_buf_i2;output n3030_lo_buf_i2;output n3042_lo_buf_i2;output n3090_lo_buf_i2;output G370_i2;output G447_i2;output G455_i2;output G459_i2;output G497_i2;output G503_i2;output G511_i2;output G515_i2;output G1036_i2;output G1062_i2;output G1067_i2;output G1014_i2;output G1171_i2;output G1166_i2;output n3018_lo_buf_i2;output G766_i2;output G451_i2;output G463_i2;output G467_i2;output G475_i2;output G479_i2;output G507_i2;output G1017_i2;output G1008_i2;output G1176_i2;output G1144_i2;output n2910_lo_buf_i2;output G471_i2;output G2138_i2;output G2147_i2;output G1148_i2;output G1137_i2;output G1329_i2;output G374_i2;output G386_i2;output G663_i2;output G674_i2;output G578_i2;output G575_i2;output G2505_i2;output G2508_i2;output G987_i2;output G984_i2;output G1862_i2;output G1859_i2;output G1260_i2;output G1865_i2;output G2073_i2;output G1402_i2;output G2048_i2;output G2276_i2;output G366_i2;output G2141_i2;output G2008_i2;output G2011_i2;output G2150_i2;output G2026_i2;output G2029_i2;output G2023_i2;output G2041_i2;output G2017_i2;output G2020_i2;output G2035_i2;output G2038_i2;output G2228_i2;output G2231_i2;output G2234_i2;output G2237_i2;output G1904_i2;output G1907_i2;output G1928_i2;output G1931_i2;output G1893_i2;output G1896_i2;output G1899_i2;output G1937_i2;output G1940_i2;output G1943_i2;output G1336_i2;output G1996_i2;output G1999_i2;output G2002_i2;output G2005_i2;output G2014_i2;output G2032_i2;output G1076_i2;output G1002_i2;output G998_i2;output G1890_i2;output G1934_i2;output G1044_i2;output G1039_i2;output n1770_lo_buf_i2;output G342_i2;output G354_i2;output G1193_i2;output n3234_lo_buf_i2;output n3246_lo_buf_i2;output G783_i2;output G786_i2;output G792_i2;output G795_i2;output G815_i2;output G818_i2;output G824_i2;output G827_i2;output G789_i2;output G798_i2;output G801_i2;output G807_i2;output G812_i2;output G821_i2;output G804_i2;output G780_i2;output G1231_i2;output G1572_i2;output G1377_i2;output G1253_i2;output G1359_i2;output G1258_i2;output G1367_i2;output G1358_i2;output G1366_i2;output G2057_i2;output G2117_i2;output G2118_i2;output G1254_i2;output G1259_i2;output G2058_i2;output G405_i2;output G417_i2;output G1269_i2;output G1275_i2;output G1287_i2;output G1266_i2;output G1272_i2;output G1278_i2;output G1281_i2;output G1284_i2;output G1290_i2;output G1293_i2;output G1299_i2;output G1305_i2;output G1296_i2;output G1302_i2;output G1308_i2;output G1311_i2;output G811_i2;output G810_i2;output G1728_i2;output G2512_i2;output G1114_i2;output G1113_i2;output G1992_i2;output G1991_i2;output G1426_i2;output G1966_i2;output G2211_i2;output G1509_i2;output G2153_i2;output G2329_i2;output G1540_i2;output G2167_i2;output G2191_i2;output G1234_i2;output G1132_i2;output G1129_i2;output G2088_i2;output G2106_i2;output G1314_i2;output G636_i2;output G647_i2;output n3186_lo_buf_i2;output n3198_lo_buf_i2;output n3210_lo_buf_i2;output n3222_lo_buf_i2;output G1225_i2;output G1342_i2;output G1222_i2;output G1228_i2;output G1348_i2;output G1345_i2;output G1351_i2;output G2242_i2;output G2260_i2;output G1374_i2;output G1537_i2;output G301_i2;output G313_i2;output G2365_i2;output G2255_i2;output G2253_i2;output G2395_i2;output G2272_i2;output G2270_i2;output G2245_i2;output G2262_i2;output G2249_i2;output G2247_i2;output G2266_i2;output G2264_i2;output G2403_i2;output G2401_i2;output G2410_i2;output G2408_i2;output G2306_i2;output G2305_i2;output G2314_i2;output G2313_i2;output G2303_i2;output G2302_i2;output G2301_i2;output G2311_i2;output G2310_i2;output G2309_i2;output G2404_i2;output G2411_i2;output G2420_i2;output G2419_i2;output G2433_i2;output G2432_i2;output G402_i2;output G403_i2;output G1053_i2;output G1049_i2;output G1058_i2;output G1364_i2;output G1079_i2;output G1478_i2;output G707_i2;output G718_i2;output G2417_i2;output G2414_i2;output G2431_i2;output G2428_i2;output G1653_i2;output G2213_i2;output G2221_i2;output G2250_i2;output G2267_i2;output G1365_i2;output G1368_i2;output G1371_i2;output G2218_i2;output G2225_i2;output n1503_lo_buf_i2;output n1863_lo_buf_i2;output n1887_lo_buf_i2;output n1983_lo_buf_i2;output n2007_lo_buf_i2;output n2115_lo_buf_i2;output n2139_lo_buf_i2;output n2247_lo_buf_i2;output n2271_lo_buf_i2;output n2919_lo_buf_i2;output n2943_lo_buf_i2;output n2967_lo_buf_i2;output n2979_lo_buf_i2;output n3063_lo_buf_i2;output n3075_lo_buf_i2;output n3099_lo_buf_i2;output n3111_lo_buf_i2;output G878_i2;output G875_i2;output G661_i2;output G660_i2;output G879_i2;output G876_i2;output G1320_i2;output G941_i2;output G732_i2;output G942_i2;output G1493_i2;output G1498_i2;output G877_i2;output G874_i2;output n1806_lo_buf_i2;output n1878_lo_buf_i2;output n1938_lo_buf_i2;output n1998_lo_buf_i2;output n2058_lo_buf_i2;output n2130_lo_buf_i2;output n2190_lo_buf_i2;output n2262_lo_buf_i2;output n2310_lo_buf_i2;output n2406_lo_buf_i2;output n2430_lo_buf_i2;output n2526_lo_buf_i2;output n2550_lo_buf_i2;output n2646_lo_buf_i2;output n2670_lo_buf_i2;output n2766_lo_buf_i2;output G603_i2;output G614_i2;output G1026_i2;output G1021_i2;output G940_i2;output G1636_i2;output G1684_i2;output n2352_lo_buf_i2;output n2364_lo_buf_i2;output n2472_lo_buf_i2;output n2484_lo_buf_i2;output n2592_lo_buf_i2;output n2604_lo_buf_i2;output n2712_lo_buf_i2;output n2724_lo_buf_i2;output n3150_lo_buf_i2;output n3162_lo_buf_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire G51_p;
  wire G51_n;
  wire G52_p;
  wire G52_n;
  wire G53_p;
  wire G53_n;
  wire G54_p;
  wire G54_n;
  wire G55_p;
  wire G55_n;
  wire G56_p;
  wire G56_n;
  wire G57_p;
  wire G57_n;
  wire G58_p;
  wire G58_n;
  wire G59_p;
  wire G59_n;
  wire G60_p;
  wire G60_n;
  wire G61_p;
  wire G61_n;
  wire G62_p;
  wire G62_n;
  wire G63_p;
  wire G63_n;
  wire G64_p;
  wire G64_n;
  wire G65_p;
  wire G65_n;
  wire G66_p;
  wire G66_n;
  wire G67_p;
  wire G67_n;
  wire G68_p;
  wire G68_n;
  wire G69_p;
  wire G69_n;
  wire G70_p;
  wire G70_n;
  wire G71_p;
  wire G71_n;
  wire G72_p;
  wire G72_n;
  wire G73_p;
  wire G73_n;
  wire G74_p;
  wire G74_n;
  wire G75_p;
  wire G75_n;
  wire G76_p;
  wire G76_n;
  wire G77_p;
  wire G77_n;
  wire G78_p;
  wire G78_n;
  wire G79_p;
  wire G79_n;
  wire G80_p;
  wire G80_n;
  wire G81_p;
  wire G81_n;
  wire G82_p;
  wire G82_n;
  wire G83_p;
  wire G83_n;
  wire G84_p;
  wire G84_n;
  wire G85_p;
  wire G85_n;
  wire G86_p;
  wire G86_n;
  wire G87_p;
  wire G87_n;
  wire G88_p;
  wire G88_n;
  wire G89_p;
  wire G89_n;
  wire G90_p;
  wire G90_n;
  wire G91_p;
  wire G91_n;
  wire G92_p;
  wire G92_n;
  wire G93_p;
  wire G93_n;
  wire G94_p;
  wire G94_n;
  wire G95_p;
  wire G95_n;
  wire G96_p;
  wire G96_n;
  wire G97_p;
  wire G97_n;
  wire G98_p;
  wire G98_n;
  wire G99_p;
  wire G99_n;
  wire G100_p;
  wire G100_n;
  wire G101_p;
  wire G101_n;
  wire G102_p;
  wire G102_n;
  wire G103_p;
  wire G103_n;
  wire G104_p;
  wire G104_n;
  wire G105_p;
  wire G105_n;
  wire G106_p;
  wire G106_n;
  wire G107_p;
  wire G107_n;
  wire G108_p;
  wire G108_n;
  wire G109_p;
  wire G109_n;
  wire G110_p;
  wire G110_n;
  wire G111_p;
  wire G111_n;
  wire G112_p;
  wire G112_n;
  wire G113_p;
  wire G113_n;
  wire G114_p;
  wire G114_n;
  wire G115_p;
  wire G115_n;
  wire G116_p;
  wire G116_n;
  wire G117_p;
  wire G117_n;
  wire G118_p;
  wire G118_n;
  wire G119_p;
  wire G119_n;
  wire G120_p;
  wire G120_n;
  wire G121_p;
  wire G121_n;
  wire G122_p;
  wire G122_n;
  wire G123_p;
  wire G123_n;
  wire G124_p;
  wire G124_n;
  wire G125_p;
  wire G125_n;
  wire G126_p;
  wire G126_n;
  wire G127_p;
  wire G127_n;
  wire G128_p;
  wire G128_n;
  wire G129_p;
  wire G129_n;
  wire G130_p;
  wire G130_n;
  wire G131_p;
  wire G131_n;
  wire G132_p;
  wire G132_n;
  wire G133_p;
  wire G133_n;
  wire G134_p;
  wire G134_n;
  wire G135_p;
  wire G135_n;
  wire G136_p;
  wire G136_n;
  wire G137_p;
  wire G137_n;
  wire G138_p;
  wire G138_n;
  wire G139_p;
  wire G139_n;
  wire G140_p;
  wire G140_n;
  wire G141_p;
  wire G141_n;
  wire G142_p;
  wire G142_n;
  wire G143_p;
  wire G143_n;
  wire G144_p;
  wire G144_n;
  wire G145_p;
  wire G145_n;
  wire G146_p;
  wire G146_n;
  wire G147_p;
  wire G147_n;
  wire G148_p;
  wire G148_n;
  wire G149_p;
  wire G149_n;
  wire G150_p;
  wire G150_n;
  wire G151_p;
  wire G151_n;
  wire G152_p;
  wire G152_n;
  wire G153_p;
  wire G153_n;
  wire G154_p;
  wire G154_n;
  wire G155_p;
  wire G155_n;
  wire G156_p;
  wire G156_n;
  wire G157_p;
  wire G157_n;
  wire n1416_lo_p;
  wire n1416_lo_n;
  wire n1419_lo_p;
  wire n1419_lo_n;
  wire n1422_lo_p;
  wire n1422_lo_n;
  wire n1425_lo_p;
  wire n1425_lo_n;
  wire n1428_lo_p;
  wire n1428_lo_n;
  wire n1431_lo_p;
  wire n1431_lo_n;
  wire n1434_lo_p;
  wire n1434_lo_n;
  wire n1437_lo_p;
  wire n1437_lo_n;
  wire n1440_lo_p;
  wire n1440_lo_n;
  wire n1443_lo_p;
  wire n1443_lo_n;
  wire n1446_lo_p;
  wire n1446_lo_n;
  wire n1449_lo_p;
  wire n1449_lo_n;
  wire n1452_lo_p;
  wire n1452_lo_n;
  wire n1455_lo_p;
  wire n1455_lo_n;
  wire n1458_lo_p;
  wire n1458_lo_n;
  wire n1464_lo_p;
  wire n1464_lo_n;
  wire n1467_lo_p;
  wire n1467_lo_n;
  wire n1470_lo_p;
  wire n1470_lo_n;
  wire n1476_lo_p;
  wire n1476_lo_n;
  wire n1479_lo_p;
  wire n1479_lo_n;
  wire n1482_lo_p;
  wire n1482_lo_n;
  wire n1488_lo_p;
  wire n1488_lo_n;
  wire n1491_lo_p;
  wire n1491_lo_n;
  wire n1494_lo_p;
  wire n1494_lo_n;
  wire n1497_lo_p;
  wire n1497_lo_n;
  wire n1500_lo_p;
  wire n1500_lo_n;
  wire n1512_lo_p;
  wire n1512_lo_n;
  wire n1515_lo_p;
  wire n1515_lo_n;
  wire n1518_lo_p;
  wire n1518_lo_n;
  wire n1521_lo_p;
  wire n1521_lo_n;
  wire n1524_lo_p;
  wire n1524_lo_n;
  wire n1527_lo_p;
  wire n1527_lo_n;
  wire n1530_lo_p;
  wire n1530_lo_n;
  wire n1533_lo_p;
  wire n1533_lo_n;
  wire n1536_lo_p;
  wire n1536_lo_n;
  wire n1539_lo_p;
  wire n1539_lo_n;
  wire n1542_lo_p;
  wire n1542_lo_n;
  wire n1545_lo_p;
  wire n1545_lo_n;
  wire n1548_lo_p;
  wire n1548_lo_n;
  wire n1551_lo_p;
  wire n1551_lo_n;
  wire n1554_lo_p;
  wire n1554_lo_n;
  wire n1560_lo_p;
  wire n1560_lo_n;
  wire n1563_lo_p;
  wire n1563_lo_n;
  wire n1566_lo_p;
  wire n1566_lo_n;
  wire n1572_lo_p;
  wire n1572_lo_n;
  wire n1575_lo_p;
  wire n1575_lo_n;
  wire n1578_lo_p;
  wire n1578_lo_n;
  wire n1584_lo_p;
  wire n1584_lo_n;
  wire n1587_lo_p;
  wire n1587_lo_n;
  wire n1590_lo_p;
  wire n1590_lo_n;
  wire n1596_lo_p;
  wire n1596_lo_n;
  wire n1599_lo_p;
  wire n1599_lo_n;
  wire n1602_lo_p;
  wire n1602_lo_n;
  wire n1608_lo_p;
  wire n1608_lo_n;
  wire n1611_lo_p;
  wire n1611_lo_n;
  wire n1614_lo_p;
  wire n1614_lo_n;
  wire n1620_lo_p;
  wire n1620_lo_n;
  wire n1623_lo_p;
  wire n1623_lo_n;
  wire n1626_lo_p;
  wire n1626_lo_n;
  wire n1632_lo_p;
  wire n1632_lo_n;
  wire n1635_lo_p;
  wire n1635_lo_n;
  wire n1638_lo_p;
  wire n1638_lo_n;
  wire n1644_lo_p;
  wire n1644_lo_n;
  wire n1647_lo_p;
  wire n1647_lo_n;
  wire n1650_lo_p;
  wire n1650_lo_n;
  wire n1656_lo_p;
  wire n1656_lo_n;
  wire n1659_lo_p;
  wire n1659_lo_n;
  wire n1662_lo_p;
  wire n1662_lo_n;
  wire n1668_lo_p;
  wire n1668_lo_n;
  wire n1671_lo_p;
  wire n1671_lo_n;
  wire n1674_lo_p;
  wire n1674_lo_n;
  wire n1677_lo_p;
  wire n1677_lo_n;
  wire n1680_lo_p;
  wire n1680_lo_n;
  wire n1683_lo_p;
  wire n1683_lo_n;
  wire n1686_lo_p;
  wire n1686_lo_n;
  wire n1692_lo_p;
  wire n1692_lo_n;
  wire n1695_lo_p;
  wire n1695_lo_n;
  wire n1698_lo_p;
  wire n1698_lo_n;
  wire n1704_lo_p;
  wire n1704_lo_n;
  wire n1707_lo_p;
  wire n1707_lo_n;
  wire n1710_lo_p;
  wire n1710_lo_n;
  wire n1716_lo_p;
  wire n1716_lo_n;
  wire n1719_lo_p;
  wire n1719_lo_n;
  wire n1722_lo_p;
  wire n1722_lo_n;
  wire n1728_lo_p;
  wire n1728_lo_n;
  wire n1731_lo_p;
  wire n1731_lo_n;
  wire n1734_lo_p;
  wire n1734_lo_n;
  wire n1740_lo_p;
  wire n1740_lo_n;
  wire n1743_lo_p;
  wire n1743_lo_n;
  wire n1746_lo_p;
  wire n1746_lo_n;
  wire n1749_lo_p;
  wire n1749_lo_n;
  wire n1752_lo_p;
  wire n1752_lo_n;
  wire n1755_lo_p;
  wire n1755_lo_n;
  wire n1758_lo_p;
  wire n1758_lo_n;
  wire n1761_lo_p;
  wire n1761_lo_n;
  wire n1764_lo_p;
  wire n1764_lo_n;
  wire n1776_lo_p;
  wire n1776_lo_n;
  wire n1779_lo_p;
  wire n1779_lo_n;
  wire n1788_lo_p;
  wire n1788_lo_n;
  wire n1791_lo_p;
  wire n1791_lo_n;
  wire n1794_lo_p;
  wire n1794_lo_n;
  wire n1797_lo_p;
  wire n1797_lo_n;
  wire n1800_lo_p;
  wire n1800_lo_n;
  wire n1812_lo_p;
  wire n1812_lo_n;
  wire n1824_lo_p;
  wire n1824_lo_n;
  wire n1836_lo_p;
  wire n1836_lo_n;
  wire n1848_lo_p;
  wire n1848_lo_n;
  wire n1860_lo_p;
  wire n1860_lo_n;
  wire n1872_lo_p;
  wire n1872_lo_n;
  wire n1884_lo_p;
  wire n1884_lo_n;
  wire n1896_lo_p;
  wire n1896_lo_n;
  wire n1899_lo_p;
  wire n1899_lo_n;
  wire n1908_lo_p;
  wire n1908_lo_n;
  wire n1911_lo_p;
  wire n1911_lo_n;
  wire n1920_lo_p;
  wire n1920_lo_n;
  wire n1923_lo_p;
  wire n1923_lo_n;
  wire n1926_lo_p;
  wire n1926_lo_n;
  wire n1929_lo_p;
  wire n1929_lo_n;
  wire n1932_lo_p;
  wire n1932_lo_n;
  wire n1944_lo_p;
  wire n1944_lo_n;
  wire n1956_lo_p;
  wire n1956_lo_n;
  wire n1968_lo_p;
  wire n1968_lo_n;
  wire n1980_lo_p;
  wire n1980_lo_n;
  wire n1992_lo_p;
  wire n1992_lo_n;
  wire n2004_lo_p;
  wire n2004_lo_n;
  wire n2016_lo_p;
  wire n2016_lo_n;
  wire n2019_lo_p;
  wire n2019_lo_n;
  wire n2028_lo_p;
  wire n2028_lo_n;
  wire n2031_lo_p;
  wire n2031_lo_n;
  wire n2040_lo_p;
  wire n2040_lo_n;
  wire n2043_lo_p;
  wire n2043_lo_n;
  wire n2046_lo_p;
  wire n2046_lo_n;
  wire n2049_lo_p;
  wire n2049_lo_n;
  wire n2052_lo_p;
  wire n2052_lo_n;
  wire n2064_lo_p;
  wire n2064_lo_n;
  wire n2076_lo_p;
  wire n2076_lo_n;
  wire n2088_lo_p;
  wire n2088_lo_n;
  wire n2100_lo_p;
  wire n2100_lo_n;
  wire n2112_lo_p;
  wire n2112_lo_n;
  wire n2124_lo_p;
  wire n2124_lo_n;
  wire n2136_lo_p;
  wire n2136_lo_n;
  wire n2148_lo_p;
  wire n2148_lo_n;
  wire n2151_lo_p;
  wire n2151_lo_n;
  wire n2160_lo_p;
  wire n2160_lo_n;
  wire n2163_lo_p;
  wire n2163_lo_n;
  wire n2172_lo_p;
  wire n2172_lo_n;
  wire n2175_lo_p;
  wire n2175_lo_n;
  wire n2178_lo_p;
  wire n2178_lo_n;
  wire n2181_lo_p;
  wire n2181_lo_n;
  wire n2184_lo_p;
  wire n2184_lo_n;
  wire n2196_lo_p;
  wire n2196_lo_n;
  wire n2208_lo_p;
  wire n2208_lo_n;
  wire n2220_lo_p;
  wire n2220_lo_n;
  wire n2232_lo_p;
  wire n2232_lo_n;
  wire n2244_lo_p;
  wire n2244_lo_n;
  wire n2256_lo_p;
  wire n2256_lo_n;
  wire n2268_lo_p;
  wire n2268_lo_n;
  wire n2280_lo_p;
  wire n2280_lo_n;
  wire n2283_lo_p;
  wire n2283_lo_n;
  wire n2292_lo_p;
  wire n2292_lo_n;
  wire n2295_lo_p;
  wire n2295_lo_n;
  wire n2298_lo_p;
  wire n2298_lo_n;
  wire n2301_lo_p;
  wire n2301_lo_n;
  wire n2304_lo_p;
  wire n2304_lo_n;
  wire n2316_lo_p;
  wire n2316_lo_n;
  wire n2319_lo_p;
  wire n2319_lo_n;
  wire n2322_lo_p;
  wire n2322_lo_n;
  wire n2325_lo_p;
  wire n2325_lo_n;
  wire n2328_lo_p;
  wire n2328_lo_n;
  wire n2331_lo_p;
  wire n2331_lo_n;
  wire n2340_lo_p;
  wire n2340_lo_n;
  wire n2343_lo_p;
  wire n2343_lo_n;
  wire n2376_lo_p;
  wire n2376_lo_n;
  wire n2379_lo_p;
  wire n2379_lo_n;
  wire n2388_lo_p;
  wire n2388_lo_n;
  wire n2400_lo_p;
  wire n2400_lo_n;
  wire n2412_lo_p;
  wire n2412_lo_n;
  wire n2415_lo_p;
  wire n2415_lo_n;
  wire n2424_lo_p;
  wire n2424_lo_n;
  wire n2436_lo_p;
  wire n2436_lo_n;
  wire n2439_lo_p;
  wire n2439_lo_n;
  wire n2442_lo_p;
  wire n2442_lo_n;
  wire n2445_lo_p;
  wire n2445_lo_n;
  wire n2448_lo_p;
  wire n2448_lo_n;
  wire n2451_lo_p;
  wire n2451_lo_n;
  wire n2460_lo_p;
  wire n2460_lo_n;
  wire n2463_lo_p;
  wire n2463_lo_n;
  wire n2496_lo_p;
  wire n2496_lo_n;
  wire n2499_lo_p;
  wire n2499_lo_n;
  wire n2508_lo_p;
  wire n2508_lo_n;
  wire n2520_lo_p;
  wire n2520_lo_n;
  wire n2532_lo_p;
  wire n2532_lo_n;
  wire n2535_lo_p;
  wire n2535_lo_n;
  wire n2544_lo_p;
  wire n2544_lo_n;
  wire n2556_lo_p;
  wire n2556_lo_n;
  wire n2559_lo_p;
  wire n2559_lo_n;
  wire n2562_lo_p;
  wire n2562_lo_n;
  wire n2565_lo_p;
  wire n2565_lo_n;
  wire n2568_lo_p;
  wire n2568_lo_n;
  wire n2571_lo_p;
  wire n2571_lo_n;
  wire n2580_lo_p;
  wire n2580_lo_n;
  wire n2583_lo_p;
  wire n2583_lo_n;
  wire n2616_lo_p;
  wire n2616_lo_n;
  wire n2619_lo_p;
  wire n2619_lo_n;
  wire n2628_lo_p;
  wire n2628_lo_n;
  wire n2640_lo_p;
  wire n2640_lo_n;
  wire n2652_lo_p;
  wire n2652_lo_n;
  wire n2655_lo_p;
  wire n2655_lo_n;
  wire n2664_lo_p;
  wire n2664_lo_n;
  wire n2676_lo_p;
  wire n2676_lo_n;
  wire n2679_lo_p;
  wire n2679_lo_n;
  wire n2682_lo_p;
  wire n2682_lo_n;
  wire n2685_lo_p;
  wire n2685_lo_n;
  wire n2688_lo_p;
  wire n2688_lo_n;
  wire n2691_lo_p;
  wire n2691_lo_n;
  wire n2700_lo_p;
  wire n2700_lo_n;
  wire n2703_lo_p;
  wire n2703_lo_n;
  wire n2736_lo_p;
  wire n2736_lo_n;
  wire n2739_lo_p;
  wire n2739_lo_n;
  wire n2748_lo_p;
  wire n2748_lo_n;
  wire n2760_lo_p;
  wire n2760_lo_n;
  wire n2772_lo_p;
  wire n2772_lo_n;
  wire n2775_lo_p;
  wire n2775_lo_n;
  wire n2784_lo_p;
  wire n2784_lo_n;
  wire n2787_lo_p;
  wire n2787_lo_n;
  wire n2790_lo_p;
  wire n2790_lo_n;
  wire n2793_lo_p;
  wire n2793_lo_n;
  wire n2796_lo_p;
  wire n2796_lo_n;
  wire n2799_lo_p;
  wire n2799_lo_n;
  wire n2802_lo_p;
  wire n2802_lo_n;
  wire n2805_lo_p;
  wire n2805_lo_n;
  wire n2808_lo_p;
  wire n2808_lo_n;
  wire n2820_lo_p;
  wire n2820_lo_n;
  wire n2823_lo_p;
  wire n2823_lo_n;
  wire n2826_lo_p;
  wire n2826_lo_n;
  wire n2832_lo_p;
  wire n2832_lo_n;
  wire n2835_lo_p;
  wire n2835_lo_n;
  wire n2838_lo_p;
  wire n2838_lo_n;
  wire n2841_lo_p;
  wire n2841_lo_n;
  wire n2844_lo_p;
  wire n2844_lo_n;
  wire n2856_lo_p;
  wire n2856_lo_n;
  wire n2859_lo_p;
  wire n2859_lo_n;
  wire n2862_lo_p;
  wire n2862_lo_n;
  wire n2865_lo_p;
  wire n2865_lo_n;
  wire n2868_lo_p;
  wire n2868_lo_n;
  wire n2871_lo_p;
  wire n2871_lo_n;
  wire n2874_lo_p;
  wire n2874_lo_n;
  wire n2877_lo_p;
  wire n2877_lo_n;
  wire n2880_lo_p;
  wire n2880_lo_n;
  wire n2883_lo_p;
  wire n2883_lo_n;
  wire n2886_lo_p;
  wire n2886_lo_n;
  wire n2889_lo_p;
  wire n2889_lo_n;
  wire n2892_lo_p;
  wire n2892_lo_n;
  wire n2895_lo_p;
  wire n2895_lo_n;
  wire n2898_lo_p;
  wire n2898_lo_n;
  wire n2901_lo_p;
  wire n2901_lo_n;
  wire n2904_lo_p;
  wire n2904_lo_n;
  wire n2907_lo_p;
  wire n2907_lo_n;
  wire n2916_lo_p;
  wire n2916_lo_n;
  wire n2928_lo_p;
  wire n2928_lo_n;
  wire n2940_lo_p;
  wire n2940_lo_n;
  wire n2952_lo_p;
  wire n2952_lo_n;
  wire n2955_lo_p;
  wire n2955_lo_n;
  wire n2964_lo_p;
  wire n2964_lo_n;
  wire n2976_lo_p;
  wire n2976_lo_n;
  wire n2988_lo_p;
  wire n2988_lo_n;
  wire n2991_lo_p;
  wire n2991_lo_n;
  wire n3000_lo_p;
  wire n3000_lo_n;
  wire n3003_lo_p;
  wire n3003_lo_n;
  wire n3012_lo_p;
  wire n3012_lo_n;
  wire n3015_lo_p;
  wire n3015_lo_n;
  wire n3024_lo_p;
  wire n3024_lo_n;
  wire n3027_lo_p;
  wire n3027_lo_n;
  wire n3036_lo_p;
  wire n3036_lo_n;
  wire n3039_lo_p;
  wire n3039_lo_n;
  wire n3048_lo_p;
  wire n3048_lo_n;
  wire n3051_lo_p;
  wire n3051_lo_n;
  wire n3054_lo_p;
  wire n3054_lo_n;
  wire n3057_lo_p;
  wire n3057_lo_n;
  wire n3060_lo_p;
  wire n3060_lo_n;
  wire n3072_lo_p;
  wire n3072_lo_n;
  wire n3081_lo_p;
  wire n3081_lo_n;
  wire n3084_lo_p;
  wire n3084_lo_n;
  wire n3087_lo_p;
  wire n3087_lo_n;
  wire n3093_lo_p;
  wire n3093_lo_n;
  wire n3096_lo_p;
  wire n3096_lo_n;
  wire n3105_lo_p;
  wire n3105_lo_n;
  wire n3108_lo_p;
  wire n3108_lo_n;
  wire n3117_lo_p;
  wire n3117_lo_n;
  wire n3120_lo_p;
  wire n3120_lo_n;
  wire n3123_lo_p;
  wire n3123_lo_n;
  wire n3126_lo_p;
  wire n3126_lo_n;
  wire n3129_lo_p;
  wire n3129_lo_n;
  wire n3132_lo_p;
  wire n3132_lo_n;
  wire n3135_lo_p;
  wire n3135_lo_n;
  wire n3138_lo_p;
  wire n3138_lo_n;
  wire n3141_lo_p;
  wire n3141_lo_n;
  wire n3168_lo_p;
  wire n3168_lo_n;
  wire n3171_lo_p;
  wire n3171_lo_n;
  wire n3174_lo_p;
  wire n3174_lo_n;
  wire n3177_lo_p;
  wire n3177_lo_n;
  wire n3180_lo_p;
  wire n3180_lo_n;
  wire n3183_lo_p;
  wire n3183_lo_n;
  wire n3192_lo_p;
  wire n3192_lo_n;
  wire n3195_lo_p;
  wire n3195_lo_n;
  wire n3204_lo_p;
  wire n3204_lo_n;
  wire n3207_lo_p;
  wire n3207_lo_n;
  wire n3216_lo_p;
  wire n3216_lo_n;
  wire n3219_lo_p;
  wire n3219_lo_n;
  wire n3228_lo_p;
  wire n3228_lo_n;
  wire n3231_lo_p;
  wire n3231_lo_n;
  wire n3240_lo_p;
  wire n3240_lo_n;
  wire n3243_lo_p;
  wire n3243_lo_n;
  wire n3252_lo_p;
  wire n3252_lo_n;
  wire n3255_lo_p;
  wire n3255_lo_n;
  wire n3258_lo_p;
  wire n3258_lo_n;
  wire n3264_lo_p;
  wire n3264_lo_n;
  wire n3267_lo_p;
  wire n3267_lo_n;
  wire n3270_lo_p;
  wire n3270_lo_n;
  wire n3276_lo_p;
  wire n3276_lo_n;
  wire n3279_lo_p;
  wire n3279_lo_n;
  wire n3282_lo_p;
  wire n3282_lo_n;
  wire n3288_lo_p;
  wire n3288_lo_n;
  wire n3291_lo_p;
  wire n3291_lo_n;
  wire n3294_lo_p;
  wire n3294_lo_n;
  wire n4537_o2_p;
  wire n4537_o2_n;
  wire n4538_o2_p;
  wire n4538_o2_n;
  wire n4710_o2_p;
  wire n4710_o2_n;
  wire n4711_o2_p;
  wire n4711_o2_n;
  wire n1211_inv_p;
  wire n1211_inv_n;
  wire n1214_inv_p;
  wire n1214_inv_n;
  wire n1217_inv_p;
  wire n1217_inv_n;
  wire n1220_inv_p;
  wire n1220_inv_n;
  wire n4927_o2_p;
  wire n4927_o2_n;
  wire n4928_o2_p;
  wire n4928_o2_n;
  wire n1229_inv_p;
  wire n1229_inv_n;
  wire n1232_inv_p;
  wire n1232_inv_n;
  wire n1235_inv_p;
  wire n1235_inv_n;
  wire n5178_o2_p;
  wire n5178_o2_n;
  wire n5179_o2_p;
  wire n5179_o2_n;
  wire n5477_o2_p;
  wire n5477_o2_n;
  wire n5478_o2_p;
  wire n5478_o2_n;
  wire n5479_o2_p;
  wire n5479_o2_n;
  wire n5222_o2_p;
  wire n5222_o2_n;
  wire n5223_o2_p;
  wire n5223_o2_n;
  wire n5553_o2_p;
  wire n5553_o2_n;
  wire n5554_o2_p;
  wire n5554_o2_n;
  wire G491_o2_p;
  wire G491_o2_n;
  wire n2922_lo_buf_o2_p;
  wire n2922_lo_buf_o2_n;
  wire n2946_lo_buf_o2_p;
  wire n2946_lo_buf_o2_n;
  wire n2970_lo_buf_o2_p;
  wire n2970_lo_buf_o2_n;
  wire n2982_lo_buf_o2_p;
  wire n2982_lo_buf_o2_n;
  wire n3066_lo_buf_o2_p;
  wire n3066_lo_buf_o2_n;
  wire n3078_lo_buf_o2_p;
  wire n3078_lo_buf_o2_n;
  wire n3102_lo_buf_o2_p;
  wire n3102_lo_buf_o2_n;
  wire n3114_lo_buf_o2_p;
  wire n3114_lo_buf_o2_n;
  wire G1321_o2_p;
  wire G1321_o2_n;
  wire G1033_o2_p;
  wire G1033_o2_n;
  wire G1030_o2_p;
  wire G1030_o2_n;
  wire G1072_o2_p;
  wire G1072_o2_n;
  wire n1304_inv_p;
  wire n1304_inv_n;
  wire n1307_inv_p;
  wire n1307_inv_n;
  wire n2958_lo_buf_o2_p;
  wire n2958_lo_buf_o2_n;
  wire n2994_lo_buf_o2_p;
  wire n2994_lo_buf_o2_n;
  wire n3006_lo_buf_o2_p;
  wire n3006_lo_buf_o2_n;
  wire n3030_lo_buf_o2_p;
  wire n3030_lo_buf_o2_n;
  wire n3042_lo_buf_o2_p;
  wire n3042_lo_buf_o2_n;
  wire n3090_lo_buf_o2_p;
  wire n3090_lo_buf_o2_n;
  wire n1328_inv_p;
  wire n1328_inv_n;
  wire n1331_inv_p;
  wire n1331_inv_n;
  wire n1334_inv_p;
  wire n1334_inv_n;
  wire n1337_inv_p;
  wire n1337_inv_n;
  wire n1340_inv_p;
  wire n1340_inv_n;
  wire n1343_inv_p;
  wire n1343_inv_n;
  wire n1346_inv_p;
  wire n1346_inv_n;
  wire n1349_inv_p;
  wire n1349_inv_n;
  wire G1036_o2_p;
  wire G1036_o2_n;
  wire G1062_o2_p;
  wire G1062_o2_n;
  wire G1067_o2_p;
  wire G1067_o2_n;
  wire G1014_o2_p;
  wire G1014_o2_n;
  wire n1364_inv_p;
  wire n1364_inv_n;
  wire n1367_inv_p;
  wire n1367_inv_n;
  wire n3018_lo_buf_o2_p;
  wire n3018_lo_buf_o2_n;
  wire G766_o2_p;
  wire G766_o2_n;
  wire n1376_inv_p;
  wire n1376_inv_n;
  wire n1379_inv_p;
  wire n1379_inv_n;
  wire n1382_inv_p;
  wire n1382_inv_n;
  wire n1385_inv_p;
  wire n1385_inv_n;
  wire n1388_inv_p;
  wire n1388_inv_n;
  wire n1391_inv_p;
  wire n1391_inv_n;
  wire G1017_o2_p;
  wire G1017_o2_n;
  wire G1008_o2_p;
  wire G1008_o2_n;
  wire n1400_inv_p;
  wire n1400_inv_n;
  wire n1403_inv_p;
  wire n1403_inv_n;
  wire n2910_lo_buf_o2_p;
  wire n2910_lo_buf_o2_n;
  wire n1409_inv_p;
  wire n1409_inv_n;
  wire G2138_o2_p;
  wire G2138_o2_n;
  wire G2147_o2_p;
  wire G2147_o2_n;
  wire n1418_inv_p;
  wire n1418_inv_n;
  wire G1137_o2_p;
  wire G1137_o2_n;
  wire G1329_o2_p;
  wire G1329_o2_n;
  wire G374_o2_p;
  wire G374_o2_n;
  wire G386_o2_p;
  wire G386_o2_n;
  wire G663_o2_p;
  wire G663_o2_n;
  wire G674_o2_p;
  wire G674_o2_n;
  wire G578_o2_p;
  wire G578_o2_n;
  wire G575_o2_p;
  wire G575_o2_n;
  wire G2505_o2_p;
  wire G2505_o2_n;
  wire n1448_inv_p;
  wire n1448_inv_n;
  wire G987_o2_p;
  wire G987_o2_n;
  wire G984_o2_p;
  wire G984_o2_n;
  wire G1862_o2_p;
  wire G1862_o2_n;
  wire G1859_o2_p;
  wire G1859_o2_n;
  wire G1260_o2_p;
  wire G1260_o2_n;
  wire G1865_o2_p;
  wire G1865_o2_n;
  wire G2073_o2_p;
  wire G2073_o2_n;
  wire G1402_o2_p;
  wire G1402_o2_n;
  wire G2048_o2_p;
  wire G2048_o2_n;
  wire G2276_o2_p;
  wire G2276_o2_n;
  wire n1481_inv_p;
  wire n1481_inv_n;
  wire G2141_o2_p;
  wire G2141_o2_n;
  wire G2008_o2_p;
  wire G2008_o2_n;
  wire G2011_o2_p;
  wire G2011_o2_n;
  wire G2150_o2_p;
  wire G2150_o2_n;
  wire G2026_o2_p;
  wire G2026_o2_n;
  wire G2029_o2_p;
  wire G2029_o2_n;
  wire G2023_o2_p;
  wire G2023_o2_n;
  wire G2041_o2_p;
  wire G2041_o2_n;
  wire G2017_o2_p;
  wire G2017_o2_n;
  wire G2020_o2_p;
  wire G2020_o2_n;
  wire G2035_o2_p;
  wire G2035_o2_n;
  wire G2038_o2_p;
  wire G2038_o2_n;
  wire G2228_o2_p;
  wire G2228_o2_n;
  wire G2231_o2_p;
  wire G2231_o2_n;
  wire G2234_o2_p;
  wire G2234_o2_n;
  wire G2237_o2_p;
  wire G2237_o2_n;
  wire G1904_o2_p;
  wire G1904_o2_n;
  wire G1907_o2_p;
  wire G1907_o2_n;
  wire G1928_o2_p;
  wire G1928_o2_n;
  wire G1931_o2_p;
  wire G1931_o2_n;
  wire G1893_o2_p;
  wire G1893_o2_n;
  wire G1896_o2_p;
  wire G1896_o2_n;
  wire G1899_o2_p;
  wire G1899_o2_n;
  wire G1937_o2_p;
  wire G1937_o2_n;
  wire G1940_o2_p;
  wire G1940_o2_n;
  wire G1943_o2_p;
  wire G1943_o2_n;
  wire G1336_o2_p;
  wire G1336_o2_n;
  wire G1996_o2_p;
  wire G1996_o2_n;
  wire G1999_o2_p;
  wire G1999_o2_n;
  wire G2002_o2_p;
  wire G2002_o2_n;
  wire G2005_o2_p;
  wire G2005_o2_n;
  wire G2014_o2_p;
  wire G2014_o2_n;
  wire G2032_o2_p;
  wire G2032_o2_n;
  wire G1076_o2_p;
  wire G1076_o2_n;
  wire G1002_o2_p;
  wire G1002_o2_n;
  wire G998_o2_p;
  wire G998_o2_n;
  wire G1890_o2_p;
  wire G1890_o2_n;
  wire G1934_o2_p;
  wire G1934_o2_n;
  wire G1044_o2_p;
  wire G1044_o2_n;
  wire G1039_o2_p;
  wire G1039_o2_n;
  wire n1770_lo_buf_o2_p;
  wire n1770_lo_buf_o2_n;
  wire G342_o2_p;
  wire G342_o2_n;
  wire G354_o2_p;
  wire G354_o2_n;
  wire G1193_o2_p;
  wire G1193_o2_n;
  wire n3234_lo_buf_o2_p;
  wire n3234_lo_buf_o2_n;
  wire n3246_lo_buf_o2_p;
  wire n3246_lo_buf_o2_n;
  wire G783_o2_p;
  wire G783_o2_n;
  wire G786_o2_p;
  wire G786_o2_n;
  wire G792_o2_p;
  wire G792_o2_n;
  wire G795_o2_p;
  wire G795_o2_n;
  wire G815_o2_p;
  wire G815_o2_n;
  wire G818_o2_p;
  wire G818_o2_n;
  wire G824_o2_p;
  wire G824_o2_n;
  wire G827_o2_p;
  wire G827_o2_n;
  wire G789_o2_p;
  wire G789_o2_n;
  wire G798_o2_p;
  wire G798_o2_n;
  wire G801_o2_p;
  wire G801_o2_n;
  wire G807_o2_p;
  wire G807_o2_n;
  wire G812_o2_p;
  wire G812_o2_n;
  wire G821_o2_p;
  wire G821_o2_n;
  wire G804_o2_p;
  wire G804_o2_n;
  wire G780_o2_p;
  wire G780_o2_n;
  wire G1231_o2_p;
  wire G1231_o2_n;
  wire G1572_o2_p;
  wire G1572_o2_n;
  wire G1377_o2_p;
  wire G1377_o2_n;
  wire G1253_o2_p;
  wire G1253_o2_n;
  wire G1359_o2_p;
  wire G1359_o2_n;
  wire G1258_o2_p;
  wire G1258_o2_n;
  wire G1367_o2_p;
  wire G1367_o2_n;
  wire G1358_o2_p;
  wire G1358_o2_n;
  wire G1366_o2_p;
  wire G1366_o2_n;
  wire G2057_o2_p;
  wire G2057_o2_n;
  wire G2117_o2_p;
  wire G2117_o2_n;
  wire G2118_o2_p;
  wire G2118_o2_n;
  wire G1254_o2_p;
  wire G1254_o2_n;
  wire G1259_o2_p;
  wire G1259_o2_n;
  wire G2058_o2_p;
  wire G2058_o2_n;
  wire G405_o2_p;
  wire G405_o2_n;
  wire G417_o2_p;
  wire G417_o2_n;
  wire G1269_o2_p;
  wire G1269_o2_n;
  wire G1275_o2_p;
  wire G1275_o2_n;
  wire G1287_o2_p;
  wire G1287_o2_n;
  wire G1266_o2_p;
  wire G1266_o2_n;
  wire G1272_o2_p;
  wire G1272_o2_n;
  wire G1278_o2_p;
  wire G1278_o2_n;
  wire G1281_o2_p;
  wire G1281_o2_n;
  wire G1284_o2_p;
  wire G1284_o2_n;
  wire G1290_o2_p;
  wire G1290_o2_n;
  wire G1293_o2_p;
  wire G1293_o2_n;
  wire G1299_o2_p;
  wire G1299_o2_n;
  wire G1305_o2_p;
  wire G1305_o2_n;
  wire G1296_o2_p;
  wire G1296_o2_n;
  wire G1302_o2_p;
  wire G1302_o2_n;
  wire G1308_o2_p;
  wire G1308_o2_n;
  wire G1311_o2_p;
  wire G1311_o2_n;
  wire G811_o2_p;
  wire G811_o2_n;
  wire G810_o2_p;
  wire G810_o2_n;
  wire G1728_o2_p;
  wire G1728_o2_n;
  wire G2512_o2_p;
  wire G2512_o2_n;
  wire G1114_o2_p;
  wire G1114_o2_n;
  wire G1113_o2_p;
  wire G1113_o2_n;
  wire G1992_o2_p;
  wire G1992_o2_n;
  wire G1991_o2_p;
  wire G1991_o2_n;
  wire G1426_o2_p;
  wire G1426_o2_n;
  wire G1966_o2_p;
  wire G1966_o2_n;
  wire G2211_o2_p;
  wire G2211_o2_n;
  wire G1509_o2_p;
  wire G1509_o2_n;
  wire G2153_o2_p;
  wire G2153_o2_n;
  wire G2329_o2_p;
  wire G2329_o2_n;
  wire G1540_o2_p;
  wire G1540_o2_n;
  wire G2167_o2_p;
  wire G2167_o2_n;
  wire G2191_o2_p;
  wire G2191_o2_n;
  wire G1234_o2_p;
  wire G1234_o2_n;
  wire G1132_o2_p;
  wire G1132_o2_n;
  wire G1129_o2_p;
  wire G1129_o2_n;
  wire G2088_o2_p;
  wire G2088_o2_n;
  wire G2106_o2_p;
  wire G2106_o2_n;
  wire G1314_o2_p;
  wire G1314_o2_n;
  wire G636_o2_p;
  wire G636_o2_n;
  wire G647_o2_p;
  wire G647_o2_n;
  wire n3186_lo_buf_o2_p;
  wire n3186_lo_buf_o2_n;
  wire n3198_lo_buf_o2_p;
  wire n3198_lo_buf_o2_n;
  wire n3210_lo_buf_o2_p;
  wire n3210_lo_buf_o2_n;
  wire n3222_lo_buf_o2_p;
  wire n3222_lo_buf_o2_n;
  wire G1225_o2_p;
  wire G1225_o2_n;
  wire G1342_o2_p;
  wire G1342_o2_n;
  wire G1222_o2_p;
  wire G1222_o2_n;
  wire G1228_o2_p;
  wire G1228_o2_n;
  wire G1348_o2_p;
  wire G1348_o2_n;
  wire G1345_o2_p;
  wire G1345_o2_n;
  wire G1351_o2_p;
  wire G1351_o2_n;
  wire G2242_o2_p;
  wire G2242_o2_n;
  wire G2260_o2_p;
  wire G2260_o2_n;
  wire G1374_o2_p;
  wire G1374_o2_n;
  wire G1537_o2_p;
  wire G1537_o2_n;
  wire G301_o2_p;
  wire G301_o2_n;
  wire G313_o2_p;
  wire G313_o2_n;
  wire G2365_o2_p;
  wire G2365_o2_n;
  wire G2255_o2_p;
  wire G2255_o2_n;
  wire G2253_o2_p;
  wire G2253_o2_n;
  wire G2395_o2_p;
  wire G2395_o2_n;
  wire G2272_o2_p;
  wire G2272_o2_n;
  wire G2270_o2_p;
  wire G2270_o2_n;
  wire G2245_o2_p;
  wire G2245_o2_n;
  wire G2262_o2_p;
  wire G2262_o2_n;
  wire G2249_o2_p;
  wire G2249_o2_n;
  wire G2247_o2_p;
  wire G2247_o2_n;
  wire G2266_o2_p;
  wire G2266_o2_n;
  wire G2264_o2_p;
  wire G2264_o2_n;
  wire G2403_o2_p;
  wire G2403_o2_n;
  wire G2401_o2_p;
  wire G2401_o2_n;
  wire G2410_o2_p;
  wire G2410_o2_n;
  wire G2408_o2_p;
  wire G2408_o2_n;
  wire G2306_o2_p;
  wire G2306_o2_n;
  wire G2305_o2_p;
  wire G2305_o2_n;
  wire G2314_o2_p;
  wire G2314_o2_n;
  wire G2313_o2_p;
  wire G2313_o2_n;
  wire G2303_o2_p;
  wire G2303_o2_n;
  wire G2302_o2_p;
  wire G2302_o2_n;
  wire G2301_o2_p;
  wire G2301_o2_n;
  wire G2311_o2_p;
  wire G2311_o2_n;
  wire G2310_o2_p;
  wire G2310_o2_n;
  wire G2309_o2_p;
  wire G2309_o2_n;
  wire G2404_o2_p;
  wire G2404_o2_n;
  wire G2411_o2_p;
  wire G2411_o2_n;
  wire G2420_o2_p;
  wire G2420_o2_n;
  wire G2419_o2_p;
  wire G2419_o2_n;
  wire G2433_o2_p;
  wire G2433_o2_n;
  wire G2432_o2_p;
  wire G2432_o2_n;
  wire G402_o2_p;
  wire G402_o2_n;
  wire G403_o2_p;
  wire G403_o2_n;
  wire G1053_o2_p;
  wire G1053_o2_n;
  wire G1049_o2_p;
  wire G1049_o2_n;
  wire n2003_inv_p;
  wire n2003_inv_n;
  wire G1364_o2_p;
  wire G1364_o2_n;
  wire G1079_o2_p;
  wire G1079_o2_n;
  wire G1478_o2_p;
  wire G1478_o2_n;
  wire G707_o2_p;
  wire G707_o2_n;
  wire G718_o2_p;
  wire G718_o2_n;
  wire G2417_o2_p;
  wire G2417_o2_n;
  wire G2414_o2_p;
  wire G2414_o2_n;
  wire G2431_o2_p;
  wire G2431_o2_n;
  wire G2428_o2_p;
  wire G2428_o2_n;
  wire G1653_o2_p;
  wire G1653_o2_n;
  wire G2213_o2_p;
  wire G2213_o2_n;
  wire G2221_o2_p;
  wire G2221_o2_n;
  wire G2250_o2_p;
  wire G2250_o2_n;
  wire G2267_o2_p;
  wire G2267_o2_n;
  wire G1365_o2_p;
  wire G1365_o2_n;
  wire G1368_o2_p;
  wire G1368_o2_n;
  wire G1371_o2_p;
  wire G1371_o2_n;
  wire G2218_o2_p;
  wire G2218_o2_n;
  wire G2225_o2_p;
  wire G2225_o2_n;
  wire n1503_lo_buf_o2_p;
  wire n1503_lo_buf_o2_n;
  wire n1863_lo_buf_o2_p;
  wire n1863_lo_buf_o2_n;
  wire n1887_lo_buf_o2_p;
  wire n1887_lo_buf_o2_n;
  wire n1983_lo_buf_o2_p;
  wire n1983_lo_buf_o2_n;
  wire n2007_lo_buf_o2_p;
  wire n2007_lo_buf_o2_n;
  wire n2115_lo_buf_o2_p;
  wire n2115_lo_buf_o2_n;
  wire n2139_lo_buf_o2_p;
  wire n2139_lo_buf_o2_n;
  wire n2247_lo_buf_o2_p;
  wire n2247_lo_buf_o2_n;
  wire n2271_lo_buf_o2_p;
  wire n2271_lo_buf_o2_n;
  wire n2919_lo_buf_o2_p;
  wire n2919_lo_buf_o2_n;
  wire n2943_lo_buf_o2_p;
  wire n2943_lo_buf_o2_n;
  wire n2967_lo_buf_o2_p;
  wire n2967_lo_buf_o2_n;
  wire n2979_lo_buf_o2_p;
  wire n2979_lo_buf_o2_n;
  wire n3063_lo_buf_o2_p;
  wire n3063_lo_buf_o2_n;
  wire n3075_lo_buf_o2_p;
  wire n3075_lo_buf_o2_n;
  wire n3099_lo_buf_o2_p;
  wire n3099_lo_buf_o2_n;
  wire n3111_lo_buf_o2_p;
  wire n3111_lo_buf_o2_n;
  wire G878_o2_p;
  wire G878_o2_n;
  wire G875_o2_p;
  wire G875_o2_n;
  wire G661_o2_p;
  wire G661_o2_n;
  wire G660_o2_p;
  wire G660_o2_n;
  wire G879_o2_p;
  wire G879_o2_n;
  wire G876_o2_p;
  wire G876_o2_n;
  wire G1320_o2_p;
  wire G1320_o2_n;
  wire G941_o2_p;
  wire G941_o2_n;
  wire G732_o2_p;
  wire G732_o2_n;
  wire G942_o2_p;
  wire G942_o2_n;
  wire G1493_o2_p;
  wire G1493_o2_n;
  wire G1498_o2_p;
  wire G1498_o2_n;
  wire G877_o2_p;
  wire G877_o2_n;
  wire G874_o2_p;
  wire G874_o2_n;
  wire n1806_lo_buf_o2_p;
  wire n1806_lo_buf_o2_n;
  wire n1878_lo_buf_o2_p;
  wire n1878_lo_buf_o2_n;
  wire n1938_lo_buf_o2_p;
  wire n1938_lo_buf_o2_n;
  wire n1998_lo_buf_o2_p;
  wire n1998_lo_buf_o2_n;
  wire n2058_lo_buf_o2_p;
  wire n2058_lo_buf_o2_n;
  wire n2130_lo_buf_o2_p;
  wire n2130_lo_buf_o2_n;
  wire n2190_lo_buf_o2_p;
  wire n2190_lo_buf_o2_n;
  wire n2262_lo_buf_o2_p;
  wire n2262_lo_buf_o2_n;
  wire n2310_lo_buf_o2_p;
  wire n2310_lo_buf_o2_n;
  wire n2406_lo_buf_o2_p;
  wire n2406_lo_buf_o2_n;
  wire n2430_lo_buf_o2_p;
  wire n2430_lo_buf_o2_n;
  wire n2526_lo_buf_o2_p;
  wire n2526_lo_buf_o2_n;
  wire n2550_lo_buf_o2_p;
  wire n2550_lo_buf_o2_n;
  wire n2646_lo_buf_o2_p;
  wire n2646_lo_buf_o2_n;
  wire n2670_lo_buf_o2_p;
  wire n2670_lo_buf_o2_n;
  wire n2766_lo_buf_o2_p;
  wire n2766_lo_buf_o2_n;
  wire G603_o2_p;
  wire G603_o2_n;
  wire G614_o2_p;
  wire G614_o2_n;
  wire G1026_o2_p;
  wire G1026_o2_n;
  wire G1021_o2_p;
  wire G1021_o2_n;
  wire G940_o2_p;
  wire G940_o2_n;
  wire G1636_o2_p;
  wire G1636_o2_n;
  wire G1684_o2_p;
  wire G1684_o2_n;
  wire n2352_lo_buf_o2_p;
  wire n2352_lo_buf_o2_n;
  wire n2364_lo_buf_o2_p;
  wire n2364_lo_buf_o2_n;
  wire n2472_lo_buf_o2_p;
  wire n2472_lo_buf_o2_n;
  wire n2484_lo_buf_o2_p;
  wire n2484_lo_buf_o2_n;
  wire n2592_lo_buf_o2_p;
  wire n2592_lo_buf_o2_n;
  wire n2604_lo_buf_o2_p;
  wire n2604_lo_buf_o2_n;
  wire n2712_lo_buf_o2_p;
  wire n2712_lo_buf_o2_n;
  wire n2724_lo_buf_o2_p;
  wire n2724_lo_buf_o2_n;
  wire n3150_lo_buf_o2_p;
  wire n3150_lo_buf_o2_n;
  wire n3162_lo_buf_o2_p;
  wire n3162_lo_buf_o2_n;
  wire g835_p;
  wire g835_n;
  wire g836_p;
  wire g836_n;
  wire g837_p;
  wire g837_n;
  wire g838_p;
  wire g838_n;
  wire g839_p;
  wire g839_n;
  wire g840_p;
  wire g840_n;
  wire g841_p;
  wire g841_n;
  wire g842_p;
  wire g842_n;
  wire g843_p;
  wire g843_n;
  wire g844_p;
  wire g844_n;
  wire g845_p;
  wire g845_n;
  wire g846_p;
  wire g846_n;
  wire g847_p;
  wire g847_n;
  wire g848_p;
  wire g848_n;
  wire g849_p;
  wire g849_n;
  wire g850_p;
  wire g850_n;
  wire g851_p;
  wire g851_n;
  wire g852_p;
  wire g852_n;
  wire g853_p;
  wire g853_n;
  wire g854_p;
  wire g854_n;
  wire g855_p;
  wire g855_n;
  wire g856_p;
  wire g856_n;
  wire g857_p;
  wire g857_n;
  wire g858_p;
  wire g858_n;
  wire g859_p;
  wire g859_n;
  wire g860_p;
  wire g860_n;
  wire g861_p;
  wire g861_n;
  wire g862_p;
  wire g862_n;
  wire g863_p;
  wire g863_n;
  wire g864_p;
  wire g864_n;
  wire g865_p;
  wire g865_n;
  wire g866_p;
  wire g866_n;
  wire g867_p;
  wire g867_n;
  wire g868_p;
  wire g868_n;
  wire g869_p;
  wire g869_n;
  wire g870_p;
  wire g870_n;
  wire g871_p;
  wire g871_n;
  wire g872_p;
  wire g872_n;
  wire g873_p;
  wire g873_n;
  wire g874_p;
  wire g874_n;
  wire g875_p;
  wire g875_n;
  wire g876_p;
  wire g876_n;
  wire g877_p;
  wire g877_n;
  wire g878_p;
  wire g878_n;
  wire g879_p;
  wire g879_n;
  wire g880_p;
  wire g880_n;
  wire g881_p;
  wire g881_n;
  wire g882_p;
  wire g882_n;
  wire g883_p;
  wire g883_n;
  wire g884_p;
  wire g884_n;
  wire g885_p;
  wire g885_n;
  wire g886_p;
  wire g886_n;
  wire g887_p;
  wire g887_n;
  wire g888_p;
  wire g888_n;
  wire g889_p;
  wire g889_n;
  wire g890_p;
  wire g890_n;
  wire g891_p;
  wire g891_n;
  wire g892_p;
  wire g892_n;
  wire g893_p;
  wire g893_n;
  wire g894_p;
  wire g894_n;
  wire g895_p;
  wire g895_n;
  wire g896_p;
  wire g896_n;
  wire g897_p;
  wire g897_n;
  wire g898_p;
  wire g898_n;
  wire g899_p;
  wire g899_n;
  wire g900_p;
  wire g900_n;
  wire g901_p;
  wire g901_n;
  wire g902_p;
  wire g902_n;
  wire g903_p;
  wire g903_n;
  wire g904_p;
  wire g904_n;
  wire g905_p;
  wire g905_n;
  wire g906_p;
  wire g906_n;
  wire g907_p;
  wire g907_n;
  wire g908_p;
  wire g908_n;
  wire g909_p;
  wire g909_n;
  wire g910_p;
  wire g910_n;
  wire g911_p;
  wire g911_n;
  wire g912_p;
  wire g912_n;
  wire g913_p;
  wire g913_n;
  wire g914_p;
  wire g914_n;
  wire g915_p;
  wire g915_n;
  wire g916_p;
  wire g916_n;
  wire g917_p;
  wire g917_n;
  wire g918_p;
  wire g918_n;
  wire g919_p;
  wire g919_n;
  wire g920_p;
  wire g920_n;
  wire g921_p;
  wire g921_n;
  wire g922_p;
  wire g922_n;
  wire g923_p;
  wire g923_n;
  wire g924_p;
  wire g924_n;
  wire g925_p;
  wire g925_n;
  wire g926_p;
  wire g926_n;
  wire g927_p;
  wire g927_n;
  wire g928_p;
  wire g928_n;
  wire g929_p;
  wire g929_n;
  wire g930_p;
  wire g930_n;
  wire g931_p;
  wire g931_n;
  wire g932_p;
  wire g932_n;
  wire g933_p;
  wire g933_n;
  wire g934_p;
  wire g934_n;
  wire g935_p;
  wire g935_n;
  wire g936_p;
  wire g936_n;
  wire g937_p;
  wire g937_n;
  wire g938_p;
  wire g938_n;
  wire g939_p;
  wire g939_n;
  wire g940_p;
  wire g940_n;
  wire g941_p;
  wire g941_n;
  wire g942_p;
  wire g942_n;
  wire g943_p;
  wire g943_n;
  wire g944_p;
  wire g944_n;
  wire g945_p;
  wire g945_n;
  wire g946_p;
  wire g946_n;
  wire g947_p;
  wire g947_n;
  wire g948_p;
  wire g948_n;
  wire g949_p;
  wire g949_n;
  wire g950_p;
  wire g950_n;
  wire g951_p;
  wire g951_n;
  wire g952_p;
  wire g952_n;
  wire g953_p;
  wire g953_n;
  wire g954_p;
  wire g954_n;
  wire g955_p;
  wire g955_n;
  wire g956_p;
  wire g956_n;
  wire g957_p;
  wire g957_n;
  wire g958_p;
  wire g958_n;
  wire g959_p;
  wire g959_n;
  wire g960_p;
  wire g960_n;
  wire g961_p;
  wire g961_n;
  wire g962_p;
  wire g962_n;
  wire g963_p;
  wire g963_n;
  wire g964_p;
  wire g964_n;
  wire g965_p;
  wire g965_n;
  wire g966_p;
  wire g966_n;
  wire g967_p;
  wire g967_n;
  wire g968_p;
  wire g968_n;
  wire g969_p;
  wire g969_n;
  wire g970_p;
  wire g970_n;
  wire g971_p;
  wire g971_n;
  wire g972_p;
  wire g972_n;
  wire g973_p;
  wire g973_n;
  wire g974_p;
  wire g974_n;
  wire g975_p;
  wire g975_n;
  wire g976_p;
  wire g976_n;
  wire g977_p;
  wire g977_n;
  wire g978_p;
  wire g978_n;
  wire g979_p;
  wire g979_n;
  wire g980_p;
  wire g980_n;
  wire g981_p;
  wire g981_n;
  wire g982_p;
  wire g982_n;
  wire g983_p;
  wire g983_n;
  wire g984_p;
  wire g984_n;
  wire g985_p;
  wire g985_n;
  wire g986_p;
  wire g986_n;
  wire g987_p;
  wire g987_n;
  wire g988_p;
  wire g988_n;
  wire g989_p;
  wire g989_n;
  wire g990_p;
  wire g990_n;
  wire g991_p;
  wire g991_n;
  wire g992_p;
  wire g992_n;
  wire g993_p;
  wire g993_n;
  wire g994_p;
  wire g994_n;
  wire g995_p;
  wire g995_n;
  wire g996_p;
  wire g996_n;
  wire g997_p;
  wire g997_n;
  wire g998_p;
  wire g998_n;
  wire g999_p;
  wire g999_n;
  wire g1000_p;
  wire g1000_n;
  wire g1001_p;
  wire g1001_n;
  wire g1002_p;
  wire g1002_n;
  wire g1003_p;
  wire g1003_n;
  wire g1004_p;
  wire g1004_n;
  wire g1005_p;
  wire g1005_n;
  wire g1006_p;
  wire g1006_n;
  wire g1007_p;
  wire g1007_n;
  wire g1008_p;
  wire g1008_n;
  wire g1009_p;
  wire g1009_n;
  wire g1010_p;
  wire g1010_n;
  wire g1011_p;
  wire g1011_n;
  wire g1012_p;
  wire g1012_n;
  wire g1013_p;
  wire g1013_n;
  wire g1014_p;
  wire g1014_n;
  wire g1015_p;
  wire g1015_n;
  wire g1016_p;
  wire g1016_n;
  wire g1017_p;
  wire g1017_n;
  wire g1018_p;
  wire g1018_n;
  wire g1019_p;
  wire g1019_n;
  wire g1020_p;
  wire g1020_n;
  wire g1021_p;
  wire g1021_n;
  wire g1022_p;
  wire g1022_n;
  wire g1023_p;
  wire g1023_n;
  wire g1024_p;
  wire g1024_n;
  wire g1025_p;
  wire g1025_n;
  wire g1026_p;
  wire g1026_n;
  wire g1027_p;
  wire g1027_n;
  wire g1028_p;
  wire g1028_n;
  wire g1029_p;
  wire g1029_n;
  wire g1030_p;
  wire g1030_n;
  wire g1031_p;
  wire g1031_n;
  wire g1032_p;
  wire g1032_n;
  wire g1033_p;
  wire g1033_n;
  wire g1034_p;
  wire g1034_n;
  wire g1035_p;
  wire g1035_n;
  wire g1036_p;
  wire g1036_n;
  wire g1037_p;
  wire g1037_n;
  wire g1038_p;
  wire g1038_n;
  wire g1039_p;
  wire g1039_n;
  wire g1040_p;
  wire g1040_n;
  wire g1041_p;
  wire g1041_n;
  wire g1042_p;
  wire g1042_n;
  wire g1043_p;
  wire g1043_n;
  wire g1044_p;
  wire g1044_n;
  wire g1045_p;
  wire g1045_n;
  wire g1046_p;
  wire g1046_n;
  wire g1047_p;
  wire g1047_n;
  wire g1048_p;
  wire g1048_n;
  wire g1049_p;
  wire g1049_n;
  wire g1050_p;
  wire g1050_n;
  wire g1051_p;
  wire g1051_n;
  wire g1052_p;
  wire g1052_n;
  wire g1053_p;
  wire g1053_n;
  wire g1054_p;
  wire g1054_n;
  wire g1055_p;
  wire g1055_n;
  wire g1056_p;
  wire g1056_n;
  wire g1057_p;
  wire g1057_n;
  wire g1058_p;
  wire g1058_n;
  wire g1059_p;
  wire g1059_n;
  wire g1060_p;
  wire g1060_n;
  wire g1061_p;
  wire g1061_n;
  wire g1062_p;
  wire g1062_n;
  wire g1063_p;
  wire g1063_n;
  wire g1064_p;
  wire g1064_n;
  wire g1065_p;
  wire g1065_n;
  wire g1066_p;
  wire g1066_n;
  wire g1067_p;
  wire g1067_n;
  wire g1068_p;
  wire g1068_n;
  wire g1069_p;
  wire g1069_n;
  wire g1070_p;
  wire g1070_n;
  wire g1071_p;
  wire g1071_n;
  wire g1072_p;
  wire g1072_n;
  wire g1073_p;
  wire g1073_n;
  wire g1074_p;
  wire g1074_n;
  wire g1075_p;
  wire g1075_n;
  wire g1076_p;
  wire g1076_n;
  wire g1077_p;
  wire g1077_n;
  wire g1078_p;
  wire g1078_n;
  wire g1079_p;
  wire g1079_n;
  wire g1080_p;
  wire g1080_n;
  wire g1081_p;
  wire g1081_n;
  wire g1082_p;
  wire g1082_n;
  wire g1083_p;
  wire g1083_n;
  wire g1084_p;
  wire g1084_n;
  wire g1085_p;
  wire g1085_n;
  wire g1086_p;
  wire g1086_n;
  wire g1087_p;
  wire g1087_n;
  wire g1088_p;
  wire g1088_n;
  wire g1089_p;
  wire g1089_n;
  wire g1090_p;
  wire g1090_n;
  wire g1091_p;
  wire g1091_n;
  wire g1092_p;
  wire g1092_n;
  wire g1093_p;
  wire g1093_n;
  wire g1094_p;
  wire g1094_n;
  wire g1095_p;
  wire g1095_n;
  wire g1096_p;
  wire g1096_n;
  wire g1097_p;
  wire g1097_n;
  wire g1098_p;
  wire g1098_n;
  wire g1099_p;
  wire g1099_n;
  wire g1100_p;
  wire g1100_n;
  wire g1101_p;
  wire g1101_n;
  wire g1102_p;
  wire g1102_n;
  wire g1103_p;
  wire g1103_n;
  wire g1104_p;
  wire g1104_n;
  wire g1105_p;
  wire g1105_n;
  wire g1106_p;
  wire g1106_n;
  wire g1107_p;
  wire g1107_n;
  wire g1108_p;
  wire g1108_n;
  wire g1109_p;
  wire g1109_n;
  wire g1110_p;
  wire g1110_n;
  wire g1111_p;
  wire g1111_n;
  wire g1112_p;
  wire g1112_n;
  wire g1113_p;
  wire g1113_n;
  wire g1114_p;
  wire g1114_n;
  wire g1115_p;
  wire g1115_n;
  wire g1116_p;
  wire g1116_n;
  wire g1117_p;
  wire g1117_n;
  wire g1118_p;
  wire g1118_n;
  wire g1119_p;
  wire g1119_n;
  wire g1120_p;
  wire g1120_n;
  wire g1121_p;
  wire g1121_n;
  wire g1122_p;
  wire g1122_n;
  wire g1123_p;
  wire g1123_n;
  wire g1124_p;
  wire g1124_n;
  wire g1125_p;
  wire g1125_n;
  wire g1126_p;
  wire g1126_n;
  wire g1127_p;
  wire g1127_n;
  wire g1128_p;
  wire g1128_n;
  wire g1129_p;
  wire g1129_n;
  wire g1130_p;
  wire g1130_n;
  wire g1131_p;
  wire g1131_n;
  wire g1132_p;
  wire g1132_n;
  wire g1133_p;
  wire g1133_n;
  wire g1134_p;
  wire g1134_n;
  wire g1135_p;
  wire g1135_n;
  wire g1136_p;
  wire g1136_n;
  wire g1137_p;
  wire g1137_n;
  wire g1138_p;
  wire g1138_n;
  wire g1139_p;
  wire g1139_n;
  wire g1140_p;
  wire g1140_n;
  wire g1141_p;
  wire g1141_n;
  wire g1142_p;
  wire g1142_n;
  wire g1143_p;
  wire g1143_n;
  wire g1144_p;
  wire g1144_n;
  wire g1145_p;
  wire g1145_n;
  wire g1146_p;
  wire g1146_n;
  wire g1147_p;
  wire g1147_n;
  wire g1148_p;
  wire g1148_n;
  wire g1149_p;
  wire g1149_n;
  wire g1150_p;
  wire g1150_n;
  wire g1151_p;
  wire g1151_n;
  wire g1152_p;
  wire g1152_n;
  wire g1153_p;
  wire g1153_n;
  wire g1154_p;
  wire g1154_n;
  wire g1155_p;
  wire g1155_n;
  wire g1156_p;
  wire g1156_n;
  wire g1157_p;
  wire g1157_n;
  wire g1158_p;
  wire g1158_n;
  wire g1159_p;
  wire g1159_n;
  wire g1160_p;
  wire g1160_n;
  wire g1161_p;
  wire g1161_n;
  wire g1162_p;
  wire g1162_n;
  wire g1163_p;
  wire g1163_n;
  wire g1164_p;
  wire g1164_n;
  wire g1165_p;
  wire g1165_n;
  wire g1166_p;
  wire g1166_n;
  wire g1167_p;
  wire g1167_n;
  wire g1168_p;
  wire g1168_n;
  wire g1169_p;
  wire g1169_n;
  wire g1170_p;
  wire g1170_n;
  wire g1171_p;
  wire g1171_n;
  wire g1172_p;
  wire g1172_n;
  wire g1173_p;
  wire g1173_n;
  wire g1174_p;
  wire g1174_n;
  wire g1175_p;
  wire g1175_n;
  wire g1176_p;
  wire g1176_n;
  wire g1177_p;
  wire g1177_n;
  wire g1178_p;
  wire g1178_n;
  wire g1179_p;
  wire g1179_n;
  wire g1180_p;
  wire g1180_n;
  wire g1181_p;
  wire g1181_n;
  wire g1182_p;
  wire g1182_n;
  wire g1183_p;
  wire g1183_n;
  wire g1184_p;
  wire g1184_n;
  wire g1185_p;
  wire g1185_n;
  wire g1186_p;
  wire g1186_n;
  wire g1187_p;
  wire g1187_n;
  wire g1188_p;
  wire g1188_n;
  wire g1189_p;
  wire g1189_n;
  wire g1190_p;
  wire g1190_n;
  wire g1191_p;
  wire g1191_n;
  wire g1192_p;
  wire g1192_n;
  wire g1193_p;
  wire g1193_n;
  wire g1194_p;
  wire g1194_n;
  wire g1195_p;
  wire g1195_n;
  wire g1196_p;
  wire g1196_n;
  wire g1197_p;
  wire g1197_n;
  wire g1198_p;
  wire g1198_n;
  wire g1199_p;
  wire g1199_n;
  wire g1200_p;
  wire g1200_n;
  wire g1201_p;
  wire g1201_n;
  wire g1202_p;
  wire g1202_n;
  wire g1203_p;
  wire g1203_n;
  wire g1204_p;
  wire g1204_n;
  wire g1205_p;
  wire g1205_n;
  wire g1206_p;
  wire g1206_n;
  wire g1207_p;
  wire g1207_n;
  wire g1208_p;
  wire g1208_n;
  wire g1209_p;
  wire g1209_n;
  wire g1210_p;
  wire g1210_n;
  wire g1211_p;
  wire g1211_n;
  wire g1212_p;
  wire g1212_n;
  wire g1213_p;
  wire g1213_n;
  wire g1214_p;
  wire g1214_n;
  wire g1215_p;
  wire g1215_n;
  wire g1216_p;
  wire g1216_n;
  wire g1217_p;
  wire g1217_n;
  wire g1218_p;
  wire g1218_n;
  wire g1219_p;
  wire g1219_n;
  wire g1220_p;
  wire g1220_n;
  wire g1221_p;
  wire g1221_n;
  wire g1222_p;
  wire g1222_n;
  wire g1223_p;
  wire g1223_n;
  wire g1224_p;
  wire g1224_n;
  wire g1225_p;
  wire g1225_n;
  wire g1226_p;
  wire g1226_n;
  wire g1227_p;
  wire g1227_n;
  wire g1228_p;
  wire g1228_n;
  wire g1229_p;
  wire g1229_n;
  wire g1230_p;
  wire g1230_n;
  wire g1231_p;
  wire g1231_n;
  wire g1232_p;
  wire g1232_n;
  wire g1233_p;
  wire g1233_n;
  wire g1234_p;
  wire g1234_n;
  wire g1235_p;
  wire g1235_n;
  wire g1236_p;
  wire g1236_n;
  wire g1237_p;
  wire g1237_n;
  wire g1238_p;
  wire g1238_n;
  wire g1239_p;
  wire g1239_n;
  wire g1240_p;
  wire g1240_n;
  wire g1241_p;
  wire g1241_n;
  wire g1242_p;
  wire g1242_n;
  wire g1243_p;
  wire g1243_n;
  wire g1244_p;
  wire g1244_n;
  wire g1245_p;
  wire g1245_n;
  wire g1246_p;
  wire g1246_n;
  wire g1247_p;
  wire g1247_n;
  wire g1248_p;
  wire g1248_n;
  wire g1249_p;
  wire g1249_n;
  wire g1250_p;
  wire g1250_n;
  wire g1251_p;
  wire g1251_n;
  wire g1252_p;
  wire g1252_n;
  wire g1253_p;
  wire g1253_n;
  wire g1254_p;
  wire g1254_n;
  wire g1255_p;
  wire g1255_n;
  wire g1256_p;
  wire g1256_n;
  wire g1257_p;
  wire g1257_n;
  wire g1258_p;
  wire g1258_n;
  wire g1259_p;
  wire g1259_n;
  wire g1260_p;
  wire g1260_n;
  wire g1261_p;
  wire g1261_n;
  wire g1262_p;
  wire g1262_n;
  wire g1263_p;
  wire g1263_n;
  wire g1264_p;
  wire g1264_n;
  wire g1265_p;
  wire g1265_n;
  wire g1266_p;
  wire g1266_n;
  wire g1267_p;
  wire g1267_n;
  wire g1268_p;
  wire g1268_n;
  wire g1269_p;
  wire g1269_n;
  wire g1270_p;
  wire g1270_n;
  wire g1271_p;
  wire g1271_n;
  wire g1272_p;
  wire g1272_n;
  wire g1273_p;
  wire g1273_n;
  wire g1274_p;
  wire g1274_n;
  wire g1275_p;
  wire g1275_n;
  wire g1276_p;
  wire g1276_n;
  wire g1277_p;
  wire g1277_n;
  wire g1278_p;
  wire g1278_n;
  wire g1279_p;
  wire g1279_n;
  wire g1280_p;
  wire g1280_n;
  wire g1281_p;
  wire g1281_n;
  wire g1282_p;
  wire g1282_n;
  wire g1283_p;
  wire g1283_n;
  wire g1284_p;
  wire g1284_n;
  wire g1285_p;
  wire g1285_n;
  wire g1286_p;
  wire g1286_n;
  wire g1287_p;
  wire g1287_n;
  wire g1288_p;
  wire g1288_n;
  wire g1289_p;
  wire g1289_n;
  wire g1290_p;
  wire g1290_n;
  wire g1291_p;
  wire g1291_n;
  wire g1292_p;
  wire g1292_n;
  wire g1293_p;
  wire g1293_n;
  wire g1294_p;
  wire g1294_n;
  wire g1295_p;
  wire g1295_n;
  wire g1296_p;
  wire g1296_n;
  wire g1297_p;
  wire g1297_n;
  wire g1298_p;
  wire g1298_n;
  wire g1299_p;
  wire g1299_n;
  wire g1300_p;
  wire g1300_n;
  wire g1301_p;
  wire g1301_n;
  wire g1302_p;
  wire g1302_n;
  wire g1303_p;
  wire g1303_n;
  wire g1304_p;
  wire g1304_n;
  wire g1305_p;
  wire g1305_n;
  wire g1306_p;
  wire g1306_n;
  wire g1307_p;
  wire g1307_n;
  wire g1308_p;
  wire g1308_n;
  wire g1309_p;
  wire g1309_n;
  wire g1310_p;
  wire g1310_n;
  wire g1311_p;
  wire g1311_n;
  wire g1312_p;
  wire g1312_n;
  wire g1313_p;
  wire g1313_n;
  wire g1314_p;
  wire g1314_n;
  wire g1315_p;
  wire g1315_n;
  wire g1316_p;
  wire g1316_n;
  wire g1317_p;
  wire g1317_n;
  wire g1318_p;
  wire g1318_n;
  wire g1319_p;
  wire g1319_n;
  wire g1320_p;
  wire g1320_n;
  wire g1321_p;
  wire g1321_n;
  wire g1322_p;
  wire g1322_n;
  wire g1323_p;
  wire g1323_n;
  wire g1324_p;
  wire g1324_n;
  wire g1325_p;
  wire g1325_n;
  wire g1326_p;
  wire g1326_n;
  wire g1327_p;
  wire g1327_n;
  wire g1328_p;
  wire g1328_n;
  wire g1329_p;
  wire g1329_n;
  wire g1330_p;
  wire g1330_n;
  wire g1331_p;
  wire g1331_n;
  wire g1332_p;
  wire g1332_n;
  wire g1333_p;
  wire g1333_n;
  wire g1334_p;
  wire g1334_n;
  wire g1335_p;
  wire g1335_n;
  wire g1336_p;
  wire g1336_n;
  wire g1337_p;
  wire g1337_n;
  wire g1338_p;
  wire g1338_n;
  wire g1339_p;
  wire g1339_n;
  wire g1340_p;
  wire g1340_n;
  wire g1341_p;
  wire g1341_n;
  wire g1342_p;
  wire g1342_n;
  wire g1343_p;
  wire g1343_n;
  wire g1344_p;
  wire g1344_n;
  wire g1345_p;
  wire g1345_n;
  wire g1346_p;
  wire g1346_n;
  wire g1347_p;
  wire g1347_n;
  wire g1348_p;
  wire g1348_n;
  wire g1349_p;
  wire g1349_n;
  wire g1350_p;
  wire g1350_n;
  wire g1351_p;
  wire g1351_n;
  wire g1352_p;
  wire g1352_n;
  wire g1353_p;
  wire g1353_n;
  wire g1354_p;
  wire g1354_n;
  wire g1355_p;
  wire g1355_n;
  wire g1356_p;
  wire g1356_n;
  wire g1357_p;
  wire g1357_n;
  wire g1358_p;
  wire g1358_n;
  wire g1359_p;
  wire g1359_n;
  wire g1360_p;
  wire g1360_n;
  wire g1361_p;
  wire g1361_n;
  wire g1362_p;
  wire g1362_n;
  wire g1363_p;
  wire g1363_n;
  wire g1364_p;
  wire g1364_n;
  wire g1365_p;
  wire g1365_n;
  wire g1366_p;
  wire g1366_n;
  wire g1367_p;
  wire g1367_n;
  wire g1368_p;
  wire g1368_n;
  wire g1369_p;
  wire g1369_n;
  wire g1370_p;
  wire g1370_n;
  wire g1371_p;
  wire g1371_n;
  wire g1372_p;
  wire g1372_n;
  wire g1373_p;
  wire g1373_n;
  wire g1374_p;
  wire g1374_n;
  wire g1375_p;
  wire g1375_n;
  wire g1376_p;
  wire g1376_n;
  wire g1377_p;
  wire g1377_n;
  wire g1378_p;
  wire g1378_n;
  wire g1379_p;
  wire g1379_n;
  wire g1380_p;
  wire g1380_n;
  wire g1381_p;
  wire g1381_n;
  wire g1382_p;
  wire g1382_n;
  wire g1383_p;
  wire g1383_n;
  wire g1384_p;
  wire g1384_n;
  wire g1385_p;
  wire g1385_n;
  wire g1386_p;
  wire g1386_n;
  wire g1387_p;
  wire g1387_n;
  wire g1388_p;
  wire g1388_n;
  wire g1389_p;
  wire g1389_n;
  wire g1390_p;
  wire g1390_n;
  wire g1391_p;
  wire g1391_n;
  wire g1392_p;
  wire g1392_n;
  wire g1393_p;
  wire g1393_n;
  wire g1394_p;
  wire g1394_n;
  wire g1395_p;
  wire g1395_n;
  wire g1396_p;
  wire g1396_n;
  wire g1397_p;
  wire g1397_n;
  wire g1398_p;
  wire g1398_n;
  wire g1399_p;
  wire g1399_n;
  wire g1400_p;
  wire g1400_n;
  wire g1401_p;
  wire g1401_n;
  wire g1402_p;
  wire g1402_n;
  wire g1403_p;
  wire g1403_n;
  wire g1404_p;
  wire g1404_n;
  wire g1405_p;
  wire g1405_n;
  wire g1406_p;
  wire g1406_n;
  wire g1407_p;
  wire g1407_n;
  wire g1408_p;
  wire g1408_n;
  wire g1409_p;
  wire g1409_n;
  wire g1410_p;
  wire g1410_n;
  wire g1411_p;
  wire g1411_n;
  wire g1412_p;
  wire g1412_n;
  wire g1413_p;
  wire g1413_n;
  wire g1414_p;
  wire g1414_n;
  wire g1415_p;
  wire g1415_n;
  wire g1416_p;
  wire g1416_n;
  wire g1417_p;
  wire g1417_n;
  wire g1418_p;
  wire g1418_n;
  wire g1419_p;
  wire g1419_n;
  wire g1420_p;
  wire g1420_n;
  wire g1421_p;
  wire g1421_n;
  wire g1422_p;
  wire g1422_n;
  wire g1423_p;
  wire g1423_n;
  wire g1424_p;
  wire g1424_n;
  wire g1425_p;
  wire g1425_n;
  wire g1426_p;
  wire g1426_n;
  wire g1427_p;
  wire g1427_n;
  wire g1428_p;
  wire g1428_n;
  wire g1429_p;
  wire g1429_n;
  wire g1430_p;
  wire g1430_n;
  wire g1431_p;
  wire g1431_n;
  wire g1432_p;
  wire g1432_n;
  wire g1433_p;
  wire g1433_n;
  wire g1434_p;
  wire g1434_n;
  wire g1435_p;
  wire g1435_n;
  wire g1436_p;
  wire g1436_n;
  wire g1437_p;
  wire g1437_n;
  wire g1438_p;
  wire g1438_n;
  wire g1439_p;
  wire g1439_n;
  wire g1440_p;
  wire g1440_n;
  wire g1441_p;
  wire g1441_n;
  wire g1442_p;
  wire g1442_n;
  wire g1443_p;
  wire g1443_n;
  wire g1444_p;
  wire g1444_n;
  wire g1445_p;
  wire g1445_n;
  wire g1446_p;
  wire g1446_n;
  wire g1447_p;
  wire g1447_n;
  wire g1448_p;
  wire g1448_n;
  wire g1449_p;
  wire g1449_n;
  wire g1450_p;
  wire g1450_n;
  wire g1451_p;
  wire g1451_n;
  wire g1452_p;
  wire g1452_n;
  wire g1453_p;
  wire g1453_n;
  wire g1454_p;
  wire g1454_n;
  wire g1455_p;
  wire g1455_n;
  wire g1456_p;
  wire g1456_n;
  wire g1457_p;
  wire g1457_n;
  wire g1458_p;
  wire g1458_n;
  wire g1459_p;
  wire g1459_n;
  wire g1460_p;
  wire g1460_n;
  wire g1461_p;
  wire g1461_n;
  wire g1462_p;
  wire g1462_n;
  wire g1463_p;
  wire g1463_n;
  wire g1464_p;
  wire g1464_n;
  wire g1465_p;
  wire g1465_n;
  wire g1466_p;
  wire g1466_n;
  wire g1467_p;
  wire g1467_n;
  wire g1468_p;
  wire g1468_n;
  wire g1469_p;
  wire g1469_n;
  wire g1470_p;
  wire g1470_n;
  wire g1471_p;
  wire g1471_n;
  wire g1472_p;
  wire g1472_n;
  wire g1473_p;
  wire g1473_n;
  wire g1474_p;
  wire g1474_n;
  wire g1475_p;
  wire g1475_n;
  wire g1476_p;
  wire g1476_n;
  wire g1477_p;
  wire g1477_n;
  wire g1478_p;
  wire g1478_n;
  wire g1479_p;
  wire g1479_n;
  wire g1480_p;
  wire g1480_n;
  wire g1481_p;
  wire g1481_n;
  wire g1482_p;
  wire g1482_n;
  wire g1483_p;
  wire g1483_n;
  wire g1484_p;
  wire g1484_n;
  wire g1485_p;
  wire g1485_n;
  wire g1486_p;
  wire g1486_n;
  wire g1487_p;
  wire g1487_n;
  wire g1488_p;
  wire g1488_n;
  wire g1489_p;
  wire g1489_n;
  wire g1490_p;
  wire g1490_n;
  wire g1491_p;
  wire g1491_n;
  wire g1492_p;
  wire g1492_n;
  wire g1493_p;
  wire g1493_n;
  wire g1494_p;
  wire g1494_n;
  wire g1495_p;
  wire g1495_n;
  wire g1496_p;
  wire g1496_n;
  wire g1497_p;
  wire g1497_n;
  wire g1498_p;
  wire g1498_n;
  wire g1499_p;
  wire g1499_n;
  wire g1500_p;
  wire g1500_n;
  wire g1501_p;
  wire g1501_n;
  wire g1502_p;
  wire g1502_n;
  wire g1503_p;
  wire g1503_n;
  wire g1504_p;
  wire g1504_n;
  wire g1505_p;
  wire g1505_n;
  wire g1506_p;
  wire g1506_n;
  wire g1507_p;
  wire g1507_n;
  wire g1508_p;
  wire g1508_n;
  wire g1509_p;
  wire g1509_n;
  wire g1510_p;
  wire g1510_n;
  wire g1511_p;
  wire g1511_n;
  wire g1512_p;
  wire g1512_n;
  wire g1513_p;
  wire g1513_n;
  wire g1514_p;
  wire g1514_n;
  wire g1515_p;
  wire g1515_n;
  wire g1516_p;
  wire g1516_n;
  wire g1517_p;
  wire g1517_n;
  wire g1518_p;
  wire g1518_n;
  wire g1519_p;
  wire g1519_n;
  wire g1520_p;
  wire g1520_n;
  wire g1521_p;
  wire g1521_n;
  wire g1522_p;
  wire g1522_n;
  wire g1523_p;
  wire g1523_n;
  wire g1524_p;
  wire g1524_n;
  wire g1525_p;
  wire g1525_n;
  wire g1526_p;
  wire g1526_n;
  wire g1527_p;
  wire g1527_n;
  wire g1528_p;
  wire g1528_n;
  wire g1529_p;
  wire g1529_n;
  wire g1530_p;
  wire g1530_n;
  wire g1531_p;
  wire g1531_n;
  wire g1532_p;
  wire g1532_n;
  wire g1533_p;
  wire g1533_n;
  wire g1534_p;
  wire g1534_n;
  wire g1535_p;
  wire g1535_n;
  wire g1536_p;
  wire g1536_n;
  wire g1537_p;
  wire g1537_n;
  wire g1538_p;
  wire g1538_n;
  wire g1539_p;
  wire g1539_n;
  wire g1540_p;
  wire g1540_n;
  wire g1541_p;
  wire g1541_n;
  wire g1542_p;
  wire g1542_n;
  wire g1543_p;
  wire g1543_n;
  wire g1544_p;
  wire g1544_n;
  wire g1545_p;
  wire g1545_n;
  wire g1546_p;
  wire g1546_n;
  wire g1547_p;
  wire g1547_n;
  wire g1548_p;
  wire g1548_n;
  wire g1549_p;
  wire g1549_n;
  wire g1550_p;
  wire g1550_n;
  wire g1551_p;
  wire g1551_n;
  wire g1552_p;
  wire g1552_n;
  wire g1553_p;
  wire g1553_n;
  wire g1554_p;
  wire g1554_n;
  wire g1555_p;
  wire g1555_n;
  wire g1556_p;
  wire g1556_n;
  wire g1557_p;
  wire g1557_n;
  wire g1558_p;
  wire g1558_n;
  wire g1559_p;
  wire g1559_n;
  wire g1560_p;
  wire g1560_n;
  wire g1561_p;
  wire g1561_n;
  wire g1562_p;
  wire g1562_n;
  wire g1563_p;
  wire g1563_n;
  wire g1564_p;
  wire g1564_n;
  wire g1565_p;
  wire g1565_n;
  wire g1566_p;
  wire g1566_n;
  wire g1567_p;
  wire g1567_n;
  wire g1568_p;
  wire g1568_n;
  wire g1569_p;
  wire g1569_n;
  wire g1570_p;
  wire g1570_n;
  wire g1571_p;
  wire g1571_n;
  wire g1572_p;
  wire g1572_n;
  wire g1573_p;
  wire g1573_n;
  wire g1574_p;
  wire g1574_n;
  wire g1575_p;
  wire g1575_n;
  wire g1576_p;
  wire g1576_n;
  wire g1577_p;
  wire g1577_n;
  wire g1578_p;
  wire g1578_n;
  wire g1579_p;
  wire g1579_n;
  wire g1580_p;
  wire g1580_n;
  wire g1581_p;
  wire g1581_n;
  wire g1582_p;
  wire g1582_n;
  wire g1583_p;
  wire g1583_n;
  wire g1584_p;
  wire g1584_n;
  wire g1585_p;
  wire g1585_n;
  wire g1586_p;
  wire g1586_n;
  wire g1587_p;
  wire g1587_n;
  wire g1588_p;
  wire g1588_n;
  wire g1589_p;
  wire g1589_n;
  wire g1590_p;
  wire g1590_n;
  wire g1591_p;
  wire g1591_n;
  wire g1592_p;
  wire g1592_n;
  wire g1593_p;
  wire g1593_n;
  wire g1594_p;
  wire g1594_n;
  wire g1595_p;
  wire g1595_n;
  wire g1596_p;
  wire g1596_n;
  wire g1597_p;
  wire g1597_n;
  wire g1598_p;
  wire g1598_n;
  wire g1599_p;
  wire g1599_n;
  wire g1600_p;
  wire g1600_n;
  wire g1601_p;
  wire g1601_n;
  wire g1602_p;
  wire g1602_n;
  wire g1603_p;
  wire g1603_n;
  wire g1604_p;
  wire g1604_n;
  wire g1605_p;
  wire g1605_n;
  wire g1606_p;
  wire g1606_n;
  wire g1607_p;
  wire g1607_n;
  wire g1608_p;
  wire g1608_n;
  wire g1609_p;
  wire g1609_n;
  wire g1610_p;
  wire g1610_n;
  wire g1611_p;
  wire g1611_n;
  wire g1612_p;
  wire g1612_n;
  wire g1613_p;
  wire g1613_n;
  wire g1614_p;
  wire g1614_n;
  wire g1615_p;
  wire g1615_n;
  wire g1616_p;
  wire g1616_n;
  wire g1617_p;
  wire g1617_n;
  wire g1618_p;
  wire g1618_n;
  wire g1619_p;
  wire g1619_n;
  wire g1620_p;
  wire g1620_n;
  wire g1621_p;
  wire g1621_n;
  wire g1622_p;
  wire g1622_n;
  wire g1623_p;
  wire g1623_n;
  wire g1624_p;
  wire g1624_n;
  wire g1625_p;
  wire g1625_n;
  wire g1626_p;
  wire g1626_n;
  wire g1627_p;
  wire g1627_n;
  wire g1628_p;
  wire g1628_n;
  wire g1629_p;
  wire g1629_n;
  wire g1630_p;
  wire g1630_n;
  wire g1631_p;
  wire g1631_n;
  wire g1632_p;
  wire g1632_n;
  wire g1633_p;
  wire g1633_n;
  wire g1634_p;
  wire g1634_n;
  wire g1635_p;
  wire g1635_n;
  wire g1636_p;
  wire g1636_n;
  wire g1637_p;
  wire g1637_n;
  wire g1638_p;
  wire g1638_n;
  wire g1639_p;
  wire g1639_n;
  wire g1640_p;
  wire g1640_n;
  wire g1641_p;
  wire g1641_n;
  wire g1642_p;
  wire g1642_n;
  wire g1643_p;
  wire g1643_n;
  wire g1644_p;
  wire g1644_n;
  wire g1645_p;
  wire g1645_n;
  wire g1646_p;
  wire g1646_n;
  wire g1647_p;
  wire g1647_n;
  wire g1648_p;
  wire g1648_n;
  wire g1649_p;
  wire g1649_n;
  wire g1650_p;
  wire g1650_n;
  wire g1651_p;
  wire g1651_n;
  wire g1652_p;
  wire g1652_n;
  wire g1653_p;
  wire g1653_n;
  wire g1654_p;
  wire g1654_n;
  wire g1655_p;
  wire g1655_n;
  wire g1656_p;
  wire g1656_n;
  wire g1657_p;
  wire g1657_n;
  wire g1658_p;
  wire g1658_n;
  wire g1659_p;
  wire g1659_n;
  wire g1660_p;
  wire g1660_n;
  wire g1661_p;
  wire g1661_n;
  wire g1662_p;
  wire g1662_n;
  wire g1663_p;
  wire g1663_n;
  wire g1664_p;
  wire g1664_n;
  wire g1665_p;
  wire g1665_n;
  wire g1666_p;
  wire g1666_n;
  wire g1667_p;
  wire g1667_n;
  wire g1668_p;
  wire g1668_n;
  wire g1669_p;
  wire g1669_n;
  wire g1670_p;
  wire g1670_n;
  wire g1671_p;
  wire g1671_n;
  wire g1672_p;
  wire g1672_n;
  wire g1673_p;
  wire g1673_n;
  wire g1674_p;
  wire g1674_n;
  wire g1675_p;
  wire g1675_n;
  wire g1676_p;
  wire g1676_n;
  wire g1677_p;
  wire g1677_n;
  wire g1678_p;
  wire g1678_n;
  wire g1679_p;
  wire g1679_n;
  wire g1680_p;
  wire g1680_n;
  wire g1681_p;
  wire g1681_n;
  wire g1682_p;
  wire g1682_n;
  wire g1683_p;
  wire g1683_n;
  wire g1684_p;
  wire g1684_n;
  wire g1685_p;
  wire g1685_n;
  wire g1686_p;
  wire g1686_n;
  wire g1687_p;
  wire g1687_n;
  wire g1688_p;
  wire g1688_n;
  wire g1689_p;
  wire g1689_n;
  wire g1690_p;
  wire g1690_n;
  wire g1691_p;
  wire g1691_n;
  wire g1692_p;
  wire g1692_n;
  wire g1693_p;
  wire g1693_n;
  wire g1694_p;
  wire g1694_n;
  wire g1695_p;
  wire g1695_n;
  wire n2865_lo_n_spl_;
  wire n2793_lo_n_spl_;
  wire n2793_lo_n_spl_0;
  wire n2793_lo_n_spl_1;
  wire g841_n_spl_;
  wire g841_n_spl_0;
  wire n2565_lo_n_spl_;
  wire n1929_lo_n_spl_;
  wire n2445_lo_n_spl_;
  wire n2049_lo_n_spl_;
  wire n2685_lo_n_spl_;
  wire n2181_lo_n_spl_;
  wire n2325_lo_n_spl_;
  wire n1797_lo_n_spl_;
  wire g849_n_spl_;
  wire g846_n_spl_;
  wire n2877_lo_p_spl_;
  wire n2877_lo_p_spl_0;
  wire n2877_lo_n_spl_;
  wire n2877_lo_n_spl_0;
  wire g856_n_spl_;
  wire g853_n_spl_;
  wire g853_n_spl_0;
  wire g853_n_spl_1;
  wire n2889_lo_p_spl_;
  wire n2889_lo_p_spl_0;
  wire n2889_lo_p_spl_00;
  wire n2889_lo_p_spl_1;
  wire n1235_inv_p_spl_;
  wire n2889_lo_n_spl_;
  wire n2889_lo_n_spl_0;
  wire n2889_lo_n_spl_00;
  wire n2889_lo_n_spl_1;
  wire n1232_inv_p_spl_;
  wire n4711_o2_n_spl_;
  wire g874_n_spl_;
  wire n5477_o2_n_spl_;
  wire g878_n_spl_;
  wire n1521_lo_n_spl_;
  wire G1728_o2_n_spl_;
  wire G1572_o2_p_spl_;
  wire G1728_o2_p_spl_;
  wire G1572_o2_n_spl_;
  wire n5179_o2_p_spl_;
  wire n5179_o2_p_spl_0;
  wire n1761_lo_n_spl_;
  wire G2512_o2_p_spl_;
  wire g1004_p_spl_;
  wire g988_p_spl_;
  wire g895_p_spl_;
  wire g904_p_spl_;
  wire g886_p_spl_;
  wire g1007_n_spl_;
  wire G1008_o2_n_spl_;
  wire G1008_o2_p_spl_;
  wire G1008_o2_p_spl_0;
  wire G1008_o2_p_spl_1;
  wire G636_o2_p_spl_;
  wire G647_o2_p_spl_;
  wire G342_o2_n_spl_;
  wire G354_o2_n_spl_;
  wire G707_o2_p_spl_;
  wire G707_o2_p_spl_0;
  wire G707_o2_p_spl_00;
  wire G707_o2_p_spl_01;
  wire G707_o2_p_spl_1;
  wire G707_o2_p_spl_10;
  wire G707_o2_p_spl_11;
  wire G718_o2_p_spl_;
  wire G718_o2_p_spl_0;
  wire G718_o2_p_spl_00;
  wire G718_o2_p_spl_01;
  wire G718_o2_p_spl_1;
  wire G718_o2_p_spl_10;
  wire G718_o2_p_spl_11;
  wire G405_o2_n_spl_;
  wire G405_o2_n_spl_0;
  wire G405_o2_n_spl_00;
  wire G405_o2_n_spl_01;
  wire G405_o2_n_spl_1;
  wire G405_o2_n_spl_10;
  wire G405_o2_n_spl_11;
  wire G417_o2_n_spl_;
  wire G417_o2_n_spl_0;
  wire G417_o2_n_spl_00;
  wire G417_o2_n_spl_01;
  wire G417_o2_n_spl_1;
  wire G417_o2_n_spl_10;
  wire G417_o2_n_spl_11;
  wire G603_o2_p_spl_;
  wire G603_o2_p_spl_0;
  wire G603_o2_p_spl_00;
  wire G603_o2_p_spl_000;
  wire G603_o2_p_spl_001;
  wire G603_o2_p_spl_01;
  wire G603_o2_p_spl_1;
  wire G603_o2_p_spl_10;
  wire G603_o2_p_spl_11;
  wire G603_o2_n_spl_;
  wire G603_o2_n_spl_0;
  wire G603_o2_n_spl_00;
  wire G603_o2_n_spl_01;
  wire G603_o2_n_spl_1;
  wire G614_o2_p_spl_;
  wire G614_o2_p_spl_0;
  wire G614_o2_p_spl_00;
  wire G614_o2_p_spl_000;
  wire G614_o2_p_spl_001;
  wire G614_o2_p_spl_01;
  wire G614_o2_p_spl_1;
  wire G614_o2_p_spl_10;
  wire G614_o2_p_spl_11;
  wire G614_o2_n_spl_;
  wire G614_o2_n_spl_0;
  wire G614_o2_n_spl_00;
  wire G614_o2_n_spl_01;
  wire G614_o2_n_spl_1;
  wire G301_o2_n_spl_;
  wire G301_o2_n_spl_0;
  wire G301_o2_n_spl_00;
  wire G301_o2_n_spl_000;
  wire G301_o2_n_spl_001;
  wire G301_o2_n_spl_01;
  wire G301_o2_n_spl_1;
  wire G301_o2_n_spl_10;
  wire G301_o2_n_spl_11;
  wire G301_o2_p_spl_;
  wire G301_o2_p_spl_0;
  wire G301_o2_p_spl_00;
  wire G301_o2_p_spl_01;
  wire G301_o2_p_spl_1;
  wire G313_o2_n_spl_;
  wire G313_o2_n_spl_0;
  wire G313_o2_n_spl_00;
  wire G313_o2_n_spl_000;
  wire G313_o2_n_spl_001;
  wire G313_o2_n_spl_01;
  wire G313_o2_n_spl_1;
  wire G313_o2_n_spl_10;
  wire G313_o2_n_spl_11;
  wire G313_o2_p_spl_;
  wire G313_o2_p_spl_0;
  wire G313_o2_p_spl_00;
  wire G313_o2_p_spl_01;
  wire G313_o2_p_spl_1;
  wire G1636_o2_p_spl_;
  wire G1636_o2_p_spl_0;
  wire G1636_o2_p_spl_00;
  wire G1636_o2_p_spl_000;
  wire G1636_o2_p_spl_001;
  wire G1636_o2_p_spl_01;
  wire G1636_o2_p_spl_010;
  wire G1636_o2_p_spl_1;
  wire G1636_o2_p_spl_10;
  wire G1636_o2_p_spl_11;
  wire n3075_lo_buf_o2_n_spl_;
  wire G1636_o2_n_spl_;
  wire G1636_o2_n_spl_0;
  wire G1636_o2_n_spl_00;
  wire G1636_o2_n_spl_000;
  wire G1636_o2_n_spl_001;
  wire G1636_o2_n_spl_01;
  wire G1636_o2_n_spl_010;
  wire G1636_o2_n_spl_1;
  wire G1636_o2_n_spl_10;
  wire G1636_o2_n_spl_11;
  wire n3075_lo_buf_o2_p_spl_;
  wire n3075_lo_buf_o2_p_spl_0;
  wire n3075_lo_buf_o2_p_spl_1;
  wire n2943_lo_buf_o2_n_spl_;
  wire n2943_lo_buf_o2_p_spl_;
  wire n2943_lo_buf_o2_p_spl_0;
  wire n2943_lo_buf_o2_p_spl_1;
  wire G1684_o2_p_spl_;
  wire G1684_o2_p_spl_0;
  wire G1684_o2_p_spl_00;
  wire G1684_o2_p_spl_000;
  wire G1684_o2_p_spl_001;
  wire G1684_o2_p_spl_01;
  wire G1684_o2_p_spl_010;
  wire G1684_o2_p_spl_1;
  wire G1684_o2_p_spl_10;
  wire G1684_o2_p_spl_11;
  wire G1684_o2_n_spl_;
  wire G1684_o2_n_spl_0;
  wire G1684_o2_n_spl_00;
  wire G1684_o2_n_spl_000;
  wire G1684_o2_n_spl_001;
  wire G1684_o2_n_spl_01;
  wire G1684_o2_n_spl_010;
  wire G1684_o2_n_spl_1;
  wire G1684_o2_n_spl_10;
  wire G1684_o2_n_spl_11;
  wire g1097_n_spl_;
  wire g1097_n_spl_0;
  wire g1097_n_spl_1;
  wire g1100_n_spl_;
  wire g1100_n_spl_0;
  wire g1104_n_spl_;
  wire g1113_n_spl_;
  wire g1113_n_spl_0;
  wire g1113_n_spl_00;
  wire g1113_n_spl_1;
  wire g1113_p_spl_;
  wire g1113_p_spl_0;
  wire g1113_p_spl_00;
  wire g1113_p_spl_1;
  wire g1116_n_spl_;
  wire g1116_n_spl_0;
  wire g1116_n_spl_1;
  wire g1116_p_spl_;
  wire g1116_p_spl_0;
  wire g1116_p_spl_1;
  wire g1120_n_spl_;
  wire g1120_n_spl_0;
  wire g1120_p_spl_;
  wire g1120_p_spl_0;
  wire G1336_o2_p_spl_;
  wire G1336_o2_n_spl_;
  wire g1125_n_spl_;
  wire g1125_p_spl_;
  wire G1329_o2_p_spl_;
  wire G1329_o2_p_spl_0;
  wire G1329_o2_n_spl_;
  wire G1329_o2_n_spl_0;
  wire G2414_o2_n_spl_;
  wire G2414_o2_p_spl_;
  wire g1111_n_spl_;
  wire g1159_n_spl_;
  wire g1159_n_spl_0;
  wire g1159_n_spl_1;
  wire g1162_n_spl_;
  wire g1162_n_spl_0;
  wire g1166_n_spl_;
  wire g1175_n_spl_;
  wire g1175_n_spl_0;
  wire g1175_n_spl_00;
  wire g1175_n_spl_1;
  wire g1175_p_spl_;
  wire g1175_p_spl_0;
  wire g1175_p_spl_00;
  wire g1175_p_spl_1;
  wire g1178_n_spl_;
  wire g1178_n_spl_0;
  wire g1178_n_spl_1;
  wire g1178_p_spl_;
  wire g1178_p_spl_0;
  wire g1178_p_spl_1;
  wire g1182_n_spl_;
  wire g1182_n_spl_0;
  wire g1182_p_spl_;
  wire g1182_p_spl_0;
  wire g1187_n_spl_;
  wire g1187_p_spl_;
  wire G2428_o2_n_spl_;
  wire G2428_o2_p_spl_;
  wire g1173_n_spl_;
  wire G1345_o2_p_spl_;
  wire G1342_o2_n_spl_;
  wire G1345_o2_n_spl_;
  wire G1342_o2_p_spl_;
  wire G1351_o2_p_spl_;
  wire G1348_o2_n_spl_;
  wire G1351_o2_n_spl_;
  wire G1348_o2_p_spl_;
  wire n3270_lo_p_spl_;
  wire n3258_lo_n_spl_;
  wire n3270_lo_n_spl_;
  wire n3258_lo_p_spl_;
  wire n2910_lo_buf_o2_n_spl_;
  wire n2922_lo_buf_o2_p_spl_;
  wire n2910_lo_buf_o2_p_spl_;
  wire n2922_lo_buf_o2_n_spl_;
  wire G1049_o2_p_spl_;
  wire G1049_o2_p_spl_0;
  wire G1049_o2_p_spl_1;
  wire n5222_o2_n_spl_;
  wire G1049_o2_n_spl_;
  wire n5222_o2_p_spl_;
  wire n5222_o2_p_spl_0;
  wire n5222_o2_p_spl_1;
  wire n2003_inv_n_spl_;
  wire G1053_o2_n_spl_;
  wire n2003_inv_p_spl_;
  wire n2003_inv_p_spl_0;
  wire G1053_o2_p_spl_;
  wire G1053_o2_p_spl_0;
  wire g1228_n_spl_;
  wire g1228_n_spl_0;
  wire g1231_n_spl_;
  wire g1231_n_spl_0;
  wire n3198_lo_buf_o2_p_spl_;
  wire n3186_lo_buf_o2_n_spl_;
  wire n3198_lo_buf_o2_n_spl_;
  wire n3186_lo_buf_o2_p_spl_;
  wire n3222_lo_buf_o2_p_spl_;
  wire n3210_lo_buf_o2_n_spl_;
  wire n3222_lo_buf_o2_n_spl_;
  wire n3210_lo_buf_o2_p_spl_;
  wire g1258_n_spl_;
  wire g1255_p_spl_;
  wire g1261_p_spl_;
  wire g1255_n_spl_;
  wire g1261_n_spl_;
  wire g1258_p_spl_;
  wire G1079_o2_p_spl_;
  wire G1222_o2_p_spl_;
  wire G1079_o2_n_spl_;
  wire G1222_o2_n_spl_;
  wire G1228_o2_n_spl_;
  wire G1225_o2_p_spl_;
  wire G1228_o2_p_spl_;
  wire G1225_o2_n_spl_;
  wire g1278_p_spl_;
  wire g1275_n_spl_;
  wire g1281_n_spl_;
  wire g1275_p_spl_;
  wire g1281_p_spl_;
  wire g1278_n_spl_;
  wire G1371_o2_p_spl_;
  wire G1368_o2_n_spl_;
  wire G1371_o2_n_spl_;
  wire G1368_o2_p_spl_;
  wire G1537_o2_p_spl_;
  wire G1374_o2_p_spl_;
  wire G1537_o2_n_spl_;
  wire G1374_o2_n_spl_;
  wire g1298_n_spl_;
  wire g1295_p_spl_;
  wire g1301_p_spl_;
  wire g1295_n_spl_;
  wire g1301_n_spl_;
  wire g1298_p_spl_;
  wire n3087_lo_n_spl_;
  wire n2955_lo_n_spl_;
  wire n2991_lo_p_spl_;
  wire n2991_lo_p_spl_0;
  wire n2991_lo_p_spl_1;
  wire n1503_lo_buf_o2_n_spl_;
  wire n1503_lo_buf_o2_n_spl_0;
  wire n1503_lo_buf_o2_n_spl_00;
  wire n1503_lo_buf_o2_n_spl_000;
  wire n1503_lo_buf_o2_n_spl_001;
  wire n1503_lo_buf_o2_n_spl_01;
  wire n1503_lo_buf_o2_n_spl_010;
  wire n1503_lo_buf_o2_n_spl_011;
  wire n1503_lo_buf_o2_n_spl_1;
  wire n1503_lo_buf_o2_n_spl_10;
  wire n1503_lo_buf_o2_n_spl_100;
  wire n1503_lo_buf_o2_n_spl_101;
  wire n1503_lo_buf_o2_n_spl_11;
  wire n1503_lo_buf_o2_n_spl_110;
  wire n1503_lo_buf_o2_n_spl_111;
  wire n3003_lo_p_spl_;
  wire n3003_lo_p_spl_0;
  wire n3003_lo_p_spl_1;
  wire n3063_lo_buf_o2_p_spl_;
  wire n3063_lo_buf_o2_p_spl_0;
  wire n3063_lo_buf_o2_p_spl_00;
  wire n3063_lo_buf_o2_p_spl_01;
  wire n3063_lo_buf_o2_p_spl_1;
  wire g1329_n_spl_;
  wire g1329_n_spl_0;
  wire g1329_n_spl_1;
  wire n3027_lo_n_spl_;
  wire g1329_p_spl_;
  wire g1329_p_spl_0;
  wire g1329_p_spl_00;
  wire g1329_p_spl_01;
  wire g1329_p_spl_1;
  wire g1329_p_spl_10;
  wire g1329_p_spl_11;
  wire n3039_lo_n_spl_;
  wire n3099_lo_buf_o2_p_spl_;
  wire n3099_lo_buf_o2_p_spl_0;
  wire n3099_lo_buf_o2_p_spl_1;
  wire n2967_lo_buf_o2_p_spl_;
  wire n2967_lo_buf_o2_p_spl_0;
  wire n2967_lo_buf_o2_p_spl_1;
  wire n3111_lo_buf_o2_p_spl_;
  wire n3111_lo_buf_o2_p_spl_0;
  wire n3111_lo_buf_o2_p_spl_1;
  wire n2979_lo_buf_o2_p_spl_;
  wire n2979_lo_buf_o2_p_spl_0;
  wire n2979_lo_buf_o2_p_spl_1;
  wire g1020_n_spl_;
  wire g1020_n_spl_0;
  wire g1020_n_spl_00;
  wire g1020_n_spl_1;
  wire G1493_o2_n_spl_;
  wire G1493_o2_n_spl_0;
  wire G1493_o2_n_spl_1;
  wire g1017_n_spl_;
  wire g1017_n_spl_0;
  wire g1017_n_spl_00;
  wire g1017_n_spl_1;
  wire G1498_o2_n_spl_;
  wire G1498_o2_n_spl_0;
  wire G1498_o2_n_spl_1;
  wire g1045_n_spl_;
  wire g1045_n_spl_0;
  wire G1314_o2_n_spl_;
  wire g1056_n_spl_;
  wire g1056_n_spl_0;
  wire g1023_n_spl_;
  wire g1023_n_spl_0;
  wire G1314_o2_p_spl_;
  wire G1021_o2_p_spl_;
  wire G1021_o2_p_spl_0;
  wire G1021_o2_p_spl_00;
  wire G1021_o2_p_spl_01;
  wire G1021_o2_p_spl_1;
  wire G1021_o2_p_spl_10;
  wire G1021_o2_p_spl_11;
  wire G1493_o2_p_spl_;
  wire G1026_o2_p_spl_;
  wire G1026_o2_p_spl_0;
  wire G1026_o2_p_spl_00;
  wire G1026_o2_p_spl_01;
  wire G1026_o2_p_spl_1;
  wire G1026_o2_p_spl_10;
  wire G1498_o2_p_spl_;
  wire n3015_lo_n_spl_;
  wire g1034_n_spl_;
  wire g1034_n_spl_0;
  wire g1034_n_spl_1;
  wire n3150_lo_buf_o2_p_spl_;
  wire n3150_lo_buf_o2_p_spl_0;
  wire n3150_lo_buf_o2_p_spl_00;
  wire n3150_lo_buf_o2_p_spl_000;
  wire n3150_lo_buf_o2_p_spl_001;
  wire n3150_lo_buf_o2_p_spl_01;
  wire n3150_lo_buf_o2_p_spl_1;
  wire n3150_lo_buf_o2_p_spl_10;
  wire n3150_lo_buf_o2_p_spl_11;
  wire n3162_lo_buf_o2_p_spl_;
  wire n3162_lo_buf_o2_p_spl_0;
  wire n3162_lo_buf_o2_p_spl_00;
  wire n3162_lo_buf_o2_p_spl_000;
  wire n3162_lo_buf_o2_p_spl_001;
  wire n3162_lo_buf_o2_p_spl_01;
  wire n3162_lo_buf_o2_p_spl_1;
  wire n3162_lo_buf_o2_p_spl_10;
  wire n3162_lo_buf_o2_p_spl_11;
  wire n3150_lo_buf_o2_n_spl_;
  wire n3150_lo_buf_o2_n_spl_0;
  wire n3150_lo_buf_o2_n_spl_00;
  wire n3150_lo_buf_o2_n_spl_01;
  wire n3150_lo_buf_o2_n_spl_1;
  wire n3162_lo_buf_o2_n_spl_;
  wire n3162_lo_buf_o2_n_spl_0;
  wire n3162_lo_buf_o2_n_spl_00;
  wire n3162_lo_buf_o2_n_spl_01;
  wire n3162_lo_buf_o2_n_spl_1;
  wire n2958_lo_buf_o2_n_spl_;
  wire n2970_lo_buf_o2_p_spl_;
  wire n2958_lo_buf_o2_p_spl_;
  wire n2970_lo_buf_o2_n_spl_;
  wire n2946_lo_buf_o2_p_spl_;
  wire n3282_lo_p_spl_;
  wire n2946_lo_buf_o2_n_spl_;
  wire n3282_lo_n_spl_;
  wire g1453_p_spl_;
  wire g1450_p_spl_;
  wire g1456_n_spl_;
  wire g1456_n_spl_0;
  wire g1456_n_spl_1;
  wire g1453_n_spl_;
  wire n3090_lo_buf_o2_p_spl_;
  wire n3090_lo_buf_o2_p_spl_0;
  wire n3078_lo_buf_o2_n_spl_;
  wire n3090_lo_buf_o2_n_spl_;
  wire n3078_lo_buf_o2_p_spl_;
  wire n3078_lo_buf_o2_p_spl_0;
  wire n3066_lo_buf_o2_p_spl_;
  wire n3294_lo_p_spl_;
  wire n3066_lo_buf_o2_n_spl_;
  wire n3294_lo_n_spl_;
  wire n3114_lo_buf_o2_p_spl_;
  wire n3102_lo_buf_o2_p_spl_;
  wire g1466_p_spl_;
  wire g1463_p_spl_;
  wire g1469_n_spl_;
  wire g1469_n_spl_0;
  wire g1469_n_spl_1;
  wire g1466_n_spl_;
  wire g1450_n_spl_;
  wire g1463_n_spl_;
  wire G1129_o2_p_spl_;
  wire G1132_o2_n_spl_;
  wire G1129_o2_n_spl_;
  wire G1132_o2_p_spl_;
  wire g1480_p_spl_;
  wire g1014_n_spl_;
  wire g1014_n_spl_0;
  wire g1014_n_spl_1;
  wire g1483_n_spl_;
  wire g1483_n_spl_0;
  wire g1483_n_spl_1;
  wire g1480_n_spl_;
  wire g1014_p_spl_;
  wire n1554_lo_p_spl_;
  wire n1554_lo_p_spl_0;
  wire n1554_lo_p_spl_00;
  wire n1554_lo_p_spl_000;
  wire n1554_lo_p_spl_01;
  wire n1554_lo_p_spl_1;
  wire n1554_lo_p_spl_10;
  wire n1554_lo_p_spl_11;
  wire n1554_lo_n_spl_;
  wire n1554_lo_n_spl_0;
  wire n1554_lo_n_spl_00;
  wire n1554_lo_n_spl_000;
  wire n1554_lo_n_spl_01;
  wire n1554_lo_n_spl_1;
  wire n1554_lo_n_spl_10;
  wire n1554_lo_n_spl_11;
  wire G1017_o2_p_spl_;
  wire G1002_o2_p_spl_;
  wire G1002_o2_p_spl_0;
  wire n5554_o2_p_spl_;
  wire n5553_o2_p_spl_;
  wire n1686_lo_p_spl_;
  wire n1686_lo_p_spl_0;
  wire n1686_lo_p_spl_00;
  wire n1686_lo_p_spl_000;
  wire n1686_lo_p_spl_01;
  wire n1686_lo_p_spl_1;
  wire n1686_lo_p_spl_10;
  wire n1686_lo_p_spl_11;
  wire n1686_lo_n_spl_;
  wire n1686_lo_n_spl_0;
  wire n1686_lo_n_spl_00;
  wire n1686_lo_n_spl_01;
  wire n1686_lo_n_spl_1;
  wire n1686_lo_n_spl_10;
  wire n5223_o2_p_spl_;
  wire g1219_n_spl_;
  wire g1157_n_spl_;
  wire g1447_p_spl_;
  wire g1548_n_spl_;
  wire g1436_n_spl_;
  wire g1436_n_spl_0;
  wire n3063_lo_buf_o2_n_spl_;
  wire n2919_lo_buf_o2_n_spl_;
  wire n2919_lo_buf_o2_p_spl_;
  wire n2919_lo_buf_o2_p_spl_0;
  wire n2919_lo_buf_o2_p_spl_1;
  wire g1553_p_spl_;
  wire g1089_n_spl_;
  wire g1089_n_spl_0;
  wire g1089_n_spl_00;
  wire g1089_n_spl_01;
  wire g1089_n_spl_1;
  wire g1089_n_spl_10;
  wire g1557_p_spl_;
  wire g1315_n_spl_;
  wire g1315_n_spl_0;
  wire g1078_p_spl_;
  wire g1078_p_spl_0;
  wire g1078_p_spl_1;
  wire g1358_n_spl_;
  wire g1358_n_spl_0;
  wire g1317_n_spl_;
  wire g1317_n_spl_0;
  wire g1360_n_spl_;
  wire g1360_n_spl_0;
  wire g1319_n_spl_;
  wire g1319_n_spl_0;
  wire g1322_n_spl_;
  wire g1322_n_spl_0;
  wire g1362_n_spl_;
  wire g1362_n_spl_0;
  wire g1324_n_spl_;
  wire g1324_n_spl_0;
  wire g1364_n_spl_;
  wire g1364_n_spl_0;
  wire g1326_n_spl_;
  wire g1326_n_spl_0;
  wire g1370_n_spl_;
  wire g1370_n_spl_0;
  wire g1370_n_spl_00;
  wire g1370_n_spl_01;
  wire g1370_n_spl_1;
  wire g1330_n_spl_;
  wire g1330_n_spl_0;
  wire g1332_n_spl_;
  wire g1332_n_spl_0;
  wire g1366_p_spl_;
  wire g1366_p_spl_0;
  wire g1366_p_spl_00;
  wire g1366_p_spl_01;
  wire g1366_p_spl_1;
  wire g1334_p_spl_;
  wire g1334_p_spl_0;
  wire g1368_p_spl_;
  wire g1368_p_spl_0;
  wire g1368_p_spl_00;
  wire g1368_p_spl_01;
  wire g1368_p_spl_1;
  wire g1336_p_spl_;
  wire g1336_p_spl_0;
  wire g1338_p_spl_;
  wire g1338_p_spl_0;
  wire g1340_p_spl_;
  wire g1340_p_spl_0;
  wire g1374_n_spl_;
  wire g1374_n_spl_0;
  wire g1344_n_spl_;
  wire g1344_n_spl_0;
  wire g1378_n_spl_;
  wire g1378_n_spl_0;
  wire g1348_n_spl_;
  wire g1348_n_spl_0;
  wire g1382_n_spl_;
  wire g1382_n_spl_0;
  wire g1352_n_spl_;
  wire g1352_n_spl_0;
  wire g1386_n_spl_;
  wire g1386_n_spl_0;
  wire g1356_n_spl_;
  wire g1356_n_spl_0;
  wire G663_o2_p_spl_;
  wire G663_o2_p_spl_0;
  wire G663_o2_p_spl_1;
  wire G674_o2_p_spl_;
  wire G674_o2_p_spl_0;
  wire G674_o2_p_spl_1;
  wire G374_o2_n_spl_;
  wire G374_o2_n_spl_0;
  wire G374_o2_n_spl_1;
  wire G386_o2_n_spl_;
  wire G386_o2_n_spl_0;
  wire G386_o2_n_spl_1;
  wire G674_o2_n_spl_;
  wire G663_o2_n_spl_;
  wire G374_o2_p_spl_;
  wire G386_o2_p_spl_;
  wire g1089_p_spl_;
  wire g1092_p_spl_;
  wire g1067_n_spl_;
  wire g1067_n_spl_0;
  wire g1067_n_spl_00;
  wire g1067_n_spl_01;
  wire g1067_n_spl_1;
  wire g1067_p_spl_;
  wire g1095_p_spl_;
  wire n3039_lo_p_spl_;
  wire n3039_lo_p_spl_0;
  wire n3039_lo_p_spl_1;
  wire n2907_lo_p_spl_;
  wire n2907_lo_p_spl_0;
  wire n2907_lo_p_spl_1;
  wire g1412_n_spl_;
  wire g1412_n_spl_0;
  wire g1412_n_spl_00;
  wire g1412_n_spl_1;
  wire n2808_lo_n_spl_;
  wire n2808_lo_n_spl_0;
  wire n2808_lo_n_spl_00;
  wire n2808_lo_n_spl_01;
  wire n2808_lo_n_spl_1;
  wire n2808_lo_n_spl_10;
  wire n2808_lo_n_spl_11;
  wire n2844_lo_p_spl_;
  wire n2844_lo_p_spl_0;
  wire n2844_lo_p_spl_00;
  wire n2844_lo_p_spl_000;
  wire n2844_lo_p_spl_001;
  wire n2844_lo_p_spl_01;
  wire n2844_lo_p_spl_010;
  wire n2844_lo_p_spl_011;
  wire n2844_lo_p_spl_1;
  wire n2844_lo_p_spl_10;
  wire n2844_lo_p_spl_11;
  wire n2844_lo_n_spl_;
  wire n2844_lo_n_spl_0;
  wire n2844_lo_n_spl_00;
  wire n2844_lo_n_spl_01;
  wire n2844_lo_n_spl_1;
  wire n2844_lo_n_spl_10;
  wire n2844_lo_n_spl_11;
  wire n2808_lo_p_spl_;
  wire n2808_lo_p_spl_0;
  wire n2808_lo_p_spl_00;
  wire n2808_lo_p_spl_000;
  wire n2808_lo_p_spl_001;
  wire n2808_lo_p_spl_01;
  wire n2808_lo_p_spl_010;
  wire n2808_lo_p_spl_011;
  wire n2808_lo_p_spl_1;
  wire n2808_lo_p_spl_10;
  wire n2808_lo_p_spl_11;
  wire n2901_lo_n_spl_;
  wire n3057_lo_n_spl_;
  wire n3057_lo_n_spl_0;
  wire g850_n_spl_;
  wire g864_p_spl_;
  wire g867_p_spl_;
  wire g873_p_spl_;
  wire g975_n_spl_;
  wire g1000_p_spl_;
  wire g1013_n_spl_;
  wire n3126_lo_p_spl_;
  wire n3126_lo_p_spl_0;
  wire n3138_lo_p_spl_;
  wire n3138_lo_p_spl_0;
  wire G1039_o2_p_spl_;
  wire G1039_o2_p_spl_0;
  wire n2955_lo_p_spl_;
  wire n3027_lo_p_spl_;
  wire n3087_lo_p_spl_;
  wire n3015_lo_p_spl_;
  wire g1078_n_spl_;
  wire g1078_n_spl_0;
  wire g1078_n_spl_00;
  wire g1078_n_spl_1;
  wire g1222_n_spl_;
  wire g1225_n_spl_;
  wire g1240_n_spl_;
  wire g1249_p_spl_;
  wire g1252_n_spl_;
  wire g1272_p_spl_;
  wire g1292_n_spl_;
  wire g1312_p_spl_;
  wire g1388_p_spl_;
  wire g1388_p_spl_0;
  wire g1390_p_spl_;
  wire g1390_p_spl_0;
  wire g1401_n_spl_;
  wire g1401_n_spl_0;
  wire g1423_n_spl_;
  wire g1423_n_spl_0;
  wire g1425_n_spl_;
  wire g1425_n_spl_0;
  wire g1425_n_spl_00;
  wire g1425_n_spl_01;
  wire g1425_n_spl_1;
  wire n3231_lo_p_spl_;
  wire n3243_lo_p_spl_;
  wire g1550_n_spl_;
  wire g1550_n_spl_0;
  wire g1550_n_spl_00;
  wire g1550_n_spl_1;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  buf

  (
    G42_p,
    G42
  );


  not

  (
    G42_n,
    G42
  );


  buf

  (
    G43_p,
    G43
  );


  not

  (
    G43_n,
    G43
  );


  buf

  (
    G44_p,
    G44
  );


  not

  (
    G44_n,
    G44
  );


  buf

  (
    G45_p,
    G45
  );


  not

  (
    G45_n,
    G45
  );


  buf

  (
    G46_p,
    G46
  );


  not

  (
    G46_n,
    G46
  );


  buf

  (
    G47_p,
    G47
  );


  not

  (
    G47_n,
    G47
  );


  buf

  (
    G48_p,
    G48
  );


  not

  (
    G48_n,
    G48
  );


  buf

  (
    G49_p,
    G49
  );


  not

  (
    G49_n,
    G49
  );


  buf

  (
    G50_p,
    G50
  );


  not

  (
    G50_n,
    G50
  );


  buf

  (
    G51_p,
    G51
  );


  not

  (
    G51_n,
    G51
  );


  buf

  (
    G52_p,
    G52
  );


  not

  (
    G52_n,
    G52
  );


  buf

  (
    G53_p,
    G53
  );


  not

  (
    G53_n,
    G53
  );


  buf

  (
    G54_p,
    G54
  );


  not

  (
    G54_n,
    G54
  );


  buf

  (
    G55_p,
    G55
  );


  not

  (
    G55_n,
    G55
  );


  buf

  (
    G56_p,
    G56
  );


  not

  (
    G56_n,
    G56
  );


  buf

  (
    G57_p,
    G57
  );


  not

  (
    G57_n,
    G57
  );


  buf

  (
    G58_p,
    G58
  );


  not

  (
    G58_n,
    G58
  );


  buf

  (
    G59_p,
    G59
  );


  not

  (
    G59_n,
    G59
  );


  buf

  (
    G60_p,
    G60
  );


  not

  (
    G60_n,
    G60
  );


  buf

  (
    G61_p,
    G61
  );


  not

  (
    G61_n,
    G61
  );


  buf

  (
    G62_p,
    G62
  );


  not

  (
    G62_n,
    G62
  );


  buf

  (
    G63_p,
    G63
  );


  not

  (
    G63_n,
    G63
  );


  buf

  (
    G64_p,
    G64
  );


  not

  (
    G64_n,
    G64
  );


  buf

  (
    G65_p,
    G65
  );


  not

  (
    G65_n,
    G65
  );


  buf

  (
    G66_p,
    G66
  );


  not

  (
    G66_n,
    G66
  );


  buf

  (
    G67_p,
    G67
  );


  not

  (
    G67_n,
    G67
  );


  buf

  (
    G68_p,
    G68
  );


  not

  (
    G68_n,
    G68
  );


  buf

  (
    G69_p,
    G69
  );


  not

  (
    G69_n,
    G69
  );


  buf

  (
    G70_p,
    G70
  );


  not

  (
    G70_n,
    G70
  );


  buf

  (
    G71_p,
    G71
  );


  not

  (
    G71_n,
    G71
  );


  buf

  (
    G72_p,
    G72
  );


  not

  (
    G72_n,
    G72
  );


  buf

  (
    G73_p,
    G73
  );


  not

  (
    G73_n,
    G73
  );


  buf

  (
    G74_p,
    G74
  );


  not

  (
    G74_n,
    G74
  );


  buf

  (
    G75_p,
    G75
  );


  not

  (
    G75_n,
    G75
  );


  buf

  (
    G76_p,
    G76
  );


  not

  (
    G76_n,
    G76
  );


  buf

  (
    G77_p,
    G77
  );


  not

  (
    G77_n,
    G77
  );


  buf

  (
    G78_p,
    G78
  );


  not

  (
    G78_n,
    G78
  );


  buf

  (
    G79_p,
    G79
  );


  not

  (
    G79_n,
    G79
  );


  buf

  (
    G80_p,
    G80
  );


  not

  (
    G80_n,
    G80
  );


  buf

  (
    G81_p,
    G81
  );


  not

  (
    G81_n,
    G81
  );


  buf

  (
    G82_p,
    G82
  );


  not

  (
    G82_n,
    G82
  );


  buf

  (
    G83_p,
    G83
  );


  not

  (
    G83_n,
    G83
  );


  buf

  (
    G84_p,
    G84
  );


  not

  (
    G84_n,
    G84
  );


  buf

  (
    G85_p,
    G85
  );


  not

  (
    G85_n,
    G85
  );


  buf

  (
    G86_p,
    G86
  );


  not

  (
    G86_n,
    G86
  );


  buf

  (
    G87_p,
    G87
  );


  not

  (
    G87_n,
    G87
  );


  buf

  (
    G88_p,
    G88
  );


  not

  (
    G88_n,
    G88
  );


  buf

  (
    G89_p,
    G89
  );


  not

  (
    G89_n,
    G89
  );


  buf

  (
    G90_p,
    G90
  );


  not

  (
    G90_n,
    G90
  );


  buf

  (
    G91_p,
    G91
  );


  not

  (
    G91_n,
    G91
  );


  buf

  (
    G92_p,
    G92
  );


  not

  (
    G92_n,
    G92
  );


  buf

  (
    G93_p,
    G93
  );


  not

  (
    G93_n,
    G93
  );


  buf

  (
    G94_p,
    G94
  );


  not

  (
    G94_n,
    G94
  );


  buf

  (
    G95_p,
    G95
  );


  not

  (
    G95_n,
    G95
  );


  buf

  (
    G96_p,
    G96
  );


  not

  (
    G96_n,
    G96
  );


  buf

  (
    G97_p,
    G97
  );


  not

  (
    G97_n,
    G97
  );


  buf

  (
    G98_p,
    G98
  );


  not

  (
    G98_n,
    G98
  );


  buf

  (
    G99_p,
    G99
  );


  not

  (
    G99_n,
    G99
  );


  buf

  (
    G100_p,
    G100
  );


  not

  (
    G100_n,
    G100
  );


  buf

  (
    G101_p,
    G101
  );


  not

  (
    G101_n,
    G101
  );


  buf

  (
    G102_p,
    G102
  );


  not

  (
    G102_n,
    G102
  );


  buf

  (
    G103_p,
    G103
  );


  not

  (
    G103_n,
    G103
  );


  buf

  (
    G104_p,
    G104
  );


  not

  (
    G104_n,
    G104
  );


  buf

  (
    G105_p,
    G105
  );


  not

  (
    G105_n,
    G105
  );


  buf

  (
    G106_p,
    G106
  );


  not

  (
    G106_n,
    G106
  );


  buf

  (
    G107_p,
    G107
  );


  not

  (
    G107_n,
    G107
  );


  buf

  (
    G108_p,
    G108
  );


  not

  (
    G108_n,
    G108
  );


  buf

  (
    G109_p,
    G109
  );


  not

  (
    G109_n,
    G109
  );


  buf

  (
    G110_p,
    G110
  );


  not

  (
    G110_n,
    G110
  );


  buf

  (
    G111_p,
    G111
  );


  not

  (
    G111_n,
    G111
  );


  buf

  (
    G112_p,
    G112
  );


  not

  (
    G112_n,
    G112
  );


  buf

  (
    G113_p,
    G113
  );


  not

  (
    G113_n,
    G113
  );


  buf

  (
    G114_p,
    G114
  );


  not

  (
    G114_n,
    G114
  );


  buf

  (
    G115_p,
    G115
  );


  not

  (
    G115_n,
    G115
  );


  buf

  (
    G116_p,
    G116
  );


  not

  (
    G116_n,
    G116
  );


  buf

  (
    G117_p,
    G117
  );


  not

  (
    G117_n,
    G117
  );


  buf

  (
    G118_p,
    G118
  );


  not

  (
    G118_n,
    G118
  );


  buf

  (
    G119_p,
    G119
  );


  not

  (
    G119_n,
    G119
  );


  buf

  (
    G120_p,
    G120
  );


  not

  (
    G120_n,
    G120
  );


  buf

  (
    G121_p,
    G121
  );


  not

  (
    G121_n,
    G121
  );


  buf

  (
    G122_p,
    G122
  );


  not

  (
    G122_n,
    G122
  );


  buf

  (
    G123_p,
    G123
  );


  not

  (
    G123_n,
    G123
  );


  buf

  (
    G124_p,
    G124
  );


  not

  (
    G124_n,
    G124
  );


  buf

  (
    G125_p,
    G125
  );


  not

  (
    G125_n,
    G125
  );


  buf

  (
    G126_p,
    G126
  );


  not

  (
    G126_n,
    G126
  );


  buf

  (
    G127_p,
    G127
  );


  not

  (
    G127_n,
    G127
  );


  buf

  (
    G128_p,
    G128
  );


  not

  (
    G128_n,
    G128
  );


  buf

  (
    G129_p,
    G129
  );


  not

  (
    G129_n,
    G129
  );


  buf

  (
    G130_p,
    G130
  );


  not

  (
    G130_n,
    G130
  );


  buf

  (
    G131_p,
    G131
  );


  not

  (
    G131_n,
    G131
  );


  buf

  (
    G132_p,
    G132
  );


  not

  (
    G132_n,
    G132
  );


  buf

  (
    G133_p,
    G133
  );


  not

  (
    G133_n,
    G133
  );


  buf

  (
    G134_p,
    G134
  );


  not

  (
    G134_n,
    G134
  );


  buf

  (
    G135_p,
    G135
  );


  not

  (
    G135_n,
    G135
  );


  buf

  (
    G136_p,
    G136
  );


  not

  (
    G136_n,
    G136
  );


  buf

  (
    G137_p,
    G137
  );


  not

  (
    G137_n,
    G137
  );


  buf

  (
    G138_p,
    G138
  );


  not

  (
    G138_n,
    G138
  );


  buf

  (
    G139_p,
    G139
  );


  not

  (
    G139_n,
    G139
  );


  buf

  (
    G140_p,
    G140
  );


  not

  (
    G140_n,
    G140
  );


  buf

  (
    G141_p,
    G141
  );


  not

  (
    G141_n,
    G141
  );


  buf

  (
    G142_p,
    G142
  );


  not

  (
    G142_n,
    G142
  );


  buf

  (
    G143_p,
    G143
  );


  not

  (
    G143_n,
    G143
  );


  buf

  (
    G144_p,
    G144
  );


  not

  (
    G144_n,
    G144
  );


  buf

  (
    G145_p,
    G145
  );


  not

  (
    G145_n,
    G145
  );


  buf

  (
    G146_p,
    G146
  );


  not

  (
    G146_n,
    G146
  );


  buf

  (
    G147_p,
    G147
  );


  not

  (
    G147_n,
    G147
  );


  buf

  (
    G148_p,
    G148
  );


  not

  (
    G148_n,
    G148
  );


  buf

  (
    G149_p,
    G149
  );


  not

  (
    G149_n,
    G149
  );


  buf

  (
    G150_p,
    G150
  );


  not

  (
    G150_n,
    G150
  );


  buf

  (
    G151_p,
    G151
  );


  not

  (
    G151_n,
    G151
  );


  buf

  (
    G152_p,
    G152
  );


  not

  (
    G152_n,
    G152
  );


  buf

  (
    G153_p,
    G153
  );


  not

  (
    G153_n,
    G153
  );


  buf

  (
    G154_p,
    G154
  );


  not

  (
    G154_n,
    G154
  );


  buf

  (
    G155_p,
    G155
  );


  not

  (
    G155_n,
    G155
  );


  buf

  (
    G156_p,
    G156
  );


  not

  (
    G156_n,
    G156
  );


  buf

  (
    G157_p,
    G157
  );


  not

  (
    G157_n,
    G157
  );


  buf

  (
    n1416_lo_p,
    n1416_lo
  );


  not

  (
    n1416_lo_n,
    n1416_lo
  );


  buf

  (
    n1419_lo_p,
    n1419_lo
  );


  not

  (
    n1419_lo_n,
    n1419_lo
  );


  buf

  (
    n1422_lo_p,
    n1422_lo
  );


  not

  (
    n1422_lo_n,
    n1422_lo
  );


  buf

  (
    n1425_lo_p,
    n1425_lo
  );


  not

  (
    n1425_lo_n,
    n1425_lo
  );


  buf

  (
    n1428_lo_p,
    n1428_lo
  );


  not

  (
    n1428_lo_n,
    n1428_lo
  );


  buf

  (
    n1431_lo_p,
    n1431_lo
  );


  not

  (
    n1431_lo_n,
    n1431_lo
  );


  buf

  (
    n1434_lo_p,
    n1434_lo
  );


  not

  (
    n1434_lo_n,
    n1434_lo
  );


  buf

  (
    n1437_lo_p,
    n1437_lo
  );


  not

  (
    n1437_lo_n,
    n1437_lo
  );


  buf

  (
    n1440_lo_p,
    n1440_lo
  );


  not

  (
    n1440_lo_n,
    n1440_lo
  );


  buf

  (
    n1443_lo_p,
    n1443_lo
  );


  not

  (
    n1443_lo_n,
    n1443_lo
  );


  buf

  (
    n1446_lo_p,
    n1446_lo
  );


  not

  (
    n1446_lo_n,
    n1446_lo
  );


  buf

  (
    n1449_lo_p,
    n1449_lo
  );


  not

  (
    n1449_lo_n,
    n1449_lo
  );


  buf

  (
    n1452_lo_p,
    n1452_lo
  );


  not

  (
    n1452_lo_n,
    n1452_lo
  );


  buf

  (
    n1455_lo_p,
    n1455_lo
  );


  not

  (
    n1455_lo_n,
    n1455_lo
  );


  buf

  (
    n1458_lo_p,
    n1458_lo
  );


  not

  (
    n1458_lo_n,
    n1458_lo
  );


  buf

  (
    n1464_lo_p,
    n1464_lo
  );


  not

  (
    n1464_lo_n,
    n1464_lo
  );


  buf

  (
    n1467_lo_p,
    n1467_lo
  );


  not

  (
    n1467_lo_n,
    n1467_lo
  );


  buf

  (
    n1470_lo_p,
    n1470_lo
  );


  not

  (
    n1470_lo_n,
    n1470_lo
  );


  buf

  (
    n1476_lo_p,
    n1476_lo
  );


  not

  (
    n1476_lo_n,
    n1476_lo
  );


  buf

  (
    n1479_lo_p,
    n1479_lo
  );


  not

  (
    n1479_lo_n,
    n1479_lo
  );


  buf

  (
    n1482_lo_p,
    n1482_lo
  );


  not

  (
    n1482_lo_n,
    n1482_lo
  );


  buf

  (
    n1488_lo_p,
    n1488_lo
  );


  not

  (
    n1488_lo_n,
    n1488_lo
  );


  buf

  (
    n1491_lo_p,
    n1491_lo
  );


  not

  (
    n1491_lo_n,
    n1491_lo
  );


  buf

  (
    n1494_lo_p,
    n1494_lo
  );


  not

  (
    n1494_lo_n,
    n1494_lo
  );


  buf

  (
    n1497_lo_p,
    n1497_lo
  );


  not

  (
    n1497_lo_n,
    n1497_lo
  );


  buf

  (
    n1500_lo_p,
    n1500_lo
  );


  not

  (
    n1500_lo_n,
    n1500_lo
  );


  buf

  (
    n1512_lo_p,
    n1512_lo
  );


  not

  (
    n1512_lo_n,
    n1512_lo
  );


  buf

  (
    n1515_lo_p,
    n1515_lo
  );


  not

  (
    n1515_lo_n,
    n1515_lo
  );


  buf

  (
    n1518_lo_p,
    n1518_lo
  );


  not

  (
    n1518_lo_n,
    n1518_lo
  );


  buf

  (
    n1521_lo_p,
    n1521_lo
  );


  not

  (
    n1521_lo_n,
    n1521_lo
  );


  buf

  (
    n1524_lo_p,
    n1524_lo
  );


  not

  (
    n1524_lo_n,
    n1524_lo
  );


  buf

  (
    n1527_lo_p,
    n1527_lo
  );


  not

  (
    n1527_lo_n,
    n1527_lo
  );


  buf

  (
    n1530_lo_p,
    n1530_lo
  );


  not

  (
    n1530_lo_n,
    n1530_lo
  );


  buf

  (
    n1533_lo_p,
    n1533_lo
  );


  not

  (
    n1533_lo_n,
    n1533_lo
  );


  buf

  (
    n1536_lo_p,
    n1536_lo
  );


  not

  (
    n1536_lo_n,
    n1536_lo
  );


  buf

  (
    n1539_lo_p,
    n1539_lo
  );


  not

  (
    n1539_lo_n,
    n1539_lo
  );


  buf

  (
    n1542_lo_p,
    n1542_lo
  );


  not

  (
    n1542_lo_n,
    n1542_lo
  );


  buf

  (
    n1545_lo_p,
    n1545_lo
  );


  not

  (
    n1545_lo_n,
    n1545_lo
  );


  buf

  (
    n1548_lo_p,
    n1548_lo
  );


  not

  (
    n1548_lo_n,
    n1548_lo
  );


  buf

  (
    n1551_lo_p,
    n1551_lo
  );


  not

  (
    n1551_lo_n,
    n1551_lo
  );


  buf

  (
    n1554_lo_p,
    n1554_lo
  );


  not

  (
    n1554_lo_n,
    n1554_lo
  );


  buf

  (
    n1560_lo_p,
    n1560_lo
  );


  not

  (
    n1560_lo_n,
    n1560_lo
  );


  buf

  (
    n1563_lo_p,
    n1563_lo
  );


  not

  (
    n1563_lo_n,
    n1563_lo
  );


  buf

  (
    n1566_lo_p,
    n1566_lo
  );


  not

  (
    n1566_lo_n,
    n1566_lo
  );


  buf

  (
    n1572_lo_p,
    n1572_lo
  );


  not

  (
    n1572_lo_n,
    n1572_lo
  );


  buf

  (
    n1575_lo_p,
    n1575_lo
  );


  not

  (
    n1575_lo_n,
    n1575_lo
  );


  buf

  (
    n1578_lo_p,
    n1578_lo
  );


  not

  (
    n1578_lo_n,
    n1578_lo
  );


  buf

  (
    n1584_lo_p,
    n1584_lo
  );


  not

  (
    n1584_lo_n,
    n1584_lo
  );


  buf

  (
    n1587_lo_p,
    n1587_lo
  );


  not

  (
    n1587_lo_n,
    n1587_lo
  );


  buf

  (
    n1590_lo_p,
    n1590_lo
  );


  not

  (
    n1590_lo_n,
    n1590_lo
  );


  buf

  (
    n1596_lo_p,
    n1596_lo
  );


  not

  (
    n1596_lo_n,
    n1596_lo
  );


  buf

  (
    n1599_lo_p,
    n1599_lo
  );


  not

  (
    n1599_lo_n,
    n1599_lo
  );


  buf

  (
    n1602_lo_p,
    n1602_lo
  );


  not

  (
    n1602_lo_n,
    n1602_lo
  );


  buf

  (
    n1608_lo_p,
    n1608_lo
  );


  not

  (
    n1608_lo_n,
    n1608_lo
  );


  buf

  (
    n1611_lo_p,
    n1611_lo
  );


  not

  (
    n1611_lo_n,
    n1611_lo
  );


  buf

  (
    n1614_lo_p,
    n1614_lo
  );


  not

  (
    n1614_lo_n,
    n1614_lo
  );


  buf

  (
    n1620_lo_p,
    n1620_lo
  );


  not

  (
    n1620_lo_n,
    n1620_lo
  );


  buf

  (
    n1623_lo_p,
    n1623_lo
  );


  not

  (
    n1623_lo_n,
    n1623_lo
  );


  buf

  (
    n1626_lo_p,
    n1626_lo
  );


  not

  (
    n1626_lo_n,
    n1626_lo
  );


  buf

  (
    n1632_lo_p,
    n1632_lo
  );


  not

  (
    n1632_lo_n,
    n1632_lo
  );


  buf

  (
    n1635_lo_p,
    n1635_lo
  );


  not

  (
    n1635_lo_n,
    n1635_lo
  );


  buf

  (
    n1638_lo_p,
    n1638_lo
  );


  not

  (
    n1638_lo_n,
    n1638_lo
  );


  buf

  (
    n1644_lo_p,
    n1644_lo
  );


  not

  (
    n1644_lo_n,
    n1644_lo
  );


  buf

  (
    n1647_lo_p,
    n1647_lo
  );


  not

  (
    n1647_lo_n,
    n1647_lo
  );


  buf

  (
    n1650_lo_p,
    n1650_lo
  );


  not

  (
    n1650_lo_n,
    n1650_lo
  );


  buf

  (
    n1656_lo_p,
    n1656_lo
  );


  not

  (
    n1656_lo_n,
    n1656_lo
  );


  buf

  (
    n1659_lo_p,
    n1659_lo
  );


  not

  (
    n1659_lo_n,
    n1659_lo
  );


  buf

  (
    n1662_lo_p,
    n1662_lo
  );


  not

  (
    n1662_lo_n,
    n1662_lo
  );


  buf

  (
    n1668_lo_p,
    n1668_lo
  );


  not

  (
    n1668_lo_n,
    n1668_lo
  );


  buf

  (
    n1671_lo_p,
    n1671_lo
  );


  not

  (
    n1671_lo_n,
    n1671_lo
  );


  buf

  (
    n1674_lo_p,
    n1674_lo
  );


  not

  (
    n1674_lo_n,
    n1674_lo
  );


  buf

  (
    n1677_lo_p,
    n1677_lo
  );


  not

  (
    n1677_lo_n,
    n1677_lo
  );


  buf

  (
    n1680_lo_p,
    n1680_lo
  );


  not

  (
    n1680_lo_n,
    n1680_lo
  );


  buf

  (
    n1683_lo_p,
    n1683_lo
  );


  not

  (
    n1683_lo_n,
    n1683_lo
  );


  buf

  (
    n1686_lo_p,
    n1686_lo
  );


  not

  (
    n1686_lo_n,
    n1686_lo
  );


  buf

  (
    n1692_lo_p,
    n1692_lo
  );


  not

  (
    n1692_lo_n,
    n1692_lo
  );


  buf

  (
    n1695_lo_p,
    n1695_lo
  );


  not

  (
    n1695_lo_n,
    n1695_lo
  );


  buf

  (
    n1698_lo_p,
    n1698_lo
  );


  not

  (
    n1698_lo_n,
    n1698_lo
  );


  buf

  (
    n1704_lo_p,
    n1704_lo
  );


  not

  (
    n1704_lo_n,
    n1704_lo
  );


  buf

  (
    n1707_lo_p,
    n1707_lo
  );


  not

  (
    n1707_lo_n,
    n1707_lo
  );


  buf

  (
    n1710_lo_p,
    n1710_lo
  );


  not

  (
    n1710_lo_n,
    n1710_lo
  );


  buf

  (
    n1716_lo_p,
    n1716_lo
  );


  not

  (
    n1716_lo_n,
    n1716_lo
  );


  buf

  (
    n1719_lo_p,
    n1719_lo
  );


  not

  (
    n1719_lo_n,
    n1719_lo
  );


  buf

  (
    n1722_lo_p,
    n1722_lo
  );


  not

  (
    n1722_lo_n,
    n1722_lo
  );


  buf

  (
    n1728_lo_p,
    n1728_lo
  );


  not

  (
    n1728_lo_n,
    n1728_lo
  );


  buf

  (
    n1731_lo_p,
    n1731_lo
  );


  not

  (
    n1731_lo_n,
    n1731_lo
  );


  buf

  (
    n1734_lo_p,
    n1734_lo
  );


  not

  (
    n1734_lo_n,
    n1734_lo
  );


  buf

  (
    n1740_lo_p,
    n1740_lo
  );


  not

  (
    n1740_lo_n,
    n1740_lo
  );


  buf

  (
    n1743_lo_p,
    n1743_lo
  );


  not

  (
    n1743_lo_n,
    n1743_lo
  );


  buf

  (
    n1746_lo_p,
    n1746_lo
  );


  not

  (
    n1746_lo_n,
    n1746_lo
  );


  buf

  (
    n1749_lo_p,
    n1749_lo
  );


  not

  (
    n1749_lo_n,
    n1749_lo
  );


  buf

  (
    n1752_lo_p,
    n1752_lo
  );


  not

  (
    n1752_lo_n,
    n1752_lo
  );


  buf

  (
    n1755_lo_p,
    n1755_lo
  );


  not

  (
    n1755_lo_n,
    n1755_lo
  );


  buf

  (
    n1758_lo_p,
    n1758_lo
  );


  not

  (
    n1758_lo_n,
    n1758_lo
  );


  buf

  (
    n1761_lo_p,
    n1761_lo
  );


  not

  (
    n1761_lo_n,
    n1761_lo
  );


  buf

  (
    n1764_lo_p,
    n1764_lo
  );


  not

  (
    n1764_lo_n,
    n1764_lo
  );


  buf

  (
    n1776_lo_p,
    n1776_lo
  );


  not

  (
    n1776_lo_n,
    n1776_lo
  );


  buf

  (
    n1779_lo_p,
    n1779_lo
  );


  not

  (
    n1779_lo_n,
    n1779_lo
  );


  buf

  (
    n1788_lo_p,
    n1788_lo
  );


  not

  (
    n1788_lo_n,
    n1788_lo
  );


  buf

  (
    n1791_lo_p,
    n1791_lo
  );


  not

  (
    n1791_lo_n,
    n1791_lo
  );


  buf

  (
    n1794_lo_p,
    n1794_lo
  );


  not

  (
    n1794_lo_n,
    n1794_lo
  );


  buf

  (
    n1797_lo_p,
    n1797_lo
  );


  not

  (
    n1797_lo_n,
    n1797_lo
  );


  buf

  (
    n1800_lo_p,
    n1800_lo
  );


  not

  (
    n1800_lo_n,
    n1800_lo
  );


  buf

  (
    n1812_lo_p,
    n1812_lo
  );


  not

  (
    n1812_lo_n,
    n1812_lo
  );


  buf

  (
    n1824_lo_p,
    n1824_lo
  );


  not

  (
    n1824_lo_n,
    n1824_lo
  );


  buf

  (
    n1836_lo_p,
    n1836_lo
  );


  not

  (
    n1836_lo_n,
    n1836_lo
  );


  buf

  (
    n1848_lo_p,
    n1848_lo
  );


  not

  (
    n1848_lo_n,
    n1848_lo
  );


  buf

  (
    n1860_lo_p,
    n1860_lo
  );


  not

  (
    n1860_lo_n,
    n1860_lo
  );


  buf

  (
    n1872_lo_p,
    n1872_lo
  );


  not

  (
    n1872_lo_n,
    n1872_lo
  );


  buf

  (
    n1884_lo_p,
    n1884_lo
  );


  not

  (
    n1884_lo_n,
    n1884_lo
  );


  buf

  (
    n1896_lo_p,
    n1896_lo
  );


  not

  (
    n1896_lo_n,
    n1896_lo
  );


  buf

  (
    n1899_lo_p,
    n1899_lo
  );


  not

  (
    n1899_lo_n,
    n1899_lo
  );


  buf

  (
    n1908_lo_p,
    n1908_lo
  );


  not

  (
    n1908_lo_n,
    n1908_lo
  );


  buf

  (
    n1911_lo_p,
    n1911_lo
  );


  not

  (
    n1911_lo_n,
    n1911_lo
  );


  buf

  (
    n1920_lo_p,
    n1920_lo
  );


  not

  (
    n1920_lo_n,
    n1920_lo
  );


  buf

  (
    n1923_lo_p,
    n1923_lo
  );


  not

  (
    n1923_lo_n,
    n1923_lo
  );


  buf

  (
    n1926_lo_p,
    n1926_lo
  );


  not

  (
    n1926_lo_n,
    n1926_lo
  );


  buf

  (
    n1929_lo_p,
    n1929_lo
  );


  not

  (
    n1929_lo_n,
    n1929_lo
  );


  buf

  (
    n1932_lo_p,
    n1932_lo
  );


  not

  (
    n1932_lo_n,
    n1932_lo
  );


  buf

  (
    n1944_lo_p,
    n1944_lo
  );


  not

  (
    n1944_lo_n,
    n1944_lo
  );


  buf

  (
    n1956_lo_p,
    n1956_lo
  );


  not

  (
    n1956_lo_n,
    n1956_lo
  );


  buf

  (
    n1968_lo_p,
    n1968_lo
  );


  not

  (
    n1968_lo_n,
    n1968_lo
  );


  buf

  (
    n1980_lo_p,
    n1980_lo
  );


  not

  (
    n1980_lo_n,
    n1980_lo
  );


  buf

  (
    n1992_lo_p,
    n1992_lo
  );


  not

  (
    n1992_lo_n,
    n1992_lo
  );


  buf

  (
    n2004_lo_p,
    n2004_lo
  );


  not

  (
    n2004_lo_n,
    n2004_lo
  );


  buf

  (
    n2016_lo_p,
    n2016_lo
  );


  not

  (
    n2016_lo_n,
    n2016_lo
  );


  buf

  (
    n2019_lo_p,
    n2019_lo
  );


  not

  (
    n2019_lo_n,
    n2019_lo
  );


  buf

  (
    n2028_lo_p,
    n2028_lo
  );


  not

  (
    n2028_lo_n,
    n2028_lo
  );


  buf

  (
    n2031_lo_p,
    n2031_lo
  );


  not

  (
    n2031_lo_n,
    n2031_lo
  );


  buf

  (
    n2040_lo_p,
    n2040_lo
  );


  not

  (
    n2040_lo_n,
    n2040_lo
  );


  buf

  (
    n2043_lo_p,
    n2043_lo
  );


  not

  (
    n2043_lo_n,
    n2043_lo
  );


  buf

  (
    n2046_lo_p,
    n2046_lo
  );


  not

  (
    n2046_lo_n,
    n2046_lo
  );


  buf

  (
    n2049_lo_p,
    n2049_lo
  );


  not

  (
    n2049_lo_n,
    n2049_lo
  );


  buf

  (
    n2052_lo_p,
    n2052_lo
  );


  not

  (
    n2052_lo_n,
    n2052_lo
  );


  buf

  (
    n2064_lo_p,
    n2064_lo
  );


  not

  (
    n2064_lo_n,
    n2064_lo
  );


  buf

  (
    n2076_lo_p,
    n2076_lo
  );


  not

  (
    n2076_lo_n,
    n2076_lo
  );


  buf

  (
    n2088_lo_p,
    n2088_lo
  );


  not

  (
    n2088_lo_n,
    n2088_lo
  );


  buf

  (
    n2100_lo_p,
    n2100_lo
  );


  not

  (
    n2100_lo_n,
    n2100_lo
  );


  buf

  (
    n2112_lo_p,
    n2112_lo
  );


  not

  (
    n2112_lo_n,
    n2112_lo
  );


  buf

  (
    n2124_lo_p,
    n2124_lo
  );


  not

  (
    n2124_lo_n,
    n2124_lo
  );


  buf

  (
    n2136_lo_p,
    n2136_lo
  );


  not

  (
    n2136_lo_n,
    n2136_lo
  );


  buf

  (
    n2148_lo_p,
    n2148_lo
  );


  not

  (
    n2148_lo_n,
    n2148_lo
  );


  buf

  (
    n2151_lo_p,
    n2151_lo
  );


  not

  (
    n2151_lo_n,
    n2151_lo
  );


  buf

  (
    n2160_lo_p,
    n2160_lo
  );


  not

  (
    n2160_lo_n,
    n2160_lo
  );


  buf

  (
    n2163_lo_p,
    n2163_lo
  );


  not

  (
    n2163_lo_n,
    n2163_lo
  );


  buf

  (
    n2172_lo_p,
    n2172_lo
  );


  not

  (
    n2172_lo_n,
    n2172_lo
  );


  buf

  (
    n2175_lo_p,
    n2175_lo
  );


  not

  (
    n2175_lo_n,
    n2175_lo
  );


  buf

  (
    n2178_lo_p,
    n2178_lo
  );


  not

  (
    n2178_lo_n,
    n2178_lo
  );


  buf

  (
    n2181_lo_p,
    n2181_lo
  );


  not

  (
    n2181_lo_n,
    n2181_lo
  );


  buf

  (
    n2184_lo_p,
    n2184_lo
  );


  not

  (
    n2184_lo_n,
    n2184_lo
  );


  buf

  (
    n2196_lo_p,
    n2196_lo
  );


  not

  (
    n2196_lo_n,
    n2196_lo
  );


  buf

  (
    n2208_lo_p,
    n2208_lo
  );


  not

  (
    n2208_lo_n,
    n2208_lo
  );


  buf

  (
    n2220_lo_p,
    n2220_lo
  );


  not

  (
    n2220_lo_n,
    n2220_lo
  );


  buf

  (
    n2232_lo_p,
    n2232_lo
  );


  not

  (
    n2232_lo_n,
    n2232_lo
  );


  buf

  (
    n2244_lo_p,
    n2244_lo
  );


  not

  (
    n2244_lo_n,
    n2244_lo
  );


  buf

  (
    n2256_lo_p,
    n2256_lo
  );


  not

  (
    n2256_lo_n,
    n2256_lo
  );


  buf

  (
    n2268_lo_p,
    n2268_lo
  );


  not

  (
    n2268_lo_n,
    n2268_lo
  );


  buf

  (
    n2280_lo_p,
    n2280_lo
  );


  not

  (
    n2280_lo_n,
    n2280_lo
  );


  buf

  (
    n2283_lo_p,
    n2283_lo
  );


  not

  (
    n2283_lo_n,
    n2283_lo
  );


  buf

  (
    n2292_lo_p,
    n2292_lo
  );


  not

  (
    n2292_lo_n,
    n2292_lo
  );


  buf

  (
    n2295_lo_p,
    n2295_lo
  );


  not

  (
    n2295_lo_n,
    n2295_lo
  );


  buf

  (
    n2298_lo_p,
    n2298_lo
  );


  not

  (
    n2298_lo_n,
    n2298_lo
  );


  buf

  (
    n2301_lo_p,
    n2301_lo
  );


  not

  (
    n2301_lo_n,
    n2301_lo
  );


  buf

  (
    n2304_lo_p,
    n2304_lo
  );


  not

  (
    n2304_lo_n,
    n2304_lo
  );


  buf

  (
    n2316_lo_p,
    n2316_lo
  );


  not

  (
    n2316_lo_n,
    n2316_lo
  );


  buf

  (
    n2319_lo_p,
    n2319_lo
  );


  not

  (
    n2319_lo_n,
    n2319_lo
  );


  buf

  (
    n2322_lo_p,
    n2322_lo
  );


  not

  (
    n2322_lo_n,
    n2322_lo
  );


  buf

  (
    n2325_lo_p,
    n2325_lo
  );


  not

  (
    n2325_lo_n,
    n2325_lo
  );


  buf

  (
    n2328_lo_p,
    n2328_lo
  );


  not

  (
    n2328_lo_n,
    n2328_lo
  );


  buf

  (
    n2331_lo_p,
    n2331_lo
  );


  not

  (
    n2331_lo_n,
    n2331_lo
  );


  buf

  (
    n2340_lo_p,
    n2340_lo
  );


  not

  (
    n2340_lo_n,
    n2340_lo
  );


  buf

  (
    n2343_lo_p,
    n2343_lo
  );


  not

  (
    n2343_lo_n,
    n2343_lo
  );


  buf

  (
    n2376_lo_p,
    n2376_lo
  );


  not

  (
    n2376_lo_n,
    n2376_lo
  );


  buf

  (
    n2379_lo_p,
    n2379_lo
  );


  not

  (
    n2379_lo_n,
    n2379_lo
  );


  buf

  (
    n2388_lo_p,
    n2388_lo
  );


  not

  (
    n2388_lo_n,
    n2388_lo
  );


  buf

  (
    n2400_lo_p,
    n2400_lo
  );


  not

  (
    n2400_lo_n,
    n2400_lo
  );


  buf

  (
    n2412_lo_p,
    n2412_lo
  );


  not

  (
    n2412_lo_n,
    n2412_lo
  );


  buf

  (
    n2415_lo_p,
    n2415_lo
  );


  not

  (
    n2415_lo_n,
    n2415_lo
  );


  buf

  (
    n2424_lo_p,
    n2424_lo
  );


  not

  (
    n2424_lo_n,
    n2424_lo
  );


  buf

  (
    n2436_lo_p,
    n2436_lo
  );


  not

  (
    n2436_lo_n,
    n2436_lo
  );


  buf

  (
    n2439_lo_p,
    n2439_lo
  );


  not

  (
    n2439_lo_n,
    n2439_lo
  );


  buf

  (
    n2442_lo_p,
    n2442_lo
  );


  not

  (
    n2442_lo_n,
    n2442_lo
  );


  buf

  (
    n2445_lo_p,
    n2445_lo
  );


  not

  (
    n2445_lo_n,
    n2445_lo
  );


  buf

  (
    n2448_lo_p,
    n2448_lo
  );


  not

  (
    n2448_lo_n,
    n2448_lo
  );


  buf

  (
    n2451_lo_p,
    n2451_lo
  );


  not

  (
    n2451_lo_n,
    n2451_lo
  );


  buf

  (
    n2460_lo_p,
    n2460_lo
  );


  not

  (
    n2460_lo_n,
    n2460_lo
  );


  buf

  (
    n2463_lo_p,
    n2463_lo
  );


  not

  (
    n2463_lo_n,
    n2463_lo
  );


  buf

  (
    n2496_lo_p,
    n2496_lo
  );


  not

  (
    n2496_lo_n,
    n2496_lo
  );


  buf

  (
    n2499_lo_p,
    n2499_lo
  );


  not

  (
    n2499_lo_n,
    n2499_lo
  );


  buf

  (
    n2508_lo_p,
    n2508_lo
  );


  not

  (
    n2508_lo_n,
    n2508_lo
  );


  buf

  (
    n2520_lo_p,
    n2520_lo
  );


  not

  (
    n2520_lo_n,
    n2520_lo
  );


  buf

  (
    n2532_lo_p,
    n2532_lo
  );


  not

  (
    n2532_lo_n,
    n2532_lo
  );


  buf

  (
    n2535_lo_p,
    n2535_lo
  );


  not

  (
    n2535_lo_n,
    n2535_lo
  );


  buf

  (
    n2544_lo_p,
    n2544_lo
  );


  not

  (
    n2544_lo_n,
    n2544_lo
  );


  buf

  (
    n2556_lo_p,
    n2556_lo
  );


  not

  (
    n2556_lo_n,
    n2556_lo
  );


  buf

  (
    n2559_lo_p,
    n2559_lo
  );


  not

  (
    n2559_lo_n,
    n2559_lo
  );


  buf

  (
    n2562_lo_p,
    n2562_lo
  );


  not

  (
    n2562_lo_n,
    n2562_lo
  );


  buf

  (
    n2565_lo_p,
    n2565_lo
  );


  not

  (
    n2565_lo_n,
    n2565_lo
  );


  buf

  (
    n2568_lo_p,
    n2568_lo
  );


  not

  (
    n2568_lo_n,
    n2568_lo
  );


  buf

  (
    n2571_lo_p,
    n2571_lo
  );


  not

  (
    n2571_lo_n,
    n2571_lo
  );


  buf

  (
    n2580_lo_p,
    n2580_lo
  );


  not

  (
    n2580_lo_n,
    n2580_lo
  );


  buf

  (
    n2583_lo_p,
    n2583_lo
  );


  not

  (
    n2583_lo_n,
    n2583_lo
  );


  buf

  (
    n2616_lo_p,
    n2616_lo
  );


  not

  (
    n2616_lo_n,
    n2616_lo
  );


  buf

  (
    n2619_lo_p,
    n2619_lo
  );


  not

  (
    n2619_lo_n,
    n2619_lo
  );


  buf

  (
    n2628_lo_p,
    n2628_lo
  );


  not

  (
    n2628_lo_n,
    n2628_lo
  );


  buf

  (
    n2640_lo_p,
    n2640_lo
  );


  not

  (
    n2640_lo_n,
    n2640_lo
  );


  buf

  (
    n2652_lo_p,
    n2652_lo
  );


  not

  (
    n2652_lo_n,
    n2652_lo
  );


  buf

  (
    n2655_lo_p,
    n2655_lo
  );


  not

  (
    n2655_lo_n,
    n2655_lo
  );


  buf

  (
    n2664_lo_p,
    n2664_lo
  );


  not

  (
    n2664_lo_n,
    n2664_lo
  );


  buf

  (
    n2676_lo_p,
    n2676_lo
  );


  not

  (
    n2676_lo_n,
    n2676_lo
  );


  buf

  (
    n2679_lo_p,
    n2679_lo
  );


  not

  (
    n2679_lo_n,
    n2679_lo
  );


  buf

  (
    n2682_lo_p,
    n2682_lo
  );


  not

  (
    n2682_lo_n,
    n2682_lo
  );


  buf

  (
    n2685_lo_p,
    n2685_lo
  );


  not

  (
    n2685_lo_n,
    n2685_lo
  );


  buf

  (
    n2688_lo_p,
    n2688_lo
  );


  not

  (
    n2688_lo_n,
    n2688_lo
  );


  buf

  (
    n2691_lo_p,
    n2691_lo
  );


  not

  (
    n2691_lo_n,
    n2691_lo
  );


  buf

  (
    n2700_lo_p,
    n2700_lo
  );


  not

  (
    n2700_lo_n,
    n2700_lo
  );


  buf

  (
    n2703_lo_p,
    n2703_lo
  );


  not

  (
    n2703_lo_n,
    n2703_lo
  );


  buf

  (
    n2736_lo_p,
    n2736_lo
  );


  not

  (
    n2736_lo_n,
    n2736_lo
  );


  buf

  (
    n2739_lo_p,
    n2739_lo
  );


  not

  (
    n2739_lo_n,
    n2739_lo
  );


  buf

  (
    n2748_lo_p,
    n2748_lo
  );


  not

  (
    n2748_lo_n,
    n2748_lo
  );


  buf

  (
    n2760_lo_p,
    n2760_lo
  );


  not

  (
    n2760_lo_n,
    n2760_lo
  );


  buf

  (
    n2772_lo_p,
    n2772_lo
  );


  not

  (
    n2772_lo_n,
    n2772_lo
  );


  buf

  (
    n2775_lo_p,
    n2775_lo
  );


  not

  (
    n2775_lo_n,
    n2775_lo
  );


  buf

  (
    n2784_lo_p,
    n2784_lo
  );


  not

  (
    n2784_lo_n,
    n2784_lo
  );


  buf

  (
    n2787_lo_p,
    n2787_lo
  );


  not

  (
    n2787_lo_n,
    n2787_lo
  );


  buf

  (
    n2790_lo_p,
    n2790_lo
  );


  not

  (
    n2790_lo_n,
    n2790_lo
  );


  buf

  (
    n2793_lo_p,
    n2793_lo
  );


  not

  (
    n2793_lo_n,
    n2793_lo
  );


  buf

  (
    n2796_lo_p,
    n2796_lo
  );


  not

  (
    n2796_lo_n,
    n2796_lo
  );


  buf

  (
    n2799_lo_p,
    n2799_lo
  );


  not

  (
    n2799_lo_n,
    n2799_lo
  );


  buf

  (
    n2802_lo_p,
    n2802_lo
  );


  not

  (
    n2802_lo_n,
    n2802_lo
  );


  buf

  (
    n2805_lo_p,
    n2805_lo
  );


  not

  (
    n2805_lo_n,
    n2805_lo
  );


  buf

  (
    n2808_lo_p,
    n2808_lo
  );


  not

  (
    n2808_lo_n,
    n2808_lo
  );


  buf

  (
    n2820_lo_p,
    n2820_lo
  );


  not

  (
    n2820_lo_n,
    n2820_lo
  );


  buf

  (
    n2823_lo_p,
    n2823_lo
  );


  not

  (
    n2823_lo_n,
    n2823_lo
  );


  buf

  (
    n2826_lo_p,
    n2826_lo
  );


  not

  (
    n2826_lo_n,
    n2826_lo
  );


  buf

  (
    n2832_lo_p,
    n2832_lo
  );


  not

  (
    n2832_lo_n,
    n2832_lo
  );


  buf

  (
    n2835_lo_p,
    n2835_lo
  );


  not

  (
    n2835_lo_n,
    n2835_lo
  );


  buf

  (
    n2838_lo_p,
    n2838_lo
  );


  not

  (
    n2838_lo_n,
    n2838_lo
  );


  buf

  (
    n2841_lo_p,
    n2841_lo
  );


  not

  (
    n2841_lo_n,
    n2841_lo
  );


  buf

  (
    n2844_lo_p,
    n2844_lo
  );


  not

  (
    n2844_lo_n,
    n2844_lo
  );


  buf

  (
    n2856_lo_p,
    n2856_lo
  );


  not

  (
    n2856_lo_n,
    n2856_lo
  );


  buf

  (
    n2859_lo_p,
    n2859_lo
  );


  not

  (
    n2859_lo_n,
    n2859_lo
  );


  buf

  (
    n2862_lo_p,
    n2862_lo
  );


  not

  (
    n2862_lo_n,
    n2862_lo
  );


  buf

  (
    n2865_lo_p,
    n2865_lo
  );


  not

  (
    n2865_lo_n,
    n2865_lo
  );


  buf

  (
    n2868_lo_p,
    n2868_lo
  );


  not

  (
    n2868_lo_n,
    n2868_lo
  );


  buf

  (
    n2871_lo_p,
    n2871_lo
  );


  not

  (
    n2871_lo_n,
    n2871_lo
  );


  buf

  (
    n2874_lo_p,
    n2874_lo
  );


  not

  (
    n2874_lo_n,
    n2874_lo
  );


  buf

  (
    n2877_lo_p,
    n2877_lo
  );


  not

  (
    n2877_lo_n,
    n2877_lo
  );


  buf

  (
    n2880_lo_p,
    n2880_lo
  );


  not

  (
    n2880_lo_n,
    n2880_lo
  );


  buf

  (
    n2883_lo_p,
    n2883_lo
  );


  not

  (
    n2883_lo_n,
    n2883_lo
  );


  buf

  (
    n2886_lo_p,
    n2886_lo
  );


  not

  (
    n2886_lo_n,
    n2886_lo
  );


  buf

  (
    n2889_lo_p,
    n2889_lo
  );


  not

  (
    n2889_lo_n,
    n2889_lo
  );


  buf

  (
    n2892_lo_p,
    n2892_lo
  );


  not

  (
    n2892_lo_n,
    n2892_lo
  );


  buf

  (
    n2895_lo_p,
    n2895_lo
  );


  not

  (
    n2895_lo_n,
    n2895_lo
  );


  buf

  (
    n2898_lo_p,
    n2898_lo
  );


  not

  (
    n2898_lo_n,
    n2898_lo
  );


  buf

  (
    n2901_lo_p,
    n2901_lo
  );


  not

  (
    n2901_lo_n,
    n2901_lo
  );


  buf

  (
    n2904_lo_p,
    n2904_lo
  );


  not

  (
    n2904_lo_n,
    n2904_lo
  );


  buf

  (
    n2907_lo_p,
    n2907_lo
  );


  not

  (
    n2907_lo_n,
    n2907_lo
  );


  buf

  (
    n2916_lo_p,
    n2916_lo
  );


  not

  (
    n2916_lo_n,
    n2916_lo
  );


  buf

  (
    n2928_lo_p,
    n2928_lo
  );


  not

  (
    n2928_lo_n,
    n2928_lo
  );


  buf

  (
    n2940_lo_p,
    n2940_lo
  );


  not

  (
    n2940_lo_n,
    n2940_lo
  );


  buf

  (
    n2952_lo_p,
    n2952_lo
  );


  not

  (
    n2952_lo_n,
    n2952_lo
  );


  buf

  (
    n2955_lo_p,
    n2955_lo
  );


  not

  (
    n2955_lo_n,
    n2955_lo
  );


  buf

  (
    n2964_lo_p,
    n2964_lo
  );


  not

  (
    n2964_lo_n,
    n2964_lo
  );


  buf

  (
    n2976_lo_p,
    n2976_lo
  );


  not

  (
    n2976_lo_n,
    n2976_lo
  );


  buf

  (
    n2988_lo_p,
    n2988_lo
  );


  not

  (
    n2988_lo_n,
    n2988_lo
  );


  buf

  (
    n2991_lo_p,
    n2991_lo
  );


  not

  (
    n2991_lo_n,
    n2991_lo
  );


  buf

  (
    n3000_lo_p,
    n3000_lo
  );


  not

  (
    n3000_lo_n,
    n3000_lo
  );


  buf

  (
    n3003_lo_p,
    n3003_lo
  );


  not

  (
    n3003_lo_n,
    n3003_lo
  );


  buf

  (
    n3012_lo_p,
    n3012_lo
  );


  not

  (
    n3012_lo_n,
    n3012_lo
  );


  buf

  (
    n3015_lo_p,
    n3015_lo
  );


  not

  (
    n3015_lo_n,
    n3015_lo
  );


  buf

  (
    n3024_lo_p,
    n3024_lo
  );


  not

  (
    n3024_lo_n,
    n3024_lo
  );


  buf

  (
    n3027_lo_p,
    n3027_lo
  );


  not

  (
    n3027_lo_n,
    n3027_lo
  );


  buf

  (
    n3036_lo_p,
    n3036_lo
  );


  not

  (
    n3036_lo_n,
    n3036_lo
  );


  buf

  (
    n3039_lo_p,
    n3039_lo
  );


  not

  (
    n3039_lo_n,
    n3039_lo
  );


  buf

  (
    n3048_lo_p,
    n3048_lo
  );


  not

  (
    n3048_lo_n,
    n3048_lo
  );


  buf

  (
    n3051_lo_p,
    n3051_lo
  );


  not

  (
    n3051_lo_n,
    n3051_lo
  );


  buf

  (
    n3054_lo_p,
    n3054_lo
  );


  not

  (
    n3054_lo_n,
    n3054_lo
  );


  buf

  (
    n3057_lo_p,
    n3057_lo
  );


  not

  (
    n3057_lo_n,
    n3057_lo
  );


  buf

  (
    n3060_lo_p,
    n3060_lo
  );


  not

  (
    n3060_lo_n,
    n3060_lo
  );


  buf

  (
    n3072_lo_p,
    n3072_lo
  );


  not

  (
    n3072_lo_n,
    n3072_lo
  );


  buf

  (
    n3081_lo_p,
    n3081_lo
  );


  not

  (
    n3081_lo_n,
    n3081_lo
  );


  buf

  (
    n3084_lo_p,
    n3084_lo
  );


  not

  (
    n3084_lo_n,
    n3084_lo
  );


  buf

  (
    n3087_lo_p,
    n3087_lo
  );


  not

  (
    n3087_lo_n,
    n3087_lo
  );


  buf

  (
    n3093_lo_p,
    n3093_lo
  );


  not

  (
    n3093_lo_n,
    n3093_lo
  );


  buf

  (
    n3096_lo_p,
    n3096_lo
  );


  not

  (
    n3096_lo_n,
    n3096_lo
  );


  buf

  (
    n3105_lo_p,
    n3105_lo
  );


  not

  (
    n3105_lo_n,
    n3105_lo
  );


  buf

  (
    n3108_lo_p,
    n3108_lo
  );


  not

  (
    n3108_lo_n,
    n3108_lo
  );


  buf

  (
    n3117_lo_p,
    n3117_lo
  );


  not

  (
    n3117_lo_n,
    n3117_lo
  );


  buf

  (
    n3120_lo_p,
    n3120_lo
  );


  not

  (
    n3120_lo_n,
    n3120_lo
  );


  buf

  (
    n3123_lo_p,
    n3123_lo
  );


  not

  (
    n3123_lo_n,
    n3123_lo
  );


  buf

  (
    n3126_lo_p,
    n3126_lo
  );


  not

  (
    n3126_lo_n,
    n3126_lo
  );


  buf

  (
    n3129_lo_p,
    n3129_lo
  );


  not

  (
    n3129_lo_n,
    n3129_lo
  );


  buf

  (
    n3132_lo_p,
    n3132_lo
  );


  not

  (
    n3132_lo_n,
    n3132_lo
  );


  buf

  (
    n3135_lo_p,
    n3135_lo
  );


  not

  (
    n3135_lo_n,
    n3135_lo
  );


  buf

  (
    n3138_lo_p,
    n3138_lo
  );


  not

  (
    n3138_lo_n,
    n3138_lo
  );


  buf

  (
    n3141_lo_p,
    n3141_lo
  );


  not

  (
    n3141_lo_n,
    n3141_lo
  );


  buf

  (
    n3168_lo_p,
    n3168_lo
  );


  not

  (
    n3168_lo_n,
    n3168_lo
  );


  buf

  (
    n3171_lo_p,
    n3171_lo
  );


  not

  (
    n3171_lo_n,
    n3171_lo
  );


  buf

  (
    n3174_lo_p,
    n3174_lo
  );


  not

  (
    n3174_lo_n,
    n3174_lo
  );


  buf

  (
    n3177_lo_p,
    n3177_lo
  );


  not

  (
    n3177_lo_n,
    n3177_lo
  );


  buf

  (
    n3180_lo_p,
    n3180_lo
  );


  not

  (
    n3180_lo_n,
    n3180_lo
  );


  buf

  (
    n3183_lo_p,
    n3183_lo
  );


  not

  (
    n3183_lo_n,
    n3183_lo
  );


  buf

  (
    n3192_lo_p,
    n3192_lo
  );


  not

  (
    n3192_lo_n,
    n3192_lo
  );


  buf

  (
    n3195_lo_p,
    n3195_lo
  );


  not

  (
    n3195_lo_n,
    n3195_lo
  );


  buf

  (
    n3204_lo_p,
    n3204_lo
  );


  not

  (
    n3204_lo_n,
    n3204_lo
  );


  buf

  (
    n3207_lo_p,
    n3207_lo
  );


  not

  (
    n3207_lo_n,
    n3207_lo
  );


  buf

  (
    n3216_lo_p,
    n3216_lo
  );


  not

  (
    n3216_lo_n,
    n3216_lo
  );


  buf

  (
    n3219_lo_p,
    n3219_lo
  );


  not

  (
    n3219_lo_n,
    n3219_lo
  );


  buf

  (
    n3228_lo_p,
    n3228_lo
  );


  not

  (
    n3228_lo_n,
    n3228_lo
  );


  buf

  (
    n3231_lo_p,
    n3231_lo
  );


  not

  (
    n3231_lo_n,
    n3231_lo
  );


  buf

  (
    n3240_lo_p,
    n3240_lo
  );


  not

  (
    n3240_lo_n,
    n3240_lo
  );


  buf

  (
    n3243_lo_p,
    n3243_lo
  );


  not

  (
    n3243_lo_n,
    n3243_lo
  );


  buf

  (
    n3252_lo_p,
    n3252_lo
  );


  not

  (
    n3252_lo_n,
    n3252_lo
  );


  buf

  (
    n3255_lo_p,
    n3255_lo
  );


  not

  (
    n3255_lo_n,
    n3255_lo
  );


  buf

  (
    n3258_lo_p,
    n3258_lo
  );


  not

  (
    n3258_lo_n,
    n3258_lo
  );


  buf

  (
    n3264_lo_p,
    n3264_lo
  );


  not

  (
    n3264_lo_n,
    n3264_lo
  );


  buf

  (
    n3267_lo_p,
    n3267_lo
  );


  not

  (
    n3267_lo_n,
    n3267_lo
  );


  buf

  (
    n3270_lo_p,
    n3270_lo
  );


  not

  (
    n3270_lo_n,
    n3270_lo
  );


  buf

  (
    n3276_lo_p,
    n3276_lo
  );


  not

  (
    n3276_lo_n,
    n3276_lo
  );


  buf

  (
    n3279_lo_p,
    n3279_lo
  );


  not

  (
    n3279_lo_n,
    n3279_lo
  );


  buf

  (
    n3282_lo_p,
    n3282_lo
  );


  not

  (
    n3282_lo_n,
    n3282_lo
  );


  buf

  (
    n3288_lo_p,
    n3288_lo
  );


  not

  (
    n3288_lo_n,
    n3288_lo
  );


  buf

  (
    n3291_lo_p,
    n3291_lo
  );


  not

  (
    n3291_lo_n,
    n3291_lo
  );


  buf

  (
    n3294_lo_p,
    n3294_lo
  );


  not

  (
    n3294_lo_n,
    n3294_lo
  );


  buf

  (
    n4537_o2_p,
    n4537_o2
  );


  not

  (
    n4537_o2_n,
    n4537_o2
  );


  buf

  (
    n4538_o2_p,
    n4538_o2
  );


  not

  (
    n4538_o2_n,
    n4538_o2
  );


  buf

  (
    n4710_o2_p,
    n4710_o2
  );


  not

  (
    n4710_o2_n,
    n4710_o2
  );


  buf

  (
    n4711_o2_p,
    n4711_o2
  );


  not

  (
    n4711_o2_n,
    n4711_o2
  );


  buf

  (
    n1211_inv_p,
    n1211_inv
  );


  not

  (
    n1211_inv_n,
    n1211_inv
  );


  buf

  (
    n1214_inv_p,
    n1214_inv
  );


  not

  (
    n1214_inv_n,
    n1214_inv
  );


  buf

  (
    n1217_inv_p,
    n1217_inv
  );


  not

  (
    n1217_inv_n,
    n1217_inv
  );


  buf

  (
    n1220_inv_p,
    n1220_inv
  );


  not

  (
    n1220_inv_n,
    n1220_inv
  );


  buf

  (
    n4927_o2_p,
    n4927_o2
  );


  not

  (
    n4927_o2_n,
    n4927_o2
  );


  buf

  (
    n4928_o2_p,
    n4928_o2
  );


  not

  (
    n4928_o2_n,
    n4928_o2
  );


  buf

  (
    n1229_inv_p,
    n1229_inv
  );


  not

  (
    n1229_inv_n,
    n1229_inv
  );


  buf

  (
    n1232_inv_p,
    n1232_inv
  );


  not

  (
    n1232_inv_n,
    n1232_inv
  );


  buf

  (
    n1235_inv_p,
    n1235_inv
  );


  not

  (
    n1235_inv_n,
    n1235_inv
  );


  buf

  (
    n5178_o2_p,
    n5178_o2
  );


  not

  (
    n5178_o2_n,
    n5178_o2
  );


  buf

  (
    n5179_o2_p,
    n5179_o2
  );


  not

  (
    n5179_o2_n,
    n5179_o2
  );


  buf

  (
    n5477_o2_p,
    n5477_o2
  );


  not

  (
    n5477_o2_n,
    n5477_o2
  );


  buf

  (
    n5478_o2_p,
    n5478_o2
  );


  not

  (
    n5478_o2_n,
    n5478_o2
  );


  buf

  (
    n5479_o2_p,
    n5479_o2
  );


  not

  (
    n5479_o2_n,
    n5479_o2
  );


  buf

  (
    n5222_o2_p,
    n5222_o2
  );


  not

  (
    n5222_o2_n,
    n5222_o2
  );


  buf

  (
    n5223_o2_p,
    n5223_o2
  );


  not

  (
    n5223_o2_n,
    n5223_o2
  );


  buf

  (
    n5553_o2_p,
    n5553_o2
  );


  not

  (
    n5553_o2_n,
    n5553_o2
  );


  buf

  (
    n5554_o2_p,
    n5554_o2
  );


  not

  (
    n5554_o2_n,
    n5554_o2
  );


  buf

  (
    G491_o2_p,
    G491_o2
  );


  not

  (
    G491_o2_n,
    G491_o2
  );


  buf

  (
    n2922_lo_buf_o2_p,
    n2922_lo_buf_o2
  );


  not

  (
    n2922_lo_buf_o2_n,
    n2922_lo_buf_o2
  );


  buf

  (
    n2946_lo_buf_o2_p,
    n2946_lo_buf_o2
  );


  not

  (
    n2946_lo_buf_o2_n,
    n2946_lo_buf_o2
  );


  buf

  (
    n2970_lo_buf_o2_p,
    n2970_lo_buf_o2
  );


  not

  (
    n2970_lo_buf_o2_n,
    n2970_lo_buf_o2
  );


  buf

  (
    n2982_lo_buf_o2_p,
    n2982_lo_buf_o2
  );


  not

  (
    n2982_lo_buf_o2_n,
    n2982_lo_buf_o2
  );


  buf

  (
    n3066_lo_buf_o2_p,
    n3066_lo_buf_o2
  );


  not

  (
    n3066_lo_buf_o2_n,
    n3066_lo_buf_o2
  );


  buf

  (
    n3078_lo_buf_o2_p,
    n3078_lo_buf_o2
  );


  not

  (
    n3078_lo_buf_o2_n,
    n3078_lo_buf_o2
  );


  buf

  (
    n3102_lo_buf_o2_p,
    n3102_lo_buf_o2
  );


  not

  (
    n3102_lo_buf_o2_n,
    n3102_lo_buf_o2
  );


  buf

  (
    n3114_lo_buf_o2_p,
    n3114_lo_buf_o2
  );


  not

  (
    n3114_lo_buf_o2_n,
    n3114_lo_buf_o2
  );


  buf

  (
    G1321_o2_p,
    G1321_o2
  );


  not

  (
    G1321_o2_n,
    G1321_o2
  );


  buf

  (
    G1033_o2_p,
    G1033_o2
  );


  not

  (
    G1033_o2_n,
    G1033_o2
  );


  buf

  (
    G1030_o2_p,
    G1030_o2
  );


  not

  (
    G1030_o2_n,
    G1030_o2
  );


  buf

  (
    G1072_o2_p,
    G1072_o2
  );


  not

  (
    G1072_o2_n,
    G1072_o2
  );


  buf

  (
    n1304_inv_p,
    n1304_inv
  );


  not

  (
    n1304_inv_n,
    n1304_inv
  );


  buf

  (
    n1307_inv_p,
    n1307_inv
  );


  not

  (
    n1307_inv_n,
    n1307_inv
  );


  buf

  (
    n2958_lo_buf_o2_p,
    n2958_lo_buf_o2
  );


  not

  (
    n2958_lo_buf_o2_n,
    n2958_lo_buf_o2
  );


  buf

  (
    n2994_lo_buf_o2_p,
    n2994_lo_buf_o2
  );


  not

  (
    n2994_lo_buf_o2_n,
    n2994_lo_buf_o2
  );


  buf

  (
    n3006_lo_buf_o2_p,
    n3006_lo_buf_o2
  );


  not

  (
    n3006_lo_buf_o2_n,
    n3006_lo_buf_o2
  );


  buf

  (
    n3030_lo_buf_o2_p,
    n3030_lo_buf_o2
  );


  not

  (
    n3030_lo_buf_o2_n,
    n3030_lo_buf_o2
  );


  buf

  (
    n3042_lo_buf_o2_p,
    n3042_lo_buf_o2
  );


  not

  (
    n3042_lo_buf_o2_n,
    n3042_lo_buf_o2
  );


  buf

  (
    n3090_lo_buf_o2_p,
    n3090_lo_buf_o2
  );


  not

  (
    n3090_lo_buf_o2_n,
    n3090_lo_buf_o2
  );


  buf

  (
    n1328_inv_p,
    n1328_inv
  );


  not

  (
    n1328_inv_n,
    n1328_inv
  );


  buf

  (
    n1331_inv_p,
    n1331_inv
  );


  not

  (
    n1331_inv_n,
    n1331_inv
  );


  buf

  (
    n1334_inv_p,
    n1334_inv
  );


  not

  (
    n1334_inv_n,
    n1334_inv
  );


  buf

  (
    n1337_inv_p,
    n1337_inv
  );


  not

  (
    n1337_inv_n,
    n1337_inv
  );


  buf

  (
    n1340_inv_p,
    n1340_inv
  );


  not

  (
    n1340_inv_n,
    n1340_inv
  );


  buf

  (
    n1343_inv_p,
    n1343_inv
  );


  not

  (
    n1343_inv_n,
    n1343_inv
  );


  buf

  (
    n1346_inv_p,
    n1346_inv
  );


  not

  (
    n1346_inv_n,
    n1346_inv
  );


  buf

  (
    n1349_inv_p,
    n1349_inv
  );


  not

  (
    n1349_inv_n,
    n1349_inv
  );


  buf

  (
    G1036_o2_p,
    G1036_o2
  );


  not

  (
    G1036_o2_n,
    G1036_o2
  );


  buf

  (
    G1062_o2_p,
    G1062_o2
  );


  not

  (
    G1062_o2_n,
    G1062_o2
  );


  buf

  (
    G1067_o2_p,
    G1067_o2
  );


  not

  (
    G1067_o2_n,
    G1067_o2
  );


  buf

  (
    G1014_o2_p,
    G1014_o2
  );


  not

  (
    G1014_o2_n,
    G1014_o2
  );


  buf

  (
    n1364_inv_p,
    n1364_inv
  );


  not

  (
    n1364_inv_n,
    n1364_inv
  );


  buf

  (
    n1367_inv_p,
    n1367_inv
  );


  not

  (
    n1367_inv_n,
    n1367_inv
  );


  buf

  (
    n3018_lo_buf_o2_p,
    n3018_lo_buf_o2
  );


  not

  (
    n3018_lo_buf_o2_n,
    n3018_lo_buf_o2
  );


  buf

  (
    G766_o2_p,
    G766_o2
  );


  not

  (
    G766_o2_n,
    G766_o2
  );


  buf

  (
    n1376_inv_p,
    n1376_inv
  );


  not

  (
    n1376_inv_n,
    n1376_inv
  );


  buf

  (
    n1379_inv_p,
    n1379_inv
  );


  not

  (
    n1379_inv_n,
    n1379_inv
  );


  buf

  (
    n1382_inv_p,
    n1382_inv
  );


  not

  (
    n1382_inv_n,
    n1382_inv
  );


  buf

  (
    n1385_inv_p,
    n1385_inv
  );


  not

  (
    n1385_inv_n,
    n1385_inv
  );


  buf

  (
    n1388_inv_p,
    n1388_inv
  );


  not

  (
    n1388_inv_n,
    n1388_inv
  );


  buf

  (
    n1391_inv_p,
    n1391_inv
  );


  not

  (
    n1391_inv_n,
    n1391_inv
  );


  buf

  (
    G1017_o2_p,
    G1017_o2
  );


  not

  (
    G1017_o2_n,
    G1017_o2
  );


  buf

  (
    G1008_o2_p,
    G1008_o2
  );


  not

  (
    G1008_o2_n,
    G1008_o2
  );


  buf

  (
    n1400_inv_p,
    n1400_inv
  );


  not

  (
    n1400_inv_n,
    n1400_inv
  );


  buf

  (
    n1403_inv_p,
    n1403_inv
  );


  not

  (
    n1403_inv_n,
    n1403_inv
  );


  buf

  (
    n2910_lo_buf_o2_p,
    n2910_lo_buf_o2
  );


  not

  (
    n2910_lo_buf_o2_n,
    n2910_lo_buf_o2
  );


  buf

  (
    n1409_inv_p,
    n1409_inv
  );


  not

  (
    n1409_inv_n,
    n1409_inv
  );


  buf

  (
    G2138_o2_p,
    G2138_o2
  );


  not

  (
    G2138_o2_n,
    G2138_o2
  );


  buf

  (
    G2147_o2_p,
    G2147_o2
  );


  not

  (
    G2147_o2_n,
    G2147_o2
  );


  buf

  (
    n1418_inv_p,
    n1418_inv
  );


  not

  (
    n1418_inv_n,
    n1418_inv
  );


  buf

  (
    G1137_o2_p,
    G1137_o2
  );


  not

  (
    G1137_o2_n,
    G1137_o2
  );


  buf

  (
    G1329_o2_p,
    G1329_o2
  );


  not

  (
    G1329_o2_n,
    G1329_o2
  );


  buf

  (
    G374_o2_p,
    G374_o2
  );


  not

  (
    G374_o2_n,
    G374_o2
  );


  buf

  (
    G386_o2_p,
    G386_o2
  );


  not

  (
    G386_o2_n,
    G386_o2
  );


  buf

  (
    G663_o2_p,
    G663_o2
  );


  not

  (
    G663_o2_n,
    G663_o2
  );


  buf

  (
    G674_o2_p,
    G674_o2
  );


  not

  (
    G674_o2_n,
    G674_o2
  );


  buf

  (
    G578_o2_p,
    G578_o2
  );


  not

  (
    G578_o2_n,
    G578_o2
  );


  buf

  (
    G575_o2_p,
    G575_o2
  );


  not

  (
    G575_o2_n,
    G575_o2
  );


  buf

  (
    G2505_o2_p,
    G2505_o2
  );


  not

  (
    G2505_o2_n,
    G2505_o2
  );


  buf

  (
    n1448_inv_p,
    n1448_inv
  );


  not

  (
    n1448_inv_n,
    n1448_inv
  );


  buf

  (
    G987_o2_p,
    G987_o2
  );


  not

  (
    G987_o2_n,
    G987_o2
  );


  buf

  (
    G984_o2_p,
    G984_o2
  );


  not

  (
    G984_o2_n,
    G984_o2
  );


  buf

  (
    G1862_o2_p,
    G1862_o2
  );


  not

  (
    G1862_o2_n,
    G1862_o2
  );


  buf

  (
    G1859_o2_p,
    G1859_o2
  );


  not

  (
    G1859_o2_n,
    G1859_o2
  );


  buf

  (
    G1260_o2_p,
    G1260_o2
  );


  not

  (
    G1260_o2_n,
    G1260_o2
  );


  buf

  (
    G1865_o2_p,
    G1865_o2
  );


  not

  (
    G1865_o2_n,
    G1865_o2
  );


  buf

  (
    G2073_o2_p,
    G2073_o2
  );


  not

  (
    G2073_o2_n,
    G2073_o2
  );


  buf

  (
    G1402_o2_p,
    G1402_o2
  );


  not

  (
    G1402_o2_n,
    G1402_o2
  );


  buf

  (
    G2048_o2_p,
    G2048_o2
  );


  not

  (
    G2048_o2_n,
    G2048_o2
  );


  buf

  (
    G2276_o2_p,
    G2276_o2
  );


  not

  (
    G2276_o2_n,
    G2276_o2
  );


  buf

  (
    n1481_inv_p,
    n1481_inv
  );


  not

  (
    n1481_inv_n,
    n1481_inv
  );


  buf

  (
    G2141_o2_p,
    G2141_o2
  );


  not

  (
    G2141_o2_n,
    G2141_o2
  );


  buf

  (
    G2008_o2_p,
    G2008_o2
  );


  not

  (
    G2008_o2_n,
    G2008_o2
  );


  buf

  (
    G2011_o2_p,
    G2011_o2
  );


  not

  (
    G2011_o2_n,
    G2011_o2
  );


  buf

  (
    G2150_o2_p,
    G2150_o2
  );


  not

  (
    G2150_o2_n,
    G2150_o2
  );


  buf

  (
    G2026_o2_p,
    G2026_o2
  );


  not

  (
    G2026_o2_n,
    G2026_o2
  );


  buf

  (
    G2029_o2_p,
    G2029_o2
  );


  not

  (
    G2029_o2_n,
    G2029_o2
  );


  buf

  (
    G2023_o2_p,
    G2023_o2
  );


  not

  (
    G2023_o2_n,
    G2023_o2
  );


  buf

  (
    G2041_o2_p,
    G2041_o2
  );


  not

  (
    G2041_o2_n,
    G2041_o2
  );


  buf

  (
    G2017_o2_p,
    G2017_o2
  );


  not

  (
    G2017_o2_n,
    G2017_o2
  );


  buf

  (
    G2020_o2_p,
    G2020_o2
  );


  not

  (
    G2020_o2_n,
    G2020_o2
  );


  buf

  (
    G2035_o2_p,
    G2035_o2
  );


  not

  (
    G2035_o2_n,
    G2035_o2
  );


  buf

  (
    G2038_o2_p,
    G2038_o2
  );


  not

  (
    G2038_o2_n,
    G2038_o2
  );


  buf

  (
    G2228_o2_p,
    G2228_o2
  );


  not

  (
    G2228_o2_n,
    G2228_o2
  );


  buf

  (
    G2231_o2_p,
    G2231_o2
  );


  not

  (
    G2231_o2_n,
    G2231_o2
  );


  buf

  (
    G2234_o2_p,
    G2234_o2
  );


  not

  (
    G2234_o2_n,
    G2234_o2
  );


  buf

  (
    G2237_o2_p,
    G2237_o2
  );


  not

  (
    G2237_o2_n,
    G2237_o2
  );


  buf

  (
    G1904_o2_p,
    G1904_o2
  );


  not

  (
    G1904_o2_n,
    G1904_o2
  );


  buf

  (
    G1907_o2_p,
    G1907_o2
  );


  not

  (
    G1907_o2_n,
    G1907_o2
  );


  buf

  (
    G1928_o2_p,
    G1928_o2
  );


  not

  (
    G1928_o2_n,
    G1928_o2
  );


  buf

  (
    G1931_o2_p,
    G1931_o2
  );


  not

  (
    G1931_o2_n,
    G1931_o2
  );


  buf

  (
    G1893_o2_p,
    G1893_o2
  );


  not

  (
    G1893_o2_n,
    G1893_o2
  );


  buf

  (
    G1896_o2_p,
    G1896_o2
  );


  not

  (
    G1896_o2_n,
    G1896_o2
  );


  buf

  (
    G1899_o2_p,
    G1899_o2
  );


  not

  (
    G1899_o2_n,
    G1899_o2
  );


  buf

  (
    G1937_o2_p,
    G1937_o2
  );


  not

  (
    G1937_o2_n,
    G1937_o2
  );


  buf

  (
    G1940_o2_p,
    G1940_o2
  );


  not

  (
    G1940_o2_n,
    G1940_o2
  );


  buf

  (
    G1943_o2_p,
    G1943_o2
  );


  not

  (
    G1943_o2_n,
    G1943_o2
  );


  buf

  (
    G1336_o2_p,
    G1336_o2
  );


  not

  (
    G1336_o2_n,
    G1336_o2
  );


  buf

  (
    G1996_o2_p,
    G1996_o2
  );


  not

  (
    G1996_o2_n,
    G1996_o2
  );


  buf

  (
    G1999_o2_p,
    G1999_o2
  );


  not

  (
    G1999_o2_n,
    G1999_o2
  );


  buf

  (
    G2002_o2_p,
    G2002_o2
  );


  not

  (
    G2002_o2_n,
    G2002_o2
  );


  buf

  (
    G2005_o2_p,
    G2005_o2
  );


  not

  (
    G2005_o2_n,
    G2005_o2
  );


  buf

  (
    G2014_o2_p,
    G2014_o2
  );


  not

  (
    G2014_o2_n,
    G2014_o2
  );


  buf

  (
    G2032_o2_p,
    G2032_o2
  );


  not

  (
    G2032_o2_n,
    G2032_o2
  );


  buf

  (
    G1076_o2_p,
    G1076_o2
  );


  not

  (
    G1076_o2_n,
    G1076_o2
  );


  buf

  (
    G1002_o2_p,
    G1002_o2
  );


  not

  (
    G1002_o2_n,
    G1002_o2
  );


  buf

  (
    G998_o2_p,
    G998_o2
  );


  not

  (
    G998_o2_n,
    G998_o2
  );


  buf

  (
    G1890_o2_p,
    G1890_o2
  );


  not

  (
    G1890_o2_n,
    G1890_o2
  );


  buf

  (
    G1934_o2_p,
    G1934_o2
  );


  not

  (
    G1934_o2_n,
    G1934_o2
  );


  buf

  (
    G1044_o2_p,
    G1044_o2
  );


  not

  (
    G1044_o2_n,
    G1044_o2
  );


  buf

  (
    G1039_o2_p,
    G1039_o2
  );


  not

  (
    G1039_o2_n,
    G1039_o2
  );


  buf

  (
    n1770_lo_buf_o2_p,
    n1770_lo_buf_o2
  );


  not

  (
    n1770_lo_buf_o2_n,
    n1770_lo_buf_o2
  );


  buf

  (
    G342_o2_p,
    G342_o2
  );


  not

  (
    G342_o2_n,
    G342_o2
  );


  buf

  (
    G354_o2_p,
    G354_o2
  );


  not

  (
    G354_o2_n,
    G354_o2
  );


  buf

  (
    G1193_o2_p,
    G1193_o2
  );


  not

  (
    G1193_o2_n,
    G1193_o2
  );


  buf

  (
    n3234_lo_buf_o2_p,
    n3234_lo_buf_o2
  );


  not

  (
    n3234_lo_buf_o2_n,
    n3234_lo_buf_o2
  );


  buf

  (
    n3246_lo_buf_o2_p,
    n3246_lo_buf_o2
  );


  not

  (
    n3246_lo_buf_o2_n,
    n3246_lo_buf_o2
  );


  buf

  (
    G783_o2_p,
    G783_o2
  );


  not

  (
    G783_o2_n,
    G783_o2
  );


  buf

  (
    G786_o2_p,
    G786_o2
  );


  not

  (
    G786_o2_n,
    G786_o2
  );


  buf

  (
    G792_o2_p,
    G792_o2
  );


  not

  (
    G792_o2_n,
    G792_o2
  );


  buf

  (
    G795_o2_p,
    G795_o2
  );


  not

  (
    G795_o2_n,
    G795_o2
  );


  buf

  (
    G815_o2_p,
    G815_o2
  );


  not

  (
    G815_o2_n,
    G815_o2
  );


  buf

  (
    G818_o2_p,
    G818_o2
  );


  not

  (
    G818_o2_n,
    G818_o2
  );


  buf

  (
    G824_o2_p,
    G824_o2
  );


  not

  (
    G824_o2_n,
    G824_o2
  );


  buf

  (
    G827_o2_p,
    G827_o2
  );


  not

  (
    G827_o2_n,
    G827_o2
  );


  buf

  (
    G789_o2_p,
    G789_o2
  );


  not

  (
    G789_o2_n,
    G789_o2
  );


  buf

  (
    G798_o2_p,
    G798_o2
  );


  not

  (
    G798_o2_n,
    G798_o2
  );


  buf

  (
    G801_o2_p,
    G801_o2
  );


  not

  (
    G801_o2_n,
    G801_o2
  );


  buf

  (
    G807_o2_p,
    G807_o2
  );


  not

  (
    G807_o2_n,
    G807_o2
  );


  buf

  (
    G812_o2_p,
    G812_o2
  );


  not

  (
    G812_o2_n,
    G812_o2
  );


  buf

  (
    G821_o2_p,
    G821_o2
  );


  not

  (
    G821_o2_n,
    G821_o2
  );


  buf

  (
    G804_o2_p,
    G804_o2
  );


  not

  (
    G804_o2_n,
    G804_o2
  );


  buf

  (
    G780_o2_p,
    G780_o2
  );


  not

  (
    G780_o2_n,
    G780_o2
  );


  buf

  (
    G1231_o2_p,
    G1231_o2
  );


  not

  (
    G1231_o2_n,
    G1231_o2
  );


  buf

  (
    G1572_o2_p,
    G1572_o2
  );


  not

  (
    G1572_o2_n,
    G1572_o2
  );


  buf

  (
    G1377_o2_p,
    G1377_o2
  );


  not

  (
    G1377_o2_n,
    G1377_o2
  );


  buf

  (
    G1253_o2_p,
    G1253_o2
  );


  not

  (
    G1253_o2_n,
    G1253_o2
  );


  buf

  (
    G1359_o2_p,
    G1359_o2
  );


  not

  (
    G1359_o2_n,
    G1359_o2
  );


  buf

  (
    G1258_o2_p,
    G1258_o2
  );


  not

  (
    G1258_o2_n,
    G1258_o2
  );


  buf

  (
    G1367_o2_p,
    G1367_o2
  );


  not

  (
    G1367_o2_n,
    G1367_o2
  );


  buf

  (
    G1358_o2_p,
    G1358_o2
  );


  not

  (
    G1358_o2_n,
    G1358_o2
  );


  buf

  (
    G1366_o2_p,
    G1366_o2
  );


  not

  (
    G1366_o2_n,
    G1366_o2
  );


  buf

  (
    G2057_o2_p,
    G2057_o2
  );


  not

  (
    G2057_o2_n,
    G2057_o2
  );


  buf

  (
    G2117_o2_p,
    G2117_o2
  );


  not

  (
    G2117_o2_n,
    G2117_o2
  );


  buf

  (
    G2118_o2_p,
    G2118_o2
  );


  not

  (
    G2118_o2_n,
    G2118_o2
  );


  buf

  (
    G1254_o2_p,
    G1254_o2
  );


  not

  (
    G1254_o2_n,
    G1254_o2
  );


  buf

  (
    G1259_o2_p,
    G1259_o2
  );


  not

  (
    G1259_o2_n,
    G1259_o2
  );


  buf

  (
    G2058_o2_p,
    G2058_o2
  );


  not

  (
    G2058_o2_n,
    G2058_o2
  );


  buf

  (
    G405_o2_p,
    G405_o2
  );


  not

  (
    G405_o2_n,
    G405_o2
  );


  buf

  (
    G417_o2_p,
    G417_o2
  );


  not

  (
    G417_o2_n,
    G417_o2
  );


  buf

  (
    G1269_o2_p,
    G1269_o2
  );


  not

  (
    G1269_o2_n,
    G1269_o2
  );


  buf

  (
    G1275_o2_p,
    G1275_o2
  );


  not

  (
    G1275_o2_n,
    G1275_o2
  );


  buf

  (
    G1287_o2_p,
    G1287_o2
  );


  not

  (
    G1287_o2_n,
    G1287_o2
  );


  buf

  (
    G1266_o2_p,
    G1266_o2
  );


  not

  (
    G1266_o2_n,
    G1266_o2
  );


  buf

  (
    G1272_o2_p,
    G1272_o2
  );


  not

  (
    G1272_o2_n,
    G1272_o2
  );


  buf

  (
    G1278_o2_p,
    G1278_o2
  );


  not

  (
    G1278_o2_n,
    G1278_o2
  );


  buf

  (
    G1281_o2_p,
    G1281_o2
  );


  not

  (
    G1281_o2_n,
    G1281_o2
  );


  buf

  (
    G1284_o2_p,
    G1284_o2
  );


  not

  (
    G1284_o2_n,
    G1284_o2
  );


  buf

  (
    G1290_o2_p,
    G1290_o2
  );


  not

  (
    G1290_o2_n,
    G1290_o2
  );


  buf

  (
    G1293_o2_p,
    G1293_o2
  );


  not

  (
    G1293_o2_n,
    G1293_o2
  );


  buf

  (
    G1299_o2_p,
    G1299_o2
  );


  not

  (
    G1299_o2_n,
    G1299_o2
  );


  buf

  (
    G1305_o2_p,
    G1305_o2
  );


  not

  (
    G1305_o2_n,
    G1305_o2
  );


  buf

  (
    G1296_o2_p,
    G1296_o2
  );


  not

  (
    G1296_o2_n,
    G1296_o2
  );


  buf

  (
    G1302_o2_p,
    G1302_o2
  );


  not

  (
    G1302_o2_n,
    G1302_o2
  );


  buf

  (
    G1308_o2_p,
    G1308_o2
  );


  not

  (
    G1308_o2_n,
    G1308_o2
  );


  buf

  (
    G1311_o2_p,
    G1311_o2
  );


  not

  (
    G1311_o2_n,
    G1311_o2
  );


  buf

  (
    G811_o2_p,
    G811_o2
  );


  not

  (
    G811_o2_n,
    G811_o2
  );


  buf

  (
    G810_o2_p,
    G810_o2
  );


  not

  (
    G810_o2_n,
    G810_o2
  );


  buf

  (
    G1728_o2_p,
    G1728_o2
  );


  not

  (
    G1728_o2_n,
    G1728_o2
  );


  buf

  (
    G2512_o2_p,
    G2512_o2
  );


  not

  (
    G2512_o2_n,
    G2512_o2
  );


  buf

  (
    G1114_o2_p,
    G1114_o2
  );


  not

  (
    G1114_o2_n,
    G1114_o2
  );


  buf

  (
    G1113_o2_p,
    G1113_o2
  );


  not

  (
    G1113_o2_n,
    G1113_o2
  );


  buf

  (
    G1992_o2_p,
    G1992_o2
  );


  not

  (
    G1992_o2_n,
    G1992_o2
  );


  buf

  (
    G1991_o2_p,
    G1991_o2
  );


  not

  (
    G1991_o2_n,
    G1991_o2
  );


  buf

  (
    G1426_o2_p,
    G1426_o2
  );


  not

  (
    G1426_o2_n,
    G1426_o2
  );


  buf

  (
    G1966_o2_p,
    G1966_o2
  );


  not

  (
    G1966_o2_n,
    G1966_o2
  );


  buf

  (
    G2211_o2_p,
    G2211_o2
  );


  not

  (
    G2211_o2_n,
    G2211_o2
  );


  buf

  (
    G1509_o2_p,
    G1509_o2
  );


  not

  (
    G1509_o2_n,
    G1509_o2
  );


  buf

  (
    G2153_o2_p,
    G2153_o2
  );


  not

  (
    G2153_o2_n,
    G2153_o2
  );


  buf

  (
    G2329_o2_p,
    G2329_o2
  );


  not

  (
    G2329_o2_n,
    G2329_o2
  );


  buf

  (
    G1540_o2_p,
    G1540_o2
  );


  not

  (
    G1540_o2_n,
    G1540_o2
  );


  buf

  (
    G2167_o2_p,
    G2167_o2
  );


  not

  (
    G2167_o2_n,
    G2167_o2
  );


  buf

  (
    G2191_o2_p,
    G2191_o2
  );


  not

  (
    G2191_o2_n,
    G2191_o2
  );


  buf

  (
    G1234_o2_p,
    G1234_o2
  );


  not

  (
    G1234_o2_n,
    G1234_o2
  );


  buf

  (
    G1132_o2_p,
    G1132_o2
  );


  not

  (
    G1132_o2_n,
    G1132_o2
  );


  buf

  (
    G1129_o2_p,
    G1129_o2
  );


  not

  (
    G1129_o2_n,
    G1129_o2
  );


  buf

  (
    G2088_o2_p,
    G2088_o2
  );


  not

  (
    G2088_o2_n,
    G2088_o2
  );


  buf

  (
    G2106_o2_p,
    G2106_o2
  );


  not

  (
    G2106_o2_n,
    G2106_o2
  );


  buf

  (
    G1314_o2_p,
    G1314_o2
  );


  not

  (
    G1314_o2_n,
    G1314_o2
  );


  buf

  (
    G636_o2_p,
    G636_o2
  );


  not

  (
    G636_o2_n,
    G636_o2
  );


  buf

  (
    G647_o2_p,
    G647_o2
  );


  not

  (
    G647_o2_n,
    G647_o2
  );


  buf

  (
    n3186_lo_buf_o2_p,
    n3186_lo_buf_o2
  );


  not

  (
    n3186_lo_buf_o2_n,
    n3186_lo_buf_o2
  );


  buf

  (
    n3198_lo_buf_o2_p,
    n3198_lo_buf_o2
  );


  not

  (
    n3198_lo_buf_o2_n,
    n3198_lo_buf_o2
  );


  buf

  (
    n3210_lo_buf_o2_p,
    n3210_lo_buf_o2
  );


  not

  (
    n3210_lo_buf_o2_n,
    n3210_lo_buf_o2
  );


  buf

  (
    n3222_lo_buf_o2_p,
    n3222_lo_buf_o2
  );


  not

  (
    n3222_lo_buf_o2_n,
    n3222_lo_buf_o2
  );


  buf

  (
    G1225_o2_p,
    G1225_o2
  );


  not

  (
    G1225_o2_n,
    G1225_o2
  );


  buf

  (
    G1342_o2_p,
    G1342_o2
  );


  not

  (
    G1342_o2_n,
    G1342_o2
  );


  buf

  (
    G1222_o2_p,
    G1222_o2
  );


  not

  (
    G1222_o2_n,
    G1222_o2
  );


  buf

  (
    G1228_o2_p,
    G1228_o2
  );


  not

  (
    G1228_o2_n,
    G1228_o2
  );


  buf

  (
    G1348_o2_p,
    G1348_o2
  );


  not

  (
    G1348_o2_n,
    G1348_o2
  );


  buf

  (
    G1345_o2_p,
    G1345_o2
  );


  not

  (
    G1345_o2_n,
    G1345_o2
  );


  buf

  (
    G1351_o2_p,
    G1351_o2
  );


  not

  (
    G1351_o2_n,
    G1351_o2
  );


  buf

  (
    G2242_o2_p,
    G2242_o2
  );


  not

  (
    G2242_o2_n,
    G2242_o2
  );


  buf

  (
    G2260_o2_p,
    G2260_o2
  );


  not

  (
    G2260_o2_n,
    G2260_o2
  );


  buf

  (
    G1374_o2_p,
    G1374_o2
  );


  not

  (
    G1374_o2_n,
    G1374_o2
  );


  buf

  (
    G1537_o2_p,
    G1537_o2
  );


  not

  (
    G1537_o2_n,
    G1537_o2
  );


  buf

  (
    G301_o2_p,
    G301_o2
  );


  not

  (
    G301_o2_n,
    G301_o2
  );


  buf

  (
    G313_o2_p,
    G313_o2
  );


  not

  (
    G313_o2_n,
    G313_o2
  );


  buf

  (
    G2365_o2_p,
    G2365_o2
  );


  not

  (
    G2365_o2_n,
    G2365_o2
  );


  buf

  (
    G2255_o2_p,
    G2255_o2
  );


  not

  (
    G2255_o2_n,
    G2255_o2
  );


  buf

  (
    G2253_o2_p,
    G2253_o2
  );


  not

  (
    G2253_o2_n,
    G2253_o2
  );


  buf

  (
    G2395_o2_p,
    G2395_o2
  );


  not

  (
    G2395_o2_n,
    G2395_o2
  );


  buf

  (
    G2272_o2_p,
    G2272_o2
  );


  not

  (
    G2272_o2_n,
    G2272_o2
  );


  buf

  (
    G2270_o2_p,
    G2270_o2
  );


  not

  (
    G2270_o2_n,
    G2270_o2
  );


  buf

  (
    G2245_o2_p,
    G2245_o2
  );


  not

  (
    G2245_o2_n,
    G2245_o2
  );


  buf

  (
    G2262_o2_p,
    G2262_o2
  );


  not

  (
    G2262_o2_n,
    G2262_o2
  );


  buf

  (
    G2249_o2_p,
    G2249_o2
  );


  not

  (
    G2249_o2_n,
    G2249_o2
  );


  buf

  (
    G2247_o2_p,
    G2247_o2
  );


  not

  (
    G2247_o2_n,
    G2247_o2
  );


  buf

  (
    G2266_o2_p,
    G2266_o2
  );


  not

  (
    G2266_o2_n,
    G2266_o2
  );


  buf

  (
    G2264_o2_p,
    G2264_o2
  );


  not

  (
    G2264_o2_n,
    G2264_o2
  );


  buf

  (
    G2403_o2_p,
    G2403_o2
  );


  not

  (
    G2403_o2_n,
    G2403_o2
  );


  buf

  (
    G2401_o2_p,
    G2401_o2
  );


  not

  (
    G2401_o2_n,
    G2401_o2
  );


  buf

  (
    G2410_o2_p,
    G2410_o2
  );


  not

  (
    G2410_o2_n,
    G2410_o2
  );


  buf

  (
    G2408_o2_p,
    G2408_o2
  );


  not

  (
    G2408_o2_n,
    G2408_o2
  );


  buf

  (
    G2306_o2_p,
    G2306_o2
  );


  not

  (
    G2306_o2_n,
    G2306_o2
  );


  buf

  (
    G2305_o2_p,
    G2305_o2
  );


  not

  (
    G2305_o2_n,
    G2305_o2
  );


  buf

  (
    G2314_o2_p,
    G2314_o2
  );


  not

  (
    G2314_o2_n,
    G2314_o2
  );


  buf

  (
    G2313_o2_p,
    G2313_o2
  );


  not

  (
    G2313_o2_n,
    G2313_o2
  );


  buf

  (
    G2303_o2_p,
    G2303_o2
  );


  not

  (
    G2303_o2_n,
    G2303_o2
  );


  buf

  (
    G2302_o2_p,
    G2302_o2
  );


  not

  (
    G2302_o2_n,
    G2302_o2
  );


  buf

  (
    G2301_o2_p,
    G2301_o2
  );


  not

  (
    G2301_o2_n,
    G2301_o2
  );


  buf

  (
    G2311_o2_p,
    G2311_o2
  );


  not

  (
    G2311_o2_n,
    G2311_o2
  );


  buf

  (
    G2310_o2_p,
    G2310_o2
  );


  not

  (
    G2310_o2_n,
    G2310_o2
  );


  buf

  (
    G2309_o2_p,
    G2309_o2
  );


  not

  (
    G2309_o2_n,
    G2309_o2
  );


  buf

  (
    G2404_o2_p,
    G2404_o2
  );


  not

  (
    G2404_o2_n,
    G2404_o2
  );


  buf

  (
    G2411_o2_p,
    G2411_o2
  );


  not

  (
    G2411_o2_n,
    G2411_o2
  );


  buf

  (
    G2420_o2_p,
    G2420_o2
  );


  not

  (
    G2420_o2_n,
    G2420_o2
  );


  buf

  (
    G2419_o2_p,
    G2419_o2
  );


  not

  (
    G2419_o2_n,
    G2419_o2
  );


  buf

  (
    G2433_o2_p,
    G2433_o2
  );


  not

  (
    G2433_o2_n,
    G2433_o2
  );


  buf

  (
    G2432_o2_p,
    G2432_o2
  );


  not

  (
    G2432_o2_n,
    G2432_o2
  );


  buf

  (
    G402_o2_p,
    G402_o2
  );


  not

  (
    G402_o2_n,
    G402_o2
  );


  buf

  (
    G403_o2_p,
    G403_o2
  );


  not

  (
    G403_o2_n,
    G403_o2
  );


  buf

  (
    G1053_o2_p,
    G1053_o2
  );


  not

  (
    G1053_o2_n,
    G1053_o2
  );


  buf

  (
    G1049_o2_p,
    G1049_o2
  );


  not

  (
    G1049_o2_n,
    G1049_o2
  );


  buf

  (
    n2003_inv_p,
    n2003_inv
  );


  not

  (
    n2003_inv_n,
    n2003_inv
  );


  buf

  (
    G1364_o2_p,
    G1364_o2
  );


  not

  (
    G1364_o2_n,
    G1364_o2
  );


  buf

  (
    G1079_o2_p,
    G1079_o2
  );


  not

  (
    G1079_o2_n,
    G1079_o2
  );


  buf

  (
    G1478_o2_p,
    G1478_o2
  );


  not

  (
    G1478_o2_n,
    G1478_o2
  );


  buf

  (
    G707_o2_p,
    G707_o2
  );


  not

  (
    G707_o2_n,
    G707_o2
  );


  buf

  (
    G718_o2_p,
    G718_o2
  );


  not

  (
    G718_o2_n,
    G718_o2
  );


  buf

  (
    G2417_o2_p,
    G2417_o2
  );


  not

  (
    G2417_o2_n,
    G2417_o2
  );


  buf

  (
    G2414_o2_p,
    G2414_o2
  );


  not

  (
    G2414_o2_n,
    G2414_o2
  );


  buf

  (
    G2431_o2_p,
    G2431_o2
  );


  not

  (
    G2431_o2_n,
    G2431_o2
  );


  buf

  (
    G2428_o2_p,
    G2428_o2
  );


  not

  (
    G2428_o2_n,
    G2428_o2
  );


  buf

  (
    G1653_o2_p,
    G1653_o2
  );


  not

  (
    G1653_o2_n,
    G1653_o2
  );


  buf

  (
    G2213_o2_p,
    G2213_o2
  );


  not

  (
    G2213_o2_n,
    G2213_o2
  );


  buf

  (
    G2221_o2_p,
    G2221_o2
  );


  not

  (
    G2221_o2_n,
    G2221_o2
  );


  buf

  (
    G2250_o2_p,
    G2250_o2
  );


  not

  (
    G2250_o2_n,
    G2250_o2
  );


  buf

  (
    G2267_o2_p,
    G2267_o2
  );


  not

  (
    G2267_o2_n,
    G2267_o2
  );


  buf

  (
    G1365_o2_p,
    G1365_o2
  );


  not

  (
    G1365_o2_n,
    G1365_o2
  );


  buf

  (
    G1368_o2_p,
    G1368_o2
  );


  not

  (
    G1368_o2_n,
    G1368_o2
  );


  buf

  (
    G1371_o2_p,
    G1371_o2
  );


  not

  (
    G1371_o2_n,
    G1371_o2
  );


  buf

  (
    G2218_o2_p,
    G2218_o2
  );


  not

  (
    G2218_o2_n,
    G2218_o2
  );


  buf

  (
    G2225_o2_p,
    G2225_o2
  );


  not

  (
    G2225_o2_n,
    G2225_o2
  );


  buf

  (
    n1503_lo_buf_o2_p,
    n1503_lo_buf_o2
  );


  not

  (
    n1503_lo_buf_o2_n,
    n1503_lo_buf_o2
  );


  buf

  (
    n1863_lo_buf_o2_p,
    n1863_lo_buf_o2
  );


  not

  (
    n1863_lo_buf_o2_n,
    n1863_lo_buf_o2
  );


  buf

  (
    n1887_lo_buf_o2_p,
    n1887_lo_buf_o2
  );


  not

  (
    n1887_lo_buf_o2_n,
    n1887_lo_buf_o2
  );


  buf

  (
    n1983_lo_buf_o2_p,
    n1983_lo_buf_o2
  );


  not

  (
    n1983_lo_buf_o2_n,
    n1983_lo_buf_o2
  );


  buf

  (
    n2007_lo_buf_o2_p,
    n2007_lo_buf_o2
  );


  not

  (
    n2007_lo_buf_o2_n,
    n2007_lo_buf_o2
  );


  buf

  (
    n2115_lo_buf_o2_p,
    n2115_lo_buf_o2
  );


  not

  (
    n2115_lo_buf_o2_n,
    n2115_lo_buf_o2
  );


  buf

  (
    n2139_lo_buf_o2_p,
    n2139_lo_buf_o2
  );


  not

  (
    n2139_lo_buf_o2_n,
    n2139_lo_buf_o2
  );


  buf

  (
    n2247_lo_buf_o2_p,
    n2247_lo_buf_o2
  );


  not

  (
    n2247_lo_buf_o2_n,
    n2247_lo_buf_o2
  );


  buf

  (
    n2271_lo_buf_o2_p,
    n2271_lo_buf_o2
  );


  not

  (
    n2271_lo_buf_o2_n,
    n2271_lo_buf_o2
  );


  buf

  (
    n2919_lo_buf_o2_p,
    n2919_lo_buf_o2
  );


  not

  (
    n2919_lo_buf_o2_n,
    n2919_lo_buf_o2
  );


  buf

  (
    n2943_lo_buf_o2_p,
    n2943_lo_buf_o2
  );


  not

  (
    n2943_lo_buf_o2_n,
    n2943_lo_buf_o2
  );


  buf

  (
    n2967_lo_buf_o2_p,
    n2967_lo_buf_o2
  );


  not

  (
    n2967_lo_buf_o2_n,
    n2967_lo_buf_o2
  );


  buf

  (
    n2979_lo_buf_o2_p,
    n2979_lo_buf_o2
  );


  not

  (
    n2979_lo_buf_o2_n,
    n2979_lo_buf_o2
  );


  buf

  (
    n3063_lo_buf_o2_p,
    n3063_lo_buf_o2
  );


  not

  (
    n3063_lo_buf_o2_n,
    n3063_lo_buf_o2
  );


  buf

  (
    n3075_lo_buf_o2_p,
    n3075_lo_buf_o2
  );


  not

  (
    n3075_lo_buf_o2_n,
    n3075_lo_buf_o2
  );


  buf

  (
    n3099_lo_buf_o2_p,
    n3099_lo_buf_o2
  );


  not

  (
    n3099_lo_buf_o2_n,
    n3099_lo_buf_o2
  );


  buf

  (
    n3111_lo_buf_o2_p,
    n3111_lo_buf_o2
  );


  not

  (
    n3111_lo_buf_o2_n,
    n3111_lo_buf_o2
  );


  buf

  (
    G878_o2_p,
    G878_o2
  );


  not

  (
    G878_o2_n,
    G878_o2
  );


  buf

  (
    G875_o2_p,
    G875_o2
  );


  not

  (
    G875_o2_n,
    G875_o2
  );


  buf

  (
    G661_o2_p,
    G661_o2
  );


  not

  (
    G661_o2_n,
    G661_o2
  );


  buf

  (
    G660_o2_p,
    G660_o2
  );


  not

  (
    G660_o2_n,
    G660_o2
  );


  buf

  (
    G879_o2_p,
    G879_o2
  );


  not

  (
    G879_o2_n,
    G879_o2
  );


  buf

  (
    G876_o2_p,
    G876_o2
  );


  not

  (
    G876_o2_n,
    G876_o2
  );


  buf

  (
    G1320_o2_p,
    G1320_o2
  );


  not

  (
    G1320_o2_n,
    G1320_o2
  );


  buf

  (
    G941_o2_p,
    G941_o2
  );


  not

  (
    G941_o2_n,
    G941_o2
  );


  buf

  (
    G732_o2_p,
    G732_o2
  );


  not

  (
    G732_o2_n,
    G732_o2
  );


  buf

  (
    G942_o2_p,
    G942_o2
  );


  not

  (
    G942_o2_n,
    G942_o2
  );


  buf

  (
    G1493_o2_p,
    G1493_o2
  );


  not

  (
    G1493_o2_n,
    G1493_o2
  );


  buf

  (
    G1498_o2_p,
    G1498_o2
  );


  not

  (
    G1498_o2_n,
    G1498_o2
  );


  buf

  (
    G877_o2_p,
    G877_o2
  );


  not

  (
    G877_o2_n,
    G877_o2
  );


  buf

  (
    G874_o2_p,
    G874_o2
  );


  not

  (
    G874_o2_n,
    G874_o2
  );


  buf

  (
    n1806_lo_buf_o2_p,
    n1806_lo_buf_o2
  );


  not

  (
    n1806_lo_buf_o2_n,
    n1806_lo_buf_o2
  );


  buf

  (
    n1878_lo_buf_o2_p,
    n1878_lo_buf_o2
  );


  not

  (
    n1878_lo_buf_o2_n,
    n1878_lo_buf_o2
  );


  buf

  (
    n1938_lo_buf_o2_p,
    n1938_lo_buf_o2
  );


  not

  (
    n1938_lo_buf_o2_n,
    n1938_lo_buf_o2
  );


  buf

  (
    n1998_lo_buf_o2_p,
    n1998_lo_buf_o2
  );


  not

  (
    n1998_lo_buf_o2_n,
    n1998_lo_buf_o2
  );


  buf

  (
    n2058_lo_buf_o2_p,
    n2058_lo_buf_o2
  );


  not

  (
    n2058_lo_buf_o2_n,
    n2058_lo_buf_o2
  );


  buf

  (
    n2130_lo_buf_o2_p,
    n2130_lo_buf_o2
  );


  not

  (
    n2130_lo_buf_o2_n,
    n2130_lo_buf_o2
  );


  buf

  (
    n2190_lo_buf_o2_p,
    n2190_lo_buf_o2
  );


  not

  (
    n2190_lo_buf_o2_n,
    n2190_lo_buf_o2
  );


  buf

  (
    n2262_lo_buf_o2_p,
    n2262_lo_buf_o2
  );


  not

  (
    n2262_lo_buf_o2_n,
    n2262_lo_buf_o2
  );


  buf

  (
    n2310_lo_buf_o2_p,
    n2310_lo_buf_o2
  );


  not

  (
    n2310_lo_buf_o2_n,
    n2310_lo_buf_o2
  );


  buf

  (
    n2406_lo_buf_o2_p,
    n2406_lo_buf_o2
  );


  not

  (
    n2406_lo_buf_o2_n,
    n2406_lo_buf_o2
  );


  buf

  (
    n2430_lo_buf_o2_p,
    n2430_lo_buf_o2
  );


  not

  (
    n2430_lo_buf_o2_n,
    n2430_lo_buf_o2
  );


  buf

  (
    n2526_lo_buf_o2_p,
    n2526_lo_buf_o2
  );


  not

  (
    n2526_lo_buf_o2_n,
    n2526_lo_buf_o2
  );


  buf

  (
    n2550_lo_buf_o2_p,
    n2550_lo_buf_o2
  );


  not

  (
    n2550_lo_buf_o2_n,
    n2550_lo_buf_o2
  );


  buf

  (
    n2646_lo_buf_o2_p,
    n2646_lo_buf_o2
  );


  not

  (
    n2646_lo_buf_o2_n,
    n2646_lo_buf_o2
  );


  buf

  (
    n2670_lo_buf_o2_p,
    n2670_lo_buf_o2
  );


  not

  (
    n2670_lo_buf_o2_n,
    n2670_lo_buf_o2
  );


  buf

  (
    n2766_lo_buf_o2_p,
    n2766_lo_buf_o2
  );


  not

  (
    n2766_lo_buf_o2_n,
    n2766_lo_buf_o2
  );


  buf

  (
    G603_o2_p,
    G603_o2
  );


  not

  (
    G603_o2_n,
    G603_o2
  );


  buf

  (
    G614_o2_p,
    G614_o2
  );


  not

  (
    G614_o2_n,
    G614_o2
  );


  buf

  (
    G1026_o2_p,
    G1026_o2
  );


  not

  (
    G1026_o2_n,
    G1026_o2
  );


  buf

  (
    G1021_o2_p,
    G1021_o2
  );


  not

  (
    G1021_o2_n,
    G1021_o2
  );


  buf

  (
    G940_o2_p,
    G940_o2
  );


  not

  (
    G940_o2_n,
    G940_o2
  );


  buf

  (
    G1636_o2_p,
    G1636_o2
  );


  not

  (
    G1636_o2_n,
    G1636_o2
  );


  buf

  (
    G1684_o2_p,
    G1684_o2
  );


  not

  (
    G1684_o2_n,
    G1684_o2
  );


  buf

  (
    n2352_lo_buf_o2_p,
    n2352_lo_buf_o2
  );


  not

  (
    n2352_lo_buf_o2_n,
    n2352_lo_buf_o2
  );


  buf

  (
    n2364_lo_buf_o2_p,
    n2364_lo_buf_o2
  );


  not

  (
    n2364_lo_buf_o2_n,
    n2364_lo_buf_o2
  );


  buf

  (
    n2472_lo_buf_o2_p,
    n2472_lo_buf_o2
  );


  not

  (
    n2472_lo_buf_o2_n,
    n2472_lo_buf_o2
  );


  buf

  (
    n2484_lo_buf_o2_p,
    n2484_lo_buf_o2
  );


  not

  (
    n2484_lo_buf_o2_n,
    n2484_lo_buf_o2
  );


  buf

  (
    n2592_lo_buf_o2_p,
    n2592_lo_buf_o2
  );


  not

  (
    n2592_lo_buf_o2_n,
    n2592_lo_buf_o2
  );


  buf

  (
    n2604_lo_buf_o2_p,
    n2604_lo_buf_o2
  );


  not

  (
    n2604_lo_buf_o2_n,
    n2604_lo_buf_o2
  );


  buf

  (
    n2712_lo_buf_o2_p,
    n2712_lo_buf_o2
  );


  not

  (
    n2712_lo_buf_o2_n,
    n2712_lo_buf_o2
  );


  buf

  (
    n2724_lo_buf_o2_p,
    n2724_lo_buf_o2
  );


  not

  (
    n2724_lo_buf_o2_n,
    n2724_lo_buf_o2
  );


  buf

  (
    n3150_lo_buf_o2_p,
    n3150_lo_buf_o2
  );


  not

  (
    n3150_lo_buf_o2_n,
    n3150_lo_buf_o2
  );


  buf

  (
    n3162_lo_buf_o2_p,
    n3162_lo_buf_o2
  );


  not

  (
    n3162_lo_buf_o2_n,
    n3162_lo_buf_o2
  );


  or

  (
    g835_n,
    n3117_lo_n,
    n3105_lo_n
  );


  or

  (
    g836_n,
    g835_n,
    n3093_lo_n
  );


  or

  (
    g837_n,
    g836_n,
    n3081_lo_n
  );


  or

  (
    g838_n,
    n1545_lo_n,
    n1437_lo_n
  );


  or

  (
    g839_n,
    g838_n,
    n2865_lo_n_spl_
  );


  and

  (
    g840_p,
    n2793_lo_n_spl_0,
    n2301_lo_p
  );


  or

  (
    g841_n,
    n2865_lo_n_spl_,
    n1497_lo_n
  );


  or

  (
    g842_n,
    g841_n_spl_0,
    n2841_lo_n
  );


  or

  (
    g843_n,
    g841_n_spl_0,
    n3177_lo_n
  );


  or

  (
    g844_n,
    n2565_lo_n_spl_,
    n1929_lo_n_spl_
  );


  or

  (
    g845_n,
    g844_n,
    n2445_lo_n_spl_
  );


  or

  (
    g846_n,
    g845_n,
    n2049_lo_n_spl_
  );


  or

  (
    g847_n,
    n2685_lo_n_spl_,
    n2181_lo_n_spl_
  );


  or

  (
    g848_n,
    g847_n,
    n2325_lo_n_spl_
  );


  or

  (
    g849_n,
    g848_n,
    n1797_lo_n_spl_
  );


  or

  (
    g850_n,
    g849_n_spl_,
    g846_n_spl_
  );


  and

  (
    g851_p,
    g849_n_spl_,
    n3177_lo_p
  );


  and

  (
    g852_p,
    g846_n_spl_,
    n2841_lo_p
  );


  or

  (
    g853_n,
    g852_p,
    g851_p
  );


  and

  (
    g854_p,
    n5178_o2_p,
    n2877_lo_p_spl_0
  );


  or

  (
    g855_n,
    g854_p,
    n2877_lo_n_spl_0
  );


  or

  (
    g856_n,
    n2865_lo_p,
    n2805_lo_n
  );


  or

  (
    g857_n,
    g856_n_spl_,
    n1749_lo_n
  );


  or

  (
    g858_n,
    g857_n,
    g853_n_spl_0
  );


  and

  (
    g859_p,
    n1449_lo_p,
    n1425_lo_p
  );


  or

  (
    g860_n,
    g856_n_spl_,
    g853_n_spl_0
  );


  or

  (
    g861_n,
    g860_n,
    g859_p
  );


  or

  (
    g862_n,
    n4928_o2_n,
    n2889_lo_p_spl_00
  );


  or

  (
    g863_n,
    n1235_inv_p_spl_,
    n2889_lo_n_spl_00
  );


  and

  (
    g864_p,
    g863_n,
    g862_n
  );


  or

  (
    g865_n,
    n1232_inv_p_spl_,
    n2889_lo_p_spl_00
  );


  or

  (
    g866_n,
    n4711_o2_n_spl_,
    n2889_lo_n_spl_00
  );


  and

  (
    g867_p,
    g866_n,
    g865_n
  );


  and

  (
    g868_p,
    G1321_o2_p,
    n2877_lo_n_spl_0
  );


  and

  (
    g869_p,
    n4928_o2_p,
    n2877_lo_p_spl_0
  );


  or

  (
    g870_n,
    g869_p,
    g868_p
  );


  or

  (
    g871_n,
    n5178_o2_n,
    n2889_lo_p_spl_0
  );


  or

  (
    g872_n,
    G1321_o2_n,
    n2889_lo_n_spl_0
  );


  and

  (
    g873_p,
    g872_n,
    g871_n
  );


  or

  (
    g874_n,
    n5479_o2_p,
    n3141_lo_p
  );


  and

  (
    g875_p,
    g874_n_spl_,
    n3141_lo_n
  );


  and

  (
    g876_p,
    g874_n_spl_,
    n5479_o2_n
  );


  or

  (
    g877_n,
    g876_p,
    g875_p
  );


  or

  (
    g878_n,
    n5477_o2_n_spl_,
    n3129_lo_p
  );


  and

  (
    g879_p,
    g878_n_spl_,
    n3129_lo_n
  );


  and

  (
    g880_p,
    g878_n_spl_,
    n5477_o2_p
  );


  or

  (
    g881_n,
    g880_p,
    g879_p
  );


  or

  (
    g882_n,
    g881_n,
    g877_n
  );


  or

  (
    g883_n,
    G1509_o2_n,
    G1260_o2_n
  );


  or

  (
    g884_n,
    G1426_o2_p,
    G1402_o2_p
  );


  and

  (
    g885_p,
    g884_n,
    g883_n
  );


  and

  (
    g886_p,
    g885_p,
    n1533_lo_p
  );


  and

  (
    g887_p,
    G810_o2_p,
    G578_o2_n
  );


  or

  (
    g887_n,
    G810_o2_n,
    G578_o2_p
  );


  and

  (
    g888_p,
    G811_o2_p,
    G575_o2_n
  );


  or

  (
    g888_n,
    G811_o2_n,
    G575_o2_p
  );


  and

  (
    g889_p,
    g888_n,
    g887_n
  );


  or

  (
    g889_n,
    g888_p,
    g887_p
  );


  and

  (
    g890_p,
    G1259_o2_n,
    G1367_o2_n
  );


  or

  (
    g890_n,
    G1259_o2_p,
    G1367_o2_p
  );


  and

  (
    g891_p,
    G1366_o2_n,
    G1258_o2_n
  );


  or

  (
    g891_n,
    G1366_o2_p,
    G1258_o2_p
  );


  and

  (
    g892_p,
    g891_p,
    g890_p
  );


  or

  (
    g892_n,
    g891_n,
    g890_n
  );


  or

  (
    g893_n,
    g892_n,
    g889_p
  );


  or

  (
    g894_n,
    g892_p,
    g889_n
  );


  and

  (
    g895_p,
    g894_n,
    g893_n
  );


  and

  (
    g896_p,
    G1113_o2_n,
    G987_o2_p
  );


  or

  (
    g896_n,
    G1113_o2_p,
    G987_o2_n
  );


  and

  (
    g897_p,
    G1114_o2_n,
    G984_o2_p
  );


  or

  (
    g897_n,
    G1114_o2_p,
    G984_o2_n
  );


  and

  (
    g898_p,
    g897_n,
    g896_n
  );


  or

  (
    g898_n,
    g897_p,
    g896_p
  );


  and

  (
    g899_p,
    G1254_o2_n,
    G1359_o2_n
  );


  or

  (
    g899_n,
    G1254_o2_p,
    G1359_o2_p
  );


  and

  (
    g900_p,
    G1358_o2_n,
    G1253_o2_n
  );


  or

  (
    g900_n,
    G1358_o2_p,
    G1253_o2_p
  );


  and

  (
    g901_p,
    g900_p,
    g899_p
  );


  or

  (
    g901_n,
    g900_n,
    g899_n
  );


  or

  (
    g902_n,
    g901_n,
    g898_p
  );


  or

  (
    g903_n,
    g901_p,
    g898_n
  );


  and

  (
    g904_p,
    g903_n,
    g902_n
  );


  and

  (
    g905_p,
    G1293_o2_p,
    G807_o2_n
  );


  and

  (
    g906_p,
    G1293_o2_n,
    G807_o2_p
  );


  or

  (
    g907_n,
    g906_p,
    g905_p
  );


  and

  (
    g908_p,
    G1290_o2_p,
    G804_o2_n
  );


  and

  (
    g909_p,
    G1290_o2_n,
    G804_o2_p
  );


  or

  (
    g910_n,
    g909_p,
    g908_p
  );


  and

  (
    g911_p,
    G1287_o2_p,
    G801_o2_n
  );


  and

  (
    g912_p,
    G1287_o2_n,
    G801_o2_p
  );


  or

  (
    g913_n,
    g912_p,
    g911_p
  );


  and

  (
    g914_p,
    G1284_o2_p,
    G798_o2_n
  );


  and

  (
    g915_p,
    G1284_o2_n,
    G798_o2_p
  );


  or

  (
    g916_n,
    g915_p,
    g914_p
  );


  and

  (
    g917_p,
    G1281_o2_p,
    G795_o2_n
  );


  and

  (
    g918_p,
    G1281_o2_n,
    G795_o2_p
  );


  or

  (
    g919_n,
    g918_p,
    g917_p
  );


  or

  (
    g920_n,
    g910_n,
    g907_n
  );


  or

  (
    g921_n,
    g920_n,
    g913_n
  );


  or

  (
    g922_n,
    g921_n,
    g916_n
  );


  or

  (
    g923_n,
    g922_n,
    g919_n
  );


  and

  (
    g924_p,
    G1278_o2_p,
    G792_o2_n
  );


  and

  (
    g925_p,
    G1278_o2_n,
    G792_o2_p
  );


  or

  (
    g926_n,
    g925_p,
    g924_p
  );


  and

  (
    g927_p,
    G1275_o2_p,
    G789_o2_n
  );


  and

  (
    g928_p,
    G1275_o2_n,
    G789_o2_p
  );


  or

  (
    g929_n,
    g928_p,
    g927_p
  );


  and

  (
    g930_p,
    G1272_o2_p,
    G786_o2_n
  );


  and

  (
    g931_p,
    G1272_o2_n,
    G786_o2_p
  );


  or

  (
    g932_n,
    g931_p,
    g930_p
  );


  and

  (
    g933_p,
    G1269_o2_p,
    G783_o2_n
  );


  and

  (
    g934_p,
    G1269_o2_n,
    G783_o2_p
  );


  or

  (
    g935_n,
    g934_p,
    g933_p
  );


  and

  (
    g936_p,
    G1266_o2_p,
    G780_o2_n
  );


  and

  (
    g937_p,
    G1266_o2_n,
    G780_o2_p
  );


  or

  (
    g938_n,
    g937_p,
    g936_p
  );


  or

  (
    g939_n,
    g929_n,
    g926_n
  );


  or

  (
    g940_n,
    g939_n,
    g932_n
  );


  or

  (
    g941_n,
    g940_n,
    g935_n
  );


  or

  (
    g942_n,
    g941_n,
    g938_n
  );


  or

  (
    g943_n,
    g942_n,
    g923_n
  );


  or

  (
    g944_n,
    G766_o2_n,
    n1677_lo_n
  );


  or

  (
    g945_n,
    G491_o2_p,
    n5477_o2_n_spl_
  );


  and

  (
    g946_p,
    g945_n,
    g944_n
  );


  and

  (
    g947_p,
    G1311_o2_p,
    G827_o2_n
  );


  and

  (
    g948_p,
    G1311_o2_n,
    G827_o2_p
  );


  or

  (
    g949_n,
    g948_p,
    g947_p
  );


  or

  (
    g950_n,
    g949_n,
    g946_p
  );


  and

  (
    g951_p,
    G1308_o2_p,
    G824_o2_n
  );


  and

  (
    g952_p,
    G1308_o2_n,
    G824_o2_p
  );


  or

  (
    g953_n,
    g952_p,
    g951_p
  );


  and

  (
    g954_p,
    G1305_o2_p,
    G821_o2_n
  );


  and

  (
    g955_p,
    G1305_o2_n,
    G821_o2_p
  );


  or

  (
    g956_n,
    g955_p,
    g954_p
  );


  and

  (
    g957_p,
    G1302_o2_p,
    G818_o2_n
  );


  and

  (
    g958_p,
    G1302_o2_n,
    G818_o2_p
  );


  or

  (
    g959_n,
    g958_p,
    g957_p
  );


  and

  (
    g960_p,
    G1299_o2_p,
    G815_o2_n
  );


  and

  (
    g961_p,
    G1299_o2_n,
    G815_o2_p
  );


  or

  (
    g962_n,
    g961_p,
    g960_p
  );


  and

  (
    g963_p,
    G1296_o2_p,
    G812_o2_n
  );


  and

  (
    g964_p,
    G1296_o2_n,
    G812_o2_p
  );


  or

  (
    g965_n,
    g964_p,
    g963_p
  );


  or

  (
    g966_n,
    g956_n,
    g953_n
  );


  or

  (
    g967_n,
    g966_n,
    g959_n
  );


  or

  (
    g968_n,
    g967_n,
    g962_n
  );


  or

  (
    g969_n,
    g968_n,
    g965_n
  );


  or

  (
    g970_n,
    g969_n,
    g950_n
  );


  or

  (
    g971_n,
    n2889_lo_p_spl_1,
    n1521_lo_n_spl_
  );


  or

  (
    g972_n,
    n2889_lo_n_spl_1,
    n1521_lo_n_spl_
  );


  and

  (
    g973_p,
    g972_n,
    g971_n
  );


  or

  (
    g974_n,
    g970_n,
    g943_n
  );


  or

  (
    g975_n,
    g974_n,
    g973_p
  );


  and

  (
    g976_p,
    G1728_o2_n_spl_,
    G1572_o2_p_spl_
  );


  or

  (
    g976_n,
    G1728_o2_p_spl_,
    G1572_o2_n_spl_
  );


  and

  (
    g977_p,
    G1728_o2_p_spl_,
    G1572_o2_n_spl_
  );


  or

  (
    g977_n,
    G1728_o2_n_spl_,
    G1572_o2_p_spl_
  );


  and

  (
    g978_p,
    g977_n,
    g976_n
  );


  or

  (
    g978_n,
    g977_p,
    g976_p
  );


  and

  (
    g979_p,
    g978_n,
    n5179_o2_n
  );


  and

  (
    g980_p,
    g978_p,
    n5179_o2_p_spl_0
  );


  or

  (
    g981_n,
    g980_p,
    g979_p
  );


  and

  (
    g982_p,
    g981_n,
    n2877_lo_n_spl_
  );


  and

  (
    g983_p,
    n5179_o2_p_spl_0,
    n2877_lo_p_spl_
  );


  or

  (
    g984_n,
    g983_p,
    g982_p
  );


  or

  (
    g985_n,
    G2153_o2_p,
    G1865_o2_p
  );


  or

  (
    g986_n,
    G1966_o2_n,
    G2048_o2_n
  );


  and

  (
    g987_p,
    g986_n,
    g985_n
  );


  and

  (
    g988_p,
    g987_p,
    n1761_lo_n_spl_
  );


  or

  (
    g989_n,
    n5179_o2_p_spl_,
    n2889_lo_p_spl_1
  );


  and

  (
    g990_p,
    G1991_o2_n,
    G1862_o2_p
  );


  or

  (
    g990_n,
    G1991_o2_p,
    G1862_o2_n
  );


  and

  (
    g991_p,
    G1992_o2_n,
    G1859_o2_p
  );


  or

  (
    g991_n,
    G1992_o2_p,
    G1859_o2_n
  );


  and

  (
    g992_p,
    g991_n,
    g990_n
  );


  or

  (
    g992_n,
    g991_p,
    g990_p
  );


  and

  (
    g993_p,
    G2058_o2_n,
    G2118_o2_p
  );


  or

  (
    g993_n,
    G2058_o2_p,
    G2118_o2_n
  );


  and

  (
    g994_p,
    G2117_o2_n,
    G2057_o2_n
  );


  or

  (
    g994_n,
    G2117_o2_p,
    G2057_o2_p
  );


  and

  (
    g995_p,
    g994_p,
    g993_p
  );


  or

  (
    g995_n,
    g994_n,
    g993_n
  );


  or

  (
    g996_n,
    g995_n,
    g992_p
  );


  or

  (
    g997_n,
    g995_p,
    g992_n
  );


  and

  (
    g998_p,
    g997_n,
    g996_n
  );


  or

  (
    g999_n,
    g998_p,
    n2889_lo_n_spl_1
  );


  and

  (
    g1000_p,
    g999_n,
    g989_n
  );


  or

  (
    g1001_n,
    G2329_o2_n,
    G2073_o2_n
  );


  or

  (
    g1002_n,
    G2211_o2_p,
    G2276_o2_p
  );


  and

  (
    g1003_p,
    g1002_n,
    g1001_n
  );


  and

  (
    g1004_p,
    g1003_p,
    n1761_lo_n_spl_
  );


  and

  (
    g1005_p,
    G2512_o2_p_spl_,
    n1448_inv_n
  );


  and

  (
    g1006_p,
    G2512_o2_p_spl_,
    G2505_o2_n
  );


  or

  (
    g1007_n,
    g1006_p,
    g1005_p
  );


  or

  (
    g1008_n,
    g1004_p_spl_,
    g988_p_spl_
  );


  or

  (
    g1009_n,
    g1008_n,
    g895_p_spl_
  );


  or

  (
    g1010_n,
    g904_p_spl_,
    g886_p_spl_
  );


  or

  (
    g1011_n,
    g1010_n,
    g1007_n_spl_
  );


  or

  (
    g1012_n,
    g1011_n,
    g1009_n
  );


  or

  (
    g1013_n,
    g1012_n,
    g853_n_spl_1
  );


  and

  (
    g1014_p,
    G1008_o2_n_spl_,
    n2826_lo_n
  );


  or

  (
    g1014_n,
    G1008_o2_p_spl_0,
    n2826_lo_p
  );


  or

  (
    g1015_n,
    G877_o2_p,
    G878_o2_p
  );


  or

  (
    g1016_n,
    g1015_n,
    G879_o2_p
  );


  or

  (
    g1017_n,
    g1016_n,
    G661_o2_p
  );


  or

  (
    g1018_n,
    G874_o2_p,
    G875_o2_p
  );


  or

  (
    g1019_n,
    g1018_n,
    G876_o2_p
  );


  or

  (
    g1020_n,
    g1019_n,
    G660_o2_p
  );


  or

  (
    g1021_n,
    G940_o2_p,
    G941_o2_p
  );


  or

  (
    g1022_n,
    g1021_n,
    G942_o2_p
  );


  or

  (
    g1023_n,
    g1022_n,
    G732_o2_p
  );


  and

  (
    g1024_p,
    n2190_lo_buf_o2_p,
    G636_o2_p_spl_
  );


  and

  (
    g1025_p,
    g1024_p,
    G647_o2_p_spl_
  );


  and

  (
    g1026_p,
    n1806_lo_buf_o2_p,
    G342_o2_n_spl_
  );


  and

  (
    g1027_p,
    g1026_p,
    G647_o2_p_spl_
  );


  and

  (
    g1028_p,
    n1938_lo_buf_o2_p,
    G636_o2_p_spl_
  );


  and

  (
    g1029_p,
    g1028_p,
    G354_o2_n_spl_
  );


  and

  (
    g1030_p,
    n2058_lo_buf_o2_p,
    G342_o2_n_spl_
  );


  and

  (
    g1031_p,
    g1030_p,
    G354_o2_n_spl_
  );


  or

  (
    g1032_n,
    g1027_p,
    g1025_p
  );


  or

  (
    g1033_n,
    g1032_n,
    g1029_p
  );


  or

  (
    g1034_n,
    g1033_n,
    g1031_p
  );


  and

  (
    g1035_p,
    n2670_lo_buf_o2_p,
    G707_o2_p_spl_00
  );


  and

  (
    g1036_p,
    g1035_p,
    G718_o2_p_spl_00
  );


  and

  (
    g1037_p,
    n2310_lo_buf_o2_p,
    G405_o2_n_spl_00
  );


  and

  (
    g1038_p,
    g1037_p,
    G718_o2_p_spl_00
  );


  and

  (
    g1039_p,
    n2550_lo_buf_o2_p,
    G707_o2_p_spl_00
  );


  and

  (
    g1040_p,
    g1039_p,
    G417_o2_n_spl_00
  );


  and

  (
    g1041_p,
    n2430_lo_buf_o2_p,
    G405_o2_n_spl_00
  );


  and

  (
    g1042_p,
    g1041_p,
    G417_o2_n_spl_00
  );


  or

  (
    g1043_n,
    g1038_p,
    g1036_p
  );


  or

  (
    g1044_n,
    g1043_n,
    g1040_p
  );


  or

  (
    g1045_n,
    g1044_n,
    g1042_p
  );


  and

  (
    g1046_p,
    n2766_lo_buf_o2_p,
    G707_o2_p_spl_01
  );


  and

  (
    g1047_p,
    g1046_p,
    G718_o2_p_spl_01
  );


  and

  (
    g1048_p,
    n2406_lo_buf_o2_p,
    G405_o2_n_spl_01
  );


  and

  (
    g1049_p,
    g1048_p,
    G718_o2_p_spl_01
  );


  and

  (
    g1050_p,
    n2646_lo_buf_o2_p,
    G707_o2_p_spl_01
  );


  and

  (
    g1051_p,
    g1050_p,
    G417_o2_n_spl_01
  );


  and

  (
    g1052_p,
    n2526_lo_buf_o2_p,
    G405_o2_n_spl_01
  );


  and

  (
    g1053_p,
    g1052_p,
    G417_o2_n_spl_01
  );


  or

  (
    g1054_n,
    g1049_p,
    g1047_p
  );


  or

  (
    g1055_n,
    g1054_n,
    g1051_p
  );


  or

  (
    g1056_n,
    g1055_n,
    g1053_p
  );


  and

  (
    g1057_p,
    G603_o2_p_spl_000,
    n2262_lo_buf_o2_p
  );


  or

  (
    g1057_n,
    G603_o2_n_spl_00,
    n2262_lo_buf_o2_n
  );


  and

  (
    g1058_p,
    g1057_p,
    G614_o2_p_spl_000
  );


  or

  (
    g1058_n,
    g1057_n,
    G614_o2_n_spl_00
  );


  and

  (
    g1059_p,
    n1878_lo_buf_o2_p,
    G301_o2_n_spl_000
  );


  or

  (
    g1059_n,
    n1878_lo_buf_o2_n,
    G301_o2_p_spl_00
  );


  and

  (
    g1060_p,
    g1059_p,
    G614_o2_p_spl_000
  );


  or

  (
    g1060_n,
    g1059_n,
    G614_o2_n_spl_00
  );


  and

  (
    g1061_p,
    G603_o2_p_spl_000,
    n1998_lo_buf_o2_p
  );


  or

  (
    g1061_n,
    G603_o2_n_spl_00,
    n1998_lo_buf_o2_n
  );


  and

  (
    g1062_p,
    g1061_p,
    G313_o2_n_spl_000
  );


  or

  (
    g1062_n,
    g1061_n,
    G313_o2_p_spl_00
  );


  and

  (
    g1063_p,
    n2130_lo_buf_o2_p,
    G301_o2_n_spl_000
  );


  or

  (
    g1063_n,
    n2130_lo_buf_o2_n,
    G301_o2_p_spl_00
  );


  and

  (
    g1064_p,
    g1063_p,
    G313_o2_n_spl_000
  );


  or

  (
    g1064_n,
    g1063_n,
    G313_o2_p_spl_00
  );


  and

  (
    g1065_p,
    g1060_n,
    g1058_n
  );


  or

  (
    g1065_n,
    g1060_p,
    g1058_p
  );


  and

  (
    g1066_p,
    g1065_p,
    g1062_n
  );


  or

  (
    g1066_n,
    g1065_n,
    g1062_p
  );


  and

  (
    g1067_p,
    g1066_p,
    g1064_n
  );


  or

  (
    g1067_n,
    g1066_n,
    g1064_p
  );


  and

  (
    g1068_p,
    G603_o2_p_spl_001,
    n2247_lo_buf_o2_p
  );


  or

  (
    g1068_n,
    G603_o2_n_spl_01,
    n2247_lo_buf_o2_n
  );


  and

  (
    g1069_p,
    g1068_p,
    G614_o2_p_spl_001
  );


  or

  (
    g1069_n,
    g1068_n,
    G614_o2_n_spl_01
  );


  and

  (
    g1070_p,
    n1863_lo_buf_o2_p,
    G301_o2_n_spl_001
  );


  or

  (
    g1070_n,
    n1863_lo_buf_o2_n,
    G301_o2_p_spl_01
  );


  and

  (
    g1071_p,
    g1070_p,
    G614_o2_p_spl_001
  );


  or

  (
    g1071_n,
    g1070_n,
    G614_o2_n_spl_01
  );


  and

  (
    g1072_p,
    G603_o2_p_spl_001,
    n1983_lo_buf_o2_p
  );


  or

  (
    g1072_n,
    G603_o2_n_spl_01,
    n1983_lo_buf_o2_n
  );


  and

  (
    g1073_p,
    g1072_p,
    G313_o2_n_spl_001
  );


  or

  (
    g1073_n,
    g1072_n,
    G313_o2_p_spl_01
  );


  and

  (
    g1074_p,
    n2115_lo_buf_o2_p,
    G301_o2_n_spl_001
  );


  or

  (
    g1074_n,
    n2115_lo_buf_o2_n,
    G301_o2_p_spl_01
  );


  and

  (
    g1075_p,
    g1074_p,
    G313_o2_n_spl_001
  );


  or

  (
    g1075_n,
    g1074_n,
    G313_o2_p_spl_01
  );


  and

  (
    g1076_p,
    g1071_n,
    g1069_n
  );


  or

  (
    g1076_n,
    g1071_p,
    g1069_p
  );


  and

  (
    g1077_p,
    g1076_p,
    g1073_n
  );


  or

  (
    g1077_n,
    g1076_n,
    g1073_p
  );


  and

  (
    g1078_p,
    g1077_p,
    g1075_n
  );


  or

  (
    g1078_n,
    g1077_n,
    g1075_p
  );


  and

  (
    g1079_p,
    G603_o2_p_spl_01,
    n2271_lo_buf_o2_p
  );


  or

  (
    g1079_n,
    G603_o2_n_spl_1,
    n2271_lo_buf_o2_n
  );


  and

  (
    g1080_p,
    g1079_p,
    G614_o2_p_spl_01
  );


  or

  (
    g1080_n,
    g1079_n,
    G614_o2_n_spl_1
  );


  and

  (
    g1081_p,
    n1887_lo_buf_o2_p,
    G301_o2_n_spl_01
  );


  or

  (
    g1081_n,
    n1887_lo_buf_o2_n,
    G301_o2_p_spl_1
  );


  and

  (
    g1082_p,
    g1081_p,
    G614_o2_p_spl_01
  );


  or

  (
    g1082_n,
    g1081_n,
    G614_o2_n_spl_1
  );


  and

  (
    g1083_p,
    G603_o2_p_spl_01,
    n2007_lo_buf_o2_p
  );


  or

  (
    g1083_n,
    G603_o2_n_spl_1,
    n2007_lo_buf_o2_n
  );


  and

  (
    g1084_p,
    g1083_p,
    G313_o2_n_spl_01
  );


  or

  (
    g1084_n,
    g1083_n,
    G313_o2_p_spl_1
  );


  and

  (
    g1085_p,
    n2139_lo_buf_o2_p,
    G301_o2_n_spl_01
  );


  or

  (
    g1085_n,
    n2139_lo_buf_o2_n,
    G301_o2_p_spl_1
  );


  and

  (
    g1086_p,
    g1085_p,
    G313_o2_n_spl_01
  );


  or

  (
    g1086_n,
    g1085_n,
    G313_o2_p_spl_1
  );


  and

  (
    g1087_p,
    g1082_n,
    g1080_n
  );


  or

  (
    g1087_n,
    g1082_p,
    g1080_p
  );


  and

  (
    g1088_p,
    g1087_p,
    g1084_n
  );


  or

  (
    g1088_n,
    g1087_n,
    g1084_p
  );


  and

  (
    g1089_p,
    g1088_p,
    g1086_n
  );


  or

  (
    g1089_n,
    g1088_n,
    g1086_p
  );


  and

  (
    g1090_p,
    G1636_o2_p_spl_000,
    n3075_lo_buf_o2_n_spl_
  );


  or

  (
    g1090_n,
    G1636_o2_n_spl_000,
    n3075_lo_buf_o2_p_spl_0
  );


  and

  (
    g1091_p,
    G1636_o2_n_spl_000,
    n2943_lo_buf_o2_n_spl_
  );


  or

  (
    g1091_n,
    G1636_o2_p_spl_000,
    n2943_lo_buf_o2_p_spl_0
  );


  and

  (
    g1092_p,
    g1091_n,
    g1090_n
  );


  or

  (
    g1092_n,
    g1091_p,
    g1090_p
  );


  and

  (
    g1093_p,
    G1684_o2_p_spl_000,
    n3075_lo_buf_o2_n_spl_
  );


  or

  (
    g1093_n,
    G1684_o2_n_spl_000,
    n3075_lo_buf_o2_p_spl_0
  );


  and

  (
    g1094_p,
    G1684_o2_n_spl_000,
    n2943_lo_buf_o2_n_spl_
  );


  or

  (
    g1094_n,
    G1684_o2_p_spl_000,
    n2943_lo_buf_o2_p_spl_0
  );


  and

  (
    g1095_p,
    g1094_n,
    g1093_n
  );


  or

  (
    g1095_n,
    g1094_p,
    g1093_p
  );


  and

  (
    g1096_p,
    G1899_o2_n,
    G2023_o2_p
  );


  or

  (
    g1097_n,
    G2301_o2_p,
    G2245_o2_n
  );


  and

  (
    g1098_p,
    G1896_o2_n,
    G2020_o2_p
  );


  and

  (
    g1099_p,
    g1098_p,
    g1097_n_spl_0
  );


  or

  (
    g1100_n,
    G2302_o2_p,
    G2247_o2_n
  );


  and

  (
    g1101_p,
    G1893_o2_n,
    G2017_o2_p
  );


  and

  (
    g1102_p,
    g1100_n_spl_0,
    g1097_n_spl_0
  );


  and

  (
    g1103_p,
    g1102_p,
    g1101_p
  );


  or

  (
    g1104_n,
    G2303_o2_p,
    G2249_o2_n
  );


  and

  (
    g1105_p,
    G1890_o2_n,
    G2014_o2_p
  );


  and

  (
    g1106_p,
    g1104_n_spl_,
    g1097_n_spl_1
  );


  and

  (
    g1107_p,
    g1106_p,
    g1105_p
  );


  and

  (
    g1108_p,
    g1107_p,
    g1100_n_spl_0
  );


  or

  (
    g1109_n,
    g1099_p,
    g1096_p
  );


  or

  (
    g1110_n,
    g1109_n,
    g1103_p
  );


  or

  (
    g1111_n,
    g1110_n,
    g1108_p
  );


  and

  (
    g1112_p,
    G1907_o2_n,
    G2011_o2_p
  );


  or

  (
    g1112_n,
    G1907_o2_p,
    G2011_o2_n
  );


  and

  (
    g1113_p,
    G2305_o2_n,
    G2253_o2_p
  );


  or

  (
    g1113_n,
    G2305_o2_p,
    G2253_o2_n
  );


  and

  (
    g1114_p,
    G1904_o2_n,
    G2008_o2_p
  );


  or

  (
    g1114_n,
    G1904_o2_p,
    G2008_o2_n
  );


  and

  (
    g1115_p,
    g1114_p,
    g1113_n_spl_00
  );


  or

  (
    g1115_n,
    g1114_n,
    g1113_p_spl_00
  );


  and

  (
    g1116_p,
    G2306_o2_n,
    G2255_o2_p
  );


  or

  (
    g1116_n,
    G2306_o2_p,
    G2255_o2_n
  );


  and

  (
    g1117_p,
    G1999_o2_n,
    G2231_o2_p
  );


  or

  (
    g1117_n,
    G1999_o2_p,
    G2231_o2_n
  );


  and

  (
    g1118_p,
    g1116_n_spl_0,
    g1113_n_spl_00
  );


  or

  (
    g1118_n,
    g1116_p_spl_0,
    g1113_p_spl_00
  );


  and

  (
    g1119_p,
    g1118_p,
    g1117_p
  );


  or

  (
    g1119_n,
    g1118_n,
    g1117_n
  );


  and

  (
    g1120_p,
    G2419_o2_n,
    G2401_o2_p
  );


  or

  (
    g1120_n,
    G2419_o2_p,
    G2401_o2_n
  );


  and

  (
    g1121_p,
    G1996_o2_n,
    G2228_o2_p
  );


  or

  (
    g1121_n,
    G1996_o2_p,
    G2228_o2_n
  );


  and

  (
    g1122_p,
    g1120_n_spl_0,
    g1113_n_spl_0
  );


  or

  (
    g1122_n,
    g1120_p_spl_0,
    g1113_p_spl_0
  );


  and

  (
    g1123_p,
    g1122_p,
    g1121_p
  );


  or

  (
    g1123_n,
    g1122_n,
    g1121_n
  );


  and

  (
    g1124_p,
    g1123_p,
    g1116_n_spl_0
  );


  or

  (
    g1124_n,
    g1123_n,
    g1116_p_spl_0
  );


  and

  (
    g1125_p,
    G2420_o2_n,
    G2403_o2_p
  );


  or

  (
    g1125_n,
    G2420_o2_p,
    G2403_o2_n
  );


  and

  (
    g1126_p,
    G1336_o2_p_spl_,
    G2141_o2_n
  );


  or

  (
    g1126_n,
    G1336_o2_n_spl_,
    G2141_o2_p
  );


  and

  (
    g1127_p,
    g1125_n_spl_,
    g1120_n_spl_0
  );


  or

  (
    g1127_n,
    g1125_p_spl_,
    g1120_p_spl_0
  );


  and

  (
    g1128_p,
    g1127_p,
    g1113_n_spl_1
  );


  or

  (
    g1128_n,
    g1127_n,
    g1113_p_spl_1
  );


  and

  (
    g1129_p,
    g1128_p,
    g1126_p
  );


  or

  (
    g1129_n,
    g1128_n,
    g1126_n
  );


  and

  (
    g1130_p,
    g1129_p,
    g1116_n_spl_1
  );


  or

  (
    g1130_n,
    g1129_n,
    g1116_p_spl_1
  );


  and

  (
    g1131_p,
    g1115_n,
    g1112_n
  );


  or

  (
    g1131_n,
    g1115_p,
    g1112_p
  );


  and

  (
    g1132_p,
    g1131_p,
    g1119_n
  );


  or

  (
    g1132_n,
    g1131_n,
    g1119_p
  );


  and

  (
    g1133_p,
    g1132_p,
    g1124_n
  );


  or

  (
    g1133_n,
    g1132_n,
    g1124_p
  );


  and

  (
    g1134_p,
    g1133_p,
    g1130_n
  );


  or

  (
    g1134_n,
    g1133_n,
    g1130_p
  );


  and

  (
    g1135_p,
    G2404_o2_p,
    G2365_o2_n
  );


  or

  (
    g1135_n,
    G2404_o2_n,
    G2365_o2_p
  );


  and

  (
    g1136_p,
    g1135_n,
    g1116_n_spl_1
  );


  or

  (
    g1136_n,
    g1135_p,
    g1116_p_spl_1
  );


  and

  (
    g1137_p,
    g1136_p,
    g1120_n_spl_
  );


  or

  (
    g1137_n,
    g1136_n,
    g1120_p_spl_
  );


  and

  (
    g1138_p,
    g1137_p,
    g1113_n_spl_1
  );


  or

  (
    g1138_n,
    g1137_n,
    g1113_p_spl_1
  );


  and

  (
    g1139_p,
    g1138_p,
    g1125_n_spl_
  );


  or

  (
    g1139_n,
    g1138_n,
    g1125_p_spl_
  );


  and

  (
    g1140_p,
    G1329_o2_p_spl_0,
    G2138_o2_n
  );


  or

  (
    g1140_n,
    G1329_o2_n_spl_0,
    G2138_o2_p
  );


  and

  (
    g1141_p,
    G2414_o2_n_spl_,
    G2242_o2_n
  );


  or

  (
    g1141_n,
    G2414_o2_p_spl_,
    G2242_o2_p
  );


  and

  (
    g1142_p,
    G2414_o2_n_spl_,
    G2417_o2_p
  );


  or

  (
    g1142_n,
    G2414_o2_p_spl_,
    G2417_o2_n
  );


  and

  (
    g1143_p,
    g1142_p,
    G2213_o2_n
  );


  or

  (
    g1143_n,
    g1142_n,
    G2213_o2_p
  );


  and

  (
    g1144_p,
    g1141_n,
    g1140_n
  );


  or

  (
    g1144_n,
    g1141_p,
    g1140_p
  );


  and

  (
    g1145_p,
    g1144_p,
    g1143_n
  );


  or

  (
    g1145_n,
    g1144_n,
    g1143_p
  );


  and

  (
    g1146_p,
    g1145_n,
    g1139_p
  );


  or

  (
    g1146_n,
    g1145_p,
    g1139_n
  );


  and

  (
    g1147_p,
    g1146_n,
    g1134_p
  );


  or

  (
    g1147_n,
    g1146_p,
    g1134_n
  );


  and

  (
    g1148_p,
    g1147_p,
    g1111_n_spl_
  );


  and

  (
    g1149_p,
    G2250_o2_p,
    G2088_o2_p
  );


  and

  (
    g1150_p,
    G2218_o2_n,
    G2167_o2_n
  );


  or

  (
    g1151_n,
    g1150_p,
    g1149_p
  );


  and

  (
    g1152_p,
    g1151_n,
    g1100_n_spl_
  );


  and

  (
    g1153_p,
    g1152_p,
    g1104_n_spl_
  );


  and

  (
    g1154_p,
    g1153_p,
    g1097_n_spl_1
  );


  or

  (
    g1155_n,
    g1154_p,
    g1111_n_spl_
  );


  and

  (
    g1156_p,
    g1155_n,
    g1147_n
  );


  or

  (
    g1157_n,
    g1156_p,
    g1148_p
  );


  and

  (
    g1158_p,
    G1943_o2_n,
    G2041_o2_p
  );


  or

  (
    g1159_n,
    G2309_o2_p,
    G2262_o2_n
  );


  and

  (
    g1160_p,
    G1940_o2_n,
    G2038_o2_p
  );


  and

  (
    g1161_p,
    g1160_p,
    g1159_n_spl_0
  );


  or

  (
    g1162_n,
    G2310_o2_p,
    G2264_o2_n
  );


  and

  (
    g1163_p,
    G1937_o2_n,
    G2035_o2_p
  );


  and

  (
    g1164_p,
    g1162_n_spl_0,
    g1159_n_spl_0
  );


  and

  (
    g1165_p,
    g1164_p,
    g1163_p
  );


  or

  (
    g1166_n,
    G2311_o2_p,
    G2266_o2_n
  );


  and

  (
    g1167_p,
    G1934_o2_n,
    G2032_o2_p
  );


  and

  (
    g1168_p,
    g1166_n_spl_,
    g1159_n_spl_1
  );


  and

  (
    g1169_p,
    g1168_p,
    g1167_p
  );


  and

  (
    g1170_p,
    g1169_p,
    g1162_n_spl_0
  );


  or

  (
    g1171_n,
    g1161_p,
    g1158_p
  );


  or

  (
    g1172_n,
    g1171_n,
    g1165_p
  );


  or

  (
    g1173_n,
    g1172_n,
    g1170_p
  );


  and

  (
    g1174_p,
    G1931_o2_n,
    G2029_o2_p
  );


  or

  (
    g1174_n,
    G1931_o2_p,
    G2029_o2_n
  );


  and

  (
    g1175_p,
    G2313_o2_n,
    G2270_o2_p
  );


  or

  (
    g1175_n,
    G2313_o2_p,
    G2270_o2_n
  );


  and

  (
    g1176_p,
    G1928_o2_n,
    G2026_o2_p
  );


  or

  (
    g1176_n,
    G1928_o2_p,
    G2026_o2_n
  );


  and

  (
    g1177_p,
    g1176_p,
    g1175_n_spl_00
  );


  or

  (
    g1177_n,
    g1176_n,
    g1175_p_spl_00
  );


  and

  (
    g1178_p,
    G2314_o2_n,
    G2272_o2_p
  );


  or

  (
    g1178_n,
    G2314_o2_p,
    G2272_o2_n
  );


  and

  (
    g1179_p,
    G2005_o2_n,
    G2237_o2_p
  );


  or

  (
    g1179_n,
    G2005_o2_p,
    G2237_o2_n
  );


  and

  (
    g1180_p,
    g1178_n_spl_0,
    g1175_n_spl_00
  );


  or

  (
    g1180_n,
    g1178_p_spl_0,
    g1175_p_spl_00
  );


  and

  (
    g1181_p,
    g1180_p,
    g1179_p
  );


  or

  (
    g1181_n,
    g1180_n,
    g1179_n
  );


  and

  (
    g1182_p,
    G2432_o2_n,
    G2408_o2_p
  );


  or

  (
    g1182_n,
    G2432_o2_p,
    G2408_o2_n
  );


  and

  (
    g1183_p,
    G2002_o2_n,
    G2234_o2_p
  );


  or

  (
    g1183_n,
    G2002_o2_p,
    G2234_o2_n
  );


  and

  (
    g1184_p,
    g1182_n_spl_0,
    g1175_n_spl_0
  );


  or

  (
    g1184_n,
    g1182_p_spl_0,
    g1175_p_spl_0
  );


  and

  (
    g1185_p,
    g1184_p,
    g1183_p
  );


  or

  (
    g1185_n,
    g1184_n,
    g1183_n
  );


  and

  (
    g1186_p,
    g1185_p,
    g1178_n_spl_0
  );


  or

  (
    g1186_n,
    g1185_n,
    g1178_p_spl_0
  );


  and

  (
    g1187_p,
    G2433_o2_n,
    G2410_o2_p
  );


  or

  (
    g1187_n,
    G2433_o2_p,
    G2410_o2_n
  );


  and

  (
    g1188_p,
    G1336_o2_p_spl_,
    G2150_o2_n
  );


  or

  (
    g1188_n,
    G1336_o2_n_spl_,
    G2150_o2_p
  );


  and

  (
    g1189_p,
    g1187_n_spl_,
    g1182_n_spl_0
  );


  or

  (
    g1189_n,
    g1187_p_spl_,
    g1182_p_spl_0
  );


  and

  (
    g1190_p,
    g1189_p,
    g1175_n_spl_1
  );


  or

  (
    g1190_n,
    g1189_n,
    g1175_p_spl_1
  );


  and

  (
    g1191_p,
    g1190_p,
    g1188_p
  );


  or

  (
    g1191_n,
    g1190_n,
    g1188_n
  );


  and

  (
    g1192_p,
    g1191_p,
    g1178_n_spl_1
  );


  or

  (
    g1192_n,
    g1191_n,
    g1178_p_spl_1
  );


  and

  (
    g1193_p,
    g1177_n,
    g1174_n
  );


  or

  (
    g1193_n,
    g1177_p,
    g1174_p
  );


  and

  (
    g1194_p,
    g1193_p,
    g1181_n
  );


  or

  (
    g1194_n,
    g1193_n,
    g1181_p
  );


  and

  (
    g1195_p,
    g1194_p,
    g1186_n
  );


  or

  (
    g1195_n,
    g1194_n,
    g1186_p
  );


  and

  (
    g1196_p,
    g1195_p,
    g1192_n
  );


  or

  (
    g1196_n,
    g1195_n,
    g1192_p
  );


  and

  (
    g1197_p,
    G2411_o2_p,
    G2395_o2_n
  );


  or

  (
    g1197_n,
    G2411_o2_n,
    G2395_o2_p
  );


  and

  (
    g1198_p,
    g1197_n,
    g1178_n_spl_1
  );


  or

  (
    g1198_n,
    g1197_p,
    g1178_p_spl_1
  );


  and

  (
    g1199_p,
    g1198_p,
    g1182_n_spl_
  );


  or

  (
    g1199_n,
    g1198_n,
    g1182_p_spl_
  );


  and

  (
    g1200_p,
    g1199_p,
    g1175_n_spl_1
  );


  or

  (
    g1200_n,
    g1199_n,
    g1175_p_spl_1
  );


  and

  (
    g1201_p,
    g1200_p,
    g1187_n_spl_
  );


  or

  (
    g1201_n,
    g1200_n,
    g1187_p_spl_
  );


  and

  (
    g1202_p,
    G1329_o2_p_spl_0,
    G2147_o2_n
  );


  or

  (
    g1202_n,
    G1329_o2_n_spl_0,
    G2147_o2_p
  );


  and

  (
    g1203_p,
    G2428_o2_n_spl_,
    G2260_o2_n
  );


  or

  (
    g1203_n,
    G2428_o2_p_spl_,
    G2260_o2_p
  );


  and

  (
    g1204_p,
    G2428_o2_n_spl_,
    G2431_o2_p
  );


  or

  (
    g1204_n,
    G2428_o2_p_spl_,
    G2431_o2_n
  );


  and

  (
    g1205_p,
    g1204_p,
    G2221_o2_n
  );


  or

  (
    g1205_n,
    g1204_n,
    G2221_o2_p
  );


  and

  (
    g1206_p,
    g1203_n,
    g1202_n
  );


  or

  (
    g1206_n,
    g1203_p,
    g1202_p
  );


  and

  (
    g1207_p,
    g1206_p,
    g1205_n
  );


  or

  (
    g1207_n,
    g1206_n,
    g1205_p
  );


  and

  (
    g1208_p,
    g1207_n,
    g1201_p
  );


  or

  (
    g1208_n,
    g1207_p,
    g1201_n
  );


  and

  (
    g1209_p,
    g1208_n,
    g1196_p
  );


  or

  (
    g1209_n,
    g1208_p,
    g1196_n
  );


  and

  (
    g1210_p,
    g1209_p,
    g1173_n_spl_
  );


  and

  (
    g1211_p,
    G2267_o2_p,
    G2106_o2_p
  );


  and

  (
    g1212_p,
    G2225_o2_n,
    G2191_o2_n
  );


  or

  (
    g1213_n,
    g1212_p,
    g1211_p
  );


  and

  (
    g1214_p,
    g1213_n,
    g1162_n_spl_
  );


  and

  (
    g1215_p,
    g1214_p,
    g1166_n_spl_
  );


  and

  (
    g1216_p,
    g1215_p,
    g1159_n_spl_1
  );


  or

  (
    g1217_n,
    g1216_p,
    g1173_n_spl_
  );


  and

  (
    g1218_p,
    g1217_n,
    g1209_n
  );


  or

  (
    g1219_n,
    g1218_p,
    g1210_p
  );


  and

  (
    g1220_p,
    n3018_lo_buf_o2_p,
    n3006_lo_buf_o2_n
  );


  and

  (
    g1221_p,
    n3018_lo_buf_o2_n,
    n3006_lo_buf_o2_p
  );


  or

  (
    g1222_n,
    g1221_p,
    g1220_p
  );


  and

  (
    g1223_p,
    n3042_lo_buf_o2_p,
    n3030_lo_buf_o2_n
  );


  and

  (
    g1224_p,
    n3042_lo_buf_o2_n,
    n3030_lo_buf_o2_p
  );


  or

  (
    g1225_n,
    g1224_p,
    g1223_p
  );


  and

  (
    g1226_p,
    G1345_o2_p_spl_,
    G1342_o2_n_spl_
  );


  or

  (
    g1226_n,
    G1345_o2_n_spl_,
    G1342_o2_p_spl_
  );


  and

  (
    g1227_p,
    G1345_o2_n_spl_,
    G1342_o2_p_spl_
  );


  or

  (
    g1227_n,
    G1345_o2_p_spl_,
    G1342_o2_n_spl_
  );


  and

  (
    g1228_p,
    g1227_n,
    g1226_n
  );


  or

  (
    g1228_n,
    g1227_p,
    g1226_p
  );


  and

  (
    g1229_p,
    G1351_o2_p_spl_,
    G1348_o2_n_spl_
  );


  or

  (
    g1229_n,
    G1351_o2_n_spl_,
    G1348_o2_p_spl_
  );


  and

  (
    g1230_p,
    G1351_o2_n_spl_,
    G1348_o2_p_spl_
  );


  or

  (
    g1230_n,
    G1351_o2_p_spl_,
    G1348_o2_n_spl_
  );


  and

  (
    g1231_p,
    g1230_n,
    g1229_n
  );


  or

  (
    g1231_n,
    g1230_p,
    g1229_p
  );


  and

  (
    g1232_p,
    n3270_lo_p_spl_,
    n3258_lo_n_spl_
  );


  or

  (
    g1232_n,
    n3270_lo_n_spl_,
    n3258_lo_p_spl_
  );


  and

  (
    g1233_p,
    n3270_lo_n_spl_,
    n3258_lo_p_spl_
  );


  or

  (
    g1233_n,
    n3270_lo_p_spl_,
    n3258_lo_n_spl_
  );


  and

  (
    g1234_p,
    g1233_n,
    g1232_n
  );


  or

  (
    g1234_n,
    g1233_p,
    g1232_p
  );


  and

  (
    g1235_p,
    n2910_lo_buf_o2_n_spl_,
    n2922_lo_buf_o2_p_spl_
  );


  or

  (
    g1235_n,
    n2910_lo_buf_o2_p_spl_,
    n2922_lo_buf_o2_n_spl_
  );


  and

  (
    g1236_p,
    n2910_lo_buf_o2_p_spl_,
    n2922_lo_buf_o2_n_spl_
  );


  or

  (
    g1236_n,
    n2910_lo_buf_o2_n_spl_,
    n2922_lo_buf_o2_p_spl_
  );


  and

  (
    g1237_p,
    g1236_n,
    g1235_n
  );


  or

  (
    g1237_n,
    g1236_p,
    g1235_p
  );


  and

  (
    g1238_p,
    g1237_p,
    g1234_n
  );


  and

  (
    g1239_p,
    g1237_n,
    g1234_p
  );


  or

  (
    g1240_n,
    g1239_p,
    g1238_p
  );


  and

  (
    g1241_p,
    G1049_o2_p_spl_0,
    n5222_o2_n_spl_
  );


  or

  (
    g1241_n,
    G1049_o2_n_spl_,
    n5222_o2_p_spl_0
  );


  and

  (
    g1242_p,
    G1049_o2_n_spl_,
    n5222_o2_p_spl_0
  );


  or

  (
    g1242_n,
    G1049_o2_p_spl_0,
    n5222_o2_n_spl_
  );


  and

  (
    g1243_p,
    g1242_n,
    g1241_n
  );


  or

  (
    g1243_n,
    g1242_p,
    g1241_p
  );


  and

  (
    g1244_p,
    n2003_inv_n_spl_,
    G1053_o2_n_spl_
  );


  or

  (
    g1244_n,
    n2003_inv_p_spl_0,
    G1053_o2_p_spl_0
  );


  and

  (
    g1245_p,
    n2003_inv_p_spl_0,
    G1053_o2_p_spl_0
  );


  or

  (
    g1245_n,
    n2003_inv_n_spl_,
    G1053_o2_n_spl_
  );


  and

  (
    g1246_p,
    g1245_n,
    g1244_n
  );


  or

  (
    g1246_n,
    g1245_p,
    g1244_p
  );


  or

  (
    g1247_n,
    g1246_n,
    g1243_p
  );


  or

  (
    g1248_n,
    g1246_p,
    g1243_n
  );


  and

  (
    g1249_p,
    g1248_n,
    g1247_n
  );


  and

  (
    g1250_p,
    g1231_p,
    g1228_n_spl_0
  );


  and

  (
    g1251_p,
    g1231_n_spl_0,
    g1228_p
  );


  or

  (
    g1252_n,
    g1251_p,
    g1250_p
  );


  and

  (
    g1253_p,
    n3198_lo_buf_o2_p_spl_,
    n3186_lo_buf_o2_n_spl_
  );


  or

  (
    g1253_n,
    n3198_lo_buf_o2_n_spl_,
    n3186_lo_buf_o2_p_spl_
  );


  and

  (
    g1254_p,
    n3198_lo_buf_o2_n_spl_,
    n3186_lo_buf_o2_p_spl_
  );


  or

  (
    g1254_n,
    n3198_lo_buf_o2_p_spl_,
    n3186_lo_buf_o2_n_spl_
  );


  and

  (
    g1255_p,
    g1254_n,
    g1253_n
  );


  or

  (
    g1255_n,
    g1254_p,
    g1253_p
  );


  and

  (
    g1256_p,
    n3222_lo_buf_o2_p_spl_,
    n3210_lo_buf_o2_n_spl_
  );


  or

  (
    g1256_n,
    n3222_lo_buf_o2_n_spl_,
    n3210_lo_buf_o2_p_spl_
  );


  and

  (
    g1257_p,
    n3222_lo_buf_o2_n_spl_,
    n3210_lo_buf_o2_p_spl_
  );


  or

  (
    g1257_n,
    n3222_lo_buf_o2_p_spl_,
    n3210_lo_buf_o2_n_spl_
  );


  and

  (
    g1258_p,
    g1257_n,
    g1256_n
  );


  or

  (
    g1258_n,
    g1257_p,
    g1256_p
  );


  and

  (
    g1259_p,
    G402_o2_n,
    n3246_lo_buf_o2_p
  );


  or

  (
    g1259_n,
    G402_o2_p,
    n3246_lo_buf_o2_n
  );


  and

  (
    g1260_p,
    G403_o2_n,
    n3234_lo_buf_o2_p
  );


  or

  (
    g1260_n,
    G403_o2_p,
    n3234_lo_buf_o2_n
  );


  and

  (
    g1261_p,
    g1260_n,
    g1259_n
  );


  or

  (
    g1261_n,
    g1260_p,
    g1259_p
  );


  or

  (
    g1262_n,
    g1258_n_spl_,
    g1255_p_spl_
  );


  or

  (
    g1263_n,
    g1262_n,
    g1261_p_spl_
  );


  or

  (
    g1264_n,
    g1258_n_spl_,
    g1255_n_spl_
  );


  or

  (
    g1265_n,
    g1264_n,
    g1261_n_spl_
  );


  and

  (
    g1266_p,
    g1265_n,
    g1263_n
  );


  or

  (
    g1267_n,
    g1258_p_spl_,
    g1255_n_spl_
  );


  or

  (
    g1268_n,
    g1267_n,
    g1261_p_spl_
  );


  or

  (
    g1269_n,
    g1258_p_spl_,
    g1255_p_spl_
  );


  or

  (
    g1270_n,
    g1269_n,
    g1261_n_spl_
  );


  and

  (
    g1271_p,
    g1270_n,
    g1268_n
  );


  and

  (
    g1272_p,
    g1271_p,
    g1266_p
  );


  and

  (
    g1273_p,
    G1079_o2_p_spl_,
    G1222_o2_p_spl_
  );


  or

  (
    g1273_n,
    G1079_o2_n_spl_,
    G1222_o2_n_spl_
  );


  and

  (
    g1274_p,
    G1079_o2_n_spl_,
    G1222_o2_n_spl_
  );


  or

  (
    g1274_n,
    G1079_o2_p_spl_,
    G1222_o2_p_spl_
  );


  and

  (
    g1275_p,
    g1274_n,
    g1273_n
  );


  or

  (
    g1275_n,
    g1274_p,
    g1273_p
  );


  and

  (
    g1276_p,
    G1228_o2_n_spl_,
    G1225_o2_p_spl_
  );


  or

  (
    g1276_n,
    G1228_o2_p_spl_,
    G1225_o2_n_spl_
  );


  and

  (
    g1277_p,
    G1228_o2_p_spl_,
    G1225_o2_n_spl_
  );


  or

  (
    g1277_n,
    G1228_o2_n_spl_,
    G1225_o2_p_spl_
  );


  and

  (
    g1278_p,
    g1277_n,
    g1276_n
  );


  or

  (
    g1278_n,
    g1277_p,
    g1276_p
  );


  and

  (
    g1279_p,
    G1364_o2_p,
    G1234_o2_n
  );


  or

  (
    g1279_n,
    G1364_o2_n,
    G1234_o2_p
  );


  and

  (
    g1280_p,
    G1365_o2_p,
    G1231_o2_n
  );


  or

  (
    g1280_n,
    G1365_o2_n,
    G1231_o2_p
  );


  and

  (
    g1281_p,
    g1280_n,
    g1279_n
  );


  or

  (
    g1281_n,
    g1280_p,
    g1279_p
  );


  and

  (
    g1282_p,
    g1278_p_spl_,
    g1275_n_spl_
  );


  and

  (
    g1283_p,
    g1282_p,
    g1281_n_spl_
  );


  and

  (
    g1284_p,
    g1278_p_spl_,
    g1275_p_spl_
  );


  and

  (
    g1285_p,
    g1284_p,
    g1281_p_spl_
  );


  or

  (
    g1286_n,
    g1285_p,
    g1283_p
  );


  and

  (
    g1287_p,
    g1278_n_spl_,
    g1275_p_spl_
  );


  and

  (
    g1288_p,
    g1287_p,
    g1281_n_spl_
  );


  and

  (
    g1289_p,
    g1278_n_spl_,
    g1275_n_spl_
  );


  and

  (
    g1290_p,
    g1289_p,
    g1281_p_spl_
  );


  or

  (
    g1291_n,
    g1290_p,
    g1288_p
  );


  or

  (
    g1292_n,
    g1291_n,
    g1286_n
  );


  and

  (
    g1293_p,
    G1371_o2_p_spl_,
    G1368_o2_n_spl_
  );


  or

  (
    g1293_n,
    G1371_o2_n_spl_,
    G1368_o2_p_spl_
  );


  and

  (
    g1294_p,
    G1371_o2_n_spl_,
    G1368_o2_p_spl_
  );


  or

  (
    g1294_n,
    G1371_o2_p_spl_,
    G1368_o2_n_spl_
  );


  and

  (
    g1295_p,
    g1294_n,
    g1293_n
  );


  or

  (
    g1295_n,
    g1294_p,
    g1293_p
  );


  and

  (
    g1296_p,
    G1537_o2_p_spl_,
    G1374_o2_p_spl_
  );


  or

  (
    g1296_n,
    G1537_o2_n_spl_,
    G1374_o2_n_spl_
  );


  and

  (
    g1297_p,
    G1537_o2_n_spl_,
    G1374_o2_n_spl_
  );


  or

  (
    g1297_n,
    G1537_o2_p_spl_,
    G1374_o2_p_spl_
  );


  and

  (
    g1298_p,
    g1297_n,
    g1296_n
  );


  or

  (
    g1298_n,
    g1297_p,
    g1296_p
  );


  and

  (
    g1299_p,
    G1478_o2_n,
    G1540_o2_n
  );


  or

  (
    g1299_n,
    G1478_o2_p,
    G1540_o2_p
  );


  and

  (
    g1300_p,
    G1653_o2_p,
    G1377_o2_p
  );


  or

  (
    g1300_n,
    G1653_o2_n,
    G1377_o2_n
  );


  and

  (
    g1301_p,
    g1300_n,
    g1299_n
  );


  or

  (
    g1301_n,
    g1300_p,
    g1299_p
  );


  or

  (
    g1302_n,
    g1298_n_spl_,
    g1295_p_spl_
  );


  or

  (
    g1303_n,
    g1302_n,
    g1301_p_spl_
  );


  or

  (
    g1304_n,
    g1298_n_spl_,
    g1295_n_spl_
  );


  or

  (
    g1305_n,
    g1304_n,
    g1301_n_spl_
  );


  and

  (
    g1306_p,
    g1305_n,
    g1303_n
  );


  or

  (
    g1307_n,
    g1298_p_spl_,
    g1295_n_spl_
  );


  or

  (
    g1308_n,
    g1307_n,
    g1301_p_spl_
  );


  or

  (
    g1309_n,
    g1298_p_spl_,
    g1295_p_spl_
  );


  or

  (
    g1310_n,
    g1309_n,
    g1301_n_spl_
  );


  and

  (
    g1311_p,
    g1310_n,
    g1308_n
  );


  and

  (
    g1312_p,
    g1311_p,
    g1306_p
  );


  and

  (
    g1313_p,
    G1636_o2_p_spl_001,
    n3087_lo_n_spl_
  );


  and

  (
    g1314_p,
    G1636_o2_n_spl_001,
    n2955_lo_n_spl_
  );


  or

  (
    g1315_n,
    g1314_p,
    g1313_p
  );


  or

  (
    g1316_n,
    G1636_o2_p_spl_001,
    n2991_lo_p_spl_0
  );


  or

  (
    g1317_n,
    g1316_n,
    n1503_lo_buf_o2_n_spl_000
  );


  or

  (
    g1318_n,
    G1636_o2_p_spl_010,
    n3003_lo_p_spl_0
  );


  or

  (
    g1319_n,
    g1318_n,
    n1503_lo_buf_o2_n_spl_000
  );


  and

  (
    g1320_p,
    G1684_o2_p_spl_001,
    n3087_lo_n_spl_
  );


  and

  (
    g1321_p,
    G1684_o2_n_spl_001,
    n2955_lo_n_spl_
  );


  or

  (
    g1322_n,
    g1321_p,
    g1320_p
  );


  or

  (
    g1323_n,
    G1684_o2_p_spl_001,
    n2991_lo_p_spl_0
  );


  or

  (
    g1324_n,
    g1323_n,
    n1503_lo_buf_o2_n_spl_001
  );


  or

  (
    g1325_n,
    G1684_o2_p_spl_010,
    n3003_lo_p_spl_0
  );


  or

  (
    g1326_n,
    g1325_n,
    n1503_lo_buf_o2_n_spl_001
  );


  or

  (
    g1327_n,
    G1636_o2_p_spl_010,
    n3063_lo_buf_o2_p_spl_00
  );


  and

  (
    g1328_p,
    G1193_o2_n,
    n1770_lo_buf_o2_p
  );


  or

  (
    g1328_n,
    G1193_o2_p,
    n1770_lo_buf_o2_n
  );


  and

  (
    g1329_p,
    g1328_p,
    G1320_o2_n
  );


  or

  (
    g1329_n,
    g1328_n,
    G1320_o2_p
  );


  or

  (
    g1330_n,
    g1329_n_spl_0,
    g1327_n
  );


  or

  (
    g1331_n,
    G1684_o2_p_spl_010,
    n3063_lo_buf_o2_p_spl_00
  );


  or

  (
    g1332_n,
    g1331_n,
    g1329_n_spl_0
  );


  and

  (
    g1333_p,
    G1636_o2_n_spl_001,
    n3027_lo_n_spl_
  );


  and

  (
    g1334_p,
    g1333_p,
    g1329_p_spl_00
  );


  and

  (
    g1335_p,
    G1636_o2_n_spl_010,
    n3039_lo_n_spl_
  );


  and

  (
    g1336_p,
    g1335_p,
    g1329_p_spl_00
  );


  and

  (
    g1337_p,
    G1684_o2_n_spl_001,
    n3027_lo_n_spl_
  );


  and

  (
    g1338_p,
    g1337_p,
    g1329_p_spl_01
  );


  and

  (
    g1339_p,
    G1684_o2_n_spl_010,
    n3039_lo_n_spl_
  );


  and

  (
    g1340_p,
    g1339_p,
    g1329_p_spl_01
  );


  or

  (
    g1341_n,
    G1636_o2_n_spl_010,
    n3099_lo_buf_o2_p_spl_0
  );


  or

  (
    g1342_n,
    G1636_o2_p_spl_01,
    n2967_lo_buf_o2_p_spl_0
  );


  and

  (
    g1343_p,
    g1342_n,
    g1341_n
  );


  or

  (
    g1344_n,
    g1343_p,
    n1503_lo_buf_o2_n_spl_010
  );


  or

  (
    g1345_n,
    G1636_o2_n_spl_01,
    n3111_lo_buf_o2_p_spl_0
  );


  or

  (
    g1346_n,
    G1636_o2_p_spl_10,
    n2979_lo_buf_o2_p_spl_0
  );


  and

  (
    g1347_p,
    g1346_n,
    g1345_n
  );


  or

  (
    g1348_n,
    g1347_p,
    n1503_lo_buf_o2_n_spl_010
  );


  or

  (
    g1349_n,
    G1684_o2_n_spl_010,
    n3099_lo_buf_o2_p_spl_0
  );


  or

  (
    g1350_n,
    G1684_o2_p_spl_01,
    n2967_lo_buf_o2_p_spl_0
  );


  and

  (
    g1351_p,
    g1350_n,
    g1349_n
  );


  or

  (
    g1352_n,
    g1351_p,
    n1503_lo_buf_o2_n_spl_011
  );


  or

  (
    g1353_n,
    G1684_o2_n_spl_01,
    n3111_lo_buf_o2_p_spl_0
  );


  or

  (
    g1354_n,
    G1684_o2_p_spl_10,
    n2979_lo_buf_o2_p_spl_0
  );


  and

  (
    g1355_p,
    g1354_n,
    g1353_n
  );


  or

  (
    g1356_n,
    g1355_p,
    n1503_lo_buf_o2_n_spl_011
  );


  or

  (
    g1357_n,
    g1020_n_spl_00,
    G1493_o2_n_spl_0
  );


  or

  (
    g1358_n,
    g1357_n,
    n1503_lo_buf_o2_n_spl_100
  );


  or

  (
    g1359_n,
    g1017_n_spl_00,
    G1493_o2_n_spl_0
  );


  or

  (
    g1360_n,
    g1359_n,
    n1503_lo_buf_o2_n_spl_100
  );


  or

  (
    g1361_n,
    g1020_n_spl_00,
    G1498_o2_n_spl_0
  );


  or

  (
    g1362_n,
    g1361_n,
    n1503_lo_buf_o2_n_spl_101
  );


  or

  (
    g1363_n,
    g1017_n_spl_00,
    G1498_o2_n_spl_0
  );


  or

  (
    g1364_n,
    g1363_n,
    n1503_lo_buf_o2_n_spl_101
  );


  and

  (
    g1365_p,
    g1045_n_spl_0,
    G1314_o2_n_spl_
  );


  and

  (
    g1366_p,
    g1365_p,
    g1329_p_spl_10
  );


  and

  (
    g1367_p,
    g1056_n_spl_0,
    G1314_o2_n_spl_
  );


  and

  (
    g1368_p,
    g1367_p,
    g1329_p_spl_10
  );


  or

  (
    g1369_n,
    g1023_n_spl_0,
    G1314_o2_p_spl_
  );


  or

  (
    g1370_n,
    g1369_n,
    g1329_n_spl_1
  );


  or

  (
    g1371_n,
    G1021_o2_p_spl_00,
    G1493_o2_n_spl_1
  );


  or

  (
    g1372_n,
    G1021_o2_p_spl_00,
    G1493_o2_p_spl_
  );


  and

  (
    g1373_p,
    g1372_n,
    g1371_n
  );


  or

  (
    g1374_n,
    g1373_p,
    n1503_lo_buf_o2_n_spl_110
  );


  or

  (
    g1375_n,
    G1026_o2_p_spl_00,
    G1493_o2_n_spl_1
  );


  or

  (
    g1376_n,
    G1026_o2_p_spl_00,
    G1493_o2_p_spl_
  );


  and

  (
    g1377_p,
    g1376_n,
    g1375_n
  );


  or

  (
    g1378_n,
    g1377_p,
    n1503_lo_buf_o2_n_spl_110
  );


  or

  (
    g1379_n,
    G1021_o2_p_spl_01,
    G1498_o2_n_spl_1
  );


  or

  (
    g1380_n,
    G1021_o2_p_spl_01,
    G1498_o2_p_spl_
  );


  and

  (
    g1381_p,
    g1380_n,
    g1379_n
  );


  or

  (
    g1382_n,
    g1381_p,
    n1503_lo_buf_o2_n_spl_111
  );


  or

  (
    g1383_n,
    G1026_o2_p_spl_01,
    G1498_o2_n_spl_1
  );


  or

  (
    g1384_n,
    G1026_o2_p_spl_01,
    G1498_o2_p_spl_
  );


  and

  (
    g1385_p,
    g1384_n,
    g1383_n
  );


  or

  (
    g1386_n,
    g1385_p,
    n1503_lo_buf_o2_n_spl_111
  );


  and

  (
    g1387_p,
    G1636_o2_n_spl_10,
    n3015_lo_n_spl_
  );


  and

  (
    g1388_p,
    g1387_p,
    g1329_p_spl_11
  );


  and

  (
    g1389_p,
    G1684_o2_n_spl_10,
    n3015_lo_n_spl_
  );


  and

  (
    g1390_p,
    g1389_p,
    g1329_p_spl_11
  );


  and

  (
    g1391_p,
    G707_o2_p_spl_10,
    n2739_lo_p
  );


  and

  (
    g1392_p,
    g1391_p,
    G718_o2_p_spl_10
  );


  and

  (
    g1393_p,
    G405_o2_n_spl_10,
    n2379_lo_p
  );


  and

  (
    g1394_p,
    g1393_p,
    G718_o2_p_spl_10
  );


  and

  (
    g1395_p,
    G707_o2_p_spl_10,
    n2619_lo_p
  );


  and

  (
    g1396_p,
    g1395_p,
    G417_o2_n_spl_10
  );


  and

  (
    g1397_p,
    G405_o2_n_spl_10,
    n2499_lo_p
  );


  and

  (
    g1398_p,
    g1397_p,
    G417_o2_n_spl_10
  );


  or

  (
    g1399_n,
    g1394_p,
    g1392_p
  );


  or

  (
    g1400_n,
    g1399_n,
    g1396_p
  );


  or

  (
    g1401_n,
    g1400_n,
    g1398_p
  );


  and

  (
    g1402_p,
    G603_o2_p_spl_10,
    n2163_lo_p
  );


  and

  (
    g1403_p,
    g1402_p,
    G614_o2_p_spl_10
  );


  and

  (
    g1404_p,
    G301_o2_n_spl_10,
    n1779_lo_p
  );


  and

  (
    g1405_p,
    g1404_p,
    G614_o2_p_spl_10
  );


  and

  (
    g1406_p,
    G603_o2_p_spl_10,
    n1911_lo_p
  );


  and

  (
    g1407_p,
    g1406_p,
    G313_o2_n_spl_10
  );


  and

  (
    g1408_p,
    G301_o2_n_spl_10,
    n2031_lo_p
  );


  and

  (
    g1409_p,
    g1408_p,
    G313_o2_n_spl_10
  );


  or

  (
    g1410_n,
    g1405_p,
    g1403_p
  );


  or

  (
    g1411_n,
    g1410_n,
    g1407_p
  );


  or

  (
    g1412_n,
    g1411_n,
    g1409_p
  );


  and

  (
    g1413_p,
    G603_o2_p_spl_11,
    n2283_lo_p
  );


  and

  (
    g1414_p,
    g1413_p,
    G614_o2_p_spl_11
  );


  and

  (
    g1415_p,
    G301_o2_n_spl_11,
    n1899_lo_p
  );


  and

  (
    g1416_p,
    g1415_p,
    G614_o2_p_spl_11
  );


  and

  (
    g1417_p,
    G603_o2_p_spl_11,
    n2019_lo_p
  );


  and

  (
    g1418_p,
    g1417_p,
    G313_o2_n_spl_11
  );


  and

  (
    g1419_p,
    G301_o2_n_spl_11,
    n2151_lo_p
  );


  and

  (
    g1420_p,
    g1419_p,
    G313_o2_n_spl_11
  );


  or

  (
    g1421_n,
    g1416_p,
    g1414_p
  );


  or

  (
    g1422_n,
    g1421_n,
    g1418_p
  );


  or

  (
    g1423_n,
    g1422_n,
    g1420_p
  );


  or

  (
    g1424_n,
    g1034_n_spl_0,
    G1314_o2_p_spl_
  );


  or

  (
    g1425_n,
    g1424_n,
    g1329_n_spl_1
  );


  and

  (
    g1426_p,
    n3150_lo_buf_o2_p_spl_000,
    n2712_lo_buf_o2_p
  );


  and

  (
    g1427_p,
    g1426_p,
    n3162_lo_buf_o2_p_spl_000
  );


  and

  (
    g1428_p,
    n3150_lo_buf_o2_n_spl_00,
    n2352_lo_buf_o2_p
  );


  and

  (
    g1429_p,
    g1428_p,
    n3162_lo_buf_o2_p_spl_000
  );


  and

  (
    g1430_p,
    n3150_lo_buf_o2_p_spl_000,
    n2592_lo_buf_o2_p
  );


  and

  (
    g1431_p,
    g1430_p,
    n3162_lo_buf_o2_n_spl_00
  );


  and

  (
    g1432_p,
    n3150_lo_buf_o2_n_spl_00,
    n2472_lo_buf_o2_p
  );


  and

  (
    g1433_p,
    g1432_p,
    n3162_lo_buf_o2_n_spl_00
  );


  or

  (
    g1434_n,
    g1429_p,
    g1427_p
  );


  or

  (
    g1435_n,
    g1434_n,
    g1431_p
  );


  or

  (
    g1436_n,
    g1435_n,
    g1433_p
  );


  or

  (
    g1437_n,
    n3150_lo_buf_o2_n_spl_01,
    n2724_lo_buf_o2_n
  );


  or

  (
    g1438_n,
    g1437_n,
    n3162_lo_buf_o2_n_spl_01
  );


  or

  (
    g1439_n,
    n3150_lo_buf_o2_p_spl_001,
    n2364_lo_buf_o2_n
  );


  or

  (
    g1440_n,
    g1439_n,
    n3162_lo_buf_o2_n_spl_01
  );


  or

  (
    g1441_n,
    n3150_lo_buf_o2_n_spl_01,
    n2604_lo_buf_o2_n
  );


  or

  (
    g1442_n,
    g1441_n,
    n3162_lo_buf_o2_p_spl_001
  );


  or

  (
    g1443_n,
    n3150_lo_buf_o2_p_spl_001,
    n2484_lo_buf_o2_n
  );


  or

  (
    g1444_n,
    g1443_n,
    n3162_lo_buf_o2_p_spl_001
  );


  and

  (
    g1445_p,
    g1440_n,
    g1438_n
  );


  and

  (
    g1446_p,
    g1445_p,
    g1442_n
  );


  and

  (
    g1447_p,
    g1446_p,
    g1444_n
  );


  and

  (
    g1448_p,
    n2958_lo_buf_o2_n_spl_,
    n2970_lo_buf_o2_p_spl_
  );


  or

  (
    g1448_n,
    n2958_lo_buf_o2_p_spl_,
    n2970_lo_buf_o2_n_spl_
  );


  and

  (
    g1449_p,
    n2958_lo_buf_o2_p_spl_,
    n2970_lo_buf_o2_n_spl_
  );


  or

  (
    g1449_n,
    n2958_lo_buf_o2_n_spl_,
    n2970_lo_buf_o2_p_spl_
  );


  and

  (
    g1450_p,
    g1449_n,
    g1448_n
  );


  or

  (
    g1450_n,
    g1449_p,
    g1448_p
  );


  and

  (
    g1451_p,
    n2946_lo_buf_o2_p_spl_,
    n3282_lo_p_spl_
  );


  or

  (
    g1451_n,
    n2946_lo_buf_o2_n_spl_,
    n3282_lo_n_spl_
  );


  and

  (
    g1452_p,
    n2946_lo_buf_o2_n_spl_,
    n3282_lo_n_spl_
  );


  or

  (
    g1452_n,
    n2946_lo_buf_o2_p_spl_,
    n3282_lo_p_spl_
  );


  and

  (
    g1453_p,
    g1452_n,
    g1451_n
  );


  or

  (
    g1453_n,
    g1452_p,
    g1451_p
  );


  and

  (
    g1454_p,
    n2994_lo_buf_o2_p,
    n2982_lo_buf_o2_n
  );


  and

  (
    g1455_p,
    n2994_lo_buf_o2_n,
    n2982_lo_buf_o2_p
  );


  or

  (
    g1456_n,
    g1455_p,
    g1454_p
  );


  or

  (
    g1457_n,
    g1453_p_spl_,
    g1450_p_spl_
  );


  or

  (
    g1458_n,
    g1457_n,
    g1456_n_spl_0
  );


  and

  (
    g1459_p,
    g1453_n_spl_,
    g1450_p_spl_
  );


  and

  (
    g1460_p,
    g1459_p,
    g1456_n_spl_0
  );


  and

  (
    g1461_p,
    n3090_lo_buf_o2_p_spl_0,
    n3078_lo_buf_o2_n_spl_
  );


  or

  (
    g1461_n,
    n3090_lo_buf_o2_n_spl_,
    n3078_lo_buf_o2_p_spl_0
  );


  and

  (
    g1462_p,
    n3090_lo_buf_o2_n_spl_,
    n3078_lo_buf_o2_p_spl_0
  );


  or

  (
    g1462_n,
    n3090_lo_buf_o2_p_spl_0,
    n3078_lo_buf_o2_n_spl_
  );


  and

  (
    g1463_p,
    g1462_n,
    g1461_n
  );


  or

  (
    g1463_n,
    g1462_p,
    g1461_p
  );


  and

  (
    g1464_p,
    n3066_lo_buf_o2_p_spl_,
    n3294_lo_p_spl_
  );


  or

  (
    g1464_n,
    n3066_lo_buf_o2_n_spl_,
    n3294_lo_n_spl_
  );


  and

  (
    g1465_p,
    n3066_lo_buf_o2_n_spl_,
    n3294_lo_n_spl_
  );


  or

  (
    g1465_n,
    n3066_lo_buf_o2_p_spl_,
    n3294_lo_p_spl_
  );


  and

  (
    g1466_p,
    g1465_n,
    g1464_n
  );


  or

  (
    g1466_n,
    g1465_p,
    g1464_p
  );


  and

  (
    g1467_p,
    n3114_lo_buf_o2_p_spl_,
    n3102_lo_buf_o2_n
  );


  and

  (
    g1468_p,
    n3114_lo_buf_o2_n,
    n3102_lo_buf_o2_p_spl_
  );


  or

  (
    g1469_n,
    g1468_p,
    g1467_p
  );


  or

  (
    g1470_n,
    g1466_p_spl_,
    g1463_p_spl_
  );


  or

  (
    g1471_n,
    g1470_n,
    g1469_n_spl_0
  );


  and

  (
    g1472_p,
    g1466_n_spl_,
    g1463_p_spl_
  );


  and

  (
    g1473_p,
    g1472_p,
    g1469_n_spl_0
  );


  and

  (
    g1474_p,
    g1453_p_spl_,
    g1450_n_spl_
  );


  and

  (
    g1475_p,
    g1474_p,
    g1456_n_spl_1
  );


  and

  (
    g1476_p,
    g1466_p_spl_,
    g1463_n_spl_
  );


  and

  (
    g1477_p,
    g1476_p,
    g1469_n_spl_1
  );


  and

  (
    g1478_p,
    G1129_o2_p_spl_,
    G1132_o2_n_spl_
  );


  or

  (
    g1478_n,
    G1129_o2_n_spl_,
    G1132_o2_p_spl_
  );


  and

  (
    g1479_p,
    G1129_o2_n_spl_,
    G1132_o2_p_spl_
  );


  or

  (
    g1479_n,
    G1129_o2_p_spl_,
    G1132_o2_n_spl_
  );


  and

  (
    g1480_p,
    g1479_n,
    g1478_n
  );


  or

  (
    g1480_n,
    g1479_p,
    g1478_p
  );


  and

  (
    g1481_p,
    G1329_o2_p_spl_,
    G1137_o2_p
  );


  and

  (
    g1482_p,
    G1329_o2_n_spl_,
    G1137_o2_n
  );


  or

  (
    g1483_n,
    g1482_p,
    g1481_p
  );


  or

  (
    g1484_n,
    g1480_p_spl_,
    g1014_n_spl_0
  );


  or

  (
    g1485_n,
    g1484_n,
    g1483_n_spl_0
  );


  and

  (
    g1486_p,
    g1480_n_spl_,
    g1014_n_spl_0
  );


  and

  (
    g1487_p,
    g1486_p,
    g1483_n_spl_0
  );


  and

  (
    g1488_p,
    g1480_p_spl_,
    g1014_p_spl_
  );


  and

  (
    g1489_p,
    g1488_p,
    g1483_n_spl_1
  );


  or

  (
    g1490_n,
    g1453_n_spl_,
    g1450_n_spl_
  );


  or

  (
    g1491_n,
    g1490_n,
    g1456_n_spl_1
  );


  or

  (
    g1492_n,
    g1466_n_spl_,
    g1463_n_spl_
  );


  or

  (
    g1493_n,
    g1492_n,
    g1469_n_spl_1
  );


  or

  (
    g1494_n,
    g1480_n_spl_,
    g1014_p_spl_
  );


  or

  (
    g1495_n,
    g1494_n,
    g1483_n_spl_1
  );


  and

  (
    g1496_p,
    n1554_lo_p_spl_000,
    n1458_lo_p
  );


  and

  (
    g1497_p,
    G1008_o2_p_spl_0,
    n1554_lo_n_spl_000
  );


  or

  (
    g1498_n,
    g1497_p,
    g1496_p
  );


  and

  (
    g1499_p,
    n1554_lo_p_spl_000,
    n1470_lo_p
  );


  and

  (
    g1500_p,
    G1017_o2_p_spl_,
    n1554_lo_n_spl_000
  );


  or

  (
    g1501_n,
    g1500_p,
    g1499_p
  );


  and

  (
    g1502_p,
    n1554_lo_p_spl_00,
    n1482_lo_p
  );


  and

  (
    g1503_p,
    G1033_o2_p,
    n1554_lo_n_spl_00
  );


  or

  (
    g1504_n,
    g1503_p,
    g1502_p
  );


  and

  (
    g1505_p,
    n1566_lo_p,
    n1554_lo_p_spl_01
  );


  and

  (
    g1506_p,
    G1002_o2_p_spl_0,
    n1554_lo_n_spl_01
  );


  or

  (
    g1507_n,
    g1506_p,
    g1505_p
  );


  and

  (
    g1508_p,
    n1578_lo_p,
    n1554_lo_p_spl_01
  );


  and

  (
    g1509_p,
    G1014_o2_p,
    n1554_lo_n_spl_01
  );


  or

  (
    g1510_n,
    g1509_p,
    g1508_p
  );


  and

  (
    g1511_p,
    n1590_lo_p,
    n1554_lo_p_spl_10
  );


  and

  (
    g1512_p,
    n5554_o2_p_spl_,
    n1554_lo_n_spl_10
  );


  or

  (
    g1513_n,
    g1512_p,
    g1511_p
  );


  and

  (
    g1514_p,
    n1602_lo_p,
    n1554_lo_p_spl_10
  );


  and

  (
    g1515_p,
    n5553_o2_p_spl_,
    n1554_lo_n_spl_10
  );


  or

  (
    g1516_n,
    g1515_p,
    g1514_p
  );


  and

  (
    g1517_p,
    n1614_lo_p,
    n1554_lo_p_spl_11
  );


  and

  (
    g1518_p,
    G1030_o2_p,
    n1554_lo_n_spl_11
  );


  or

  (
    g1519_n,
    g1518_p,
    g1517_p
  );


  and

  (
    g1520_p,
    n1626_lo_p,
    n1554_lo_p_spl_11
  );


  and

  (
    g1521_p,
    G1036_o2_p,
    n1554_lo_n_spl_11
  );


  or

  (
    g1522_n,
    g1521_p,
    g1520_p
  );


  and

  (
    g1523_p,
    n1686_lo_p_spl_000,
    n1638_lo_p
  );


  and

  (
    g1524_p,
    G1062_o2_p,
    n1686_lo_n_spl_00
  );


  or

  (
    g1525_n,
    g1524_p,
    g1523_p
  );


  and

  (
    g1526_p,
    n1686_lo_p_spl_000,
    n1650_lo_p
  );


  and

  (
    g1527_p,
    G1072_o2_p,
    n1686_lo_n_spl_00
  );


  or

  (
    g1528_n,
    g1527_p,
    g1526_p
  );


  and

  (
    g1529_p,
    n1686_lo_p_spl_00,
    n1662_lo_p
  );


  and

  (
    g1530_p,
    n5223_o2_p_spl_,
    n1686_lo_n_spl_01
  );


  or

  (
    g1531_n,
    g1530_p,
    g1529_p
  );


  and

  (
    g1532_p,
    n1698_lo_p,
    n1686_lo_p_spl_01
  );


  and

  (
    g1533_p,
    G1067_o2_p,
    n1686_lo_n_spl_01
  );


  or

  (
    g1534_n,
    g1533_p,
    g1532_p
  );


  and

  (
    g1535_p,
    n1710_lo_p,
    n1686_lo_p_spl_01
  );


  and

  (
    g1536_p,
    G1076_o2_p,
    n1686_lo_n_spl_10
  );


  or

  (
    g1537_n,
    g1536_p,
    g1535_p
  );


  and

  (
    g1538_p,
    n1722_lo_p,
    n1686_lo_p_spl_10
  );


  and

  (
    g1539_p,
    n5222_o2_p_spl_1,
    n1686_lo_n_spl_10
  );


  or

  (
    g1540_n,
    g1539_p,
    g1538_p
  );


  and

  (
    g1541_p,
    n1734_lo_p,
    n1686_lo_p_spl_10
  );


  and

  (
    g1542_p,
    G1049_o2_p_spl_1,
    n1686_lo_n_spl_1
  );


  or

  (
    g1543_n,
    g1542_p,
    g1541_p
  );


  or

  (
    g1544_n,
    G1002_o2_p_spl_0,
    G1008_o2_p_spl_1
  );


  or

  (
    g1545_n,
    G1002_o2_n,
    G1008_o2_n_spl_
  );


  and

  (
    g1546_p,
    g1545_n,
    g1544_n
  );


  and

  (
    g1547_p,
    g1219_n_spl_,
    g1157_n_spl_
  );


  or

  (
    g1548_n,
    g1447_p_spl_,
    n2928_lo_p
  );


  or

  (
    g1549_n,
    g1548_n_spl_,
    g1436_n_spl_0
  );


  or

  (
    g1550_n,
    g1549_n,
    n1764_lo_n
  );


  and

  (
    g1551_p,
    G1636_o2_p_spl_10,
    n3063_lo_buf_o2_n_spl_
  );


  or

  (
    g1551_n,
    G1636_o2_n_spl_10,
    n3063_lo_buf_o2_p_spl_01
  );


  and

  (
    g1552_p,
    G1636_o2_n_spl_11,
    n2919_lo_buf_o2_n_spl_
  );


  or

  (
    g1552_n,
    G1636_o2_p_spl_11,
    n2919_lo_buf_o2_p_spl_0
  );


  and

  (
    g1553_p,
    g1552_n,
    g1551_n
  );


  or

  (
    g1553_n,
    g1552_p,
    g1551_p
  );


  or

  (
    g1554_n,
    g1553_p_spl_,
    g1089_n_spl_00
  );


  and

  (
    g1555_p,
    G1684_o2_p_spl_10,
    n3063_lo_buf_o2_n_spl_
  );


  or

  (
    g1555_n,
    G1684_o2_n_spl_10,
    n3063_lo_buf_o2_p_spl_01
  );


  and

  (
    g1556_p,
    G1684_o2_n_spl_11,
    n2919_lo_buf_o2_n_spl_
  );


  or

  (
    g1556_n,
    G1684_o2_p_spl_11,
    n2919_lo_buf_o2_p_spl_0
  );


  and

  (
    g1557_p,
    g1556_n,
    g1555_n
  );


  or

  (
    g1557_n,
    g1556_p,
    g1555_p
  );


  or

  (
    g1558_n,
    g1557_p_spl_,
    g1089_n_spl_00
  );


  or

  (
    g1559_n,
    g1315_n_spl_0,
    g1078_p_spl_0
  );


  and

  (
    g1560_p,
    g1358_n_spl_0,
    g1317_n_spl_0
  );


  and

  (
    g1561_p,
    g1360_n_spl_0,
    g1319_n_spl_0
  );


  or

  (
    g1562_n,
    g1322_n_spl_0,
    g1078_p_spl_0
  );


  and

  (
    g1563_p,
    g1362_n_spl_0,
    g1324_n_spl_0
  );


  and

  (
    g1564_p,
    g1364_n_spl_0,
    g1326_n_spl_0
  );


  and

  (
    g1565_p,
    g1370_n_spl_00,
    g1330_n_spl_0
  );


  and

  (
    g1566_p,
    g1370_n_spl_00,
    g1332_n_spl_0
  );


  or

  (
    g1567_n,
    g1366_p_spl_00,
    g1334_p_spl_0
  );


  or

  (
    g1568_n,
    g1368_p_spl_00,
    g1336_p_spl_0
  );


  or

  (
    g1569_n,
    g1366_p_spl_00,
    g1338_p_spl_0
  );


  or

  (
    g1570_n,
    g1368_p_spl_00,
    g1340_p_spl_0
  );


  and

  (
    g1571_p,
    g1374_n_spl_0,
    g1344_n_spl_0
  );


  and

  (
    g1572_p,
    g1378_n_spl_0,
    g1348_n_spl_0
  );


  and

  (
    g1573_p,
    g1382_n_spl_0,
    g1352_n_spl_0
  );


  and

  (
    g1574_p,
    g1386_n_spl_0,
    g1356_n_spl_0
  );


  or

  (
    g1575_n,
    g1358_n_spl_0,
    g1317_n_spl_0
  );


  or

  (
    g1576_n,
    g1360_n_spl_0,
    g1319_n_spl_0
  );


  or

  (
    g1577_n,
    g1362_n_spl_0,
    g1324_n_spl_0
  );


  or

  (
    g1578_n,
    g1364_n_spl_0,
    g1326_n_spl_0
  );


  and

  (
    g1579_p,
    g1366_p_spl_01,
    g1334_p_spl_0
  );


  and

  (
    g1580_p,
    g1368_p_spl_01,
    g1336_p_spl_0
  );


  or

  (
    g1581_n,
    g1370_n_spl_01,
    g1330_n_spl_0
  );


  and

  (
    g1582_p,
    g1366_p_spl_01,
    g1338_p_spl_0
  );


  and

  (
    g1583_p,
    g1368_p_spl_01,
    g1340_p_spl_0
  );


  or

  (
    g1584_n,
    g1370_n_spl_01,
    g1332_n_spl_0
  );


  and

  (
    g1585_p,
    g1315_n_spl_0,
    g1078_p_spl_1
  );


  and

  (
    g1586_p,
    g1322_n_spl_0,
    g1078_p_spl_1
  );


  or

  (
    g1587_n,
    g1374_n_spl_0,
    g1344_n_spl_0
  );


  or

  (
    g1588_n,
    g1378_n_spl_0,
    g1348_n_spl_0
  );


  or

  (
    g1589_n,
    g1382_n_spl_0,
    g1352_n_spl_0
  );


  or

  (
    g1590_n,
    g1386_n_spl_0,
    g1356_n_spl_0
  );


  and

  (
    g1591_p,
    G663_o2_p_spl_0,
    n2691_lo_p
  );


  and

  (
    g1592_p,
    g1591_p,
    G674_o2_p_spl_0
  );


  and

  (
    g1593_p,
    G374_o2_n_spl_0,
    n2331_lo_p
  );


  and

  (
    g1594_p,
    g1593_p,
    G674_o2_p_spl_0
  );


  and

  (
    g1595_p,
    G663_o2_p_spl_0,
    n2571_lo_p
  );


  and

  (
    g1596_p,
    g1595_p,
    G386_o2_n_spl_0
  );


  and

  (
    g1597_p,
    G374_o2_n_spl_0,
    n2451_lo_p
  );


  and

  (
    g1598_p,
    g1597_p,
    G386_o2_n_spl_0
  );


  or

  (
    g1599_n,
    g1594_p,
    g1592_p
  );


  or

  (
    g1600_n,
    g1599_n,
    g1596_p
  );


  or

  (
    g1601_n,
    g1600_n,
    g1598_p
  );


  and

  (
    g1602_p,
    G663_o2_p_spl_1,
    n2703_lo_p
  );


  and

  (
    g1603_p,
    g1602_p,
    G674_o2_p_spl_1
  );


  and

  (
    g1604_p,
    G374_o2_n_spl_1,
    n2343_lo_p
  );


  and

  (
    g1605_p,
    g1604_p,
    G674_o2_p_spl_1
  );


  and

  (
    g1606_p,
    G663_o2_p_spl_1,
    n2583_lo_p
  );


  and

  (
    g1607_p,
    g1606_p,
    G386_o2_n_spl_1
  );


  and

  (
    g1608_p,
    G374_o2_n_spl_1,
    n2463_lo_p
  );


  and

  (
    g1609_p,
    g1608_p,
    G386_o2_n_spl_1
  );


  or

  (
    g1610_n,
    g1605_p,
    g1603_p
  );


  or

  (
    g1611_n,
    g1610_n,
    g1607_p
  );


  or

  (
    g1612_n,
    g1611_n,
    g1609_p
  );


  or

  (
    g1613_n,
    G674_o2_n_spl_,
    G663_o2_n_spl_
  );


  or

  (
    g1614_n,
    G674_o2_n_spl_,
    G374_o2_p_spl_
  );


  or

  (
    g1615_n,
    G663_o2_n_spl_,
    G386_o2_p_spl_
  );


  or

  (
    g1616_n,
    G386_o2_p_spl_,
    G374_o2_p_spl_
  );


  and

  (
    g1617_p,
    g1614_n,
    g1613_n
  );


  and

  (
    g1618_p,
    g1617_p,
    g1615_n
  );


  and

  (
    g1619_p,
    g1618_p,
    g1616_n
  );


  and

  (
    g1620_p,
    G707_o2_p_spl_11,
    n2775_lo_p
  );


  and

  (
    g1621_p,
    g1620_p,
    G718_o2_p_spl_11
  );


  and

  (
    g1622_p,
    G405_o2_n_spl_11,
    n2415_lo_p
  );


  and

  (
    g1623_p,
    g1622_p,
    G718_o2_p_spl_11
  );


  and

  (
    g1624_p,
    G707_o2_p_spl_11,
    n2655_lo_p
  );


  and

  (
    g1625_p,
    g1624_p,
    G417_o2_n_spl_11
  );


  and

  (
    g1626_p,
    G405_o2_n_spl_11,
    n2535_lo_p
  );


  and

  (
    g1627_p,
    g1626_p,
    G417_o2_n_spl_11
  );


  or

  (
    g1628_n,
    g1623_p,
    g1621_p
  );


  or

  (
    g1629_n,
    g1628_n,
    g1625_p
  );


  or

  (
    g1630_n,
    g1629_n,
    g1627_p
  );


  and

  (
    g1631_p,
    g1553_n,
    g1089_n_spl_01
  );


  and

  (
    g1632_p,
    g1553_p_spl_,
    g1089_p_spl_
  );


  or

  (
    g1633_n,
    g1632_p,
    g1631_p
  );


  or

  (
    g1634_n,
    g1092_p_spl_,
    g1067_n_spl_00
  );


  or

  (
    g1635_n,
    g1092_n,
    g1067_p_spl_
  );


  and

  (
    g1636_p,
    g1635_n,
    g1634_n
  );


  and

  (
    g1637_p,
    g1557_n,
    g1089_n_spl_01
  );


  and

  (
    g1638_p,
    g1557_p_spl_,
    g1089_p_spl_
  );


  or

  (
    g1639_n,
    g1638_p,
    g1637_p
  );


  or

  (
    g1640_n,
    g1095_p_spl_,
    g1067_n_spl_00
  );


  or

  (
    g1641_n,
    g1095_n,
    g1067_p_spl_
  );


  and

  (
    g1642_p,
    g1641_n,
    g1640_n
  );


  or

  (
    g1643_n,
    G1636_o2_n_spl_11,
    n3039_lo_p_spl_0
  );


  or

  (
    g1644_n,
    G1636_o2_p_spl_11,
    n2907_lo_p_spl_0
  );


  and

  (
    g1645_p,
    g1644_n,
    g1643_n
  );


  or

  (
    g1646_n,
    g1645_p,
    g1412_n_spl_00
  );


  or

  (
    g1647_n,
    G1684_o2_n_spl_11,
    n3039_lo_p_spl_0
  );


  or

  (
    g1648_n,
    G1684_o2_p_spl_11,
    n2907_lo_p_spl_0
  );


  and

  (
    g1649_p,
    g1648_n,
    g1647_n
  );


  or

  (
    g1650_n,
    g1649_p,
    g1412_n_spl_00
  );


  and

  (
    g1651_p,
    n2808_lo_n_spl_00,
    n1812_lo_p
  );


  and

  (
    g1652_p,
    g1651_p,
    n2844_lo_p_spl_000
  );


  and

  (
    g1653_p,
    n2808_lo_n_spl_00,
    n1824_lo_p
  );


  and

  (
    g1654_p,
    g1653_p,
    n2844_lo_p_spl_000
  );


  and

  (
    g1655_p,
    n2808_lo_n_spl_01,
    n2064_lo_p
  );


  and

  (
    g1656_p,
    g1655_p,
    n2844_lo_n_spl_00
  );


  and

  (
    g1657_p,
    n2808_lo_n_spl_01,
    n2076_lo_p
  );


  and

  (
    g1658_p,
    g1657_p,
    n2844_lo_n_spl_00
  );


  and

  (
    g1659_p,
    n2808_lo_p_spl_000,
    n1944_lo_p
  );


  and

  (
    g1660_p,
    g1659_p,
    n2844_lo_n_spl_01
  );


  and

  (
    g1661_p,
    n2844_lo_n_spl_01,
    n2808_lo_p_spl_000
  );


  and

  (
    g1662_p,
    n3150_lo_buf_o2_n_spl_1,
    n2388_lo_p
  );


  and

  (
    g1663_p,
    g1662_p,
    n3162_lo_buf_o2_p_spl_01
  );


  and

  (
    g1664_p,
    n3150_lo_buf_o2_n_spl_1,
    n2508_lo_p
  );


  and

  (
    g1665_p,
    g1664_p,
    n3162_lo_buf_o2_n_spl_1
  );


  and

  (
    g1666_p,
    n3150_lo_buf_o2_p_spl_01,
    n2628_lo_p
  );


  and

  (
    g1667_p,
    g1666_p,
    n3162_lo_buf_o2_n_spl_1
  );


  and

  (
    g1668_p,
    n2808_lo_p_spl_001,
    n2196_lo_p
  );


  and

  (
    g1669_p,
    g1668_p,
    n2844_lo_p_spl_001
  );


  and

  (
    g1670_p,
    n2808_lo_p_spl_001,
    n2208_lo_p
  );


  and

  (
    g1671_p,
    g1670_p,
    n2844_lo_p_spl_001
  );


  and

  (
    g1672_p,
    n2808_lo_p_spl_010,
    n2220_lo_p
  );


  and

  (
    g1673_p,
    g1672_p,
    n2844_lo_p_spl_010
  );


  and

  (
    g1674_p,
    n2808_lo_n_spl_10,
    n1836_lo_p
  );


  and

  (
    g1675_p,
    g1674_p,
    n2844_lo_p_spl_010
  );


  and

  (
    g1676_p,
    n2808_lo_p_spl_010,
    n1956_lo_p
  );


  and

  (
    g1677_p,
    g1676_p,
    n2844_lo_n_spl_10
  );


  and

  (
    g1678_p,
    n2808_lo_n_spl_10,
    n2088_lo_p
  );


  and

  (
    g1679_p,
    g1678_p,
    n2844_lo_n_spl_10
  );


  or

  (
    g1680_n,
    g1675_p,
    g1673_p
  );


  or

  (
    g1681_n,
    g1680_n,
    g1677_p
  );


  or

  (
    g1682_n,
    g1681_n,
    g1679_p
  );


  and

  (
    g1683_p,
    n2808_lo_p_spl_011,
    n2232_lo_p
  );


  and

  (
    g1684_p,
    g1683_p,
    n2844_lo_p_spl_011
  );


  and

  (
    g1685_p,
    n2808_lo_n_spl_11,
    n1848_lo_p
  );


  and

  (
    g1686_p,
    g1685_p,
    n2844_lo_p_spl_011
  );


  and

  (
    g1687_p,
    n2808_lo_p_spl_011,
    n1968_lo_p
  );


  and

  (
    g1688_p,
    g1687_p,
    n2844_lo_n_spl_11
  );


  and

  (
    g1689_p,
    n2808_lo_n_spl_11,
    n2100_lo_p
  );


  and

  (
    g1690_p,
    g1689_p,
    n2844_lo_n_spl_11
  );


  or

  (
    g1691_n,
    g1686_p,
    g1684_p
  );


  or

  (
    g1692_n,
    g1691_n,
    g1688_p
  );


  or

  (
    g1693_n,
    g1692_n,
    g1690_p
  );


  and

  (
    g1694_p,
    n3150_lo_buf_o2_p_spl_01,
    n2748_lo_p
  );


  and

  (
    g1695_p,
    g1694_p,
    n3162_lo_buf_o2_p_spl_01
  );


  buf

  (
    G2531,
    n2793_lo_n_spl_0
  );


  buf

  (
    G2532,
    n2793_lo_n_spl_1
  );


  buf

  (
    G2533,
    n2793_lo_n_spl_1
  );


  buf

  (
    G2534,
    n2901_lo_n_spl_
  );


  buf

  (
    G2535,
    n2901_lo_n_spl_
  );


  buf

  (
    G2536,
    n3057_lo_n_spl_0
  );


  buf

  (
    G2537,
    n3057_lo_n_spl_0
  );


  buf

  (
    G2538,
    n3057_lo_n_spl_
  );


  buf

  (
    G2539,
    n1797_lo_n_spl_
  );


  buf

  (
    G2540,
    n2685_lo_n_spl_
  );


  buf

  (
    G2541,
    n2181_lo_n_spl_
  );


  buf

  (
    G2542,
    n2325_lo_n_spl_
  );


  buf

  (
    G2543,
    n2049_lo_n_spl_
  );


  buf

  (
    G2544,
    n2565_lo_n_spl_
  );


  buf

  (
    G2545,
    n1929_lo_n_spl_
  );


  buf

  (
    G2546,
    n2445_lo_n_spl_
  );


  buf

  (
    G2547,
    g837_n
  );


  buf

  (
    G2548,
    g839_n
  );


  buf

  (
    G2549,
    n2793_lo_p
  );


  buf

  (
    G2550,
    g840_p
  );


  buf

  (
    G2551,
    g841_n_spl_
  );


  buf

  (
    G2552,
    g842_n
  );


  buf

  (
    G2553,
    g843_n
  );


  buf

  (
    G2554,
    g850_n_spl_
  );


  buf

  (
    G2555,
    g850_n_spl_
  );


  buf

  (
    G2556,
    g853_n_spl_1
  );


  buf

  (
    G2557,
    n4537_o2_n
  );


  buf

  (
    G2558,
    n5478_o2_n
  );


  buf

  (
    G2559,
    n4538_o2_n
  );


  buf

  (
    G2560,
    n4710_o2_n
  );


  buf

  (
    G2561,
    n4711_o2_n_spl_
  );


  buf

  (
    G2562,
    n4927_o2_n
  );


  buf

  (
    G2563,
    g855_n
  );


  buf

  (
    G2564,
    g858_n
  );


  buf

  (
    G2565,
    g861_n
  );


  buf

  (
    G2566,
    n1232_inv_p_spl_
  );


  buf

  (
    G2567,
    n1235_inv_p_spl_
  );


  buf

  (
    G2568,
    n1214_inv_p
  );


  buf

  (
    G2569,
    n1211_inv_p
  );


  buf

  (
    G2570,
    n1220_inv_p
  );


  buf

  (
    G2571,
    n1217_inv_p
  );


  buf

  (
    G2572,
    n1229_inv_p
  );


  buf

  (
    G2573,
    g864_p_spl_
  );


  buf

  (
    G2574,
    g864_p_spl_
  );


  buf

  (
    G2575,
    g867_p_spl_
  );


  buf

  (
    G2576,
    g867_p_spl_
  );


  buf

  (
    G2577,
    g870_n
  );


  buf

  (
    G2578,
    g873_p_spl_
  );


  buf

  (
    G2579,
    g873_p_spl_
  );


  buf

  (
    G2580,
    g882_n
  );


  not

  (
    G2581,
    g886_p_spl_
  );


  buf

  (
    G2582,
    g895_p_spl_
  );


  buf

  (
    G2583,
    g904_p_spl_
  );


  buf

  (
    G2584,
    g975_n_spl_
  );


  buf

  (
    G2585,
    g975_n_spl_
  );


  buf

  (
    G2586,
    g984_n
  );


  not

  (
    G2587,
    g988_p_spl_
  );


  buf

  (
    G2588,
    g1000_p_spl_
  );


  buf

  (
    G2589,
    g1000_p_spl_
  );


  not

  (
    G2590,
    g1004_p_spl_
  );


  buf

  (
    G2591,
    n1448_inv_p
  );


  buf

  (
    G2592,
    g1007_n_spl_
  );


  buf

  (
    G2593,
    g1013_n_spl_
  );


  buf

  (
    G2594,
    g1013_n_spl_
  );


  buf

  (
    n1416_li,
    G1_p
  );


  buf

  (
    n1419_li,
    n1416_lo_p
  );


  buf

  (
    n1422_li,
    n1419_lo_p
  );


  buf

  (
    n1425_li,
    n1422_lo_p
  );


  buf

  (
    n1428_li,
    G2_p
  );


  buf

  (
    n1431_li,
    n1428_lo_p
  );


  buf

  (
    n1434_li,
    n1431_lo_p
  );


  buf

  (
    n1437_li,
    n1434_lo_p
  );


  buf

  (
    n1440_li,
    G3_p
  );


  buf

  (
    n1443_li,
    n1440_lo_p
  );


  buf

  (
    n1446_li,
    n1443_lo_p
  );


  buf

  (
    n1449_li,
    n1446_lo_p
  );


  buf

  (
    n1452_li,
    G4_p
  );


  buf

  (
    n1455_li,
    n1452_lo_p
  );


  buf

  (
    n1458_li,
    n1455_lo_p
  );


  buf

  (
    n1464_li,
    G5_p
  );


  buf

  (
    n1467_li,
    n1464_lo_p
  );


  buf

  (
    n1470_li,
    n1467_lo_p
  );


  buf

  (
    n1476_li,
    G6_p
  );


  buf

  (
    n1479_li,
    n1476_lo_p
  );


  buf

  (
    n1482_li,
    n1479_lo_p
  );


  buf

  (
    n1488_li,
    G7_p
  );


  buf

  (
    n1491_li,
    n1488_lo_p
  );


  buf

  (
    n1494_li,
    n1491_lo_p
  );


  buf

  (
    n1497_li,
    n1494_lo_p
  );


  buf

  (
    n1500_li,
    G8_p
  );


  buf

  (
    n1512_li,
    G9_p
  );


  buf

  (
    n1515_li,
    n1512_lo_p
  );


  buf

  (
    n1518_li,
    n1515_lo_p
  );


  buf

  (
    n1521_li,
    n1518_lo_p
  );


  buf

  (
    n1524_li,
    G10_p
  );


  buf

  (
    n1527_li,
    n1524_lo_p
  );


  buf

  (
    n1530_li,
    n1527_lo_p
  );


  buf

  (
    n1533_li,
    n1530_lo_p
  );


  buf

  (
    n1536_li,
    G11_p
  );


  buf

  (
    n1539_li,
    n1536_lo_p
  );


  buf

  (
    n1542_li,
    n1539_lo_p
  );


  buf

  (
    n1545_li,
    n1542_lo_p
  );


  buf

  (
    n1548_li,
    G12_p
  );


  buf

  (
    n1551_li,
    n1548_lo_p
  );


  buf

  (
    n1554_li,
    n1551_lo_p
  );


  buf

  (
    n1560_li,
    G13_p
  );


  buf

  (
    n1563_li,
    n1560_lo_p
  );


  buf

  (
    n1566_li,
    n1563_lo_p
  );


  buf

  (
    n1572_li,
    G14_p
  );


  buf

  (
    n1575_li,
    n1572_lo_p
  );


  buf

  (
    n1578_li,
    n1575_lo_p
  );


  buf

  (
    n1584_li,
    G15_p
  );


  buf

  (
    n1587_li,
    n1584_lo_p
  );


  buf

  (
    n1590_li,
    n1587_lo_p
  );


  buf

  (
    n1596_li,
    G16_p
  );


  buf

  (
    n1599_li,
    n1596_lo_p
  );


  buf

  (
    n1602_li,
    n1599_lo_p
  );


  buf

  (
    n1608_li,
    G17_p
  );


  buf

  (
    n1611_li,
    n1608_lo_p
  );


  buf

  (
    n1614_li,
    n1611_lo_p
  );


  buf

  (
    n1620_li,
    G18_p
  );


  buf

  (
    n1623_li,
    n1620_lo_p
  );


  buf

  (
    n1626_li,
    n1623_lo_p
  );


  buf

  (
    n1632_li,
    G19_p
  );


  buf

  (
    n1635_li,
    n1632_lo_p
  );


  buf

  (
    n1638_li,
    n1635_lo_p
  );


  buf

  (
    n1644_li,
    G20_p
  );


  buf

  (
    n1647_li,
    n1644_lo_p
  );


  buf

  (
    n1650_li,
    n1647_lo_p
  );


  buf

  (
    n1656_li,
    G21_p
  );


  buf

  (
    n1659_li,
    n1656_lo_p
  );


  buf

  (
    n1662_li,
    n1659_lo_p
  );


  buf

  (
    n1668_li,
    G22_p
  );


  buf

  (
    n1671_li,
    n1668_lo_p
  );


  buf

  (
    n1674_li,
    n1671_lo_p
  );


  buf

  (
    n1677_li,
    n1674_lo_p
  );


  buf

  (
    n1680_li,
    G23_p
  );


  buf

  (
    n1683_li,
    n1680_lo_p
  );


  buf

  (
    n1686_li,
    n1683_lo_p
  );


  buf

  (
    n1692_li,
    G24_p
  );


  buf

  (
    n1695_li,
    n1692_lo_p
  );


  buf

  (
    n1698_li,
    n1695_lo_p
  );


  buf

  (
    n1704_li,
    G25_p
  );


  buf

  (
    n1707_li,
    n1704_lo_p
  );


  buf

  (
    n1710_li,
    n1707_lo_p
  );


  buf

  (
    n1716_li,
    G26_p
  );


  buf

  (
    n1719_li,
    n1716_lo_p
  );


  buf

  (
    n1722_li,
    n1719_lo_p
  );


  buf

  (
    n1728_li,
    G27_p
  );


  buf

  (
    n1731_li,
    n1728_lo_p
  );


  buf

  (
    n1734_li,
    n1731_lo_p
  );


  buf

  (
    n1740_li,
    G28_p
  );


  buf

  (
    n1743_li,
    n1740_lo_p
  );


  buf

  (
    n1746_li,
    n1743_lo_p
  );


  buf

  (
    n1749_li,
    n1746_lo_p
  );


  buf

  (
    n1752_li,
    G29_p
  );


  buf

  (
    n1755_li,
    n1752_lo_p
  );


  buf

  (
    n1758_li,
    n1755_lo_p
  );


  buf

  (
    n1761_li,
    n1758_lo_p
  );


  buf

  (
    n1764_li,
    G30_p
  );


  buf

  (
    n1776_li,
    G31_p
  );


  buf

  (
    n1779_li,
    n1776_lo_p
  );


  buf

  (
    n1788_li,
    G32_p
  );


  buf

  (
    n1791_li,
    n1788_lo_p
  );


  buf

  (
    n1794_li,
    n1791_lo_p
  );


  buf

  (
    n1797_li,
    n1794_lo_p
  );


  buf

  (
    n1800_li,
    G33_p
  );


  buf

  (
    n1812_li,
    G34_p
  );


  buf

  (
    n1824_li,
    G35_p
  );


  buf

  (
    n1836_li,
    G36_p
  );


  buf

  (
    n1848_li,
    G37_p
  );


  buf

  (
    n1860_li,
    G38_p
  );


  buf

  (
    n1872_li,
    G39_p
  );


  buf

  (
    n1884_li,
    G40_p
  );


  buf

  (
    n1896_li,
    G41_p
  );


  buf

  (
    n1899_li,
    n1896_lo_p
  );


  buf

  (
    n1908_li,
    G42_p
  );


  buf

  (
    n1911_li,
    n1908_lo_p
  );


  buf

  (
    n1920_li,
    G43_p
  );


  buf

  (
    n1923_li,
    n1920_lo_p
  );


  buf

  (
    n1926_li,
    n1923_lo_p
  );


  buf

  (
    n1929_li,
    n1926_lo_p
  );


  buf

  (
    n1932_li,
    G44_p
  );


  buf

  (
    n1944_li,
    G45_p
  );


  buf

  (
    n1956_li,
    G46_p
  );


  buf

  (
    n1968_li,
    G47_p
  );


  buf

  (
    n1980_li,
    G48_p
  );


  buf

  (
    n1992_li,
    G49_p
  );


  buf

  (
    n2004_li,
    G50_p
  );


  buf

  (
    n2016_li,
    G51_p
  );


  buf

  (
    n2019_li,
    n2016_lo_p
  );


  buf

  (
    n2028_li,
    G52_p
  );


  buf

  (
    n2031_li,
    n2028_lo_p
  );


  buf

  (
    n2040_li,
    G53_p
  );


  buf

  (
    n2043_li,
    n2040_lo_p
  );


  buf

  (
    n2046_li,
    n2043_lo_p
  );


  buf

  (
    n2049_li,
    n2046_lo_p
  );


  buf

  (
    n2052_li,
    G54_p
  );


  buf

  (
    n2064_li,
    G55_p
  );


  buf

  (
    n2076_li,
    G56_p
  );


  buf

  (
    n2088_li,
    G57_p
  );


  buf

  (
    n2100_li,
    G58_p
  );


  buf

  (
    n2112_li,
    G59_p
  );


  buf

  (
    n2124_li,
    G60_p
  );


  buf

  (
    n2136_li,
    G61_p
  );


  buf

  (
    n2148_li,
    G62_p
  );


  buf

  (
    n2151_li,
    n2148_lo_p
  );


  buf

  (
    n2160_li,
    G63_p
  );


  buf

  (
    n2163_li,
    n2160_lo_p
  );


  buf

  (
    n2172_li,
    G64_p
  );


  buf

  (
    n2175_li,
    n2172_lo_p
  );


  buf

  (
    n2178_li,
    n2175_lo_p
  );


  buf

  (
    n2181_li,
    n2178_lo_p
  );


  buf

  (
    n2184_li,
    G65_p
  );


  buf

  (
    n2196_li,
    G66_p
  );


  buf

  (
    n2208_li,
    G67_p
  );


  buf

  (
    n2220_li,
    G68_p
  );


  buf

  (
    n2232_li,
    G69_p
  );


  buf

  (
    n2244_li,
    G70_p
  );


  buf

  (
    n2256_li,
    G71_p
  );


  buf

  (
    n2268_li,
    G72_p
  );


  buf

  (
    n2280_li,
    G73_p
  );


  buf

  (
    n2283_li,
    n2280_lo_p
  );


  buf

  (
    n2292_li,
    G74_p
  );


  buf

  (
    n2295_li,
    n2292_lo_p
  );


  buf

  (
    n2298_li,
    n2295_lo_p
  );


  buf

  (
    n2301_li,
    n2298_lo_p
  );


  buf

  (
    n2304_li,
    G75_p
  );


  buf

  (
    n2316_li,
    G76_p
  );


  buf

  (
    n2319_li,
    n2316_lo_p
  );


  buf

  (
    n2322_li,
    n2319_lo_p
  );


  buf

  (
    n2325_li,
    n2322_lo_p
  );


  buf

  (
    n2328_li,
    G77_p
  );


  buf

  (
    n2331_li,
    n2328_lo_p
  );


  buf

  (
    n2340_li,
    G78_p
  );


  buf

  (
    n2343_li,
    n2340_lo_p
  );


  buf

  (
    n2376_li,
    G81_p
  );


  buf

  (
    n2379_li,
    n2376_lo_p
  );


  buf

  (
    n2388_li,
    G82_p
  );


  buf

  (
    n2400_li,
    G83_p
  );


  buf

  (
    n2412_li,
    G84_p
  );


  buf

  (
    n2415_li,
    n2412_lo_p
  );


  buf

  (
    n2424_li,
    G85_p
  );


  buf

  (
    n2436_li,
    G86_p
  );


  buf

  (
    n2439_li,
    n2436_lo_p
  );


  buf

  (
    n2442_li,
    n2439_lo_p
  );


  buf

  (
    n2445_li,
    n2442_lo_p
  );


  buf

  (
    n2448_li,
    G87_p
  );


  buf

  (
    n2451_li,
    n2448_lo_p
  );


  buf

  (
    n2460_li,
    G88_p
  );


  buf

  (
    n2463_li,
    n2460_lo_p
  );


  buf

  (
    n2496_li,
    G91_p
  );


  buf

  (
    n2499_li,
    n2496_lo_p
  );


  buf

  (
    n2508_li,
    G92_p
  );


  buf

  (
    n2520_li,
    G93_p
  );


  buf

  (
    n2532_li,
    G94_p
  );


  buf

  (
    n2535_li,
    n2532_lo_p
  );


  buf

  (
    n2544_li,
    G95_p
  );


  buf

  (
    n2556_li,
    G96_p
  );


  buf

  (
    n2559_li,
    n2556_lo_p
  );


  buf

  (
    n2562_li,
    n2559_lo_p
  );


  buf

  (
    n2565_li,
    n2562_lo_p
  );


  buf

  (
    n2568_li,
    G97_p
  );


  buf

  (
    n2571_li,
    n2568_lo_p
  );


  buf

  (
    n2580_li,
    G98_p
  );


  buf

  (
    n2583_li,
    n2580_lo_p
  );


  buf

  (
    n2616_li,
    G101_p
  );


  buf

  (
    n2619_li,
    n2616_lo_p
  );


  buf

  (
    n2628_li,
    G102_p
  );


  buf

  (
    n2640_li,
    G103_p
  );


  buf

  (
    n2652_li,
    G104_p
  );


  buf

  (
    n2655_li,
    n2652_lo_p
  );


  buf

  (
    n2664_li,
    G105_p
  );


  buf

  (
    n2676_li,
    G106_p
  );


  buf

  (
    n2679_li,
    n2676_lo_p
  );


  buf

  (
    n2682_li,
    n2679_lo_p
  );


  buf

  (
    n2685_li,
    n2682_lo_p
  );


  buf

  (
    n2688_li,
    G107_p
  );


  buf

  (
    n2691_li,
    n2688_lo_p
  );


  buf

  (
    n2700_li,
    G108_p
  );


  buf

  (
    n2703_li,
    n2700_lo_p
  );


  buf

  (
    n2736_li,
    G111_p
  );


  buf

  (
    n2739_li,
    n2736_lo_p
  );


  buf

  (
    n2748_li,
    G112_p
  );


  buf

  (
    n2760_li,
    G113_p
  );


  buf

  (
    n2772_li,
    G114_p
  );


  buf

  (
    n2775_li,
    n2772_lo_p
  );


  buf

  (
    n2784_li,
    G115_p
  );


  buf

  (
    n2787_li,
    n2784_lo_p
  );


  buf

  (
    n2790_li,
    n2787_lo_p
  );


  buf

  (
    n2793_li,
    n2790_lo_p
  );


  buf

  (
    n2796_li,
    G116_p
  );


  buf

  (
    n2799_li,
    n2796_lo_p
  );


  buf

  (
    n2802_li,
    n2799_lo_p
  );


  buf

  (
    n2805_li,
    n2802_lo_p
  );


  buf

  (
    n2808_li,
    G117_p
  );


  buf

  (
    n2820_li,
    G118_p
  );


  buf

  (
    n2823_li,
    n2820_lo_p
  );


  buf

  (
    n2826_li,
    n2823_lo_p
  );


  buf

  (
    n2832_li,
    G119_p
  );


  buf

  (
    n2835_li,
    n2832_lo_p
  );


  buf

  (
    n2838_li,
    n2835_lo_p
  );


  buf

  (
    n2841_li,
    n2838_lo_p
  );


  buf

  (
    n2844_li,
    G120_p
  );


  buf

  (
    n2856_li,
    G121_p
  );


  buf

  (
    n2859_li,
    n2856_lo_p
  );


  buf

  (
    n2862_li,
    n2859_lo_p
  );


  buf

  (
    n2865_li,
    n2862_lo_p
  );


  buf

  (
    n2868_li,
    G122_p
  );


  buf

  (
    n2871_li,
    n2868_lo_p
  );


  buf

  (
    n2874_li,
    n2871_lo_p
  );


  buf

  (
    n2877_li,
    n2874_lo_p
  );


  buf

  (
    n2880_li,
    G123_p
  );


  buf

  (
    n2883_li,
    n2880_lo_p
  );


  buf

  (
    n2886_li,
    n2883_lo_p
  );


  buf

  (
    n2889_li,
    n2886_lo_p
  );


  buf

  (
    n2892_li,
    G124_p
  );


  buf

  (
    n2895_li,
    n2892_lo_p
  );


  buf

  (
    n2898_li,
    n2895_lo_p
  );


  buf

  (
    n2901_li,
    n2898_lo_p
  );


  buf

  (
    n2904_li,
    G125_p
  );


  buf

  (
    n2907_li,
    n2904_lo_p
  );


  buf

  (
    n2916_li,
    G126_p
  );


  buf

  (
    n2928_li,
    G127_p
  );


  buf

  (
    n2940_li,
    G128_p
  );


  buf

  (
    n2952_li,
    G129_p
  );


  buf

  (
    n2955_li,
    n2952_lo_p
  );


  buf

  (
    n2964_li,
    G130_p
  );


  buf

  (
    n2976_li,
    G131_p
  );


  buf

  (
    n2988_li,
    G132_p
  );


  buf

  (
    n2991_li,
    n2988_lo_p
  );


  buf

  (
    n3000_li,
    G133_p
  );


  buf

  (
    n3003_li,
    n3000_lo_p
  );


  buf

  (
    n3012_li,
    G134_p
  );


  buf

  (
    n3015_li,
    n3012_lo_p
  );


  buf

  (
    n3024_li,
    G135_p
  );


  buf

  (
    n3027_li,
    n3024_lo_p
  );


  buf

  (
    n3036_li,
    G136_p
  );


  buf

  (
    n3039_li,
    n3036_lo_p
  );


  buf

  (
    n3048_li,
    G137_p
  );


  buf

  (
    n3051_li,
    n3048_lo_p
  );


  buf

  (
    n3054_li,
    n3051_lo_p
  );


  buf

  (
    n3057_li,
    n3054_lo_p
  );


  buf

  (
    n3060_li,
    G138_p
  );


  buf

  (
    n3072_li,
    G139_p
  );


  buf

  (
    n3081_li,
    n3078_lo_buf_o2_p_spl_
  );


  buf

  (
    n3084_li,
    G140_p
  );


  buf

  (
    n3087_li,
    n3084_lo_p
  );


  buf

  (
    n3093_li,
    n3090_lo_buf_o2_p_spl_
  );


  buf

  (
    n3096_li,
    G141_p
  );


  buf

  (
    n3105_li,
    n3102_lo_buf_o2_p_spl_
  );


  buf

  (
    n3108_li,
    G142_p
  );


  buf

  (
    n3117_li,
    n3114_lo_buf_o2_p_spl_
  );


  buf

  (
    n3120_li,
    G143_p
  );


  buf

  (
    n3123_li,
    n3120_lo_p
  );


  buf

  (
    n3126_li,
    n3123_lo_p
  );


  buf

  (
    n3129_li,
    n3126_lo_p_spl_0
  );


  buf

  (
    n3132_li,
    G144_p
  );


  buf

  (
    n3135_li,
    n3132_lo_p
  );


  buf

  (
    n3138_li,
    n3135_lo_p
  );


  buf

  (
    n3141_li,
    n3138_lo_p_spl_0
  );


  buf

  (
    n3168_li,
    G147_p
  );


  buf

  (
    n3171_li,
    n3168_lo_p
  );


  buf

  (
    n3174_li,
    n3171_lo_p
  );


  buf

  (
    n3177_li,
    n3174_lo_p
  );


  buf

  (
    n3180_li,
    G148_p
  );


  buf

  (
    n3183_li,
    n3180_lo_p
  );


  buf

  (
    n3192_li,
    G149_p
  );


  buf

  (
    n3195_li,
    n3192_lo_p
  );


  buf

  (
    n3204_li,
    G150_p
  );


  buf

  (
    n3207_li,
    n3204_lo_p
  );


  buf

  (
    n3216_li,
    G151_p
  );


  buf

  (
    n3219_li,
    n3216_lo_p
  );


  buf

  (
    n3228_li,
    G152_p
  );


  buf

  (
    n3231_li,
    n3228_lo_p
  );


  buf

  (
    n3240_li,
    G153_p
  );


  buf

  (
    n3243_li,
    n3240_lo_p
  );


  buf

  (
    n3252_li,
    G154_p
  );


  buf

  (
    n3255_li,
    n3252_lo_p
  );


  buf

  (
    n3258_li,
    n3255_lo_p
  );


  buf

  (
    n3264_li,
    G155_p
  );


  buf

  (
    n3267_li,
    n3264_lo_p
  );


  buf

  (
    n3270_li,
    n3267_lo_p
  );


  buf

  (
    n3276_li,
    G156_p
  );


  buf

  (
    n3279_li,
    n3276_lo_p
  );


  buf

  (
    n3282_li,
    n3279_lo_p
  );


  buf

  (
    n3288_li,
    G157_p
  );


  buf

  (
    n3291_li,
    n3288_lo_p
  );


  buf

  (
    n3294_li,
    n3291_lo_p
  );


  buf

  (
    n4537_i2,
    n5222_o2_p_spl_1
  );


  buf

  (
    n4538_i2,
    n5223_o2_p_spl_
  );


  buf

  (
    n4710_i2,
    n5553_o2_p_spl_
  );


  buf

  (
    n4711_i2,
    n5554_o2_p_spl_
  );


  buf

  (
    n4803_i2,
    n1304_inv_p
  );


  buf

  (
    n4804_i2,
    n1307_inv_p
  );


  buf

  (
    n4843_i2,
    n1364_inv_p
  );


  buf

  (
    n4844_i2,
    n1367_inv_p
  );


  buf

  (
    n4927_i2,
    G1017_o2_p_spl_
  );


  buf

  (
    n4928_i2,
    G1008_o2_p_spl_1
  );


  buf

  (
    n4945_i2,
    n1400_inv_p
  );


  buf

  (
    n4946_i2,
    n1403_inv_p
  );


  buf

  (
    n5009_i2,
    n1418_inv_p
  );


  buf

  (
    n5178_i2,
    G1002_o2_p_spl_
  );


  buf

  (
    n5179_i2,
    G998_o2_p
  );


  buf

  (
    n5477_i2,
    G1053_o2_p_spl_
  );


  buf

  (
    n5478_i2,
    G1049_o2_p_spl_1
  );


  buf

  (
    n5479_i2,
    n2003_inv_p_spl_
  );


  buf

  (
    n5222_i2,
    G1044_o2_p
  );


  buf

  (
    n5223_i2,
    G1039_o2_p_spl_0
  );


  buf

  (
    n5553_i2,
    G1026_o2_p_spl_10
  );


  buf

  (
    n5554_i2,
    G1021_o2_p_spl_10
  );


  buf

  (
    G491_i2,
    n1686_lo_p_spl_11
  );


  buf

  (
    n2922_lo_buf_i2,
    n2919_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2946_lo_buf_i2,
    n2943_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2970_lo_buf_i2,
    n2967_lo_buf_o2_p_spl_1
  );


  buf

  (
    n2982_lo_buf_i2,
    n2979_lo_buf_o2_p_spl_1
  );


  buf

  (
    n3066_lo_buf_i2,
    n3063_lo_buf_o2_p_spl_1
  );


  buf

  (
    n3078_lo_buf_i2,
    n3075_lo_buf_o2_p_spl_1
  );


  buf

  (
    n3102_lo_buf_i2,
    n3099_lo_buf_o2_p_spl_1
  );


  buf

  (
    n3114_lo_buf_i2,
    n3111_lo_buf_o2_p_spl_1
  );


  buf

  (
    G1321_i2,
    g1014_n_spl_1
  );


  buf

  (
    G1033_i2,
    g1017_n_spl_0
  );


  buf

  (
    G1030_i2,
    g1020_n_spl_0
  );


  buf

  (
    G1072_i2,
    g1023_n_spl_0
  );


  buf

  (
    G1159_i2,
    G1026_o2_p_spl_10
  );


  buf

  (
    G1152_i2,
    G1021_o2_p_spl_10
  );


  buf

  (
    n2958_lo_buf_i2,
    n2955_lo_p_spl_
  );


  buf

  (
    n2994_lo_buf_i2,
    n2991_lo_p_spl_1
  );


  buf

  (
    n3006_lo_buf_i2,
    n3003_lo_p_spl_1
  );


  buf

  (
    n3030_lo_buf_i2,
    n3027_lo_p_spl_
  );


  buf

  (
    n3042_lo_buf_i2,
    n3039_lo_p_spl_1
  );


  buf

  (
    n3090_lo_buf_i2,
    n3087_lo_p_spl_
  );


  buf

  (
    G370_i2,
    n2919_lo_buf_o2_p_spl_1
  );


  buf

  (
    G447_i2,
    n2943_lo_buf_o2_p_spl_1
  );


  buf

  (
    G455_i2,
    n2967_lo_buf_o2_p_spl_1
  );


  buf

  (
    G459_i2,
    n2979_lo_buf_o2_p_spl_1
  );


  buf

  (
    G497_i2,
    n3063_lo_buf_o2_p_spl_1
  );


  buf

  (
    G503_i2,
    n3075_lo_buf_o2_p_spl_1
  );


  buf

  (
    G511_i2,
    n3099_lo_buf_o2_p_spl_1
  );


  buf

  (
    G515_i2,
    n3111_lo_buf_o2_p_spl_1
  );


  buf

  (
    G1036_i2,
    g1034_n_spl_0
  );


  buf

  (
    G1062_i2,
    g1045_n_spl_0
  );


  buf

  (
    G1067_i2,
    g1056_n_spl_0
  );


  buf

  (
    G1014_i2,
    g1067_n_spl_01
  );


  buf

  (
    G1171_i2,
    g1017_n_spl_1
  );


  buf

  (
    G1166_i2,
    g1020_n_spl_1
  );


  buf

  (
    n3018_lo_buf_i2,
    n3015_lo_p_spl_
  );


  buf

  (
    G766_i2,
    n1686_lo_p_spl_11
  );


  buf

  (
    G451_i2,
    n2955_lo_p_spl_
  );


  buf

  (
    G463_i2,
    n2991_lo_p_spl_1
  );


  buf

  (
    G467_i2,
    n3003_lo_p_spl_1
  );


  buf

  (
    G475_i2,
    n3027_lo_p_spl_
  );


  buf

  (
    G479_i2,
    n3039_lo_p_spl_1
  );


  buf

  (
    G507_i2,
    n3087_lo_p_spl_
  );


  buf

  (
    G1017_i2,
    g1078_n_spl_00
  );


  buf

  (
    G1008_i2,
    g1089_n_spl_10
  );


  buf

  (
    G1176_i2,
    g1034_n_spl_1
  );


  buf

  (
    G1144_i2,
    g1067_n_spl_01
  );


  buf

  (
    n2910_lo_buf_i2,
    n2907_lo_p_spl_1
  );


  buf

  (
    G471_i2,
    n3015_lo_p_spl_
  );


  buf

  (
    G2138_i2,
    g1092_p_spl_
  );


  buf

  (
    G2147_i2,
    g1095_p_spl_
  );


  buf

  (
    G1148_i2,
    g1078_n_spl_00
  );


  buf

  (
    G1137_i2,
    g1089_n_spl_10
  );


  buf

  (
    G1329_i2,
    g1067_n_spl_1
  );


  buf

  (
    G374_i2,
    n3150_lo_buf_o2_p_spl_10
  );


  buf

  (
    G386_i2,
    n3162_lo_buf_o2_p_spl_10
  );


  buf

  (
    G663_i2,
    n3150_lo_buf_o2_p_spl_10
  );


  buf

  (
    G674_i2,
    n3162_lo_buf_o2_p_spl_10
  );


  buf

  (
    G578_i2,
    n3126_lo_p_spl_0
  );


  buf

  (
    G575_i2,
    n3138_lo_p_spl_0
  );


  not

  (
    G2505_i2,
    g1157_n_spl_
  );


  not

  (
    G2508_i2,
    g1219_n_spl_
  );


  buf

  (
    G987_i2,
    g1222_n_spl_
  );


  buf

  (
    G984_i2,
    g1225_n_spl_
  );


  buf

  (
    G1862_i2,
    g1228_n_spl_0
  );


  buf

  (
    G1859_i2,
    g1231_n_spl_0
  );


  buf

  (
    G1260_i2,
    g1240_n_spl_
  );


  buf

  (
    G1865_i2,
    g1249_p_spl_
  );


  buf

  (
    G2073_i2,
    g1252_n_spl_
  );


  buf

  (
    G1402_i2,
    g1272_p_spl_
  );


  buf

  (
    G2048_i2,
    g1292_n_spl_
  );


  buf

  (
    G2276_i2,
    g1312_p_spl_
  );


  buf

  (
    G366_i2,
    n2907_lo_p_spl_1
  );


  not

  (
    G2141_i2,
    g1315_n_spl_
  );


  not

  (
    G2008_i2,
    g1317_n_spl_
  );


  not

  (
    G2011_i2,
    g1319_n_spl_
  );


  not

  (
    G2150_i2,
    g1322_n_spl_
  );


  not

  (
    G2026_i2,
    g1324_n_spl_
  );


  not

  (
    G2029_i2,
    g1326_n_spl_
  );


  not

  (
    G2023_i2,
    g1330_n_spl_
  );


  not

  (
    G2041_i2,
    g1332_n_spl_
  );


  buf

  (
    G2017_i2,
    g1334_p_spl_
  );


  buf

  (
    G2020_i2,
    g1336_p_spl_
  );


  buf

  (
    G2035_i2,
    g1338_p_spl_
  );


  buf

  (
    G2038_i2,
    g1340_p_spl_
  );


  not

  (
    G2228_i2,
    g1344_n_spl_
  );


  not

  (
    G2231_i2,
    g1348_n_spl_
  );


  not

  (
    G2234_i2,
    g1352_n_spl_
  );


  not

  (
    G2237_i2,
    g1356_n_spl_
  );


  not

  (
    G1904_i2,
    g1358_n_spl_
  );


  not

  (
    G1907_i2,
    g1360_n_spl_
  );


  not

  (
    G1928_i2,
    g1362_n_spl_
  );


  not

  (
    G1931_i2,
    g1364_n_spl_
  );


  buf

  (
    G1893_i2,
    g1366_p_spl_1
  );


  buf

  (
    G1896_i2,
    g1368_p_spl_1
  );


  not

  (
    G1899_i2,
    g1370_n_spl_1
  );


  buf

  (
    G1937_i2,
    g1366_p_spl_1
  );


  buf

  (
    G1940_i2,
    g1368_p_spl_1
  );


  not

  (
    G1943_i2,
    g1370_n_spl_1
  );


  buf

  (
    G1336_i2,
    g1078_n_spl_0
  );


  not

  (
    G1996_i2,
    g1374_n_spl_
  );


  not

  (
    G1999_i2,
    g1378_n_spl_
  );


  not

  (
    G2002_i2,
    g1382_n_spl_
  );


  not

  (
    G2005_i2,
    g1386_n_spl_
  );


  buf

  (
    G2014_i2,
    g1388_p_spl_0
  );


  buf

  (
    G2032_i2,
    g1390_p_spl_0
  );


  buf

  (
    G1076_i2,
    g1401_n_spl_0
  );


  buf

  (
    G1002_i2,
    g1412_n_spl_0
  );


  buf

  (
    G998_i2,
    g1423_n_spl_0
  );


  not

  (
    G1890_i2,
    g1425_n_spl_00
  );


  not

  (
    G1934_i2,
    g1425_n_spl_00
  );


  buf

  (
    G1044_i2,
    g1436_n_spl_0
  );


  not

  (
    G1039_i2,
    g1447_p_spl_
  );


  buf

  (
    n1770_lo_buf_i2,
    n1764_lo_p
  );


  buf

  (
    G342_i2,
    n2808_lo_p_spl_10
  );


  buf

  (
    G354_i2,
    n2844_lo_p_spl_10
  );


  buf

  (
    G1193_i2,
    g1436_n_spl_
  );


  buf

  (
    n3234_lo_buf_i2,
    n3231_lo_p_spl_
  );


  buf

  (
    n3246_lo_buf_i2,
    n3243_lo_p_spl_
  );


  buf

  (
    G783_i2,
    n1328_inv_p
  );


  buf

  (
    G786_i2,
    n1331_inv_p
  );


  buf

  (
    G792_i2,
    n1334_inv_p
  );


  buf

  (
    G795_i2,
    n1337_inv_p
  );


  buf

  (
    G815_i2,
    n1340_inv_p
  );


  buf

  (
    G818_i2,
    n1343_inv_p
  );


  buf

  (
    G824_i2,
    n1346_inv_p
  );


  buf

  (
    G827_i2,
    n1349_inv_p
  );


  buf

  (
    G789_i2,
    n1376_inv_p
  );


  buf

  (
    G798_i2,
    n1379_inv_p
  );


  buf

  (
    G801_i2,
    n1382_inv_p
  );


  buf

  (
    G807_i2,
    n1385_inv_p
  );


  buf

  (
    G812_i2,
    n1388_inv_p
  );


  buf

  (
    G821_i2,
    n1391_inv_p
  );


  buf

  (
    G804_i2,
    n1409_inv_p
  );


  buf

  (
    G780_i2,
    n1481_inv_p
  );


  buf

  (
    G1231_i2,
    G1039_o2_p_spl_0
  );


  buf

  (
    G1572_i2,
    g1014_n_spl_1
  );


  buf

  (
    G1377_i2,
    G1021_o2_p_spl_11
  );


  not

  (
    G1253_i2,
    g1458_n
  );


  buf

  (
    G1359_i2,
    g1460_p
  );


  not

  (
    G1258_i2,
    g1471_n
  );


  buf

  (
    G1367_i2,
    g1473_p
  );


  buf

  (
    G1358_i2,
    g1475_p
  );


  buf

  (
    G1366_i2,
    g1477_p
  );


  not

  (
    G2057_i2,
    g1485_n
  );


  buf

  (
    G2117_i2,
    g1487_p
  );


  not

  (
    G2118_i2,
    g1489_p
  );


  not

  (
    G1254_i2,
    g1491_n
  );


  not

  (
    G1259_i2,
    g1493_n
  );


  not

  (
    G2058_i2,
    g1495_n
  );


  buf

  (
    G405_i2,
    n3150_lo_buf_o2_p_spl_11
  );


  buf

  (
    G417_i2,
    n3162_lo_buf_o2_p_spl_11
  );


  buf

  (
    G1269_i2,
    g1498_n
  );


  buf

  (
    G1275_i2,
    g1501_n
  );


  buf

  (
    G1287_i2,
    g1504_n
  );


  buf

  (
    G1266_i2,
    g1507_n
  );


  buf

  (
    G1272_i2,
    g1510_n
  );


  buf

  (
    G1278_i2,
    g1513_n
  );


  buf

  (
    G1281_i2,
    g1516_n
  );


  buf

  (
    G1284_i2,
    g1519_n
  );


  buf

  (
    G1290_i2,
    g1522_n
  );


  buf

  (
    G1293_i2,
    g1525_n
  );


  buf

  (
    G1299_i2,
    g1528_n
  );


  buf

  (
    G1305_i2,
    g1531_n
  );


  buf

  (
    G1296_i2,
    g1534_n
  );


  buf

  (
    G1302_i2,
    g1537_n
  );


  buf

  (
    G1308_i2,
    g1540_n
  );


  buf

  (
    G1311_i2,
    g1543_n
  );


  buf

  (
    G811_i2,
    n3126_lo_p_spl_
  );


  buf

  (
    G810_i2,
    n3138_lo_p_spl_
  );


  buf

  (
    G1728_i2,
    g1546_p
  );


  not

  (
    G2512_i2,
    g1547_p
  );


  buf

  (
    G1114_i2,
    g1222_n_spl_
  );


  buf

  (
    G1113_i2,
    g1225_n_spl_
  );


  buf

  (
    G1992_i2,
    g1228_n_spl_
  );


  buf

  (
    G1991_i2,
    g1231_n_spl_
  );


  buf

  (
    G1426_i2,
    g1240_n_spl_
  );


  buf

  (
    G1966_i2,
    g1249_p_spl_
  );


  buf

  (
    G2211_i2,
    g1252_n_spl_
  );


  buf

  (
    G1509_i2,
    g1272_p_spl_
  );


  buf

  (
    G2153_i2,
    g1292_n_spl_
  );


  buf

  (
    G2329_i2,
    g1312_p_spl_
  );


  buf

  (
    G1540_i2,
    g1078_n_spl_1
  );


  buf

  (
    G2167_i2,
    g1388_p_spl_0
  );


  buf

  (
    G2191_i2,
    g1390_p_spl_0
  );


  buf

  (
    G1234_i2,
    g1401_n_spl_0
  );


  buf

  (
    G1132_i2,
    g1412_n_spl_1
  );


  buf

  (
    G1129_i2,
    g1423_n_spl_0
  );


  not

  (
    G2088_i2,
    g1425_n_spl_01
  );


  not

  (
    G2106_i2,
    g1425_n_spl_01
  );


  not

  (
    G1314_i2,
    g1550_n_spl_00
  );


  buf

  (
    G636_i2,
    n2808_lo_p_spl_10
  );


  buf

  (
    G647_i2,
    n2844_lo_p_spl_10
  );


  buf

  (
    n3186_lo_buf_i2,
    n3183_lo_p
  );


  buf

  (
    n3198_lo_buf_i2,
    n3195_lo_p
  );


  buf

  (
    n3210_lo_buf_i2,
    n3207_lo_p
  );


  buf

  (
    n3222_lo_buf_i2,
    n3219_lo_p
  );


  buf

  (
    G1225_i2,
    g1023_n_spl_
  );


  buf

  (
    G1342_i2,
    G1026_o2_p_spl_1
  );


  buf

  (
    G1222_i2,
    g1045_n_spl_
  );


  buf

  (
    G1228_i2,
    g1056_n_spl_
  );


  buf

  (
    G1348_i2,
    g1017_n_spl_1
  );


  buf

  (
    G1345_i2,
    g1020_n_spl_1
  );


  buf

  (
    G1351_i2,
    g1034_n_spl_1
  );


  buf

  (
    G2242_i2,
    g1554_n
  );


  buf

  (
    G2260_i2,
    g1558_n
  );


  buf

  (
    G1374_i2,
    g1089_n_spl_1
  );


  buf

  (
    G1537_i2,
    g1067_n_spl_1
  );


  buf

  (
    G301_i2,
    n2808_lo_p_spl_11
  );


  buf

  (
    G313_i2,
    n2844_lo_p_spl_11
  );


  not

  (
    G2365_i2,
    g1559_n
  );


  not

  (
    G2255_i2,
    g1560_p
  );


  not

  (
    G2253_i2,
    g1561_p
  );


  not

  (
    G2395_i2,
    g1562_n
  );


  not

  (
    G2272_i2,
    g1563_p
  );


  not

  (
    G2270_i2,
    g1564_p
  );


  not

  (
    G2245_i2,
    g1565_p
  );


  not

  (
    G2262_i2,
    g1566_p
  );


  buf

  (
    G2249_i2,
    g1567_n
  );


  buf

  (
    G2247_i2,
    g1568_n
  );


  buf

  (
    G2266_i2,
    g1569_n
  );


  buf

  (
    G2264_i2,
    g1570_n
  );


  not

  (
    G2403_i2,
    g1571_p
  );


  not

  (
    G2401_i2,
    g1572_p
  );


  not

  (
    G2410_i2,
    g1573_p
  );


  not

  (
    G2408_i2,
    g1574_p
  );


  not

  (
    G2306_i2,
    g1575_n
  );


  not

  (
    G2305_i2,
    g1576_n
  );


  not

  (
    G2314_i2,
    g1577_n
  );


  not

  (
    G2313_i2,
    g1578_n
  );


  buf

  (
    G2303_i2,
    g1579_p
  );


  buf

  (
    G2302_i2,
    g1580_p
  );


  not

  (
    G2301_i2,
    g1581_n
  );


  buf

  (
    G2311_i2,
    g1582_p
  );


  buf

  (
    G2310_i2,
    g1583_p
  );


  not

  (
    G2309_i2,
    g1584_n
  );


  not

  (
    G2404_i2,
    g1585_p
  );


  not

  (
    G2411_i2,
    g1586_p
  );


  not

  (
    G2420_i2,
    g1587_n
  );


  not

  (
    G2419_i2,
    g1588_n
  );


  not

  (
    G2433_i2,
    g1589_n
  );


  not

  (
    G2432_i2,
    g1590_n
  );


  buf

  (
    G402_i2,
    n3231_lo_p_spl_
  );


  buf

  (
    G403_i2,
    n3243_lo_p_spl_
  );


  buf

  (
    G1053_i2,
    g1601_n
  );


  buf

  (
    G1049_i2,
    g1612_n
  );


  buf

  (
    G1058_i2,
    g1619_p
  );


  buf

  (
    G1364_i2,
    G1039_o2_p_spl_
  );


  buf

  (
    G1079_i2,
    g1630_n
  );


  buf

  (
    G1478_i2,
    G1021_o2_p_spl_11
  );


  buf

  (
    G707_i2,
    n3150_lo_buf_o2_p_spl_11
  );


  buf

  (
    G718_i2,
    n3162_lo_buf_o2_p_spl_11
  );


  buf

  (
    G2417_i2,
    g1633_n
  );


  buf

  (
    G2414_i2,
    g1636_p
  );


  buf

  (
    G2431_i2,
    g1639_n
  );


  buf

  (
    G2428_i2,
    g1642_p
  );


  buf

  (
    G1653_i2,
    g1078_n_spl_1
  );


  buf

  (
    G2213_i2,
    g1646_n
  );


  buf

  (
    G2221_i2,
    g1650_n
  );


  buf

  (
    G2250_i2,
    g1388_p_spl_
  );


  buf

  (
    G2267_i2,
    g1390_p_spl_
  );


  buf

  (
    G1365_i2,
    g1401_n_spl_
  );


  buf

  (
    G1368_i2,
    g1412_n_spl_1
  );


  buf

  (
    G1371_i2,
    g1423_n_spl_
  );


  not

  (
    G2218_i2,
    g1425_n_spl_1
  );


  not

  (
    G2225_i2,
    g1425_n_spl_1
  );


  buf

  (
    n1503_lo_buf_i2,
    n1500_lo_p
  );


  buf

  (
    n1863_lo_buf_i2,
    n1860_lo_p
  );


  buf

  (
    n1887_lo_buf_i2,
    n1884_lo_p
  );


  buf

  (
    n1983_lo_buf_i2,
    n1980_lo_p
  );


  buf

  (
    n2007_lo_buf_i2,
    n2004_lo_p
  );


  buf

  (
    n2115_lo_buf_i2,
    n2112_lo_p
  );


  buf

  (
    n2139_lo_buf_i2,
    n2136_lo_p
  );


  buf

  (
    n2247_lo_buf_i2,
    n2244_lo_p
  );


  buf

  (
    n2271_lo_buf_i2,
    n2268_lo_p
  );


  buf

  (
    n2919_lo_buf_i2,
    n2916_lo_p
  );


  buf

  (
    n2943_lo_buf_i2,
    n2940_lo_p
  );


  buf

  (
    n2967_lo_buf_i2,
    n2964_lo_p
  );


  buf

  (
    n2979_lo_buf_i2,
    n2976_lo_p
  );


  buf

  (
    n3063_lo_buf_i2,
    n3060_lo_p
  );


  buf

  (
    n3075_lo_buf_i2,
    n3072_lo_p
  );


  buf

  (
    n3099_lo_buf_i2,
    n3096_lo_p
  );


  buf

  (
    n3111_lo_buf_i2,
    n3108_lo_p
  );


  buf

  (
    G878_i2,
    g1652_p
  );


  buf

  (
    G875_i2,
    g1654_p
  );


  buf

  (
    G661_i2,
    g1656_p
  );


  buf

  (
    G660_i2,
    g1658_p
  );


  buf

  (
    G879_i2,
    g1660_p
  );


  buf

  (
    G876_i2,
    g1661_p
  );


  not

  (
    G1320_i2,
    g1548_n_spl_
  );


  buf

  (
    G941_i2,
    g1663_p
  );


  buf

  (
    G732_i2,
    g1665_p
  );


  buf

  (
    G942_i2,
    g1667_p
  );


  not

  (
    G1493_i2,
    g1550_n_spl_00
  );


  not

  (
    G1498_i2,
    g1550_n_spl_0
  );


  buf

  (
    G877_i2,
    g1669_p
  );


  buf

  (
    G874_i2,
    g1671_p
  );


  buf

  (
    n1806_lo_buf_i2,
    n1800_lo_p
  );


  buf

  (
    n1878_lo_buf_i2,
    n1872_lo_p
  );


  buf

  (
    n1938_lo_buf_i2,
    n1932_lo_p
  );


  buf

  (
    n1998_lo_buf_i2,
    n1992_lo_p
  );


  buf

  (
    n2058_lo_buf_i2,
    n2052_lo_p
  );


  buf

  (
    n2130_lo_buf_i2,
    n2124_lo_p
  );


  buf

  (
    n2190_lo_buf_i2,
    n2184_lo_p
  );


  buf

  (
    n2262_lo_buf_i2,
    n2256_lo_p
  );


  buf

  (
    n2310_lo_buf_i2,
    n2304_lo_p
  );


  buf

  (
    n2406_lo_buf_i2,
    n2400_lo_p
  );


  buf

  (
    n2430_lo_buf_i2,
    n2424_lo_p
  );


  buf

  (
    n2526_lo_buf_i2,
    n2520_lo_p
  );


  buf

  (
    n2550_lo_buf_i2,
    n2544_lo_p
  );


  buf

  (
    n2646_lo_buf_i2,
    n2640_lo_p
  );


  buf

  (
    n2670_lo_buf_i2,
    n2664_lo_p
  );


  buf

  (
    n2766_lo_buf_i2,
    n2760_lo_p
  );


  buf

  (
    G603_i2,
    n2808_lo_p_spl_11
  );


  buf

  (
    G614_i2,
    n2844_lo_p_spl_11
  );


  buf

  (
    G1026_i2,
    g1682_n
  );


  buf

  (
    G1021_i2,
    g1693_n
  );


  buf

  (
    G940_i2,
    g1695_p
  );


  not

  (
    G1636_i2,
    g1550_n_spl_1
  );


  not

  (
    G1684_i2,
    g1550_n_spl_1
  );


  buf

  (
    n2352_lo_buf_i2,
    G79_p
  );


  buf

  (
    n2364_lo_buf_i2,
    G80_p
  );


  buf

  (
    n2472_lo_buf_i2,
    G89_p
  );


  buf

  (
    n2484_lo_buf_i2,
    G90_p
  );


  buf

  (
    n2592_lo_buf_i2,
    G99_p
  );


  buf

  (
    n2604_lo_buf_i2,
    G100_p
  );


  buf

  (
    n2712_lo_buf_i2,
    G109_p
  );


  buf

  (
    n2724_lo_buf_i2,
    G110_p
  );


  buf

  (
    n3150_lo_buf_i2,
    G145_p
  );


  buf

  (
    n3162_lo_buf_i2,
    G146_p
  );


  buf

  (
    n2865_lo_n_spl_,
    n2865_lo_n
  );


  buf

  (
    n2793_lo_n_spl_,
    n2793_lo_n
  );


  buf

  (
    n2793_lo_n_spl_0,
    n2793_lo_n_spl_
  );


  buf

  (
    n2793_lo_n_spl_1,
    n2793_lo_n_spl_
  );


  buf

  (
    g841_n_spl_,
    g841_n
  );


  buf

  (
    g841_n_spl_0,
    g841_n_spl_
  );


  buf

  (
    n2565_lo_n_spl_,
    n2565_lo_n
  );


  buf

  (
    n1929_lo_n_spl_,
    n1929_lo_n
  );


  buf

  (
    n2445_lo_n_spl_,
    n2445_lo_n
  );


  buf

  (
    n2049_lo_n_spl_,
    n2049_lo_n
  );


  buf

  (
    n2685_lo_n_spl_,
    n2685_lo_n
  );


  buf

  (
    n2181_lo_n_spl_,
    n2181_lo_n
  );


  buf

  (
    n2325_lo_n_spl_,
    n2325_lo_n
  );


  buf

  (
    n1797_lo_n_spl_,
    n1797_lo_n
  );


  buf

  (
    g849_n_spl_,
    g849_n
  );


  buf

  (
    g846_n_spl_,
    g846_n
  );


  buf

  (
    n2877_lo_p_spl_,
    n2877_lo_p
  );


  buf

  (
    n2877_lo_p_spl_0,
    n2877_lo_p_spl_
  );


  buf

  (
    n2877_lo_n_spl_,
    n2877_lo_n
  );


  buf

  (
    n2877_lo_n_spl_0,
    n2877_lo_n_spl_
  );


  buf

  (
    g856_n_spl_,
    g856_n
  );


  buf

  (
    g853_n_spl_,
    g853_n
  );


  buf

  (
    g853_n_spl_0,
    g853_n_spl_
  );


  buf

  (
    g853_n_spl_1,
    g853_n_spl_
  );


  buf

  (
    n2889_lo_p_spl_,
    n2889_lo_p
  );


  buf

  (
    n2889_lo_p_spl_0,
    n2889_lo_p_spl_
  );


  buf

  (
    n2889_lo_p_spl_00,
    n2889_lo_p_spl_0
  );


  buf

  (
    n2889_lo_p_spl_1,
    n2889_lo_p_spl_
  );


  buf

  (
    n1235_inv_p_spl_,
    n1235_inv_p
  );


  buf

  (
    n2889_lo_n_spl_,
    n2889_lo_n
  );


  buf

  (
    n2889_lo_n_spl_0,
    n2889_lo_n_spl_
  );


  buf

  (
    n2889_lo_n_spl_00,
    n2889_lo_n_spl_0
  );


  buf

  (
    n2889_lo_n_spl_1,
    n2889_lo_n_spl_
  );


  buf

  (
    n1232_inv_p_spl_,
    n1232_inv_p
  );


  buf

  (
    n4711_o2_n_spl_,
    n4711_o2_n
  );


  buf

  (
    g874_n_spl_,
    g874_n
  );


  buf

  (
    n5477_o2_n_spl_,
    n5477_o2_n
  );


  buf

  (
    g878_n_spl_,
    g878_n
  );


  buf

  (
    n1521_lo_n_spl_,
    n1521_lo_n
  );


  buf

  (
    G1728_o2_n_spl_,
    G1728_o2_n
  );


  buf

  (
    G1572_o2_p_spl_,
    G1572_o2_p
  );


  buf

  (
    G1728_o2_p_spl_,
    G1728_o2_p
  );


  buf

  (
    G1572_o2_n_spl_,
    G1572_o2_n
  );


  buf

  (
    n5179_o2_p_spl_,
    n5179_o2_p
  );


  buf

  (
    n5179_o2_p_spl_0,
    n5179_o2_p_spl_
  );


  buf

  (
    n1761_lo_n_spl_,
    n1761_lo_n
  );


  buf

  (
    G2512_o2_p_spl_,
    G2512_o2_p
  );


  buf

  (
    g1004_p_spl_,
    g1004_p
  );


  buf

  (
    g988_p_spl_,
    g988_p
  );


  buf

  (
    g895_p_spl_,
    g895_p
  );


  buf

  (
    g904_p_spl_,
    g904_p
  );


  buf

  (
    g886_p_spl_,
    g886_p
  );


  buf

  (
    g1007_n_spl_,
    g1007_n
  );


  buf

  (
    G1008_o2_n_spl_,
    G1008_o2_n
  );


  buf

  (
    G1008_o2_p_spl_,
    G1008_o2_p
  );


  buf

  (
    G1008_o2_p_spl_0,
    G1008_o2_p_spl_
  );


  buf

  (
    G1008_o2_p_spl_1,
    G1008_o2_p_spl_
  );


  buf

  (
    G636_o2_p_spl_,
    G636_o2_p
  );


  buf

  (
    G647_o2_p_spl_,
    G647_o2_p
  );


  buf

  (
    G342_o2_n_spl_,
    G342_o2_n
  );


  buf

  (
    G354_o2_n_spl_,
    G354_o2_n
  );


  buf

  (
    G707_o2_p_spl_,
    G707_o2_p
  );


  buf

  (
    G707_o2_p_spl_0,
    G707_o2_p_spl_
  );


  buf

  (
    G707_o2_p_spl_00,
    G707_o2_p_spl_0
  );


  buf

  (
    G707_o2_p_spl_01,
    G707_o2_p_spl_0
  );


  buf

  (
    G707_o2_p_spl_1,
    G707_o2_p_spl_
  );


  buf

  (
    G707_o2_p_spl_10,
    G707_o2_p_spl_1
  );


  buf

  (
    G707_o2_p_spl_11,
    G707_o2_p_spl_1
  );


  buf

  (
    G718_o2_p_spl_,
    G718_o2_p
  );


  buf

  (
    G718_o2_p_spl_0,
    G718_o2_p_spl_
  );


  buf

  (
    G718_o2_p_spl_00,
    G718_o2_p_spl_0
  );


  buf

  (
    G718_o2_p_spl_01,
    G718_o2_p_spl_0
  );


  buf

  (
    G718_o2_p_spl_1,
    G718_o2_p_spl_
  );


  buf

  (
    G718_o2_p_spl_10,
    G718_o2_p_spl_1
  );


  buf

  (
    G718_o2_p_spl_11,
    G718_o2_p_spl_1
  );


  buf

  (
    G405_o2_n_spl_,
    G405_o2_n
  );


  buf

  (
    G405_o2_n_spl_0,
    G405_o2_n_spl_
  );


  buf

  (
    G405_o2_n_spl_00,
    G405_o2_n_spl_0
  );


  buf

  (
    G405_o2_n_spl_01,
    G405_o2_n_spl_0
  );


  buf

  (
    G405_o2_n_spl_1,
    G405_o2_n_spl_
  );


  buf

  (
    G405_o2_n_spl_10,
    G405_o2_n_spl_1
  );


  buf

  (
    G405_o2_n_spl_11,
    G405_o2_n_spl_1
  );


  buf

  (
    G417_o2_n_spl_,
    G417_o2_n
  );


  buf

  (
    G417_o2_n_spl_0,
    G417_o2_n_spl_
  );


  buf

  (
    G417_o2_n_spl_00,
    G417_o2_n_spl_0
  );


  buf

  (
    G417_o2_n_spl_01,
    G417_o2_n_spl_0
  );


  buf

  (
    G417_o2_n_spl_1,
    G417_o2_n_spl_
  );


  buf

  (
    G417_o2_n_spl_10,
    G417_o2_n_spl_1
  );


  buf

  (
    G417_o2_n_spl_11,
    G417_o2_n_spl_1
  );


  buf

  (
    G603_o2_p_spl_,
    G603_o2_p
  );


  buf

  (
    G603_o2_p_spl_0,
    G603_o2_p_spl_
  );


  buf

  (
    G603_o2_p_spl_00,
    G603_o2_p_spl_0
  );


  buf

  (
    G603_o2_p_spl_000,
    G603_o2_p_spl_00
  );


  buf

  (
    G603_o2_p_spl_001,
    G603_o2_p_spl_00
  );


  buf

  (
    G603_o2_p_spl_01,
    G603_o2_p_spl_0
  );


  buf

  (
    G603_o2_p_spl_1,
    G603_o2_p_spl_
  );


  buf

  (
    G603_o2_p_spl_10,
    G603_o2_p_spl_1
  );


  buf

  (
    G603_o2_p_spl_11,
    G603_o2_p_spl_1
  );


  buf

  (
    G603_o2_n_spl_,
    G603_o2_n
  );


  buf

  (
    G603_o2_n_spl_0,
    G603_o2_n_spl_
  );


  buf

  (
    G603_o2_n_spl_00,
    G603_o2_n_spl_0
  );


  buf

  (
    G603_o2_n_spl_01,
    G603_o2_n_spl_0
  );


  buf

  (
    G603_o2_n_spl_1,
    G603_o2_n_spl_
  );


  buf

  (
    G614_o2_p_spl_,
    G614_o2_p
  );


  buf

  (
    G614_o2_p_spl_0,
    G614_o2_p_spl_
  );


  buf

  (
    G614_o2_p_spl_00,
    G614_o2_p_spl_0
  );


  buf

  (
    G614_o2_p_spl_000,
    G614_o2_p_spl_00
  );


  buf

  (
    G614_o2_p_spl_001,
    G614_o2_p_spl_00
  );


  buf

  (
    G614_o2_p_spl_01,
    G614_o2_p_spl_0
  );


  buf

  (
    G614_o2_p_spl_1,
    G614_o2_p_spl_
  );


  buf

  (
    G614_o2_p_spl_10,
    G614_o2_p_spl_1
  );


  buf

  (
    G614_o2_p_spl_11,
    G614_o2_p_spl_1
  );


  buf

  (
    G614_o2_n_spl_,
    G614_o2_n
  );


  buf

  (
    G614_o2_n_spl_0,
    G614_o2_n_spl_
  );


  buf

  (
    G614_o2_n_spl_00,
    G614_o2_n_spl_0
  );


  buf

  (
    G614_o2_n_spl_01,
    G614_o2_n_spl_0
  );


  buf

  (
    G614_o2_n_spl_1,
    G614_o2_n_spl_
  );


  buf

  (
    G301_o2_n_spl_,
    G301_o2_n
  );


  buf

  (
    G301_o2_n_spl_0,
    G301_o2_n_spl_
  );


  buf

  (
    G301_o2_n_spl_00,
    G301_o2_n_spl_0
  );


  buf

  (
    G301_o2_n_spl_000,
    G301_o2_n_spl_00
  );


  buf

  (
    G301_o2_n_spl_001,
    G301_o2_n_spl_00
  );


  buf

  (
    G301_o2_n_spl_01,
    G301_o2_n_spl_0
  );


  buf

  (
    G301_o2_n_spl_1,
    G301_o2_n_spl_
  );


  buf

  (
    G301_o2_n_spl_10,
    G301_o2_n_spl_1
  );


  buf

  (
    G301_o2_n_spl_11,
    G301_o2_n_spl_1
  );


  buf

  (
    G301_o2_p_spl_,
    G301_o2_p
  );


  buf

  (
    G301_o2_p_spl_0,
    G301_o2_p_spl_
  );


  buf

  (
    G301_o2_p_spl_00,
    G301_o2_p_spl_0
  );


  buf

  (
    G301_o2_p_spl_01,
    G301_o2_p_spl_0
  );


  buf

  (
    G301_o2_p_spl_1,
    G301_o2_p_spl_
  );


  buf

  (
    G313_o2_n_spl_,
    G313_o2_n
  );


  buf

  (
    G313_o2_n_spl_0,
    G313_o2_n_spl_
  );


  buf

  (
    G313_o2_n_spl_00,
    G313_o2_n_spl_0
  );


  buf

  (
    G313_o2_n_spl_000,
    G313_o2_n_spl_00
  );


  buf

  (
    G313_o2_n_spl_001,
    G313_o2_n_spl_00
  );


  buf

  (
    G313_o2_n_spl_01,
    G313_o2_n_spl_0
  );


  buf

  (
    G313_o2_n_spl_1,
    G313_o2_n_spl_
  );


  buf

  (
    G313_o2_n_spl_10,
    G313_o2_n_spl_1
  );


  buf

  (
    G313_o2_n_spl_11,
    G313_o2_n_spl_1
  );


  buf

  (
    G313_o2_p_spl_,
    G313_o2_p
  );


  buf

  (
    G313_o2_p_spl_0,
    G313_o2_p_spl_
  );


  buf

  (
    G313_o2_p_spl_00,
    G313_o2_p_spl_0
  );


  buf

  (
    G313_o2_p_spl_01,
    G313_o2_p_spl_0
  );


  buf

  (
    G313_o2_p_spl_1,
    G313_o2_p_spl_
  );


  buf

  (
    G1636_o2_p_spl_,
    G1636_o2_p
  );


  buf

  (
    G1636_o2_p_spl_0,
    G1636_o2_p_spl_
  );


  buf

  (
    G1636_o2_p_spl_00,
    G1636_o2_p_spl_0
  );


  buf

  (
    G1636_o2_p_spl_000,
    G1636_o2_p_spl_00
  );


  buf

  (
    G1636_o2_p_spl_001,
    G1636_o2_p_spl_00
  );


  buf

  (
    G1636_o2_p_spl_01,
    G1636_o2_p_spl_0
  );


  buf

  (
    G1636_o2_p_spl_010,
    G1636_o2_p_spl_01
  );


  buf

  (
    G1636_o2_p_spl_1,
    G1636_o2_p_spl_
  );


  buf

  (
    G1636_o2_p_spl_10,
    G1636_o2_p_spl_1
  );


  buf

  (
    G1636_o2_p_spl_11,
    G1636_o2_p_spl_1
  );


  buf

  (
    n3075_lo_buf_o2_n_spl_,
    n3075_lo_buf_o2_n
  );


  buf

  (
    G1636_o2_n_spl_,
    G1636_o2_n
  );


  buf

  (
    G1636_o2_n_spl_0,
    G1636_o2_n_spl_
  );


  buf

  (
    G1636_o2_n_spl_00,
    G1636_o2_n_spl_0
  );


  buf

  (
    G1636_o2_n_spl_000,
    G1636_o2_n_spl_00
  );


  buf

  (
    G1636_o2_n_spl_001,
    G1636_o2_n_spl_00
  );


  buf

  (
    G1636_o2_n_spl_01,
    G1636_o2_n_spl_0
  );


  buf

  (
    G1636_o2_n_spl_010,
    G1636_o2_n_spl_01
  );


  buf

  (
    G1636_o2_n_spl_1,
    G1636_o2_n_spl_
  );


  buf

  (
    G1636_o2_n_spl_10,
    G1636_o2_n_spl_1
  );


  buf

  (
    G1636_o2_n_spl_11,
    G1636_o2_n_spl_1
  );


  buf

  (
    n3075_lo_buf_o2_p_spl_,
    n3075_lo_buf_o2_p
  );


  buf

  (
    n3075_lo_buf_o2_p_spl_0,
    n3075_lo_buf_o2_p_spl_
  );


  buf

  (
    n3075_lo_buf_o2_p_spl_1,
    n3075_lo_buf_o2_p_spl_
  );


  buf

  (
    n2943_lo_buf_o2_n_spl_,
    n2943_lo_buf_o2_n
  );


  buf

  (
    n2943_lo_buf_o2_p_spl_,
    n2943_lo_buf_o2_p
  );


  buf

  (
    n2943_lo_buf_o2_p_spl_0,
    n2943_lo_buf_o2_p_spl_
  );


  buf

  (
    n2943_lo_buf_o2_p_spl_1,
    n2943_lo_buf_o2_p_spl_
  );


  buf

  (
    G1684_o2_p_spl_,
    G1684_o2_p
  );


  buf

  (
    G1684_o2_p_spl_0,
    G1684_o2_p_spl_
  );


  buf

  (
    G1684_o2_p_spl_00,
    G1684_o2_p_spl_0
  );


  buf

  (
    G1684_o2_p_spl_000,
    G1684_o2_p_spl_00
  );


  buf

  (
    G1684_o2_p_spl_001,
    G1684_o2_p_spl_00
  );


  buf

  (
    G1684_o2_p_spl_01,
    G1684_o2_p_spl_0
  );


  buf

  (
    G1684_o2_p_spl_010,
    G1684_o2_p_spl_01
  );


  buf

  (
    G1684_o2_p_spl_1,
    G1684_o2_p_spl_
  );


  buf

  (
    G1684_o2_p_spl_10,
    G1684_o2_p_spl_1
  );


  buf

  (
    G1684_o2_p_spl_11,
    G1684_o2_p_spl_1
  );


  buf

  (
    G1684_o2_n_spl_,
    G1684_o2_n
  );


  buf

  (
    G1684_o2_n_spl_0,
    G1684_o2_n_spl_
  );


  buf

  (
    G1684_o2_n_spl_00,
    G1684_o2_n_spl_0
  );


  buf

  (
    G1684_o2_n_spl_000,
    G1684_o2_n_spl_00
  );


  buf

  (
    G1684_o2_n_spl_001,
    G1684_o2_n_spl_00
  );


  buf

  (
    G1684_o2_n_spl_01,
    G1684_o2_n_spl_0
  );


  buf

  (
    G1684_o2_n_spl_010,
    G1684_o2_n_spl_01
  );


  buf

  (
    G1684_o2_n_spl_1,
    G1684_o2_n_spl_
  );


  buf

  (
    G1684_o2_n_spl_10,
    G1684_o2_n_spl_1
  );


  buf

  (
    G1684_o2_n_spl_11,
    G1684_o2_n_spl_1
  );


  buf

  (
    g1097_n_spl_,
    g1097_n
  );


  buf

  (
    g1097_n_spl_0,
    g1097_n_spl_
  );


  buf

  (
    g1097_n_spl_1,
    g1097_n_spl_
  );


  buf

  (
    g1100_n_spl_,
    g1100_n
  );


  buf

  (
    g1100_n_spl_0,
    g1100_n_spl_
  );


  buf

  (
    g1104_n_spl_,
    g1104_n
  );


  buf

  (
    g1113_n_spl_,
    g1113_n
  );


  buf

  (
    g1113_n_spl_0,
    g1113_n_spl_
  );


  buf

  (
    g1113_n_spl_00,
    g1113_n_spl_0
  );


  buf

  (
    g1113_n_spl_1,
    g1113_n_spl_
  );


  buf

  (
    g1113_p_spl_,
    g1113_p
  );


  buf

  (
    g1113_p_spl_0,
    g1113_p_spl_
  );


  buf

  (
    g1113_p_spl_00,
    g1113_p_spl_0
  );


  buf

  (
    g1113_p_spl_1,
    g1113_p_spl_
  );


  buf

  (
    g1116_n_spl_,
    g1116_n
  );


  buf

  (
    g1116_n_spl_0,
    g1116_n_spl_
  );


  buf

  (
    g1116_n_spl_1,
    g1116_n_spl_
  );


  buf

  (
    g1116_p_spl_,
    g1116_p
  );


  buf

  (
    g1116_p_spl_0,
    g1116_p_spl_
  );


  buf

  (
    g1116_p_spl_1,
    g1116_p_spl_
  );


  buf

  (
    g1120_n_spl_,
    g1120_n
  );


  buf

  (
    g1120_n_spl_0,
    g1120_n_spl_
  );


  buf

  (
    g1120_p_spl_,
    g1120_p
  );


  buf

  (
    g1120_p_spl_0,
    g1120_p_spl_
  );


  buf

  (
    G1336_o2_p_spl_,
    G1336_o2_p
  );


  buf

  (
    G1336_o2_n_spl_,
    G1336_o2_n
  );


  buf

  (
    g1125_n_spl_,
    g1125_n
  );


  buf

  (
    g1125_p_spl_,
    g1125_p
  );


  buf

  (
    G1329_o2_p_spl_,
    G1329_o2_p
  );


  buf

  (
    G1329_o2_p_spl_0,
    G1329_o2_p_spl_
  );


  buf

  (
    G1329_o2_n_spl_,
    G1329_o2_n
  );


  buf

  (
    G1329_o2_n_spl_0,
    G1329_o2_n_spl_
  );


  buf

  (
    G2414_o2_n_spl_,
    G2414_o2_n
  );


  buf

  (
    G2414_o2_p_spl_,
    G2414_o2_p
  );


  buf

  (
    g1111_n_spl_,
    g1111_n
  );


  buf

  (
    g1159_n_spl_,
    g1159_n
  );


  buf

  (
    g1159_n_spl_0,
    g1159_n_spl_
  );


  buf

  (
    g1159_n_spl_1,
    g1159_n_spl_
  );


  buf

  (
    g1162_n_spl_,
    g1162_n
  );


  buf

  (
    g1162_n_spl_0,
    g1162_n_spl_
  );


  buf

  (
    g1166_n_spl_,
    g1166_n
  );


  buf

  (
    g1175_n_spl_,
    g1175_n
  );


  buf

  (
    g1175_n_spl_0,
    g1175_n_spl_
  );


  buf

  (
    g1175_n_spl_00,
    g1175_n_spl_0
  );


  buf

  (
    g1175_n_spl_1,
    g1175_n_spl_
  );


  buf

  (
    g1175_p_spl_,
    g1175_p
  );


  buf

  (
    g1175_p_spl_0,
    g1175_p_spl_
  );


  buf

  (
    g1175_p_spl_00,
    g1175_p_spl_0
  );


  buf

  (
    g1175_p_spl_1,
    g1175_p_spl_
  );


  buf

  (
    g1178_n_spl_,
    g1178_n
  );


  buf

  (
    g1178_n_spl_0,
    g1178_n_spl_
  );


  buf

  (
    g1178_n_spl_1,
    g1178_n_spl_
  );


  buf

  (
    g1178_p_spl_,
    g1178_p
  );


  buf

  (
    g1178_p_spl_0,
    g1178_p_spl_
  );


  buf

  (
    g1178_p_spl_1,
    g1178_p_spl_
  );


  buf

  (
    g1182_n_spl_,
    g1182_n
  );


  buf

  (
    g1182_n_spl_0,
    g1182_n_spl_
  );


  buf

  (
    g1182_p_spl_,
    g1182_p
  );


  buf

  (
    g1182_p_spl_0,
    g1182_p_spl_
  );


  buf

  (
    g1187_n_spl_,
    g1187_n
  );


  buf

  (
    g1187_p_spl_,
    g1187_p
  );


  buf

  (
    G2428_o2_n_spl_,
    G2428_o2_n
  );


  buf

  (
    G2428_o2_p_spl_,
    G2428_o2_p
  );


  buf

  (
    g1173_n_spl_,
    g1173_n
  );


  buf

  (
    G1345_o2_p_spl_,
    G1345_o2_p
  );


  buf

  (
    G1342_o2_n_spl_,
    G1342_o2_n
  );


  buf

  (
    G1345_o2_n_spl_,
    G1345_o2_n
  );


  buf

  (
    G1342_o2_p_spl_,
    G1342_o2_p
  );


  buf

  (
    G1351_o2_p_spl_,
    G1351_o2_p
  );


  buf

  (
    G1348_o2_n_spl_,
    G1348_o2_n
  );


  buf

  (
    G1351_o2_n_spl_,
    G1351_o2_n
  );


  buf

  (
    G1348_o2_p_spl_,
    G1348_o2_p
  );


  buf

  (
    n3270_lo_p_spl_,
    n3270_lo_p
  );


  buf

  (
    n3258_lo_n_spl_,
    n3258_lo_n
  );


  buf

  (
    n3270_lo_n_spl_,
    n3270_lo_n
  );


  buf

  (
    n3258_lo_p_spl_,
    n3258_lo_p
  );


  buf

  (
    n2910_lo_buf_o2_n_spl_,
    n2910_lo_buf_o2_n
  );


  buf

  (
    n2922_lo_buf_o2_p_spl_,
    n2922_lo_buf_o2_p
  );


  buf

  (
    n2910_lo_buf_o2_p_spl_,
    n2910_lo_buf_o2_p
  );


  buf

  (
    n2922_lo_buf_o2_n_spl_,
    n2922_lo_buf_o2_n
  );


  buf

  (
    G1049_o2_p_spl_,
    G1049_o2_p
  );


  buf

  (
    G1049_o2_p_spl_0,
    G1049_o2_p_spl_
  );


  buf

  (
    G1049_o2_p_spl_1,
    G1049_o2_p_spl_
  );


  buf

  (
    n5222_o2_n_spl_,
    n5222_o2_n
  );


  buf

  (
    G1049_o2_n_spl_,
    G1049_o2_n
  );


  buf

  (
    n5222_o2_p_spl_,
    n5222_o2_p
  );


  buf

  (
    n5222_o2_p_spl_0,
    n5222_o2_p_spl_
  );


  buf

  (
    n5222_o2_p_spl_1,
    n5222_o2_p_spl_
  );


  buf

  (
    n2003_inv_n_spl_,
    n2003_inv_n
  );


  buf

  (
    G1053_o2_n_spl_,
    G1053_o2_n
  );


  buf

  (
    n2003_inv_p_spl_,
    n2003_inv_p
  );


  buf

  (
    n2003_inv_p_spl_0,
    n2003_inv_p_spl_
  );


  buf

  (
    G1053_o2_p_spl_,
    G1053_o2_p
  );


  buf

  (
    G1053_o2_p_spl_0,
    G1053_o2_p_spl_
  );


  buf

  (
    g1228_n_spl_,
    g1228_n
  );


  buf

  (
    g1228_n_spl_0,
    g1228_n_spl_
  );


  buf

  (
    g1231_n_spl_,
    g1231_n
  );


  buf

  (
    g1231_n_spl_0,
    g1231_n_spl_
  );


  buf

  (
    n3198_lo_buf_o2_p_spl_,
    n3198_lo_buf_o2_p
  );


  buf

  (
    n3186_lo_buf_o2_n_spl_,
    n3186_lo_buf_o2_n
  );


  buf

  (
    n3198_lo_buf_o2_n_spl_,
    n3198_lo_buf_o2_n
  );


  buf

  (
    n3186_lo_buf_o2_p_spl_,
    n3186_lo_buf_o2_p
  );


  buf

  (
    n3222_lo_buf_o2_p_spl_,
    n3222_lo_buf_o2_p
  );


  buf

  (
    n3210_lo_buf_o2_n_spl_,
    n3210_lo_buf_o2_n
  );


  buf

  (
    n3222_lo_buf_o2_n_spl_,
    n3222_lo_buf_o2_n
  );


  buf

  (
    n3210_lo_buf_o2_p_spl_,
    n3210_lo_buf_o2_p
  );


  buf

  (
    g1258_n_spl_,
    g1258_n
  );


  buf

  (
    g1255_p_spl_,
    g1255_p
  );


  buf

  (
    g1261_p_spl_,
    g1261_p
  );


  buf

  (
    g1255_n_spl_,
    g1255_n
  );


  buf

  (
    g1261_n_spl_,
    g1261_n
  );


  buf

  (
    g1258_p_spl_,
    g1258_p
  );


  buf

  (
    G1079_o2_p_spl_,
    G1079_o2_p
  );


  buf

  (
    G1222_o2_p_spl_,
    G1222_o2_p
  );


  buf

  (
    G1079_o2_n_spl_,
    G1079_o2_n
  );


  buf

  (
    G1222_o2_n_spl_,
    G1222_o2_n
  );


  buf

  (
    G1228_o2_n_spl_,
    G1228_o2_n
  );


  buf

  (
    G1225_o2_p_spl_,
    G1225_o2_p
  );


  buf

  (
    G1228_o2_p_spl_,
    G1228_o2_p
  );


  buf

  (
    G1225_o2_n_spl_,
    G1225_o2_n
  );


  buf

  (
    g1278_p_spl_,
    g1278_p
  );


  buf

  (
    g1275_n_spl_,
    g1275_n
  );


  buf

  (
    g1281_n_spl_,
    g1281_n
  );


  buf

  (
    g1275_p_spl_,
    g1275_p
  );


  buf

  (
    g1281_p_spl_,
    g1281_p
  );


  buf

  (
    g1278_n_spl_,
    g1278_n
  );


  buf

  (
    G1371_o2_p_spl_,
    G1371_o2_p
  );


  buf

  (
    G1368_o2_n_spl_,
    G1368_o2_n
  );


  buf

  (
    G1371_o2_n_spl_,
    G1371_o2_n
  );


  buf

  (
    G1368_o2_p_spl_,
    G1368_o2_p
  );


  buf

  (
    G1537_o2_p_spl_,
    G1537_o2_p
  );


  buf

  (
    G1374_o2_p_spl_,
    G1374_o2_p
  );


  buf

  (
    G1537_o2_n_spl_,
    G1537_o2_n
  );


  buf

  (
    G1374_o2_n_spl_,
    G1374_o2_n
  );


  buf

  (
    g1298_n_spl_,
    g1298_n
  );


  buf

  (
    g1295_p_spl_,
    g1295_p
  );


  buf

  (
    g1301_p_spl_,
    g1301_p
  );


  buf

  (
    g1295_n_spl_,
    g1295_n
  );


  buf

  (
    g1301_n_spl_,
    g1301_n
  );


  buf

  (
    g1298_p_spl_,
    g1298_p
  );


  buf

  (
    n3087_lo_n_spl_,
    n3087_lo_n
  );


  buf

  (
    n2955_lo_n_spl_,
    n2955_lo_n
  );


  buf

  (
    n2991_lo_p_spl_,
    n2991_lo_p
  );


  buf

  (
    n2991_lo_p_spl_0,
    n2991_lo_p_spl_
  );


  buf

  (
    n2991_lo_p_spl_1,
    n2991_lo_p_spl_
  );


  buf

  (
    n1503_lo_buf_o2_n_spl_,
    n1503_lo_buf_o2_n
  );


  buf

  (
    n1503_lo_buf_o2_n_spl_0,
    n1503_lo_buf_o2_n_spl_
  );


  buf

  (
    n1503_lo_buf_o2_n_spl_00,
    n1503_lo_buf_o2_n_spl_0
  );


  buf

  (
    n1503_lo_buf_o2_n_spl_000,
    n1503_lo_buf_o2_n_spl_00
  );


  buf

  (
    n1503_lo_buf_o2_n_spl_001,
    n1503_lo_buf_o2_n_spl_00
  );


  buf

  (
    n1503_lo_buf_o2_n_spl_01,
    n1503_lo_buf_o2_n_spl_0
  );


  buf

  (
    n1503_lo_buf_o2_n_spl_010,
    n1503_lo_buf_o2_n_spl_01
  );


  buf

  (
    n1503_lo_buf_o2_n_spl_011,
    n1503_lo_buf_o2_n_spl_01
  );


  buf

  (
    n1503_lo_buf_o2_n_spl_1,
    n1503_lo_buf_o2_n_spl_
  );


  buf

  (
    n1503_lo_buf_o2_n_spl_10,
    n1503_lo_buf_o2_n_spl_1
  );


  buf

  (
    n1503_lo_buf_o2_n_spl_100,
    n1503_lo_buf_o2_n_spl_10
  );


  buf

  (
    n1503_lo_buf_o2_n_spl_101,
    n1503_lo_buf_o2_n_spl_10
  );


  buf

  (
    n1503_lo_buf_o2_n_spl_11,
    n1503_lo_buf_o2_n_spl_1
  );


  buf

  (
    n1503_lo_buf_o2_n_spl_110,
    n1503_lo_buf_o2_n_spl_11
  );


  buf

  (
    n1503_lo_buf_o2_n_spl_111,
    n1503_lo_buf_o2_n_spl_11
  );


  buf

  (
    n3003_lo_p_spl_,
    n3003_lo_p
  );


  buf

  (
    n3003_lo_p_spl_0,
    n3003_lo_p_spl_
  );


  buf

  (
    n3003_lo_p_spl_1,
    n3003_lo_p_spl_
  );


  buf

  (
    n3063_lo_buf_o2_p_spl_,
    n3063_lo_buf_o2_p
  );


  buf

  (
    n3063_lo_buf_o2_p_spl_0,
    n3063_lo_buf_o2_p_spl_
  );


  buf

  (
    n3063_lo_buf_o2_p_spl_00,
    n3063_lo_buf_o2_p_spl_0
  );


  buf

  (
    n3063_lo_buf_o2_p_spl_01,
    n3063_lo_buf_o2_p_spl_0
  );


  buf

  (
    n3063_lo_buf_o2_p_spl_1,
    n3063_lo_buf_o2_p_spl_
  );


  buf

  (
    g1329_n_spl_,
    g1329_n
  );


  buf

  (
    g1329_n_spl_0,
    g1329_n_spl_
  );


  buf

  (
    g1329_n_spl_1,
    g1329_n_spl_
  );


  buf

  (
    n3027_lo_n_spl_,
    n3027_lo_n
  );


  buf

  (
    g1329_p_spl_,
    g1329_p
  );


  buf

  (
    g1329_p_spl_0,
    g1329_p_spl_
  );


  buf

  (
    g1329_p_spl_00,
    g1329_p_spl_0
  );


  buf

  (
    g1329_p_spl_01,
    g1329_p_spl_0
  );


  buf

  (
    g1329_p_spl_1,
    g1329_p_spl_
  );


  buf

  (
    g1329_p_spl_10,
    g1329_p_spl_1
  );


  buf

  (
    g1329_p_spl_11,
    g1329_p_spl_1
  );


  buf

  (
    n3039_lo_n_spl_,
    n3039_lo_n
  );


  buf

  (
    n3099_lo_buf_o2_p_spl_,
    n3099_lo_buf_o2_p
  );


  buf

  (
    n3099_lo_buf_o2_p_spl_0,
    n3099_lo_buf_o2_p_spl_
  );


  buf

  (
    n3099_lo_buf_o2_p_spl_1,
    n3099_lo_buf_o2_p_spl_
  );


  buf

  (
    n2967_lo_buf_o2_p_spl_,
    n2967_lo_buf_o2_p
  );


  buf

  (
    n2967_lo_buf_o2_p_spl_0,
    n2967_lo_buf_o2_p_spl_
  );


  buf

  (
    n2967_lo_buf_o2_p_spl_1,
    n2967_lo_buf_o2_p_spl_
  );


  buf

  (
    n3111_lo_buf_o2_p_spl_,
    n3111_lo_buf_o2_p
  );


  buf

  (
    n3111_lo_buf_o2_p_spl_0,
    n3111_lo_buf_o2_p_spl_
  );


  buf

  (
    n3111_lo_buf_o2_p_spl_1,
    n3111_lo_buf_o2_p_spl_
  );


  buf

  (
    n2979_lo_buf_o2_p_spl_,
    n2979_lo_buf_o2_p
  );


  buf

  (
    n2979_lo_buf_o2_p_spl_0,
    n2979_lo_buf_o2_p_spl_
  );


  buf

  (
    n2979_lo_buf_o2_p_spl_1,
    n2979_lo_buf_o2_p_spl_
  );


  buf

  (
    g1020_n_spl_,
    g1020_n
  );


  buf

  (
    g1020_n_spl_0,
    g1020_n_spl_
  );


  buf

  (
    g1020_n_spl_00,
    g1020_n_spl_0
  );


  buf

  (
    g1020_n_spl_1,
    g1020_n_spl_
  );


  buf

  (
    G1493_o2_n_spl_,
    G1493_o2_n
  );


  buf

  (
    G1493_o2_n_spl_0,
    G1493_o2_n_spl_
  );


  buf

  (
    G1493_o2_n_spl_1,
    G1493_o2_n_spl_
  );


  buf

  (
    g1017_n_spl_,
    g1017_n
  );


  buf

  (
    g1017_n_spl_0,
    g1017_n_spl_
  );


  buf

  (
    g1017_n_spl_00,
    g1017_n_spl_0
  );


  buf

  (
    g1017_n_spl_1,
    g1017_n_spl_
  );


  buf

  (
    G1498_o2_n_spl_,
    G1498_o2_n
  );


  buf

  (
    G1498_o2_n_spl_0,
    G1498_o2_n_spl_
  );


  buf

  (
    G1498_o2_n_spl_1,
    G1498_o2_n_spl_
  );


  buf

  (
    g1045_n_spl_,
    g1045_n
  );


  buf

  (
    g1045_n_spl_0,
    g1045_n_spl_
  );


  buf

  (
    G1314_o2_n_spl_,
    G1314_o2_n
  );


  buf

  (
    g1056_n_spl_,
    g1056_n
  );


  buf

  (
    g1056_n_spl_0,
    g1056_n_spl_
  );


  buf

  (
    g1023_n_spl_,
    g1023_n
  );


  buf

  (
    g1023_n_spl_0,
    g1023_n_spl_
  );


  buf

  (
    G1314_o2_p_spl_,
    G1314_o2_p
  );


  buf

  (
    G1021_o2_p_spl_,
    G1021_o2_p
  );


  buf

  (
    G1021_o2_p_spl_0,
    G1021_o2_p_spl_
  );


  buf

  (
    G1021_o2_p_spl_00,
    G1021_o2_p_spl_0
  );


  buf

  (
    G1021_o2_p_spl_01,
    G1021_o2_p_spl_0
  );


  buf

  (
    G1021_o2_p_spl_1,
    G1021_o2_p_spl_
  );


  buf

  (
    G1021_o2_p_spl_10,
    G1021_o2_p_spl_1
  );


  buf

  (
    G1021_o2_p_spl_11,
    G1021_o2_p_spl_1
  );


  buf

  (
    G1493_o2_p_spl_,
    G1493_o2_p
  );


  buf

  (
    G1026_o2_p_spl_,
    G1026_o2_p
  );


  buf

  (
    G1026_o2_p_spl_0,
    G1026_o2_p_spl_
  );


  buf

  (
    G1026_o2_p_spl_00,
    G1026_o2_p_spl_0
  );


  buf

  (
    G1026_o2_p_spl_01,
    G1026_o2_p_spl_0
  );


  buf

  (
    G1026_o2_p_spl_1,
    G1026_o2_p_spl_
  );


  buf

  (
    G1026_o2_p_spl_10,
    G1026_o2_p_spl_1
  );


  buf

  (
    G1498_o2_p_spl_,
    G1498_o2_p
  );


  buf

  (
    n3015_lo_n_spl_,
    n3015_lo_n
  );


  buf

  (
    g1034_n_spl_,
    g1034_n
  );


  buf

  (
    g1034_n_spl_0,
    g1034_n_spl_
  );


  buf

  (
    g1034_n_spl_1,
    g1034_n_spl_
  );


  buf

  (
    n3150_lo_buf_o2_p_spl_,
    n3150_lo_buf_o2_p
  );


  buf

  (
    n3150_lo_buf_o2_p_spl_0,
    n3150_lo_buf_o2_p_spl_
  );


  buf

  (
    n3150_lo_buf_o2_p_spl_00,
    n3150_lo_buf_o2_p_spl_0
  );


  buf

  (
    n3150_lo_buf_o2_p_spl_000,
    n3150_lo_buf_o2_p_spl_00
  );


  buf

  (
    n3150_lo_buf_o2_p_spl_001,
    n3150_lo_buf_o2_p_spl_00
  );


  buf

  (
    n3150_lo_buf_o2_p_spl_01,
    n3150_lo_buf_o2_p_spl_0
  );


  buf

  (
    n3150_lo_buf_o2_p_spl_1,
    n3150_lo_buf_o2_p_spl_
  );


  buf

  (
    n3150_lo_buf_o2_p_spl_10,
    n3150_lo_buf_o2_p_spl_1
  );


  buf

  (
    n3150_lo_buf_o2_p_spl_11,
    n3150_lo_buf_o2_p_spl_1
  );


  buf

  (
    n3162_lo_buf_o2_p_spl_,
    n3162_lo_buf_o2_p
  );


  buf

  (
    n3162_lo_buf_o2_p_spl_0,
    n3162_lo_buf_o2_p_spl_
  );


  buf

  (
    n3162_lo_buf_o2_p_spl_00,
    n3162_lo_buf_o2_p_spl_0
  );


  buf

  (
    n3162_lo_buf_o2_p_spl_000,
    n3162_lo_buf_o2_p_spl_00
  );


  buf

  (
    n3162_lo_buf_o2_p_spl_001,
    n3162_lo_buf_o2_p_spl_00
  );


  buf

  (
    n3162_lo_buf_o2_p_spl_01,
    n3162_lo_buf_o2_p_spl_0
  );


  buf

  (
    n3162_lo_buf_o2_p_spl_1,
    n3162_lo_buf_o2_p_spl_
  );


  buf

  (
    n3162_lo_buf_o2_p_spl_10,
    n3162_lo_buf_o2_p_spl_1
  );


  buf

  (
    n3162_lo_buf_o2_p_spl_11,
    n3162_lo_buf_o2_p_spl_1
  );


  buf

  (
    n3150_lo_buf_o2_n_spl_,
    n3150_lo_buf_o2_n
  );


  buf

  (
    n3150_lo_buf_o2_n_spl_0,
    n3150_lo_buf_o2_n_spl_
  );


  buf

  (
    n3150_lo_buf_o2_n_spl_00,
    n3150_lo_buf_o2_n_spl_0
  );


  buf

  (
    n3150_lo_buf_o2_n_spl_01,
    n3150_lo_buf_o2_n_spl_0
  );


  buf

  (
    n3150_lo_buf_o2_n_spl_1,
    n3150_lo_buf_o2_n_spl_
  );


  buf

  (
    n3162_lo_buf_o2_n_spl_,
    n3162_lo_buf_o2_n
  );


  buf

  (
    n3162_lo_buf_o2_n_spl_0,
    n3162_lo_buf_o2_n_spl_
  );


  buf

  (
    n3162_lo_buf_o2_n_spl_00,
    n3162_lo_buf_o2_n_spl_0
  );


  buf

  (
    n3162_lo_buf_o2_n_spl_01,
    n3162_lo_buf_o2_n_spl_0
  );


  buf

  (
    n3162_lo_buf_o2_n_spl_1,
    n3162_lo_buf_o2_n_spl_
  );


  buf

  (
    n2958_lo_buf_o2_n_spl_,
    n2958_lo_buf_o2_n
  );


  buf

  (
    n2970_lo_buf_o2_p_spl_,
    n2970_lo_buf_o2_p
  );


  buf

  (
    n2958_lo_buf_o2_p_spl_,
    n2958_lo_buf_o2_p
  );


  buf

  (
    n2970_lo_buf_o2_n_spl_,
    n2970_lo_buf_o2_n
  );


  buf

  (
    n2946_lo_buf_o2_p_spl_,
    n2946_lo_buf_o2_p
  );


  buf

  (
    n3282_lo_p_spl_,
    n3282_lo_p
  );


  buf

  (
    n2946_lo_buf_o2_n_spl_,
    n2946_lo_buf_o2_n
  );


  buf

  (
    n3282_lo_n_spl_,
    n3282_lo_n
  );


  buf

  (
    g1453_p_spl_,
    g1453_p
  );


  buf

  (
    g1450_p_spl_,
    g1450_p
  );


  buf

  (
    g1456_n_spl_,
    g1456_n
  );


  buf

  (
    g1456_n_spl_0,
    g1456_n_spl_
  );


  buf

  (
    g1456_n_spl_1,
    g1456_n_spl_
  );


  buf

  (
    g1453_n_spl_,
    g1453_n
  );


  buf

  (
    n3090_lo_buf_o2_p_spl_,
    n3090_lo_buf_o2_p
  );


  buf

  (
    n3090_lo_buf_o2_p_spl_0,
    n3090_lo_buf_o2_p_spl_
  );


  buf

  (
    n3078_lo_buf_o2_n_spl_,
    n3078_lo_buf_o2_n
  );


  buf

  (
    n3090_lo_buf_o2_n_spl_,
    n3090_lo_buf_o2_n
  );


  buf

  (
    n3078_lo_buf_o2_p_spl_,
    n3078_lo_buf_o2_p
  );


  buf

  (
    n3078_lo_buf_o2_p_spl_0,
    n3078_lo_buf_o2_p_spl_
  );


  buf

  (
    n3066_lo_buf_o2_p_spl_,
    n3066_lo_buf_o2_p
  );


  buf

  (
    n3294_lo_p_spl_,
    n3294_lo_p
  );


  buf

  (
    n3066_lo_buf_o2_n_spl_,
    n3066_lo_buf_o2_n
  );


  buf

  (
    n3294_lo_n_spl_,
    n3294_lo_n
  );


  buf

  (
    n3114_lo_buf_o2_p_spl_,
    n3114_lo_buf_o2_p
  );


  buf

  (
    n3102_lo_buf_o2_p_spl_,
    n3102_lo_buf_o2_p
  );


  buf

  (
    g1466_p_spl_,
    g1466_p
  );


  buf

  (
    g1463_p_spl_,
    g1463_p
  );


  buf

  (
    g1469_n_spl_,
    g1469_n
  );


  buf

  (
    g1469_n_spl_0,
    g1469_n_spl_
  );


  buf

  (
    g1469_n_spl_1,
    g1469_n_spl_
  );


  buf

  (
    g1466_n_spl_,
    g1466_n
  );


  buf

  (
    g1450_n_spl_,
    g1450_n
  );


  buf

  (
    g1463_n_spl_,
    g1463_n
  );


  buf

  (
    G1129_o2_p_spl_,
    G1129_o2_p
  );


  buf

  (
    G1132_o2_n_spl_,
    G1132_o2_n
  );


  buf

  (
    G1129_o2_n_spl_,
    G1129_o2_n
  );


  buf

  (
    G1132_o2_p_spl_,
    G1132_o2_p
  );


  buf

  (
    g1480_p_spl_,
    g1480_p
  );


  buf

  (
    g1014_n_spl_,
    g1014_n
  );


  buf

  (
    g1014_n_spl_0,
    g1014_n_spl_
  );


  buf

  (
    g1014_n_spl_1,
    g1014_n_spl_
  );


  buf

  (
    g1483_n_spl_,
    g1483_n
  );


  buf

  (
    g1483_n_spl_0,
    g1483_n_spl_
  );


  buf

  (
    g1483_n_spl_1,
    g1483_n_spl_
  );


  buf

  (
    g1480_n_spl_,
    g1480_n
  );


  buf

  (
    g1014_p_spl_,
    g1014_p
  );


  buf

  (
    n1554_lo_p_spl_,
    n1554_lo_p
  );


  buf

  (
    n1554_lo_p_spl_0,
    n1554_lo_p_spl_
  );


  buf

  (
    n1554_lo_p_spl_00,
    n1554_lo_p_spl_0
  );


  buf

  (
    n1554_lo_p_spl_000,
    n1554_lo_p_spl_00
  );


  buf

  (
    n1554_lo_p_spl_01,
    n1554_lo_p_spl_0
  );


  buf

  (
    n1554_lo_p_spl_1,
    n1554_lo_p_spl_
  );


  buf

  (
    n1554_lo_p_spl_10,
    n1554_lo_p_spl_1
  );


  buf

  (
    n1554_lo_p_spl_11,
    n1554_lo_p_spl_1
  );


  buf

  (
    n1554_lo_n_spl_,
    n1554_lo_n
  );


  buf

  (
    n1554_lo_n_spl_0,
    n1554_lo_n_spl_
  );


  buf

  (
    n1554_lo_n_spl_00,
    n1554_lo_n_spl_0
  );


  buf

  (
    n1554_lo_n_spl_000,
    n1554_lo_n_spl_00
  );


  buf

  (
    n1554_lo_n_spl_01,
    n1554_lo_n_spl_0
  );


  buf

  (
    n1554_lo_n_spl_1,
    n1554_lo_n_spl_
  );


  buf

  (
    n1554_lo_n_spl_10,
    n1554_lo_n_spl_1
  );


  buf

  (
    n1554_lo_n_spl_11,
    n1554_lo_n_spl_1
  );


  buf

  (
    G1017_o2_p_spl_,
    G1017_o2_p
  );


  buf

  (
    G1002_o2_p_spl_,
    G1002_o2_p
  );


  buf

  (
    G1002_o2_p_spl_0,
    G1002_o2_p_spl_
  );


  buf

  (
    n5554_o2_p_spl_,
    n5554_o2_p
  );


  buf

  (
    n5553_o2_p_spl_,
    n5553_o2_p
  );


  buf

  (
    n1686_lo_p_spl_,
    n1686_lo_p
  );


  buf

  (
    n1686_lo_p_spl_0,
    n1686_lo_p_spl_
  );


  buf

  (
    n1686_lo_p_spl_00,
    n1686_lo_p_spl_0
  );


  buf

  (
    n1686_lo_p_spl_000,
    n1686_lo_p_spl_00
  );


  buf

  (
    n1686_lo_p_spl_01,
    n1686_lo_p_spl_0
  );


  buf

  (
    n1686_lo_p_spl_1,
    n1686_lo_p_spl_
  );


  buf

  (
    n1686_lo_p_spl_10,
    n1686_lo_p_spl_1
  );


  buf

  (
    n1686_lo_p_spl_11,
    n1686_lo_p_spl_1
  );


  buf

  (
    n1686_lo_n_spl_,
    n1686_lo_n
  );


  buf

  (
    n1686_lo_n_spl_0,
    n1686_lo_n_spl_
  );


  buf

  (
    n1686_lo_n_spl_00,
    n1686_lo_n_spl_0
  );


  buf

  (
    n1686_lo_n_spl_01,
    n1686_lo_n_spl_0
  );


  buf

  (
    n1686_lo_n_spl_1,
    n1686_lo_n_spl_
  );


  buf

  (
    n1686_lo_n_spl_10,
    n1686_lo_n_spl_1
  );


  buf

  (
    n5223_o2_p_spl_,
    n5223_o2_p
  );


  buf

  (
    g1219_n_spl_,
    g1219_n
  );


  buf

  (
    g1157_n_spl_,
    g1157_n
  );


  buf

  (
    g1447_p_spl_,
    g1447_p
  );


  buf

  (
    g1548_n_spl_,
    g1548_n
  );


  buf

  (
    g1436_n_spl_,
    g1436_n
  );


  buf

  (
    g1436_n_spl_0,
    g1436_n_spl_
  );


  buf

  (
    n3063_lo_buf_o2_n_spl_,
    n3063_lo_buf_o2_n
  );


  buf

  (
    n2919_lo_buf_o2_n_spl_,
    n2919_lo_buf_o2_n
  );


  buf

  (
    n2919_lo_buf_o2_p_spl_,
    n2919_lo_buf_o2_p
  );


  buf

  (
    n2919_lo_buf_o2_p_spl_0,
    n2919_lo_buf_o2_p_spl_
  );


  buf

  (
    n2919_lo_buf_o2_p_spl_1,
    n2919_lo_buf_o2_p_spl_
  );


  buf

  (
    g1553_p_spl_,
    g1553_p
  );


  buf

  (
    g1089_n_spl_,
    g1089_n
  );


  buf

  (
    g1089_n_spl_0,
    g1089_n_spl_
  );


  buf

  (
    g1089_n_spl_00,
    g1089_n_spl_0
  );


  buf

  (
    g1089_n_spl_01,
    g1089_n_spl_0
  );


  buf

  (
    g1089_n_spl_1,
    g1089_n_spl_
  );


  buf

  (
    g1089_n_spl_10,
    g1089_n_spl_1
  );


  buf

  (
    g1557_p_spl_,
    g1557_p
  );


  buf

  (
    g1315_n_spl_,
    g1315_n
  );


  buf

  (
    g1315_n_spl_0,
    g1315_n_spl_
  );


  buf

  (
    g1078_p_spl_,
    g1078_p
  );


  buf

  (
    g1078_p_spl_0,
    g1078_p_spl_
  );


  buf

  (
    g1078_p_spl_1,
    g1078_p_spl_
  );


  buf

  (
    g1358_n_spl_,
    g1358_n
  );


  buf

  (
    g1358_n_spl_0,
    g1358_n_spl_
  );


  buf

  (
    g1317_n_spl_,
    g1317_n
  );


  buf

  (
    g1317_n_spl_0,
    g1317_n_spl_
  );


  buf

  (
    g1360_n_spl_,
    g1360_n
  );


  buf

  (
    g1360_n_spl_0,
    g1360_n_spl_
  );


  buf

  (
    g1319_n_spl_,
    g1319_n
  );


  buf

  (
    g1319_n_spl_0,
    g1319_n_spl_
  );


  buf

  (
    g1322_n_spl_,
    g1322_n
  );


  buf

  (
    g1322_n_spl_0,
    g1322_n_spl_
  );


  buf

  (
    g1362_n_spl_,
    g1362_n
  );


  buf

  (
    g1362_n_spl_0,
    g1362_n_spl_
  );


  buf

  (
    g1324_n_spl_,
    g1324_n
  );


  buf

  (
    g1324_n_spl_0,
    g1324_n_spl_
  );


  buf

  (
    g1364_n_spl_,
    g1364_n
  );


  buf

  (
    g1364_n_spl_0,
    g1364_n_spl_
  );


  buf

  (
    g1326_n_spl_,
    g1326_n
  );


  buf

  (
    g1326_n_spl_0,
    g1326_n_spl_
  );


  buf

  (
    g1370_n_spl_,
    g1370_n
  );


  buf

  (
    g1370_n_spl_0,
    g1370_n_spl_
  );


  buf

  (
    g1370_n_spl_00,
    g1370_n_spl_0
  );


  buf

  (
    g1370_n_spl_01,
    g1370_n_spl_0
  );


  buf

  (
    g1370_n_spl_1,
    g1370_n_spl_
  );


  buf

  (
    g1330_n_spl_,
    g1330_n
  );


  buf

  (
    g1330_n_spl_0,
    g1330_n_spl_
  );


  buf

  (
    g1332_n_spl_,
    g1332_n
  );


  buf

  (
    g1332_n_spl_0,
    g1332_n_spl_
  );


  buf

  (
    g1366_p_spl_,
    g1366_p
  );


  buf

  (
    g1366_p_spl_0,
    g1366_p_spl_
  );


  buf

  (
    g1366_p_spl_00,
    g1366_p_spl_0
  );


  buf

  (
    g1366_p_spl_01,
    g1366_p_spl_0
  );


  buf

  (
    g1366_p_spl_1,
    g1366_p_spl_
  );


  buf

  (
    g1334_p_spl_,
    g1334_p
  );


  buf

  (
    g1334_p_spl_0,
    g1334_p_spl_
  );


  buf

  (
    g1368_p_spl_,
    g1368_p
  );


  buf

  (
    g1368_p_spl_0,
    g1368_p_spl_
  );


  buf

  (
    g1368_p_spl_00,
    g1368_p_spl_0
  );


  buf

  (
    g1368_p_spl_01,
    g1368_p_spl_0
  );


  buf

  (
    g1368_p_spl_1,
    g1368_p_spl_
  );


  buf

  (
    g1336_p_spl_,
    g1336_p
  );


  buf

  (
    g1336_p_spl_0,
    g1336_p_spl_
  );


  buf

  (
    g1338_p_spl_,
    g1338_p
  );


  buf

  (
    g1338_p_spl_0,
    g1338_p_spl_
  );


  buf

  (
    g1340_p_spl_,
    g1340_p
  );


  buf

  (
    g1340_p_spl_0,
    g1340_p_spl_
  );


  buf

  (
    g1374_n_spl_,
    g1374_n
  );


  buf

  (
    g1374_n_spl_0,
    g1374_n_spl_
  );


  buf

  (
    g1344_n_spl_,
    g1344_n
  );


  buf

  (
    g1344_n_spl_0,
    g1344_n_spl_
  );


  buf

  (
    g1378_n_spl_,
    g1378_n
  );


  buf

  (
    g1378_n_spl_0,
    g1378_n_spl_
  );


  buf

  (
    g1348_n_spl_,
    g1348_n
  );


  buf

  (
    g1348_n_spl_0,
    g1348_n_spl_
  );


  buf

  (
    g1382_n_spl_,
    g1382_n
  );


  buf

  (
    g1382_n_spl_0,
    g1382_n_spl_
  );


  buf

  (
    g1352_n_spl_,
    g1352_n
  );


  buf

  (
    g1352_n_spl_0,
    g1352_n_spl_
  );


  buf

  (
    g1386_n_spl_,
    g1386_n
  );


  buf

  (
    g1386_n_spl_0,
    g1386_n_spl_
  );


  buf

  (
    g1356_n_spl_,
    g1356_n
  );


  buf

  (
    g1356_n_spl_0,
    g1356_n_spl_
  );


  buf

  (
    G663_o2_p_spl_,
    G663_o2_p
  );


  buf

  (
    G663_o2_p_spl_0,
    G663_o2_p_spl_
  );


  buf

  (
    G663_o2_p_spl_1,
    G663_o2_p_spl_
  );


  buf

  (
    G674_o2_p_spl_,
    G674_o2_p
  );


  buf

  (
    G674_o2_p_spl_0,
    G674_o2_p_spl_
  );


  buf

  (
    G674_o2_p_spl_1,
    G674_o2_p_spl_
  );


  buf

  (
    G374_o2_n_spl_,
    G374_o2_n
  );


  buf

  (
    G374_o2_n_spl_0,
    G374_o2_n_spl_
  );


  buf

  (
    G374_o2_n_spl_1,
    G374_o2_n_spl_
  );


  buf

  (
    G386_o2_n_spl_,
    G386_o2_n
  );


  buf

  (
    G386_o2_n_spl_0,
    G386_o2_n_spl_
  );


  buf

  (
    G386_o2_n_spl_1,
    G386_o2_n_spl_
  );


  buf

  (
    G674_o2_n_spl_,
    G674_o2_n
  );


  buf

  (
    G663_o2_n_spl_,
    G663_o2_n
  );


  buf

  (
    G374_o2_p_spl_,
    G374_o2_p
  );


  buf

  (
    G386_o2_p_spl_,
    G386_o2_p
  );


  buf

  (
    g1089_p_spl_,
    g1089_p
  );


  buf

  (
    g1092_p_spl_,
    g1092_p
  );


  buf

  (
    g1067_n_spl_,
    g1067_n
  );


  buf

  (
    g1067_n_spl_0,
    g1067_n_spl_
  );


  buf

  (
    g1067_n_spl_00,
    g1067_n_spl_0
  );


  buf

  (
    g1067_n_spl_01,
    g1067_n_spl_0
  );


  buf

  (
    g1067_n_spl_1,
    g1067_n_spl_
  );


  buf

  (
    g1067_p_spl_,
    g1067_p
  );


  buf

  (
    g1095_p_spl_,
    g1095_p
  );


  buf

  (
    n3039_lo_p_spl_,
    n3039_lo_p
  );


  buf

  (
    n3039_lo_p_spl_0,
    n3039_lo_p_spl_
  );


  buf

  (
    n3039_lo_p_spl_1,
    n3039_lo_p_spl_
  );


  buf

  (
    n2907_lo_p_spl_,
    n2907_lo_p
  );


  buf

  (
    n2907_lo_p_spl_0,
    n2907_lo_p_spl_
  );


  buf

  (
    n2907_lo_p_spl_1,
    n2907_lo_p_spl_
  );


  buf

  (
    g1412_n_spl_,
    g1412_n
  );


  buf

  (
    g1412_n_spl_0,
    g1412_n_spl_
  );


  buf

  (
    g1412_n_spl_00,
    g1412_n_spl_0
  );


  buf

  (
    g1412_n_spl_1,
    g1412_n_spl_
  );


  buf

  (
    n2808_lo_n_spl_,
    n2808_lo_n
  );


  buf

  (
    n2808_lo_n_spl_0,
    n2808_lo_n_spl_
  );


  buf

  (
    n2808_lo_n_spl_00,
    n2808_lo_n_spl_0
  );


  buf

  (
    n2808_lo_n_spl_01,
    n2808_lo_n_spl_0
  );


  buf

  (
    n2808_lo_n_spl_1,
    n2808_lo_n_spl_
  );


  buf

  (
    n2808_lo_n_spl_10,
    n2808_lo_n_spl_1
  );


  buf

  (
    n2808_lo_n_spl_11,
    n2808_lo_n_spl_1
  );


  buf

  (
    n2844_lo_p_spl_,
    n2844_lo_p
  );


  buf

  (
    n2844_lo_p_spl_0,
    n2844_lo_p_spl_
  );


  buf

  (
    n2844_lo_p_spl_00,
    n2844_lo_p_spl_0
  );


  buf

  (
    n2844_lo_p_spl_000,
    n2844_lo_p_spl_00
  );


  buf

  (
    n2844_lo_p_spl_001,
    n2844_lo_p_spl_00
  );


  buf

  (
    n2844_lo_p_spl_01,
    n2844_lo_p_spl_0
  );


  buf

  (
    n2844_lo_p_spl_010,
    n2844_lo_p_spl_01
  );


  buf

  (
    n2844_lo_p_spl_011,
    n2844_lo_p_spl_01
  );


  buf

  (
    n2844_lo_p_spl_1,
    n2844_lo_p_spl_
  );


  buf

  (
    n2844_lo_p_spl_10,
    n2844_lo_p_spl_1
  );


  buf

  (
    n2844_lo_p_spl_11,
    n2844_lo_p_spl_1
  );


  buf

  (
    n2844_lo_n_spl_,
    n2844_lo_n
  );


  buf

  (
    n2844_lo_n_spl_0,
    n2844_lo_n_spl_
  );


  buf

  (
    n2844_lo_n_spl_00,
    n2844_lo_n_spl_0
  );


  buf

  (
    n2844_lo_n_spl_01,
    n2844_lo_n_spl_0
  );


  buf

  (
    n2844_lo_n_spl_1,
    n2844_lo_n_spl_
  );


  buf

  (
    n2844_lo_n_spl_10,
    n2844_lo_n_spl_1
  );


  buf

  (
    n2844_lo_n_spl_11,
    n2844_lo_n_spl_1
  );


  buf

  (
    n2808_lo_p_spl_,
    n2808_lo_p
  );


  buf

  (
    n2808_lo_p_spl_0,
    n2808_lo_p_spl_
  );


  buf

  (
    n2808_lo_p_spl_00,
    n2808_lo_p_spl_0
  );


  buf

  (
    n2808_lo_p_spl_000,
    n2808_lo_p_spl_00
  );


  buf

  (
    n2808_lo_p_spl_001,
    n2808_lo_p_spl_00
  );


  buf

  (
    n2808_lo_p_spl_01,
    n2808_lo_p_spl_0
  );


  buf

  (
    n2808_lo_p_spl_010,
    n2808_lo_p_spl_01
  );


  buf

  (
    n2808_lo_p_spl_011,
    n2808_lo_p_spl_01
  );


  buf

  (
    n2808_lo_p_spl_1,
    n2808_lo_p_spl_
  );


  buf

  (
    n2808_lo_p_spl_10,
    n2808_lo_p_spl_1
  );


  buf

  (
    n2808_lo_p_spl_11,
    n2808_lo_p_spl_1
  );


  buf

  (
    n2901_lo_n_spl_,
    n2901_lo_n
  );


  buf

  (
    n3057_lo_n_spl_,
    n3057_lo_n
  );


  buf

  (
    n3057_lo_n_spl_0,
    n3057_lo_n_spl_
  );


  buf

  (
    g850_n_spl_,
    g850_n
  );


  buf

  (
    g864_p_spl_,
    g864_p
  );


  buf

  (
    g867_p_spl_,
    g867_p
  );


  buf

  (
    g873_p_spl_,
    g873_p
  );


  buf

  (
    g975_n_spl_,
    g975_n
  );


  buf

  (
    g1000_p_spl_,
    g1000_p
  );


  buf

  (
    g1013_n_spl_,
    g1013_n
  );


  buf

  (
    n3126_lo_p_spl_,
    n3126_lo_p
  );


  buf

  (
    n3126_lo_p_spl_0,
    n3126_lo_p_spl_
  );


  buf

  (
    n3138_lo_p_spl_,
    n3138_lo_p
  );


  buf

  (
    n3138_lo_p_spl_0,
    n3138_lo_p_spl_
  );


  buf

  (
    G1039_o2_p_spl_,
    G1039_o2_p
  );


  buf

  (
    G1039_o2_p_spl_0,
    G1039_o2_p_spl_
  );


  buf

  (
    n2955_lo_p_spl_,
    n2955_lo_p
  );


  buf

  (
    n3027_lo_p_spl_,
    n3027_lo_p
  );


  buf

  (
    n3087_lo_p_spl_,
    n3087_lo_p
  );


  buf

  (
    n3015_lo_p_spl_,
    n3015_lo_p
  );


  buf

  (
    g1078_n_spl_,
    g1078_n
  );


  buf

  (
    g1078_n_spl_0,
    g1078_n_spl_
  );


  buf

  (
    g1078_n_spl_00,
    g1078_n_spl_0
  );


  buf

  (
    g1078_n_spl_1,
    g1078_n_spl_
  );


  buf

  (
    g1222_n_spl_,
    g1222_n
  );


  buf

  (
    g1225_n_spl_,
    g1225_n
  );


  buf

  (
    g1240_n_spl_,
    g1240_n
  );


  buf

  (
    g1249_p_spl_,
    g1249_p
  );


  buf

  (
    g1252_n_spl_,
    g1252_n
  );


  buf

  (
    g1272_p_spl_,
    g1272_p
  );


  buf

  (
    g1292_n_spl_,
    g1292_n
  );


  buf

  (
    g1312_p_spl_,
    g1312_p
  );


  buf

  (
    g1388_p_spl_,
    g1388_p
  );


  buf

  (
    g1388_p_spl_0,
    g1388_p_spl_
  );


  buf

  (
    g1390_p_spl_,
    g1390_p
  );


  buf

  (
    g1390_p_spl_0,
    g1390_p_spl_
  );


  buf

  (
    g1401_n_spl_,
    g1401_n
  );


  buf

  (
    g1401_n_spl_0,
    g1401_n_spl_
  );


  buf

  (
    g1423_n_spl_,
    g1423_n
  );


  buf

  (
    g1423_n_spl_0,
    g1423_n_spl_
  );


  buf

  (
    g1425_n_spl_,
    g1425_n
  );


  buf

  (
    g1425_n_spl_0,
    g1425_n_spl_
  );


  buf

  (
    g1425_n_spl_00,
    g1425_n_spl_0
  );


  buf

  (
    g1425_n_spl_01,
    g1425_n_spl_0
  );


  buf

  (
    g1425_n_spl_1,
    g1425_n_spl_
  );


  buf

  (
    n3231_lo_p_spl_,
    n3231_lo_p
  );


  buf

  (
    n3243_lo_p_spl_,
    n3243_lo_p
  );


  buf

  (
    g1550_n_spl_,
    g1550_n
  );


  buf

  (
    g1550_n_spl_0,
    g1550_n_spl_
  );


  buf

  (
    g1550_n_spl_00,
    g1550_n_spl_0
  );


  buf

  (
    g1550_n_spl_1,
    g1550_n_spl_
  );


endmodule
