// Benchmark "mymod" written by ABC on Wed Nov  1 23:37:39 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41,
    G468, G469, G470, G471, G472, G473, G474, G475, G476, G477, G478, G479,
    G480, G481, G482, G483, G484, G485, G486, G487, G488, G489, G490, G491,
    G492, G493, G494, G495, G496, G497, G498, G499  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41;
  output G468, G469, G470, G471, G472, G473, G474, G475, G476, G477, G478,
    G479, G480, G481, G482, G483, G484, G485, G486, G487, G488, G489, G490,
    G491, G492, G493, G494, G495, G496, G497, G498, G499;
  reg n286_lo, n298_lo, n310_lo, n322_lo, n334_lo, n346_lo, n358_lo,
    n370_lo, n382_lo, n394_lo, n406_lo, n418_lo, n430_lo, n442_lo, n454_lo,
    n466_lo, n478_lo, n490_lo, n502_lo, n514_lo, n526_lo, n538_lo, n550_lo,
    n562_lo, n574_lo, n586_lo, n598_lo, n610_lo, n622_lo, n634_lo, n646_lo,
    n658_lo, n661_lo, n673_lo, n685_lo, n697_lo, n709_lo, n721_lo, n733_lo,
    n745_lo, n757_lo, n1589_o2, n1590_o2, n1591_o2, n1592_o2, n1593_o2,
    n1594_o2, n1595_o2, n1596_o2, n1597_o2, n1598_o2, n1599_o2, n1600_o2,
    n1601_o2, n1602_o2, n1603_o2, n1604_o2, n1605_o2, n1606_o2, n1607_o2,
    n1608_o2, n1609_o2, n1610_o2, n1611_o2, n1612_o2, n1613_o2, n1614_o2,
    n1615_o2, n1616_o2, n1617_o2, n1618_o2, n1619_o2, n1620_o2, n602_o2,
    n639_o2, n678_o2, n658_o2, n783_o2, n802_o2, n726_o2, n763_o2, n685_o2,
    n680_o2, n822_o2, n843_o2, n842_o2, n681_o2, n684_o2, n686_o2, n823_o2,
    lo002_buf_o2, lo006_buf_o2, lo010_buf_o2, lo014_buf_o2, lo018_buf_o2,
    lo022_buf_o2, lo026_buf_o2, lo030_buf_o2, lo034_buf_o2, lo038_buf_o2,
    lo042_buf_o2, lo046_buf_o2, lo050_buf_o2, lo054_buf_o2, lo058_buf_o2,
    lo062_buf_o2, lo066_buf_o2, lo070_buf_o2, lo074_buf_o2, lo078_buf_o2,
    lo082_buf_o2, lo086_buf_o2, lo090_buf_o2, lo094_buf_o2, lo098_buf_o2,
    lo102_buf_o2, lo106_buf_o2, lo110_buf_o2, lo114_buf_o2, lo118_buf_o2,
    lo122_buf_o2, lo126_buf_o2, n683_o2, n688_o2, n803_o2, n862_o2,
    n764_o2, n863_o2, n886_o2, n600_o2, n601_o2, n637_o2, n638_o2, n676_o2,
    n677_o2, n656_o2, n657_o2, n781_o2, n782_o2, n800_o2, n801_o2, n724_o2,
    n725_o2, n761_o2, n762_o2, lo129_buf_o2, lo133_buf_o2, lo137_buf_o2,
    lo141_buf_o2, lo145_buf_o2, lo149_buf_o2, lo153_buf_o2, lo157_buf_o2,
    lo161_buf_o2, n708_o2, n745_o2, n717_o2, n754_o2, n584_o2, n593_o2,
    n630_o2, n621_o2, lo001_buf_o2, lo005_buf_o2, lo009_buf_o2,
    lo013_buf_o2, lo017_buf_o2, lo021_buf_o2, lo025_buf_o2, lo029_buf_o2,
    lo033_buf_o2, lo037_buf_o2, lo041_buf_o2, lo045_buf_o2, lo049_buf_o2,
    lo053_buf_o2, lo057_buf_o2, lo061_buf_o2, lo065_buf_o2, lo069_buf_o2,
    lo073_buf_o2, lo077_buf_o2, lo081_buf_o2, lo085_buf_o2, lo089_buf_o2,
    lo093_buf_o2, lo097_buf_o2, lo101_buf_o2, lo105_buf_o2, lo109_buf_o2,
    lo113_buf_o2, lo117_buf_o2, lo121_buf_o2, lo125_buf_o2;
  wire new_n462_, new_n464_, new_n466_, new_n468_, new_n470_, new_n472_,
    new_n474_, new_n476_, new_n478_, new_n480_, new_n482_, new_n484_,
    new_n486_, new_n488_, new_n490_, new_n492_, new_n494_, new_n496_,
    new_n498_, new_n500_, new_n502_, new_n504_, new_n506_, new_n508_,
    new_n510_, new_n512_, new_n514_, new_n516_, new_n518_, new_n520_,
    new_n522_, new_n524_, new_n526_, new_n528_, new_n530_, new_n532_,
    new_n534_, new_n536_, new_n538_, new_n540_, new_n542_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n612_,
    new_n614_, new_n616_, new_n618_, new_n620_, new_n622_, new_n624_,
    new_n626_, new_n628_, new_n630_, new_n632_, new_n634_, new_n636_,
    new_n638_, new_n640_, new_n642_, new_n644_, new_n646_, new_n648_,
    new_n650_, new_n652_, new_n654_, new_n656_, new_n658_, new_n660_,
    new_n662_, new_n664_, new_n666_, new_n668_, new_n670_, new_n672_,
    new_n674_, new_n676_, new_n678_, new_n680_, new_n682_, new_n684_,
    new_n686_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1738_, new_n1739_, new_n1740_, new_n1741_,
    new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_,
    new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_,
    new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_,
    new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_,
    new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_,
    new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_,
    new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_,
    new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_,
    new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_,
    new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_,
    new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_,
    new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_,
    new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_,
    new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_,
    new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_,
    new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_,
    new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_,
    new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_,
    new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_,
    new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_,
    new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_,
    new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_,
    new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_,
    new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_,
    new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_,
    new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_,
    new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_,
    new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_,
    new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_,
    new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_,
    new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_,
    new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_,
    new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_,
    new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_,
    new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_,
    new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_,
    new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_,
    new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_,
    new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_,
    new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_,
    new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_,
    new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_,
    new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_,
    new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_,
    new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_,
    new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_,
    new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_,
    new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_,
    new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_,
    new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_,
    new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_,
    new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_,
    new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_,
    new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_,
    new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_,
    new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_,
    new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_,
    new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_,
    new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_,
    new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_,
    new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_,
    new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_,
    new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_,
    n1020_li003_li003, n1032_li007_li007, n1044_li011_li011,
    n1056_li015_li015, n1068_li019_li019, n1080_li023_li023,
    n1092_li027_li027, n1104_li031_li031, n1116_li035_li035,
    n1128_li039_li039, n1140_li043_li043, n1152_li047_li047,
    n1164_li051_li051, n1176_li055_li055, n1188_li059_li059,
    n1200_li063_li063, n1212_li067_li067, n1224_li071_li071,
    n1236_li075_li075, n1248_li079_li079, n1260_li083_li083,
    n1272_li087_li087, n1284_li091_li091, n1296_li095_li095,
    n1308_li099_li099, n1320_li103_li103, n1332_li107_li107,
    n1344_li111_li111, n1356_li115_li115, n1368_li119_li119,
    n1380_li123_li123, n1392_li127_li127, n1395_li128_li128,
    n1407_li132_li132, n1419_li136_li136, n1431_li140_li140,
    n1443_li144_li144, n1455_li148_li148, n1467_li152_li152,
    n1479_li156_li156, n1491_li160_li160, n1589_i2, n1590_i2, n1591_i2,
    n1592_i2, n1593_i2, n1594_i2, n1595_i2, n1596_i2, n1597_i2, n1598_i2,
    n1599_i2, n1600_i2, n1601_i2, n1602_i2, n1603_i2, n1604_i2, n1605_i2,
    n1606_i2, n1607_i2, n1608_i2, n1609_i2, n1610_i2, n1611_i2, n1612_i2,
    n1613_i2, n1614_i2, n1615_i2, n1616_i2, n1617_i2, n1618_i2, n1619_i2,
    n1620_i2, n602_i2, n639_i2, n678_i2, n658_i2, n783_i2, n802_i2,
    n726_i2, n763_i2, n685_i2, n680_i2, n822_i2, n843_i2, n842_i2, n681_i2,
    n684_i2, n686_i2, n823_i2, lo002_buf_i2, lo006_buf_i2, lo010_buf_i2,
    lo014_buf_i2, lo018_buf_i2, lo022_buf_i2, lo026_buf_i2, lo030_buf_i2,
    lo034_buf_i2, lo038_buf_i2, lo042_buf_i2, lo046_buf_i2, lo050_buf_i2,
    lo054_buf_i2, lo058_buf_i2, lo062_buf_i2, lo066_buf_i2, lo070_buf_i2,
    lo074_buf_i2, lo078_buf_i2, lo082_buf_i2, lo086_buf_i2, lo090_buf_i2,
    lo094_buf_i2, lo098_buf_i2, lo102_buf_i2, lo106_buf_i2, lo110_buf_i2,
    lo114_buf_i2, lo118_buf_i2, lo122_buf_i2, lo126_buf_i2, n683_i2,
    n688_i2, n803_i2, n862_i2, n764_i2, n863_i2, n886_i2, n600_i2, n601_i2,
    n637_i2, n638_i2, n676_i2, n677_i2, n656_i2, n657_i2, n781_i2, n782_i2,
    n800_i2, n801_i2, n724_i2, n725_i2, n761_i2, n762_i2, lo129_buf_i2,
    lo133_buf_i2, lo137_buf_i2, lo141_buf_i2, lo145_buf_i2, lo149_buf_i2,
    lo153_buf_i2, lo157_buf_i2, lo161_buf_i2, n708_i2, n745_i2, n717_i2,
    n754_i2, n584_i2, n593_i2, n630_i2, n621_i2, lo001_buf_i2,
    lo005_buf_i2, lo009_buf_i2, lo013_buf_i2, lo017_buf_i2, lo021_buf_i2,
    lo025_buf_i2, lo029_buf_i2, lo033_buf_i2, lo037_buf_i2, lo041_buf_i2,
    lo045_buf_i2, lo049_buf_i2, lo053_buf_i2, lo057_buf_i2, lo061_buf_i2,
    lo065_buf_i2, lo069_buf_i2, lo073_buf_i2, lo077_buf_i2, lo081_buf_i2,
    lo085_buf_i2, lo089_buf_i2, lo093_buf_i2, lo097_buf_i2, lo101_buf_i2,
    lo105_buf_i2, lo109_buf_i2, lo113_buf_i2, lo117_buf_i2, lo121_buf_i2,
    lo125_buf_i2;
  assign new_n462_ = G1;
  assign new_n464_ = G2;
  assign new_n466_ = G3;
  assign new_n468_ = G4;
  assign new_n470_ = G5;
  assign new_n472_ = G6;
  assign new_n474_ = G7;
  assign new_n476_ = G8;
  assign new_n478_ = G9;
  assign new_n480_ = G10;
  assign new_n482_ = G11;
  assign new_n484_ = G12;
  assign new_n486_ = G13;
  assign new_n488_ = G14;
  assign new_n490_ = G15;
  assign new_n492_ = G16;
  assign new_n494_ = G17;
  assign new_n496_ = G18;
  assign new_n498_ = G19;
  assign new_n500_ = G20;
  assign new_n502_ = G21;
  assign new_n504_ = G22;
  assign new_n506_ = G23;
  assign new_n508_ = G24;
  assign new_n510_ = G25;
  assign new_n512_ = G26;
  assign new_n514_ = G27;
  assign new_n516_ = G28;
  assign new_n518_ = G29;
  assign new_n520_ = G30;
  assign new_n522_ = G31;
  assign new_n524_ = G32;
  assign new_n526_ = G33;
  assign new_n528_ = G34;
  assign new_n530_ = G35;
  assign new_n532_ = G36;
  assign new_n534_ = G37;
  assign new_n536_ = G38;
  assign new_n538_ = G39;
  assign new_n540_ = G40;
  assign new_n542_ = G41;
  assign new_n544_ = n286_lo;
  assign new_n545_ = ~n286_lo;
  assign new_n546_ = n298_lo;
  assign new_n547_ = ~n298_lo;
  assign new_n548_ = n310_lo;
  assign new_n549_ = ~n310_lo;
  assign new_n550_ = n322_lo;
  assign new_n551_ = ~n322_lo;
  assign new_n552_ = n334_lo;
  assign new_n553_ = ~n334_lo;
  assign new_n554_ = n346_lo;
  assign new_n555_ = ~n346_lo;
  assign new_n556_ = n358_lo;
  assign new_n557_ = ~n358_lo;
  assign new_n558_ = n370_lo;
  assign new_n559_ = ~n370_lo;
  assign new_n560_ = n382_lo;
  assign new_n561_ = ~n382_lo;
  assign new_n562_ = n394_lo;
  assign new_n563_ = ~n394_lo;
  assign new_n564_ = n406_lo;
  assign new_n565_ = ~n406_lo;
  assign new_n566_ = n418_lo;
  assign new_n567_ = ~n418_lo;
  assign new_n568_ = n430_lo;
  assign new_n569_ = ~n430_lo;
  assign new_n570_ = n442_lo;
  assign new_n571_ = ~n442_lo;
  assign new_n572_ = n454_lo;
  assign new_n573_ = ~n454_lo;
  assign new_n574_ = n466_lo;
  assign new_n575_ = ~n466_lo;
  assign new_n576_ = n478_lo;
  assign new_n577_ = ~n478_lo;
  assign new_n578_ = n490_lo;
  assign new_n579_ = ~n490_lo;
  assign new_n580_ = n502_lo;
  assign new_n581_ = ~n502_lo;
  assign new_n582_ = n514_lo;
  assign new_n583_ = ~n514_lo;
  assign new_n584_ = n526_lo;
  assign new_n585_ = ~n526_lo;
  assign new_n586_ = n538_lo;
  assign new_n587_ = ~n538_lo;
  assign new_n588_ = n550_lo;
  assign new_n589_ = ~n550_lo;
  assign new_n590_ = n562_lo;
  assign new_n591_ = ~n562_lo;
  assign new_n592_ = n574_lo;
  assign new_n593_ = ~n574_lo;
  assign new_n594_ = n586_lo;
  assign new_n595_ = ~n586_lo;
  assign new_n596_ = n598_lo;
  assign new_n597_ = ~n598_lo;
  assign new_n598_ = n610_lo;
  assign new_n599_ = ~n610_lo;
  assign new_n600_ = n622_lo;
  assign new_n601_ = ~n622_lo;
  assign new_n602_ = n634_lo;
  assign new_n603_ = ~n634_lo;
  assign new_n604_ = n646_lo;
  assign new_n605_ = ~n646_lo;
  assign new_n606_ = n658_lo;
  assign new_n607_ = ~n658_lo;
  assign new_n608_ = n661_lo;
  assign new_n610_ = n673_lo;
  assign new_n612_ = n685_lo;
  assign new_n614_ = n697_lo;
  assign new_n616_ = n709_lo;
  assign new_n618_ = n721_lo;
  assign new_n620_ = n733_lo;
  assign new_n622_ = n745_lo;
  assign new_n624_ = n757_lo;
  assign new_n626_ = n1589_o2;
  assign new_n628_ = n1590_o2;
  assign new_n630_ = n1591_o2;
  assign new_n632_ = n1592_o2;
  assign new_n634_ = n1593_o2;
  assign new_n636_ = n1594_o2;
  assign new_n638_ = n1595_o2;
  assign new_n640_ = n1596_o2;
  assign new_n642_ = n1597_o2;
  assign new_n644_ = n1598_o2;
  assign new_n646_ = n1599_o2;
  assign new_n648_ = n1600_o2;
  assign new_n650_ = n1601_o2;
  assign new_n652_ = n1602_o2;
  assign new_n654_ = n1603_o2;
  assign new_n656_ = n1604_o2;
  assign new_n658_ = n1605_o2;
  assign new_n660_ = n1606_o2;
  assign new_n662_ = n1607_o2;
  assign new_n664_ = n1608_o2;
  assign new_n666_ = n1609_o2;
  assign new_n668_ = n1610_o2;
  assign new_n670_ = n1611_o2;
  assign new_n672_ = n1612_o2;
  assign new_n674_ = n1613_o2;
  assign new_n676_ = n1614_o2;
  assign new_n678_ = n1615_o2;
  assign new_n680_ = n1616_o2;
  assign new_n682_ = n1617_o2;
  assign new_n684_ = n1618_o2;
  assign new_n686_ = n1619_o2;
  assign new_n688_ = n1620_o2;
  assign new_n690_ = n602_o2;
  assign new_n691_ = ~n602_o2;
  assign new_n692_ = n639_o2;
  assign new_n693_ = ~n639_o2;
  assign new_n694_ = n678_o2;
  assign new_n695_ = ~n678_o2;
  assign new_n696_ = n658_o2;
  assign new_n697_ = ~n658_o2;
  assign new_n698_ = n783_o2;
  assign new_n699_ = ~n783_o2;
  assign new_n700_ = n802_o2;
  assign new_n701_ = ~n802_o2;
  assign new_n702_ = n726_o2;
  assign new_n703_ = ~n726_o2;
  assign new_n704_ = n763_o2;
  assign new_n705_ = ~n763_o2;
  assign new_n706_ = n685_o2;
  assign new_n707_ = ~n685_o2;
  assign new_n708_ = n680_o2;
  assign new_n709_ = ~n680_o2;
  assign new_n710_ = n822_o2;
  assign new_n711_ = ~n822_o2;
  assign new_n712_ = n843_o2;
  assign new_n713_ = ~n843_o2;
  assign new_n714_ = n842_o2;
  assign new_n715_ = ~n842_o2;
  assign new_n716_ = n681_o2;
  assign new_n717_ = ~n681_o2;
  assign new_n718_ = n684_o2;
  assign new_n719_ = ~n684_o2;
  assign new_n720_ = n686_o2;
  assign new_n721_ = ~n686_o2;
  assign new_n722_ = n823_o2;
  assign new_n723_ = ~n823_o2;
  assign new_n724_ = lo002_buf_o2;
  assign new_n725_ = ~lo002_buf_o2;
  assign new_n726_ = lo006_buf_o2;
  assign new_n727_ = ~lo006_buf_o2;
  assign new_n728_ = lo010_buf_o2;
  assign new_n729_ = ~lo010_buf_o2;
  assign new_n730_ = lo014_buf_o2;
  assign new_n731_ = ~lo014_buf_o2;
  assign new_n732_ = lo018_buf_o2;
  assign new_n733_ = ~lo018_buf_o2;
  assign new_n734_ = lo022_buf_o2;
  assign new_n735_ = ~lo022_buf_o2;
  assign new_n736_ = lo026_buf_o2;
  assign new_n737_ = ~lo026_buf_o2;
  assign new_n738_ = lo030_buf_o2;
  assign new_n739_ = ~lo030_buf_o2;
  assign new_n740_ = lo034_buf_o2;
  assign new_n741_ = ~lo034_buf_o2;
  assign new_n742_ = lo038_buf_o2;
  assign new_n743_ = ~lo038_buf_o2;
  assign new_n744_ = lo042_buf_o2;
  assign new_n745_ = ~lo042_buf_o2;
  assign new_n746_ = lo046_buf_o2;
  assign new_n747_ = ~lo046_buf_o2;
  assign new_n748_ = lo050_buf_o2;
  assign new_n749_ = ~lo050_buf_o2;
  assign new_n750_ = lo054_buf_o2;
  assign new_n751_ = ~lo054_buf_o2;
  assign new_n752_ = lo058_buf_o2;
  assign new_n753_ = ~lo058_buf_o2;
  assign new_n754_ = lo062_buf_o2;
  assign new_n755_ = ~lo062_buf_o2;
  assign new_n756_ = lo066_buf_o2;
  assign new_n757_ = ~lo066_buf_o2;
  assign new_n758_ = lo070_buf_o2;
  assign new_n759_ = ~lo070_buf_o2;
  assign new_n760_ = lo074_buf_o2;
  assign new_n761_ = ~lo074_buf_o2;
  assign new_n762_ = lo078_buf_o2;
  assign new_n763_ = ~lo078_buf_o2;
  assign new_n764_ = lo082_buf_o2;
  assign new_n765_ = ~lo082_buf_o2;
  assign new_n766_ = lo086_buf_o2;
  assign new_n767_ = ~lo086_buf_o2;
  assign new_n768_ = lo090_buf_o2;
  assign new_n769_ = ~lo090_buf_o2;
  assign new_n770_ = lo094_buf_o2;
  assign new_n771_ = ~lo094_buf_o2;
  assign new_n772_ = lo098_buf_o2;
  assign new_n773_ = ~lo098_buf_o2;
  assign new_n774_ = lo102_buf_o2;
  assign new_n775_ = ~lo102_buf_o2;
  assign new_n776_ = lo106_buf_o2;
  assign new_n777_ = ~lo106_buf_o2;
  assign new_n778_ = lo110_buf_o2;
  assign new_n779_ = ~lo110_buf_o2;
  assign new_n780_ = lo114_buf_o2;
  assign new_n781_ = ~lo114_buf_o2;
  assign new_n782_ = lo118_buf_o2;
  assign new_n783_ = ~lo118_buf_o2;
  assign new_n784_ = lo122_buf_o2;
  assign new_n785_ = ~lo122_buf_o2;
  assign new_n786_ = lo126_buf_o2;
  assign new_n787_ = ~lo126_buf_o2;
  assign new_n788_ = n683_o2;
  assign new_n789_ = ~n683_o2;
  assign new_n790_ = n688_o2;
  assign new_n791_ = ~n688_o2;
  assign new_n792_ = n803_o2;
  assign new_n793_ = ~n803_o2;
  assign new_n794_ = n862_o2;
  assign new_n795_ = ~n862_o2;
  assign new_n796_ = n764_o2;
  assign new_n797_ = ~n764_o2;
  assign new_n798_ = n863_o2;
  assign new_n799_ = ~n863_o2;
  assign new_n800_ = n886_o2;
  assign new_n801_ = ~n886_o2;
  assign new_n802_ = n600_o2;
  assign new_n803_ = ~n600_o2;
  assign new_n804_ = n601_o2;
  assign new_n805_ = ~n601_o2;
  assign new_n806_ = n637_o2;
  assign new_n807_ = ~n637_o2;
  assign new_n808_ = n638_o2;
  assign new_n809_ = ~n638_o2;
  assign new_n810_ = n676_o2;
  assign new_n811_ = ~n676_o2;
  assign new_n812_ = n677_o2;
  assign new_n813_ = ~n677_o2;
  assign new_n814_ = n656_o2;
  assign new_n815_ = ~n656_o2;
  assign new_n816_ = n657_o2;
  assign new_n817_ = ~n657_o2;
  assign new_n818_ = n781_o2;
  assign new_n819_ = ~n781_o2;
  assign new_n820_ = n782_o2;
  assign new_n821_ = ~n782_o2;
  assign new_n822_ = n800_o2;
  assign new_n823_ = ~n800_o2;
  assign new_n824_ = n801_o2;
  assign new_n825_ = ~n801_o2;
  assign new_n826_ = n724_o2;
  assign new_n827_ = ~n724_o2;
  assign new_n828_ = n725_o2;
  assign new_n829_ = ~n725_o2;
  assign new_n830_ = n761_o2;
  assign new_n831_ = ~n761_o2;
  assign new_n832_ = n762_o2;
  assign new_n833_ = ~n762_o2;
  assign new_n834_ = lo129_buf_o2;
  assign new_n835_ = ~lo129_buf_o2;
  assign new_n836_ = lo133_buf_o2;
  assign new_n837_ = ~lo133_buf_o2;
  assign new_n838_ = lo137_buf_o2;
  assign new_n839_ = ~lo137_buf_o2;
  assign new_n840_ = lo141_buf_o2;
  assign new_n841_ = ~lo141_buf_o2;
  assign new_n842_ = lo145_buf_o2;
  assign new_n843_ = ~lo145_buf_o2;
  assign new_n844_ = lo149_buf_o2;
  assign new_n845_ = ~lo149_buf_o2;
  assign new_n846_ = lo153_buf_o2;
  assign new_n847_ = ~lo153_buf_o2;
  assign new_n848_ = lo157_buf_o2;
  assign new_n849_ = ~lo157_buf_o2;
  assign new_n850_ = lo161_buf_o2;
  assign new_n851_ = ~lo161_buf_o2;
  assign new_n852_ = n708_o2;
  assign new_n853_ = ~n708_o2;
  assign new_n854_ = n745_o2;
  assign new_n855_ = ~n745_o2;
  assign new_n856_ = n717_o2;
  assign new_n857_ = ~n717_o2;
  assign new_n858_ = n754_o2;
  assign new_n859_ = ~n754_o2;
  assign new_n860_ = n584_o2;
  assign new_n861_ = ~n584_o2;
  assign new_n862_ = n593_o2;
  assign new_n863_ = ~n593_o2;
  assign new_n864_ = n630_o2;
  assign new_n865_ = ~n630_o2;
  assign new_n866_ = n621_o2;
  assign new_n867_ = ~n621_o2;
  assign new_n868_ = lo001_buf_o2;
  assign new_n869_ = ~lo001_buf_o2;
  assign new_n870_ = lo005_buf_o2;
  assign new_n871_ = ~lo005_buf_o2;
  assign new_n872_ = lo009_buf_o2;
  assign new_n873_ = ~lo009_buf_o2;
  assign new_n874_ = lo013_buf_o2;
  assign new_n875_ = ~lo013_buf_o2;
  assign new_n876_ = lo017_buf_o2;
  assign new_n877_ = ~lo017_buf_o2;
  assign new_n878_ = lo021_buf_o2;
  assign new_n879_ = ~lo021_buf_o2;
  assign new_n880_ = lo025_buf_o2;
  assign new_n881_ = ~lo025_buf_o2;
  assign new_n882_ = lo029_buf_o2;
  assign new_n883_ = ~lo029_buf_o2;
  assign new_n884_ = lo033_buf_o2;
  assign new_n885_ = ~lo033_buf_o2;
  assign new_n886_ = lo037_buf_o2;
  assign new_n887_ = ~lo037_buf_o2;
  assign new_n888_ = lo041_buf_o2;
  assign new_n889_ = ~lo041_buf_o2;
  assign new_n890_ = lo045_buf_o2;
  assign new_n891_ = ~lo045_buf_o2;
  assign new_n892_ = lo049_buf_o2;
  assign new_n893_ = ~lo049_buf_o2;
  assign new_n894_ = lo053_buf_o2;
  assign new_n895_ = ~lo053_buf_o2;
  assign new_n896_ = lo057_buf_o2;
  assign new_n897_ = ~lo057_buf_o2;
  assign new_n898_ = lo061_buf_o2;
  assign new_n899_ = ~lo061_buf_o2;
  assign new_n900_ = lo065_buf_o2;
  assign new_n901_ = ~lo065_buf_o2;
  assign new_n902_ = lo069_buf_o2;
  assign new_n903_ = ~lo069_buf_o2;
  assign new_n904_ = lo073_buf_o2;
  assign new_n905_ = ~lo073_buf_o2;
  assign new_n906_ = lo077_buf_o2;
  assign new_n907_ = ~lo077_buf_o2;
  assign new_n908_ = lo081_buf_o2;
  assign new_n909_ = ~lo081_buf_o2;
  assign new_n910_ = lo085_buf_o2;
  assign new_n911_ = ~lo085_buf_o2;
  assign new_n912_ = lo089_buf_o2;
  assign new_n913_ = ~lo089_buf_o2;
  assign new_n914_ = lo093_buf_o2;
  assign new_n915_ = ~lo093_buf_o2;
  assign new_n916_ = lo097_buf_o2;
  assign new_n917_ = ~lo097_buf_o2;
  assign new_n918_ = lo101_buf_o2;
  assign new_n919_ = ~lo101_buf_o2;
  assign new_n920_ = lo105_buf_o2;
  assign new_n921_ = ~lo105_buf_o2;
  assign new_n922_ = lo109_buf_o2;
  assign new_n923_ = ~lo109_buf_o2;
  assign new_n924_ = lo113_buf_o2;
  assign new_n925_ = ~lo113_buf_o2;
  assign new_n926_ = lo117_buf_o2;
  assign new_n927_ = ~lo117_buf_o2;
  assign new_n928_ = lo121_buf_o2;
  assign new_n929_ = ~lo121_buf_o2;
  assign new_n930_ = lo125_buf_o2;
  assign new_n931_ = ~lo125_buf_o2;
  assign new_n932_ = new_n789_ & new_n791_;
  assign new_n933_ = new_n788_ | new_n790_;
  assign new_n934_ = new_n792_ & new_n796_;
  assign new_n935_ = new_n793_ | new_n797_;
  assign new_n936_ = new_n1739_ & new_n934_;
  assign new_n937_ = new_n1742_ | new_n935_;
  assign new_n938_ = new_n1745_ & new_n1748_;
  assign new_n939_ = new_n1751_ | new_n1754_;
  assign new_n940_ = new_n545_ & new_n938_;
  assign new_n941_ = new_n544_ & new_n939_;
  assign new_n942_ = new_n940_ | new_n941_;
  assign new_n943_ = new_n1758_ & new_n1748_;
  assign new_n944_ = new_n1762_ | new_n1754_;
  assign new_n945_ = new_n547_ & new_n943_;
  assign new_n946_ = new_n546_ & new_n944_;
  assign new_n947_ = new_n945_ | new_n946_;
  assign new_n948_ = new_n1766_ & new_n1749_;
  assign new_n949_ = new_n1771_ | new_n1755_;
  assign new_n950_ = new_n549_ & new_n948_;
  assign new_n951_ = new_n548_ & new_n949_;
  assign new_n952_ = new_n950_ | new_n951_;
  assign new_n953_ = new_n1775_ & new_n1749_;
  assign new_n954_ = new_n1778_ | new_n1755_;
  assign new_n955_ = new_n551_ & new_n953_;
  assign new_n956_ = new_n550_ & new_n954_;
  assign new_n957_ = new_n955_ | new_n956_;
  assign new_n958_ = new_n710_ & new_n723_;
  assign new_n959_ = new_n711_ | new_n722_;
  assign new_n960_ = new_n1739_ & new_n958_;
  assign new_n961_ = new_n1742_ | new_n959_;
  assign new_n962_ = new_n1745_ & new_n1781_;
  assign new_n963_ = new_n1751_ | new_n1784_;
  assign new_n964_ = new_n553_ & new_n962_;
  assign new_n965_ = new_n552_ & new_n963_;
  assign new_n966_ = new_n964_ | new_n965_;
  assign new_n967_ = new_n1758_ & new_n1781_;
  assign new_n968_ = new_n1762_ | new_n1784_;
  assign new_n969_ = new_n555_ & new_n967_;
  assign new_n970_ = new_n554_ & new_n968_;
  assign new_n971_ = new_n969_ | new_n970_;
  assign new_n972_ = new_n1766_ & new_n1782_;
  assign new_n973_ = new_n1771_ | new_n1785_;
  assign new_n974_ = new_n557_ & new_n972_;
  assign new_n975_ = new_n556_ & new_n973_;
  assign new_n976_ = new_n974_ | new_n975_;
  assign new_n977_ = new_n1775_ & new_n1782_;
  assign new_n978_ = new_n1778_ | new_n1785_;
  assign new_n979_ = new_n559_ & new_n977_;
  assign new_n980_ = new_n558_ & new_n978_;
  assign new_n981_ = new_n979_ | new_n980_;
  assign new_n982_ = new_n713_ & new_n714_;
  assign new_n983_ = new_n712_ | new_n715_;
  assign new_n984_ = new_n1740_ & new_n982_;
  assign new_n985_ = new_n1743_ | new_n983_;
  assign new_n986_ = new_n1746_ & new_n1787_;
  assign new_n987_ = new_n1752_ | new_n1790_;
  assign new_n988_ = new_n561_ & new_n986_;
  assign new_n989_ = new_n560_ & new_n987_;
  assign new_n990_ = new_n988_ | new_n989_;
  assign new_n991_ = new_n1757_ & new_n1787_;
  assign new_n992_ = new_n1761_ | new_n1790_;
  assign new_n993_ = new_n563_ & new_n991_;
  assign new_n994_ = new_n562_ & new_n992_;
  assign new_n995_ = new_n993_ | new_n994_;
  assign new_n996_ = new_n1767_ & new_n1788_;
  assign new_n997_ = new_n1772_ | new_n1791_;
  assign new_n998_ = new_n565_ & new_n996_;
  assign new_n999_ = new_n564_ & new_n997_;
  assign new_n1000_ = new_n998_ | new_n999_;
  assign new_n1001_ = new_n1776_ & new_n1788_;
  assign new_n1002_ = new_n1779_ | new_n1791_;
  assign new_n1003_ = new_n567_ & new_n1001_;
  assign new_n1004_ = new_n566_ & new_n1002_;
  assign new_n1005_ = new_n1003_ | new_n1004_;
  assign new_n1006_ = new_n794_ & new_n798_;
  assign new_n1007_ = new_n795_ | new_n799_;
  assign new_n1008_ = new_n1740_ & new_n1006_;
  assign new_n1009_ = new_n1743_ | new_n1007_;
  assign new_n1010_ = new_n1746_ & new_n1793_;
  assign new_n1011_ = new_n1752_ | new_n1796_;
  assign new_n1012_ = new_n569_ & new_n1010_;
  assign new_n1013_ = new_n568_ & new_n1011_;
  assign new_n1014_ = new_n1012_ | new_n1013_;
  assign new_n1015_ = new_n1759_ & new_n1793_;
  assign new_n1016_ = new_n1763_ | new_n1796_;
  assign new_n1017_ = new_n571_ & new_n1015_;
  assign new_n1018_ = new_n570_ & new_n1016_;
  assign new_n1019_ = new_n1017_ | new_n1018_;
  assign new_n1020_ = new_n1767_ & new_n1794_;
  assign new_n1021_ = new_n1772_ | new_n1797_;
  assign new_n1022_ = new_n573_ & new_n1020_;
  assign new_n1023_ = new_n572_ & new_n1021_;
  assign new_n1024_ = new_n1022_ | new_n1023_;
  assign new_n1025_ = new_n1776_ & new_n1794_;
  assign new_n1026_ = new_n1779_ | new_n1797_;
  assign new_n1027_ = new_n575_ & new_n1025_;
  assign new_n1028_ = new_n574_ & new_n1026_;
  assign new_n1029_ = new_n1027_ | new_n1028_;
  assign new_n1030_ = new_n720_ & new_n1799_;
  assign new_n1031_ = new_n721_ | new_n1802_;
  assign new_n1032_ = new_n1768_ & new_n1030_;
  assign new_n1033_ = new_n1773_ | new_n1031_;
  assign new_n1034_ = new_n1805_ & new_n1808_;
  assign new_n1035_ = new_n1811_ | new_n1814_;
  assign new_n1036_ = new_n577_ & new_n1034_;
  assign new_n1037_ = new_n576_ & new_n1035_;
  assign new_n1038_ = new_n1036_ | new_n1037_;
  assign new_n1039_ = new_n1817_ & new_n1808_;
  assign new_n1040_ = new_n1820_ | new_n1814_;
  assign new_n1041_ = new_n579_ & new_n1039_;
  assign new_n1042_ = new_n578_ & new_n1040_;
  assign new_n1043_ = new_n1041_ | new_n1042_;
  assign new_n1044_ = new_n1823_ & new_n1809_;
  assign new_n1045_ = new_n1826_ | new_n1815_;
  assign new_n1046_ = new_n581_ & new_n1044_;
  assign new_n1047_ = new_n580_ & new_n1045_;
  assign new_n1048_ = new_n1046_ | new_n1047_;
  assign new_n1049_ = new_n1829_ & new_n1809_;
  assign new_n1050_ = new_n1832_ | new_n1815_;
  assign new_n1051_ = new_n583_ & new_n1049_;
  assign new_n1052_ = new_n582_ & new_n1050_;
  assign new_n1053_ = new_n1051_ | new_n1052_;
  assign new_n1054_ = new_n706_ & new_n708_;
  assign new_n1055_ = new_n707_ | new_n709_;
  assign new_n1056_ = new_n1799_ & new_n1054_;
  assign new_n1057_ = new_n1802_ | new_n1055_;
  assign new_n1058_ = new_n1805_ & new_n1835_;
  assign new_n1059_ = new_n1811_ | new_n1838_;
  assign new_n1060_ = new_n585_ & new_n1058_;
  assign new_n1061_ = new_n584_ & new_n1059_;
  assign new_n1062_ = new_n1060_ | new_n1061_;
  assign new_n1063_ = new_n1817_ & new_n1835_;
  assign new_n1064_ = new_n1820_ | new_n1838_;
  assign new_n1065_ = new_n587_ & new_n1063_;
  assign new_n1066_ = new_n586_ & new_n1064_;
  assign new_n1067_ = new_n1065_ | new_n1066_;
  assign new_n1068_ = new_n1823_ & new_n1836_;
  assign new_n1069_ = new_n1826_ | new_n1839_;
  assign new_n1070_ = new_n589_ & new_n1068_;
  assign new_n1071_ = new_n588_ & new_n1069_;
  assign new_n1072_ = new_n1070_ | new_n1071_;
  assign new_n1073_ = new_n1829_ & new_n1836_;
  assign new_n1074_ = new_n1832_ | new_n1839_;
  assign new_n1075_ = new_n591_ & new_n1073_;
  assign new_n1076_ = new_n590_ & new_n1074_;
  assign new_n1077_ = new_n1075_ | new_n1076_;
  assign new_n1078_ = new_n1768_ & new_n718_;
  assign new_n1079_ = new_n1773_ | new_n719_;
  assign new_n1080_ = new_n1800_ & new_n1078_;
  assign new_n1081_ = new_n1803_ | new_n1079_;
  assign new_n1082_ = new_n1806_ & new_n1841_;
  assign new_n1083_ = new_n1812_ | new_n1844_;
  assign new_n1084_ = new_n593_ & new_n1082_;
  assign new_n1085_ = new_n592_ & new_n1083_;
  assign new_n1086_ = new_n1084_ | new_n1085_;
  assign new_n1087_ = new_n1818_ & new_n1841_;
  assign new_n1088_ = new_n1821_ | new_n1844_;
  assign new_n1089_ = new_n595_ & new_n1087_;
  assign new_n1090_ = new_n594_ & new_n1088_;
  assign new_n1091_ = new_n1089_ | new_n1090_;
  assign new_n1092_ = new_n1824_ & new_n1842_;
  assign new_n1093_ = new_n1827_ | new_n1845_;
  assign new_n1094_ = new_n597_ & new_n1092_;
  assign new_n1095_ = new_n596_ & new_n1093_;
  assign new_n1096_ = new_n1094_ | new_n1095_;
  assign new_n1097_ = new_n1830_ & new_n1842_;
  assign new_n1098_ = new_n1833_ | new_n1845_;
  assign new_n1099_ = new_n599_ & new_n1097_;
  assign new_n1100_ = new_n598_ & new_n1098_;
  assign new_n1101_ = new_n1099_ | new_n1100_;
  assign new_n1102_ = new_n1759_ & new_n716_;
  assign new_n1103_ = new_n1763_ | new_n717_;
  assign new_n1104_ = new_n1800_ & new_n1102_;
  assign new_n1105_ = new_n1803_ | new_n1103_;
  assign new_n1106_ = new_n1806_ & new_n1847_;
  assign new_n1107_ = new_n1812_ | new_n1850_;
  assign new_n1108_ = new_n601_ & new_n1106_;
  assign new_n1109_ = new_n600_ & new_n1107_;
  assign new_n1110_ = new_n1108_ | new_n1109_;
  assign new_n1111_ = new_n1818_ & new_n1847_;
  assign new_n1112_ = new_n1821_ | new_n1850_;
  assign new_n1113_ = new_n603_ & new_n1111_;
  assign new_n1114_ = new_n602_ & new_n1112_;
  assign new_n1115_ = new_n1113_ | new_n1114_;
  assign new_n1116_ = new_n1824_ & new_n1848_;
  assign new_n1117_ = new_n1827_ | new_n1851_;
  assign new_n1118_ = new_n605_ & new_n1116_;
  assign new_n1119_ = new_n604_ & new_n1117_;
  assign new_n1120_ = new_n1118_ | new_n1119_;
  assign new_n1121_ = new_n1830_ & new_n1848_;
  assign new_n1122_ = new_n1833_ | new_n1851_;
  assign new_n1123_ = new_n607_ & new_n1121_;
  assign new_n1124_ = new_n606_ & new_n1122_;
  assign new_n1125_ = new_n1123_ | new_n1124_;
  assign new_n1126_ = new_n803_ & new_n805_;
  assign new_n1127_ = new_n802_ | new_n804_;
  assign new_n1128_ = new_n807_ & new_n809_;
  assign new_n1129_ = new_n806_ | new_n808_;
  assign new_n1130_ = new_n811_ & new_n813_;
  assign new_n1131_ = new_n810_ | new_n812_;
  assign new_n1132_ = new_n815_ & new_n817_;
  assign new_n1133_ = new_n814_ | new_n816_;
  assign new_n1134_ = new_n819_ & new_n821_;
  assign new_n1135_ = new_n818_ | new_n820_;
  assign new_n1136_ = new_n823_ & new_n825_;
  assign new_n1137_ = new_n822_ | new_n824_;
  assign new_n1138_ = new_n827_ & new_n829_;
  assign new_n1139_ = new_n826_ | new_n828_;
  assign new_n1140_ = new_n831_ & new_n833_;
  assign new_n1141_ = new_n830_ | new_n832_;
  assign new_n1142_ = new_n1126_ | new_n1853_;
  assign new_n1143_ = new_n1855_ | new_n1132_;
  assign new_n1144_ = new_n1857_ | new_n1859_;
  assign new_n1145_ = new_n1857_ & new_n1859_;
  assign new_n1146_ = new_n1861_ | new_n1863_;
  assign new_n1147_ = new_n1865_ | new_n1867_;
  assign new_n1148_ = new_n1869_ | new_n1870_;
  assign new_n1149_ = new_n1869_ | new_n1872_;
  assign new_n1150_ = new_n1128_ | new_n1873_;
  assign new_n1151_ = new_n1872_ | new_n1874_;
  assign new_n1152_ = new_n1865_ & new_n1867_;
  assign new_n1153_ = new_n1876_ | new_n1878_;
  assign new_n1154_ = new_n1130_ | new_n1873_;
  assign new_n1155_ = new_n1879_ & new_n1154_;
  assign new_n1156_ = new_n1853_ | new_n1155_;
  assign new_n1157_ = new_n1880_ & new_n1881_;
  assign new_n1158_ = new_n1855_ | new_n1157_;
  assign new_n1159_ = new_n1861_ & new_n1864_;
  assign new_n1160_ = new_n1856_ & new_n1876_;
  assign new_n1161_ = new_n1878_ & new_n1858_;
  assign new_n1162_ = new_n1866_ & new_n1863_;
  assign new_n1163_ = new_n1882_ & new_n1883_;
  assign new_n1164_ = new_n1884_ | new_n1163_;
  assign new_n1165_ = new_n1145_ & new_n1885_;
  assign new_n1166_ = new_n1152_ | new_n1165_;
  assign new_n1167_ = new_n1164_ & new_n1166_;
  assign new_n1168_ = new_n1887_ & new_n1888_;
  assign new_n1169_ = new_n1889_ | new_n1891_;
  assign new_n1170_ = new_n1889_ & new_n1891_;
  assign new_n1171_ = new_n1887_ | new_n1888_;
  assign new_n1172_ = new_n1169_ & new_n1171_;
  assign new_n1173_ = new_n1168_ | new_n1170_;
  assign new_n1174_ = new_n1893_ & new_n1894_;
  assign new_n1175_ = new_n1895_ | new_n1897_;
  assign new_n1176_ = new_n1895_ & new_n1897_;
  assign new_n1177_ = new_n1893_ | new_n1894_;
  assign new_n1178_ = new_n1175_ & new_n1177_;
  assign new_n1179_ = new_n1174_ | new_n1176_;
  assign new_n1180_ = new_n1172_ & new_n1179_;
  assign new_n1181_ = new_n1173_ & new_n1178_;
  assign new_n1182_ = new_n1180_ | new_n1181_;
  assign new_n1183_ = new_n834_ & new_n1900_;
  assign new_n1184_ = new_n835_ | new_n1907_;
  assign new_n1185_ = new_n1913_ & new_n1916_;
  assign new_n1186_ = new_n1919_ | new_n1922_;
  assign new_n1187_ = new_n1919_ & new_n1922_;
  assign new_n1188_ = new_n1913_ | new_n1916_;
  assign new_n1189_ = new_n1186_ & new_n1188_;
  assign new_n1190_ = new_n1185_ | new_n1187_;
  assign new_n1191_ = new_n1183_ | new_n1189_;
  assign new_n1192_ = new_n1184_ | new_n1190_;
  assign new_n1193_ = new_n1191_ & new_n1192_;
  assign new_n1194_ = new_n1924_ | new_n1925_;
  assign new_n1195_ = new_n1924_ & new_n1925_;
  assign new_n1196_ = new_n1927_ & new_n1928_;
  assign new_n1197_ = new_n1929_ | new_n1931_;
  assign new_n1198_ = new_n1929_ & new_n1931_;
  assign new_n1199_ = new_n1927_ | new_n1928_;
  assign new_n1200_ = new_n1197_ & new_n1199_;
  assign new_n1201_ = new_n1196_ | new_n1198_;
  assign new_n1202_ = new_n1933_ & new_n1934_;
  assign new_n1203_ = new_n1935_ | new_n1937_;
  assign new_n1204_ = new_n1935_ & new_n1937_;
  assign new_n1205_ = new_n1933_ | new_n1934_;
  assign new_n1206_ = new_n1203_ & new_n1205_;
  assign new_n1207_ = new_n1202_ | new_n1204_;
  assign new_n1208_ = new_n1200_ & new_n1207_;
  assign new_n1209_ = new_n1201_ & new_n1206_;
  assign new_n1210_ = new_n1208_ | new_n1209_;
  assign new_n1211_ = new_n836_ & new_n1900_;
  assign new_n1212_ = new_n837_ | new_n1907_;
  assign new_n1213_ = new_n1939_ & new_n1942_;
  assign new_n1214_ = new_n1945_ | new_n1948_;
  assign new_n1215_ = new_n1945_ & new_n1948_;
  assign new_n1216_ = new_n1939_ | new_n1942_;
  assign new_n1217_ = new_n1214_ & new_n1216_;
  assign new_n1218_ = new_n1213_ | new_n1215_;
  assign new_n1219_ = new_n1211_ | new_n1217_;
  assign new_n1220_ = new_n1212_ | new_n1218_;
  assign new_n1221_ = new_n1219_ & new_n1220_;
  assign new_n1222_ = new_n1950_ | new_n1951_;
  assign new_n1223_ = new_n1950_ & new_n1951_;
  assign new_n1224_ = new_n1953_ & new_n1954_;
  assign new_n1225_ = new_n1955_ | new_n1957_;
  assign new_n1226_ = new_n1955_ & new_n1957_;
  assign new_n1227_ = new_n1953_ | new_n1954_;
  assign new_n1228_ = new_n1225_ & new_n1227_;
  assign new_n1229_ = new_n1224_ | new_n1226_;
  assign new_n1230_ = new_n1959_ & new_n1960_;
  assign new_n1231_ = new_n1961_ | new_n1963_;
  assign new_n1232_ = new_n1961_ & new_n1963_;
  assign new_n1233_ = new_n1959_ | new_n1960_;
  assign new_n1234_ = new_n1231_ & new_n1233_;
  assign new_n1235_ = new_n1230_ | new_n1232_;
  assign new_n1236_ = new_n1228_ & new_n1235_;
  assign new_n1237_ = new_n1229_ & new_n1234_;
  assign new_n1238_ = new_n1236_ | new_n1237_;
  assign new_n1239_ = new_n838_ & new_n1901_;
  assign new_n1240_ = new_n839_ | new_n1908_;
  assign new_n1241_ = new_n1914_ & new_n1940_;
  assign new_n1242_ = new_n1920_ | new_n1946_;
  assign new_n1243_ = new_n1920_ & new_n1946_;
  assign new_n1244_ = new_n1914_ | new_n1940_;
  assign new_n1245_ = new_n1242_ & new_n1244_;
  assign new_n1246_ = new_n1241_ | new_n1243_;
  assign new_n1247_ = new_n1239_ | new_n1245_;
  assign new_n1248_ = new_n1240_ | new_n1246_;
  assign new_n1249_ = new_n1247_ & new_n1248_;
  assign new_n1250_ = new_n1964_ | new_n1965_;
  assign new_n1251_ = new_n1964_ & new_n1965_;
  assign new_n1252_ = new_n1967_ & new_n1968_;
  assign new_n1253_ = new_n1969_ | new_n1971_;
  assign new_n1254_ = new_n1969_ & new_n1971_;
  assign new_n1255_ = new_n1967_ | new_n1968_;
  assign new_n1256_ = new_n1253_ & new_n1255_;
  assign new_n1257_ = new_n1252_ | new_n1254_;
  assign new_n1258_ = new_n1973_ & new_n1974_;
  assign new_n1259_ = new_n1975_ | new_n1977_;
  assign new_n1260_ = new_n1975_ & new_n1977_;
  assign new_n1261_ = new_n1973_ | new_n1974_;
  assign new_n1262_ = new_n1259_ & new_n1261_;
  assign new_n1263_ = new_n1258_ | new_n1260_;
  assign new_n1264_ = new_n1256_ & new_n1263_;
  assign new_n1265_ = new_n1257_ & new_n1262_;
  assign new_n1266_ = new_n1264_ | new_n1265_;
  assign new_n1267_ = new_n840_ & new_n1901_;
  assign new_n1268_ = new_n841_ | new_n1908_;
  assign new_n1269_ = new_n1923_ & new_n1949_;
  assign new_n1270_ = new_n1917_ | new_n1943_;
  assign new_n1271_ = new_n1917_ & new_n1943_;
  assign new_n1272_ = new_n1923_ | new_n1949_;
  assign new_n1273_ = new_n1270_ & new_n1272_;
  assign new_n1274_ = new_n1269_ | new_n1271_;
  assign new_n1275_ = new_n1267_ | new_n1273_;
  assign new_n1276_ = new_n1268_ | new_n1274_;
  assign new_n1277_ = new_n1275_ & new_n1276_;
  assign new_n1278_ = new_n1978_ | new_n1979_;
  assign new_n1279_ = new_n1978_ & new_n1979_;
  assign new_n1280_ = new_n1981_ & new_n1982_;
  assign new_n1281_ = new_n1983_ | new_n1985_;
  assign new_n1282_ = new_n1983_ & new_n1985_;
  assign new_n1283_ = new_n1981_ | new_n1982_;
  assign new_n1284_ = new_n1281_ & new_n1283_;
  assign new_n1285_ = new_n1280_ | new_n1282_;
  assign new_n1286_ = new_n1987_ & new_n1988_;
  assign new_n1287_ = new_n1989_ | new_n1991_;
  assign new_n1288_ = new_n1989_ & new_n1991_;
  assign new_n1289_ = new_n1987_ | new_n1988_;
  assign new_n1290_ = new_n1287_ & new_n1289_;
  assign new_n1291_ = new_n1286_ | new_n1288_;
  assign new_n1292_ = new_n1284_ & new_n1291_;
  assign new_n1293_ = new_n1285_ & new_n1290_;
  assign new_n1294_ = new_n1292_ | new_n1293_;
  assign new_n1295_ = new_n842_ & new_n1903_;
  assign new_n1296_ = new_n843_ | new_n1910_;
  assign new_n1297_ = new_n1993_ & new_n1996_;
  assign new_n1298_ = new_n1999_ | new_n2002_;
  assign new_n1299_ = new_n1999_ & new_n2002_;
  assign new_n1300_ = new_n1993_ | new_n1996_;
  assign new_n1301_ = new_n1298_ & new_n1300_;
  assign new_n1302_ = new_n1297_ | new_n1299_;
  assign new_n1303_ = new_n1295_ | new_n1301_;
  assign new_n1304_ = new_n1296_ | new_n1302_;
  assign new_n1305_ = new_n1303_ & new_n1304_;
  assign new_n1306_ = new_n2004_ | new_n2005_;
  assign new_n1307_ = new_n2004_ & new_n2005_;
  assign new_n1308_ = new_n2007_ & new_n2008_;
  assign new_n1309_ = new_n2009_ | new_n2011_;
  assign new_n1310_ = new_n2009_ & new_n2011_;
  assign new_n1311_ = new_n2007_ | new_n2008_;
  assign new_n1312_ = new_n1309_ & new_n1311_;
  assign new_n1313_ = new_n1308_ | new_n1310_;
  assign new_n1314_ = new_n2013_ & new_n2014_;
  assign new_n1315_ = new_n2015_ | new_n2017_;
  assign new_n1316_ = new_n2015_ & new_n2017_;
  assign new_n1317_ = new_n2013_ | new_n2014_;
  assign new_n1318_ = new_n1315_ & new_n1317_;
  assign new_n1319_ = new_n1314_ | new_n1316_;
  assign new_n1320_ = new_n1312_ & new_n1319_;
  assign new_n1321_ = new_n1313_ & new_n1318_;
  assign new_n1322_ = new_n1320_ | new_n1321_;
  assign new_n1323_ = new_n844_ & new_n1903_;
  assign new_n1324_ = new_n845_ | new_n1910_;
  assign new_n1325_ = new_n2019_ & new_n2022_;
  assign new_n1326_ = new_n2025_ | new_n2028_;
  assign new_n1327_ = new_n2025_ & new_n2028_;
  assign new_n1328_ = new_n2019_ | new_n2022_;
  assign new_n1329_ = new_n1326_ & new_n1328_;
  assign new_n1330_ = new_n1325_ | new_n1327_;
  assign new_n1331_ = new_n1323_ | new_n1329_;
  assign new_n1332_ = new_n1324_ | new_n1330_;
  assign new_n1333_ = new_n1331_ & new_n1332_;
  assign new_n1334_ = new_n2030_ | new_n2031_;
  assign new_n1335_ = new_n2030_ & new_n2031_;
  assign new_n1336_ = new_n2033_ & new_n2034_;
  assign new_n1337_ = new_n2035_ | new_n2037_;
  assign new_n1338_ = new_n2035_ & new_n2037_;
  assign new_n1339_ = new_n2033_ | new_n2034_;
  assign new_n1340_ = new_n1337_ & new_n1339_;
  assign new_n1341_ = new_n1336_ | new_n1338_;
  assign new_n1342_ = new_n2039_ & new_n2040_;
  assign new_n1343_ = new_n2041_ | new_n2043_;
  assign new_n1344_ = new_n2041_ & new_n2043_;
  assign new_n1345_ = new_n2039_ | new_n2040_;
  assign new_n1346_ = new_n1343_ & new_n1345_;
  assign new_n1347_ = new_n1342_ | new_n1344_;
  assign new_n1348_ = new_n1340_ & new_n1347_;
  assign new_n1349_ = new_n1341_ & new_n1346_;
  assign new_n1350_ = new_n1348_ | new_n1349_;
  assign new_n1351_ = new_n846_ & new_n1904_;
  assign new_n1352_ = new_n847_ | new_n1911_;
  assign new_n1353_ = new_n1994_ & new_n2026_;
  assign new_n1354_ = new_n2000_ | new_n2020_;
  assign new_n1355_ = new_n2000_ & new_n2020_;
  assign new_n1356_ = new_n1994_ | new_n2026_;
  assign new_n1357_ = new_n1354_ & new_n1356_;
  assign new_n1358_ = new_n1353_ | new_n1355_;
  assign new_n1359_ = new_n1351_ | new_n1357_;
  assign new_n1360_ = new_n1352_ | new_n1358_;
  assign new_n1361_ = new_n1359_ & new_n1360_;
  assign new_n1362_ = new_n2044_ | new_n2045_;
  assign new_n1363_ = new_n2044_ & new_n2045_;
  assign new_n1364_ = new_n2047_ & new_n2048_;
  assign new_n1365_ = new_n2049_ | new_n2051_;
  assign new_n1366_ = new_n2049_ & new_n2051_;
  assign new_n1367_ = new_n2047_ | new_n2048_;
  assign new_n1368_ = new_n1365_ & new_n1367_;
  assign new_n1369_ = new_n1364_ | new_n1366_;
  assign new_n1370_ = new_n2053_ & new_n2054_;
  assign new_n1371_ = new_n2055_ | new_n2057_;
  assign new_n1372_ = new_n2055_ & new_n2057_;
  assign new_n1373_ = new_n2053_ | new_n2054_;
  assign new_n1374_ = new_n1371_ & new_n1373_;
  assign new_n1375_ = new_n1370_ | new_n1372_;
  assign new_n1376_ = new_n1368_ & new_n1375_;
  assign new_n1377_ = new_n1369_ & new_n1374_;
  assign new_n1378_ = new_n1376_ | new_n1377_;
  assign new_n1379_ = new_n848_ & new_n1904_;
  assign new_n1380_ = new_n849_ | new_n1911_;
  assign new_n1381_ = new_n2003_ & new_n2023_;
  assign new_n1382_ = new_n1997_ | new_n2029_;
  assign new_n1383_ = new_n1997_ & new_n2029_;
  assign new_n1384_ = new_n2003_ | new_n2023_;
  assign new_n1385_ = new_n1382_ & new_n1384_;
  assign new_n1386_ = new_n1381_ | new_n1383_;
  assign new_n1387_ = new_n1379_ | new_n1385_;
  assign new_n1388_ = new_n1380_ | new_n1386_;
  assign new_n1389_ = new_n1387_ & new_n1388_;
  assign new_n1390_ = new_n2058_ | new_n2059_;
  assign new_n1391_ = new_n2058_ & new_n2059_;
  assign new_n1392_ = new_n2061_ & new_n2062_;
  assign new_n1393_ = new_n2063_ | new_n2065_;
  assign new_n1394_ = new_n2063_ & new_n2065_;
  assign new_n1395_ = new_n2061_ | new_n2062_;
  assign new_n1396_ = new_n1393_ & new_n1395_;
  assign new_n1397_ = new_n1392_ | new_n1394_;
  assign new_n1398_ = new_n2067_ & new_n2068_;
  assign new_n1399_ = new_n2069_ | new_n2071_;
  assign new_n1400_ = new_n2069_ & new_n2071_;
  assign new_n1401_ = new_n2067_ | new_n2068_;
  assign new_n1402_ = new_n1399_ & new_n1401_;
  assign new_n1403_ = new_n1398_ | new_n1400_;
  assign new_n1404_ = new_n1396_ & new_n1403_;
  assign new_n1405_ = new_n1397_ & new_n1402_;
  assign new_n1406_ = new_n1404_ | new_n1405_;
  assign new_n1407_ = new_n2073_ & new_n2074_;
  assign new_n1408_ = new_n2075_ | new_n2077_;
  assign new_n1409_ = new_n2075_ & new_n2077_;
  assign new_n1410_ = new_n2073_ | new_n2074_;
  assign new_n1411_ = new_n1408_ & new_n1410_;
  assign new_n1412_ = new_n1407_ | new_n1409_;
  assign new_n1413_ = new_n2079_ & new_n2080_;
  assign new_n1414_ = new_n2081_ | new_n2083_;
  assign new_n1415_ = new_n2081_ & new_n2083_;
  assign new_n1416_ = new_n2079_ | new_n2080_;
  assign new_n1417_ = new_n1414_ & new_n1416_;
  assign new_n1418_ = new_n1413_ | new_n1415_;
  assign new_n1419_ = new_n1411_ & new_n1418_;
  assign new_n1420_ = new_n1412_ & new_n1417_;
  assign new_n1421_ = new_n1419_ | new_n1420_;
  assign new_n1422_ = new_n2085_ & new_n2086_;
  assign new_n1423_ = new_n2087_ | new_n2089_;
  assign new_n1424_ = new_n2087_ & new_n2089_;
  assign new_n1425_ = new_n2085_ | new_n2086_;
  assign new_n1426_ = new_n1423_ & new_n1425_;
  assign new_n1427_ = new_n1422_ | new_n1424_;
  assign new_n1428_ = new_n2091_ & new_n2092_;
  assign new_n1429_ = new_n2093_ | new_n2095_;
  assign new_n1430_ = new_n2093_ & new_n2095_;
  assign new_n1431_ = new_n2091_ | new_n2092_;
  assign new_n1432_ = new_n1429_ & new_n1431_;
  assign new_n1433_ = new_n1428_ | new_n1430_;
  assign new_n1434_ = new_n1426_ & new_n1433_;
  assign new_n1435_ = new_n1427_ & new_n1432_;
  assign new_n1436_ = new_n1434_ | new_n1435_;
  assign new_n1437_ = new_n2097_ & new_n2098_;
  assign new_n1438_ = new_n2099_ | new_n2101_;
  assign new_n1439_ = new_n2099_ & new_n2101_;
  assign new_n1440_ = new_n2097_ | new_n2098_;
  assign new_n1441_ = new_n1438_ & new_n1440_;
  assign new_n1442_ = new_n1437_ | new_n1439_;
  assign new_n1443_ = new_n2103_ & new_n2104_;
  assign new_n1444_ = new_n2105_ | new_n2107_;
  assign new_n1445_ = new_n2105_ & new_n2107_;
  assign new_n1446_ = new_n2103_ | new_n2104_;
  assign new_n1447_ = new_n1444_ & new_n1446_;
  assign new_n1448_ = new_n1443_ | new_n1445_;
  assign new_n1449_ = new_n1441_ & new_n1448_;
  assign new_n1450_ = new_n1442_ & new_n1447_;
  assign new_n1451_ = new_n1449_ | new_n1450_;
  assign new_n1452_ = new_n2109_ & new_n2110_;
  assign new_n1453_ = new_n2111_ | new_n2113_;
  assign new_n1454_ = new_n2111_ & new_n2113_;
  assign new_n1455_ = new_n2109_ | new_n2110_;
  assign new_n1456_ = new_n1453_ & new_n1455_;
  assign new_n1457_ = new_n1452_ | new_n1454_;
  assign new_n1458_ = new_n2115_ & new_n2116_;
  assign new_n1459_ = new_n2117_ | new_n2119_;
  assign new_n1460_ = new_n2117_ & new_n2119_;
  assign new_n1461_ = new_n2115_ | new_n2116_;
  assign new_n1462_ = new_n1459_ & new_n1461_;
  assign new_n1463_ = new_n1458_ | new_n1460_;
  assign new_n1464_ = new_n1456_ & new_n1463_;
  assign new_n1465_ = new_n1457_ & new_n1462_;
  assign new_n1466_ = new_n1464_ | new_n1465_;
  assign new_n1467_ = new_n2121_ & new_n2122_;
  assign new_n1468_ = new_n2123_ | new_n2125_;
  assign new_n1469_ = new_n2123_ & new_n2125_;
  assign new_n1470_ = new_n2121_ | new_n2122_;
  assign new_n1471_ = new_n1468_ & new_n1470_;
  assign new_n1472_ = new_n1467_ | new_n1469_;
  assign new_n1473_ = new_n2127_ & new_n2128_;
  assign new_n1474_ = new_n2129_ | new_n2131_;
  assign new_n1475_ = new_n2129_ & new_n2131_;
  assign new_n1476_ = new_n2127_ | new_n2128_;
  assign new_n1477_ = new_n1474_ & new_n1476_;
  assign new_n1478_ = new_n1473_ | new_n1475_;
  assign new_n1479_ = new_n1471_ & new_n1478_;
  assign new_n1480_ = new_n1472_ & new_n1477_;
  assign new_n1481_ = new_n1479_ | new_n1480_;
  assign new_n1482_ = new_n2133_ & new_n2134_;
  assign new_n1483_ = new_n2135_ | new_n2137_;
  assign new_n1484_ = new_n2135_ & new_n2137_;
  assign new_n1485_ = new_n2133_ | new_n2134_;
  assign new_n1486_ = new_n1483_ & new_n1485_;
  assign new_n1487_ = new_n1482_ | new_n1484_;
  assign new_n1488_ = new_n2139_ & new_n2140_;
  assign new_n1489_ = new_n2141_ | new_n2143_;
  assign new_n1490_ = new_n2141_ & new_n2143_;
  assign new_n1491_ = new_n2139_ | new_n2140_;
  assign new_n1492_ = new_n1489_ & new_n1491_;
  assign new_n1493_ = new_n1488_ | new_n1490_;
  assign new_n1494_ = new_n1486_ & new_n1493_;
  assign new_n1495_ = new_n1487_ & new_n1492_;
  assign new_n1496_ = new_n1494_ | new_n1495_;
  assign new_n1497_ = new_n2145_ & new_n2146_;
  assign new_n1498_ = new_n2147_ | new_n2149_;
  assign new_n1499_ = new_n2147_ & new_n2149_;
  assign new_n1500_ = new_n2145_ | new_n2146_;
  assign new_n1501_ = new_n1498_ & new_n1500_;
  assign new_n1502_ = new_n1497_ | new_n1499_;
  assign new_n1503_ = new_n2151_ & new_n2152_;
  assign new_n1504_ = new_n2153_ | new_n2155_;
  assign new_n1505_ = new_n2153_ & new_n2155_;
  assign new_n1506_ = new_n2151_ | new_n2152_;
  assign new_n1507_ = new_n1504_ & new_n1506_;
  assign new_n1508_ = new_n1503_ | new_n1505_;
  assign new_n1509_ = new_n1501_ & new_n1508_;
  assign new_n1510_ = new_n1502_ & new_n1507_;
  assign new_n1511_ = new_n1509_ | new_n1510_;
  assign G468 = new_n942_;
  assign G469 = new_n947_;
  assign G470 = new_n952_;
  assign G471 = new_n957_;
  assign G472 = new_n966_;
  assign G473 = new_n971_;
  assign G474 = new_n976_;
  assign G475 = new_n981_;
  assign G476 = new_n990_;
  assign G477 = new_n995_;
  assign G478 = new_n1000_;
  assign G479 = new_n1005_;
  assign G480 = new_n1014_;
  assign G481 = new_n1019_;
  assign G482 = new_n1024_;
  assign G483 = new_n1029_;
  assign G484 = new_n1038_;
  assign G485 = new_n1043_;
  assign G486 = new_n1048_;
  assign G487 = new_n1053_;
  assign G488 = new_n1062_;
  assign G489 = new_n1067_;
  assign G490 = new_n1072_;
  assign G491 = new_n1077_;
  assign G492 = new_n1086_;
  assign G493 = new_n1091_;
  assign G494 = new_n1096_;
  assign G495 = new_n1101_;
  assign G496 = new_n1110_;
  assign G497 = new_n1115_;
  assign G498 = new_n1120_;
  assign G499 = new_n1125_;
  assign n1020_li003_li003 = new_n626_;
  assign n1032_li007_li007 = new_n628_;
  assign n1044_li011_li011 = new_n630_;
  assign n1056_li015_li015 = new_n632_;
  assign n1068_li019_li019 = new_n634_;
  assign n1080_li023_li023 = new_n636_;
  assign n1092_li027_li027 = new_n638_;
  assign n1104_li031_li031 = new_n640_;
  assign n1116_li035_li035 = new_n642_;
  assign n1128_li039_li039 = new_n644_;
  assign n1140_li043_li043 = new_n646_;
  assign n1152_li047_li047 = new_n648_;
  assign n1164_li051_li051 = new_n650_;
  assign n1176_li055_li055 = new_n652_;
  assign n1188_li059_li059 = new_n654_;
  assign n1200_li063_li063 = new_n656_;
  assign n1212_li067_li067 = new_n658_;
  assign n1224_li071_li071 = new_n660_;
  assign n1236_li075_li075 = new_n662_;
  assign n1248_li079_li079 = new_n664_;
  assign n1260_li083_li083 = new_n666_;
  assign n1272_li087_li087 = new_n668_;
  assign n1284_li091_li091 = new_n670_;
  assign n1296_li095_li095 = new_n672_;
  assign n1308_li099_li099 = new_n674_;
  assign n1320_li103_li103 = new_n676_;
  assign n1332_li107_li107 = new_n678_;
  assign n1344_li111_li111 = new_n680_;
  assign n1356_li115_li115 = new_n682_;
  assign n1368_li119_li119 = new_n684_;
  assign n1380_li123_li123 = new_n686_;
  assign n1392_li127_li127 = new_n688_;
  assign n1395_li128_li128 = new_n526_;
  assign n1407_li132_li132 = new_n528_;
  assign n1419_li136_li136 = new_n530_;
  assign n1431_li140_li140 = new_n532_;
  assign n1443_li144_li144 = new_n534_;
  assign n1455_li148_li148 = new_n536_;
  assign n1467_li152_li152 = new_n538_;
  assign n1479_li156_li156 = new_n540_;
  assign n1491_li160_li160 = new_n542_;
  assign n1589_i2 = new_n1886_;
  assign n1590_i2 = new_n1926_;
  assign n1591_i2 = new_n1952_;
  assign n1592_i2 = new_n1966_;
  assign n1593_i2 = new_n1890_;
  assign n1594_i2 = new_n1930_;
  assign n1595_i2 = new_n1956_;
  assign n1596_i2 = new_n1970_;
  assign n1597_i2 = new_n1892_;
  assign n1598_i2 = new_n1932_;
  assign n1599_i2 = new_n1958_;
  assign n1600_i2 = new_n1972_;
  assign n1601_i2 = new_n1896_;
  assign n1602_i2 = new_n1936_;
  assign n1603_i2 = new_n1962_;
  assign n1604_i2 = new_n1976_;
  assign n1605_i2 = new_n1980_;
  assign n1606_i2 = new_n2006_;
  assign n1607_i2 = new_n2032_;
  assign n1608_i2 = new_n2046_;
  assign n1609_i2 = new_n1984_;
  assign n1610_i2 = new_n2010_;
  assign n1611_i2 = new_n2036_;
  assign n1612_i2 = new_n2050_;
  assign n1613_i2 = new_n1986_;
  assign n1614_i2 = new_n2012_;
  assign n1615_i2 = new_n2038_;
  assign n1616_i2 = new_n2052_;
  assign n1617_i2 = new_n1990_;
  assign n1618_i2 = new_n2016_;
  assign n1619_i2 = new_n2042_;
  assign n1620_i2 = new_n2056_;
  assign n602_i2 = new_n1868_;
  assign n639_i2 = new_n1852_;
  assign n678_i2 = new_n1854_;
  assign n658_i2 = new_n1871_;
  assign n783_i2 = new_n1860_;
  assign n802_i2 = new_n1875_;
  assign n726_i2 = new_n1877_;
  assign n763_i2 = new_n1862_;
  assign n685_i2 = ~new_n1874_;
  assign n680_i2 = ~new_n1870_;
  assign n822_i2 = ~new_n1882_;
  assign n843_i2 = new_n1883_;
  assign n842_i2 = ~new_n1885_;
  assign n681_i2 = ~new_n1879_;
  assign n684_i2 = ~new_n1880_;
  assign n686_i2 = ~new_n1881_;
  assign n823_i2 = new_n1884_;
  assign lo002_buf_i2 = new_n2060_;
  assign lo006_buf_i2 = new_n2064_;
  assign lo010_buf_i2 = new_n2066_;
  assign lo014_buf_i2 = new_n2070_;
  assign lo018_buf_i2 = new_n2072_;
  assign lo022_buf_i2 = new_n2076_;
  assign lo026_buf_i2 = new_n2078_;
  assign lo030_buf_i2 = new_n2082_;
  assign lo034_buf_i2 = new_n2084_;
  assign lo038_buf_i2 = new_n2088_;
  assign lo042_buf_i2 = new_n2090_;
  assign lo046_buf_i2 = new_n2094_;
  assign lo050_buf_i2 = new_n2096_;
  assign lo054_buf_i2 = new_n2100_;
  assign lo058_buf_i2 = new_n2102_;
  assign lo062_buf_i2 = new_n2106_;
  assign lo066_buf_i2 = new_n2108_;
  assign lo070_buf_i2 = new_n2112_;
  assign lo074_buf_i2 = new_n2114_;
  assign lo078_buf_i2 = new_n2118_;
  assign lo082_buf_i2 = new_n2120_;
  assign lo086_buf_i2 = new_n2124_;
  assign lo090_buf_i2 = new_n2126_;
  assign lo094_buf_i2 = new_n2130_;
  assign lo098_buf_i2 = new_n2132_;
  assign lo102_buf_i2 = new_n2136_;
  assign lo106_buf_i2 = new_n2138_;
  assign lo110_buf_i2 = new_n2142_;
  assign lo114_buf_i2 = new_n2144_;
  assign lo118_buf_i2 = new_n2148_;
  assign lo122_buf_i2 = new_n2150_;
  assign lo126_buf_i2 = new_n2154_;
  assign n683_i2 = ~new_n1156_;
  assign n688_i2 = ~new_n1158_;
  assign n803_i2 = new_n1159_;
  assign n862_i2 = new_n1160_;
  assign n764_i2 = new_n1161_;
  assign n863_i2 = new_n1162_;
  assign n886_i2 = new_n1167_;
  assign n600_i2 = ~new_n1194_;
  assign n601_i2 = new_n1195_;
  assign n637_i2 = ~new_n1222_;
  assign n638_i2 = new_n1223_;
  assign n676_i2 = ~new_n1250_;
  assign n677_i2 = new_n1251_;
  assign n656_i2 = ~new_n1278_;
  assign n657_i2 = new_n1279_;
  assign n781_i2 = ~new_n1306_;
  assign n782_i2 = new_n1307_;
  assign n800_i2 = ~new_n1334_;
  assign n801_i2 = new_n1335_;
  assign n724_i2 = ~new_n1362_;
  assign n725_i2 = new_n1363_;
  assign n761_i2 = ~new_n1390_;
  assign n762_i2 = new_n1391_;
  assign lo129_buf_i2 = new_n608_;
  assign lo133_buf_i2 = new_n610_;
  assign lo137_buf_i2 = new_n612_;
  assign lo141_buf_i2 = new_n614_;
  assign lo145_buf_i2 = new_n616_;
  assign lo149_buf_i2 = new_n618_;
  assign lo153_buf_i2 = new_n620_;
  assign lo157_buf_i2 = new_n622_;
  assign lo161_buf_i2 = new_n624_;
  assign n708_i2 = new_n1406_;
  assign n745_i2 = new_n1421_;
  assign n717_i2 = new_n1436_;
  assign n754_i2 = new_n1451_;
  assign n584_i2 = new_n1466_;
  assign n593_i2 = new_n1481_;
  assign n630_i2 = new_n1496_;
  assign n621_i2 = new_n1511_;
  assign lo001_buf_i2 = new_n462_;
  assign lo005_buf_i2 = new_n464_;
  assign lo009_buf_i2 = new_n466_;
  assign lo013_buf_i2 = new_n468_;
  assign lo017_buf_i2 = new_n470_;
  assign lo021_buf_i2 = new_n472_;
  assign lo025_buf_i2 = new_n474_;
  assign lo029_buf_i2 = new_n476_;
  assign lo033_buf_i2 = new_n478_;
  assign lo037_buf_i2 = new_n480_;
  assign lo041_buf_i2 = new_n482_;
  assign lo045_buf_i2 = new_n484_;
  assign lo049_buf_i2 = new_n486_;
  assign lo053_buf_i2 = new_n488_;
  assign lo057_buf_i2 = new_n490_;
  assign lo061_buf_i2 = new_n492_;
  assign lo065_buf_i2 = new_n494_;
  assign lo069_buf_i2 = new_n496_;
  assign lo073_buf_i2 = new_n498_;
  assign lo077_buf_i2 = new_n500_;
  assign lo081_buf_i2 = new_n502_;
  assign lo085_buf_i2 = new_n504_;
  assign lo089_buf_i2 = new_n506_;
  assign lo093_buf_i2 = new_n508_;
  assign lo097_buf_i2 = new_n510_;
  assign lo101_buf_i2 = new_n512_;
  assign lo105_buf_i2 = new_n514_;
  assign lo109_buf_i2 = new_n516_;
  assign lo113_buf_i2 = new_n518_;
  assign lo117_buf_i2 = new_n520_;
  assign lo121_buf_i2 = new_n522_;
  assign lo125_buf_i2 = new_n524_;
  assign new_n1738_ = new_n933_;
  assign new_n1739_ = new_n1738_;
  assign new_n1740_ = new_n1738_;
  assign new_n1741_ = new_n932_;
  assign new_n1742_ = new_n1741_;
  assign new_n1743_ = new_n1741_;
  assign new_n1744_ = new_n690_;
  assign new_n1745_ = new_n1744_;
  assign new_n1746_ = new_n1744_;
  assign new_n1747_ = new_n936_;
  assign new_n1748_ = new_n1747_;
  assign new_n1749_ = new_n1747_;
  assign new_n1750_ = new_n691_;
  assign new_n1751_ = new_n1750_;
  assign new_n1752_ = new_n1750_;
  assign new_n1753_ = new_n937_;
  assign new_n1754_ = new_n1753_;
  assign new_n1755_ = new_n1753_;
  assign new_n1756_ = new_n692_;
  assign new_n1757_ = new_n1756_;
  assign new_n1758_ = new_n1757_;
  assign new_n1759_ = new_n1756_;
  assign new_n1760_ = new_n693_;
  assign new_n1761_ = new_n1760_;
  assign new_n1762_ = new_n1761_;
  assign new_n1763_ = new_n1760_;
  assign new_n1764_ = new_n694_;
  assign new_n1765_ = new_n1764_;
  assign new_n1766_ = new_n1765_;
  assign new_n1767_ = new_n1765_;
  assign new_n1768_ = new_n1764_;
  assign new_n1769_ = new_n695_;
  assign new_n1770_ = new_n1769_;
  assign new_n1771_ = new_n1770_;
  assign new_n1772_ = new_n1770_;
  assign new_n1773_ = new_n1769_;
  assign new_n1774_ = new_n696_;
  assign new_n1775_ = new_n1774_;
  assign new_n1776_ = new_n1774_;
  assign new_n1777_ = new_n697_;
  assign new_n1778_ = new_n1777_;
  assign new_n1779_ = new_n1777_;
  assign new_n1780_ = new_n960_;
  assign new_n1781_ = new_n1780_;
  assign new_n1782_ = new_n1780_;
  assign new_n1783_ = new_n961_;
  assign new_n1784_ = new_n1783_;
  assign new_n1785_ = new_n1783_;
  assign new_n1786_ = new_n984_;
  assign new_n1787_ = new_n1786_;
  assign new_n1788_ = new_n1786_;
  assign new_n1789_ = new_n985_;
  assign new_n1790_ = new_n1789_;
  assign new_n1791_ = new_n1789_;
  assign new_n1792_ = new_n1008_;
  assign new_n1793_ = new_n1792_;
  assign new_n1794_ = new_n1792_;
  assign new_n1795_ = new_n1009_;
  assign new_n1796_ = new_n1795_;
  assign new_n1797_ = new_n1795_;
  assign new_n1798_ = new_n800_;
  assign new_n1799_ = new_n1798_;
  assign new_n1800_ = new_n1798_;
  assign new_n1801_ = new_n801_;
  assign new_n1802_ = new_n1801_;
  assign new_n1803_ = new_n1801_;
  assign new_n1804_ = new_n698_;
  assign new_n1805_ = new_n1804_;
  assign new_n1806_ = new_n1804_;
  assign new_n1807_ = new_n1032_;
  assign new_n1808_ = new_n1807_;
  assign new_n1809_ = new_n1807_;
  assign new_n1810_ = new_n699_;
  assign new_n1811_ = new_n1810_;
  assign new_n1812_ = new_n1810_;
  assign new_n1813_ = new_n1033_;
  assign new_n1814_ = new_n1813_;
  assign new_n1815_ = new_n1813_;
  assign new_n1816_ = new_n700_;
  assign new_n1817_ = new_n1816_;
  assign new_n1818_ = new_n1816_;
  assign new_n1819_ = new_n701_;
  assign new_n1820_ = new_n1819_;
  assign new_n1821_ = new_n1819_;
  assign new_n1822_ = new_n702_;
  assign new_n1823_ = new_n1822_;
  assign new_n1824_ = new_n1822_;
  assign new_n1825_ = new_n703_;
  assign new_n1826_ = new_n1825_;
  assign new_n1827_ = new_n1825_;
  assign new_n1828_ = new_n704_;
  assign new_n1829_ = new_n1828_;
  assign new_n1830_ = new_n1828_;
  assign new_n1831_ = new_n705_;
  assign new_n1832_ = new_n1831_;
  assign new_n1833_ = new_n1831_;
  assign new_n1834_ = new_n1056_;
  assign new_n1835_ = new_n1834_;
  assign new_n1836_ = new_n1834_;
  assign new_n1837_ = new_n1057_;
  assign new_n1838_ = new_n1837_;
  assign new_n1839_ = new_n1837_;
  assign new_n1840_ = new_n1080_;
  assign new_n1841_ = new_n1840_;
  assign new_n1842_ = new_n1840_;
  assign new_n1843_ = new_n1081_;
  assign new_n1844_ = new_n1843_;
  assign new_n1845_ = new_n1843_;
  assign new_n1846_ = new_n1104_;
  assign new_n1847_ = new_n1846_;
  assign new_n1848_ = new_n1846_;
  assign new_n1849_ = new_n1105_;
  assign new_n1850_ = new_n1849_;
  assign new_n1851_ = new_n1849_;
  assign new_n1852_ = new_n1129_;
  assign new_n1853_ = new_n1852_;
  assign new_n1854_ = new_n1131_;
  assign new_n1855_ = new_n1854_;
  assign new_n1856_ = new_n1134_;
  assign new_n1857_ = new_n1856_;
  assign new_n1858_ = new_n1140_;
  assign new_n1859_ = new_n1858_;
  assign new_n1860_ = new_n1135_;
  assign new_n1861_ = new_n1860_;
  assign new_n1862_ = new_n1141_;
  assign new_n1863_ = new_n1862_;
  assign new_n1864_ = new_n1136_;
  assign new_n1865_ = new_n1864_;
  assign new_n1866_ = new_n1138_;
  assign new_n1867_ = new_n1866_;
  assign new_n1868_ = new_n1127_;
  assign new_n1869_ = new_n1868_;
  assign new_n1870_ = new_n1143_;
  assign new_n1871_ = new_n1133_;
  assign new_n1872_ = new_n1871_;
  assign new_n1873_ = new_n1149_;
  assign new_n1874_ = new_n1142_;
  assign new_n1875_ = new_n1137_;
  assign new_n1876_ = new_n1875_;
  assign new_n1877_ = new_n1139_;
  assign new_n1878_ = new_n1877_;
  assign new_n1879_ = new_n1148_;
  assign new_n1880_ = new_n1150_;
  assign new_n1881_ = new_n1151_;
  assign new_n1882_ = new_n1144_;
  assign new_n1883_ = new_n1146_;
  assign new_n1884_ = new_n1153_;
  assign new_n1885_ = new_n1147_;
  assign new_n1886_ = new_n724_;
  assign new_n1887_ = new_n1886_;
  assign new_n1888_ = new_n733_;
  assign new_n1889_ = new_n725_;
  assign new_n1890_ = new_n732_;
  assign new_n1891_ = new_n1890_;
  assign new_n1892_ = new_n740_;
  assign new_n1893_ = new_n1892_;
  assign new_n1894_ = new_n749_;
  assign new_n1895_ = new_n741_;
  assign new_n1896_ = new_n748_;
  assign new_n1897_ = new_n1896_;
  assign new_n1898_ = new_n850_;
  assign new_n1899_ = new_n1898_;
  assign new_n1900_ = new_n1899_;
  assign new_n1901_ = new_n1899_;
  assign new_n1902_ = new_n1898_;
  assign new_n1903_ = new_n1902_;
  assign new_n1904_ = new_n1902_;
  assign new_n1905_ = new_n851_;
  assign new_n1906_ = new_n1905_;
  assign new_n1907_ = new_n1906_;
  assign new_n1908_ = new_n1906_;
  assign new_n1909_ = new_n1905_;
  assign new_n1910_ = new_n1909_;
  assign new_n1911_ = new_n1909_;
  assign new_n1912_ = new_n861_;
  assign new_n1913_ = new_n1912_;
  assign new_n1914_ = new_n1912_;
  assign new_n1915_ = new_n862_;
  assign new_n1916_ = new_n1915_;
  assign new_n1917_ = new_n1915_;
  assign new_n1918_ = new_n860_;
  assign new_n1919_ = new_n1918_;
  assign new_n1920_ = new_n1918_;
  assign new_n1921_ = new_n863_;
  assign new_n1922_ = new_n1921_;
  assign new_n1923_ = new_n1921_;
  assign new_n1924_ = new_n1182_;
  assign new_n1925_ = new_n1193_;
  assign new_n1926_ = new_n726_;
  assign new_n1927_ = new_n1926_;
  assign new_n1928_ = new_n735_;
  assign new_n1929_ = new_n727_;
  assign new_n1930_ = new_n734_;
  assign new_n1931_ = new_n1930_;
  assign new_n1932_ = new_n742_;
  assign new_n1933_ = new_n1932_;
  assign new_n1934_ = new_n751_;
  assign new_n1935_ = new_n743_;
  assign new_n1936_ = new_n750_;
  assign new_n1937_ = new_n1936_;
  assign new_n1938_ = new_n864_;
  assign new_n1939_ = new_n1938_;
  assign new_n1940_ = new_n1938_;
  assign new_n1941_ = new_n867_;
  assign new_n1942_ = new_n1941_;
  assign new_n1943_ = new_n1941_;
  assign new_n1944_ = new_n865_;
  assign new_n1945_ = new_n1944_;
  assign new_n1946_ = new_n1944_;
  assign new_n1947_ = new_n866_;
  assign new_n1948_ = new_n1947_;
  assign new_n1949_ = new_n1947_;
  assign new_n1950_ = new_n1210_;
  assign new_n1951_ = new_n1221_;
  assign new_n1952_ = new_n728_;
  assign new_n1953_ = new_n1952_;
  assign new_n1954_ = new_n737_;
  assign new_n1955_ = new_n729_;
  assign new_n1956_ = new_n736_;
  assign new_n1957_ = new_n1956_;
  assign new_n1958_ = new_n744_;
  assign new_n1959_ = new_n1958_;
  assign new_n1960_ = new_n753_;
  assign new_n1961_ = new_n745_;
  assign new_n1962_ = new_n752_;
  assign new_n1963_ = new_n1962_;
  assign new_n1964_ = new_n1238_;
  assign new_n1965_ = new_n1249_;
  assign new_n1966_ = new_n730_;
  assign new_n1967_ = new_n1966_;
  assign new_n1968_ = new_n739_;
  assign new_n1969_ = new_n731_;
  assign new_n1970_ = new_n738_;
  assign new_n1971_ = new_n1970_;
  assign new_n1972_ = new_n746_;
  assign new_n1973_ = new_n1972_;
  assign new_n1974_ = new_n755_;
  assign new_n1975_ = new_n747_;
  assign new_n1976_ = new_n754_;
  assign new_n1977_ = new_n1976_;
  assign new_n1978_ = new_n1266_;
  assign new_n1979_ = new_n1277_;
  assign new_n1980_ = new_n756_;
  assign new_n1981_ = new_n1980_;
  assign new_n1982_ = new_n765_;
  assign new_n1983_ = new_n757_;
  assign new_n1984_ = new_n764_;
  assign new_n1985_ = new_n1984_;
  assign new_n1986_ = new_n772_;
  assign new_n1987_ = new_n1986_;
  assign new_n1988_ = new_n781_;
  assign new_n1989_ = new_n773_;
  assign new_n1990_ = new_n780_;
  assign new_n1991_ = new_n1990_;
  assign new_n1992_ = new_n853_;
  assign new_n1993_ = new_n1992_;
  assign new_n1994_ = new_n1992_;
  assign new_n1995_ = new_n854_;
  assign new_n1996_ = new_n1995_;
  assign new_n1997_ = new_n1995_;
  assign new_n1998_ = new_n852_;
  assign new_n1999_ = new_n1998_;
  assign new_n2000_ = new_n1998_;
  assign new_n2001_ = new_n855_;
  assign new_n2002_ = new_n2001_;
  assign new_n2003_ = new_n2001_;
  assign new_n2004_ = new_n1294_;
  assign new_n2005_ = new_n1305_;
  assign new_n2006_ = new_n758_;
  assign new_n2007_ = new_n2006_;
  assign new_n2008_ = new_n767_;
  assign new_n2009_ = new_n759_;
  assign new_n2010_ = new_n766_;
  assign new_n2011_ = new_n2010_;
  assign new_n2012_ = new_n774_;
  assign new_n2013_ = new_n2012_;
  assign new_n2014_ = new_n783_;
  assign new_n2015_ = new_n775_;
  assign new_n2016_ = new_n782_;
  assign new_n2017_ = new_n2016_;
  assign new_n2018_ = new_n857_;
  assign new_n2019_ = new_n2018_;
  assign new_n2020_ = new_n2018_;
  assign new_n2021_ = new_n858_;
  assign new_n2022_ = new_n2021_;
  assign new_n2023_ = new_n2021_;
  assign new_n2024_ = new_n856_;
  assign new_n2025_ = new_n2024_;
  assign new_n2026_ = new_n2024_;
  assign new_n2027_ = new_n859_;
  assign new_n2028_ = new_n2027_;
  assign new_n2029_ = new_n2027_;
  assign new_n2030_ = new_n1322_;
  assign new_n2031_ = new_n1333_;
  assign new_n2032_ = new_n760_;
  assign new_n2033_ = new_n2032_;
  assign new_n2034_ = new_n769_;
  assign new_n2035_ = new_n761_;
  assign new_n2036_ = new_n768_;
  assign new_n2037_ = new_n2036_;
  assign new_n2038_ = new_n776_;
  assign new_n2039_ = new_n2038_;
  assign new_n2040_ = new_n785_;
  assign new_n2041_ = new_n777_;
  assign new_n2042_ = new_n784_;
  assign new_n2043_ = new_n2042_;
  assign new_n2044_ = new_n1350_;
  assign new_n2045_ = new_n1361_;
  assign new_n2046_ = new_n762_;
  assign new_n2047_ = new_n2046_;
  assign new_n2048_ = new_n771_;
  assign new_n2049_ = new_n763_;
  assign new_n2050_ = new_n770_;
  assign new_n2051_ = new_n2050_;
  assign new_n2052_ = new_n778_;
  assign new_n2053_ = new_n2052_;
  assign new_n2054_ = new_n787_;
  assign new_n2055_ = new_n779_;
  assign new_n2056_ = new_n786_;
  assign new_n2057_ = new_n2056_;
  assign new_n2058_ = new_n1378_;
  assign new_n2059_ = new_n1389_;
  assign new_n2060_ = new_n868_;
  assign new_n2061_ = new_n2060_;
  assign new_n2062_ = new_n871_;
  assign new_n2063_ = new_n869_;
  assign new_n2064_ = new_n870_;
  assign new_n2065_ = new_n2064_;
  assign new_n2066_ = new_n872_;
  assign new_n2067_ = new_n2066_;
  assign new_n2068_ = new_n875_;
  assign new_n2069_ = new_n873_;
  assign new_n2070_ = new_n874_;
  assign new_n2071_ = new_n2070_;
  assign new_n2072_ = new_n876_;
  assign new_n2073_ = new_n2072_;
  assign new_n2074_ = new_n879_;
  assign new_n2075_ = new_n877_;
  assign new_n2076_ = new_n878_;
  assign new_n2077_ = new_n2076_;
  assign new_n2078_ = new_n880_;
  assign new_n2079_ = new_n2078_;
  assign new_n2080_ = new_n883_;
  assign new_n2081_ = new_n881_;
  assign new_n2082_ = new_n882_;
  assign new_n2083_ = new_n2082_;
  assign new_n2084_ = new_n884_;
  assign new_n2085_ = new_n2084_;
  assign new_n2086_ = new_n887_;
  assign new_n2087_ = new_n885_;
  assign new_n2088_ = new_n886_;
  assign new_n2089_ = new_n2088_;
  assign new_n2090_ = new_n888_;
  assign new_n2091_ = new_n2090_;
  assign new_n2092_ = new_n891_;
  assign new_n2093_ = new_n889_;
  assign new_n2094_ = new_n890_;
  assign new_n2095_ = new_n2094_;
  assign new_n2096_ = new_n892_;
  assign new_n2097_ = new_n2096_;
  assign new_n2098_ = new_n895_;
  assign new_n2099_ = new_n893_;
  assign new_n2100_ = new_n894_;
  assign new_n2101_ = new_n2100_;
  assign new_n2102_ = new_n896_;
  assign new_n2103_ = new_n2102_;
  assign new_n2104_ = new_n899_;
  assign new_n2105_ = new_n897_;
  assign new_n2106_ = new_n898_;
  assign new_n2107_ = new_n2106_;
  assign new_n2108_ = new_n900_;
  assign new_n2109_ = new_n2108_;
  assign new_n2110_ = new_n903_;
  assign new_n2111_ = new_n901_;
  assign new_n2112_ = new_n902_;
  assign new_n2113_ = new_n2112_;
  assign new_n2114_ = new_n904_;
  assign new_n2115_ = new_n2114_;
  assign new_n2116_ = new_n907_;
  assign new_n2117_ = new_n905_;
  assign new_n2118_ = new_n906_;
  assign new_n2119_ = new_n2118_;
  assign new_n2120_ = new_n908_;
  assign new_n2121_ = new_n2120_;
  assign new_n2122_ = new_n911_;
  assign new_n2123_ = new_n909_;
  assign new_n2124_ = new_n910_;
  assign new_n2125_ = new_n2124_;
  assign new_n2126_ = new_n912_;
  assign new_n2127_ = new_n2126_;
  assign new_n2128_ = new_n915_;
  assign new_n2129_ = new_n913_;
  assign new_n2130_ = new_n914_;
  assign new_n2131_ = new_n2130_;
  assign new_n2132_ = new_n916_;
  assign new_n2133_ = new_n2132_;
  assign new_n2134_ = new_n919_;
  assign new_n2135_ = new_n917_;
  assign new_n2136_ = new_n918_;
  assign new_n2137_ = new_n2136_;
  assign new_n2138_ = new_n920_;
  assign new_n2139_ = new_n2138_;
  assign new_n2140_ = new_n923_;
  assign new_n2141_ = new_n921_;
  assign new_n2142_ = new_n922_;
  assign new_n2143_ = new_n2142_;
  assign new_n2144_ = new_n924_;
  assign new_n2145_ = new_n2144_;
  assign new_n2146_ = new_n927_;
  assign new_n2147_ = new_n925_;
  assign new_n2148_ = new_n926_;
  assign new_n2149_ = new_n2148_;
  assign new_n2150_ = new_n928_;
  assign new_n2151_ = new_n2150_;
  assign new_n2152_ = new_n931_;
  assign new_n2153_ = new_n929_;
  assign new_n2154_ = new_n930_;
  assign new_n2155_ = new_n2154_;
  always @ (posedge clock) begin
    n286_lo <= n1020_li003_li003;
    n298_lo <= n1032_li007_li007;
    n310_lo <= n1044_li011_li011;
    n322_lo <= n1056_li015_li015;
    n334_lo <= n1068_li019_li019;
    n346_lo <= n1080_li023_li023;
    n358_lo <= n1092_li027_li027;
    n370_lo <= n1104_li031_li031;
    n382_lo <= n1116_li035_li035;
    n394_lo <= n1128_li039_li039;
    n406_lo <= n1140_li043_li043;
    n418_lo <= n1152_li047_li047;
    n430_lo <= n1164_li051_li051;
    n442_lo <= n1176_li055_li055;
    n454_lo <= n1188_li059_li059;
    n466_lo <= n1200_li063_li063;
    n478_lo <= n1212_li067_li067;
    n490_lo <= n1224_li071_li071;
    n502_lo <= n1236_li075_li075;
    n514_lo <= n1248_li079_li079;
    n526_lo <= n1260_li083_li083;
    n538_lo <= n1272_li087_li087;
    n550_lo <= n1284_li091_li091;
    n562_lo <= n1296_li095_li095;
    n574_lo <= n1308_li099_li099;
    n586_lo <= n1320_li103_li103;
    n598_lo <= n1332_li107_li107;
    n610_lo <= n1344_li111_li111;
    n622_lo <= n1356_li115_li115;
    n634_lo <= n1368_li119_li119;
    n646_lo <= n1380_li123_li123;
    n658_lo <= n1392_li127_li127;
    n661_lo <= n1395_li128_li128;
    n673_lo <= n1407_li132_li132;
    n685_lo <= n1419_li136_li136;
    n697_lo <= n1431_li140_li140;
    n709_lo <= n1443_li144_li144;
    n721_lo <= n1455_li148_li148;
    n733_lo <= n1467_li152_li152;
    n745_lo <= n1479_li156_li156;
    n757_lo <= n1491_li160_li160;
    n1589_o2 <= n1589_i2;
    n1590_o2 <= n1590_i2;
    n1591_o2 <= n1591_i2;
    n1592_o2 <= n1592_i2;
    n1593_o2 <= n1593_i2;
    n1594_o2 <= n1594_i2;
    n1595_o2 <= n1595_i2;
    n1596_o2 <= n1596_i2;
    n1597_o2 <= n1597_i2;
    n1598_o2 <= n1598_i2;
    n1599_o2 <= n1599_i2;
    n1600_o2 <= n1600_i2;
    n1601_o2 <= n1601_i2;
    n1602_o2 <= n1602_i2;
    n1603_o2 <= n1603_i2;
    n1604_o2 <= n1604_i2;
    n1605_o2 <= n1605_i2;
    n1606_o2 <= n1606_i2;
    n1607_o2 <= n1607_i2;
    n1608_o2 <= n1608_i2;
    n1609_o2 <= n1609_i2;
    n1610_o2 <= n1610_i2;
    n1611_o2 <= n1611_i2;
    n1612_o2 <= n1612_i2;
    n1613_o2 <= n1613_i2;
    n1614_o2 <= n1614_i2;
    n1615_o2 <= n1615_i2;
    n1616_o2 <= n1616_i2;
    n1617_o2 <= n1617_i2;
    n1618_o2 <= n1618_i2;
    n1619_o2 <= n1619_i2;
    n1620_o2 <= n1620_i2;
    n602_o2 <= n602_i2;
    n639_o2 <= n639_i2;
    n678_o2 <= n678_i2;
    n658_o2 <= n658_i2;
    n783_o2 <= n783_i2;
    n802_o2 <= n802_i2;
    n726_o2 <= n726_i2;
    n763_o2 <= n763_i2;
    n685_o2 <= n685_i2;
    n680_o2 <= n680_i2;
    n822_o2 <= n822_i2;
    n843_o2 <= n843_i2;
    n842_o2 <= n842_i2;
    n681_o2 <= n681_i2;
    n684_o2 <= n684_i2;
    n686_o2 <= n686_i2;
    n823_o2 <= n823_i2;
    lo002_buf_o2 <= lo002_buf_i2;
    lo006_buf_o2 <= lo006_buf_i2;
    lo010_buf_o2 <= lo010_buf_i2;
    lo014_buf_o2 <= lo014_buf_i2;
    lo018_buf_o2 <= lo018_buf_i2;
    lo022_buf_o2 <= lo022_buf_i2;
    lo026_buf_o2 <= lo026_buf_i2;
    lo030_buf_o2 <= lo030_buf_i2;
    lo034_buf_o2 <= lo034_buf_i2;
    lo038_buf_o2 <= lo038_buf_i2;
    lo042_buf_o2 <= lo042_buf_i2;
    lo046_buf_o2 <= lo046_buf_i2;
    lo050_buf_o2 <= lo050_buf_i2;
    lo054_buf_o2 <= lo054_buf_i2;
    lo058_buf_o2 <= lo058_buf_i2;
    lo062_buf_o2 <= lo062_buf_i2;
    lo066_buf_o2 <= lo066_buf_i2;
    lo070_buf_o2 <= lo070_buf_i2;
    lo074_buf_o2 <= lo074_buf_i2;
    lo078_buf_o2 <= lo078_buf_i2;
    lo082_buf_o2 <= lo082_buf_i2;
    lo086_buf_o2 <= lo086_buf_i2;
    lo090_buf_o2 <= lo090_buf_i2;
    lo094_buf_o2 <= lo094_buf_i2;
    lo098_buf_o2 <= lo098_buf_i2;
    lo102_buf_o2 <= lo102_buf_i2;
    lo106_buf_o2 <= lo106_buf_i2;
    lo110_buf_o2 <= lo110_buf_i2;
    lo114_buf_o2 <= lo114_buf_i2;
    lo118_buf_o2 <= lo118_buf_i2;
    lo122_buf_o2 <= lo122_buf_i2;
    lo126_buf_o2 <= lo126_buf_i2;
    n683_o2 <= n683_i2;
    n688_o2 <= n688_i2;
    n803_o2 <= n803_i2;
    n862_o2 <= n862_i2;
    n764_o2 <= n764_i2;
    n863_o2 <= n863_i2;
    n886_o2 <= n886_i2;
    n600_o2 <= n600_i2;
    n601_o2 <= n601_i2;
    n637_o2 <= n637_i2;
    n638_o2 <= n638_i2;
    n676_o2 <= n676_i2;
    n677_o2 <= n677_i2;
    n656_o2 <= n656_i2;
    n657_o2 <= n657_i2;
    n781_o2 <= n781_i2;
    n782_o2 <= n782_i2;
    n800_o2 <= n800_i2;
    n801_o2 <= n801_i2;
    n724_o2 <= n724_i2;
    n725_o2 <= n725_i2;
    n761_o2 <= n761_i2;
    n762_o2 <= n762_i2;
    lo129_buf_o2 <= lo129_buf_i2;
    lo133_buf_o2 <= lo133_buf_i2;
    lo137_buf_o2 <= lo137_buf_i2;
    lo141_buf_o2 <= lo141_buf_i2;
    lo145_buf_o2 <= lo145_buf_i2;
    lo149_buf_o2 <= lo149_buf_i2;
    lo153_buf_o2 <= lo153_buf_i2;
    lo157_buf_o2 <= lo157_buf_i2;
    lo161_buf_o2 <= lo161_buf_i2;
    n708_o2 <= n708_i2;
    n745_o2 <= n745_i2;
    n717_o2 <= n717_i2;
    n754_o2 <= n754_i2;
    n584_o2 <= n584_i2;
    n593_o2 <= n593_i2;
    n630_o2 <= n630_i2;
    n621_o2 <= n621_i2;
    lo001_buf_o2 <= lo001_buf_i2;
    lo005_buf_o2 <= lo005_buf_i2;
    lo009_buf_o2 <= lo009_buf_i2;
    lo013_buf_o2 <= lo013_buf_i2;
    lo017_buf_o2 <= lo017_buf_i2;
    lo021_buf_o2 <= lo021_buf_i2;
    lo025_buf_o2 <= lo025_buf_i2;
    lo029_buf_o2 <= lo029_buf_i2;
    lo033_buf_o2 <= lo033_buf_i2;
    lo037_buf_o2 <= lo037_buf_i2;
    lo041_buf_o2 <= lo041_buf_i2;
    lo045_buf_o2 <= lo045_buf_i2;
    lo049_buf_o2 <= lo049_buf_i2;
    lo053_buf_o2 <= lo053_buf_i2;
    lo057_buf_o2 <= lo057_buf_i2;
    lo061_buf_o2 <= lo061_buf_i2;
    lo065_buf_o2 <= lo065_buf_i2;
    lo069_buf_o2 <= lo069_buf_i2;
    lo073_buf_o2 <= lo073_buf_i2;
    lo077_buf_o2 <= lo077_buf_i2;
    lo081_buf_o2 <= lo081_buf_i2;
    lo085_buf_o2 <= lo085_buf_i2;
    lo089_buf_o2 <= lo089_buf_i2;
    lo093_buf_o2 <= lo093_buf_i2;
    lo097_buf_o2 <= lo097_buf_i2;
    lo101_buf_o2 <= lo101_buf_i2;
    lo105_buf_o2 <= lo105_buf_i2;
    lo109_buf_o2 <= lo109_buf_i2;
    lo113_buf_o2 <= lo113_buf_i2;
    lo117_buf_o2 <= lo117_buf_i2;
    lo121_buf_o2 <= lo121_buf_i2;
    lo125_buf_o2 <= lo125_buf_i2;
  end
  initial begin
    n286_lo <= 1'b0;
    n298_lo <= 1'b0;
    n310_lo <= 1'b0;
    n322_lo <= 1'b0;
    n334_lo <= 1'b0;
    n346_lo <= 1'b0;
    n358_lo <= 1'b0;
    n370_lo <= 1'b0;
    n382_lo <= 1'b0;
    n394_lo <= 1'b0;
    n406_lo <= 1'b0;
    n418_lo <= 1'b0;
    n430_lo <= 1'b0;
    n442_lo <= 1'b0;
    n454_lo <= 1'b0;
    n466_lo <= 1'b0;
    n478_lo <= 1'b0;
    n490_lo <= 1'b0;
    n502_lo <= 1'b0;
    n514_lo <= 1'b0;
    n526_lo <= 1'b0;
    n538_lo <= 1'b0;
    n550_lo <= 1'b0;
    n562_lo <= 1'b0;
    n574_lo <= 1'b0;
    n586_lo <= 1'b0;
    n598_lo <= 1'b0;
    n610_lo <= 1'b0;
    n622_lo <= 1'b0;
    n634_lo <= 1'b0;
    n646_lo <= 1'b0;
    n658_lo <= 1'b0;
    n661_lo <= 1'b0;
    n673_lo <= 1'b0;
    n685_lo <= 1'b0;
    n697_lo <= 1'b0;
    n709_lo <= 1'b0;
    n721_lo <= 1'b0;
    n733_lo <= 1'b0;
    n745_lo <= 1'b0;
    n757_lo <= 1'b0;
    n1589_o2 <= 1'b0;
    n1590_o2 <= 1'b0;
    n1591_o2 <= 1'b0;
    n1592_o2 <= 1'b0;
    n1593_o2 <= 1'b0;
    n1594_o2 <= 1'b0;
    n1595_o2 <= 1'b0;
    n1596_o2 <= 1'b0;
    n1597_o2 <= 1'b0;
    n1598_o2 <= 1'b0;
    n1599_o2 <= 1'b0;
    n1600_o2 <= 1'b0;
    n1601_o2 <= 1'b0;
    n1602_o2 <= 1'b0;
    n1603_o2 <= 1'b0;
    n1604_o2 <= 1'b0;
    n1605_o2 <= 1'b0;
    n1606_o2 <= 1'b0;
    n1607_o2 <= 1'b0;
    n1608_o2 <= 1'b0;
    n1609_o2 <= 1'b0;
    n1610_o2 <= 1'b0;
    n1611_o2 <= 1'b0;
    n1612_o2 <= 1'b0;
    n1613_o2 <= 1'b0;
    n1614_o2 <= 1'b0;
    n1615_o2 <= 1'b0;
    n1616_o2 <= 1'b0;
    n1617_o2 <= 1'b0;
    n1618_o2 <= 1'b0;
    n1619_o2 <= 1'b0;
    n1620_o2 <= 1'b0;
    n602_o2 <= 1'b0;
    n639_o2 <= 1'b0;
    n678_o2 <= 1'b0;
    n658_o2 <= 1'b0;
    n783_o2 <= 1'b0;
    n802_o2 <= 1'b0;
    n726_o2 <= 1'b0;
    n763_o2 <= 1'b0;
    n685_o2 <= 1'b0;
    n680_o2 <= 1'b0;
    n822_o2 <= 1'b0;
    n843_o2 <= 1'b0;
    n842_o2 <= 1'b0;
    n681_o2 <= 1'b0;
    n684_o2 <= 1'b0;
    n686_o2 <= 1'b0;
    n823_o2 <= 1'b0;
    lo002_buf_o2 <= 1'b0;
    lo006_buf_o2 <= 1'b0;
    lo010_buf_o2 <= 1'b0;
    lo014_buf_o2 <= 1'b0;
    lo018_buf_o2 <= 1'b0;
    lo022_buf_o2 <= 1'b0;
    lo026_buf_o2 <= 1'b0;
    lo030_buf_o2 <= 1'b0;
    lo034_buf_o2 <= 1'b0;
    lo038_buf_o2 <= 1'b0;
    lo042_buf_o2 <= 1'b0;
    lo046_buf_o2 <= 1'b0;
    lo050_buf_o2 <= 1'b0;
    lo054_buf_o2 <= 1'b0;
    lo058_buf_o2 <= 1'b0;
    lo062_buf_o2 <= 1'b0;
    lo066_buf_o2 <= 1'b0;
    lo070_buf_o2 <= 1'b0;
    lo074_buf_o2 <= 1'b0;
    lo078_buf_o2 <= 1'b0;
    lo082_buf_o2 <= 1'b0;
    lo086_buf_o2 <= 1'b0;
    lo090_buf_o2 <= 1'b0;
    lo094_buf_o2 <= 1'b0;
    lo098_buf_o2 <= 1'b0;
    lo102_buf_o2 <= 1'b0;
    lo106_buf_o2 <= 1'b0;
    lo110_buf_o2 <= 1'b0;
    lo114_buf_o2 <= 1'b0;
    lo118_buf_o2 <= 1'b0;
    lo122_buf_o2 <= 1'b0;
    lo126_buf_o2 <= 1'b0;
    n683_o2 <= 1'b0;
    n688_o2 <= 1'b0;
    n803_o2 <= 1'b0;
    n862_o2 <= 1'b0;
    n764_o2 <= 1'b0;
    n863_o2 <= 1'b0;
    n886_o2 <= 1'b0;
    n600_o2 <= 1'b0;
    n601_o2 <= 1'b0;
    n637_o2 <= 1'b0;
    n638_o2 <= 1'b0;
    n676_o2 <= 1'b0;
    n677_o2 <= 1'b0;
    n656_o2 <= 1'b0;
    n657_o2 <= 1'b0;
    n781_o2 <= 1'b0;
    n782_o2 <= 1'b0;
    n800_o2 <= 1'b0;
    n801_o2 <= 1'b0;
    n724_o2 <= 1'b0;
    n725_o2 <= 1'b0;
    n761_o2 <= 1'b0;
    n762_o2 <= 1'b0;
    lo129_buf_o2 <= 1'b0;
    lo133_buf_o2 <= 1'b0;
    lo137_buf_o2 <= 1'b0;
    lo141_buf_o2 <= 1'b0;
    lo145_buf_o2 <= 1'b0;
    lo149_buf_o2 <= 1'b0;
    lo153_buf_o2 <= 1'b0;
    lo157_buf_o2 <= 1'b0;
    lo161_buf_o2 <= 1'b0;
    n708_o2 <= 1'b0;
    n745_o2 <= 1'b0;
    n717_o2 <= 1'b0;
    n754_o2 <= 1'b0;
    n584_o2 <= 1'b0;
    n593_o2 <= 1'b0;
    n630_o2 <= 1'b0;
    n621_o2 <= 1'b0;
    lo001_buf_o2 <= 1'b0;
    lo005_buf_o2 <= 1'b0;
    lo009_buf_o2 <= 1'b0;
    lo013_buf_o2 <= 1'b0;
    lo017_buf_o2 <= 1'b0;
    lo021_buf_o2 <= 1'b0;
    lo025_buf_o2 <= 1'b0;
    lo029_buf_o2 <= 1'b0;
    lo033_buf_o2 <= 1'b0;
    lo037_buf_o2 <= 1'b0;
    lo041_buf_o2 <= 1'b0;
    lo045_buf_o2 <= 1'b0;
    lo049_buf_o2 <= 1'b0;
    lo053_buf_o2 <= 1'b0;
    lo057_buf_o2 <= 1'b0;
    lo061_buf_o2 <= 1'b0;
    lo065_buf_o2 <= 1'b0;
    lo069_buf_o2 <= 1'b0;
    lo073_buf_o2 <= 1'b0;
    lo077_buf_o2 <= 1'b0;
    lo081_buf_o2 <= 1'b0;
    lo085_buf_o2 <= 1'b0;
    lo089_buf_o2 <= 1'b0;
    lo093_buf_o2 <= 1'b0;
    lo097_buf_o2 <= 1'b0;
    lo101_buf_o2 <= 1'b0;
    lo105_buf_o2 <= 1'b0;
    lo109_buf_o2 <= 1'b0;
    lo113_buf_o2 <= 1'b0;
    lo117_buf_o2 <= 1'b0;
    lo121_buf_o2 <= 1'b0;
    lo125_buf_o2 <= 1'b0;
  end
endmodule


