
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  G42,
  G43,
  G44,
  G45,
  G46,
  G47,
  G48,
  G49,
  G50,
  G51,
  G52,
  G53,
  G54,
  G55,
  G56,
  G57,
  G58,
  G59,
  G60,
  G61,
  G62,
  G63,
  G64,
  G65,
  G66,
  G67,
  G68,
  G69,
  G70,
  G71,
  G72,
  G73,
  G74,
  G75,
  G76,
  G77,
  G78,
  G79,
  G80,
  G81,
  G82,
  G83,
  G84,
  G85,
  G86,
  G87,
  G88,
  G89,
  G90,
  G91,
  G92,
  G93,
  G94,
  G95,
  G96,
  G97,
  G98,
  G99,
  G100,
  G101,
  G102,
  G103,
  G104,
  G105,
  G106,
  G107,
  G108,
  G109,
  G110,
  G111,
  G112,
  G113,
  G114,
  G115,
  G116,
  G117,
  G118,
  G119,
  G120,
  G121,
  G122,
  G123,
  G124,
  G125,
  G126,
  G127,
  G128,
  G129,
  G130,
  G131,
  G132,
  G133,
  G134,
  G135,
  G136,
  G137,
  G138,
  G139,
  G140,
  G141,
  G142,
  G143,
  G144,
  G145,
  G146,
  G147,
  G148,
  G149,
  G150,
  G151,
  G152,
  G153,
  G154,
  G155,
  G156,
  G157,
  G158,
  G159,
  G160,
  G161,
  G162,
  G163,
  G164,
  G165,
  G166,
  G167,
  G168,
  G169,
  G170,
  G171,
  G172,
  G173,
  G174,
  G175,
  G176,
  G177,
  G178,
  G5193,
  G5194,
  G5195,
  G5196,
  G5197,
  G5198,
  G5199,
  G5200,
  G5201,
  G5202,
  G5203,
  G5204,
  G5205,
  G5206,
  G5207,
  G5208,
  G5209,
  G5210,
  G5211,
  G5212,
  G5213,
  G5214,
  G5215,
  G5216,
  G5217,
  G5218,
  G5219,
  G5220,
  G5221,
  G5222,
  G5223,
  G5224,
  G5225,
  G5226,
  G5227,
  G5228,
  G5229,
  G5230,
  G5231,
  G5232,
  G5233,
  G5234,
  G5235,
  G5236,
  G5237,
  G5238,
  G5239,
  G5240,
  G5241,
  G5242,
  G5243,
  G5244,
  G5245,
  G5246,
  G5247,
  G5248,
  G5249,
  G5250,
  G5251,
  G5252,
  G5253,
  G5254,
  G5255,
  G5256,
  G5257,
  G5258,
  G5259,
  G5260,
  G5261,
  G5262,
  G5263,
  G5264,
  G5265,
  G5266,
  G5267,
  G5268,
  G5269,
  G5270,
  G5271,
  G5272,
  G5273,
  G5274,
  G5275,
  G5276,
  G5277,
  G5278,
  G5279,
  G5280,
  G5281,
  G5282,
  G5283,
  G5284,
  G5285,
  G5286,
  G5287,
  G5288,
  G5289,
  G5290,
  G5291,
  G5292,
  G5293,
  G5294,
  G5295,
  G5296,
  G5297,
  G5298,
  G5299,
  G5300,
  G5301,
  G5302,
  G5303,
  G5304,
  G5305,
  G5306,
  G5307,
  G5308,
  G5309,
  G5310,
  G5311,
  G5312,
  G5313,
  G5314,
  G5315
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input G42;input G43;input G44;input G45;input G46;input G47;input G48;input G49;input G50;input G51;input G52;input G53;input G54;input G55;input G56;input G57;input G58;input G59;input G60;input G61;input G62;input G63;input G64;input G65;input G66;input G67;input G68;input G69;input G70;input G71;input G72;input G73;input G74;input G75;input G76;input G77;input G78;input G79;input G80;input G81;input G82;input G83;input G84;input G85;input G86;input G87;input G88;input G89;input G90;input G91;input G92;input G93;input G94;input G95;input G96;input G97;input G98;input G99;input G100;input G101;input G102;input G103;input G104;input G105;input G106;input G107;input G108;input G109;input G110;input G111;input G112;input G113;input G114;input G115;input G116;input G117;input G118;input G119;input G120;input G121;input G122;input G123;input G124;input G125;input G126;input G127;input G128;input G129;input G130;input G131;input G132;input G133;input G134;input G135;input G136;input G137;input G138;input G139;input G140;input G141;input G142;input G143;input G144;input G145;input G146;input G147;input G148;input G149;input G150;input G151;input G152;input G153;input G154;input G155;input G156;input G157;input G158;input G159;input G160;input G161;input G162;input G163;input G164;input G165;input G166;input G167;input G168;input G169;input G170;input G171;input G172;input G173;input G174;input G175;input G176;input G177;input G178;
  output G5193;output G5194;output G5195;output G5196;output G5197;output G5198;output G5199;output G5200;output G5201;output G5202;output G5203;output G5204;output G5205;output G5206;output G5207;output G5208;output G5209;output G5210;output G5211;output G5212;output G5213;output G5214;output G5215;output G5216;output G5217;output G5218;output G5219;output G5220;output G5221;output G5222;output G5223;output G5224;output G5225;output G5226;output G5227;output G5228;output G5229;output G5230;output G5231;output G5232;output G5233;output G5234;output G5235;output G5236;output G5237;output G5238;output G5239;output G5240;output G5241;output G5242;output G5243;output G5244;output G5245;output G5246;output G5247;output G5248;output G5249;output G5250;output G5251;output G5252;output G5253;output G5254;output G5255;output G5256;output G5257;output G5258;output G5259;output G5260;output G5261;output G5262;output G5263;output G5264;output G5265;output G5266;output G5267;output G5268;output G5269;output G5270;output G5271;output G5272;output G5273;output G5274;output G5275;output G5276;output G5277;output G5278;output G5279;output G5280;output G5281;output G5282;output G5283;output G5284;output G5285;output G5286;output G5287;output G5288;output G5289;output G5290;output G5291;output G5292;output G5293;output G5294;output G5295;output G5296;output G5297;output G5298;output G5299;output G5300;output G5301;output G5302;output G5303;output G5304;output G5305;output G5306;output G5307;output G5308;output G5309;output G5310;output G5311;output G5312;output G5313;output G5314;output G5315;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire G51_p;
  wire G51_n;
  wire G52_p;
  wire G52_n;
  wire G53_p;
  wire G53_n;
  wire G54_p;
  wire G54_n;
  wire G55_p;
  wire G55_n;
  wire G56_p;
  wire G56_n;
  wire G57_p;
  wire G57_n;
  wire G58_p;
  wire G58_n;
  wire G59_p;
  wire G59_n;
  wire G60_p;
  wire G60_n;
  wire G61_p;
  wire G61_n;
  wire G62_p;
  wire G62_n;
  wire G63_p;
  wire G63_n;
  wire G64_p;
  wire G64_n;
  wire G65_p;
  wire G65_n;
  wire G66_p;
  wire G66_n;
  wire G67_p;
  wire G67_n;
  wire G68_p;
  wire G68_n;
  wire G69_p;
  wire G69_n;
  wire G70_p;
  wire G70_n;
  wire G71_p;
  wire G71_n;
  wire G72_p;
  wire G72_n;
  wire G73_p;
  wire G73_n;
  wire G74_p;
  wire G74_n;
  wire G75_p;
  wire G75_n;
  wire G76_p;
  wire G76_n;
  wire G77_p;
  wire G77_n;
  wire G78_p;
  wire G78_n;
  wire G79_p;
  wire G79_n;
  wire G80_p;
  wire G80_n;
  wire G81_p;
  wire G81_n;
  wire G82_p;
  wire G82_n;
  wire G83_p;
  wire G83_n;
  wire G84_p;
  wire G84_n;
  wire G85_p;
  wire G85_n;
  wire G86_p;
  wire G86_n;
  wire G87_p;
  wire G87_n;
  wire G88_p;
  wire G88_n;
  wire G89_p;
  wire G89_n;
  wire G90_p;
  wire G90_n;
  wire G91_p;
  wire G91_n;
  wire G92_p;
  wire G92_n;
  wire G93_p;
  wire G93_n;
  wire G94_p;
  wire G94_n;
  wire G95_p;
  wire G95_n;
  wire G96_p;
  wire G96_n;
  wire G97_p;
  wire G97_n;
  wire G98_p;
  wire G98_n;
  wire G99_p;
  wire G99_n;
  wire G100_p;
  wire G100_n;
  wire G101_p;
  wire G101_n;
  wire G102_p;
  wire G102_n;
  wire G103_p;
  wire G103_n;
  wire G104_p;
  wire G104_n;
  wire G105_p;
  wire G105_n;
  wire G106_p;
  wire G106_n;
  wire G107_p;
  wire G107_n;
  wire G108_p;
  wire G108_n;
  wire G109_p;
  wire G109_n;
  wire G110_p;
  wire G110_n;
  wire G111_p;
  wire G111_n;
  wire G112_p;
  wire G112_n;
  wire G113_p;
  wire G113_n;
  wire G114_p;
  wire G114_n;
  wire G115_p;
  wire G115_n;
  wire G116_p;
  wire G116_n;
  wire G117_p;
  wire G117_n;
  wire G118_p;
  wire G118_n;
  wire G119_p;
  wire G119_n;
  wire G120_p;
  wire G120_n;
  wire G121_p;
  wire G121_n;
  wire G122_p;
  wire G122_n;
  wire G123_p;
  wire G123_n;
  wire G124_p;
  wire G124_n;
  wire G125_p;
  wire G125_n;
  wire G126_p;
  wire G126_n;
  wire G127_p;
  wire G127_n;
  wire G128_p;
  wire G128_n;
  wire G129_p;
  wire G129_n;
  wire G130_p;
  wire G130_n;
  wire G131_p;
  wire G131_n;
  wire G132_p;
  wire G132_n;
  wire G133_p;
  wire G133_n;
  wire G134_p;
  wire G134_n;
  wire G135_p;
  wire G135_n;
  wire G136_p;
  wire G136_n;
  wire G137_p;
  wire G137_n;
  wire G138_p;
  wire G138_n;
  wire G139_p;
  wire G139_n;
  wire G140_p;
  wire G140_n;
  wire G141_p;
  wire G141_n;
  wire G142_p;
  wire G142_n;
  wire G143_p;
  wire G143_n;
  wire G144_p;
  wire G144_n;
  wire G145_p;
  wire G145_n;
  wire G146_p;
  wire G146_n;
  wire G147_p;
  wire G147_n;
  wire G148_p;
  wire G148_n;
  wire G149_p;
  wire G149_n;
  wire G150_p;
  wire G150_n;
  wire G151_p;
  wire G151_n;
  wire G152_p;
  wire G152_n;
  wire G153_p;
  wire G153_n;
  wire G154_p;
  wire G154_n;
  wire G155_p;
  wire G155_n;
  wire G156_p;
  wire G156_n;
  wire G157_p;
  wire G157_n;
  wire G158_p;
  wire G158_n;
  wire G159_p;
  wire G159_n;
  wire G160_p;
  wire G160_n;
  wire G161_p;
  wire G161_n;
  wire G162_p;
  wire G162_n;
  wire G163_p;
  wire G163_n;
  wire G164_p;
  wire G164_n;
  wire G165_p;
  wire G165_n;
  wire G166_p;
  wire G166_n;
  wire G167_p;
  wire G167_n;
  wire G168_p;
  wire G168_n;
  wire G169_p;
  wire G169_n;
  wire G170_p;
  wire G170_n;
  wire G171_p;
  wire G171_n;
  wire G172_p;
  wire G172_n;
  wire G173_p;
  wire G173_n;
  wire G174_p;
  wire G174_n;
  wire G175_p;
  wire G175_n;
  wire G176_p;
  wire G176_n;
  wire G177_p;
  wire G177_n;
  wire G178_p;
  wire G178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire g693_p;
  wire g693_n;
  wire g694_p;
  wire g694_n;
  wire g695_p;
  wire g695_n;
  wire g696_p;
  wire g696_n;
  wire g697_p;
  wire g697_n;
  wire g698_p;
  wire g698_n;
  wire g699_p;
  wire g699_n;
  wire g700_p;
  wire g700_n;
  wire g701_p;
  wire g701_n;
  wire g702_p;
  wire g702_n;
  wire g703_p;
  wire g703_n;
  wire g704_p;
  wire g704_n;
  wire g705_p;
  wire g705_n;
  wire g706_p;
  wire g706_n;
  wire g707_p;
  wire g707_n;
  wire g708_p;
  wire g708_n;
  wire g709_p;
  wire g709_n;
  wire g710_p;
  wire g710_n;
  wire g711_p;
  wire g711_n;
  wire g712_p;
  wire g712_n;
  wire g713_p;
  wire g713_n;
  wire g714_p;
  wire g714_n;
  wire g715_p;
  wire g715_n;
  wire g716_p;
  wire g716_n;
  wire g717_p;
  wire g717_n;
  wire g718_p;
  wire g718_n;
  wire g719_p;
  wire g719_n;
  wire g720_p;
  wire g720_n;
  wire g721_p;
  wire g721_n;
  wire g722_p;
  wire g722_n;
  wire g723_p;
  wire g723_n;
  wire g724_p;
  wire g724_n;
  wire g725_p;
  wire g725_n;
  wire g726_p;
  wire g726_n;
  wire g727_p;
  wire g727_n;
  wire g728_p;
  wire g728_n;
  wire g729_p;
  wire g729_n;
  wire g730_p;
  wire g730_n;
  wire g731_p;
  wire g731_n;
  wire g732_p;
  wire g732_n;
  wire g733_p;
  wire g733_n;
  wire g734_p;
  wire g734_n;
  wire g735_p;
  wire g735_n;
  wire g736_p;
  wire g736_n;
  wire g737_p;
  wire g737_n;
  wire g738_p;
  wire g738_n;
  wire g739_p;
  wire g739_n;
  wire g740_p;
  wire g740_n;
  wire g741_p;
  wire g741_n;
  wire g742_p;
  wire g742_n;
  wire g743_p;
  wire g743_n;
  wire g744_p;
  wire g744_n;
  wire g745_p;
  wire g745_n;
  wire g746_p;
  wire g746_n;
  wire g747_p;
  wire g747_n;
  wire g748_p;
  wire g748_n;
  wire g749_p;
  wire g749_n;
  wire g750_p;
  wire g750_n;
  wire g751_p;
  wire g751_n;
  wire g752_p;
  wire g752_n;
  wire g753_p;
  wire g753_n;
  wire g754_p;
  wire g754_n;
  wire g755_p;
  wire g755_n;
  wire g756_p;
  wire g756_n;
  wire g757_p;
  wire g757_n;
  wire g758_p;
  wire g758_n;
  wire g759_p;
  wire g759_n;
  wire g760_p;
  wire g760_n;
  wire g761_p;
  wire g761_n;
  wire g762_p;
  wire g762_n;
  wire g763_p;
  wire g763_n;
  wire g764_p;
  wire g764_n;
  wire g765_p;
  wire g765_n;
  wire g766_p;
  wire g766_n;
  wire g767_p;
  wire g767_n;
  wire g768_p;
  wire g768_n;
  wire g769_p;
  wire g769_n;
  wire g770_p;
  wire g770_n;
  wire g771_p;
  wire g771_n;
  wire g772_p;
  wire g772_n;
  wire g773_p;
  wire g773_n;
  wire g774_p;
  wire g774_n;
  wire g775_p;
  wire g775_n;
  wire g776_p;
  wire g776_n;
  wire g777_p;
  wire g777_n;
  wire g778_p;
  wire g778_n;
  wire g779_p;
  wire g779_n;
  wire g780_p;
  wire g780_n;
  wire g781_p;
  wire g781_n;
  wire g782_p;
  wire g782_n;
  wire g783_p;
  wire g783_n;
  wire g784_p;
  wire g784_n;
  wire g785_p;
  wire g785_n;
  wire g786_p;
  wire g786_n;
  wire g787_p;
  wire g787_n;
  wire g788_p;
  wire g788_n;
  wire g789_p;
  wire g789_n;
  wire g790_p;
  wire g790_n;
  wire g791_p;
  wire g791_n;
  wire g792_p;
  wire g792_n;
  wire g793_p;
  wire g793_n;
  wire g794_p;
  wire g794_n;
  wire g795_p;
  wire g795_n;
  wire g796_p;
  wire g796_n;
  wire g797_p;
  wire g797_n;
  wire g798_p;
  wire g798_n;
  wire g799_p;
  wire g799_n;
  wire g800_p;
  wire g800_n;
  wire g801_p;
  wire g801_n;
  wire g802_p;
  wire g802_n;
  wire g803_p;
  wire g803_n;
  wire g804_p;
  wire g804_n;
  wire g805_p;
  wire g805_n;
  wire g806_p;
  wire g806_n;
  wire g807_p;
  wire g807_n;
  wire g808_p;
  wire g808_n;
  wire g809_p;
  wire g809_n;
  wire g810_p;
  wire g810_n;
  wire g811_p;
  wire g811_n;
  wire g812_p;
  wire g812_n;
  wire g813_p;
  wire g813_n;
  wire g814_p;
  wire g814_n;
  wire g815_p;
  wire g815_n;
  wire g816_p;
  wire g816_n;
  wire g817_p;
  wire g817_n;
  wire g818_p;
  wire g818_n;
  wire g819_p;
  wire g819_n;
  wire g820_p;
  wire g820_n;
  wire g821_p;
  wire g821_n;
  wire g822_p;
  wire g822_n;
  wire g823_p;
  wire g823_n;
  wire g824_p;
  wire g824_n;
  wire g825_p;
  wire g825_n;
  wire g826_p;
  wire g826_n;
  wire g827_p;
  wire g827_n;
  wire g828_p;
  wire g828_n;
  wire g829_p;
  wire g829_n;
  wire g830_p;
  wire g830_n;
  wire g831_p;
  wire g831_n;
  wire g832_p;
  wire g832_n;
  wire g833_p;
  wire g833_n;
  wire g834_p;
  wire g834_n;
  wire g835_p;
  wire g835_n;
  wire g836_p;
  wire g836_n;
  wire g837_p;
  wire g837_n;
  wire g838_p;
  wire g838_n;
  wire g839_p;
  wire g839_n;
  wire g840_p;
  wire g840_n;
  wire g841_p;
  wire g841_n;
  wire g842_p;
  wire g842_n;
  wire g843_p;
  wire g843_n;
  wire g844_p;
  wire g844_n;
  wire g845_p;
  wire g845_n;
  wire g846_p;
  wire g846_n;
  wire g847_p;
  wire g847_n;
  wire g848_p;
  wire g848_n;
  wire g849_p;
  wire g849_n;
  wire g850_p;
  wire g850_n;
  wire g851_p;
  wire g851_n;
  wire g852_p;
  wire g852_n;
  wire g853_p;
  wire g853_n;
  wire g854_p;
  wire g854_n;
  wire g855_p;
  wire g855_n;
  wire g856_p;
  wire g856_n;
  wire g857_p;
  wire g857_n;
  wire g858_p;
  wire g858_n;
  wire g859_p;
  wire g859_n;
  wire g860_p;
  wire g860_n;
  wire g861_p;
  wire g861_n;
  wire g862_p;
  wire g862_n;
  wire g863_p;
  wire g863_n;
  wire g864_p;
  wire g864_n;
  wire g865_p;
  wire g865_n;
  wire g866_p;
  wire g866_n;
  wire g867_p;
  wire g867_n;
  wire g868_p;
  wire g868_n;
  wire g869_p;
  wire g869_n;
  wire g870_p;
  wire g870_n;
  wire g871_p;
  wire g871_n;
  wire g872_p;
  wire g872_n;
  wire g873_p;
  wire g873_n;
  wire g874_p;
  wire g874_n;
  wire g875_p;
  wire g875_n;
  wire g876_p;
  wire g876_n;
  wire g877_p;
  wire g877_n;
  wire g878_p;
  wire g878_n;
  wire g879_p;
  wire g879_n;
  wire g880_p;
  wire g880_n;
  wire g881_p;
  wire g881_n;
  wire g882_p;
  wire g882_n;
  wire g883_p;
  wire g883_n;
  wire g884_p;
  wire g884_n;
  wire g885_p;
  wire g885_n;
  wire g886_p;
  wire g886_n;
  wire g887_p;
  wire g887_n;
  wire g888_p;
  wire g888_n;
  wire g889_p;
  wire g889_n;
  wire g890_p;
  wire g890_n;
  wire g891_p;
  wire g891_n;
  wire g892_p;
  wire g892_n;
  wire g893_p;
  wire g893_n;
  wire g894_p;
  wire g894_n;
  wire g895_p;
  wire g895_n;
  wire g896_p;
  wire g896_n;
  wire g897_p;
  wire g897_n;
  wire g898_p;
  wire g898_n;
  wire g899_p;
  wire g899_n;
  wire g900_p;
  wire g900_n;
  wire g901_p;
  wire g901_n;
  wire g902_p;
  wire g902_n;
  wire g903_p;
  wire g903_n;
  wire g904_p;
  wire g904_n;
  wire g905_p;
  wire g905_n;
  wire g906_p;
  wire g906_n;
  wire g907_p;
  wire g907_n;
  wire g908_p;
  wire g908_n;
  wire g909_p;
  wire g909_n;
  wire g910_p;
  wire g910_n;
  wire g911_p;
  wire g911_n;
  wire g912_p;
  wire g912_n;
  wire g913_p;
  wire g913_n;
  wire g914_p;
  wire g914_n;
  wire g915_p;
  wire g915_n;
  wire g916_p;
  wire g916_n;
  wire g917_p;
  wire g917_n;
  wire g918_p;
  wire g918_n;
  wire g919_p;
  wire g919_n;
  wire g920_p;
  wire g920_n;
  wire g921_p;
  wire g921_n;
  wire g922_p;
  wire g922_n;
  wire g923_p;
  wire g923_n;
  wire g924_p;
  wire g924_n;
  wire g925_p;
  wire g925_n;
  wire g926_p;
  wire g926_n;
  wire g927_p;
  wire g927_n;
  wire g928_p;
  wire g928_n;
  wire g929_p;
  wire g929_n;
  wire g930_p;
  wire g930_n;
  wire g931_p;
  wire g931_n;
  wire g932_p;
  wire g932_n;
  wire g933_p;
  wire g933_n;
  wire g934_p;
  wire g934_n;
  wire g935_p;
  wire g935_n;
  wire g936_p;
  wire g936_n;
  wire g937_p;
  wire g937_n;
  wire g938_p;
  wire g938_n;
  wire g939_p;
  wire g939_n;
  wire g940_p;
  wire g940_n;
  wire g941_p;
  wire g941_n;
  wire g942_p;
  wire g942_n;
  wire g943_p;
  wire g943_n;
  wire g944_p;
  wire g944_n;
  wire g945_p;
  wire g945_n;
  wire g946_p;
  wire g946_n;
  wire g947_p;
  wire g947_n;
  wire g948_p;
  wire g948_n;
  wire g949_p;
  wire g949_n;
  wire g950_p;
  wire g950_n;
  wire g951_p;
  wire g951_n;
  wire g952_p;
  wire g952_n;
  wire g953_p;
  wire g953_n;
  wire g954_p;
  wire g954_n;
  wire g955_p;
  wire g955_n;
  wire g956_p;
  wire g956_n;
  wire g957_p;
  wire g957_n;
  wire g958_p;
  wire g958_n;
  wire g959_p;
  wire g959_n;
  wire g960_p;
  wire g960_n;
  wire g961_p;
  wire g961_n;
  wire g962_p;
  wire g962_n;
  wire g963_p;
  wire g963_n;
  wire g964_p;
  wire g964_n;
  wire g965_p;
  wire g965_n;
  wire g966_p;
  wire g966_n;
  wire g967_p;
  wire g967_n;
  wire g968_p;
  wire g968_n;
  wire g969_p;
  wire g969_n;
  wire g970_p;
  wire g970_n;
  wire g971_p;
  wire g971_n;
  wire g972_p;
  wire g972_n;
  wire g973_p;
  wire g973_n;
  wire g974_p;
  wire g974_n;
  wire g975_p;
  wire g975_n;
  wire g976_p;
  wire g976_n;
  wire g977_p;
  wire g977_n;
  wire g978_p;
  wire g978_n;
  wire g979_p;
  wire g979_n;
  wire g980_p;
  wire g980_n;
  wire g981_p;
  wire g981_n;
  wire g982_p;
  wire g982_n;
  wire g983_p;
  wire g983_n;
  wire g984_p;
  wire g984_n;
  wire g985_p;
  wire g985_n;
  wire g986_p;
  wire g986_n;
  wire g987_p;
  wire g987_n;
  wire g988_p;
  wire g988_n;
  wire g989_p;
  wire g989_n;
  wire g990_p;
  wire g990_n;
  wire g991_p;
  wire g991_n;
  wire g992_p;
  wire g992_n;
  wire g993_p;
  wire g993_n;
  wire g994_p;
  wire g994_n;
  wire g995_p;
  wire g995_n;
  wire g996_p;
  wire g996_n;
  wire g997_p;
  wire g997_n;
  wire g998_p;
  wire g998_n;
  wire g999_p;
  wire g999_n;
  wire g1000_p;
  wire g1000_n;
  wire g1001_p;
  wire g1001_n;
  wire g1002_p;
  wire g1002_n;
  wire g1003_p;
  wire g1003_n;
  wire g1004_p;
  wire g1004_n;
  wire g1005_p;
  wire g1005_n;
  wire g1006_p;
  wire g1006_n;
  wire g1007_p;
  wire g1007_n;
  wire g1008_p;
  wire g1008_n;
  wire g1009_p;
  wire g1009_n;
  wire g1010_p;
  wire g1010_n;
  wire g1011_p;
  wire g1011_n;
  wire g1012_p;
  wire g1012_n;
  wire g1013_p;
  wire g1013_n;
  wire g1014_p;
  wire g1014_n;
  wire g1015_p;
  wire g1015_n;
  wire g1016_p;
  wire g1016_n;
  wire g1017_p;
  wire g1017_n;
  wire g1018_p;
  wire g1018_n;
  wire g1019_p;
  wire g1019_n;
  wire g1020_p;
  wire g1020_n;
  wire g1021_p;
  wire g1021_n;
  wire g1022_p;
  wire g1022_n;
  wire g1023_p;
  wire g1023_n;
  wire g1024_p;
  wire g1024_n;
  wire g1025_p;
  wire g1025_n;
  wire g1026_p;
  wire g1026_n;
  wire g1027_p;
  wire g1027_n;
  wire g1028_p;
  wire g1028_n;
  wire g1029_p;
  wire g1029_n;
  wire g1030_p;
  wire g1030_n;
  wire g1031_p;
  wire g1031_n;
  wire g1032_p;
  wire g1032_n;
  wire g1033_p;
  wire g1033_n;
  wire g1034_p;
  wire g1034_n;
  wire g1035_p;
  wire g1035_n;
  wire g1036_p;
  wire g1036_n;
  wire g1037_p;
  wire g1037_n;
  wire g1038_p;
  wire g1038_n;
  wire g1039_p;
  wire g1039_n;
  wire g1040_p;
  wire g1040_n;
  wire g1041_p;
  wire g1041_n;
  wire g1042_p;
  wire g1042_n;
  wire g1043_p;
  wire g1043_n;
  wire g1044_p;
  wire g1044_n;
  wire g1045_p;
  wire g1045_n;
  wire g1046_p;
  wire g1046_n;
  wire g1047_p;
  wire g1047_n;
  wire g1048_p;
  wire g1048_n;
  wire g1049_p;
  wire g1049_n;
  wire g1050_p;
  wire g1050_n;
  wire g1051_p;
  wire g1051_n;
  wire g1052_p;
  wire g1052_n;
  wire g1053_p;
  wire g1053_n;
  wire g1054_p;
  wire g1054_n;
  wire g1055_p;
  wire g1055_n;
  wire g1056_p;
  wire g1056_n;
  wire g1057_p;
  wire g1057_n;
  wire g1058_p;
  wire g1058_n;
  wire g1059_p;
  wire g1059_n;
  wire g1060_p;
  wire g1060_n;
  wire g1061_p;
  wire g1061_n;
  wire g1062_p;
  wire g1062_n;
  wire g1063_p;
  wire g1063_n;
  wire g1064_p;
  wire g1064_n;
  wire g1065_p;
  wire g1065_n;
  wire g1066_p;
  wire g1066_n;
  wire g1067_p;
  wire g1067_n;
  wire g1068_p;
  wire g1068_n;
  wire g1069_p;
  wire g1069_n;
  wire g1070_p;
  wire g1070_n;
  wire g1071_p;
  wire g1071_n;
  wire g1072_p;
  wire g1072_n;
  wire g1073_p;
  wire g1073_n;
  wire g1074_p;
  wire g1074_n;
  wire g1075_p;
  wire g1075_n;
  wire g1076_p;
  wire g1076_n;
  wire g1077_p;
  wire g1077_n;
  wire g1078_p;
  wire g1078_n;
  wire g1079_p;
  wire g1079_n;
  wire g1080_p;
  wire g1080_n;
  wire g1081_p;
  wire g1081_n;
  wire g1082_p;
  wire g1082_n;
  wire g1083_p;
  wire g1083_n;
  wire g1084_p;
  wire g1084_n;
  wire g1085_p;
  wire g1085_n;
  wire g1086_p;
  wire g1086_n;
  wire g1087_p;
  wire g1087_n;
  wire g1088_p;
  wire g1088_n;
  wire g1089_p;
  wire g1089_n;
  wire g1090_p;
  wire g1090_n;
  wire g1091_p;
  wire g1091_n;
  wire g1092_p;
  wire g1092_n;
  wire g1093_p;
  wire g1093_n;
  wire g1094_p;
  wire g1094_n;
  wire g1095_p;
  wire g1095_n;
  wire g1096_p;
  wire g1096_n;
  wire g1097_p;
  wire g1097_n;
  wire g1098_p;
  wire g1098_n;
  wire g1099_p;
  wire g1099_n;
  wire g1100_p;
  wire g1100_n;
  wire g1101_p;
  wire g1101_n;
  wire g1102_p;
  wire g1102_n;
  wire g1103_p;
  wire g1103_n;
  wire g1104_p;
  wire g1104_n;
  wire g1105_p;
  wire g1105_n;
  wire g1106_p;
  wire g1106_n;
  wire g1107_p;
  wire g1107_n;
  wire g1108_p;
  wire g1108_n;
  wire g1109_p;
  wire g1109_n;
  wire g1110_p;
  wire g1110_n;
  wire g1111_p;
  wire g1111_n;
  wire g1112_p;
  wire g1112_n;
  wire g1113_p;
  wire g1113_n;
  wire g1114_p;
  wire g1114_n;
  wire g1115_p;
  wire g1115_n;
  wire g1116_p;
  wire g1116_n;
  wire g1117_p;
  wire g1117_n;
  wire g1118_p;
  wire g1118_n;
  wire g1119_p;
  wire g1119_n;
  wire g1120_p;
  wire g1120_n;
  wire g1121_p;
  wire g1121_n;
  wire g1122_p;
  wire g1122_n;
  wire g1123_p;
  wire g1123_n;
  wire g1124_p;
  wire g1124_n;
  wire g1125_p;
  wire g1125_n;
  wire g1126_p;
  wire g1126_n;
  wire g1127_p;
  wire g1127_n;
  wire g1128_p;
  wire g1128_n;
  wire g1129_p;
  wire g1129_n;
  wire g1130_p;
  wire g1130_n;
  wire g1131_p;
  wire g1131_n;
  wire g1132_p;
  wire g1132_n;
  wire g1133_p;
  wire g1133_n;
  wire g1134_p;
  wire g1134_n;
  wire g1135_p;
  wire g1135_n;
  wire g1136_p;
  wire g1136_n;
  wire g1137_p;
  wire g1137_n;
  wire g1138_p;
  wire g1138_n;
  wire g1139_p;
  wire g1139_n;
  wire g1140_p;
  wire g1140_n;
  wire g1141_p;
  wire g1141_n;
  wire g1142_p;
  wire g1142_n;
  wire g1143_p;
  wire g1143_n;
  wire g1144_p;
  wire g1144_n;
  wire g1145_p;
  wire g1145_n;
  wire g1146_p;
  wire g1146_n;
  wire g1147_p;
  wire g1147_n;
  wire g1148_p;
  wire g1148_n;
  wire g1149_p;
  wire g1149_n;
  wire g1150_p;
  wire g1150_n;
  wire g1151_p;
  wire g1151_n;
  wire g1152_p;
  wire g1152_n;
  wire g1153_p;
  wire g1153_n;
  wire g1154_p;
  wire g1154_n;
  wire g1155_p;
  wire g1155_n;
  wire g1156_p;
  wire g1156_n;
  wire g1157_p;
  wire g1157_n;
  wire g1158_p;
  wire g1158_n;
  wire g1159_p;
  wire g1159_n;
  wire g1160_p;
  wire g1160_n;
  wire g1161_p;
  wire g1161_n;
  wire g1162_p;
  wire g1162_n;
  wire g1163_p;
  wire g1163_n;
  wire g1164_p;
  wire g1164_n;
  wire g1165_p;
  wire g1165_n;
  wire g1166_p;
  wire g1166_n;
  wire g1167_p;
  wire g1167_n;
  wire g1168_p;
  wire g1168_n;
  wire g1169_p;
  wire g1169_n;
  wire g1170_p;
  wire g1170_n;
  wire g1171_p;
  wire g1171_n;
  wire g1172_p;
  wire g1172_n;
  wire g1173_p;
  wire g1173_n;
  wire g1174_p;
  wire g1174_n;
  wire g1175_p;
  wire g1175_n;
  wire g1176_p;
  wire g1176_n;
  wire g1177_p;
  wire g1177_n;
  wire g1178_p;
  wire g1178_n;
  wire g1179_p;
  wire g1179_n;
  wire g1180_p;
  wire g1180_n;
  wire g1181_p;
  wire g1181_n;
  wire g1182_p;
  wire g1182_n;
  wire g1183_p;
  wire g1183_n;
  wire g1184_p;
  wire g1184_n;
  wire g1185_p;
  wire g1185_n;
  wire g1186_p;
  wire g1186_n;
  wire g1187_p;
  wire g1187_n;
  wire g1188_p;
  wire g1188_n;
  wire g1189_p;
  wire g1189_n;
  wire g1190_p;
  wire g1190_n;
  wire g1191_p;
  wire g1191_n;
  wire g1192_p;
  wire g1192_n;
  wire g1193_p;
  wire g1193_n;
  wire g1194_p;
  wire g1194_n;
  wire g1195_p;
  wire g1195_n;
  wire g1196_p;
  wire g1196_n;
  wire g1197_p;
  wire g1197_n;
  wire g1198_p;
  wire g1198_n;
  wire g1199_p;
  wire g1199_n;
  wire g1200_p;
  wire g1200_n;
  wire g1201_p;
  wire g1201_n;
  wire g1202_p;
  wire g1202_n;
  wire g1203_p;
  wire g1203_n;
  wire g1204_p;
  wire g1204_n;
  wire g1205_p;
  wire g1205_n;
  wire g1206_p;
  wire g1206_n;
  wire g1207_p;
  wire g1207_n;
  wire g1208_p;
  wire g1208_n;
  wire g1209_p;
  wire g1209_n;
  wire g1210_p;
  wire g1210_n;
  wire g1211_p;
  wire g1211_n;
  wire g1212_p;
  wire g1212_n;
  wire g1213_p;
  wire g1213_n;
  wire g1214_p;
  wire g1214_n;
  wire g1215_p;
  wire g1215_n;
  wire g1216_p;
  wire g1216_n;
  wire g1217_p;
  wire g1217_n;
  wire g1218_p;
  wire g1218_n;
  wire g1219_p;
  wire g1219_n;
  wire g1220_p;
  wire g1220_n;
  wire g1221_p;
  wire g1221_n;
  wire g1222_p;
  wire g1222_n;
  wire g1223_p;
  wire g1223_n;
  wire g1224_p;
  wire g1224_n;
  wire g1225_p;
  wire g1225_n;
  wire g1226_p;
  wire g1226_n;
  wire g1227_p;
  wire g1227_n;
  wire g1228_p;
  wire g1228_n;
  wire g1229_p;
  wire g1229_n;
  wire g1230_p;
  wire g1230_n;
  wire g1231_p;
  wire g1231_n;
  wire g1232_p;
  wire g1232_n;
  wire g1233_p;
  wire g1233_n;
  wire g1234_p;
  wire g1234_n;
  wire g1235_p;
  wire g1235_n;
  wire g1236_p;
  wire g1236_n;
  wire g1237_p;
  wire g1237_n;
  wire g1238_p;
  wire g1238_n;
  wire g1239_p;
  wire g1239_n;
  wire g1240_p;
  wire g1240_n;
  wire g1241_p;
  wire g1241_n;
  wire g1242_p;
  wire g1242_n;
  wire g1243_p;
  wire g1243_n;
  wire g1244_p;
  wire g1244_n;
  wire g1245_p;
  wire g1245_n;
  wire g1246_p;
  wire g1246_n;
  wire g1247_p;
  wire g1247_n;
  wire g1248_p;
  wire g1248_n;
  wire g1249_p;
  wire g1249_n;
  wire g1250_p;
  wire g1250_n;
  wire g1251_p;
  wire g1251_n;
  wire g1252_p;
  wire g1252_n;
  wire g1253_p;
  wire g1253_n;
  wire g1254_p;
  wire g1254_n;
  wire g1255_p;
  wire g1255_n;
  wire g1256_p;
  wire g1256_n;
  wire g1257_p;
  wire g1257_n;
  wire g1258_p;
  wire g1258_n;
  wire g1259_p;
  wire g1259_n;
  wire g1260_p;
  wire g1260_n;
  wire g1261_p;
  wire g1261_n;
  wire g1262_p;
  wire g1262_n;
  wire g1263_p;
  wire g1263_n;
  wire g1264_p;
  wire g1264_n;
  wire g1265_p;
  wire g1265_n;
  wire g1266_p;
  wire g1266_n;
  wire g1267_p;
  wire g1267_n;
  wire g1268_p;
  wire g1268_n;
  wire g1269_p;
  wire g1269_n;
  wire g1270_p;
  wire g1270_n;
  wire g1271_p;
  wire g1271_n;
  wire g1272_p;
  wire g1272_n;
  wire g1273_p;
  wire g1273_n;
  wire g1274_p;
  wire g1274_n;
  wire g1275_p;
  wire g1275_n;
  wire g1276_p;
  wire g1276_n;
  wire g1277_p;
  wire g1277_n;
  wire g1278_p;
  wire g1278_n;
  wire g1279_p;
  wire g1279_n;
  wire g1280_p;
  wire g1280_n;
  wire g1281_p;
  wire g1281_n;
  wire g1282_p;
  wire g1282_n;
  wire g1283_p;
  wire g1283_n;
  wire g1284_p;
  wire g1284_n;
  wire g1285_p;
  wire g1285_n;
  wire g1286_p;
  wire g1286_n;
  wire g1287_p;
  wire g1287_n;
  wire g1288_p;
  wire g1288_n;
  wire g1289_p;
  wire g1289_n;
  wire g1290_p;
  wire g1290_n;
  wire g1291_p;
  wire g1291_n;
  wire g1292_p;
  wire g1292_n;
  wire g1293_p;
  wire g1293_n;
  wire g1294_p;
  wire g1294_n;
  wire g1295_p;
  wire g1295_n;
  wire g1296_p;
  wire g1296_n;
  wire g1297_p;
  wire g1297_n;
  wire g1298_p;
  wire g1298_n;
  wire g1299_p;
  wire g1299_n;
  wire g1300_p;
  wire g1300_n;
  wire g1301_p;
  wire g1301_n;
  wire g1302_p;
  wire g1302_n;
  wire g1303_p;
  wire g1303_n;
  wire g1304_p;
  wire g1304_n;
  wire g1305_p;
  wire g1305_n;
  wire g1306_p;
  wire g1306_n;
  wire g1307_p;
  wire g1307_n;
  wire g1308_p;
  wire g1308_n;
  wire g1309_p;
  wire g1309_n;
  wire g1310_p;
  wire g1310_n;
  wire g1311_p;
  wire g1311_n;
  wire g1312_p;
  wire g1312_n;
  wire g1313_p;
  wire g1313_n;
  wire g1314_p;
  wire g1314_n;
  wire g1315_p;
  wire g1315_n;
  wire g1316_p;
  wire g1316_n;
  wire g1317_p;
  wire g1317_n;
  wire g1318_p;
  wire g1318_n;
  wire g1319_p;
  wire g1319_n;
  wire g1320_p;
  wire g1320_n;
  wire g1321_p;
  wire g1321_n;
  wire g1322_p;
  wire g1322_n;
  wire g1323_p;
  wire g1323_n;
  wire g1324_p;
  wire g1324_n;
  wire g1325_p;
  wire g1325_n;
  wire g1326_p;
  wire g1326_n;
  wire g1327_p;
  wire g1327_n;
  wire g1328_p;
  wire g1328_n;
  wire g1329_p;
  wire g1329_n;
  wire g1330_p;
  wire g1330_n;
  wire g1331_p;
  wire g1331_n;
  wire g1332_p;
  wire g1332_n;
  wire g1333_p;
  wire g1333_n;
  wire g1334_p;
  wire g1334_n;
  wire g1335_p;
  wire g1335_n;
  wire g1336_p;
  wire g1336_n;
  wire g1337_p;
  wire g1337_n;
  wire g1338_p;
  wire g1338_n;
  wire g1339_p;
  wire g1339_n;
  wire g1340_p;
  wire g1340_n;
  wire g1341_p;
  wire g1341_n;
  wire g1342_p;
  wire g1342_n;
  wire g1343_p;
  wire g1343_n;
  wire g1344_p;
  wire g1344_n;
  wire g1345_p;
  wire g1345_n;
  wire g1346_p;
  wire g1346_n;
  wire g1347_p;
  wire g1347_n;
  wire g1348_p;
  wire g1348_n;
  wire g1349_p;
  wire g1349_n;
  wire g1350_p;
  wire g1350_n;
  wire g1351_p;
  wire g1351_n;
  wire g1352_p;
  wire g1352_n;
  wire g1353_p;
  wire g1353_n;
  wire g1354_p;
  wire g1354_n;
  wire g1355_p;
  wire g1355_n;
  wire g1356_p;
  wire g1356_n;
  wire g1357_p;
  wire g1357_n;
  wire g1358_p;
  wire g1358_n;
  wire g1359_p;
  wire g1359_n;
  wire g1360_p;
  wire g1360_n;
  wire g1361_p;
  wire g1361_n;
  wire g1362_p;
  wire g1362_n;
  wire g1363_p;
  wire g1363_n;
  wire g1364_p;
  wire g1364_n;
  wire g1365_p;
  wire g1365_n;
  wire g1366_p;
  wire g1366_n;
  wire g1367_p;
  wire g1367_n;
  wire g1368_p;
  wire g1368_n;
  wire g1369_p;
  wire g1369_n;
  wire g1370_p;
  wire g1370_n;
  wire g1371_p;
  wire g1371_n;
  wire g1372_p;
  wire g1372_n;
  wire g1373_p;
  wire g1373_n;
  wire g1374_p;
  wire g1374_n;
  wire g1375_p;
  wire g1375_n;
  wire g1376_p;
  wire g1376_n;
  wire g1377_p;
  wire g1377_n;
  wire g1378_p;
  wire g1378_n;
  wire g1379_p;
  wire g1379_n;
  wire g1380_p;
  wire g1380_n;
  wire g1381_p;
  wire g1381_n;
  wire g1382_p;
  wire g1382_n;
  wire g1383_p;
  wire g1383_n;
  wire g1384_p;
  wire g1384_n;
  wire g1385_p;
  wire g1385_n;
  wire g1386_p;
  wire g1386_n;
  wire g1387_p;
  wire g1387_n;
  wire g1388_p;
  wire g1388_n;
  wire g1389_p;
  wire g1389_n;
  wire g1390_p;
  wire g1390_n;
  wire g1391_p;
  wire g1391_n;
  wire g1392_p;
  wire g1392_n;
  wire g1393_p;
  wire g1393_n;
  wire g1394_p;
  wire g1394_n;
  wire g1395_p;
  wire g1395_n;
  wire g1396_p;
  wire g1396_n;
  wire g1397_p;
  wire g1397_n;
  wire g1398_p;
  wire g1398_n;
  wire g1399_p;
  wire g1399_n;
  wire g1400_p;
  wire g1400_n;
  wire g1401_p;
  wire g1401_n;
  wire g1402_p;
  wire g1402_n;
  wire g1403_p;
  wire g1403_n;
  wire g1404_p;
  wire g1404_n;
  wire g1405_p;
  wire g1405_n;
  wire g1406_p;
  wire g1406_n;
  wire g1407_p;
  wire g1407_n;
  wire g1408_p;
  wire g1408_n;
  wire g1409_p;
  wire g1409_n;
  wire g1410_p;
  wire g1410_n;
  wire g1411_p;
  wire g1411_n;
  wire g1412_p;
  wire g1412_n;
  wire g1413_p;
  wire g1413_n;
  wire g1414_p;
  wire g1414_n;
  wire g1415_p;
  wire g1415_n;
  wire g1416_p;
  wire g1416_n;
  wire g1417_p;
  wire g1417_n;
  wire g1418_p;
  wire g1418_n;
  wire g1419_p;
  wire g1419_n;
  wire g1420_p;
  wire g1420_n;
  wire g1421_p;
  wire g1421_n;
  wire g1422_p;
  wire g1422_n;
  wire g1423_p;
  wire g1423_n;
  wire g1424_p;
  wire g1424_n;
  wire g1425_p;
  wire g1425_n;
  wire g1426_p;
  wire g1426_n;
  wire g1427_p;
  wire g1427_n;
  wire g1428_p;
  wire g1428_n;
  wire g1429_p;
  wire g1429_n;
  wire g1430_p;
  wire g1430_n;
  wire g1431_p;
  wire g1431_n;
  wire g1432_p;
  wire g1432_n;
  wire g1433_p;
  wire g1433_n;
  wire g1434_p;
  wire g1434_n;
  wire g1435_p;
  wire g1435_n;
  wire g1436_p;
  wire g1436_n;
  wire g1437_p;
  wire g1437_n;
  wire g1438_p;
  wire g1438_n;
  wire g1439_p;
  wire g1439_n;
  wire g1440_p;
  wire g1440_n;
  wire g1441_p;
  wire g1441_n;
  wire g1442_p;
  wire g1442_n;
  wire g1443_p;
  wire g1443_n;
  wire g1444_p;
  wire g1444_n;
  wire g1445_p;
  wire g1445_n;
  wire g1446_p;
  wire g1446_n;
  wire g1447_p;
  wire g1447_n;
  wire g1448_p;
  wire g1448_n;
  wire g1449_p;
  wire g1449_n;
  wire g1450_p;
  wire g1450_n;
  wire g1451_p;
  wire g1451_n;
  wire g1452_p;
  wire g1452_n;
  wire g1453_p;
  wire g1453_n;
  wire g1454_p;
  wire g1454_n;
  wire g1455_p;
  wire g1455_n;
  wire g1456_p;
  wire g1456_n;
  wire g1457_p;
  wire g1457_n;
  wire g1458_p;
  wire g1458_n;
  wire g1459_p;
  wire g1459_n;
  wire g1460_p;
  wire g1460_n;
  wire g1461_p;
  wire g1461_n;
  wire g1462_p;
  wire g1462_n;
  wire g1463_p;
  wire g1463_n;
  wire g1464_p;
  wire g1464_n;
  wire g1465_p;
  wire g1465_n;
  wire g1466_p;
  wire g1466_n;
  wire g1467_p;
  wire g1467_n;
  wire g1468_p;
  wire g1468_n;
  wire g1469_p;
  wire g1469_n;
  wire g1470_p;
  wire g1470_n;
  wire g1471_p;
  wire g1471_n;
  wire g1472_p;
  wire g1472_n;
  wire g1473_p;
  wire g1473_n;
  wire g1474_p;
  wire g1474_n;
  wire g1475_p;
  wire g1475_n;
  wire g1476_p;
  wire g1476_n;
  wire g1477_p;
  wire g1477_n;
  wire g1478_p;
  wire g1478_n;
  wire g1479_p;
  wire g1479_n;
  wire g1480_p;
  wire g1480_n;
  wire g1481_p;
  wire g1481_n;
  wire g1482_p;
  wire g1482_n;
  wire g1483_p;
  wire g1483_n;
  wire g1484_p;
  wire g1484_n;
  wire g1485_p;
  wire g1485_n;
  wire g1486_p;
  wire g1486_n;
  wire g1487_p;
  wire g1487_n;
  wire g1488_p;
  wire g1488_n;
  wire g1489_p;
  wire g1489_n;
  wire g1490_p;
  wire g1490_n;
  wire g1491_p;
  wire g1491_n;
  wire g1492_p;
  wire g1492_n;
  wire g1493_p;
  wire g1493_n;
  wire g1494_p;
  wire g1494_n;
  wire g1495_p;
  wire g1495_n;
  wire g1496_p;
  wire g1496_n;
  wire g1497_p;
  wire g1497_n;
  wire g1498_p;
  wire g1498_n;
  wire g1499_p;
  wire g1499_n;
  wire g1500_p;
  wire g1500_n;
  wire g1501_p;
  wire g1501_n;
  wire g1502_p;
  wire g1502_n;
  wire g1503_p;
  wire g1503_n;
  wire g1504_p;
  wire g1504_n;
  wire g1505_p;
  wire g1505_n;
  wire g1506_p;
  wire g1506_n;
  wire g1507_p;
  wire g1507_n;
  wire g1508_p;
  wire g1508_n;
  wire g1509_p;
  wire g1509_n;
  wire g1510_p;
  wire g1510_n;
  wire g1511_p;
  wire g1511_n;
  wire g1512_p;
  wire g1512_n;
  wire g1513_p;
  wire g1513_n;
  wire g1514_p;
  wire g1514_n;
  wire g1515_p;
  wire g1515_n;
  wire g1516_p;
  wire g1516_n;
  wire g1517_p;
  wire g1517_n;
  wire g1518_p;
  wire g1518_n;
  wire g1519_p;
  wire g1519_n;
  wire g1520_p;
  wire g1520_n;
  wire g1521_p;
  wire g1521_n;
  wire g1522_p;
  wire g1522_n;
  wire g1523_p;
  wire g1523_n;
  wire g1524_p;
  wire g1524_n;
  wire g1525_p;
  wire g1525_n;
  wire g1526_p;
  wire g1526_n;
  wire g1527_p;
  wire g1527_n;
  wire g1528_p;
  wire g1528_n;
  wire g1529_p;
  wire g1529_n;
  wire g1530_p;
  wire g1530_n;
  wire g1531_p;
  wire g1531_n;
  wire g1532_p;
  wire g1532_n;
  wire g1533_p;
  wire g1533_n;
  wire g1534_p;
  wire g1534_n;
  wire g1535_p;
  wire g1535_n;
  wire g1536_p;
  wire g1536_n;
  wire g1537_p;
  wire g1537_n;
  wire g1538_p;
  wire g1538_n;
  wire g1539_p;
  wire g1539_n;
  wire g1540_p;
  wire g1540_n;
  wire g1541_p;
  wire g1541_n;
  wire g1542_p;
  wire g1542_n;
  wire g1543_p;
  wire g1543_n;
  wire g1544_p;
  wire g1544_n;
  wire g1545_p;
  wire g1545_n;
  wire G156_n_spl_;
  wire G153_n_spl_;
  wire G66_p_spl_;
  wire G66_p_spl_0;
  wire G66_p_spl_00;
  wire G66_p_spl_01;
  wire G66_p_spl_1;
  wire G1_p_spl_;
  wire G165_n_spl_;
  wire G11_n_spl_;
  wire g185_n_spl_;
  wire g185_n_spl_0;
  wire g185_n_spl_00;
  wire g185_n_spl_000;
  wire g185_n_spl_01;
  wire g185_n_spl_1;
  wire g185_n_spl_10;
  wire g185_n_spl_11;
  wire G163_n_spl_;
  wire G163_n_spl_0;
  wire G163_n_spl_00;
  wire G163_n_spl_01;
  wire G163_n_spl_1;
  wire G163_p_spl_;
  wire G163_p_spl_0;
  wire G163_p_spl_00;
  wire G163_p_spl_01;
  wire G163_p_spl_1;
  wire G168_p_spl_;
  wire G168_p_spl_0;
  wire G168_p_spl_00;
  wire G168_p_spl_000;
  wire G168_p_spl_001;
  wire G168_p_spl_01;
  wire G168_p_spl_010;
  wire G168_p_spl_1;
  wire G168_p_spl_10;
  wire G168_p_spl_11;
  wire G128_p_spl_;
  wire G128_p_spl_0;
  wire G128_p_spl_00;
  wire G128_p_spl_000;
  wire G128_p_spl_01;
  wire G128_p_spl_1;
  wire G128_p_spl_10;
  wire G128_p_spl_11;
  wire G169_p_spl_;
  wire G169_p_spl_0;
  wire G169_p_spl_00;
  wire G169_p_spl_000;
  wire G169_p_spl_001;
  wire G169_p_spl_01;
  wire G169_p_spl_010;
  wire G169_p_spl_011;
  wire G169_p_spl_1;
  wire G169_p_spl_10;
  wire G169_p_spl_11;
  wire G128_n_spl_;
  wire G128_n_spl_0;
  wire G128_n_spl_00;
  wire G128_n_spl_000;
  wire G128_n_spl_01;
  wire G128_n_spl_1;
  wire G128_n_spl_10;
  wire G128_n_spl_11;
  wire G150_p_spl_;
  wire G150_p_spl_0;
  wire G150_p_spl_00;
  wire G150_p_spl_1;
  wire G167_n_spl_;
  wire G167_n_spl_0;
  wire G167_n_spl_00;
  wire G167_n_spl_000;
  wire G167_n_spl_001;
  wire G167_n_spl_01;
  wire G167_n_spl_010;
  wire G167_n_spl_1;
  wire G167_n_spl_10;
  wire G167_n_spl_11;
  wire G166_n_spl_;
  wire G166_n_spl_0;
  wire G166_n_spl_00;
  wire G166_n_spl_000;
  wire G166_n_spl_001;
  wire G166_n_spl_01;
  wire G166_n_spl_010;
  wire G166_n_spl_011;
  wire G166_n_spl_1;
  wire G166_n_spl_10;
  wire G166_n_spl_11;
  wire G150_n_spl_;
  wire G150_n_spl_0;
  wire G150_n_spl_00;
  wire G150_n_spl_1;
  wire G126_p_spl_;
  wire G126_p_spl_0;
  wire G126_p_spl_00;
  wire G126_p_spl_000;
  wire G126_p_spl_01;
  wire G126_p_spl_1;
  wire G126_p_spl_10;
  wire G126_p_spl_11;
  wire G126_n_spl_;
  wire G126_n_spl_0;
  wire G126_n_spl_00;
  wire G126_n_spl_000;
  wire G126_n_spl_01;
  wire G126_n_spl_1;
  wire G126_n_spl_10;
  wire G126_n_spl_11;
  wire G149_p_spl_;
  wire G149_p_spl_0;
  wire G149_p_spl_00;
  wire G149_p_spl_1;
  wire G149_n_spl_;
  wire G149_n_spl_0;
  wire G149_n_spl_00;
  wire G149_n_spl_1;
  wire g233_n_spl_;
  wire g224_n_spl_;
  wire G113_p_spl_;
  wire G113_p_spl_0;
  wire G113_p_spl_00;
  wire G113_p_spl_1;
  wire G102_p_spl_;
  wire G102_p_spl_0;
  wire G102_p_spl_00;
  wire G102_p_spl_000;
  wire G102_p_spl_001;
  wire G102_p_spl_01;
  wire G102_p_spl_010;
  wire G102_p_spl_011;
  wire G102_p_spl_1;
  wire G102_p_spl_10;
  wire G102_p_spl_100;
  wire G102_p_spl_101;
  wire G102_p_spl_11;
  wire G102_p_spl_110;
  wire G113_n_spl_;
  wire G113_n_spl_0;
  wire G113_n_spl_00;
  wire G113_n_spl_01;
  wire G113_n_spl_1;
  wire G102_n_spl_;
  wire G102_n_spl_0;
  wire G102_n_spl_00;
  wire G102_n_spl_000;
  wire G102_n_spl_001;
  wire G102_n_spl_01;
  wire G102_n_spl_010;
  wire G102_n_spl_011;
  wire G102_n_spl_1;
  wire G102_n_spl_10;
  wire G102_n_spl_100;
  wire G102_n_spl_101;
  wire G102_n_spl_11;
  wire G102_n_spl_110;
  wire G98_p_spl_;
  wire G98_p_spl_0;
  wire G98_p_spl_00;
  wire G98_p_spl_000;
  wire G98_p_spl_001;
  wire G98_p_spl_01;
  wire G98_p_spl_010;
  wire G98_p_spl_011;
  wire G98_p_spl_1;
  wire G98_p_spl_10;
  wire G98_p_spl_100;
  wire G98_p_spl_101;
  wire G98_p_spl_11;
  wire G98_p_spl_110;
  wire G98_p_spl_111;
  wire G98_n_spl_;
  wire G98_n_spl_0;
  wire G98_n_spl_00;
  wire G98_n_spl_000;
  wire G98_n_spl_001;
  wire G98_n_spl_01;
  wire G98_n_spl_010;
  wire G98_n_spl_011;
  wire G98_n_spl_1;
  wire G98_n_spl_10;
  wire G98_n_spl_100;
  wire G98_n_spl_101;
  wire G98_n_spl_11;
  wire G98_n_spl_110;
  wire G98_n_spl_111;
  wire G115_p_spl_;
  wire G115_p_spl_0;
  wire G115_p_spl_00;
  wire G115_p_spl_1;
  wire G101_p_spl_;
  wire G101_p_spl_0;
  wire G101_p_spl_00;
  wire G101_p_spl_000;
  wire G101_p_spl_001;
  wire G101_p_spl_01;
  wire G101_p_spl_010;
  wire G101_p_spl_011;
  wire G101_p_spl_1;
  wire G101_p_spl_10;
  wire G101_p_spl_100;
  wire G101_p_spl_101;
  wire G101_p_spl_11;
  wire G101_p_spl_110;
  wire G101_p_spl_111;
  wire G115_n_spl_;
  wire G115_n_spl_0;
  wire G115_n_spl_00;
  wire G115_n_spl_1;
  wire G101_n_spl_;
  wire G101_n_spl_0;
  wire G101_n_spl_00;
  wire G101_n_spl_000;
  wire G101_n_spl_001;
  wire G101_n_spl_01;
  wire G101_n_spl_010;
  wire G101_n_spl_011;
  wire G101_n_spl_1;
  wire G101_n_spl_10;
  wire G101_n_spl_100;
  wire G101_n_spl_101;
  wire G101_n_spl_11;
  wire G101_n_spl_110;
  wire G101_n_spl_111;
  wire G100_p_spl_;
  wire G100_p_spl_0;
  wire G100_p_spl_00;
  wire G100_p_spl_000;
  wire G100_p_spl_0000;
  wire G100_p_spl_001;
  wire G100_p_spl_01;
  wire G100_p_spl_010;
  wire G100_p_spl_011;
  wire G100_p_spl_1;
  wire G100_p_spl_10;
  wire G100_p_spl_100;
  wire G100_p_spl_101;
  wire G100_p_spl_11;
  wire G100_p_spl_110;
  wire G100_p_spl_111;
  wire G100_n_spl_;
  wire G100_n_spl_0;
  wire G100_n_spl_00;
  wire G100_n_spl_000;
  wire G100_n_spl_0000;
  wire G100_n_spl_001;
  wire G100_n_spl_01;
  wire G100_n_spl_010;
  wire G100_n_spl_011;
  wire G100_n_spl_1;
  wire G100_n_spl_10;
  wire G100_n_spl_100;
  wire G100_n_spl_101;
  wire G100_n_spl_11;
  wire G100_n_spl_110;
  wire G100_n_spl_111;
  wire g240_p_spl_;
  wire g237_n_spl_;
  wire g237_n_spl_0;
  wire g237_n_spl_1;
  wire g240_n_spl_;
  wire g240_n_spl_0;
  wire g237_p_spl_;
  wire g241_n_spl_;
  wire G130_p_spl_;
  wire G130_p_spl_0;
  wire G130_p_spl_00;
  wire G130_p_spl_1;
  wire G130_n_spl_;
  wire G130_n_spl_0;
  wire G130_n_spl_00;
  wire G130_n_spl_1;
  wire G148_n_spl_;
  wire G148_n_spl_0;
  wire G148_n_spl_00;
  wire G148_n_spl_1;
  wire G148_p_spl_;
  wire G148_p_spl_0;
  wire G148_p_spl_00;
  wire G148_p_spl_1;
  wire g248_n_spl_;
  wire g245_n_spl_;
  wire g245_n_spl_0;
  wire g245_n_spl_1;
  wire G119_p_spl_;
  wire G119_p_spl_0;
  wire G119_p_spl_00;
  wire G119_p_spl_01;
  wire G119_p_spl_1;
  wire G119_p_spl_10;
  wire G119_n_spl_;
  wire G119_n_spl_0;
  wire G119_n_spl_00;
  wire G119_n_spl_01;
  wire G119_n_spl_1;
  wire G119_n_spl_10;
  wire G146_p_spl_;
  wire G146_p_spl_0;
  wire G146_p_spl_1;
  wire G146_n_spl_;
  wire G146_n_spl_0;
  wire G146_n_spl_1;
  wire G117_p_spl_;
  wire G117_p_spl_0;
  wire G117_p_spl_00;
  wire G117_p_spl_01;
  wire G117_p_spl_1;
  wire G117_p_spl_10;
  wire G117_n_spl_;
  wire G117_n_spl_0;
  wire G117_n_spl_00;
  wire G117_n_spl_01;
  wire G117_n_spl_1;
  wire G117_n_spl_10;
  wire G145_p_spl_;
  wire G145_p_spl_0;
  wire G145_p_spl_1;
  wire G145_n_spl_;
  wire G145_n_spl_0;
  wire G145_n_spl_1;
  wire g267_p_spl_;
  wire g258_p_spl_;
  wire g267_n_spl_;
  wire g267_n_spl_0;
  wire g258_n_spl_;
  wire g258_n_spl_0;
  wire G121_p_spl_;
  wire G121_p_spl_0;
  wire G121_p_spl_00;
  wire G121_p_spl_000;
  wire G121_p_spl_01;
  wire G121_p_spl_1;
  wire G121_p_spl_10;
  wire G121_p_spl_11;
  wire G121_n_spl_;
  wire G121_n_spl_0;
  wire G121_n_spl_00;
  wire G121_n_spl_000;
  wire G121_n_spl_01;
  wire G121_n_spl_1;
  wire G121_n_spl_10;
  wire G121_n_spl_11;
  wire G147_p_spl_;
  wire G147_p_spl_0;
  wire G147_p_spl_00;
  wire G147_p_spl_1;
  wire G147_n_spl_;
  wire G147_n_spl_0;
  wire G147_n_spl_00;
  wire G147_n_spl_1;
  wire g277_n_spl_;
  wire g268_n_spl_;
  wire G107_p_spl_;
  wire G107_p_spl_0;
  wire G107_p_spl_00;
  wire G107_p_spl_000;
  wire G107_p_spl_01;
  wire G107_p_spl_1;
  wire G107_p_spl_10;
  wire G107_p_spl_11;
  wire G107_n_spl_;
  wire G107_n_spl_0;
  wire G107_n_spl_00;
  wire G107_n_spl_000;
  wire G107_n_spl_01;
  wire G107_n_spl_1;
  wire G107_n_spl_10;
  wire G107_n_spl_11;
  wire G139_p_spl_;
  wire G139_p_spl_0;
  wire G139_p_spl_00;
  wire G139_p_spl_1;
  wire G139_n_spl_;
  wire G139_n_spl_0;
  wire G139_n_spl_00;
  wire G139_n_spl_1;
  wire G105_p_spl_;
  wire G105_p_spl_0;
  wire G105_p_spl_00;
  wire G105_p_spl_000;
  wire G105_p_spl_01;
  wire G105_p_spl_1;
  wire G105_p_spl_10;
  wire G105_p_spl_11;
  wire G105_n_spl_;
  wire G105_n_spl_0;
  wire G105_n_spl_00;
  wire G105_n_spl_000;
  wire G105_n_spl_01;
  wire G105_n_spl_1;
  wire G105_n_spl_10;
  wire G105_n_spl_11;
  wire G138_p_spl_;
  wire G138_p_spl_0;
  wire G138_p_spl_00;
  wire G138_p_spl_1;
  wire G138_n_spl_;
  wire G138_n_spl_0;
  wire G138_n_spl_00;
  wire G138_n_spl_1;
  wire g298_n_spl_;
  wire g289_n_spl_;
  wire G109_p_spl_;
  wire G109_p_spl_0;
  wire G109_p_spl_00;
  wire G109_p_spl_000;
  wire G109_p_spl_01;
  wire G109_p_spl_1;
  wire G109_p_spl_10;
  wire G109_p_spl_11;
  wire G109_n_spl_;
  wire G109_n_spl_0;
  wire G109_n_spl_00;
  wire G109_n_spl_000;
  wire G109_n_spl_01;
  wire G109_n_spl_1;
  wire G109_n_spl_10;
  wire G109_n_spl_11;
  wire G135_p_spl_;
  wire G135_p_spl_0;
  wire G135_p_spl_00;
  wire G135_p_spl_1;
  wire G135_n_spl_;
  wire G135_n_spl_0;
  wire G135_n_spl_00;
  wire G135_n_spl_1;
  wire G88_p_spl_;
  wire G88_p_spl_0;
  wire G88_p_spl_00;
  wire G88_p_spl_01;
  wire G88_p_spl_1;
  wire G88_p_spl_10;
  wire G88_n_spl_;
  wire G88_n_spl_0;
  wire G88_n_spl_00;
  wire G88_n_spl_01;
  wire G88_n_spl_1;
  wire G88_n_spl_10;
  wire G142_p_spl_;
  wire G142_p_spl_0;
  wire G142_p_spl_1;
  wire G142_n_spl_;
  wire G142_n_spl_0;
  wire G142_n_spl_1;
  wire g317_n_spl_;
  wire g317_n_spl_0;
  wire g317_n_spl_1;
  wire g308_n_spl_;
  wire G90_p_spl_;
  wire G90_p_spl_0;
  wire G90_p_spl_00;
  wire G90_p_spl_000;
  wire G90_p_spl_01;
  wire G90_p_spl_1;
  wire G90_p_spl_10;
  wire G90_p_spl_11;
  wire G90_n_spl_;
  wire G90_n_spl_0;
  wire G90_n_spl_00;
  wire G90_n_spl_000;
  wire G90_n_spl_01;
  wire G90_n_spl_1;
  wire G90_n_spl_10;
  wire G90_n_spl_11;
  wire G143_p_spl_;
  wire G143_p_spl_0;
  wire G143_p_spl_00;
  wire G143_p_spl_1;
  wire G143_n_spl_;
  wire G143_n_spl_0;
  wire G143_n_spl_00;
  wire G143_n_spl_1;
  wire G92_p_spl_;
  wire G92_p_spl_0;
  wire G92_p_spl_00;
  wire G92_p_spl_000;
  wire G92_p_spl_01;
  wire G92_p_spl_1;
  wire G92_p_spl_10;
  wire G92_p_spl_11;
  wire G92_n_spl_;
  wire G92_n_spl_0;
  wire G92_n_spl_00;
  wire G92_n_spl_000;
  wire G92_n_spl_01;
  wire G92_n_spl_1;
  wire G92_n_spl_10;
  wire G92_n_spl_11;
  wire G144_p_spl_;
  wire G144_p_spl_0;
  wire G144_p_spl_00;
  wire G144_p_spl_1;
  wire G144_n_spl_;
  wire G144_n_spl_0;
  wire G144_n_spl_00;
  wire G144_n_spl_1;
  wire g337_n_spl_;
  wire g328_n_spl_;
  wire G94_p_spl_;
  wire G94_p_spl_0;
  wire G94_p_spl_00;
  wire G94_p_spl_000;
  wire G94_p_spl_01;
  wire G94_p_spl_1;
  wire G94_p_spl_10;
  wire G94_p_spl_11;
  wire G94_n_spl_;
  wire G94_n_spl_0;
  wire G94_n_spl_00;
  wire G94_n_spl_000;
  wire G94_n_spl_01;
  wire G94_n_spl_1;
  wire G94_n_spl_10;
  wire G94_n_spl_11;
  wire G140_p_spl_;
  wire G140_p_spl_0;
  wire G140_p_spl_00;
  wire G140_p_spl_1;
  wire G140_n_spl_;
  wire G140_n_spl_0;
  wire G140_n_spl_00;
  wire G140_n_spl_1;
  wire G96_p_spl_;
  wire G96_p_spl_0;
  wire G96_p_spl_00;
  wire G96_p_spl_000;
  wire G96_p_spl_01;
  wire G96_p_spl_1;
  wire G96_p_spl_10;
  wire G96_p_spl_11;
  wire G96_n_spl_;
  wire G96_n_spl_0;
  wire G96_n_spl_00;
  wire G96_n_spl_000;
  wire G96_n_spl_01;
  wire G96_n_spl_1;
  wire G96_n_spl_10;
  wire G96_n_spl_11;
  wire G141_p_spl_;
  wire G141_p_spl_0;
  wire G141_p_spl_00;
  wire G141_p_spl_1;
  wire G141_n_spl_;
  wire G141_n_spl_0;
  wire G141_n_spl_00;
  wire G141_n_spl_1;
  wire G103_p_spl_;
  wire G103_p_spl_0;
  wire G103_p_spl_00;
  wire G103_p_spl_000;
  wire G103_p_spl_01;
  wire G103_p_spl_1;
  wire G103_p_spl_10;
  wire G103_p_spl_11;
  wire G103_n_spl_;
  wire G103_n_spl_0;
  wire G103_n_spl_00;
  wire G103_n_spl_000;
  wire G103_n_spl_01;
  wire G103_n_spl_1;
  wire G103_n_spl_10;
  wire G103_n_spl_11;
  wire G137_p_spl_;
  wire G137_p_spl_0;
  wire G137_p_spl_00;
  wire G137_p_spl_1;
  wire G137_n_spl_;
  wire G137_n_spl_0;
  wire G137_n_spl_00;
  wire G137_n_spl_1;
  wire g365_n_spl_;
  wire g356_n_spl_;
  wire g347_n_spl_;
  wire G124_n_spl_;
  wire G124_n_spl_0;
  wire G124_n_spl_00;
  wire G124_n_spl_000;
  wire G124_n_spl_0000;
  wire G124_n_spl_0001;
  wire G124_n_spl_001;
  wire G124_n_spl_0010;
  wire G124_n_spl_0011;
  wire G124_n_spl_01;
  wire G124_n_spl_010;
  wire G124_n_spl_011;
  wire G124_n_spl_1;
  wire G124_n_spl_10;
  wire G124_n_spl_100;
  wire G124_n_spl_101;
  wire G124_n_spl_11;
  wire G124_n_spl_110;
  wire G124_n_spl_111;
  wire G124_p_spl_;
  wire G124_p_spl_0;
  wire G124_p_spl_00;
  wire G124_p_spl_000;
  wire G124_p_spl_0000;
  wire G124_p_spl_0001;
  wire G124_p_spl_001;
  wire G124_p_spl_0010;
  wire G124_p_spl_0011;
  wire G124_p_spl_01;
  wire G124_p_spl_010;
  wire G124_p_spl_011;
  wire G124_p_spl_1;
  wire G124_p_spl_10;
  wire G124_p_spl_100;
  wire G124_p_spl_101;
  wire G124_p_spl_11;
  wire G124_p_spl_110;
  wire G124_p_spl_111;
  wire g372_p_spl_;
  wire g372_p_spl_0;
  wire g372_p_spl_1;
  wire g372_n_spl_;
  wire g372_n_spl_0;
  wire g372_n_spl_1;
  wire g374_n_spl_;
  wire g374_n_spl_0;
  wire g374_n_spl_1;
  wire g373_n_spl_;
  wire g373_n_spl_0;
  wire g374_p_spl_;
  wire g374_p_spl_0;
  wire g374_p_spl_1;
  wire g373_p_spl_;
  wire g373_p_spl_0;
  wire g378_p_spl_;
  wire g378_p_spl_0;
  wire g378_p_spl_1;
  wire g378_n_spl_;
  wire g378_n_spl_0;
  wire g378_n_spl_1;
  wire g380_n_spl_;
  wire g379_n_spl_;
  wire g380_p_spl_;
  wire g379_p_spl_;
  wire g381_p_spl_;
  wire g381_p_spl_0;
  wire g381_p_spl_00;
  wire g381_p_spl_01;
  wire g381_p_spl_1;
  wire g381_p_spl_10;
  wire g375_p_spl_;
  wire g375_p_spl_0;
  wire g375_p_spl_00;
  wire g375_p_spl_1;
  wire g381_n_spl_;
  wire g381_n_spl_0;
  wire g381_n_spl_00;
  wire g381_n_spl_01;
  wire g381_n_spl_1;
  wire g381_n_spl_10;
  wire g375_n_spl_;
  wire g375_n_spl_0;
  wire g375_n_spl_00;
  wire g375_n_spl_1;
  wire g385_p_spl_;
  wire g385_p_spl_0;
  wire g385_p_spl_1;
  wire g385_n_spl_;
  wire g385_n_spl_0;
  wire g385_n_spl_1;
  wire g387_n_spl_;
  wire g386_n_spl_;
  wire g387_p_spl_;
  wire g386_p_spl_;
  wire g388_p_spl_;
  wire g388_p_spl_0;
  wire g388_p_spl_00;
  wire g388_p_spl_01;
  wire g388_p_spl_1;
  wire g382_p_spl_;
  wire g388_n_spl_;
  wire g388_n_spl_0;
  wire g388_n_spl_00;
  wire g388_n_spl_01;
  wire g388_n_spl_1;
  wire g382_n_spl_;
  wire g392_p_spl_;
  wire g392_p_spl_0;
  wire g392_p_spl_1;
  wire g392_n_spl_;
  wire g392_n_spl_0;
  wire g392_n_spl_1;
  wire g393_n_spl_;
  wire g395_n_spl_;
  wire g395_n_spl_0;
  wire g395_n_spl_00;
  wire g395_n_spl_01;
  wire g395_n_spl_1;
  wire g395_n_spl_10;
  wire g389_n_spl_;
  wire g389_n_spl_0;
  wire g399_p_spl_;
  wire g399_p_spl_0;
  wire g399_p_spl_1;
  wire g399_n_spl_;
  wire g399_n_spl_0;
  wire g399_n_spl_1;
  wire g401_n_spl_;
  wire g401_n_spl_0;
  wire g400_n_spl_;
  wire g400_n_spl_0;
  wire g400_n_spl_00;
  wire g400_n_spl_1;
  wire g401_p_spl_;
  wire g401_p_spl_0;
  wire g400_p_spl_;
  wire g400_p_spl_0;
  wire g400_p_spl_00;
  wire g400_p_spl_1;
  wire g405_p_spl_;
  wire g405_p_spl_0;
  wire g405_p_spl_1;
  wire g405_n_spl_;
  wire g405_n_spl_0;
  wire g405_n_spl_1;
  wire g406_n_spl_;
  wire g406_n_spl_0;
  wire g406_p_spl_;
  wire g406_p_spl_0;
  wire g408_p_spl_;
  wire g408_p_spl_0;
  wire g408_p_spl_1;
  wire g402_p_spl_;
  wire g402_p_spl_0;
  wire g402_p_spl_1;
  wire g408_n_spl_;
  wire g408_n_spl_0;
  wire g408_n_spl_00;
  wire g408_n_spl_1;
  wire g402_n_spl_;
  wire g402_n_spl_0;
  wire g412_p_spl_;
  wire g412_p_spl_0;
  wire g412_p_spl_1;
  wire g412_n_spl_;
  wire g412_n_spl_0;
  wire g412_n_spl_1;
  wire g413_n_spl_;
  wire g413_p_spl_;
  wire g415_p_spl_;
  wire g415_p_spl_0;
  wire g415_p_spl_00;
  wire g415_p_spl_1;
  wire g409_p_spl_;
  wire g409_p_spl_0;
  wire g415_n_spl_;
  wire g415_n_spl_0;
  wire g415_n_spl_00;
  wire g415_n_spl_1;
  wire g409_n_spl_;
  wire g409_n_spl_0;
  wire g419_p_spl_;
  wire g419_p_spl_0;
  wire g419_p_spl_1;
  wire g419_n_spl_;
  wire g419_n_spl_0;
  wire g419_n_spl_1;
  wire g420_n_spl_;
  wire g420_n_spl_0;
  wire g420_p_spl_;
  wire g420_p_spl_0;
  wire g422_p_spl_;
  wire g422_p_spl_0;
  wire g422_p_spl_00;
  wire g422_p_spl_1;
  wire g416_p_spl_;
  wire g416_p_spl_0;
  wire g422_n_spl_;
  wire g422_n_spl_0;
  wire g422_n_spl_00;
  wire g422_n_spl_01;
  wire g422_n_spl_1;
  wire g416_n_spl_;
  wire g416_n_spl_0;
  wire g426_p_spl_;
  wire g426_p_spl_0;
  wire g426_p_spl_1;
  wire g426_n_spl_;
  wire g426_n_spl_0;
  wire g426_n_spl_1;
  wire g427_n_spl_;
  wire g427_p_spl_;
  wire g429_p_spl_;
  wire g429_p_spl_0;
  wire g429_p_spl_00;
  wire g429_p_spl_01;
  wire g429_p_spl_1;
  wire g429_p_spl_10;
  wire g423_p_spl_;
  wire g429_n_spl_;
  wire g429_n_spl_0;
  wire g429_n_spl_00;
  wire g429_n_spl_01;
  wire g429_n_spl_1;
  wire g429_n_spl_10;
  wire g423_n_spl_;
  wire g430_n_spl_;
  wire g430_n_spl_0;
  wire g430_n_spl_1;
  wire g396_n_spl_;
  wire G123_n_spl_;
  wire G123_n_spl_0;
  wire G123_n_spl_00;
  wire G123_n_spl_000;
  wire G123_n_spl_0000;
  wire G123_n_spl_0001;
  wire G123_n_spl_001;
  wire G123_n_spl_0010;
  wire G123_n_spl_01;
  wire G123_n_spl_010;
  wire G123_n_spl_011;
  wire G123_n_spl_1;
  wire G123_n_spl_10;
  wire G123_n_spl_100;
  wire G123_n_spl_101;
  wire G123_n_spl_11;
  wire G123_n_spl_110;
  wire G123_n_spl_111;
  wire G123_p_spl_;
  wire G123_p_spl_0;
  wire G123_p_spl_00;
  wire G123_p_spl_000;
  wire G123_p_spl_0000;
  wire G123_p_spl_0001;
  wire G123_p_spl_001;
  wire G123_p_spl_0010;
  wire G123_p_spl_01;
  wire G123_p_spl_010;
  wire G123_p_spl_011;
  wire G123_p_spl_1;
  wire G123_p_spl_10;
  wire G123_p_spl_100;
  wire G123_p_spl_101;
  wire G123_p_spl_11;
  wire G123_p_spl_110;
  wire G123_p_spl_111;
  wire g434_p_spl_;
  wire g434_p_spl_0;
  wire g434_p_spl_1;
  wire g434_n_spl_;
  wire g434_n_spl_0;
  wire g434_n_spl_1;
  wire g435_n_spl_;
  wire g435_p_spl_;
  wire g440_p_spl_;
  wire g440_p_spl_0;
  wire g440_p_spl_1;
  wire g440_n_spl_;
  wire g440_n_spl_0;
  wire g440_n_spl_1;
  wire g442_n_spl_;
  wire g442_n_spl_0;
  wire g442_n_spl_1;
  wire g441_n_spl_;
  wire g441_n_spl_0;
  wire g441_n_spl_00;
  wire g441_n_spl_1;
  wire g442_p_spl_;
  wire g442_p_spl_0;
  wire g442_p_spl_1;
  wire g441_p_spl_;
  wire g441_p_spl_0;
  wire g441_p_spl_00;
  wire g441_p_spl_1;
  wire g443_p_spl_;
  wire g443_p_spl_0;
  wire g443_p_spl_00;
  wire g443_p_spl_1;
  wire g437_p_spl_;
  wire g437_p_spl_0;
  wire g437_p_spl_00;
  wire g437_p_spl_01;
  wire g437_p_spl_1;
  wire g443_n_spl_;
  wire g443_n_spl_0;
  wire g443_n_spl_00;
  wire g443_n_spl_1;
  wire g437_n_spl_;
  wire g437_n_spl_0;
  wire g437_n_spl_00;
  wire g437_n_spl_01;
  wire g437_n_spl_1;
  wire g447_p_spl_;
  wire g447_p_spl_0;
  wire g447_p_spl_1;
  wire g447_n_spl_;
  wire g447_n_spl_0;
  wire g447_n_spl_1;
  wire g448_n_spl_;
  wire g448_p_spl_;
  wire G125_n_spl_;
  wire g451_n_spl_;
  wire g451_n_spl_0;
  wire g451_n_spl_1;
  wire g451_p_spl_;
  wire g451_p_spl_0;
  wire g451_p_spl_1;
  wire g452_n_spl_;
  wire g452_n_spl_0;
  wire g452_p_spl_;
  wire g452_p_spl_0;
  wire g454_p_spl_;
  wire g454_p_spl_0;
  wire g454_p_spl_1;
  wire g450_p_spl_;
  wire g450_p_spl_0;
  wire g450_p_spl_1;
  wire g454_n_spl_;
  wire g454_n_spl_0;
  wire g454_n_spl_00;
  wire g454_n_spl_1;
  wire g450_n_spl_;
  wire g450_n_spl_0;
  wire g450_n_spl_1;
  wire G129_n_spl_;
  wire g458_p_spl_;
  wire g458_p_spl_0;
  wire g458_p_spl_1;
  wire g458_n_spl_;
  wire g458_n_spl_0;
  wire g458_n_spl_1;
  wire g459_n_spl_;
  wire g459_n_spl_0;
  wire g459_p_spl_;
  wire g459_p_spl_0;
  wire G131_n_spl_;
  wire g464_n_spl_;
  wire g464_n_spl_0;
  wire g464_n_spl_00;
  wire g464_n_spl_01;
  wire g464_n_spl_1;
  wire g464_n_spl_10;
  wire g461_p_spl_;
  wire g461_p_spl_0;
  wire g464_p_spl_;
  wire g464_p_spl_0;
  wire g464_p_spl_00;
  wire g464_p_spl_01;
  wire g464_p_spl_1;
  wire g464_p_spl_10;
  wire g461_n_spl_;
  wire g461_n_spl_0;
  wire G127_n_spl_;
  wire g468_p_spl_;
  wire g468_p_spl_0;
  wire g468_p_spl_1;
  wire g468_n_spl_;
  wire g468_n_spl_0;
  wire g468_n_spl_1;
  wire g469_n_spl_;
  wire g469_n_spl_0;
  wire g469_p_spl_;
  wire g469_p_spl_0;
  wire g471_p_spl_;
  wire g471_p_spl_0;
  wire g471_p_spl_1;
  wire g465_p_spl_;
  wire g465_p_spl_0;
  wire g471_n_spl_;
  wire g471_n_spl_0;
  wire g471_n_spl_00;
  wire g471_n_spl_1;
  wire g465_n_spl_;
  wire g465_n_spl_0;
  wire g472_p_spl_;
  wire g455_p_spl_;
  wire g472_n_spl_;
  wire g455_n_spl_;
  wire G114_n_spl_;
  wire G114_n_spl_0;
  wire G114_p_spl_;
  wire g479_n_spl_;
  wire g479_n_spl_0;
  wire g479_n_spl_00;
  wire g479_n_spl_01;
  wire g479_n_spl_1;
  wire g479_n_spl_10;
  wire g476_n_spl_;
  wire g476_n_spl_0;
  wire g476_n_spl_1;
  wire g479_p_spl_;
  wire g479_p_spl_0;
  wire g479_p_spl_00;
  wire g479_p_spl_01;
  wire g479_p_spl_1;
  wire g479_p_spl_10;
  wire g476_p_spl_;
  wire g476_p_spl_0;
  wire g476_p_spl_00;
  wire g476_p_spl_1;
  wire g480_p_spl_;
  wire g480_p_spl_0;
  wire g473_p_spl_;
  wire g444_p_spl_;
  wire g444_p_spl_0;
  wire g488_n_spl_;
  wire g485_p_spl_;
  wire g488_p_spl_;
  wire g485_n_spl_;
  wire G132_n_spl_;
  wire G132_n_spl_0;
  wire G132_p_spl_;
  wire G132_p_spl_0;
  wire g494_n_spl_;
  wire g494_p_spl_;
  wire g500_n_spl_;
  wire g497_n_spl_;
  wire g500_p_spl_;
  wire g497_p_spl_;
  wire g512_n_spl_;
  wire g509_p_spl_;
  wire g512_p_spl_;
  wire g509_n_spl_;
  wire G111_n_spl_;
  wire G111_n_spl_0;
  wire G111_p_spl_;
  wire G111_p_spl_0;
  wire g521_n_spl_;
  wire g518_n_spl_;
  wire g521_p_spl_;
  wire g518_p_spl_;
  wire g527_n_spl_;
  wire g524_n_spl_;
  wire g527_p_spl_;
  wire g524_p_spl_;
  wire g535_n_spl_;
  wire g535_n_spl_0;
  wire g535_n_spl_1;
  wire g535_p_spl_;
  wire g535_p_spl_0;
  wire g535_p_spl_1;
  wire g537_n_spl_;
  wire g537_n_spl_0;
  wire g537_n_spl_00;
  wire g537_n_spl_1;
  wire g537_p_spl_;
  wire g537_p_spl_0;
  wire g537_p_spl_00;
  wire g537_p_spl_1;
  wire g539_n_spl_;
  wire g539_n_spl_0;
  wire g539_n_spl_1;
  wire g539_p_spl_;
  wire g539_p_spl_0;
  wire g539_p_spl_1;
  wire g541_p_spl_;
  wire g541_p_spl_0;
  wire g541_p_spl_00;
  wire g541_p_spl_1;
  wire g544_n_spl_;
  wire g544_n_spl_0;
  wire g544_n_spl_1;
  wire g544_p_spl_;
  wire g544_p_spl_0;
  wire g544_p_spl_1;
  wire g545_n_spl_;
  wire g545_p_spl_;
  wire g546_p_spl_;
  wire g546_p_spl_0;
  wire g546_p_spl_1;
  wire g553_p_spl_;
  wire G177_p_spl_;
  wire G177_p_spl_0;
  wire G177_p_spl_00;
  wire G177_p_spl_000;
  wire G177_p_spl_0000;
  wire G177_p_spl_0001;
  wire G177_p_spl_001;
  wire G177_p_spl_0010;
  wire G177_p_spl_0011;
  wire G177_p_spl_01;
  wire G177_p_spl_010;
  wire G177_p_spl_0100;
  wire G177_p_spl_0101;
  wire G177_p_spl_011;
  wire G177_p_spl_0110;
  wire G177_p_spl_0111;
  wire G177_p_spl_1;
  wire G177_p_spl_10;
  wire G177_p_spl_100;
  wire G177_p_spl_1000;
  wire G177_p_spl_1001;
  wire G177_p_spl_101;
  wire G177_p_spl_11;
  wire G177_p_spl_110;
  wire G177_p_spl_111;
  wire G176_p_spl_;
  wire G176_p_spl_0;
  wire G176_p_spl_00;
  wire G176_p_spl_000;
  wire G176_p_spl_0000;
  wire G176_p_spl_00000;
  wire G176_p_spl_00001;
  wire G176_p_spl_0001;
  wire G176_p_spl_001;
  wire G176_p_spl_0010;
  wire G176_p_spl_0011;
  wire G176_p_spl_01;
  wire G176_p_spl_010;
  wire G176_p_spl_0100;
  wire G176_p_spl_0101;
  wire G176_p_spl_011;
  wire G176_p_spl_0110;
  wire G176_p_spl_0111;
  wire G176_p_spl_1;
  wire G176_p_spl_10;
  wire G176_p_spl_100;
  wire G176_p_spl_1000;
  wire G176_p_spl_1001;
  wire G176_p_spl_101;
  wire G176_p_spl_1010;
  wire G176_p_spl_1011;
  wire G176_p_spl_11;
  wire G176_p_spl_110;
  wire G176_p_spl_1100;
  wire G176_p_spl_1101;
  wire G176_p_spl_111;
  wire G176_p_spl_1110;
  wire G176_p_spl_1111;
  wire G177_n_spl_;
  wire G177_n_spl_0;
  wire G177_n_spl_00;
  wire G177_n_spl_000;
  wire G177_n_spl_0000;
  wire G177_n_spl_0001;
  wire G177_n_spl_001;
  wire G177_n_spl_0010;
  wire G177_n_spl_0011;
  wire G177_n_spl_01;
  wire G177_n_spl_010;
  wire G177_n_spl_011;
  wire G177_n_spl_1;
  wire G177_n_spl_10;
  wire G177_n_spl_100;
  wire G177_n_spl_101;
  wire G177_n_spl_11;
  wire G177_n_spl_110;
  wire G177_n_spl_111;
  wire G176_n_spl_;
  wire G176_n_spl_0;
  wire G176_n_spl_00;
  wire G176_n_spl_000;
  wire G176_n_spl_0000;
  wire G176_n_spl_0001;
  wire G176_n_spl_001;
  wire G176_n_spl_0010;
  wire G176_n_spl_0011;
  wire G176_n_spl_01;
  wire G176_n_spl_010;
  wire G176_n_spl_0100;
  wire G176_n_spl_0101;
  wire G176_n_spl_011;
  wire G176_n_spl_1;
  wire G176_n_spl_10;
  wire G176_n_spl_100;
  wire G176_n_spl_101;
  wire G176_n_spl_11;
  wire G176_n_spl_110;
  wire G176_n_spl_111;
  wire g562_n_spl_;
  wire g562_n_spl_0;
  wire G2_p_spl_;
  wire G2_p_spl_0;
  wire G2_p_spl_1;
  wire G2_n_spl_;
  wire G2_n_spl_0;
  wire g570_n_spl_;
  wire g572_p_spl_;
  wire G173_n_spl_;
  wire G173_n_spl_0;
  wire G173_n_spl_00;
  wire G173_n_spl_000;
  wire G173_n_spl_0000;
  wire G173_n_spl_0001;
  wire G173_n_spl_001;
  wire G173_n_spl_0010;
  wire G173_n_spl_0011;
  wire G173_n_spl_01;
  wire G173_n_spl_010;
  wire G173_n_spl_011;
  wire G173_n_spl_1;
  wire G173_n_spl_10;
  wire G173_n_spl_100;
  wire G173_n_spl_101;
  wire G173_n_spl_11;
  wire G173_n_spl_110;
  wire G173_n_spl_111;
  wire G22_p_spl_;
  wire G173_p_spl_;
  wire G173_p_spl_0;
  wire G173_p_spl_00;
  wire G173_p_spl_000;
  wire G173_p_spl_0000;
  wire G173_p_spl_0001;
  wire G173_p_spl_001;
  wire G173_p_spl_0010;
  wire G173_p_spl_0011;
  wire G173_p_spl_01;
  wire G173_p_spl_010;
  wire G173_p_spl_011;
  wire G173_p_spl_1;
  wire G173_p_spl_10;
  wire G173_p_spl_100;
  wire G173_p_spl_101;
  wire G173_p_spl_11;
  wire G173_p_spl_110;
  wire G173_p_spl_111;
  wire G3_p_spl_;
  wire G172_n_spl_;
  wire G172_n_spl_0;
  wire G172_n_spl_00;
  wire G172_n_spl_000;
  wire G172_n_spl_001;
  wire G172_n_spl_01;
  wire G172_n_spl_1;
  wire G172_n_spl_10;
  wire G172_n_spl_11;
  wire g579_p_spl_;
  wire g579_p_spl_0;
  wire g579_p_spl_00;
  wire g579_p_spl_1;
  wire g560_p_spl_;
  wire g560_p_spl_0;
  wire g560_p_spl_00;
  wire g560_p_spl_1;
  wire G172_p_spl_;
  wire G172_p_spl_0;
  wire G172_p_spl_00;
  wire G172_p_spl_000;
  wire G172_p_spl_001;
  wire G172_p_spl_01;
  wire G172_p_spl_1;
  wire G172_p_spl_10;
  wire G172_p_spl_11;
  wire g594_n_spl_;
  wire g594_p_spl_;
  wire g595_n_spl_;
  wire g596_n_spl_;
  wire g596_n_spl_0;
  wire g596_p_spl_;
  wire g596_p_spl_0;
  wire g596_p_spl_1;
  wire g597_p_spl_;
  wire g598_p_spl_;
  wire g598_p_spl_0;
  wire g598_n_spl_;
  wire g598_n_spl_0;
  wire g601_p_spl_;
  wire g610_n_spl_;
  wire g617_p_spl_;
  wire g617_p_spl_0;
  wire g619_n_spl_;
  wire G174_n_spl_;
  wire G174_n_spl_0;
  wire G174_n_spl_00;
  wire G174_n_spl_000;
  wire G174_n_spl_0000;
  wire G174_n_spl_0001;
  wire G174_n_spl_001;
  wire G174_n_spl_0010;
  wire G174_n_spl_0011;
  wire G174_n_spl_01;
  wire G174_n_spl_010;
  wire G174_n_spl_011;
  wire G174_n_spl_1;
  wire G174_n_spl_10;
  wire G174_n_spl_100;
  wire G174_n_spl_101;
  wire G174_n_spl_11;
  wire G174_n_spl_110;
  wire G174_n_spl_111;
  wire G174_p_spl_;
  wire G174_p_spl_0;
  wire G174_p_spl_00;
  wire G174_p_spl_000;
  wire G174_p_spl_0000;
  wire G174_p_spl_0001;
  wire G174_p_spl_001;
  wire G174_p_spl_0010;
  wire G174_p_spl_0011;
  wire G174_p_spl_01;
  wire G174_p_spl_010;
  wire G174_p_spl_011;
  wire G174_p_spl_1;
  wire G174_p_spl_10;
  wire G174_p_spl_100;
  wire G174_p_spl_101;
  wire G174_p_spl_11;
  wire G174_p_spl_110;
  wire G174_p_spl_111;
  wire G175_n_spl_;
  wire G175_n_spl_0;
  wire G175_n_spl_00;
  wire G175_n_spl_000;
  wire G175_n_spl_001;
  wire G175_n_spl_01;
  wire G175_n_spl_1;
  wire G175_n_spl_10;
  wire G175_n_spl_11;
  wire G175_p_spl_;
  wire G175_p_spl_0;
  wire G175_p_spl_00;
  wire G175_p_spl_000;
  wire G175_p_spl_001;
  wire G175_p_spl_01;
  wire G175_p_spl_1;
  wire G175_p_spl_10;
  wire G175_p_spl_11;
  wire g638_p_spl_;
  wire g639_p_spl_;
  wire g643_n_spl_;
  wire g652_n_spl_;
  wire g659_p_spl_;
  wire g660_p_spl_;
  wire g664_n_spl_;
  wire g673_n_spl_;
  wire g681_p_spl_;
  wire g581_n_spl_;
  wire g581_n_spl_0;
  wire g581_n_spl_00;
  wire g581_n_spl_01;
  wire g581_n_spl_1;
  wire g581_n_spl_10;
  wire g581_n_spl_11;
  wire g681_n_spl_;
  wire g581_p_spl_;
  wire g581_p_spl_0;
  wire g581_p_spl_00;
  wire g581_p_spl_01;
  wire g581_p_spl_1;
  wire g687_n_spl_;
  wire g687_p_spl_;
  wire g696_n_spl_;
  wire g693_n_spl_;
  wire g696_p_spl_;
  wire g693_p_spl_;
  wire g699_n_spl_;
  wire g690_p_spl_;
  wire g699_p_spl_;
  wire g690_n_spl_;
  wire g711_n_spl_;
  wire g708_p_spl_;
  wire g711_p_spl_;
  wire g708_n_spl_;
  wire g717_n_spl_;
  wire g717_p_spl_;
  wire g723_n_spl_;
  wire g720_p_spl_;
  wire g723_p_spl_;
  wire g720_n_spl_;
  wire g729_n_spl_;
  wire g726_n_spl_;
  wire g729_p_spl_;
  wire g726_p_spl_;
  wire g430_p_spl_;
  wire g430_p_spl_0;
  wire g541_n_spl_;
  wire g541_n_spl_0;
  wire g541_n_spl_1;
  wire g737_p_spl_;
  wire g737_p_spl_0;
  wire g737_p_spl_00;
  wire g737_p_spl_1;
  wire g737_n_spl_;
  wire g737_n_spl_0;
  wire g737_n_spl_00;
  wire g737_n_spl_1;
  wire g743_p_spl_;
  wire g747_p_spl_;
  wire g389_p_spl_;
  wire g546_n_spl_;
  wire g546_n_spl_0;
  wire g395_p_spl_;
  wire g395_p_spl_0;
  wire g395_p_spl_00;
  wire g395_p_spl_1;
  wire g760_p_spl_;
  wire g755_p_spl_;
  wire g774_p_spl_;
  wire g774_p_spl_0;
  wire g774_p_spl_00;
  wire g774_p_spl_01;
  wire g774_p_spl_1;
  wire g774_n_spl_;
  wire g774_n_spl_0;
  wire g774_n_spl_00;
  wire g774_n_spl_01;
  wire g774_n_spl_1;
  wire g777_p_spl_;
  wire g444_n_spl_;
  wire g780_p_spl_;
  wire g780_p_spl_0;
  wire g780_p_spl_1;
  wire g780_n_spl_;
  wire g780_n_spl_0;
  wire g780_n_spl_1;
  wire g791_p_spl_;
  wire g785_p_spl_;
  wire G158_n_spl_;
  wire G158_n_spl_0;
  wire G158_n_spl_00;
  wire G158_n_spl_000;
  wire G158_n_spl_0000;
  wire G158_n_spl_0001;
  wire G158_n_spl_001;
  wire G158_n_spl_0010;
  wire G158_n_spl_0011;
  wire G158_n_spl_01;
  wire G158_n_spl_010;
  wire G158_n_spl_011;
  wire G158_n_spl_1;
  wire G158_n_spl_10;
  wire G158_n_spl_100;
  wire G158_n_spl_101;
  wire G158_n_spl_11;
  wire G158_n_spl_110;
  wire G158_n_spl_111;
  wire G81_p_spl_;
  wire G158_p_spl_;
  wire G158_p_spl_0;
  wire G158_p_spl_00;
  wire G158_p_spl_000;
  wire G158_p_spl_0000;
  wire G158_p_spl_0001;
  wire G158_p_spl_001;
  wire G158_p_spl_0010;
  wire G158_p_spl_0011;
  wire G158_p_spl_01;
  wire G158_p_spl_010;
  wire G158_p_spl_011;
  wire G158_p_spl_1;
  wire G158_p_spl_10;
  wire G158_p_spl_100;
  wire G158_p_spl_101;
  wire G158_p_spl_11;
  wire G158_p_spl_110;
  wire G158_p_spl_111;
  wire G80_p_spl_;
  wire G159_n_spl_;
  wire G159_n_spl_0;
  wire G159_n_spl_00;
  wire G159_n_spl_000;
  wire G159_n_spl_001;
  wire G159_n_spl_01;
  wire G159_n_spl_1;
  wire G159_n_spl_10;
  wire G159_n_spl_11;
  wire G159_p_spl_;
  wire G159_p_spl_0;
  wire G159_p_spl_00;
  wire G159_p_spl_000;
  wire G159_p_spl_001;
  wire G159_p_spl_01;
  wire G159_p_spl_1;
  wire G159_p_spl_10;
  wire G159_p_spl_11;
  wire G64_p_spl_;
  wire G64_p_spl_0;
  wire G64_p_spl_00;
  wire G64_p_spl_000;
  wire G64_p_spl_0000;
  wire G64_p_spl_0001;
  wire G64_p_spl_001;
  wire G64_p_spl_0010;
  wire G64_p_spl_01;
  wire G64_p_spl_010;
  wire G64_p_spl_011;
  wire G64_p_spl_1;
  wire G64_p_spl_10;
  wire G64_p_spl_100;
  wire G64_p_spl_101;
  wire G64_p_spl_11;
  wire G64_p_spl_110;
  wire G64_p_spl_111;
  wire G160_n_spl_;
  wire G160_n_spl_0;
  wire G160_n_spl_00;
  wire G160_n_spl_000;
  wire G160_n_spl_0000;
  wire G160_n_spl_0001;
  wire G160_n_spl_001;
  wire G160_n_spl_0010;
  wire G160_n_spl_0011;
  wire G160_n_spl_01;
  wire G160_n_spl_010;
  wire G160_n_spl_011;
  wire G160_n_spl_1;
  wire G160_n_spl_10;
  wire G160_n_spl_100;
  wire G160_n_spl_101;
  wire G160_n_spl_11;
  wire G160_n_spl_110;
  wire G160_n_spl_111;
  wire G160_p_spl_;
  wire G160_p_spl_0;
  wire G160_p_spl_00;
  wire G160_p_spl_000;
  wire G160_p_spl_0000;
  wire G160_p_spl_0001;
  wire G160_p_spl_001;
  wire G160_p_spl_0010;
  wire G160_p_spl_0011;
  wire G160_p_spl_01;
  wire G160_p_spl_010;
  wire G160_p_spl_011;
  wire G160_p_spl_1;
  wire G160_p_spl_10;
  wire G160_p_spl_100;
  wire G160_p_spl_101;
  wire G160_p_spl_11;
  wire G160_p_spl_110;
  wire G160_p_spl_111;
  wire G161_n_spl_;
  wire G161_n_spl_0;
  wire G161_n_spl_00;
  wire G161_n_spl_000;
  wire G161_n_spl_001;
  wire G161_n_spl_01;
  wire G161_n_spl_1;
  wire G161_n_spl_10;
  wire G161_n_spl_11;
  wire G161_p_spl_;
  wire G161_p_spl_0;
  wire G161_p_spl_00;
  wire G161_p_spl_000;
  wire G161_p_spl_001;
  wire G161_p_spl_01;
  wire G161_p_spl_1;
  wire G161_p_spl_10;
  wire G161_p_spl_11;
  wire G14_p_spl_;
  wire G16_p_spl_;
  wire g647_n_spl_;
  wire g647_n_spl_0;
  wire g647_n_spl_00;
  wire g647_n_spl_1;
  wire g605_n_spl_;
  wire g605_n_spl_0;
  wire g605_n_spl_00;
  wire g605_n_spl_1;
  wire G6_p_spl_;
  wire G27_p_spl_;
  wire g656_n_spl_;
  wire g656_n_spl_0;
  wire g656_n_spl_00;
  wire g656_n_spl_1;
  wire g614_n_spl_;
  wire g614_n_spl_0;
  wire g614_n_spl_00;
  wire g614_n_spl_1;
  wire G5_p_spl_;
  wire G26_p_spl_;
  wire g669_n_spl_;
  wire g669_n_spl_0;
  wire g669_n_spl_00;
  wire g669_n_spl_1;
  wire g624_n_spl_;
  wire g624_n_spl_0;
  wire g624_n_spl_00;
  wire g624_n_spl_1;
  wire G25_p_spl_;
  wire G24_p_spl_;
  wire g678_n_spl_;
  wire g678_n_spl_0;
  wire g678_n_spl_00;
  wire g678_n_spl_1;
  wire g569_p_spl_;
  wire g569_p_spl_0;
  wire g569_p_spl_00;
  wire g569_p_spl_1;
  wire G76_p_spl_;
  wire G86_p_spl_;
  wire G72_p_spl_;
  wire G82_p_spl_;
  wire G70_p_spl_;
  wire G71_p_spl_;
  wire G68_p_spl_;
  wire G69_p_spl_;
  wire G171_p_spl_;
  wire G171_n_spl_;
  wire G54_p_spl_;
  wire G61_n_spl_;
  wire G61_p_spl_;
  wire g975_p_spl_;
  wire g533_n_spl_;
  wire G99_n_spl_;
  wire g735_n_spl_;
  wire g184_n_spl_;
  wire G155_n_spl_;
  wire g179_n_spl_;
  wire g705_n_spl_;
  wire g506_n_spl_;
  wire g1025_n_spl_;
  wire g1025_n_spl_0;
  wire g1025_n_spl_00;
  wire g1025_n_spl_1;
  wire g990_p_spl_;
  wire g990_p_spl_0;
  wire g990_p_spl_00;
  wire g990_p_spl_1;
  wire G41_p_spl_;
  wire G42_p_spl_;
  wire G18_p_spl_;
  wire G17_p_spl_;
  wire g1032_n_spl_;
  wire g1032_n_spl_0;
  wire g1032_n_spl_00;
  wire g1032_n_spl_1;
  wire g997_n_spl_;
  wire g997_n_spl_0;
  wire g997_n_spl_00;
  wire g997_n_spl_1;
  wire G40_p_spl_;
  wire G39_p_spl_;
  wire g1039_n_spl_;
  wire g1039_n_spl_0;
  wire g1039_n_spl_00;
  wire g1039_n_spl_1;
  wire g1004_n_spl_;
  wire g1004_n_spl_0;
  wire g1004_n_spl_00;
  wire g1004_n_spl_1;
  wire G15_p_spl_;
  wire G36_p_spl_;
  wire g1046_n_spl_;
  wire g1046_n_spl_0;
  wire g1046_n_spl_00;
  wire g1046_n_spl_1;
  wire g1011_n_spl_;
  wire g1011_n_spl_0;
  wire g1011_n_spl_00;
  wire g1011_n_spl_1;
  wire G77_p_spl_;
  wire G87_p_spl_;
  wire G75_p_spl_;
  wire G85_p_spl_;
  wire G74_p_spl_;
  wire G84_p_spl_;
  wire G73_p_spl_;
  wire G83_p_spl_;
  wire g1202_n_spl_;
  wire g1200_p_spl_;
  wire g1202_p_spl_;
  wire g1200_n_spl_;
  wire g1223_p_spl_;
  wire g1214_n_spl_;
  wire g1223_n_spl_;
  wire g1214_p_spl_;
  wire g1238_p_spl_;
  wire g1229_n_spl_;
  wire g1238_n_spl_;
  wire g1229_p_spl_;
  wire g1241_p_spl_;
  wire g1241_n_spl_;
  wire g245_p_spl_;
  wire g1244_n_spl_;
  wire g1226_p_spl_;
  wire g1244_p_spl_;
  wire g1226_n_spl_;
  wire g1254_n_spl_;
  wire g1254_p_spl_;
  wire g617_n_spl_;
  wire g1257_p_spl_;
  wire g1257_n_spl_;
  wire G162_n_spl_;
  wire G162_p_spl_;
  wire g1263_p_spl_;
  wire g1260_p_spl_;
  wire g1263_n_spl_;
  wire g1260_n_spl_;
  wire g1268_n_spl_;
  wire g1268_p_spl_;
  wire g1271_n_spl_;
  wire g1266_n_spl_;
  wire g1271_p_spl_;
  wire g1266_p_spl_;
  wire g1275_n_spl_;
  wire g1275_p_spl_;
  wire g1278_p_spl_;
  wire g1278_n_spl_;
  wire g1281_p_spl_;
  wire g1281_n_spl_;
  wire g1282_n_spl_;
  wire g1282_p_spl_;
  wire g1284_n_spl_;
  wire g1284_p_spl_;
  wire g1288_n_spl_;
  wire g1288_p_spl_;
  wire g1299_p_spl_;
  wire g1299_n_spl_;
  wire g1308_n_spl_;
  wire g1329_p_spl_;
  wire g1320_n_spl_;
  wire g1329_n_spl_;
  wire g1320_p_spl_;
  wire g1341_n_spl_;
  wire g1341_p_spl_;
  wire g317_p_spl_;
  wire g1344_p_spl_;
  wire g1332_n_spl_;
  wire g1344_n_spl_;
  wire g1332_p_spl_;
  wire g1365_p_spl_;
  wire g1356_n_spl_;
  wire g1365_n_spl_;
  wire g1356_p_spl_;
  wire g1386_p_spl_;
  wire g1377_n_spl_;
  wire g1386_n_spl_;
  wire g1377_p_spl_;
  wire g1398_n_spl_;
  wire g1389_p_spl_;
  wire g1398_p_spl_;
  wire g1389_n_spl_;
  wire g1401_n_spl_;
  wire g1368_p_spl_;
  wire g1401_p_spl_;
  wire g1368_n_spl_;
  wire g1412_n_spl_;
  wire g1409_n_spl_;
  wire g1412_p_spl_;
  wire g1409_p_spl_;
  wire g1415_p_spl_;
  wire g1415_n_spl_;
  wire g1416_n_spl_;
  wire g1416_p_spl_;
  wire g1420_p_spl_;
  wire g1420_n_spl_;
  wire g1423_p_spl_;
  wire g1423_n_spl_;
  wire g1426_p_spl_;
  wire g1426_n_spl_;
  wire g1432_p_spl_;
  wire g1432_n_spl_;
  wire g1435_p_spl_;
  wire g1435_n_spl_;
  wire g1438_p_spl_;
  wire g1438_n_spl_;
  wire g1441_n_spl_;
  wire g1441_p_spl_;
  wire g1430_n_spl_;
  wire g1430_p_spl_;
  wire G157_n_spl_;
  wire G157_n_spl_0;
  wire G157_n_spl_1;
  wire G157_p_spl_;
  wire G157_p_spl_0;
  wire G157_p_spl_1;
  wire g1453_n_spl_;
  wire g1453_p_spl_;
  wire g1458_n_spl_;
  wire g1458_n_spl_0;
  wire g1458_n_spl_1;
  wire g1458_p_spl_;
  wire g1458_p_spl_0;
  wire g1458_p_spl_1;
  wire g1461_p_spl_;
  wire g1456_n_spl_;
  wire g1461_n_spl_;
  wire g1456_p_spl_;
  wire g1464_n_spl_;
  wire g1464_p_spl_;
  wire g1471_n_spl_;
  wire g1471_p_spl_;
  wire g1474_p_spl_;
  wire g1470_n_spl_;
  wire g1474_n_spl_;
  wire g1470_p_spl_;
  wire g1477_p_spl_;
  wire g1469_n_spl_;
  wire g1477_n_spl_;
  wire g1469_p_spl_;
  wire g1483_p_spl_;
  wire g1480_n_spl_;
  wire g1483_n_spl_;
  wire g1480_p_spl_;
  wire g1488_p_spl_;
  wire g1488_n_spl_;
  wire g1491_n_spl_;
  wire g1491_p_spl_;
  wire g1500_n_spl_;
  wire G23_n_spl_;
  wire G4_n_spl_;
  wire g1509_p_spl_;
  wire g1509_p_spl_0;
  wire g1509_p_spl_1;
  wire g1512_p_spl_;
  wire g1512_p_spl_0;
  wire g1512_p_spl_1;
  wire G79_n_spl_;
  wire G78_n_spl_;
  wire G64_n_spl_;
  wire G151_n_spl_;
  wire G151_n_spl_0;
  wire G152_p_spl_;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire G1_n_spl_1;
  wire g194_n_spl_;
  wire g431_n_spl_;
  wire g482_p_spl_;
  wire g549_p_spl_;
  wire g550_n_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  buf

  (
    G42_p,
    G42
  );


  not

  (
    G42_n,
    G42
  );


  buf

  (
    G43_p,
    G43
  );


  not

  (
    G43_n,
    G43
  );


  buf

  (
    G44_p,
    G44
  );


  not

  (
    G44_n,
    G44
  );


  buf

  (
    G45_p,
    G45
  );


  not

  (
    G45_n,
    G45
  );


  buf

  (
    G46_p,
    G46
  );


  not

  (
    G46_n,
    G46
  );


  buf

  (
    G47_p,
    G47
  );


  not

  (
    G47_n,
    G47
  );


  buf

  (
    G48_p,
    G48
  );


  not

  (
    G48_n,
    G48
  );


  buf

  (
    G49_p,
    G49
  );


  not

  (
    G49_n,
    G49
  );


  buf

  (
    G50_p,
    G50
  );


  not

  (
    G50_n,
    G50
  );


  buf

  (
    G51_p,
    G51
  );


  not

  (
    G51_n,
    G51
  );


  buf

  (
    G52_p,
    G52
  );


  not

  (
    G52_n,
    G52
  );


  buf

  (
    G53_p,
    G53
  );


  not

  (
    G53_n,
    G53
  );


  buf

  (
    G54_p,
    G54
  );


  not

  (
    G54_n,
    G54
  );


  buf

  (
    G55_p,
    G55
  );


  not

  (
    G55_n,
    G55
  );


  buf

  (
    G56_p,
    G56
  );


  not

  (
    G56_n,
    G56
  );


  buf

  (
    G57_p,
    G57
  );


  not

  (
    G57_n,
    G57
  );


  buf

  (
    G58_p,
    G58
  );


  not

  (
    G58_n,
    G58
  );


  buf

  (
    G59_p,
    G59
  );


  not

  (
    G59_n,
    G59
  );


  buf

  (
    G60_p,
    G60
  );


  not

  (
    G60_n,
    G60
  );


  buf

  (
    G61_p,
    G61
  );


  not

  (
    G61_n,
    G61
  );


  buf

  (
    G62_p,
    G62
  );


  not

  (
    G62_n,
    G62
  );


  buf

  (
    G63_p,
    G63
  );


  not

  (
    G63_n,
    G63
  );


  buf

  (
    G64_p,
    G64
  );


  not

  (
    G64_n,
    G64
  );


  buf

  (
    G65_p,
    G65
  );


  not

  (
    G65_n,
    G65
  );


  buf

  (
    G66_p,
    G66
  );


  not

  (
    G66_n,
    G66
  );


  buf

  (
    G67_p,
    G67
  );


  not

  (
    G67_n,
    G67
  );


  buf

  (
    G68_p,
    G68
  );


  not

  (
    G68_n,
    G68
  );


  buf

  (
    G69_p,
    G69
  );


  not

  (
    G69_n,
    G69
  );


  buf

  (
    G70_p,
    G70
  );


  not

  (
    G70_n,
    G70
  );


  buf

  (
    G71_p,
    G71
  );


  not

  (
    G71_n,
    G71
  );


  buf

  (
    G72_p,
    G72
  );


  not

  (
    G72_n,
    G72
  );


  buf

  (
    G73_p,
    G73
  );


  not

  (
    G73_n,
    G73
  );


  buf

  (
    G74_p,
    G74
  );


  not

  (
    G74_n,
    G74
  );


  buf

  (
    G75_p,
    G75
  );


  not

  (
    G75_n,
    G75
  );


  buf

  (
    G76_p,
    G76
  );


  not

  (
    G76_n,
    G76
  );


  buf

  (
    G77_p,
    G77
  );


  not

  (
    G77_n,
    G77
  );


  buf

  (
    G78_p,
    G78
  );


  not

  (
    G78_n,
    G78
  );


  buf

  (
    G79_p,
    G79
  );


  not

  (
    G79_n,
    G79
  );


  buf

  (
    G80_p,
    G80
  );


  not

  (
    G80_n,
    G80
  );


  buf

  (
    G81_p,
    G81
  );


  not

  (
    G81_n,
    G81
  );


  buf

  (
    G82_p,
    G82
  );


  not

  (
    G82_n,
    G82
  );


  buf

  (
    G83_p,
    G83
  );


  not

  (
    G83_n,
    G83
  );


  buf

  (
    G84_p,
    G84
  );


  not

  (
    G84_n,
    G84
  );


  buf

  (
    G85_p,
    G85
  );


  not

  (
    G85_n,
    G85
  );


  buf

  (
    G86_p,
    G86
  );


  not

  (
    G86_n,
    G86
  );


  buf

  (
    G87_p,
    G87
  );


  not

  (
    G87_n,
    G87
  );


  buf

  (
    G88_p,
    G88
  );


  not

  (
    G88_n,
    G88
  );


  buf

  (
    G89_p,
    G89
  );


  not

  (
    G89_n,
    G89
  );


  buf

  (
    G90_p,
    G90
  );


  not

  (
    G90_n,
    G90
  );


  buf

  (
    G91_p,
    G91
  );


  not

  (
    G91_n,
    G91
  );


  buf

  (
    G92_p,
    G92
  );


  not

  (
    G92_n,
    G92
  );


  buf

  (
    G93_p,
    G93
  );


  not

  (
    G93_n,
    G93
  );


  buf

  (
    G94_p,
    G94
  );


  not

  (
    G94_n,
    G94
  );


  buf

  (
    G95_p,
    G95
  );


  not

  (
    G95_n,
    G95
  );


  buf

  (
    G96_p,
    G96
  );


  not

  (
    G96_n,
    G96
  );


  buf

  (
    G97_p,
    G97
  );


  not

  (
    G97_n,
    G97
  );


  buf

  (
    G98_p,
    G98
  );


  not

  (
    G98_n,
    G98
  );


  buf

  (
    G99_p,
    G99
  );


  not

  (
    G99_n,
    G99
  );


  buf

  (
    G100_p,
    G100
  );


  not

  (
    G100_n,
    G100
  );


  buf

  (
    G101_p,
    G101
  );


  not

  (
    G101_n,
    G101
  );


  buf

  (
    G102_p,
    G102
  );


  not

  (
    G102_n,
    G102
  );


  buf

  (
    G103_p,
    G103
  );


  not

  (
    G103_n,
    G103
  );


  buf

  (
    G104_p,
    G104
  );


  not

  (
    G104_n,
    G104
  );


  buf

  (
    G105_p,
    G105
  );


  not

  (
    G105_n,
    G105
  );


  buf

  (
    G106_p,
    G106
  );


  not

  (
    G106_n,
    G106
  );


  buf

  (
    G107_p,
    G107
  );


  not

  (
    G107_n,
    G107
  );


  buf

  (
    G108_p,
    G108
  );


  not

  (
    G108_n,
    G108
  );


  buf

  (
    G109_p,
    G109
  );


  not

  (
    G109_n,
    G109
  );


  buf

  (
    G110_p,
    G110
  );


  not

  (
    G110_n,
    G110
  );


  buf

  (
    G111_p,
    G111
  );


  not

  (
    G111_n,
    G111
  );


  buf

  (
    G112_p,
    G112
  );


  not

  (
    G112_n,
    G112
  );


  buf

  (
    G113_p,
    G113
  );


  not

  (
    G113_n,
    G113
  );


  buf

  (
    G114_p,
    G114
  );


  not

  (
    G114_n,
    G114
  );


  buf

  (
    G115_p,
    G115
  );


  not

  (
    G115_n,
    G115
  );


  buf

  (
    G116_p,
    G116
  );


  not

  (
    G116_n,
    G116
  );


  buf

  (
    G117_p,
    G117
  );


  not

  (
    G117_n,
    G117
  );


  buf

  (
    G118_p,
    G118
  );


  not

  (
    G118_n,
    G118
  );


  buf

  (
    G119_p,
    G119
  );


  not

  (
    G119_n,
    G119
  );


  buf

  (
    G120_p,
    G120
  );


  not

  (
    G120_n,
    G120
  );


  buf

  (
    G121_p,
    G121
  );


  not

  (
    G121_n,
    G121
  );


  buf

  (
    G122_p,
    G122
  );


  not

  (
    G122_n,
    G122
  );


  buf

  (
    G123_p,
    G123
  );


  not

  (
    G123_n,
    G123
  );


  buf

  (
    G124_p,
    G124
  );


  not

  (
    G124_n,
    G124
  );


  buf

  (
    G125_p,
    G125
  );


  not

  (
    G125_n,
    G125
  );


  buf

  (
    G126_p,
    G126
  );


  not

  (
    G126_n,
    G126
  );


  buf

  (
    G127_p,
    G127
  );


  not

  (
    G127_n,
    G127
  );


  buf

  (
    G128_p,
    G128
  );


  not

  (
    G128_n,
    G128
  );


  buf

  (
    G129_p,
    G129
  );


  not

  (
    G129_n,
    G129
  );


  buf

  (
    G130_p,
    G130
  );


  not

  (
    G130_n,
    G130
  );


  buf

  (
    G131_p,
    G131
  );


  not

  (
    G131_n,
    G131
  );


  buf

  (
    G132_p,
    G132
  );


  not

  (
    G132_n,
    G132
  );


  buf

  (
    G133_p,
    G133
  );


  not

  (
    G133_n,
    G133
  );


  buf

  (
    G134_p,
    G134
  );


  not

  (
    G134_n,
    G134
  );


  buf

  (
    G135_p,
    G135
  );


  not

  (
    G135_n,
    G135
  );


  buf

  (
    G136_p,
    G136
  );


  not

  (
    G136_n,
    G136
  );


  buf

  (
    G137_p,
    G137
  );


  not

  (
    G137_n,
    G137
  );


  buf

  (
    G138_p,
    G138
  );


  not

  (
    G138_n,
    G138
  );


  buf

  (
    G139_p,
    G139
  );


  not

  (
    G139_n,
    G139
  );


  buf

  (
    G140_p,
    G140
  );


  not

  (
    G140_n,
    G140
  );


  buf

  (
    G141_p,
    G141
  );


  not

  (
    G141_n,
    G141
  );


  buf

  (
    G142_p,
    G142
  );


  not

  (
    G142_n,
    G142
  );


  buf

  (
    G143_p,
    G143
  );


  not

  (
    G143_n,
    G143
  );


  buf

  (
    G144_p,
    G144
  );


  not

  (
    G144_n,
    G144
  );


  buf

  (
    G145_p,
    G145
  );


  not

  (
    G145_n,
    G145
  );


  buf

  (
    G146_p,
    G146
  );


  not

  (
    G146_n,
    G146
  );


  buf

  (
    G147_p,
    G147
  );


  not

  (
    G147_n,
    G147
  );


  buf

  (
    G148_p,
    G148
  );


  not

  (
    G148_n,
    G148
  );


  buf

  (
    G149_p,
    G149
  );


  not

  (
    G149_n,
    G149
  );


  buf

  (
    G150_p,
    G150
  );


  not

  (
    G150_n,
    G150
  );


  buf

  (
    G151_p,
    G151
  );


  not

  (
    G151_n,
    G151
  );


  buf

  (
    G152_p,
    G152
  );


  not

  (
    G152_n,
    G152
  );


  buf

  (
    G153_p,
    G153
  );


  not

  (
    G153_n,
    G153
  );


  buf

  (
    G154_p,
    G154
  );


  not

  (
    G154_n,
    G154
  );


  buf

  (
    G155_p,
    G155
  );


  not

  (
    G155_n,
    G155
  );


  buf

  (
    G156_p,
    G156
  );


  not

  (
    G156_n,
    G156
  );


  buf

  (
    G157_p,
    G157
  );


  not

  (
    G157_n,
    G157
  );


  buf

  (
    G158_p,
    G158
  );


  not

  (
    G158_n,
    G158
  );


  buf

  (
    G159_p,
    G159
  );


  not

  (
    G159_n,
    G159
  );


  buf

  (
    G160_p,
    G160
  );


  not

  (
    G160_n,
    G160
  );


  buf

  (
    G161_p,
    G161
  );


  not

  (
    G161_n,
    G161
  );


  buf

  (
    G162_p,
    G162
  );


  not

  (
    G162_n,
    G162
  );


  buf

  (
    G163_p,
    G163
  );


  not

  (
    G163_n,
    G163
  );


  buf

  (
    G164_p,
    G164
  );


  not

  (
    G164_n,
    G164
  );


  buf

  (
    G165_p,
    G165
  );


  not

  (
    G165_n,
    G165
  );


  buf

  (
    G166_p,
    G166
  );


  not

  (
    G166_n,
    G166
  );


  buf

  (
    G167_p,
    G167
  );


  not

  (
    G167_n,
    G167
  );


  buf

  (
    G168_p,
    G168
  );


  not

  (
    G168_n,
    G168
  );


  buf

  (
    G169_p,
    G169
  );


  not

  (
    G169_n,
    G169
  );


  buf

  (
    G170_p,
    G170
  );


  not

  (
    G170_n,
    G170
  );


  buf

  (
    G171_p,
    G171
  );


  not

  (
    G171_n,
    G171
  );


  buf

  (
    G172_p,
    G172
  );


  not

  (
    G172_n,
    G172
  );


  buf

  (
    G173_p,
    G173
  );


  not

  (
    G173_n,
    G173
  );


  buf

  (
    G174_p,
    G174
  );


  not

  (
    G174_n,
    G174
  );


  buf

  (
    G175_p,
    G175
  );


  not

  (
    G175_n,
    G175
  );


  buf

  (
    G176_p,
    G176
  );


  not

  (
    G176_n,
    G176
  );


  buf

  (
    G177_p,
    G177
  );


  not

  (
    G177_n,
    G177
  );


  buf

  (
    G178_p,
    G178
  );


  not

  (
    G178_n,
    G178
  );


  or

  (
    g179_n,
    G156_n_spl_,
    G153_n_spl_
  );


  and

  (
    g180_p,
    G67_p,
    G66_p_spl_00
  );


  and

  (
    g181_p,
    G134_p,
    G1_p_spl_
  );


  and

  (
    g182_p,
    G165_n_spl_,
    G63_p
  );


  or

  (
    g183_n,
    G164_p,
    G11_n_spl_
  );


  or

  (
    g184_n,
    G154_n,
    G136_n
  );


  or

  (
    g185_n,
    G12_n,
    G11_n_spl_
  );


  or

  (
    g186_n,
    g185_n_spl_000,
    G65_n
  );


  or

  (
    g187_n,
    G163_n_spl_00,
    G34_n
  );


  or

  (
    g188_n,
    G163_p_spl_00,
    G33_n
  );


  and

  (
    g189_p,
    g188_n,
    g187_n
  );


  or

  (
    g190_n,
    g189_p,
    g185_n_spl_000
  );


  or

  (
    g191_n,
    G163_n_spl_00,
    G13_n
  );


  or

  (
    g192_n,
    G163_p_spl_00,
    G35_n
  );


  and

  (
    g193_p,
    g192_n,
    g191_n
  );


  or

  (
    g194_n,
    g193_p,
    g185_n_spl_00
  );


  or

  (
    g195_n,
    g185_n_spl_01,
    G32_n
  );


  and

  (
    g196_p,
    G163_p_spl_01,
    G8_p
  );


  and

  (
    g197_p,
    G163_n_spl_01,
    G9_p
  );


  or

  (
    g198_n,
    g197_p,
    g185_n_spl_01
  );


  or

  (
    g199_n,
    g198_n,
    g196_p
  );


  and

  (
    g200_p,
    g199_n,
    G66_p_spl_00
  );


  and

  (
    g201_p,
    G163_p_spl_01,
    G10_p
  );


  and

  (
    g202_p,
    G163_n_spl_01,
    G30_p
  );


  or

  (
    g203_n,
    g202_p,
    g185_n_spl_10
  );


  or

  (
    g204_n,
    g203_n,
    g201_p
  );


  and

  (
    g205_p,
    g204_n,
    G66_p_spl_01
  );


  and

  (
    g206_p,
    G163_p_spl_1,
    G28_p
  );


  and

  (
    g207_p,
    G163_n_spl_1,
    G7_p
  );


  or

  (
    g208_n,
    g207_p,
    g185_n_spl_10
  );


  or

  (
    g209_n,
    g208_n,
    g206_p
  );


  and

  (
    g210_p,
    g209_n,
    G66_p_spl_01
  );


  and

  (
    g211_p,
    G163_p_spl_1,
    G31_p
  );


  and

  (
    g212_p,
    G163_n_spl_1,
    G29_p
  );


  or

  (
    g213_n,
    g212_p,
    g185_n_spl_11
  );


  or

  (
    g214_n,
    g213_n,
    g211_p
  );


  and

  (
    g215_p,
    g214_n,
    G66_p_spl_1
  );


  and

  (
    g216_p,
    G168_p_spl_000,
    G128_p_spl_000
  );


  and

  (
    g217_p,
    G169_p_spl_000,
    G128_n_spl_000
  );


  or

  (
    g218_n,
    g217_p,
    g216_p
  );


  and

  (
    g219_p,
    g218_n,
    G150_p_spl_00
  );


  and

  (
    g220_p,
    G167_n_spl_000,
    G128_p_spl_000
  );


  and

  (
    g221_p,
    G166_n_spl_000,
    G128_n_spl_000
  );


  or

  (
    g222_n,
    g221_p,
    g220_p
  );


  and

  (
    g223_p,
    g222_n,
    G150_n_spl_00
  );


  or

  (
    g224_n,
    g223_p,
    g219_p
  );


  and

  (
    g225_p,
    G168_p_spl_000,
    G126_p_spl_000
  );


  and

  (
    g226_p,
    G169_p_spl_000,
    G126_n_spl_000
  );


  or

  (
    g227_n,
    g226_p,
    g225_p
  );


  and

  (
    g228_p,
    g227_n,
    G149_p_spl_00
  );


  and

  (
    g229_p,
    G167_n_spl_000,
    G126_p_spl_000
  );


  and

  (
    g230_p,
    G166_n_spl_000,
    G126_n_spl_000
  );


  or

  (
    g231_n,
    g230_p,
    g229_p
  );


  and

  (
    g232_p,
    g231_n,
    G149_n_spl_00
  );


  or

  (
    g233_n,
    g232_p,
    g228_p
  );


  or

  (
    g234_n,
    g233_n_spl_,
    g224_n_spl_
  );


  and

  (
    g235_p,
    G113_p_spl_00,
    G102_p_spl_000
  );


  or

  (
    g235_n,
    G113_n_spl_00,
    G102_n_spl_000
  );


  and

  (
    g236_p,
    G113_n_spl_00,
    G98_p_spl_000
  );


  or

  (
    g236_n,
    G113_p_spl_00,
    G98_n_spl_000
  );


  and

  (
    g237_p,
    g236_n,
    g235_n
  );


  or

  (
    g237_n,
    g236_p,
    g235_p
  );


  and

  (
    g238_p,
    G115_p_spl_00,
    G101_p_spl_000
  );


  or

  (
    g238_n,
    G115_n_spl_00,
    G101_n_spl_000
  );


  and

  (
    g239_p,
    G115_n_spl_00,
    G100_p_spl_0000
  );


  or

  (
    g239_n,
    G115_p_spl_00,
    G100_n_spl_0000
  );


  and

  (
    g240_p,
    g239_n,
    g238_n
  );


  or

  (
    g240_n,
    g239_p,
    g238_p
  );


  and

  (
    g241_p,
    g240_p_spl_,
    g237_n_spl_0
  );


  or

  (
    g241_n,
    g240_n_spl_0,
    g237_p_spl_
  );


  or

  (
    g242_n,
    g241_n_spl_,
    g234_n
  );


  and

  (
    g243_p,
    G130_p_spl_00,
    G101_p_spl_000
  );


  or

  (
    g243_n,
    G130_n_spl_00,
    G101_n_spl_000
  );


  and

  (
    g244_p,
    G130_n_spl_00,
    G100_p_spl_0000
  );


  or

  (
    g244_n,
    G130_p_spl_00,
    G100_n_spl_0000
  );


  and

  (
    g245_p,
    g244_n,
    g243_n
  );


  or

  (
    g245_n,
    g244_p,
    g243_p
  );


  and

  (
    g246_p,
    G166_n_spl_001,
    G148_n_spl_00
  );


  and

  (
    g247_p,
    G169_p_spl_001,
    G148_p_spl_00
  );


  or

  (
    g248_n,
    g247_p,
    g246_p
  );


  or

  (
    g249_n,
    g248_n_spl_,
    g245_n_spl_0
  );


  and

  (
    g250_p,
    G119_p_spl_00,
    G101_p_spl_001
  );


  or

  (
    g250_n,
    G119_n_spl_00,
    G101_n_spl_001
  );


  and

  (
    g251_p,
    G119_n_spl_00,
    G100_p_spl_000
  );


  or

  (
    g251_n,
    G119_p_spl_00,
    G100_n_spl_000
  );


  and

  (
    g252_p,
    g251_n,
    g250_n
  );


  or

  (
    g252_n,
    g251_p,
    g250_p
  );


  and

  (
    g253_p,
    g252_n,
    G146_p_spl_0
  );


  or

  (
    g253_n,
    g252_p,
    G146_n_spl_0
  );


  and

  (
    g254_p,
    G119_p_spl_01,
    G102_n_spl_000
  );


  or

  (
    g254_n,
    G119_n_spl_01,
    G102_p_spl_000
  );


  and

  (
    g255_p,
    G119_n_spl_01,
    G98_n_spl_000
  );


  or

  (
    g255_n,
    G119_p_spl_01,
    G98_p_spl_000
  );


  and

  (
    g256_p,
    g255_n,
    g254_n
  );


  or

  (
    g256_n,
    g255_p,
    g254_p
  );


  and

  (
    g257_p,
    g256_n,
    G146_n_spl_0
  );


  or

  (
    g257_n,
    g256_p,
    G146_p_spl_0
  );


  and

  (
    g258_p,
    g257_n,
    g253_n
  );


  or

  (
    g258_n,
    g257_p,
    g253_p
  );


  and

  (
    g259_p,
    G117_p_spl_00,
    G101_p_spl_001
  );


  or

  (
    g259_n,
    G117_n_spl_00,
    G101_n_spl_001
  );


  and

  (
    g260_p,
    G117_n_spl_00,
    G100_p_spl_001
  );


  or

  (
    g260_n,
    G117_p_spl_00,
    G100_n_spl_001
  );


  and

  (
    g261_p,
    g260_n,
    g259_n
  );


  or

  (
    g261_n,
    g260_p,
    g259_p
  );


  and

  (
    g262_p,
    g261_n,
    G145_p_spl_0
  );


  or

  (
    g262_n,
    g261_p,
    G145_n_spl_0
  );


  and

  (
    g263_p,
    G117_p_spl_01,
    G102_n_spl_001
  );


  or

  (
    g263_n,
    G117_n_spl_01,
    G102_p_spl_001
  );


  and

  (
    g264_p,
    G117_n_spl_01,
    G98_n_spl_001
  );


  or

  (
    g264_n,
    G117_p_spl_01,
    G98_p_spl_001
  );


  and

  (
    g265_p,
    g264_n,
    g263_n
  );


  or

  (
    g265_n,
    g264_p,
    g263_p
  );


  and

  (
    g266_p,
    g265_n,
    G145_n_spl_0
  );


  or

  (
    g266_n,
    g265_p,
    G145_p_spl_0
  );


  and

  (
    g267_p,
    g266_n,
    g262_n
  );


  or

  (
    g267_n,
    g266_p,
    g262_p
  );


  and

  (
    g268_p,
    g267_p_spl_,
    g258_p_spl_
  );


  or

  (
    g268_n,
    g267_n_spl_0,
    g258_n_spl_0
  );


  and

  (
    g269_p,
    G168_p_spl_001,
    G121_p_spl_000
  );


  and

  (
    g270_p,
    G169_p_spl_001,
    G121_n_spl_000
  );


  or

  (
    g271_n,
    g270_p,
    g269_p
  );


  and

  (
    g272_p,
    g271_n,
    G147_p_spl_00
  );


  and

  (
    g273_p,
    G167_n_spl_001,
    G121_p_spl_000
  );


  and

  (
    g274_p,
    G166_n_spl_001,
    G121_n_spl_000
  );


  or

  (
    g275_n,
    g274_p,
    g273_p
  );


  and

  (
    g276_p,
    g275_n,
    G147_n_spl_00
  );


  or

  (
    g277_n,
    g276_p,
    g272_p
  );


  or

  (
    g278_n,
    g277_n_spl_,
    g268_n_spl_
  );


  or

  (
    g279_n,
    g278_n,
    g249_n
  );


  or

  (
    g280_n,
    g279_n,
    g242_n
  );


  and

  (
    g281_p,
    G168_p_spl_001,
    G107_p_spl_000
  );


  and

  (
    g282_p,
    G169_p_spl_010,
    G107_n_spl_000
  );


  or

  (
    g283_n,
    g282_p,
    g281_p
  );


  and

  (
    g284_p,
    g283_n,
    G139_p_spl_00
  );


  and

  (
    g285_p,
    G167_n_spl_001,
    G107_p_spl_000
  );


  and

  (
    g286_p,
    G166_n_spl_010,
    G107_n_spl_000
  );


  or

  (
    g287_n,
    g286_p,
    g285_p
  );


  and

  (
    g288_p,
    g287_n,
    G139_n_spl_00
  );


  or

  (
    g289_n,
    g288_p,
    g284_p
  );


  and

  (
    g290_p,
    G168_p_spl_010,
    G105_p_spl_000
  );


  and

  (
    g291_p,
    G169_p_spl_010,
    G105_n_spl_000
  );


  or

  (
    g292_n,
    g291_p,
    g290_p
  );


  and

  (
    g293_p,
    g292_n,
    G138_p_spl_00
  );


  and

  (
    g294_p,
    G167_n_spl_010,
    G105_p_spl_000
  );


  and

  (
    g295_p,
    G166_n_spl_010,
    G105_n_spl_000
  );


  or

  (
    g296_n,
    g295_p,
    g294_p
  );


  and

  (
    g297_p,
    g296_n,
    G138_n_spl_00
  );


  or

  (
    g298_n,
    g297_p,
    g293_p
  );


  or

  (
    g299_n,
    g298_n_spl_,
    g289_n_spl_
  );


  and

  (
    g300_p,
    G168_p_spl_010,
    G109_p_spl_000
  );


  and

  (
    g301_p,
    G169_p_spl_011,
    G109_n_spl_000
  );


  or

  (
    g302_n,
    g301_p,
    g300_p
  );


  and

  (
    g303_p,
    g302_n,
    G135_p_spl_00
  );


  and

  (
    g304_p,
    G167_n_spl_010,
    G109_p_spl_000
  );


  and

  (
    g305_p,
    G166_n_spl_011,
    G109_n_spl_000
  );


  or

  (
    g306_n,
    g305_p,
    g304_p
  );


  and

  (
    g307_p,
    g306_n,
    G135_n_spl_00
  );


  or

  (
    g308_n,
    g307_p,
    g303_p
  );


  and

  (
    g309_p,
    G100_p_spl_001,
    G88_p_spl_00
  );


  or

  (
    g309_n,
    G100_n_spl_001,
    G88_n_spl_00
  );


  and

  (
    g310_p,
    G101_p_spl_010,
    G88_n_spl_00
  );


  or

  (
    g310_n,
    G101_n_spl_010,
    G88_p_spl_00
  );


  and

  (
    g311_p,
    g310_n,
    g309_n
  );


  or

  (
    g311_n,
    g310_p,
    g309_p
  );


  and

  (
    g312_p,
    g311_n,
    G142_p_spl_0
  );


  or

  (
    g312_n,
    g311_p,
    G142_n_spl_0
  );


  and

  (
    g313_p,
    G102_n_spl_001,
    G88_n_spl_01
  );


  or

  (
    g313_n,
    G102_p_spl_001,
    G88_p_spl_01
  );


  and

  (
    g314_p,
    G98_n_spl_001,
    G88_p_spl_01
  );


  or

  (
    g314_n,
    G98_p_spl_001,
    G88_n_spl_01
  );


  and

  (
    g315_p,
    g314_n,
    g313_n
  );


  or

  (
    g315_n,
    g314_p,
    g313_p
  );


  and

  (
    g316_p,
    g315_n,
    G142_n_spl_0
  );


  or

  (
    g316_n,
    g315_p,
    G142_p_spl_0
  );


  and

  (
    g317_p,
    g316_n,
    g312_n
  );


  or

  (
    g317_n,
    g316_p,
    g312_p
  );


  or

  (
    g318_n,
    g317_n_spl_0,
    g308_n_spl_
  );


  or

  (
    g319_n,
    g318_n,
    g299_n
  );


  and

  (
    g320_p,
    G168_p_spl_01,
    G90_p_spl_000
  );


  and

  (
    g321_p,
    G169_p_spl_011,
    G90_n_spl_000
  );


  or

  (
    g322_n,
    g321_p,
    g320_p
  );


  and

  (
    g323_p,
    g322_n,
    G143_p_spl_00
  );


  and

  (
    g324_p,
    G167_n_spl_01,
    G90_p_spl_000
  );


  and

  (
    g325_p,
    G166_n_spl_011,
    G90_n_spl_000
  );


  or

  (
    g326_n,
    g325_p,
    g324_p
  );


  and

  (
    g327_p,
    g326_n,
    G143_n_spl_00
  );


  or

  (
    g328_n,
    g327_p,
    g323_p
  );


  and

  (
    g329_p,
    G168_p_spl_10,
    G92_p_spl_000
  );


  and

  (
    g330_p,
    G169_p_spl_10,
    G92_n_spl_000
  );


  or

  (
    g331_n,
    g330_p,
    g329_p
  );


  and

  (
    g332_p,
    g331_n,
    G144_p_spl_00
  );


  and

  (
    g333_p,
    G167_n_spl_10,
    G92_p_spl_000
  );


  and

  (
    g334_p,
    G166_n_spl_10,
    G92_n_spl_000
  );


  or

  (
    g335_n,
    g334_p,
    g333_p
  );


  and

  (
    g336_p,
    g335_n,
    G144_n_spl_00
  );


  or

  (
    g337_n,
    g336_p,
    g332_p
  );


  or

  (
    g338_n,
    g337_n_spl_,
    g328_n_spl_
  );


  and

  (
    g339_p,
    G168_p_spl_10,
    G94_p_spl_000
  );


  and

  (
    g340_p,
    G169_p_spl_10,
    G94_n_spl_000
  );


  or

  (
    g341_n,
    g340_p,
    g339_p
  );


  and

  (
    g342_p,
    g341_n,
    G140_p_spl_00
  );


  and

  (
    g343_p,
    G167_n_spl_10,
    G94_p_spl_000
  );


  and

  (
    g344_p,
    G166_n_spl_10,
    G94_n_spl_000
  );


  or

  (
    g345_n,
    g344_p,
    g343_p
  );


  and

  (
    g346_p,
    g345_n,
    G140_n_spl_00
  );


  or

  (
    g347_n,
    g346_p,
    g342_p
  );


  and

  (
    g348_p,
    G168_p_spl_11,
    G96_p_spl_000
  );


  and

  (
    g349_p,
    G169_p_spl_11,
    G96_n_spl_000
  );


  or

  (
    g350_n,
    g349_p,
    g348_p
  );


  and

  (
    g351_p,
    g350_n,
    G141_p_spl_00
  );


  and

  (
    g352_p,
    G167_n_spl_11,
    G96_p_spl_000
  );


  and

  (
    g353_p,
    G166_n_spl_11,
    G96_n_spl_000
  );


  or

  (
    g354_n,
    g353_p,
    g352_p
  );


  and

  (
    g355_p,
    g354_n,
    G141_n_spl_00
  );


  or

  (
    g356_n,
    g355_p,
    g351_p
  );


  and

  (
    g357_p,
    G168_p_spl_11,
    G103_p_spl_000
  );


  and

  (
    g358_p,
    G169_p_spl_11,
    G103_n_spl_000
  );


  or

  (
    g359_n,
    g358_p,
    g357_p
  );


  and

  (
    g360_p,
    g359_n,
    G137_p_spl_00
  );


  and

  (
    g361_p,
    G167_n_spl_11,
    G103_p_spl_000
  );


  and

  (
    g362_p,
    G166_n_spl_11,
    G103_n_spl_000
  );


  or

  (
    g363_n,
    g362_p,
    g361_p
  );


  and

  (
    g364_p,
    g363_n,
    G137_n_spl_00
  );


  or

  (
    g365_n,
    g364_p,
    g360_p
  );


  or

  (
    g366_n,
    g365_n_spl_,
    g356_n_spl_
  );


  or

  (
    g367_n,
    g366_n,
    g347_n_spl_
  );


  or

  (
    g368_n,
    g367_n,
    g338_n
  );


  or

  (
    g369_n,
    g368_n,
    g319_n
  );


  and

  (
    g370_p,
    G124_n_spl_0000,
    G95_n
  );


  or

  (
    g370_n,
    G124_p_spl_0000,
    G95_p
  );


  and

  (
    g371_p,
    G124_p_spl_0000,
    G94_n_spl_00
  );


  or

  (
    g371_n,
    G124_n_spl_0000,
    G94_p_spl_00
  );


  and

  (
    g372_p,
    g371_n,
    g370_n
  );


  or

  (
    g372_n,
    g371_p,
    g370_p
  );


  and

  (
    g373_p,
    g372_p_spl_0,
    G140_p_spl_00
  );


  or

  (
    g373_n,
    g372_n_spl_0,
    G140_n_spl_00
  );


  and

  (
    g374_p,
    g372_n_spl_0,
    G140_n_spl_0
  );


  or

  (
    g374_n,
    g372_p_spl_0,
    G140_p_spl_0
  );


  and

  (
    g375_p,
    g374_n_spl_0,
    g373_n_spl_0
  );


  or

  (
    g375_n,
    g374_p_spl_0,
    g373_p_spl_0
  );


  and

  (
    g376_p,
    G124_n_spl_0001,
    G93_n
  );


  or

  (
    g376_n,
    G124_p_spl_0001,
    G93_p
  );


  and

  (
    g377_p,
    G124_p_spl_0001,
    G92_n_spl_00
  );


  or

  (
    g377_n,
    G124_n_spl_0001,
    G92_p_spl_00
  );


  and

  (
    g378_p,
    g377_n,
    g376_n
  );


  or

  (
    g378_n,
    g377_p,
    g376_p
  );


  and

  (
    g379_p,
    g378_p_spl_0,
    G144_p_spl_00
  );


  or

  (
    g379_n,
    g378_n_spl_0,
    G144_n_spl_00
  );


  and

  (
    g380_p,
    g378_n_spl_0,
    G144_n_spl_0
  );


  or

  (
    g380_n,
    g378_p_spl_0,
    G144_p_spl_0
  );


  and

  (
    g381_p,
    g380_n_spl_,
    g379_n_spl_
  );


  or

  (
    g381_n,
    g380_p_spl_,
    g379_p_spl_
  );


  and

  (
    g382_p,
    g381_p_spl_00,
    g375_p_spl_00
  );


  or

  (
    g382_n,
    g381_n_spl_00,
    g375_n_spl_00
  );


  and

  (
    g383_p,
    G124_n_spl_0010,
    G91_n
  );


  or

  (
    g383_n,
    G124_p_spl_0010,
    G91_p
  );


  and

  (
    g384_p,
    G124_p_spl_0010,
    G90_n_spl_00
  );


  or

  (
    g384_n,
    G124_n_spl_0010,
    G90_p_spl_00
  );


  and

  (
    g385_p,
    g384_n,
    g383_n
  );


  or

  (
    g385_n,
    g384_p,
    g383_p
  );


  and

  (
    g386_p,
    g385_p_spl_0,
    G143_p_spl_00
  );


  or

  (
    g386_n,
    g385_n_spl_0,
    G143_n_spl_00
  );


  and

  (
    g387_p,
    g385_n_spl_0,
    G143_n_spl_0
  );


  or

  (
    g387_n,
    g385_p_spl_0,
    G143_p_spl_0
  );


  and

  (
    g388_p,
    g387_n_spl_,
    g386_n_spl_
  );


  or

  (
    g388_n,
    g387_p_spl_,
    g386_p_spl_
  );


  and

  (
    g389_p,
    g388_p_spl_00,
    g382_p_spl_
  );


  or

  (
    g389_n,
    g388_n_spl_00,
    g382_n_spl_
  );


  and

  (
    g390_p,
    G124_n_spl_0011,
    G89_n
  );


  or

  (
    g390_n,
    G124_p_spl_0011,
    G89_p
  );


  and

  (
    g391_p,
    G124_p_spl_0011,
    G88_n_spl_10
  );


  or

  (
    g391_n,
    G124_n_spl_0011,
    G88_p_spl_10
  );


  and

  (
    g392_p,
    g391_n,
    g390_n
  );


  or

  (
    g392_n,
    g391_p,
    g390_p
  );


  and

  (
    g393_p,
    g392_p_spl_0,
    G142_p_spl_1
  );


  or

  (
    g393_n,
    g392_n_spl_0,
    G142_n_spl_1
  );


  and

  (
    g394_p,
    g392_n_spl_0,
    G142_n_spl_1
  );


  or

  (
    g394_n,
    g392_p_spl_0,
    G142_p_spl_1
  );


  and

  (
    g395_p,
    g394_n,
    g393_n_spl_
  );


  or

  (
    g395_n,
    g394_p,
    g393_p
  );


  or

  (
    g396_n,
    g395_n_spl_00,
    g389_n_spl_0
  );


  and

  (
    g397_p,
    G124_n_spl_010,
    G110_n
  );


  or

  (
    g397_n,
    G124_p_spl_010,
    G110_p
  );


  and

  (
    g398_p,
    G124_p_spl_010,
    G109_n_spl_00
  );


  or

  (
    g398_n,
    G124_n_spl_010,
    G109_p_spl_00
  );


  and

  (
    g399_p,
    g398_n,
    g397_n
  );


  or

  (
    g399_n,
    g398_p,
    g397_p
  );


  and

  (
    g400_p,
    g399_p_spl_0,
    G135_p_spl_00
  );


  or

  (
    g400_n,
    g399_n_spl_0,
    G135_n_spl_00
  );


  and

  (
    g401_p,
    g399_n_spl_0,
    G135_n_spl_0
  );


  or

  (
    g401_n,
    g399_p_spl_0,
    G135_p_spl_0
  );


  and

  (
    g402_p,
    g401_n_spl_0,
    g400_n_spl_00
  );


  or

  (
    g402_n,
    g401_p_spl_0,
    g400_p_spl_00
  );


  and

  (
    g403_p,
    G124_n_spl_011,
    G108_n
  );


  or

  (
    g403_n,
    G124_p_spl_011,
    G108_p
  );


  and

  (
    g404_p,
    G124_p_spl_011,
    G107_n_spl_00
  );


  or

  (
    g404_n,
    G124_n_spl_011,
    G107_p_spl_00
  );


  and

  (
    g405_p,
    g404_n,
    g403_n
  );


  or

  (
    g405_n,
    g404_p,
    g403_p
  );


  and

  (
    g406_p,
    g405_p_spl_0,
    G139_p_spl_00
  );


  or

  (
    g406_n,
    g405_n_spl_0,
    G139_n_spl_00
  );


  and

  (
    g407_p,
    g405_n_spl_0,
    G139_n_spl_0
  );


  or

  (
    g407_n,
    g405_p_spl_0,
    G139_p_spl_0
  );


  and

  (
    g408_p,
    g407_n,
    g406_n_spl_0
  );


  or

  (
    g408_n,
    g407_p,
    g406_p_spl_0
  );


  and

  (
    g409_p,
    g408_p_spl_0,
    g402_p_spl_0
  );


  or

  (
    g409_n,
    g408_n_spl_00,
    g402_n_spl_0
  );


  and

  (
    g410_p,
    G124_n_spl_100,
    G106_n
  );


  or

  (
    g410_n,
    G124_p_spl_100,
    G106_p
  );


  and

  (
    g411_p,
    G124_p_spl_100,
    G105_n_spl_00
  );


  or

  (
    g411_n,
    G124_n_spl_100,
    G105_p_spl_00
  );


  and

  (
    g412_p,
    g411_n,
    g410_n
  );


  or

  (
    g412_n,
    g411_p,
    g410_p
  );


  and

  (
    g413_p,
    g412_p_spl_0,
    G138_p_spl_00
  );


  or

  (
    g413_n,
    g412_n_spl_0,
    G138_n_spl_00
  );


  and

  (
    g414_p,
    g412_n_spl_0,
    G138_n_spl_0
  );


  or

  (
    g414_n,
    g412_p_spl_0,
    G138_p_spl_0
  );


  and

  (
    g415_p,
    g414_n,
    g413_n_spl_
  );


  or

  (
    g415_n,
    g414_p,
    g413_p_spl_
  );


  and

  (
    g416_p,
    g415_p_spl_00,
    g409_p_spl_0
  );


  or

  (
    g416_n,
    g415_n_spl_00,
    g409_n_spl_0
  );


  and

  (
    g417_p,
    G124_n_spl_101,
    G104_n
  );


  or

  (
    g417_n,
    G124_p_spl_101,
    G104_p
  );


  and

  (
    g418_p,
    G124_p_spl_101,
    G103_n_spl_00
  );


  or

  (
    g418_n,
    G124_n_spl_101,
    G103_p_spl_00
  );


  and

  (
    g419_p,
    g418_n,
    g417_n
  );


  or

  (
    g419_n,
    g418_p,
    g417_p
  );


  and

  (
    g420_p,
    g419_p_spl_0,
    G137_p_spl_00
  );


  or

  (
    g420_n,
    g419_n_spl_0,
    G137_n_spl_00
  );


  and

  (
    g421_p,
    g419_n_spl_0,
    G137_n_spl_0
  );


  or

  (
    g421_n,
    g419_p_spl_0,
    G137_p_spl_0
  );


  and

  (
    g422_p,
    g421_n,
    g420_n_spl_0
  );


  or

  (
    g422_n,
    g421_p,
    g420_p_spl_0
  );


  and

  (
    g423_p,
    g422_p_spl_00,
    g416_p_spl_0
  );


  or

  (
    g423_n,
    g422_n_spl_00,
    g416_n_spl_0
  );


  and

  (
    g424_p,
    G124_n_spl_110,
    G97_n
  );


  or

  (
    g424_n,
    G124_p_spl_110,
    G97_p
  );


  and

  (
    g425_p,
    G124_p_spl_110,
    G96_n_spl_00
  );


  or

  (
    g425_n,
    G124_n_spl_110,
    G96_p_spl_00
  );


  and

  (
    g426_p,
    g425_n,
    g424_n
  );


  or

  (
    g426_n,
    g425_p,
    g424_p
  );


  and

  (
    g427_p,
    g426_p_spl_0,
    G141_p_spl_00
  );


  or

  (
    g427_n,
    g426_n_spl_0,
    G141_n_spl_00
  );


  and

  (
    g428_p,
    g426_n_spl_0,
    G141_n_spl_0
  );


  or

  (
    g428_n,
    g426_p_spl_0,
    G141_p_spl_0
  );


  and

  (
    g429_p,
    g428_n,
    g427_n_spl_
  );


  or

  (
    g429_n,
    g428_p,
    g427_p_spl_
  );


  and

  (
    g430_p,
    g429_p_spl_00,
    g423_p_spl_
  );


  or

  (
    g430_n,
    g429_n_spl_00,
    g423_n_spl_
  );


  or

  (
    g431_n,
    g430_n_spl_0,
    g396_n_spl_
  );


  and

  (
    g432_p,
    G123_n_spl_0000,
    G118_n
  );


  or

  (
    g432_n,
    G123_p_spl_0000,
    G118_p
  );


  and

  (
    g433_p,
    G123_p_spl_0000,
    G117_n_spl_10
  );


  or

  (
    g433_n,
    G123_n_spl_0000,
    G117_p_spl_10
  );


  and

  (
    g434_p,
    g433_n,
    g432_n
  );


  or

  (
    g434_n,
    g433_p,
    g432_p
  );


  and

  (
    g435_p,
    g434_p_spl_0,
    G145_p_spl_1
  );


  or

  (
    g435_n,
    g434_n_spl_0,
    G145_n_spl_1
  );


  and

  (
    g436_p,
    g434_n_spl_0,
    G145_n_spl_1
  );


  or

  (
    g436_n,
    g434_p_spl_0,
    G145_p_spl_1
  );


  and

  (
    g437_p,
    g436_n,
    g435_n_spl_
  );


  or

  (
    g437_n,
    g436_p,
    g435_p_spl_
  );


  and

  (
    g438_p,
    G123_n_spl_0001,
    G120_n
  );


  or

  (
    g438_n,
    G123_p_spl_0001,
    G120_p
  );


  and

  (
    g439_p,
    G123_p_spl_0001,
    G119_n_spl_10
  );


  or

  (
    g439_n,
    G123_n_spl_0001,
    G119_p_spl_10
  );


  and

  (
    g440_p,
    g439_n,
    g438_n
  );


  or

  (
    g440_n,
    g439_p,
    g438_p
  );


  and

  (
    g441_p,
    g440_p_spl_0,
    G146_p_spl_1
  );


  or

  (
    g441_n,
    g440_n_spl_0,
    G146_n_spl_1
  );


  and

  (
    g442_p,
    g440_n_spl_0,
    G146_n_spl_1
  );


  or

  (
    g442_n,
    g440_p_spl_0,
    G146_p_spl_1
  );


  and

  (
    g443_p,
    g442_n_spl_0,
    g441_n_spl_00
  );


  or

  (
    g443_n,
    g442_p_spl_0,
    g441_p_spl_00
  );


  and

  (
    g444_p,
    g443_p_spl_00,
    g437_p_spl_00
  );


  or

  (
    g444_n,
    g443_n_spl_00,
    g437_n_spl_00
  );


  and

  (
    g445_p,
    G123_n_spl_0010,
    G122_n
  );


  or

  (
    g445_n,
    G123_p_spl_0010,
    G122_p
  );


  and

  (
    g446_p,
    G123_p_spl_0010,
    G121_n_spl_00
  );


  or

  (
    g446_n,
    G123_n_spl_0010,
    G121_p_spl_00
  );


  and

  (
    g447_p,
    g446_n,
    g445_n
  );


  or

  (
    g447_n,
    g446_p,
    g445_p
  );


  and

  (
    g448_p,
    g447_p_spl_0,
    G147_p_spl_00
  );


  or

  (
    g448_n,
    g447_n_spl_0,
    G147_n_spl_00
  );


  and

  (
    g449_p,
    g447_n_spl_0,
    G147_n_spl_0
  );


  or

  (
    g449_n,
    g447_p_spl_0,
    G147_p_spl_0
  );


  and

  (
    g450_p,
    g449_n,
    g448_n_spl_
  );


  or

  (
    g450_n,
    g449_p,
    g448_p_spl_
  );


  and

  (
    g451_p,
    G125_n_spl_,
    G123_n_spl_001
  );


  or

  (
    g451_n,
    G125_p,
    G123_p_spl_001
  );


  and

  (
    g452_p,
    g451_n_spl_0,
    G148_p_spl_00
  );


  or

  (
    g452_n,
    g451_p_spl_0,
    G148_n_spl_00
  );


  and

  (
    g453_p,
    g451_p_spl_0,
    G148_n_spl_0
  );


  or

  (
    g453_n,
    g451_n_spl_0,
    G148_p_spl_0
  );


  and

  (
    g454_p,
    g453_n,
    g452_n_spl_0
  );


  or

  (
    g454_n,
    g453_p,
    g452_p_spl_0
  );


  and

  (
    g455_p,
    g454_p_spl_0,
    g450_p_spl_0
  );


  or

  (
    g455_n,
    g454_n_spl_00,
    g450_n_spl_0
  );


  and

  (
    g456_p,
    G129_n_spl_,
    G123_n_spl_010
  );


  or

  (
    g456_n,
    G129_p,
    G123_p_spl_010
  );


  and

  (
    g457_p,
    G128_n_spl_00,
    G123_p_spl_010
  );


  or

  (
    g457_n,
    G128_p_spl_00,
    G123_n_spl_010
  );


  and

  (
    g458_p,
    g457_n,
    g456_n
  );


  or

  (
    g458_n,
    g457_p,
    g456_p
  );


  and

  (
    g459_p,
    g458_p_spl_0,
    G150_p_spl_00
  );


  or

  (
    g459_n,
    g458_n_spl_0,
    G150_n_spl_00
  );


  and

  (
    g460_p,
    g458_n_spl_0,
    G150_n_spl_0
  );


  or

  (
    g460_n,
    g458_p_spl_0,
    G150_p_spl_0
  );


  and

  (
    g461_p,
    g460_n,
    g459_n_spl_0
  );


  or

  (
    g461_n,
    g460_p,
    g459_p_spl_0
  );


  and

  (
    g462_p,
    G131_n_spl_,
    G123_n_spl_011
  );


  or

  (
    g462_n,
    G131_p,
    G123_p_spl_011
  );


  and

  (
    g463_p,
    G130_n_spl_0,
    G123_p_spl_011
  );


  or

  (
    g463_n,
    G130_p_spl_0,
    G123_n_spl_011
  );


  and

  (
    g464_p,
    g463_n,
    g462_n
  );


  or

  (
    g464_n,
    g463_p,
    g462_p
  );


  and

  (
    g465_p,
    g464_n_spl_00,
    g461_p_spl_0
  );


  or

  (
    g465_n,
    g464_p_spl_00,
    g461_n_spl_0
  );


  and

  (
    g466_p,
    G127_n_spl_,
    G123_n_spl_100
  );


  or

  (
    g466_n,
    G127_p,
    G123_p_spl_100
  );


  and

  (
    g467_p,
    G126_n_spl_00,
    G123_p_spl_100
  );


  or

  (
    g467_n,
    G126_p_spl_00,
    G123_n_spl_100
  );


  and

  (
    g468_p,
    g467_n,
    g466_n
  );


  or

  (
    g468_n,
    g467_p,
    g466_p
  );


  and

  (
    g469_p,
    g468_p_spl_0,
    G149_p_spl_00
  );


  or

  (
    g469_n,
    g468_n_spl_0,
    G149_n_spl_00
  );


  and

  (
    g470_p,
    g468_n_spl_0,
    G149_n_spl_0
  );


  or

  (
    g470_n,
    g468_p_spl_0,
    G149_p_spl_0
  );


  and

  (
    g471_p,
    g470_n,
    g469_n_spl_0
  );


  or

  (
    g471_n,
    g470_p,
    g469_p_spl_0
  );


  and

  (
    g472_p,
    g471_p_spl_0,
    g465_p_spl_0
  );


  or

  (
    g472_n,
    g471_n_spl_00,
    g465_n_spl_0
  );


  and

  (
    g473_p,
    g472_p_spl_,
    g455_p_spl_
  );


  or

  (
    g473_n,
    g472_n_spl_,
    g455_n_spl_
  );


  and

  (
    g474_p,
    G123_n_spl_101,
    G114_n_spl_0
  );


  or

  (
    g474_n,
    G123_p_spl_101,
    G114_p_spl_
  );


  and

  (
    g475_p,
    G123_p_spl_101,
    G113_n_spl_01
  );


  or

  (
    g475_n,
    G123_n_spl_101,
    G113_p_spl_0
  );


  and

  (
    g476_p,
    g475_n,
    g474_n
  );


  or

  (
    g476_n,
    g475_p,
    g474_p
  );


  and

  (
    g477_p,
    G123_n_spl_110,
    G116_n
  );


  or

  (
    g477_n,
    G123_p_spl_110,
    G116_p
  );


  and

  (
    g478_p,
    G123_p_spl_110,
    G115_n_spl_0
  );


  or

  (
    g478_n,
    G123_n_spl_110,
    G115_p_spl_0
  );


  and

  (
    g479_p,
    g478_n,
    g477_n
  );


  or

  (
    g479_n,
    g478_p,
    g477_p
  );


  and

  (
    g480_p,
    g479_n_spl_00,
    g476_n_spl_0
  );


  or

  (
    g480_n,
    g479_p_spl_00,
    g476_p_spl_00
  );


  and

  (
    g481_p,
    g480_p_spl_0,
    g473_p_spl_
  );


  and

  (
    g482_p,
    g481_p,
    g444_p_spl_0
  );


  and

  (
    g483_p,
    G119_n_spl_10,
    G117_n_spl_10
  );


  or

  (
    g483_n,
    G119_p_spl_10,
    G117_p_spl_10
  );


  and

  (
    g484_p,
    G119_p_spl_1,
    G117_p_spl_1
  );


  or

  (
    g484_n,
    G119_n_spl_1,
    G117_n_spl_1
  );


  and

  (
    g485_p,
    g484_n,
    g483_n
  );


  or

  (
    g485_n,
    g484_p,
    g483_p
  );


  and

  (
    g486_p,
    G115_n_spl_1,
    G113_n_spl_01
  );


  or

  (
    g486_n,
    G115_p_spl_1,
    G113_p_spl_1
  );


  and

  (
    g487_p,
    G115_p_spl_1,
    G113_p_spl_1
  );


  or

  (
    g487_n,
    G115_n_spl_1,
    G113_n_spl_1
  );


  and

  (
    g488_p,
    g487_n,
    g486_n
  );


  or

  (
    g488_n,
    g487_p,
    g486_p
  );


  and

  (
    g489_p,
    g488_n_spl_,
    g485_p_spl_
  );


  or

  (
    g489_n,
    g488_p_spl_,
    g485_n_spl_
  );


  and

  (
    g490_p,
    g488_p_spl_,
    g485_n_spl_
  );


  or

  (
    g490_n,
    g488_n_spl_,
    g485_p_spl_
  );


  and

  (
    g491_p,
    g490_n,
    g489_n
  );


  or

  (
    g491_n,
    g490_p,
    g489_p
  );


  and

  (
    g492_p,
    G132_n_spl_0,
    G130_n_spl_1
  );


  or

  (
    g492_n,
    G132_p_spl_0,
    G130_p_spl_1
  );


  and

  (
    g493_p,
    G132_p_spl_0,
    G130_p_spl_1
  );


  or

  (
    g493_n,
    G132_n_spl_0,
    G130_n_spl_1
  );


  and

  (
    g494_p,
    g493_n,
    g492_n
  );


  or

  (
    g494_n,
    g493_p,
    g492_p
  );


  and

  (
    g495_p,
    g494_n_spl_,
    G121_p_spl_01
  );


  or

  (
    g495_n,
    g494_p_spl_,
    G121_n_spl_01
  );


  and

  (
    g496_p,
    g494_p_spl_,
    G121_n_spl_01
  );


  or

  (
    g496_n,
    g494_n_spl_,
    G121_p_spl_01
  );


  and

  (
    g497_p,
    g496_n,
    g495_n
  );


  or

  (
    g497_n,
    g496_p,
    g495_p
  );


  and

  (
    g498_p,
    G128_n_spl_01,
    G126_n_spl_01
  );


  or

  (
    g498_n,
    G128_p_spl_01,
    G126_p_spl_01
  );


  and

  (
    g499_p,
    G128_p_spl_01,
    G126_p_spl_01
  );


  or

  (
    g499_n,
    G128_n_spl_01,
    G126_n_spl_01
  );


  and

  (
    g500_p,
    g499_n,
    g498_n
  );


  or

  (
    g500_n,
    g499_p,
    g498_p
  );


  and

  (
    g501_p,
    g500_n_spl_,
    g497_n_spl_
  );


  or

  (
    g501_n,
    g500_p_spl_,
    g497_p_spl_
  );


  and

  (
    g502_p,
    g500_p_spl_,
    g497_p_spl_
  );


  or

  (
    g502_n,
    g500_n_spl_,
    g497_n_spl_
  );


  and

  (
    g503_p,
    g502_n,
    g501_n
  );


  or

  (
    g503_n,
    g502_p,
    g501_p
  );


  and

  (
    g504_p,
    g503_p,
    g491_n
  );


  and

  (
    g505_p,
    g503_n,
    g491_p
  );


  or

  (
    g506_n,
    g505_p,
    g504_p
  );


  and

  (
    g507_p,
    G94_n_spl_01,
    G92_n_spl_01
  );


  or

  (
    g507_n,
    G94_p_spl_01,
    G92_p_spl_01
  );


  and

  (
    g508_p,
    G94_p_spl_01,
    G92_p_spl_01
  );


  or

  (
    g508_n,
    G94_n_spl_01,
    G92_n_spl_01
  );


  and

  (
    g509_p,
    g508_n,
    g507_n
  );


  or

  (
    g509_n,
    g508_p,
    g507_p
  );


  and

  (
    g510_p,
    G90_n_spl_01,
    G88_p_spl_10
  );


  or

  (
    g510_n,
    G90_p_spl_01,
    G88_n_spl_10
  );


  and

  (
    g511_p,
    G90_p_spl_01,
    G88_n_spl_1
  );


  or

  (
    g511_n,
    G90_n_spl_01,
    G88_p_spl_1
  );


  and

  (
    g512_p,
    g511_n,
    g510_n
  );


  or

  (
    g512_n,
    g511_p,
    g510_p
  );


  and

  (
    g513_p,
    g512_n_spl_,
    g509_p_spl_
  );


  or

  (
    g513_n,
    g512_p_spl_,
    g509_n_spl_
  );


  and

  (
    g514_p,
    g512_p_spl_,
    g509_n_spl_
  );


  or

  (
    g514_n,
    g512_n_spl_,
    g509_p_spl_
  );


  and

  (
    g515_p,
    g514_n,
    g513_n
  );


  or

  (
    g515_n,
    g514_p,
    g513_p
  );


  and

  (
    g516_p,
    G103_n_spl_01,
    G96_n_spl_01
  );


  or

  (
    g516_n,
    G103_p_spl_01,
    G96_p_spl_01
  );


  and

  (
    g517_p,
    G103_p_spl_01,
    G96_p_spl_01
  );


  or

  (
    g517_n,
    G103_n_spl_01,
    G96_n_spl_01
  );


  and

  (
    g518_p,
    g517_n,
    g516_n
  );


  or

  (
    g518_n,
    g517_p,
    g516_p
  );


  and

  (
    g519_p,
    G111_n_spl_0,
    G109_n_spl_01
  );


  or

  (
    g519_n,
    G111_p_spl_0,
    G109_p_spl_01
  );


  and

  (
    g520_p,
    G111_p_spl_0,
    G109_p_spl_01
  );


  or

  (
    g520_n,
    G111_n_spl_0,
    G109_n_spl_01
  );


  and

  (
    g521_p,
    g520_n,
    g519_n
  );


  or

  (
    g521_n,
    g520_p,
    g519_p
  );


  and

  (
    g522_p,
    g521_n_spl_,
    g518_n_spl_
  );


  or

  (
    g522_n,
    g521_p_spl_,
    g518_p_spl_
  );


  and

  (
    g523_p,
    g521_p_spl_,
    g518_p_spl_
  );


  or

  (
    g523_n,
    g521_n_spl_,
    g518_n_spl_
  );


  and

  (
    g524_p,
    g523_n,
    g522_n
  );


  or

  (
    g524_n,
    g523_p,
    g522_p
  );


  and

  (
    g525_p,
    G107_n_spl_01,
    G105_n_spl_01
  );


  or

  (
    g525_n,
    G107_p_spl_01,
    G105_p_spl_01
  );


  and

  (
    g526_p,
    G107_p_spl_01,
    G105_p_spl_01
  );


  or

  (
    g526_n,
    G107_n_spl_01,
    G105_n_spl_01
  );


  and

  (
    g527_p,
    g526_n,
    g525_n
  );


  or

  (
    g527_n,
    g526_p,
    g525_p
  );


  and

  (
    g528_p,
    g527_n_spl_,
    g524_n_spl_
  );


  or

  (
    g528_n,
    g527_p_spl_,
    g524_p_spl_
  );


  and

  (
    g529_p,
    g527_p_spl_,
    g524_p_spl_
  );


  or

  (
    g529_n,
    g527_n_spl_,
    g524_n_spl_
  );


  and

  (
    g530_p,
    g529_n,
    g528_n
  );


  or

  (
    g530_n,
    g529_p,
    g528_p
  );


  and

  (
    g531_p,
    g530_p,
    g515_n
  );


  and

  (
    g532_p,
    g530_n,
    g515_p
  );


  or

  (
    g533_n,
    g532_p,
    g531_p
  );


  and

  (
    g534_p,
    g408_p_spl_0,
    g400_p_spl_00
  );


  or

  (
    g534_n,
    g408_n_spl_00,
    g400_n_spl_00
  );


  and

  (
    g535_p,
    g534_n,
    g406_n_spl_0
  );


  or

  (
    g535_n,
    g534_p,
    g406_p_spl_0
  );


  and

  (
    g536_p,
    g535_n_spl_0,
    g415_p_spl_00
  );


  or

  (
    g536_n,
    g535_p_spl_0,
    g415_n_spl_00
  );


  and

  (
    g537_p,
    g536_n,
    g413_n_spl_
  );


  or

  (
    g537_n,
    g536_p,
    g413_p_spl_
  );


  and

  (
    g538_p,
    g537_n_spl_00,
    g422_p_spl_00
  );


  or

  (
    g538_n,
    g537_p_spl_00,
    g422_n_spl_00
  );


  and

  (
    g539_p,
    g538_n,
    g420_n_spl_0
  );


  or

  (
    g539_n,
    g538_p,
    g420_p_spl_0
  );


  and

  (
    g540_p,
    g539_n_spl_0,
    g429_p_spl_00
  );


  or

  (
    g540_n,
    g539_p_spl_0,
    g429_n_spl_00
  );


  and

  (
    g541_p,
    g540_n,
    g427_n_spl_
  );


  or

  (
    g541_n,
    g540_p,
    g427_p_spl_
  );


  or

  (
    g542_n,
    g541_p_spl_00,
    g396_n_spl_
  );


  and

  (
    g543_p,
    g381_p_spl_00,
    g373_p_spl_0
  );


  or

  (
    g543_n,
    g381_n_spl_00,
    g373_n_spl_0
  );


  and

  (
    g544_p,
    g543_n,
    g379_n_spl_
  );


  or

  (
    g544_n,
    g543_p,
    g379_p_spl_
  );


  and

  (
    g545_p,
    g544_n_spl_0,
    g387_n_spl_
  );


  or

  (
    g545_n,
    g544_p_spl_0,
    g387_p_spl_
  );


  and

  (
    g546_p,
    g545_n_spl_,
    g386_n_spl_
  );


  or

  (
    g546_n,
    g545_p_spl_,
    g386_p_spl_
  );


  or

  (
    g547_n,
    g546_p_spl_0,
    g395_n_spl_00
  );


  and

  (
    g548_p,
    g547_n,
    g542_n
  );


  and

  (
    g549_p,
    g548_p,
    g393_n_spl_
  );


  or

  (
    g550_n,
    g480_p_spl_0,
    g476_p_spl_00
  );


  or

  (
    g551_n,
    g464_p_spl_00,
    G21_n
  );


  or

  (
    g552_n,
    g464_n_spl_00,
    G21_p
  );


  and

  (
    g553_p,
    g552_n,
    g551_n
  );


  and

  (
    g554_p,
    g553_p_spl_,
    G177_p_spl_0000
  );


  or

  (
    g555_n,
    g554_p,
    G176_p_spl_00000
  );


  or

  (
    g556_n,
    g245_n_spl_0,
    G177_n_spl_0000
  );


  or

  (
    g557_n,
    g556_n,
    G176_n_spl_0000
  );


  or

  (
    g558_n,
    G177_p_spl_0000,
    G60_p
  );


  and

  (
    g559_p,
    g558_n,
    g557_n
  );


  and

  (
    g560_p,
    g559_p,
    g555_n
  );


  and

  (
    g561_p,
    g464_p_spl_01,
    g461_n_spl_0
  );


  or

  (
    g561_n,
    g464_n_spl_01,
    g461_p_spl_0
  );


  and

  (
    g562_p,
    g561_n,
    g465_n_spl_0
  );


  or

  (
    g562_n,
    g561_p,
    g465_p_spl_0
  );


  and

  (
    g563_p,
    g562_n_spl_0,
    G177_p_spl_0001
  );


  or

  (
    g564_n,
    g563_p,
    G176_p_spl_00000
  );


  or

  (
    g565_n,
    g224_n_spl_,
    G177_n_spl_0000
  );


  or

  (
    g566_n,
    g565_n,
    G176_n_spl_0000
  );


  or

  (
    g567_n,
    G177_p_spl_0001,
    G58_p
  );


  and

  (
    g568_p,
    g567_n,
    g566_n
  );


  and

  (
    g569_p,
    g568_p,
    g564_n
  );


  and

  (
    g570_p,
    g402_p_spl_0,
    G2_p_spl_0
  );


  or

  (
    g570_n,
    g402_n_spl_0,
    G2_n_spl_0
  );


  or

  (
    g571_n,
    g402_p_spl_1,
    G2_p_spl_0
  );


  and

  (
    g572_p,
    g571_n,
    g570_n_spl_
  );


  and

  (
    g573_p,
    g572_p_spl_,
    G177_p_spl_0010
  );


  or

  (
    g574_n,
    g573_p,
    G176_p_spl_00001
  );


  or

  (
    g575_n,
    g308_n_spl_,
    G177_n_spl_0001
  );


  or

  (
    g576_n,
    g575_n,
    G176_n_spl_0001
  );


  or

  (
    g577_n,
    G177_p_spl_0010,
    G48_p
  );


  and

  (
    g578_p,
    g577_n,
    g576_n
  );


  and

  (
    g579_p,
    g578_p,
    g574_n
  );


  and

  (
    g580_p,
    g479_p_spl_00,
    g476_p_spl_0
  );


  or

  (
    g580_n,
    g479_n_spl_00,
    g476_n_spl_0
  );


  and

  (
    g581_p,
    g580_n,
    g480_n
  );


  or

  (
    g581_n,
    g580_p,
    g480_p_spl_
  );


  and

  (
    g582_p,
    G173_n_spl_0000,
    G22_p_spl_
  );


  and

  (
    g583_p,
    G173_p_spl_0000,
    G3_p_spl_
  );


  or

  (
    g584_n,
    g583_p,
    g582_p
  );


  and

  (
    g585_p,
    g584_n,
    G172_n_spl_000
  );


  or

  (
    g586_n,
    g579_p_spl_00,
    G173_p_spl_0000
  );


  or

  (
    g587_n,
    g560_p_spl_00,
    G173_n_spl_0000
  );


  and

  (
    g588_p,
    g587_n,
    G172_p_spl_000
  );


  and

  (
    g589_p,
    g588_p,
    g586_n
  );


  or

  (
    g590_n,
    g589_p,
    g585_p
  );


  and

  (
    g591_p,
    G177_n_spl_0001,
    G19_p
  );


  and

  (
    g592_p,
    g591_p,
    G176_p_spl_00001
  );


  and

  (
    g593_p,
    g277_n_spl_,
    G176_p_spl_0001
  );


  and

  (
    g594_p,
    g471_p_spl_0,
    g459_p_spl_0
  );


  or

  (
    g594_n,
    g471_n_spl_00,
    g459_n_spl_0
  );


  and

  (
    g595_p,
    g594_n_spl_,
    g472_n_spl_
  );


  or

  (
    g595_n,
    g594_p_spl_,
    g472_p_spl_
  );


  and

  (
    g596_p,
    g595_p,
    g469_n_spl_0
  );


  or

  (
    g596_n,
    g595_n_spl_,
    g469_p_spl_0
  );


  and

  (
    g597_p,
    g596_n_spl_0,
    g454_p_spl_0
  );


  or

  (
    g597_n,
    g596_p_spl_0,
    g454_n_spl_00
  );


  and

  (
    g598_p,
    g597_n,
    g452_n_spl_0
  );


  or

  (
    g598_n,
    g597_p_spl_,
    g452_p_spl_0
  );


  or

  (
    g599_n,
    g598_p_spl_0,
    g450_p_spl_0
  );


  or

  (
    g600_n,
    g598_n_spl_0,
    g450_n_spl_0
  );


  and

  (
    g601_p,
    g600_n,
    g599_n
  );


  and

  (
    g602_p,
    g601_p_spl_,
    G176_n_spl_0001
  );


  or

  (
    g603_n,
    g602_p,
    g593_p
  );


  and

  (
    g604_p,
    g603_n,
    G177_p_spl_0011
  );


  or

  (
    g605_n,
    g604_p,
    g592_p
  );


  and

  (
    g606_p,
    G177_n_spl_0010,
    G59_p
  );


  and

  (
    g607_p,
    g606_p,
    G176_p_spl_0001
  );


  and

  (
    g608_p,
    g248_n_spl_,
    G176_p_spl_0010
  );


  and

  (
    g609_p,
    g596_p_spl_0,
    g454_n_spl_0
  );


  or

  (
    g610_n,
    g609_p,
    g597_p_spl_
  );


  and

  (
    g611_p,
    g610_n_spl_,
    G176_n_spl_0010
  );


  or

  (
    g612_n,
    g611_p,
    g608_p
  );


  and

  (
    g613_p,
    g612_n,
    G177_p_spl_0011
  );


  or

  (
    g614_n,
    g613_p,
    g607_p
  );


  and

  (
    g615_p,
    G177_n_spl_0010,
    G50_p
  );


  and

  (
    g616_p,
    g615_p,
    G176_p_spl_0010
  );


  and

  (
    g617_p,
    g465_n_spl_,
    g459_n_spl_
  );


  or

  (
    g617_n,
    g465_p_spl_,
    g459_p_spl_
  );


  and

  (
    g618_p,
    g617_p_spl_0,
    g471_n_spl_0
  );


  or

  (
    g619_n,
    g618_p,
    g595_n_spl_
  );


  or

  (
    g620_n,
    g619_n_spl_,
    G176_p_spl_0011
  );


  or

  (
    g621_n,
    g233_n_spl_,
    G176_n_spl_0010
  );


  and

  (
    g622_p,
    g621_n,
    G177_p_spl_0100
  );


  and

  (
    g623_p,
    g622_p,
    g620_n
  );


  or

  (
    g624_n,
    g623_p,
    g616_p
  );


  and

  (
    g625_p,
    G174_n_spl_0000,
    G22_p_spl_
  );


  and

  (
    g626_p,
    G174_p_spl_0000,
    G3_p_spl_
  );


  or

  (
    g627_n,
    g626_p,
    g625_p
  );


  and

  (
    g628_p,
    g627_n,
    G175_n_spl_000
  );


  or

  (
    g629_n,
    g579_p_spl_00,
    G174_p_spl_0000
  );


  or

  (
    g630_n,
    g560_p_spl_00,
    G174_n_spl_0000
  );


  and

  (
    g631_p,
    g630_n,
    G175_p_spl_000
  );


  and

  (
    g632_p,
    g631_p,
    g629_n
  );


  or

  (
    g633_n,
    g632_p,
    g628_p
  );


  and

  (
    g634_p,
    G177_n_spl_0011,
    G53_p
  );


  and

  (
    g635_p,
    g634_p,
    G176_p_spl_0011
  );


  or

  (
    g636_n,
    g356_n_spl_,
    G176_n_spl_0011
  );


  and

  (
    g637_p,
    g416_p_spl_0,
    G2_p_spl_1
  );


  or

  (
    g637_n,
    g416_n_spl_0,
    G2_n_spl_0
  );


  and

  (
    g638_p,
    g637_n,
    g537_p_spl_00
  );


  or

  (
    g638_n,
    g637_p,
    g537_n_spl_00
  );


  and

  (
    g639_p,
    g638_n,
    g422_p_spl_0
  );


  or

  (
    g639_n,
    g638_p_spl_,
    g422_n_spl_01
  );


  and

  (
    g640_p,
    g639_n,
    g420_n_spl_
  );


  or

  (
    g640_n,
    g639_p_spl_,
    g420_p_spl_
  );


  and

  (
    g641_p,
    g640_p,
    g429_n_spl_01
  );


  and

  (
    g642_p,
    g640_n,
    g429_p_spl_01
  );


  or

  (
    g643_n,
    g642_p,
    g641_p
  );


  or

  (
    g644_n,
    g643_n_spl_,
    G176_p_spl_0100
  );


  and

  (
    g645_p,
    g644_n,
    G177_p_spl_0100
  );


  and

  (
    g646_p,
    g645_p,
    g636_n
  );


  or

  (
    g647_n,
    g646_p,
    g635_p
  );


  and

  (
    g648_p,
    G177_n_spl_0011,
    G57_p
  );


  and

  (
    g649_p,
    g648_p,
    G176_p_spl_0100
  );


  and

  (
    g650_p,
    g365_n_spl_,
    G176_p_spl_0101
  );


  and

  (
    g651_p,
    g638_p_spl_,
    g422_n_spl_01
  );


  or

  (
    g652_n,
    g651_p,
    g639_p_spl_
  );


  and

  (
    g653_p,
    g652_n_spl_,
    G176_n_spl_0011
  );


  or

  (
    g654_n,
    g653_p,
    g650_p
  );


  and

  (
    g655_p,
    g654_n,
    G177_p_spl_0101
  );


  or

  (
    g656_n,
    g655_p,
    g649_p
  );


  and

  (
    g657_p,
    G177_n_spl_010,
    G56_p
  );


  and

  (
    g658_p,
    g657_p,
    G176_p_spl_0101
  );


  and

  (
    g659_p,
    g570_n_spl_,
    g400_n_spl_0
  );


  or

  (
    g659_n,
    g570_p,
    g400_p_spl_0
  );


  and

  (
    g660_p,
    g659_n,
    g408_p_spl_1
  );


  or

  (
    g660_n,
    g659_p_spl_,
    g408_n_spl_0
  );


  and

  (
    g661_p,
    g660_n,
    g406_n_spl_
  );


  or

  (
    g661_n,
    g660_p_spl_,
    g406_p_spl_
  );


  and

  (
    g662_p,
    g661_p,
    g415_n_spl_0
  );


  and

  (
    g663_p,
    g661_n,
    g415_p_spl_0
  );


  or

  (
    g664_n,
    g663_p,
    g662_p
  );


  or

  (
    g665_n,
    g664_n_spl_,
    G176_p_spl_0110
  );


  or

  (
    g666_n,
    g298_n_spl_,
    G176_n_spl_0100
  );


  and

  (
    g667_p,
    g666_n,
    G177_p_spl_0101
  );


  and

  (
    g668_p,
    g667_p,
    g665_n
  );


  or

  (
    g669_n,
    g668_p,
    g658_p
  );


  and

  (
    g670_p,
    G177_n_spl_010,
    G55_p
  );


  and

  (
    g671_p,
    g670_p,
    G176_p_spl_0110
  );


  and

  (
    g672_p,
    g659_p_spl_,
    g408_n_spl_1
  );


  or

  (
    g673_n,
    g672_p,
    g660_p_spl_
  );


  or

  (
    g674_n,
    g673_n_spl_,
    G176_p_spl_0111
  );


  or

  (
    g675_n,
    g289_n_spl_,
    G176_n_spl_0100
  );


  and

  (
    g676_p,
    g675_n,
    G177_p_spl_0110
  );


  and

  (
    g677_p,
    g676_p,
    g674_n
  );


  or

  (
    g678_n,
    g677_p,
    g671_p
  );


  and

  (
    g679_p,
    g440_n_spl_1,
    g434_n_spl_1
  );


  or

  (
    g679_n,
    g440_p_spl_1,
    g434_p_spl_1
  );


  and

  (
    g680_p,
    g440_p_spl_1,
    g434_p_spl_1
  );


  or

  (
    g680_n,
    g440_n_spl_1,
    g434_n_spl_1
  );


  and

  (
    g681_p,
    g680_n,
    g679_n
  );


  or

  (
    g681_n,
    g680_p,
    g679_p
  );


  and

  (
    g682_p,
    g681_p_spl_,
    g581_n_spl_00
  );


  or

  (
    g682_n,
    g681_n_spl_,
    g581_p_spl_00
  );


  and

  (
    g683_p,
    g681_n_spl_,
    g581_p_spl_00
  );


  or

  (
    g683_n,
    g681_p_spl_,
    g581_n_spl_00
  );


  and

  (
    g684_p,
    g683_n,
    g682_n
  );


  or

  (
    g684_n,
    g683_p,
    g682_p
  );


  and

  (
    g685_p,
    G133_n,
    G123_n_spl_111
  );


  or

  (
    g685_n,
    G133_p,
    G123_p_spl_111
  );


  and

  (
    g686_p,
    G132_n_spl_,
    G123_p_spl_111
  );


  or

  (
    g686_n,
    G132_p_spl_,
    G123_n_spl_111
  );


  and

  (
    g687_p,
    g686_n,
    g685_n
  );


  or

  (
    g687_n,
    g686_p,
    g685_p
  );


  and

  (
    g688_p,
    g687_n_spl_,
    g464_n_spl_01
  );


  or

  (
    g688_n,
    g687_p_spl_,
    g464_p_spl_01
  );


  and

  (
    g689_p,
    g687_p_spl_,
    g464_p_spl_10
  );


  or

  (
    g689_n,
    g687_n_spl_,
    g464_n_spl_10
  );


  and

  (
    g690_p,
    g689_n,
    g688_n
  );


  or

  (
    g690_n,
    g689_p,
    g688_p
  );


  and

  (
    g691_p,
    g451_p_spl_1,
    g447_n_spl_1
  );


  or

  (
    g691_n,
    g451_n_spl_1,
    g447_p_spl_1
  );


  and

  (
    g692_p,
    g451_n_spl_1,
    g447_p_spl_1
  );


  or

  (
    g692_n,
    g451_p_spl_1,
    g447_n_spl_1
  );


  and

  (
    g693_p,
    g692_n,
    g691_n
  );


  or

  (
    g693_n,
    g692_p,
    g691_p
  );


  and

  (
    g694_p,
    g468_n_spl_1,
    g458_n_spl_1
  );


  or

  (
    g694_n,
    g468_p_spl_1,
    g458_p_spl_1
  );


  and

  (
    g695_p,
    g468_p_spl_1,
    g458_p_spl_1
  );


  or

  (
    g695_n,
    g468_n_spl_1,
    g458_n_spl_1
  );


  and

  (
    g696_p,
    g695_n,
    g694_n
  );


  or

  (
    g696_n,
    g695_p,
    g694_p
  );


  and

  (
    g697_p,
    g696_n_spl_,
    g693_n_spl_
  );


  or

  (
    g697_n,
    g696_p_spl_,
    g693_p_spl_
  );


  and

  (
    g698_p,
    g696_p_spl_,
    g693_p_spl_
  );


  or

  (
    g698_n,
    g696_n_spl_,
    g693_n_spl_
  );


  and

  (
    g699_p,
    g698_n,
    g697_n
  );


  or

  (
    g699_n,
    g698_p,
    g697_p
  );


  and

  (
    g700_p,
    g699_n_spl_,
    g690_p_spl_
  );


  or

  (
    g700_n,
    g699_p_spl_,
    g690_n_spl_
  );


  and

  (
    g701_p,
    g699_p_spl_,
    g690_n_spl_
  );


  or

  (
    g701_n,
    g699_n_spl_,
    g690_p_spl_
  );


  and

  (
    g702_p,
    g701_n,
    g700_n
  );


  or

  (
    g702_n,
    g701_p,
    g700_p
  );


  and

  (
    g703_p,
    g702_p,
    g684_n
  );


  and

  (
    g704_p,
    g702_n,
    g684_p
  );


  or

  (
    g705_n,
    g704_p,
    g703_p
  );


  and

  (
    g706_p,
    g405_n_spl_1,
    g399_n_spl_1
  );


  or

  (
    g706_n,
    g405_p_spl_1,
    g399_p_spl_1
  );


  and

  (
    g707_p,
    g405_p_spl_1,
    g399_p_spl_1
  );


  or

  (
    g707_n,
    g405_n_spl_1,
    g399_n_spl_1
  );


  and

  (
    g708_p,
    g707_n,
    g706_n
  );


  or

  (
    g708_n,
    g707_p,
    g706_p
  );


  and

  (
    g709_p,
    g419_n_spl_1,
    g412_n_spl_1
  );


  or

  (
    g709_n,
    g419_p_spl_1,
    g412_p_spl_1
  );


  and

  (
    g710_p,
    g419_p_spl_1,
    g412_p_spl_1
  );


  or

  (
    g710_n,
    g419_n_spl_1,
    g412_n_spl_1
  );


  and

  (
    g711_p,
    g710_n,
    g709_n
  );


  or

  (
    g711_n,
    g710_p,
    g709_p
  );


  and

  (
    g712_p,
    g711_n_spl_,
    g708_p_spl_
  );


  or

  (
    g712_n,
    g711_p_spl_,
    g708_n_spl_
  );


  and

  (
    g713_p,
    g711_p_spl_,
    g708_n_spl_
  );


  or

  (
    g713_n,
    g711_n_spl_,
    g708_p_spl_
  );


  and

  (
    g714_p,
    g713_n,
    g712_n
  );


  or

  (
    g714_n,
    g713_p,
    g712_p
  );


  and

  (
    g715_p,
    G124_n_spl_111,
    G112_n
  );


  or

  (
    g715_n,
    G124_p_spl_111,
    G112_p
  );


  and

  (
    g716_p,
    G124_p_spl_111,
    G111_n_spl_
  );


  or

  (
    g716_n,
    G124_n_spl_111,
    G111_p_spl_
  );


  and

  (
    g717_p,
    g716_n,
    g715_n
  );


  or

  (
    g717_n,
    g716_p,
    g715_p
  );


  and

  (
    g718_p,
    g717_n_spl_,
    g392_n_spl_1
  );


  or

  (
    g718_n,
    g717_p_spl_,
    g392_p_spl_1
  );


  and

  (
    g719_p,
    g717_p_spl_,
    g392_p_spl_1
  );


  or

  (
    g719_n,
    g717_n_spl_,
    g392_n_spl_1
  );


  and

  (
    g720_p,
    g719_n,
    g718_n
  );


  or

  (
    g720_n,
    g719_p,
    g718_p
  );


  and

  (
    g721_p,
    g426_n_spl_1,
    g372_n_spl_1
  );


  or

  (
    g721_n,
    g426_p_spl_1,
    g372_p_spl_1
  );


  and

  (
    g722_p,
    g426_p_spl_1,
    g372_p_spl_1
  );


  or

  (
    g722_n,
    g426_n_spl_1,
    g372_n_spl_1
  );


  and

  (
    g723_p,
    g722_n,
    g721_n
  );


  or

  (
    g723_n,
    g722_p,
    g721_p
  );


  and

  (
    g724_p,
    g723_n_spl_,
    g720_p_spl_
  );


  or

  (
    g724_n,
    g723_p_spl_,
    g720_n_spl_
  );


  and

  (
    g725_p,
    g723_p_spl_,
    g720_n_spl_
  );


  or

  (
    g725_n,
    g723_n_spl_,
    g720_p_spl_
  );


  and

  (
    g726_p,
    g725_n,
    g724_n
  );


  or

  (
    g726_n,
    g725_p,
    g724_p
  );


  and

  (
    g727_p,
    g385_n_spl_1,
    g378_n_spl_1
  );


  or

  (
    g727_n,
    g385_p_spl_1,
    g378_p_spl_1
  );


  and

  (
    g728_p,
    g385_p_spl_1,
    g378_p_spl_1
  );


  or

  (
    g728_n,
    g385_n_spl_1,
    g378_n_spl_1
  );


  and

  (
    g729_p,
    g728_n,
    g727_n
  );


  or

  (
    g729_n,
    g728_p,
    g727_p
  );


  and

  (
    g730_p,
    g729_n_spl_,
    g726_n_spl_
  );


  or

  (
    g730_n,
    g729_p_spl_,
    g726_p_spl_
  );


  and

  (
    g731_p,
    g729_p_spl_,
    g726_p_spl_
  );


  or

  (
    g731_n,
    g729_n_spl_,
    g726_n_spl_
  );


  and

  (
    g732_p,
    g731_n,
    g730_n
  );


  or

  (
    g732_n,
    g731_p,
    g730_p
  );


  and

  (
    g733_p,
    g732_p,
    g714_n
  );


  and

  (
    g734_p,
    g732_n,
    g714_p
  );


  or

  (
    g735_n,
    g734_p,
    g733_p
  );


  and

  (
    g736_p,
    g430_p_spl_0,
    G2_p_spl_1
  );


  or

  (
    g736_n,
    g430_n_spl_0,
    G2_n_spl_
  );


  and

  (
    g737_p,
    g736_n,
    g541_p_spl_00
  );


  or

  (
    g737_n,
    g736_p,
    g541_n_spl_0
  );


  and

  (
    g738_p,
    g737_p_spl_00,
    g373_p_spl_
  );


  or

  (
    g738_n,
    g737_n_spl_00,
    g373_n_spl_
  );


  and

  (
    g739_p,
    g737_n_spl_00,
    g374_p_spl_0
  );


  or

  (
    g739_n,
    g737_p_spl_00,
    g374_n_spl_0
  );


  and

  (
    g740_p,
    g739_n,
    g738_n
  );


  or

  (
    g740_n,
    g739_p,
    g738_p
  );


  or

  (
    g741_n,
    g740_p,
    g381_n_spl_01
  );


  or

  (
    g742_n,
    g740_n,
    g381_p_spl_01
  );


  and

  (
    g743_p,
    g742_n,
    g741_n
  );


  or

  (
    g744_n,
    g743_p_spl_,
    g664_n_spl_
  );


  or

  (
    g745_n,
    g737_p_spl_0,
    g375_n_spl_00
  );


  or

  (
    g746_n,
    g737_n_spl_0,
    g375_p_spl_00
  );


  and

  (
    g747_p,
    g746_n,
    g745_n
  );


  or

  (
    g748_n,
    g747_p_spl_,
    g572_p_spl_
  );


  or

  (
    g749_n,
    g748_n,
    g744_n
  );


  or

  (
    g750_n,
    g652_n_spl_,
    g643_n_spl_
  );


  and

  (
    g751_p,
    g737_n_spl_1,
    g382_p_spl_
  );


  or

  (
    g751_n,
    g737_p_spl_1,
    g382_n_spl_
  );


  and

  (
    g752_p,
    g751_n,
    g544_p_spl_0
  );


  or

  (
    g752_n,
    g751_p,
    g544_n_spl_0
  );


  or

  (
    g753_n,
    g752_n,
    g388_n_spl_00
  );


  or

  (
    g754_n,
    g752_p,
    g388_p_spl_00
  );


  and

  (
    g755_p,
    g754_n,
    g753_n
  );


  and

  (
    g756_p,
    g737_n_spl_1,
    g389_p_spl_
  );


  or

  (
    g756_n,
    g737_p_spl_1,
    g389_n_spl_0
  );


  and

  (
    g757_p,
    g756_n,
    g546_p_spl_0
  );


  or

  (
    g757_n,
    g756_p,
    g546_n_spl_0
  );


  or

  (
    g758_n,
    g757_n,
    g395_n_spl_01
  );


  or

  (
    g759_n,
    g757_p,
    g395_p_spl_00
  );


  and

  (
    g760_p,
    g759_n,
    g758_n
  );


  or

  (
    g761_n,
    g760_p_spl_,
    g755_p_spl_
  );


  or

  (
    g762_n,
    g761_n,
    g673_n_spl_
  );


  or

  (
    g763_n,
    g762_n,
    g750_n
  );


  or

  (
    g764_n,
    g763_n,
    g749_n
  );


  or

  (
    g765_n,
    g619_n_spl_,
    g601_p_spl_
  );


  or

  (
    g766_n,
    g581_n_spl_01,
    g553_p_spl_
  );


  or

  (
    g767_n,
    g766_n,
    g610_n_spl_
  );


  or

  (
    g768_n,
    g767_n,
    g765_n
  );


  and

  (
    g769_p,
    g594_n_spl_,
    g469_n_spl_
  );


  or

  (
    g769_n,
    g594_p_spl_,
    g469_p_spl_
  );


  and

  (
    g770_p,
    g769_n,
    g454_p_spl_1
  );


  or

  (
    g770_n,
    g769_p,
    g454_n_spl_1
  );


  and

  (
    g771_p,
    g770_n,
    g452_n_spl_
  );


  or

  (
    g771_n,
    g770_p,
    g452_p_spl_
  );


  and

  (
    g772_p,
    g771_n,
    g450_p_spl_1
  );


  or

  (
    g772_n,
    g771_p,
    g450_n_spl_1
  );


  and

  (
    g773_p,
    g772_n,
    g473_n
  );


  or

  (
    g773_n,
    g772_p,
    g473_p_spl_
  );


  and

  (
    g774_p,
    g773_p,
    g448_n_spl_
  );


  or

  (
    g774_n,
    g773_n,
    g448_p_spl_
  );


  or

  (
    g775_n,
    g774_p_spl_00,
    g443_n_spl_00
  );


  or

  (
    g776_n,
    g774_n_spl_00,
    g443_p_spl_00
  );


  and

  (
    g777_p,
    g776_n,
    g775_n
  );


  or

  (
    g778_n,
    g777_p_spl_,
    g562_n_spl_0
  );


  and

  (
    g779_p,
    g441_p_spl_00,
    g437_p_spl_00
  );


  or

  (
    g779_n,
    g441_n_spl_00,
    g437_n_spl_00
  );


  and

  (
    g780_p,
    g779_n,
    g435_n_spl_
  );


  or

  (
    g780_n,
    g779_p,
    g435_p_spl_
  );


  and

  (
    g781_p,
    g774_n_spl_00,
    g444_p_spl_0
  );


  or

  (
    g781_n,
    g774_p_spl_00,
    g444_n_spl_
  );


  and

  (
    g782_p,
    g781_n,
    g780_p_spl_0
  );


  or

  (
    g782_n,
    g781_p,
    g780_n_spl_0
  );


  or

  (
    g783_n,
    g782_n,
    g479_p_spl_01
  );


  or

  (
    g784_n,
    g782_p,
    g479_n_spl_01
  );


  and

  (
    g785_p,
    g784_n,
    g783_n
  );


  and

  (
    g786_p,
    g774_p_spl_01,
    g441_p_spl_0
  );


  or

  (
    g786_n,
    g774_n_spl_01,
    g441_n_spl_0
  );


  and

  (
    g787_p,
    g774_n_spl_01,
    g442_p_spl_0
  );


  or

  (
    g787_n,
    g774_p_spl_01,
    g442_n_spl_0
  );


  and

  (
    g788_p,
    g787_n,
    g786_n
  );


  or

  (
    g788_n,
    g787_p,
    g786_p
  );


  or

  (
    g789_n,
    g788_p,
    g437_n_spl_01
  );


  or

  (
    g790_n,
    g788_n,
    g437_p_spl_01
  );


  and

  (
    g791_p,
    g790_n,
    g789_n
  );


  or

  (
    g792_n,
    g791_p_spl_,
    g785_p_spl_
  );


  or

  (
    g793_n,
    g792_n,
    g778_n
  );


  or

  (
    g794_n,
    g793_n,
    g768_n
  );


  and

  (
    g795_p,
    G158_n_spl_0000,
    G81_p_spl_
  );


  and

  (
    g796_p,
    G158_p_spl_0000,
    G80_p_spl_
  );


  or

  (
    g797_n,
    g796_p,
    g795_p
  );


  and

  (
    g798_p,
    g797_n,
    G159_n_spl_000
  );


  and

  (
    g799_p,
    g560_p_spl_0,
    G158_p_spl_0000
  );


  and

  (
    g800_p,
    g579_p_spl_0,
    G158_n_spl_0000
  );


  or

  (
    g801_n,
    g800_p,
    g799_p
  );


  and

  (
    g802_p,
    g801_n,
    G159_p_spl_000
  );


  or

  (
    g803_n,
    g802_p,
    g798_p
  );


  and

  (
    g804_p,
    g803_n,
    G64_p_spl_0000
  );


  and

  (
    g805_p,
    G160_n_spl_0000,
    G81_p_spl_
  );


  and

  (
    g806_p,
    G160_p_spl_0000,
    G80_p_spl_
  );


  or

  (
    g807_n,
    g806_p,
    g805_p
  );


  and

  (
    g808_p,
    g807_n,
    G161_n_spl_000
  );


  and

  (
    g809_p,
    g560_p_spl_1,
    G160_p_spl_0000
  );


  and

  (
    g810_p,
    g579_p_spl_1,
    G160_n_spl_0000
  );


  or

  (
    g811_n,
    g810_p,
    g809_p
  );


  and

  (
    g812_p,
    g811_n,
    G161_p_spl_000
  );


  or

  (
    g813_n,
    g812_p,
    g808_p
  );


  and

  (
    g814_p,
    g813_n,
    G64_p_spl_0000
  );


  and

  (
    g815_p,
    G173_n_spl_0001,
    G14_p_spl_
  );


  and

  (
    g816_p,
    G173_p_spl_0001,
    G16_p_spl_
  );


  or

  (
    g817_n,
    g816_p,
    g815_p
  );


  and

  (
    g818_p,
    g817_n,
    G172_n_spl_000
  );


  or

  (
    g819_n,
    g647_n_spl_00,
    G173_p_spl_0001
  );


  or

  (
    g820_n,
    g605_n_spl_00,
    G173_n_spl_0001
  );


  and

  (
    g821_p,
    g820_n,
    G172_p_spl_000
  );


  and

  (
    g822_p,
    g821_p,
    g819_n
  );


  or

  (
    g823_n,
    g822_p,
    g818_p
  );


  and

  (
    g824_p,
    G173_n_spl_0010,
    G6_p_spl_
  );


  and

  (
    g825_p,
    G173_p_spl_0010,
    G27_p_spl_
  );


  or

  (
    g826_n,
    g825_p,
    g824_p
  );


  and

  (
    g827_p,
    g826_n,
    G172_n_spl_001
  );


  or

  (
    g828_n,
    g656_n_spl_00,
    G173_p_spl_0010
  );


  or

  (
    g829_n,
    g614_n_spl_00,
    G173_n_spl_0010
  );


  and

  (
    g830_p,
    g829_n,
    G172_p_spl_001
  );


  and

  (
    g831_p,
    g830_p,
    g828_n
  );


  or

  (
    g832_n,
    g831_p,
    g827_p
  );


  and

  (
    g833_p,
    G173_n_spl_0011,
    G5_p_spl_
  );


  and

  (
    g834_p,
    G173_p_spl_0011,
    G26_p_spl_
  );


  or

  (
    g835_n,
    g834_p,
    g833_p
  );


  and

  (
    g836_p,
    g835_n,
    G172_n_spl_001
  );


  or

  (
    g837_n,
    g669_n_spl_00,
    G173_p_spl_0011
  );


  or

  (
    g838_n,
    g624_n_spl_00,
    G173_n_spl_0011
  );


  and

  (
    g839_p,
    g838_n,
    G172_p_spl_001
  );


  and

  (
    g840_p,
    g839_p,
    g837_n
  );


  or

  (
    g841_n,
    g840_p,
    g836_p
  );


  and

  (
    g842_p,
    G173_n_spl_010,
    G25_p_spl_
  );


  and

  (
    g843_p,
    G173_p_spl_010,
    G24_p_spl_
  );


  or

  (
    g844_n,
    g843_p,
    g842_p
  );


  and

  (
    g845_p,
    g844_n,
    G172_n_spl_01
  );


  or

  (
    g846_n,
    g678_n_spl_00,
    G173_p_spl_010
  );


  or

  (
    g847_n,
    g569_p_spl_00,
    G173_n_spl_010
  );


  and

  (
    g848_p,
    g847_n,
    G172_p_spl_01
  );


  and

  (
    g849_p,
    g848_p,
    g846_n
  );


  or

  (
    g850_n,
    g849_p,
    g845_p
  );


  and

  (
    g851_p,
    G174_n_spl_0001,
    G14_p_spl_
  );


  and

  (
    g852_p,
    G174_p_spl_0001,
    G16_p_spl_
  );


  or

  (
    g853_n,
    g852_p,
    g851_p
  );


  and

  (
    g854_p,
    g853_n,
    G175_n_spl_000
  );


  or

  (
    g855_n,
    g647_n_spl_00,
    G174_p_spl_0001
  );


  or

  (
    g856_n,
    g605_n_spl_00,
    G174_n_spl_0001
  );


  and

  (
    g857_p,
    g856_n,
    G175_p_spl_000
  );


  and

  (
    g858_p,
    g857_p,
    g855_n
  );


  or

  (
    g859_n,
    g858_p,
    g854_p
  );


  and

  (
    g860_p,
    G174_n_spl_0010,
    G6_p_spl_
  );


  and

  (
    g861_p,
    G174_p_spl_0010,
    G27_p_spl_
  );


  or

  (
    g862_n,
    g861_p,
    g860_p
  );


  and

  (
    g863_p,
    g862_n,
    G175_n_spl_001
  );


  or

  (
    g864_n,
    g656_n_spl_00,
    G174_p_spl_0010
  );


  or

  (
    g865_n,
    g614_n_spl_00,
    G174_n_spl_0010
  );


  and

  (
    g866_p,
    g865_n,
    G175_p_spl_001
  );


  and

  (
    g867_p,
    g866_p,
    g864_n
  );


  or

  (
    g868_n,
    g867_p,
    g863_p
  );


  and

  (
    g869_p,
    G174_n_spl_0011,
    G5_p_spl_
  );


  and

  (
    g870_p,
    G174_p_spl_0011,
    G26_p_spl_
  );


  or

  (
    g871_n,
    g870_p,
    g869_p
  );


  and

  (
    g872_p,
    g871_n,
    G175_n_spl_001
  );


  or

  (
    g873_n,
    g669_n_spl_00,
    G174_p_spl_0011
  );


  or

  (
    g874_n,
    g624_n_spl_00,
    G174_n_spl_0011
  );


  and

  (
    g875_p,
    g874_n,
    G175_p_spl_001
  );


  and

  (
    g876_p,
    g875_p,
    g873_n
  );


  or

  (
    g877_n,
    g876_p,
    g872_p
  );


  and

  (
    g878_p,
    G174_n_spl_010,
    G25_p_spl_
  );


  and

  (
    g879_p,
    G174_p_spl_010,
    G24_p_spl_
  );


  or

  (
    g880_n,
    g879_p,
    g878_p
  );


  and

  (
    g881_p,
    g880_n,
    G175_n_spl_01
  );


  or

  (
    g882_n,
    g678_n_spl_00,
    G174_p_spl_010
  );


  or

  (
    g883_n,
    g569_p_spl_00,
    G174_n_spl_010
  );


  and

  (
    g884_p,
    g883_n,
    G175_p_spl_01
  );


  and

  (
    g885_p,
    g884_p,
    g882_n
  );


  or

  (
    g886_n,
    g885_p,
    g881_p
  );


  and

  (
    g887_p,
    G158_n_spl_0001,
    G76_p_spl_
  );


  and

  (
    g888_p,
    G158_p_spl_0001,
    G86_p_spl_
  );


  or

  (
    g889_n,
    g888_p,
    g887_p
  );


  and

  (
    g890_p,
    g889_n,
    G159_n_spl_000
  );


  and

  (
    g891_p,
    g605_n_spl_0,
    G158_p_spl_0001
  );


  and

  (
    g892_p,
    g647_n_spl_0,
    G158_n_spl_0001
  );


  or

  (
    g893_n,
    g892_p,
    g891_p
  );


  and

  (
    g894_p,
    g893_n,
    G159_p_spl_000
  );


  or

  (
    g895_n,
    g894_p,
    g890_p
  );


  and

  (
    g896_p,
    g895_n,
    G64_p_spl_0001
  );


  and

  (
    g897_p,
    G158_n_spl_0010,
    G72_p_spl_
  );


  and

  (
    g898_p,
    G158_p_spl_0010,
    G82_p_spl_
  );


  or

  (
    g899_n,
    g898_p,
    g897_p
  );


  and

  (
    g900_p,
    g899_n,
    G159_n_spl_001
  );


  and

  (
    g901_p,
    g569_p_spl_0,
    G158_p_spl_0010
  );


  and

  (
    g902_p,
    g678_n_spl_0,
    G158_n_spl_0010
  );


  or

  (
    g903_n,
    g902_p,
    g901_p
  );


  and

  (
    g904_p,
    g903_n,
    G159_p_spl_001
  );


  or

  (
    g905_n,
    g904_p,
    g900_p
  );


  and

  (
    g906_p,
    g905_n,
    G64_p_spl_0001
  );


  and

  (
    g907_p,
    G158_n_spl_0011,
    G70_p_spl_
  );


  and

  (
    g908_p,
    G158_p_spl_0011,
    G71_p_spl_
  );


  or

  (
    g909_n,
    g908_p,
    g907_p
  );


  and

  (
    g910_p,
    g909_n,
    G159_n_spl_001
  );


  and

  (
    g911_p,
    g624_n_spl_0,
    G158_p_spl_0011
  );


  and

  (
    g912_p,
    g669_n_spl_0,
    G158_n_spl_0011
  );


  or

  (
    g913_n,
    g912_p,
    g911_p
  );


  and

  (
    g914_p,
    g913_n,
    G159_p_spl_001
  );


  or

  (
    g915_n,
    g914_p,
    g910_p
  );


  and

  (
    g916_p,
    g915_n,
    G64_p_spl_0010
  );


  and

  (
    g917_p,
    G158_n_spl_010,
    G68_p_spl_
  );


  and

  (
    g918_p,
    G158_p_spl_010,
    G69_p_spl_
  );


  or

  (
    g919_n,
    g918_p,
    g917_p
  );


  and

  (
    g920_p,
    g919_n,
    G159_n_spl_01
  );


  and

  (
    g921_p,
    g614_n_spl_0,
    G158_p_spl_010
  );


  and

  (
    g922_p,
    g656_n_spl_0,
    G158_n_spl_010
  );


  or

  (
    g923_n,
    g922_p,
    g921_p
  );


  and

  (
    g924_p,
    g923_n,
    G159_p_spl_01
  );


  or

  (
    g925_n,
    g924_p,
    g920_p
  );


  and

  (
    g926_p,
    g925_n,
    G64_p_spl_0010
  );


  and

  (
    g927_p,
    G160_n_spl_0001,
    G76_p_spl_
  );


  and

  (
    g928_p,
    G160_p_spl_0001,
    G86_p_spl_
  );


  or

  (
    g929_n,
    g928_p,
    g927_p
  );


  and

  (
    g930_p,
    g929_n,
    G161_n_spl_000
  );


  and

  (
    g931_p,
    g605_n_spl_1,
    G160_p_spl_0001
  );


  and

  (
    g932_p,
    g647_n_spl_1,
    G160_n_spl_0001
  );


  or

  (
    g933_n,
    g932_p,
    g931_p
  );


  and

  (
    g934_p,
    g933_n,
    G161_p_spl_000
  );


  or

  (
    g935_n,
    g934_p,
    g930_p
  );


  and

  (
    g936_p,
    g935_n,
    G64_p_spl_001
  );


  and

  (
    g937_p,
    G160_n_spl_0010,
    G72_p_spl_
  );


  and

  (
    g938_p,
    G160_p_spl_0010,
    G82_p_spl_
  );


  or

  (
    g939_n,
    g938_p,
    g937_p
  );


  and

  (
    g940_p,
    g939_n,
    G161_n_spl_001
  );


  and

  (
    g941_p,
    g569_p_spl_1,
    G160_p_spl_0010
  );


  and

  (
    g942_p,
    g678_n_spl_1,
    G160_n_spl_0010
  );


  or

  (
    g943_n,
    g942_p,
    g941_p
  );


  and

  (
    g944_p,
    g943_n,
    G161_p_spl_001
  );


  or

  (
    g945_n,
    g944_p,
    g940_p
  );


  and

  (
    g946_p,
    g945_n,
    G64_p_spl_010
  );


  and

  (
    g947_p,
    G160_n_spl_0011,
    G70_p_spl_
  );


  and

  (
    g948_p,
    G160_p_spl_0011,
    G71_p_spl_
  );


  or

  (
    g949_n,
    g948_p,
    g947_p
  );


  and

  (
    g950_p,
    g949_n,
    G161_n_spl_001
  );


  and

  (
    g951_p,
    g624_n_spl_1,
    G160_p_spl_0011
  );


  and

  (
    g952_p,
    g669_n_spl_1,
    G160_n_spl_0011
  );


  or

  (
    g953_n,
    g952_p,
    g951_p
  );


  and

  (
    g954_p,
    g953_n,
    G161_p_spl_001
  );


  or

  (
    g955_n,
    g954_p,
    g950_p
  );


  and

  (
    g956_p,
    g955_n,
    G64_p_spl_010
  );


  and

  (
    g957_p,
    G160_n_spl_010,
    G68_p_spl_
  );


  and

  (
    g958_p,
    G160_p_spl_010,
    G69_p_spl_
  );


  or

  (
    g959_n,
    g958_p,
    g957_p
  );


  and

  (
    g960_p,
    g959_n,
    G161_n_spl_01
  );


  and

  (
    g961_p,
    g614_n_spl_1,
    G160_p_spl_010
  );


  and

  (
    g962_p,
    g656_n_spl_1,
    G160_n_spl_010
  );


  or

  (
    g963_n,
    g962_p,
    g961_p
  );


  and

  (
    g964_p,
    g963_n,
    G161_p_spl_01
  );


  or

  (
    g965_n,
    g964_p,
    g960_p
  );


  and

  (
    g966_p,
    g965_n,
    G64_p_spl_011
  );


  or

  (
    g967_n,
    G178_n,
    G62_n
  );


  and

  (
    g968_p,
    g581_n_spl_01,
    G171_p_spl_
  );


  and

  (
    g969_p,
    G171_n_spl_,
    G54_p_spl_
  );


  or

  (
    g970_n,
    g969_p,
    g968_p
  );


  and

  (
    g971_p,
    g970_n,
    G170_p
  );


  and

  (
    g972_p,
    g237_n_spl_0,
    G171_n_spl_
  );


  and

  (
    g973_p,
    g476_n_spl_1,
    G61_n_spl_
  );


  or

  (
    g973_n,
    g476_p_spl_1,
    G61_p_spl_
  );


  and

  (
    g974_p,
    g476_p_spl_1,
    G61_p_spl_
  );


  or

  (
    g974_n,
    g476_n_spl_1,
    G61_n_spl_
  );


  and

  (
    g975_p,
    g974_n,
    g973_n
  );


  or

  (
    g975_n,
    g974_p,
    g973_p
  );


  and

  (
    g976_p,
    g975_p_spl_,
    G171_p_spl_
  );


  or

  (
    g977_n,
    g976_p,
    g972_p
  );


  and

  (
    g978_p,
    g977_n,
    G170_n
  );


  or

  (
    g979_n,
    g978_p,
    g971_p
  );


  and

  (
    g980_p,
    g979_n,
    g967_n
  );


  and

  (
    g981_p,
    g975_n,
    g581_n_spl_10
  );


  and

  (
    g982_p,
    g975_p_spl_,
    g581_p_spl_01
  );


  or

  (
    g983_n,
    g982_p,
    g981_p
  );


  and

  (
    g984_p,
    g581_n_spl_10,
    G177_p_spl_0110
  );


  or

  (
    g985_n,
    g984_p,
    G176_p_spl_0111
  );


  or

  (
    g986_n,
    g237_n_spl_1,
    G177_n_spl_011
  );


  or

  (
    g987_n,
    g986_n,
    G176_n_spl_0101
  );


  or

  (
    g988_n,
    G177_p_spl_0111,
    G54_p_spl_
  );


  and

  (
    g989_p,
    g988_n,
    g987_n
  );


  and

  (
    g990_p,
    g989_p,
    g985_n
  );


  and

  (
    g991_p,
    G177_n_spl_011,
    G52_p
  );


  and

  (
    g992_p,
    g991_p,
    G176_p_spl_1000
  );


  or

  (
    g993_n,
    g785_p_spl_,
    G176_p_spl_1000
  );


  or

  (
    g994_n,
    g240_n_spl_0,
    G176_n_spl_0101
  );


  and

  (
    g995_p,
    g994_n,
    G177_p_spl_0111
  );


  and

  (
    g996_p,
    g995_p,
    g993_n
  );


  or

  (
    g997_n,
    g996_p,
    g992_p
  );


  and

  (
    g998_p,
    G177_n_spl_100,
    G47_p
  );


  and

  (
    g999_p,
    g998_p,
    G176_p_spl_1001
  );


  or

  (
    g1000_n,
    g791_p_spl_,
    G176_p_spl_1001
  );


  or

  (
    g1001_n,
    g267_n_spl_0,
    G176_n_spl_011
  );


  and

  (
    g1002_p,
    g1001_n,
    G177_p_spl_1000
  );


  and

  (
    g1003_p,
    g1002_p,
    g1000_n
  );


  or

  (
    g1004_n,
    g1003_p,
    g999_p
  );


  and

  (
    g1005_p,
    G177_n_spl_100,
    G43_p
  );


  and

  (
    g1006_p,
    g1005_p,
    G176_p_spl_1010
  );


  or

  (
    g1007_n,
    g258_n_spl_0,
    G176_n_spl_011
  );


  or

  (
    g1008_n,
    g777_p_spl_,
    G176_p_spl_1010
  );


  and

  (
    g1009_p,
    g1008_n,
    G177_p_spl_1000
  );


  and

  (
    g1010_p,
    g1009_p,
    g1007_n
  );


  or

  (
    g1011_n,
    g1010_p,
    g1006_p
  );


  or

  (
    g1012_n,
    g533_n_spl_,
    G99_n_spl_
  );


  or

  (
    g1013_n,
    g1012_n,
    g735_n_spl_
  );


  or

  (
    g1014_n,
    g184_n_spl_,
    G155_n_spl_
  );


  or

  (
    g1015_n,
    g1014_n,
    g179_n_spl_
  );


  or

  (
    g1016_n,
    g1015_n,
    g705_n_spl_
  );


  or

  (
    g1017_n,
    g1016_n,
    g506_n_spl_
  );


  or

  (
    g1018_n,
    g1017_n,
    g1013_n
  );


  and

  (
    g1019_p,
    G177_n_spl_101,
    G46_p
  );


  and

  (
    g1020_p,
    g1019_p,
    G176_p_spl_1011
  );


  or

  (
    g1021_n,
    g760_p_spl_,
    G176_p_spl_1011
  );


  or

  (
    g1022_n,
    g317_n_spl_0,
    G176_n_spl_100
  );


  and

  (
    g1023_p,
    g1022_n,
    G177_p_spl_1001
  );


  and

  (
    g1024_p,
    g1023_p,
    g1021_n
  );


  or

  (
    g1025_n,
    g1024_p,
    g1020_p
  );


  and

  (
    g1026_p,
    G177_n_spl_101,
    G45_p
  );


  and

  (
    g1027_p,
    g1026_p,
    G176_p_spl_1100
  );


  or

  (
    g1028_n,
    g755_p_spl_,
    G176_p_spl_1100
  );


  or

  (
    g1029_n,
    g328_n_spl_,
    G176_n_spl_100
  );


  and

  (
    g1030_p,
    g1029_n,
    G177_p_spl_1001
  );


  and

  (
    g1031_p,
    g1030_p,
    g1028_n
  );


  or

  (
    g1032_n,
    g1031_p,
    g1027_p
  );


  and

  (
    g1033_p,
    G177_n_spl_110,
    G20_p
  );


  and

  (
    g1034_p,
    g1033_p,
    G176_p_spl_1101
  );


  or

  (
    g1035_n,
    g743_p_spl_,
    G176_p_spl_1101
  );


  or

  (
    g1036_n,
    g337_n_spl_,
    G176_n_spl_101
  );


  and

  (
    g1037_p,
    g1036_n,
    G177_p_spl_101
  );


  and

  (
    g1038_p,
    g1037_p,
    g1035_n
  );


  or

  (
    g1039_n,
    g1038_p,
    g1034_p
  );


  and

  (
    g1040_p,
    G177_n_spl_110,
    G44_p
  );


  and

  (
    g1041_p,
    g1040_p,
    G176_p_spl_1110
  );


  or

  (
    g1042_n,
    g747_p_spl_,
    G176_p_spl_1110
  );


  or

  (
    g1043_n,
    g347_n_spl_,
    G176_n_spl_101
  );


  and

  (
    g1044_p,
    g1043_n,
    G177_p_spl_101
  );


  and

  (
    g1045_p,
    g1044_p,
    g1042_n
  );


  or

  (
    g1046_n,
    g1045_p,
    g1041_p
  );


  or

  (
    g1047_n,
    g1025_n_spl_00,
    G174_p_spl_011
  );


  or

  (
    g1048_n,
    g990_p_spl_00,
    G174_n_spl_011
  );


  and

  (
    g1049_p,
    g1048_n,
    G175_p_spl_01
  );


  and

  (
    g1050_p,
    g1049_p,
    g1047_n
  );


  and

  (
    g1051_p,
    G174_n_spl_011,
    G41_p_spl_
  );


  and

  (
    g1052_p,
    G174_p_spl_011,
    G42_p_spl_
  );


  or

  (
    g1053_n,
    g1052_p,
    g1051_p
  );


  and

  (
    g1054_p,
    g1053_n,
    G175_n_spl_01
  );


  or

  (
    g1055_n,
    g1054_p,
    g1050_p
  );


  or

  (
    g1056_n,
    g1025_n_spl_00,
    G173_p_spl_011
  );


  or

  (
    g1057_n,
    g990_p_spl_00,
    G173_n_spl_011
  );


  and

  (
    g1058_p,
    g1057_n,
    G172_p_spl_01
  );


  and

  (
    g1059_p,
    g1058_p,
    g1056_n
  );


  and

  (
    g1060_p,
    G173_n_spl_011,
    G41_p_spl_
  );


  and

  (
    g1061_p,
    G173_p_spl_011,
    G42_p_spl_
  );


  or

  (
    g1062_n,
    g1061_p,
    g1060_p
  );


  and

  (
    g1063_p,
    g1062_n,
    G172_n_spl_01
  );


  or

  (
    g1064_n,
    g1063_p,
    g1059_p
  );


  and

  (
    g1065_p,
    G173_n_spl_100,
    G18_p_spl_
  );


  and

  (
    g1066_p,
    G173_p_spl_100,
    G17_p_spl_
  );


  or

  (
    g1067_n,
    g1066_p,
    g1065_p
  );


  and

  (
    g1068_p,
    g1067_n,
    G172_n_spl_10
  );


  or

  (
    g1069_n,
    g1032_n_spl_00,
    G173_p_spl_100
  );


  or

  (
    g1070_n,
    g997_n_spl_00,
    G173_n_spl_100
  );


  and

  (
    g1071_p,
    g1070_n,
    G172_p_spl_10
  );


  and

  (
    g1072_p,
    g1071_p,
    g1069_n
  );


  or

  (
    g1073_n,
    g1072_p,
    g1068_p
  );


  and

  (
    g1074_p,
    G173_n_spl_101,
    G40_p_spl_
  );


  and

  (
    g1075_p,
    G173_p_spl_101,
    G39_p_spl_
  );


  or

  (
    g1076_n,
    g1075_p,
    g1074_p
  );


  and

  (
    g1077_p,
    g1076_n,
    G172_n_spl_10
  );


  or

  (
    g1078_n,
    g1039_n_spl_00,
    G173_p_spl_101
  );


  or

  (
    g1079_n,
    g1004_n_spl_00,
    G173_n_spl_101
  );


  and

  (
    g1080_p,
    g1079_n,
    G172_p_spl_10
  );


  and

  (
    g1081_p,
    g1080_p,
    g1078_n
  );


  or

  (
    g1082_n,
    g1081_p,
    g1077_p
  );


  and

  (
    g1083_p,
    G173_n_spl_110,
    G15_p_spl_
  );


  and

  (
    g1084_p,
    G173_p_spl_110,
    G36_p_spl_
  );


  or

  (
    g1085_n,
    g1084_p,
    g1083_p
  );


  and

  (
    g1086_p,
    g1085_n,
    G172_n_spl_11
  );


  or

  (
    g1087_n,
    g1046_n_spl_00,
    G173_p_spl_110
  );


  or

  (
    g1088_n,
    g1011_n_spl_00,
    G173_n_spl_110
  );


  and

  (
    g1089_p,
    g1088_n,
    G172_p_spl_11
  );


  and

  (
    g1090_p,
    g1089_p,
    g1087_n
  );


  or

  (
    g1091_n,
    g1090_p,
    g1086_p
  );


  and

  (
    g1092_p,
    G174_n_spl_100,
    G18_p_spl_
  );


  and

  (
    g1093_p,
    G174_p_spl_100,
    G17_p_spl_
  );


  or

  (
    g1094_n,
    g1093_p,
    g1092_p
  );


  and

  (
    g1095_p,
    g1094_n,
    G175_n_spl_10
  );


  or

  (
    g1096_n,
    g1032_n_spl_00,
    G174_p_spl_100
  );


  or

  (
    g1097_n,
    g997_n_spl_00,
    G174_n_spl_100
  );


  and

  (
    g1098_p,
    g1097_n,
    G175_p_spl_10
  );


  and

  (
    g1099_p,
    g1098_p,
    g1096_n
  );


  or

  (
    g1100_n,
    g1099_p,
    g1095_p
  );


  and

  (
    g1101_p,
    G174_n_spl_101,
    G40_p_spl_
  );


  and

  (
    g1102_p,
    G174_p_spl_101,
    G39_p_spl_
  );


  or

  (
    g1103_n,
    g1102_p,
    g1101_p
  );


  and

  (
    g1104_p,
    g1103_n,
    G175_n_spl_10
  );


  or

  (
    g1105_n,
    g1039_n_spl_00,
    G174_p_spl_101
  );


  or

  (
    g1106_n,
    g1004_n_spl_00,
    G174_n_spl_101
  );


  and

  (
    g1107_p,
    g1106_n,
    G175_p_spl_10
  );


  and

  (
    g1108_p,
    g1107_p,
    g1105_n
  );


  or

  (
    g1109_n,
    g1108_p,
    g1104_p
  );


  and

  (
    g1110_p,
    G174_n_spl_110,
    G15_p_spl_
  );


  and

  (
    g1111_p,
    G174_p_spl_110,
    G36_p_spl_
  );


  or

  (
    g1112_n,
    g1111_p,
    g1110_p
  );


  and

  (
    g1113_p,
    g1112_n,
    G175_n_spl_11
  );


  or

  (
    g1114_n,
    g1046_n_spl_00,
    G174_p_spl_110
  );


  or

  (
    g1115_n,
    g1011_n_spl_00,
    G174_n_spl_110
  );


  and

  (
    g1116_p,
    g1115_n,
    G175_p_spl_11
  );


  and

  (
    g1117_p,
    g1116_p,
    g1114_n
  );


  or

  (
    g1118_n,
    g1117_p,
    g1113_p
  );


  and

  (
    g1119_p,
    G158_n_spl_011,
    G77_p_spl_
  );


  and

  (
    g1120_p,
    G158_p_spl_011,
    G87_p_spl_
  );


  or

  (
    g1121_n,
    g1120_p,
    g1119_p
  );


  and

  (
    g1122_p,
    g1121_n,
    G159_n_spl_01
  );


  and

  (
    g1123_p,
    g1011_n_spl_0,
    G158_p_spl_011
  );


  and

  (
    g1124_p,
    g1046_n_spl_0,
    G158_n_spl_011
  );


  or

  (
    g1125_n,
    g1124_p,
    g1123_p
  );


  and

  (
    g1126_p,
    g1125_n,
    G159_p_spl_01
  );


  or

  (
    g1127_n,
    g1126_p,
    g1122_p
  );


  and

  (
    g1128_p,
    g1127_n,
    G64_p_spl_011
  );


  and

  (
    g1129_p,
    G158_n_spl_100,
    G75_p_spl_
  );


  and

  (
    g1130_p,
    G158_p_spl_100,
    G85_p_spl_
  );


  or

  (
    g1131_n,
    g1130_p,
    g1129_p
  );


  and

  (
    g1132_p,
    g1131_n,
    G159_n_spl_10
  );


  and

  (
    g1133_p,
    g1004_n_spl_0,
    G158_p_spl_100
  );


  and

  (
    g1134_p,
    g1039_n_spl_0,
    G158_n_spl_100
  );


  or

  (
    g1135_n,
    g1134_p,
    g1133_p
  );


  and

  (
    g1136_p,
    g1135_n,
    G159_p_spl_10
  );


  or

  (
    g1137_n,
    g1136_p,
    g1132_p
  );


  and

  (
    g1138_p,
    g1137_n,
    G64_p_spl_100
  );


  and

  (
    g1139_p,
    G158_n_spl_101,
    G74_p_spl_
  );


  and

  (
    g1140_p,
    G158_p_spl_101,
    G84_p_spl_
  );


  or

  (
    g1141_n,
    g1140_p,
    g1139_p
  );


  and

  (
    g1142_p,
    g1141_n,
    G159_n_spl_10
  );


  and

  (
    g1143_p,
    g997_n_spl_0,
    G158_p_spl_101
  );


  and

  (
    g1144_p,
    g1032_n_spl_0,
    G158_n_spl_101
  );


  or

  (
    g1145_n,
    g1144_p,
    g1143_p
  );


  and

  (
    g1146_p,
    g1145_n,
    G159_p_spl_10
  );


  or

  (
    g1147_n,
    g1146_p,
    g1142_p
  );


  and

  (
    g1148_p,
    g1147_n,
    G64_p_spl_100
  );


  or

  (
    g1149_n,
    g1025_n_spl_0,
    G158_p_spl_110
  );


  or

  (
    g1150_n,
    g990_p_spl_0,
    G158_n_spl_110
  );


  and

  (
    g1151_p,
    g1150_n,
    G159_p_spl_11
  );


  and

  (
    g1152_p,
    g1151_p,
    g1149_n
  );


  and

  (
    g1153_p,
    G158_n_spl_110,
    G73_p_spl_
  );


  and

  (
    g1154_p,
    G158_p_spl_110,
    G83_p_spl_
  );


  or

  (
    g1155_n,
    g1154_p,
    g1153_p
  );


  and

  (
    g1156_p,
    g1155_n,
    G159_n_spl_11
  );


  or

  (
    g1157_n,
    g1156_p,
    g1152_p
  );


  and

  (
    g1158_p,
    g1157_n,
    G64_p_spl_101
  );


  and

  (
    g1159_p,
    G160_n_spl_011,
    G77_p_spl_
  );


  and

  (
    g1160_p,
    G160_p_spl_011,
    G87_p_spl_
  );


  or

  (
    g1161_n,
    g1160_p,
    g1159_p
  );


  and

  (
    g1162_p,
    g1161_n,
    G161_n_spl_01
  );


  and

  (
    g1163_p,
    g1011_n_spl_1,
    G160_p_spl_011
  );


  and

  (
    g1164_p,
    g1046_n_spl_1,
    G160_n_spl_011
  );


  or

  (
    g1165_n,
    g1164_p,
    g1163_p
  );


  and

  (
    g1166_p,
    g1165_n,
    G161_p_spl_01
  );


  or

  (
    g1167_n,
    g1166_p,
    g1162_p
  );


  and

  (
    g1168_p,
    g1167_n,
    G64_p_spl_101
  );


  and

  (
    g1169_p,
    G160_n_spl_100,
    G75_p_spl_
  );


  and

  (
    g1170_p,
    G160_p_spl_100,
    G85_p_spl_
  );


  or

  (
    g1171_n,
    g1170_p,
    g1169_p
  );


  and

  (
    g1172_p,
    g1171_n,
    G161_n_spl_10
  );


  and

  (
    g1173_p,
    g1004_n_spl_1,
    G160_p_spl_100
  );


  and

  (
    g1174_p,
    g1039_n_spl_1,
    G160_n_spl_100
  );


  or

  (
    g1175_n,
    g1174_p,
    g1173_p
  );


  and

  (
    g1176_p,
    g1175_n,
    G161_p_spl_10
  );


  or

  (
    g1177_n,
    g1176_p,
    g1172_p
  );


  and

  (
    g1178_p,
    g1177_n,
    G64_p_spl_110
  );


  and

  (
    g1179_p,
    G160_n_spl_101,
    G74_p_spl_
  );


  and

  (
    g1180_p,
    G160_p_spl_101,
    G84_p_spl_
  );


  or

  (
    g1181_n,
    g1180_p,
    g1179_p
  );


  and

  (
    g1182_p,
    g1181_n,
    G161_n_spl_10
  );


  and

  (
    g1183_p,
    g997_n_spl_1,
    G160_p_spl_101
  );


  and

  (
    g1184_p,
    g1032_n_spl_1,
    G160_n_spl_101
  );


  or

  (
    g1185_n,
    g1184_p,
    g1183_p
  );


  and

  (
    g1186_p,
    g1185_n,
    G161_p_spl_10
  );


  or

  (
    g1187_n,
    g1186_p,
    g1182_p
  );


  and

  (
    g1188_p,
    g1187_n,
    G64_p_spl_110
  );


  or

  (
    g1189_n,
    g1025_n_spl_1,
    G160_p_spl_110
  );


  or

  (
    g1190_n,
    g990_p_spl_1,
    G160_n_spl_110
  );


  and

  (
    g1191_p,
    g1190_n,
    G161_p_spl_11
  );


  and

  (
    g1192_p,
    g1191_p,
    g1189_n
  );


  and

  (
    g1193_p,
    G160_n_spl_110,
    G73_p_spl_
  );


  and

  (
    g1194_p,
    G160_p_spl_110,
    G83_p_spl_
  );


  or

  (
    g1195_n,
    g1194_p,
    g1193_p
  );


  and

  (
    g1196_p,
    g1195_n,
    G161_n_spl_11
  );


  or

  (
    g1197_n,
    g1196_p,
    g1192_p
  );


  and

  (
    g1198_p,
    g1197_n,
    G64_p_spl_111
  );


  and

  (
    g1199_p,
    g267_n_spl_,
    g258_n_spl_
  );


  or

  (
    g1199_n,
    g267_p_spl_,
    g258_p_spl_
  );


  and

  (
    g1200_p,
    g1199_n,
    g268_n_spl_
  );


  or

  (
    g1200_n,
    g1199_p,
    g268_p
  );


  and

  (
    g1201_p,
    g240_n_spl_,
    g237_p_spl_
  );


  or

  (
    g1201_n,
    g240_p_spl_,
    g237_n_spl_1
  );


  and

  (
    g1202_p,
    g1201_n,
    g241_n_spl_
  );


  or

  (
    g1202_n,
    g1201_p,
    g241_p
  );


  and

  (
    g1203_p,
    g1202_n_spl_,
    g1200_p_spl_
  );


  or

  (
    g1203_n,
    g1202_p_spl_,
    g1200_n_spl_
  );


  and

  (
    g1204_p,
    g1202_p_spl_,
    g1200_n_spl_
  );


  or

  (
    g1204_n,
    g1202_n_spl_,
    g1200_p_spl_
  );


  and

  (
    g1205_p,
    g1204_n,
    g1203_n
  );


  or

  (
    g1205_n,
    g1204_p,
    g1203_p
  );


  and

  (
    g1206_p,
    G128_p_spl_10,
    G101_p_spl_010
  );


  or

  (
    g1206_n,
    G128_n_spl_10,
    G101_n_spl_010
  );


  and

  (
    g1207_p,
    G128_n_spl_10,
    G100_p_spl_010
  );


  or

  (
    g1207_n,
    G128_p_spl_10,
    G100_n_spl_010
  );


  and

  (
    g1208_p,
    g1207_n,
    g1206_n
  );


  or

  (
    g1208_n,
    g1207_p,
    g1206_p
  );


  and

  (
    g1209_p,
    g1208_n,
    G150_p_spl_1
  );


  or

  (
    g1209_n,
    g1208_p,
    G150_n_spl_1
  );


  and

  (
    g1210_p,
    G128_p_spl_11,
    G102_n_spl_010
  );


  or

  (
    g1210_n,
    G128_n_spl_11,
    G102_p_spl_010
  );


  and

  (
    g1211_p,
    G128_n_spl_11,
    G98_n_spl_010
  );


  or

  (
    g1211_n,
    G128_p_spl_11,
    G98_p_spl_010
  );


  and

  (
    g1212_p,
    g1211_n,
    g1210_n
  );


  or

  (
    g1212_n,
    g1211_p,
    g1210_p
  );


  and

  (
    g1213_p,
    g1212_n,
    G150_n_spl_1
  );


  or

  (
    g1213_n,
    g1212_p,
    G150_p_spl_1
  );


  and

  (
    g1214_p,
    g1213_n,
    g1209_n
  );


  or

  (
    g1214_n,
    g1213_p,
    g1209_p
  );


  and

  (
    g1215_p,
    G126_p_spl_10,
    G101_p_spl_011
  );


  or

  (
    g1215_n,
    G126_n_spl_10,
    G101_n_spl_011
  );


  and

  (
    g1216_p,
    G126_n_spl_10,
    G100_p_spl_010
  );


  or

  (
    g1216_n,
    G126_p_spl_10,
    G100_n_spl_010
  );


  and

  (
    g1217_p,
    g1216_n,
    g1215_n
  );


  or

  (
    g1217_n,
    g1216_p,
    g1215_p
  );


  and

  (
    g1218_p,
    g1217_n,
    G149_p_spl_1
  );


  or

  (
    g1218_n,
    g1217_p,
    G149_n_spl_1
  );


  and

  (
    g1219_p,
    G126_p_spl_11,
    G102_n_spl_010
  );


  or

  (
    g1219_n,
    G126_n_spl_11,
    G102_p_spl_010
  );


  and

  (
    g1220_p,
    G126_n_spl_11,
    G98_n_spl_010
  );


  or

  (
    g1220_n,
    G126_p_spl_11,
    G98_p_spl_010
  );


  and

  (
    g1221_p,
    g1220_n,
    g1219_n
  );


  or

  (
    g1221_n,
    g1220_p,
    g1219_p
  );


  and

  (
    g1222_p,
    g1221_n,
    G149_n_spl_1
  );


  or

  (
    g1222_n,
    g1221_p,
    G149_p_spl_1
  );


  and

  (
    g1223_p,
    g1222_n,
    g1218_n
  );


  or

  (
    g1223_n,
    g1222_p,
    g1218_p
  );


  and

  (
    g1224_p,
    g1223_p_spl_,
    g1214_n_spl_
  );


  or

  (
    g1224_n,
    g1223_n_spl_,
    g1214_p_spl_
  );


  and

  (
    g1225_p,
    g1223_n_spl_,
    g1214_p_spl_
  );


  or

  (
    g1225_n,
    g1223_p_spl_,
    g1214_n_spl_
  );


  and

  (
    g1226_p,
    g1225_n,
    g1224_n
  );


  or

  (
    g1226_n,
    g1225_p,
    g1224_p
  );


  and

  (
    g1227_p,
    G148_n_spl_1,
    G98_n_spl_011
  );


  or

  (
    g1227_n,
    G148_p_spl_1,
    G98_p_spl_011
  );


  and

  (
    g1228_p,
    G148_p_spl_1,
    G100_p_spl_011
  );


  or

  (
    g1228_n,
    G148_n_spl_1,
    G100_n_spl_011
  );


  and

  (
    g1229_p,
    g1228_n,
    g1227_n
  );


  or

  (
    g1229_n,
    g1228_p,
    g1227_p
  );


  and

  (
    g1230_p,
    G121_p_spl_10,
    G101_p_spl_011
  );


  or

  (
    g1230_n,
    G121_n_spl_10,
    G101_n_spl_011
  );


  and

  (
    g1231_p,
    G121_n_spl_10,
    G100_p_spl_011
  );


  or

  (
    g1231_n,
    G121_p_spl_10,
    G100_n_spl_011
  );


  and

  (
    g1232_p,
    g1231_n,
    g1230_n
  );


  or

  (
    g1232_n,
    g1231_p,
    g1230_p
  );


  and

  (
    g1233_p,
    g1232_n,
    G147_p_spl_1
  );


  or

  (
    g1233_n,
    g1232_p,
    G147_n_spl_1
  );


  and

  (
    g1234_p,
    G121_p_spl_11,
    G102_n_spl_011
  );


  or

  (
    g1234_n,
    G121_n_spl_11,
    G102_p_spl_011
  );


  and

  (
    g1235_p,
    G121_n_spl_11,
    G98_n_spl_011
  );


  or

  (
    g1235_n,
    G121_p_spl_11,
    G98_p_spl_011
  );


  and

  (
    g1236_p,
    g1235_n,
    g1234_n
  );


  or

  (
    g1236_n,
    g1235_p,
    g1234_p
  );


  and

  (
    g1237_p,
    g1236_n,
    G147_n_spl_1
  );


  or

  (
    g1237_n,
    g1236_p,
    G147_p_spl_1
  );


  and

  (
    g1238_p,
    g1237_n,
    g1233_n
  );


  or

  (
    g1238_n,
    g1237_p,
    g1233_p
  );


  and

  (
    g1239_p,
    g1238_p_spl_,
    g1229_n_spl_
  );


  or

  (
    g1239_n,
    g1238_n_spl_,
    g1229_p_spl_
  );


  and

  (
    g1240_p,
    g1238_n_spl_,
    g1229_p_spl_
  );


  or

  (
    g1240_n,
    g1238_p_spl_,
    g1229_n_spl_
  );


  and

  (
    g1241_p,
    g1240_n,
    g1239_n
  );


  or

  (
    g1241_n,
    g1240_p,
    g1239_p
  );


  and

  (
    g1242_p,
    g1241_p_spl_,
    g245_n_spl_1
  );


  or

  (
    g1242_n,
    g1241_n_spl_,
    g245_p_spl_
  );


  and

  (
    g1243_p,
    g1241_n_spl_,
    g245_p_spl_
  );


  or

  (
    g1243_n,
    g1241_p_spl_,
    g245_n_spl_1
  );


  and

  (
    g1244_p,
    g1243_n,
    g1242_n
  );


  or

  (
    g1244_n,
    g1243_p,
    g1242_p
  );


  and

  (
    g1245_p,
    g1244_n_spl_,
    g1226_p_spl_
  );


  or

  (
    g1245_n,
    g1244_p_spl_,
    g1226_n_spl_
  );


  and

  (
    g1246_p,
    g1244_p_spl_,
    g1226_n_spl_
  );


  or

  (
    g1246_n,
    g1244_n_spl_,
    g1226_p_spl_
  );


  and

  (
    g1247_p,
    g1246_n,
    g1245_n
  );


  or

  (
    g1247_n,
    g1246_p,
    g1245_p
  );


  or

  (
    g1248_n,
    g1247_n,
    g1205_p
  );


  or

  (
    g1249_n,
    g1247_p,
    g1205_n
  );


  and

  (
    g1250_p,
    g1249_n,
    g1248_n
  );


  or

  (
    g1251_n,
    g1250_p,
    G176_n_spl_110
  );


  and

  (
    g1252_p,
    g596_n_spl_0,
    g464_n_spl_10
  );


  or

  (
    g1252_n,
    g596_p_spl_1,
    g464_p_spl_10
  );


  and

  (
    g1253_p,
    g596_p_spl_1,
    g464_p_spl_1
  );


  or

  (
    g1253_n,
    g596_n_spl_,
    g464_n_spl_1
  );


  and

  (
    g1254_p,
    g1253_n,
    g1252_n
  );


  or

  (
    g1254_n,
    g1253_p,
    g1252_p
  );


  and

  (
    g1255_p,
    g1254_n_spl_,
    g617_p_spl_0
  );


  or

  (
    g1255_n,
    g1254_p_spl_,
    g617_n_spl_
  );


  and

  (
    g1256_p,
    g1254_p_spl_,
    g617_n_spl_
  );


  or

  (
    g1256_n,
    g1254_n_spl_,
    g617_p_spl_
  );


  and

  (
    g1257_p,
    g1256_n,
    g1255_n
  );


  or

  (
    g1257_n,
    g1256_p,
    g1255_p
  );


  and

  (
    g1258_p,
    g1257_p_spl_,
    g598_p_spl_0
  );


  or

  (
    g1258_n,
    g1257_n_spl_,
    g598_n_spl_0
  );


  and

  (
    g1259_p,
    g1257_n_spl_,
    g598_n_spl_
  );


  or

  (
    g1259_n,
    g1257_p_spl_,
    g598_p_spl_
  );


  and

  (
    g1260_p,
    g1259_n,
    g1258_n
  );


  or

  (
    g1260_n,
    g1259_p,
    g1258_p
  );


  and

  (
    g1261_p,
    g562_p,
    G162_n_spl_
  );


  or

  (
    g1261_n,
    g562_n_spl_,
    G162_p_spl_
  );


  and

  (
    g1262_p,
    g461_n_spl_,
    G162_p_spl_
  );


  or

  (
    g1262_n,
    g461_p_spl_,
    G162_n_spl_
  );


  and

  (
    g1263_p,
    g1262_n,
    g1261_n
  );


  or

  (
    g1263_n,
    g1262_p,
    g1261_p
  );


  and

  (
    g1264_p,
    g1263_p_spl_,
    g1260_p_spl_
  );


  or

  (
    g1264_n,
    g1263_n_spl_,
    g1260_n_spl_
  );


  and

  (
    g1265_p,
    g1263_n_spl_,
    g1260_n_spl_
  );


  or

  (
    g1265_n,
    g1263_p_spl_,
    g1260_p_spl_
  );


  and

  (
    g1266_p,
    g1265_n,
    g1264_n
  );


  or

  (
    g1266_n,
    g1265_p,
    g1264_p
  );


  and

  (
    g1267_p,
    g454_n_spl_1,
    g450_n_spl_1
  );


  or

  (
    g1267_n,
    g454_p_spl_1,
    g450_p_spl_1
  );


  and

  (
    g1268_p,
    g1267_n,
    g455_n_spl_
  );


  or

  (
    g1268_n,
    g1267_p,
    g455_p_spl_
  );


  and

  (
    g1269_p,
    g1268_n_spl_,
    g471_p_spl_1
  );


  or

  (
    g1269_n,
    g1268_p_spl_,
    g471_n_spl_1
  );


  and

  (
    g1270_p,
    g1268_p_spl_,
    g471_n_spl_1
  );


  or

  (
    g1270_n,
    g1268_n_spl_,
    g471_p_spl_1
  );


  and

  (
    g1271_p,
    g1270_n,
    g1269_n
  );


  or

  (
    g1271_n,
    g1270_p,
    g1269_p
  );


  and

  (
    g1272_p,
    g1271_n_spl_,
    g1266_n_spl_
  );


  or

  (
    g1272_n,
    g1271_p_spl_,
    g1266_p_spl_
  );


  and

  (
    g1273_p,
    g1271_p_spl_,
    g1266_p_spl_
  );


  or

  (
    g1273_n,
    g1271_n_spl_,
    g1266_n_spl_
  );


  and

  (
    g1274_p,
    g1273_n,
    g1272_n
  );


  or

  (
    g1274_n,
    g1273_p,
    g1272_p
  );


  and

  (
    g1275_p,
    g780_p_spl_0,
    g444_n_spl_
  );


  or

  (
    g1275_n,
    g780_n_spl_0,
    g444_p_spl_
  );


  and

  (
    g1276_p,
    g1275_n_spl_,
    g442_n_spl_1
  );


  or

  (
    g1276_n,
    g1275_p_spl_,
    g442_p_spl_1
  );


  and

  (
    g1277_p,
    g1275_p_spl_,
    g442_p_spl_1
  );


  or

  (
    g1277_n,
    g1275_n_spl_,
    g442_n_spl_1
  );


  and

  (
    g1278_p,
    g1277_n,
    g1276_n
  );


  or

  (
    g1278_n,
    g1277_p,
    g1276_p
  );


  and

  (
    g1279_p,
    g1278_p_spl_,
    g479_n_spl_01
  );


  or

  (
    g1279_n,
    g1278_n_spl_,
    g479_p_spl_01
  );


  and

  (
    g1280_p,
    g1278_n_spl_,
    g479_p_spl_10
  );


  or

  (
    g1280_n,
    g1278_p_spl_,
    g479_n_spl_10
  );


  and

  (
    g1281_p,
    g1280_n,
    g1279_n
  );


  or

  (
    g1281_n,
    g1280_p,
    g1279_p
  );


  and

  (
    g1282_p,
    g1281_p_spl_,
    g443_n_spl_0
  );


  or

  (
    g1282_n,
    g1281_n_spl_,
    g443_p_spl_0
  );


  and

  (
    g1283_p,
    g1281_n_spl_,
    g443_p_spl_1
  );


  or

  (
    g1283_n,
    g1281_p_spl_,
    g443_n_spl_1
  );


  and

  (
    g1284_p,
    g1283_n,
    g1282_n_spl_
  );


  or

  (
    g1284_n,
    g1283_p,
    g1282_p_spl_
  );


  and

  (
    g1285_p,
    g1284_n_spl_,
    g437_p_spl_01
  );


  or

  (
    g1285_n,
    g1284_p_spl_,
    g437_n_spl_01
  );


  and

  (
    g1286_p,
    g780_n_spl_1,
    g441_p_spl_1
  );


  or

  (
    g1286_n,
    g780_p_spl_1,
    g441_n_spl_1
  );


  and

  (
    g1287_p,
    g780_p_spl_1,
    g441_n_spl_1
  );


  or

  (
    g1287_n,
    g780_n_spl_1,
    g441_p_spl_1
  );


  and

  (
    g1288_p,
    g1287_n,
    g1286_n
  );


  or

  (
    g1288_n,
    g1287_p,
    g1286_p
  );


  and

  (
    g1289_p,
    g1288_n_spl_,
    g479_p_spl_10
  );


  or

  (
    g1289_n,
    g1288_p_spl_,
    g479_n_spl_10
  );


  and

  (
    g1290_p,
    g1288_p_spl_,
    g479_n_spl_1
  );


  or

  (
    g1290_n,
    g1288_n_spl_,
    g479_p_spl_1
  );


  and

  (
    g1291_p,
    g1290_n,
    g1289_n
  );


  or

  (
    g1291_n,
    g1290_p,
    g1289_p
  );


  and

  (
    g1292_p,
    g1291_n,
    g443_p_spl_1
  );


  or

  (
    g1292_n,
    g1291_p,
    g443_n_spl_1
  );


  and

  (
    g1293_p,
    g1292_n,
    g437_n_spl_1
  );


  or

  (
    g1293_n,
    g1292_p,
    g437_p_spl_1
  );


  and

  (
    g1294_p,
    g1293_p,
    g1282_n_spl_
  );


  or

  (
    g1294_n,
    g1293_n,
    g1282_p_spl_
  );


  and

  (
    g1295_p,
    g1294_p,
    g774_p_spl_1
  );


  or

  (
    g1295_n,
    g1294_n,
    g774_n_spl_1
  );


  and

  (
    g1296_p,
    g1295_n,
    g1285_n
  );


  or

  (
    g1296_n,
    g1295_p,
    g1285_p
  );


  and

  (
    g1297_p,
    g774_n_spl_1,
    g437_n_spl_1
  );


  or

  (
    g1297_n,
    g774_p_spl_1,
    g437_p_spl_1
  );


  and

  (
    g1298_p,
    g1297_p,
    g1284_p_spl_
  );


  or

  (
    g1298_n,
    g1297_n,
    g1284_n_spl_
  );


  and

  (
    g1299_p,
    g1298_n,
    g1296_p
  );


  or

  (
    g1299_n,
    g1298_p,
    g1296_n
  );


  and

  (
    g1300_p,
    g1299_p_spl_,
    g581_p_spl_01
  );


  or

  (
    g1300_n,
    g1299_n_spl_,
    g581_n_spl_11
  );


  and

  (
    g1301_p,
    g1299_n_spl_,
    g581_n_spl_11
  );


  or

  (
    g1301_n,
    g1299_p_spl_,
    g581_p_spl_1
  );


  and

  (
    g1302_p,
    g1301_n,
    g1300_n
  );


  or

  (
    g1302_n,
    g1301_p,
    g1300_p
  );


  and

  (
    g1303_p,
    g1302_n,
    g1274_p
  );


  and

  (
    g1304_p,
    g1302_p,
    g1274_n
  );


  or

  (
    g1305_n,
    g1304_p,
    G176_p_spl_1111
  );


  or

  (
    g1306_n,
    g1305_n,
    g1303_p
  );


  and

  (
    g1307_p,
    g1306_n,
    g1251_n
  );


  or

  (
    g1308_n,
    g1307_p,
    G177_n_spl_111
  );


  or

  (
    g1309_n,
    G177_p_spl_110,
    G51_p
  );


  or

  (
    g1310_n,
    g1309_n,
    G176_n_spl_110
  );


  and

  (
    g1311_p,
    g1310_n,
    g1308_n_spl_
  );


  and

  (
    g1312_p,
    G101_p_spl_100,
    G94_p_spl_10
  );


  or

  (
    g1312_n,
    G101_n_spl_100,
    G94_n_spl_10
  );


  and

  (
    g1313_p,
    G100_p_spl_100,
    G94_n_spl_10
  );


  or

  (
    g1313_n,
    G100_n_spl_100,
    G94_p_spl_10
  );


  and

  (
    g1314_p,
    g1313_n,
    g1312_n
  );


  or

  (
    g1314_n,
    g1313_p,
    g1312_p
  );


  and

  (
    g1315_p,
    g1314_n,
    G140_p_spl_1
  );


  or

  (
    g1315_n,
    g1314_p,
    G140_n_spl_1
  );


  and

  (
    g1316_p,
    G102_n_spl_011,
    G94_p_spl_11
  );


  or

  (
    g1316_n,
    G102_p_spl_011,
    G94_n_spl_11
  );


  and

  (
    g1317_p,
    G98_n_spl_100,
    G94_n_spl_11
  );


  or

  (
    g1317_n,
    G98_p_spl_100,
    G94_p_spl_11
  );


  and

  (
    g1318_p,
    g1317_n,
    g1316_n
  );


  or

  (
    g1318_n,
    g1317_p,
    g1316_p
  );


  and

  (
    g1319_p,
    g1318_n,
    G140_n_spl_1
  );


  or

  (
    g1319_n,
    g1318_p,
    G140_p_spl_1
  );


  and

  (
    g1320_p,
    g1319_n,
    g1315_n
  );


  or

  (
    g1320_n,
    g1319_p,
    g1315_p
  );


  and

  (
    g1321_p,
    G101_p_spl_100,
    G92_p_spl_10
  );


  or

  (
    g1321_n,
    G101_n_spl_100,
    G92_n_spl_10
  );


  and

  (
    g1322_p,
    G100_p_spl_100,
    G92_n_spl_10
  );


  or

  (
    g1322_n,
    G100_n_spl_100,
    G92_p_spl_10
  );


  and

  (
    g1323_p,
    g1322_n,
    g1321_n
  );


  or

  (
    g1323_n,
    g1322_p,
    g1321_p
  );


  and

  (
    g1324_p,
    g1323_n,
    G144_p_spl_1
  );


  or

  (
    g1324_n,
    g1323_p,
    G144_n_spl_1
  );


  and

  (
    g1325_p,
    G102_n_spl_100,
    G92_p_spl_11
  );


  or

  (
    g1325_n,
    G102_p_spl_100,
    G92_n_spl_11
  );


  and

  (
    g1326_p,
    G98_n_spl_100,
    G92_n_spl_11
  );


  or

  (
    g1326_n,
    G98_p_spl_100,
    G92_p_spl_11
  );


  and

  (
    g1327_p,
    g1326_n,
    g1325_n
  );


  or

  (
    g1327_n,
    g1326_p,
    g1325_p
  );


  and

  (
    g1328_p,
    g1327_n,
    G144_n_spl_1
  );


  or

  (
    g1328_n,
    g1327_p,
    G144_p_spl_1
  );


  and

  (
    g1329_p,
    g1328_n,
    g1324_n
  );


  or

  (
    g1329_n,
    g1328_p,
    g1324_p
  );


  and

  (
    g1330_p,
    g1329_p_spl_,
    g1320_n_spl_
  );


  or

  (
    g1330_n,
    g1329_n_spl_,
    g1320_p_spl_
  );


  and

  (
    g1331_p,
    g1329_n_spl_,
    g1320_p_spl_
  );


  or

  (
    g1331_n,
    g1329_p_spl_,
    g1320_n_spl_
  );


  and

  (
    g1332_p,
    g1331_n,
    g1330_n
  );


  or

  (
    g1332_n,
    g1331_p,
    g1330_p
  );


  and

  (
    g1333_p,
    G101_p_spl_101,
    G90_p_spl_10
  );


  or

  (
    g1333_n,
    G101_n_spl_101,
    G90_n_spl_10
  );


  and

  (
    g1334_p,
    G100_p_spl_101,
    G90_n_spl_10
  );


  or

  (
    g1334_n,
    G100_n_spl_101,
    G90_p_spl_10
  );


  and

  (
    g1335_p,
    g1334_n,
    g1333_n
  );


  or

  (
    g1335_n,
    g1334_p,
    g1333_p
  );


  and

  (
    g1336_p,
    g1335_n,
    G143_p_spl_1
  );


  or

  (
    g1336_n,
    g1335_p,
    G143_n_spl_1
  );


  and

  (
    g1337_p,
    G102_n_spl_100,
    G90_p_spl_11
  );


  or

  (
    g1337_n,
    G102_p_spl_100,
    G90_n_spl_11
  );


  and

  (
    g1338_p,
    G98_n_spl_101,
    G90_n_spl_11
  );


  or

  (
    g1338_n,
    G98_p_spl_101,
    G90_p_spl_11
  );


  and

  (
    g1339_p,
    g1338_n,
    g1337_n
  );


  or

  (
    g1339_n,
    g1338_p,
    g1337_p
  );


  and

  (
    g1340_p,
    g1339_n,
    G143_n_spl_1
  );


  or

  (
    g1340_n,
    g1339_p,
    G143_p_spl_1
  );


  and

  (
    g1341_p,
    g1340_n,
    g1336_n
  );


  or

  (
    g1341_n,
    g1340_p,
    g1336_p
  );


  and

  (
    g1342_p,
    g1341_n_spl_,
    g317_n_spl_1
  );


  or

  (
    g1342_n,
    g1341_p_spl_,
    g317_p_spl_
  );


  and

  (
    g1343_p,
    g1341_p_spl_,
    g317_p_spl_
  );


  or

  (
    g1343_n,
    g1341_n_spl_,
    g317_n_spl_1
  );


  and

  (
    g1344_p,
    g1343_n,
    g1342_n
  );


  or

  (
    g1344_n,
    g1343_p,
    g1342_p
  );


  and

  (
    g1345_p,
    g1344_p_spl_,
    g1332_n_spl_
  );


  or

  (
    g1345_n,
    g1344_n_spl_,
    g1332_p_spl_
  );


  and

  (
    g1346_p,
    g1344_n_spl_,
    g1332_p_spl_
  );


  or

  (
    g1346_n,
    g1344_p_spl_,
    g1332_n_spl_
  );


  and

  (
    g1347_p,
    g1346_n,
    g1345_n
  );


  or

  (
    g1347_n,
    g1346_p,
    g1345_p
  );


  and

  (
    g1348_p,
    G107_p_spl_10,
    G101_p_spl_101
  );


  or

  (
    g1348_n,
    G107_n_spl_10,
    G101_n_spl_101
  );


  and

  (
    g1349_p,
    G107_n_spl_10,
    G100_p_spl_101
  );


  or

  (
    g1349_n,
    G107_p_spl_10,
    G100_n_spl_101
  );


  and

  (
    g1350_p,
    g1349_n,
    g1348_n
  );


  or

  (
    g1350_n,
    g1349_p,
    g1348_p
  );


  and

  (
    g1351_p,
    g1350_n,
    G139_p_spl_1
  );


  or

  (
    g1351_n,
    g1350_p,
    G139_n_spl_1
  );


  and

  (
    g1352_p,
    G107_p_spl_11,
    G102_n_spl_101
  );


  or

  (
    g1352_n,
    G107_n_spl_11,
    G102_p_spl_101
  );


  and

  (
    g1353_p,
    G107_n_spl_11,
    G98_n_spl_101
  );


  or

  (
    g1353_n,
    G107_p_spl_11,
    G98_p_spl_101
  );


  and

  (
    g1354_p,
    g1353_n,
    g1352_n
  );


  or

  (
    g1354_n,
    g1353_p,
    g1352_p
  );


  and

  (
    g1355_p,
    g1354_n,
    G139_n_spl_1
  );


  or

  (
    g1355_n,
    g1354_p,
    G139_p_spl_1
  );


  and

  (
    g1356_p,
    g1355_n,
    g1351_n
  );


  or

  (
    g1356_n,
    g1355_p,
    g1351_p
  );


  and

  (
    g1357_p,
    G105_p_spl_10,
    G101_p_spl_110
  );


  or

  (
    g1357_n,
    G105_n_spl_10,
    G101_n_spl_110
  );


  and

  (
    g1358_p,
    G105_n_spl_10,
    G100_p_spl_110
  );


  or

  (
    g1358_n,
    G105_p_spl_10,
    G100_n_spl_110
  );


  and

  (
    g1359_p,
    g1358_n,
    g1357_n
  );


  or

  (
    g1359_n,
    g1358_p,
    g1357_p
  );


  and

  (
    g1360_p,
    g1359_n,
    G138_p_spl_1
  );


  or

  (
    g1360_n,
    g1359_p,
    G138_n_spl_1
  );


  and

  (
    g1361_p,
    G105_p_spl_11,
    G102_n_spl_101
  );


  or

  (
    g1361_n,
    G105_n_spl_11,
    G102_p_spl_101
  );


  and

  (
    g1362_p,
    G105_n_spl_11,
    G98_n_spl_110
  );


  or

  (
    g1362_n,
    G105_p_spl_11,
    G98_p_spl_110
  );


  and

  (
    g1363_p,
    g1362_n,
    g1361_n
  );


  or

  (
    g1363_n,
    g1362_p,
    g1361_p
  );


  and

  (
    g1364_p,
    g1363_n,
    G138_n_spl_1
  );


  or

  (
    g1364_n,
    g1363_p,
    G138_p_spl_1
  );


  and

  (
    g1365_p,
    g1364_n,
    g1360_n
  );


  or

  (
    g1365_n,
    g1364_p,
    g1360_p
  );


  and

  (
    g1366_p,
    g1365_p_spl_,
    g1356_n_spl_
  );


  or

  (
    g1366_n,
    g1365_n_spl_,
    g1356_p_spl_
  );


  and

  (
    g1367_p,
    g1365_n_spl_,
    g1356_p_spl_
  );


  or

  (
    g1367_n,
    g1365_p_spl_,
    g1356_n_spl_
  );


  and

  (
    g1368_p,
    g1367_n,
    g1366_n
  );


  or

  (
    g1368_n,
    g1367_p,
    g1366_p
  );


  and

  (
    g1369_p,
    G103_p_spl_10,
    G101_p_spl_110
  );


  or

  (
    g1369_n,
    G103_n_spl_10,
    G101_n_spl_110
  );


  and

  (
    g1370_p,
    G103_n_spl_10,
    G100_p_spl_110
  );


  or

  (
    g1370_n,
    G103_p_spl_10,
    G100_n_spl_110
  );


  and

  (
    g1371_p,
    g1370_n,
    g1369_n
  );


  or

  (
    g1371_n,
    g1370_p,
    g1369_p
  );


  and

  (
    g1372_p,
    g1371_n,
    G137_p_spl_1
  );


  or

  (
    g1372_n,
    g1371_p,
    G137_n_spl_1
  );


  and

  (
    g1373_p,
    G103_p_spl_11,
    G102_n_spl_110
  );


  or

  (
    g1373_n,
    G103_n_spl_11,
    G102_p_spl_110
  );


  and

  (
    g1374_p,
    G103_n_spl_11,
    G98_n_spl_110
  );


  or

  (
    g1374_n,
    G103_p_spl_11,
    G98_p_spl_110
  );


  and

  (
    g1375_p,
    g1374_n,
    g1373_n
  );


  or

  (
    g1375_n,
    g1374_p,
    g1373_p
  );


  and

  (
    g1376_p,
    g1375_n,
    G137_n_spl_1
  );


  or

  (
    g1376_n,
    g1375_p,
    G137_p_spl_1
  );


  and

  (
    g1377_p,
    g1376_n,
    g1372_n
  );


  or

  (
    g1377_n,
    g1376_p,
    g1372_p
  );


  and

  (
    g1378_p,
    G101_p_spl_111,
    G96_p_spl_10
  );


  or

  (
    g1378_n,
    G101_n_spl_111,
    G96_n_spl_10
  );


  and

  (
    g1379_p,
    G100_p_spl_111,
    G96_n_spl_10
  );


  or

  (
    g1379_n,
    G100_n_spl_111,
    G96_p_spl_10
  );


  and

  (
    g1380_p,
    g1379_n,
    g1378_n
  );


  or

  (
    g1380_n,
    g1379_p,
    g1378_p
  );


  and

  (
    g1381_p,
    g1380_n,
    G141_p_spl_1
  );


  or

  (
    g1381_n,
    g1380_p,
    G141_n_spl_1
  );


  and

  (
    g1382_p,
    G102_n_spl_110,
    G96_p_spl_11
  );


  or

  (
    g1382_n,
    G102_p_spl_110,
    G96_n_spl_11
  );


  and

  (
    g1383_p,
    G98_n_spl_111,
    G96_n_spl_11
  );


  or

  (
    g1383_n,
    G98_p_spl_111,
    G96_p_spl_11
  );


  and

  (
    g1384_p,
    g1383_n,
    g1382_n
  );


  or

  (
    g1384_n,
    g1383_p,
    g1382_p
  );


  and

  (
    g1385_p,
    g1384_n,
    G141_n_spl_1
  );


  or

  (
    g1385_n,
    g1384_p,
    G141_p_spl_1
  );


  and

  (
    g1386_p,
    g1385_n,
    g1381_n
  );


  or

  (
    g1386_n,
    g1385_p,
    g1381_p
  );


  and

  (
    g1387_p,
    g1386_p_spl_,
    g1377_n_spl_
  );


  or

  (
    g1387_n,
    g1386_n_spl_,
    g1377_p_spl_
  );


  and

  (
    g1388_p,
    g1386_n_spl_,
    g1377_p_spl_
  );


  or

  (
    g1388_n,
    g1386_p_spl_,
    g1377_n_spl_
  );


  and

  (
    g1389_p,
    g1388_n,
    g1387_n
  );


  or

  (
    g1389_n,
    g1388_p,
    g1387_p
  );


  and

  (
    g1390_p,
    G109_p_spl_10,
    G101_p_spl_111
  );


  or

  (
    g1390_n,
    G109_n_spl_10,
    G101_n_spl_111
  );


  and

  (
    g1391_p,
    G109_n_spl_10,
    G100_p_spl_111
  );


  or

  (
    g1391_n,
    G109_p_spl_10,
    G100_n_spl_111
  );


  and

  (
    g1392_p,
    g1391_n,
    g1390_n
  );


  or

  (
    g1392_n,
    g1391_p,
    g1390_p
  );


  and

  (
    g1393_p,
    g1392_n,
    G135_p_spl_1
  );


  or

  (
    g1393_n,
    g1392_p,
    G135_n_spl_1
  );


  and

  (
    g1394_p,
    G109_p_spl_11,
    G102_n_spl_11
  );


  or

  (
    g1394_n,
    G109_n_spl_11,
    G102_p_spl_11
  );


  and

  (
    g1395_p,
    G109_n_spl_11,
    G98_n_spl_111
  );


  or

  (
    g1395_n,
    G109_p_spl_11,
    G98_p_spl_111
  );


  and

  (
    g1396_p,
    g1395_n,
    g1394_n
  );


  or

  (
    g1396_n,
    g1395_p,
    g1394_p
  );


  and

  (
    g1397_p,
    g1396_n,
    G135_n_spl_1
  );


  or

  (
    g1397_n,
    g1396_p,
    G135_p_spl_1
  );


  and

  (
    g1398_p,
    g1397_n,
    g1393_n
  );


  or

  (
    g1398_n,
    g1397_p,
    g1393_p
  );


  and

  (
    g1399_p,
    g1398_n_spl_,
    g1389_p_spl_
  );


  or

  (
    g1399_n,
    g1398_p_spl_,
    g1389_n_spl_
  );


  and

  (
    g1400_p,
    g1398_p_spl_,
    g1389_n_spl_
  );


  or

  (
    g1400_n,
    g1398_n_spl_,
    g1389_p_spl_
  );


  and

  (
    g1401_p,
    g1400_n,
    g1399_n
  );


  or

  (
    g1401_n,
    g1400_p,
    g1399_p
  );


  and

  (
    g1402_p,
    g1401_n_spl_,
    g1368_p_spl_
  );


  or

  (
    g1402_n,
    g1401_p_spl_,
    g1368_n_spl_
  );


  and

  (
    g1403_p,
    g1401_p_spl_,
    g1368_n_spl_
  );


  or

  (
    g1403_n,
    g1401_n_spl_,
    g1368_p_spl_
  );


  and

  (
    g1404_p,
    g1403_n,
    g1402_n
  );


  or

  (
    g1404_n,
    g1403_p,
    g1402_p
  );


  or

  (
    g1405_n,
    g1404_n,
    g1347_p
  );


  or

  (
    g1406_n,
    g1404_p,
    g1347_n
  );


  and

  (
    g1407_p,
    g1406_n,
    g1405_n
  );


  or

  (
    g1408_n,
    g1407_p,
    G176_n_spl_111
  );


  and

  (
    g1409_p,
    g546_p_spl_1,
    g389_n_spl_
  );


  or

  (
    g1409_n,
    g546_n_spl_0,
    g389_p_spl_
  );


  and

  (
    g1410_p,
    g544_n_spl_1,
    g374_p_spl_1
  );


  or

  (
    g1410_n,
    g544_p_spl_1,
    g374_n_spl_1
  );


  and

  (
    g1411_p,
    g380_p_spl_,
    g374_n_spl_1
  );


  or

  (
    g1411_n,
    g380_n_spl_,
    g374_p_spl_1
  );


  and

  (
    g1412_p,
    g1411_n,
    g1410_n
  );


  or

  (
    g1412_n,
    g1411_p,
    g1410_p
  );


  and

  (
    g1413_p,
    g1412_n_spl_,
    g1409_n_spl_
  );


  or

  (
    g1413_n,
    g1412_p_spl_,
    g1409_p_spl_
  );


  and

  (
    g1414_p,
    g1412_p_spl_,
    g1409_p_spl_
  );


  or

  (
    g1414_n,
    g1412_n_spl_,
    g1409_n_spl_
  );


  and

  (
    g1415_p,
    g1414_n,
    g1413_n
  );


  or

  (
    g1415_n,
    g1414_p,
    g1413_p
  );


  and

  (
    g1416_p,
    g1415_p_spl_,
    g375_n_spl_0
  );


  or

  (
    g1416_n,
    g1415_n_spl_,
    g375_p_spl_0
  );


  and

  (
    g1417_p,
    g546_p_spl_1,
    g544_p_spl_1
  );


  or

  (
    g1417_n,
    g546_n_spl_,
    g544_n_spl_1
  );


  and

  (
    g1418_p,
    g1417_n,
    g545_n_spl_
  );


  or

  (
    g1418_n,
    g1417_p,
    g545_p_spl_
  );


  and

  (
    g1419_p,
    g1418_n,
    g375_p_spl_1
  );


  or

  (
    g1419_n,
    g1418_p,
    g375_n_spl_1
  );


  and

  (
    g1420_p,
    g1419_n,
    g1416_n_spl_
  );


  or

  (
    g1420_n,
    g1419_p,
    g1416_p_spl_
  );


  and

  (
    g1421_p,
    g1420_p_spl_,
    g381_n_spl_01
  );


  or

  (
    g1421_n,
    g1420_n_spl_,
    g381_p_spl_01
  );


  and

  (
    g1422_p,
    g1420_n_spl_,
    g381_p_spl_10
  );


  or

  (
    g1422_n,
    g1420_p_spl_,
    g381_n_spl_10
  );


  and

  (
    g1423_p,
    g1422_n,
    g1421_n
  );


  or

  (
    g1423_n,
    g1422_p,
    g1421_p
  );


  and

  (
    g1424_p,
    g1423_p_spl_,
    g395_n_spl_01
  );


  or

  (
    g1424_n,
    g1423_n_spl_,
    g395_p_spl_00
  );


  and

  (
    g1425_p,
    g1423_n_spl_,
    g395_p_spl_0
  );


  or

  (
    g1425_n,
    g1423_p_spl_,
    g395_n_spl_10
  );


  and

  (
    g1426_p,
    g1425_n,
    g1424_n
  );


  or

  (
    g1426_n,
    g1425_p,
    g1424_p
  );


  and

  (
    g1427_p,
    g1426_p_spl_,
    g388_n_spl_01
  );


  or

  (
    g1427_n,
    g1426_n_spl_,
    g388_p_spl_01
  );


  and

  (
    g1428_p,
    g1426_n_spl_,
    g388_p_spl_01
  );


  or

  (
    g1428_n,
    g1426_p_spl_,
    g388_n_spl_01
  );


  and

  (
    g1429_p,
    g1428_n,
    g1427_n
  );


  or

  (
    g1429_n,
    g1428_p,
    g1427_p
  );


  and

  (
    g1430_p,
    g1429_n,
    g541_p_spl_0
  );


  or

  (
    g1430_n,
    g1429_p,
    g541_n_spl_0
  );


  and

  (
    g1431_p,
    g1415_n_spl_,
    g375_p_spl_1
  );


  or

  (
    g1431_n,
    g1415_p_spl_,
    g375_n_spl_1
  );


  and

  (
    g1432_p,
    g1431_n,
    g1416_n_spl_
  );


  or

  (
    g1432_n,
    g1431_p,
    g1416_p_spl_
  );


  and

  (
    g1433_p,
    g1432_p_spl_,
    g381_n_spl_10
  );


  or

  (
    g1433_n,
    g1432_n_spl_,
    g381_p_spl_10
  );


  and

  (
    g1434_p,
    g1432_n_spl_,
    g381_p_spl_1
  );


  or

  (
    g1434_n,
    g1432_p_spl_,
    g381_n_spl_1
  );


  and

  (
    g1435_p,
    g1434_n,
    g1433_n
  );


  or

  (
    g1435_n,
    g1434_p,
    g1433_p
  );


  and

  (
    g1436_p,
    g1435_p_spl_,
    g395_n_spl_10
  );


  or

  (
    g1436_n,
    g1435_n_spl_,
    g395_p_spl_1
  );


  and

  (
    g1437_p,
    g1435_n_spl_,
    g395_p_spl_1
  );


  or

  (
    g1437_n,
    g1435_p_spl_,
    g395_n_spl_1
  );


  and

  (
    g1438_p,
    g1437_n,
    g1436_n
  );


  or

  (
    g1438_n,
    g1437_p,
    g1436_p
  );


  and

  (
    g1439_p,
    g1438_p_spl_,
    g388_n_spl_1
  );


  or

  (
    g1439_n,
    g1438_n_spl_,
    g388_p_spl_1
  );


  and

  (
    g1440_p,
    g1438_n_spl_,
    g388_p_spl_1
  );


  or

  (
    g1440_n,
    g1438_p_spl_,
    g388_n_spl_1
  );


  and

  (
    g1441_p,
    g1440_n,
    g1439_n
  );


  or

  (
    g1441_n,
    g1440_p,
    g1439_p
  );


  and

  (
    g1442_p,
    g1441_n_spl_,
    g541_n_spl_1
  );


  or

  (
    g1442_n,
    g1441_p_spl_,
    g541_p_spl_1
  );


  and

  (
    g1443_p,
    g1442_n,
    g1430_n_spl_
  );


  or

  (
    g1443_n,
    g1442_p,
    g1430_p_spl_
  );


  and

  (
    g1444_p,
    g1443_n,
    G157_n_spl_0
  );


  or

  (
    g1444_n,
    g1443_p,
    G157_p_spl_0
  );


  and

  (
    g1445_p,
    g541_p_spl_1,
    g430_n_spl_1
  );


  or

  (
    g1445_n,
    g541_n_spl_1,
    g430_p_spl_0
  );


  and

  (
    g1446_p,
    g1445_n,
    g1441_n_spl_
  );


  or

  (
    g1446_n,
    g1445_p,
    g1441_p_spl_
  );


  and

  (
    g1447_p,
    g1430_p_spl_,
    g430_n_spl_1
  );


  or

  (
    g1447_n,
    g1430_n_spl_,
    g430_p_spl_
  );


  and

  (
    g1448_p,
    g1447_n,
    g1446_n
  );


  or

  (
    g1448_n,
    g1447_p,
    g1446_p
  );


  and

  (
    g1449_p,
    g1448_n,
    G157_p_spl_0
  );


  or

  (
    g1449_n,
    g1448_p,
    G157_n_spl_0
  );


  and

  (
    g1450_p,
    g1449_n,
    g1444_n
  );


  or

  (
    g1450_n,
    g1449_p,
    g1444_p
  );


  and

  (
    g1451_p,
    g537_n_spl_0,
    g400_p_spl_1
  );


  or

  (
    g1451_n,
    g537_p_spl_0,
    g400_n_spl_1
  );


  and

  (
    g1452_p,
    g537_p_spl_1,
    g400_n_spl_1
  );


  or

  (
    g1452_n,
    g537_n_spl_1,
    g400_p_spl_1
  );


  and

  (
    g1453_p,
    g1452_n,
    g1451_n
  );


  or

  (
    g1453_n,
    g1452_p,
    g1451_p
  );


  and

  (
    g1454_p,
    g1453_n_spl_,
    g535_p_spl_0
  );


  or

  (
    g1454_n,
    g1453_p_spl_,
    g535_n_spl_0
  );


  and

  (
    g1455_p,
    g1453_p_spl_,
    g535_n_spl_1
  );


  or

  (
    g1455_n,
    g1453_n_spl_,
    g535_p_spl_1
  );


  and

  (
    g1456_p,
    g1455_n,
    g1454_n
  );


  or

  (
    g1456_n,
    g1455_p,
    g1454_p
  );


  and

  (
    g1457_p,
    g408_n_spl_1,
    g402_n_spl_
  );


  or

  (
    g1457_n,
    g408_p_spl_1,
    g402_p_spl_1
  );


  and

  (
    g1458_p,
    g1457_n,
    g409_n_spl_0
  );


  or

  (
    g1458_n,
    g1457_p,
    g409_p_spl_0
  );


  and

  (
    g1459_p,
    g1458_n_spl_0,
    g539_n_spl_0
  );


  or

  (
    g1459_n,
    g1458_p_spl_0,
    g539_p_spl_0
  );


  and

  (
    g1460_p,
    g1458_p_spl_0,
    g539_p_spl_1
  );


  or

  (
    g1460_n,
    g1458_n_spl_0,
    g539_n_spl_1
  );


  and

  (
    g1461_p,
    g1460_n,
    g1459_n
  );


  or

  (
    g1461_n,
    g1460_p,
    g1459_p
  );


  and

  (
    g1462_p,
    g1461_p_spl_,
    g1456_n_spl_
  );


  or

  (
    g1462_n,
    g1461_n_spl_,
    g1456_p_spl_
  );


  and

  (
    g1463_p,
    g1461_n_spl_,
    g1456_p_spl_
  );


  or

  (
    g1463_n,
    g1461_p_spl_,
    g1456_n_spl_
  );


  and

  (
    g1464_p,
    g1463_n,
    g1462_n
  );


  or

  (
    g1464_n,
    g1463_p,
    g1462_p
  );


  and

  (
    g1465_p,
    g1464_n_spl_,
    g429_n_spl_01
  );


  or

  (
    g1465_n,
    g1464_p_spl_,
    g429_p_spl_01
  );


  and

  (
    g1466_p,
    g1464_p_spl_,
    g429_p_spl_10
  );


  or

  (
    g1466_n,
    g1464_n_spl_,
    g429_n_spl_10
  );


  and

  (
    g1467_p,
    g1466_n,
    g1465_n
  );


  or

  (
    g1467_n,
    g1466_p,
    g1465_p
  );


  and

  (
    g1468_p,
    g1467_p,
    G157_n_spl_1
  );


  or

  (
    g1468_n,
    g1467_n,
    G157_p_spl_1
  );


  and

  (
    g1469_p,
    g539_p_spl_1,
    g423_n_spl_
  );


  or

  (
    g1469_n,
    g539_n_spl_1,
    g423_p_spl_
  );


  and

  (
    g1470_p,
    g535_p_spl_1,
    g409_n_spl_
  );


  or

  (
    g1470_n,
    g535_n_spl_1,
    g409_p_spl_
  );


  and

  (
    g1471_p,
    g537_p_spl_1,
    g416_n_spl_
  );


  or

  (
    g1471_n,
    g537_n_spl_1,
    g416_p_spl_
  );


  and

  (
    g1472_p,
    g1471_n_spl_,
    g401_n_spl_0
  );


  or

  (
    g1472_n,
    g1471_p_spl_,
    g401_p_spl_0
  );


  and

  (
    g1473_p,
    g1471_p_spl_,
    g401_p_spl_
  );


  or

  (
    g1473_n,
    g1471_n_spl_,
    g401_n_spl_
  );


  and

  (
    g1474_p,
    g1473_n,
    g1472_n
  );


  or

  (
    g1474_n,
    g1473_p,
    g1472_p
  );


  and

  (
    g1475_p,
    g1474_p_spl_,
    g1470_n_spl_
  );


  or

  (
    g1475_n,
    g1474_n_spl_,
    g1470_p_spl_
  );


  and

  (
    g1476_p,
    g1474_n_spl_,
    g1470_p_spl_
  );


  or

  (
    g1476_n,
    g1474_p_spl_,
    g1470_n_spl_
  );


  and

  (
    g1477_p,
    g1476_n,
    g1475_n
  );


  or

  (
    g1477_n,
    g1476_p,
    g1475_p
  );


  and

  (
    g1478_p,
    g1477_p_spl_,
    g1469_n_spl_
  );


  or

  (
    g1478_n,
    g1477_n_spl_,
    g1469_p_spl_
  );


  and

  (
    g1479_p,
    g1477_n_spl_,
    g1469_p_spl_
  );


  or

  (
    g1479_n,
    g1477_p_spl_,
    g1469_n_spl_
  );


  and

  (
    g1480_p,
    g1479_n,
    g1478_n
  );


  or

  (
    g1480_n,
    g1479_p,
    g1478_p
  );


  and

  (
    g1481_p,
    g1458_n_spl_1,
    g429_n_spl_10
  );


  or

  (
    g1481_n,
    g1458_p_spl_1,
    g429_p_spl_10
  );


  and

  (
    g1482_p,
    g1458_p_spl_1,
    g429_p_spl_1
  );


  or

  (
    g1482_n,
    g1458_n_spl_1,
    g429_n_spl_1
  );


  and

  (
    g1483_p,
    g1482_n,
    g1481_n
  );


  or

  (
    g1483_n,
    g1482_p,
    g1481_p
  );


  and

  (
    g1484_p,
    g1483_p_spl_,
    g1480_n_spl_
  );


  or

  (
    g1484_n,
    g1483_n_spl_,
    g1480_p_spl_
  );


  and

  (
    g1485_p,
    g1483_n_spl_,
    g1480_p_spl_
  );


  or

  (
    g1485_n,
    g1483_p_spl_,
    g1480_n_spl_
  );


  and

  (
    g1486_p,
    g1485_n,
    g1484_n
  );


  or

  (
    g1486_n,
    g1485_p,
    g1484_p
  );


  and

  (
    g1487_p,
    g1486_n,
    G157_p_spl_1
  );


  or

  (
    g1487_n,
    g1486_p,
    G157_n_spl_1
  );


  and

  (
    g1488_p,
    g1487_n,
    g1468_n
  );


  or

  (
    g1488_n,
    g1487_p,
    g1468_p
  );


  and

  (
    g1489_p,
    g1488_p_spl_,
    g415_p_spl_1
  );


  or

  (
    g1489_n,
    g1488_n_spl_,
    g415_n_spl_1
  );


  and

  (
    g1490_p,
    g1488_n_spl_,
    g415_n_spl_1
  );


  or

  (
    g1490_n,
    g1488_p_spl_,
    g415_p_spl_1
  );


  and

  (
    g1491_p,
    g1490_n,
    g1489_n
  );


  or

  (
    g1491_n,
    g1490_p,
    g1489_p
  );


  and

  (
    g1492_p,
    g1491_n_spl_,
    g422_p_spl_1
  );


  or

  (
    g1492_n,
    g1491_p_spl_,
    g422_n_spl_1
  );


  and

  (
    g1493_p,
    g1491_p_spl_,
    g422_n_spl_1
  );


  or

  (
    g1493_n,
    g1491_n_spl_,
    g422_p_spl_1
  );


  and

  (
    g1494_p,
    g1493_n,
    g1492_n
  );


  or

  (
    g1494_n,
    g1493_p,
    g1492_p
  );


  and

  (
    g1495_p,
    g1494_n,
    g1450_n
  );


  and

  (
    g1496_p,
    g1494_p,
    g1450_p
  );


  or

  (
    g1497_n,
    g1496_p,
    G176_p_spl_1111
  );


  or

  (
    g1498_n,
    g1497_n,
    g1495_p
  );


  and

  (
    g1499_p,
    g1498_n,
    g1408_n
  );


  or

  (
    g1500_n,
    g1499_p,
    G177_n_spl_111
  );


  or

  (
    g1501_n,
    G177_p_spl_110,
    G49_p
  );


  or

  (
    g1502_n,
    g1501_n,
    G176_n_spl_111
  );


  and

  (
    g1503_p,
    g1502_n,
    g1500_n_spl_
  );


  or

  (
    g1504_n,
    G173_p_spl_111,
    G23_n_spl_
  );


  or

  (
    g1505_n,
    G173_n_spl_111,
    G4_n_spl_
  );


  and

  (
    g1506_p,
    g1505_n,
    g1504_n
  );


  or

  (
    g1507_n,
    g1506_p,
    G172_p_spl_11
  );


  or

  (
    g1508_n,
    G177_p_spl_111,
    G38_n
  );


  and

  (
    g1509_p,
    g1508_n,
    g1500_n_spl_
  );


  and

  (
    g1510_p,
    g1509_p_spl_0,
    G173_n_spl_111
  );


  or

  (
    g1511_n,
    G177_p_spl_111,
    G37_n
  );


  and

  (
    g1512_p,
    g1511_n,
    g1308_n_spl_
  );


  and

  (
    g1513_p,
    g1512_p_spl_0,
    G173_p_spl_111
  );


  or

  (
    g1514_n,
    g1513_p,
    G172_n_spl_11
  );


  or

  (
    g1515_n,
    g1514_n,
    g1510_p
  );


  and

  (
    g1516_p,
    g1515_n,
    g1507_n
  );


  or

  (
    g1517_n,
    G174_p_spl_111,
    G23_n_spl_
  );


  or

  (
    g1518_n,
    G174_n_spl_111,
    G4_n_spl_
  );


  and

  (
    g1519_p,
    g1518_n,
    g1517_n
  );


  or

  (
    g1520_n,
    g1519_p,
    G175_p_spl_11
  );


  and

  (
    g1521_p,
    g1509_p_spl_0,
    G174_n_spl_111
  );


  and

  (
    g1522_p,
    g1512_p_spl_0,
    G174_p_spl_111
  );


  or

  (
    g1523_n,
    g1522_p,
    G175_n_spl_11
  );


  or

  (
    g1524_n,
    g1523_n,
    g1521_p
  );


  and

  (
    g1525_p,
    g1524_n,
    g1520_n
  );


  or

  (
    g1526_n,
    G158_p_spl_111,
    G79_n_spl_
  );


  or

  (
    g1527_n,
    G158_n_spl_111,
    G78_n_spl_
  );


  and

  (
    g1528_p,
    g1527_n,
    g1526_n
  );


  or

  (
    g1529_n,
    g1528_p,
    G159_p_spl_11
  );


  or

  (
    g1530_n,
    g1512_p_spl_1,
    G158_n_spl_111
  );


  or

  (
    g1531_n,
    g1509_p_spl_1,
    G158_p_spl_111
  );


  and

  (
    g1532_p,
    g1531_n,
    g1530_n
  );


  or

  (
    g1533_n,
    g1532_p,
    G159_n_spl_11
  );


  and

  (
    g1534_p,
    g1533_n,
    g1529_n
  );


  or

  (
    g1535_n,
    g1534_p,
    G64_n_spl_
  );


  or

  (
    g1536_n,
    G160_p_spl_111,
    G79_n_spl_
  );


  or

  (
    g1537_n,
    G160_n_spl_111,
    G78_n_spl_
  );


  and

  (
    g1538_p,
    g1537_n,
    g1536_n
  );


  or

  (
    g1539_n,
    g1538_p,
    G161_p_spl_11
  );


  or

  (
    g1540_n,
    g1512_p_spl_1,
    G160_n_spl_111
  );


  or

  (
    g1541_n,
    g1509_p_spl_1,
    G160_p_spl_111
  );


  and

  (
    g1542_p,
    g1541_n,
    g1540_n
  );


  or

  (
    g1543_n,
    g1542_p,
    G161_n_spl_11
  );


  and

  (
    g1544_p,
    g1543_n,
    g1539_n
  );


  or

  (
    g1545_n,
    g1544_p,
    G64_n_spl_
  );


  buf

  (
    G5193,
    G66_n
  );


  buf

  (
    G5194,
    G113_n_spl_1
  );


  buf

  (
    G5195,
    G165_n_spl_
  );


  buf

  (
    G5196,
    G151_n_spl_0
  );


  buf

  (
    G5197,
    G127_n_spl_
  );


  buf

  (
    G5198,
    G131_n_spl_
  );


  not

  (
    G5199,
    g179_n_spl_
  );


  buf

  (
    G5200,
    G152_n
  );


  buf

  (
    G5201,
    G151_n_spl_0
  );


  buf

  (
    G5202,
    G151_n_spl_
  );


  buf

  (
    G5203,
    G125_n_spl_
  );


  buf

  (
    G5204,
    G129_n_spl_
  );


  buf

  (
    G5205,
    g180_p
  );


  buf

  (
    G5206,
    G99_n_spl_
  );


  buf

  (
    G5207,
    G153_n_spl_
  );


  buf

  (
    G5208,
    G156_n_spl_
  );


  buf

  (
    G5209,
    G155_n_spl_
  );


  buf

  (
    G5210,
    g181_p
  );


  buf

  (
    G5211,
    g182_p
  );


  buf

  (
    G5212,
    g183_n
  );


  buf

  (
    G5213,
    g184_n_spl_
  );


  buf

  (
    G5214,
    G64_p_spl_111
  );


  buf

  (
    G5215,
    G66_p_spl_1
  );


  buf

  (
    G5216,
    G1_p_spl_
  );


  buf

  (
    G5217,
    G152_p_spl_
  );


  buf

  (
    G5218,
    G114_p_spl_
  );


  buf

  (
    G5219,
    G152_p_spl_
  );


  buf

  (
    G5220,
    g186_n
  );


  buf

  (
    G5221,
    g185_n_spl_11
  );


  buf

  (
    G5222,
    G1_n_spl_0
  );


  buf

  (
    G5223,
    G1_n_spl_0
  );


  buf

  (
    G5224,
    G1_n_spl_1
  );


  buf

  (
    G5225,
    G1_n_spl_1
  );


  buf

  (
    G5226,
    G114_n_spl_0
  );


  buf

  (
    G5227,
    G114_n_spl_
  );


  buf

  (
    G5228,
    g190_n
  );


  buf

  (
    G5229,
    g194_n_spl_
  );


  buf

  (
    G5230,
    g194_n_spl_
  );


  buf

  (
    G5231,
    g195_n
  );


  buf

  (
    G5232,
    g200_p
  );


  buf

  (
    G5233,
    g205_p
  );


  buf

  (
    G5234,
    g210_p
  );


  buf

  (
    G5235,
    g215_p
  );


  not

  (
    G5236,
    g280_n
  );


  not

  (
    G5237,
    g369_n
  );


  not

  (
    G5238,
    g431_n_spl_
  );


  buf

  (
    G5239,
    g482_p_spl_
  );


  buf

  (
    G5240,
    g482_p_spl_
  );


  not

  (
    G5241,
    g431_n_spl_
  );


  not

  (
    G5242,
    g506_n_spl_
  );


  not

  (
    G5243,
    g533_n_spl_
  );


  not

  (
    G5244,
    g549_p_spl_
  );


  buf

  (
    G5245,
    g550_n_spl_
  );


  not

  (
    G5246,
    g549_p_spl_
  );


  buf

  (
    G5247,
    g550_n_spl_
  );


  not

  (
    G5248,
    g560_p_spl_1
  );


  not

  (
    G5249,
    g569_p_spl_1
  );


  not

  (
    G5250,
    g579_p_spl_1
  );


  buf

  (
    G5251,
    g581_p_spl_1
  );


  buf

  (
    G5252,
    g590_n
  );


  not

  (
    G5253,
    g605_n_spl_1
  );


  not

  (
    G5254,
    g614_n_spl_1
  );


  not

  (
    G5255,
    g624_n_spl_1
  );


  buf

  (
    G5256,
    g633_n
  );


  not

  (
    G5257,
    g647_n_spl_1
  );


  not

  (
    G5258,
    g656_n_spl_1
  );


  not

  (
    G5259,
    g669_n_spl_1
  );


  not

  (
    G5260,
    g678_n_spl_1
  );


  not

  (
    G5261,
    g705_n_spl_
  );


  not

  (
    G5262,
    g735_n_spl_
  );


  not

  (
    G5263,
    g764_n
  );


  not

  (
    G5264,
    g794_n
  );


  buf

  (
    G5265,
    g804_p
  );


  buf

  (
    G5266,
    g814_p
  );


  buf

  (
    G5267,
    g823_n
  );


  buf

  (
    G5268,
    g832_n
  );


  buf

  (
    G5269,
    g841_n
  );


  buf

  (
    G5270,
    g850_n
  );


  buf

  (
    G5271,
    g859_n
  );


  buf

  (
    G5272,
    g868_n
  );


  buf

  (
    G5273,
    g877_n
  );


  buf

  (
    G5274,
    g886_n
  );


  buf

  (
    G5275,
    g896_p
  );


  buf

  (
    G5276,
    g906_p
  );


  buf

  (
    G5277,
    g916_p
  );


  buf

  (
    G5278,
    g926_p
  );


  buf

  (
    G5279,
    g936_p
  );


  buf

  (
    G5280,
    g946_p
  );


  buf

  (
    G5281,
    g956_p
  );


  buf

  (
    G5282,
    g966_p
  );


  buf

  (
    G5283,
    g980_p
  );


  buf

  (
    G5284,
    g983_n
  );


  not

  (
    G5285,
    g990_p_spl_1
  );


  not

  (
    G5286,
    g997_n_spl_1
  );


  not

  (
    G5287,
    g1004_n_spl_1
  );


  not

  (
    G5288,
    g1011_n_spl_1
  );


  not

  (
    G5289,
    g1018_n
  );


  not

  (
    G5290,
    g1025_n_spl_1
  );


  not

  (
    G5291,
    g1032_n_spl_1
  );


  not

  (
    G5292,
    g1039_n_spl_1
  );


  not

  (
    G5293,
    g1046_n_spl_1
  );


  buf

  (
    G5294,
    g1055_n
  );


  buf

  (
    G5295,
    g1064_n
  );


  buf

  (
    G5296,
    g1073_n
  );


  buf

  (
    G5297,
    g1082_n
  );


  buf

  (
    G5298,
    g1091_n
  );


  buf

  (
    G5299,
    g1100_n
  );


  buf

  (
    G5300,
    g1109_n
  );


  buf

  (
    G5301,
    g1118_n
  );


  buf

  (
    G5302,
    g1128_p
  );


  buf

  (
    G5303,
    g1138_p
  );


  buf

  (
    G5304,
    g1148_p
  );


  buf

  (
    G5305,
    g1158_p
  );


  buf

  (
    G5306,
    g1168_p
  );


  buf

  (
    G5307,
    g1178_p
  );


  buf

  (
    G5308,
    g1188_p
  );


  buf

  (
    G5309,
    g1198_p
  );


  buf

  (
    G5310,
    g1311_p
  );


  buf

  (
    G5311,
    g1503_p
  );


  not

  (
    G5312,
    g1516_p
  );


  not

  (
    G5313,
    g1525_p
  );


  buf

  (
    G5314,
    g1535_n
  );


  buf

  (
    G5315,
    g1545_n
  );


  buf

  (
    G156_n_spl_,
    G156_n
  );


  buf

  (
    G153_n_spl_,
    G153_n
  );


  buf

  (
    G66_p_spl_,
    G66_p
  );


  buf

  (
    G66_p_spl_0,
    G66_p_spl_
  );


  buf

  (
    G66_p_spl_00,
    G66_p_spl_0
  );


  buf

  (
    G66_p_spl_01,
    G66_p_spl_0
  );


  buf

  (
    G66_p_spl_1,
    G66_p_spl_
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G165_n_spl_,
    G165_n
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    g185_n_spl_,
    g185_n
  );


  buf

  (
    g185_n_spl_0,
    g185_n_spl_
  );


  buf

  (
    g185_n_spl_00,
    g185_n_spl_0
  );


  buf

  (
    g185_n_spl_000,
    g185_n_spl_00
  );


  buf

  (
    g185_n_spl_01,
    g185_n_spl_0
  );


  buf

  (
    g185_n_spl_1,
    g185_n_spl_
  );


  buf

  (
    g185_n_spl_10,
    g185_n_spl_1
  );


  buf

  (
    g185_n_spl_11,
    g185_n_spl_1
  );


  buf

  (
    G163_n_spl_,
    G163_n
  );


  buf

  (
    G163_n_spl_0,
    G163_n_spl_
  );


  buf

  (
    G163_n_spl_00,
    G163_n_spl_0
  );


  buf

  (
    G163_n_spl_01,
    G163_n_spl_0
  );


  buf

  (
    G163_n_spl_1,
    G163_n_spl_
  );


  buf

  (
    G163_p_spl_,
    G163_p
  );


  buf

  (
    G163_p_spl_0,
    G163_p_spl_
  );


  buf

  (
    G163_p_spl_00,
    G163_p_spl_0
  );


  buf

  (
    G163_p_spl_01,
    G163_p_spl_0
  );


  buf

  (
    G163_p_spl_1,
    G163_p_spl_
  );


  buf

  (
    G168_p_spl_,
    G168_p
  );


  buf

  (
    G168_p_spl_0,
    G168_p_spl_
  );


  buf

  (
    G168_p_spl_00,
    G168_p_spl_0
  );


  buf

  (
    G168_p_spl_000,
    G168_p_spl_00
  );


  buf

  (
    G168_p_spl_001,
    G168_p_spl_00
  );


  buf

  (
    G168_p_spl_01,
    G168_p_spl_0
  );


  buf

  (
    G168_p_spl_010,
    G168_p_spl_01
  );


  buf

  (
    G168_p_spl_1,
    G168_p_spl_
  );


  buf

  (
    G168_p_spl_10,
    G168_p_spl_1
  );


  buf

  (
    G168_p_spl_11,
    G168_p_spl_1
  );


  buf

  (
    G128_p_spl_,
    G128_p
  );


  buf

  (
    G128_p_spl_0,
    G128_p_spl_
  );


  buf

  (
    G128_p_spl_00,
    G128_p_spl_0
  );


  buf

  (
    G128_p_spl_000,
    G128_p_spl_00
  );


  buf

  (
    G128_p_spl_01,
    G128_p_spl_0
  );


  buf

  (
    G128_p_spl_1,
    G128_p_spl_
  );


  buf

  (
    G128_p_spl_10,
    G128_p_spl_1
  );


  buf

  (
    G128_p_spl_11,
    G128_p_spl_1
  );


  buf

  (
    G169_p_spl_,
    G169_p
  );


  buf

  (
    G169_p_spl_0,
    G169_p_spl_
  );


  buf

  (
    G169_p_spl_00,
    G169_p_spl_0
  );


  buf

  (
    G169_p_spl_000,
    G169_p_spl_00
  );


  buf

  (
    G169_p_spl_001,
    G169_p_spl_00
  );


  buf

  (
    G169_p_spl_01,
    G169_p_spl_0
  );


  buf

  (
    G169_p_spl_010,
    G169_p_spl_01
  );


  buf

  (
    G169_p_spl_011,
    G169_p_spl_01
  );


  buf

  (
    G169_p_spl_1,
    G169_p_spl_
  );


  buf

  (
    G169_p_spl_10,
    G169_p_spl_1
  );


  buf

  (
    G169_p_spl_11,
    G169_p_spl_1
  );


  buf

  (
    G128_n_spl_,
    G128_n
  );


  buf

  (
    G128_n_spl_0,
    G128_n_spl_
  );


  buf

  (
    G128_n_spl_00,
    G128_n_spl_0
  );


  buf

  (
    G128_n_spl_000,
    G128_n_spl_00
  );


  buf

  (
    G128_n_spl_01,
    G128_n_spl_0
  );


  buf

  (
    G128_n_spl_1,
    G128_n_spl_
  );


  buf

  (
    G128_n_spl_10,
    G128_n_spl_1
  );


  buf

  (
    G128_n_spl_11,
    G128_n_spl_1
  );


  buf

  (
    G150_p_spl_,
    G150_p
  );


  buf

  (
    G150_p_spl_0,
    G150_p_spl_
  );


  buf

  (
    G150_p_spl_00,
    G150_p_spl_0
  );


  buf

  (
    G150_p_spl_1,
    G150_p_spl_
  );


  buf

  (
    G167_n_spl_,
    G167_n
  );


  buf

  (
    G167_n_spl_0,
    G167_n_spl_
  );


  buf

  (
    G167_n_spl_00,
    G167_n_spl_0
  );


  buf

  (
    G167_n_spl_000,
    G167_n_spl_00
  );


  buf

  (
    G167_n_spl_001,
    G167_n_spl_00
  );


  buf

  (
    G167_n_spl_01,
    G167_n_spl_0
  );


  buf

  (
    G167_n_spl_010,
    G167_n_spl_01
  );


  buf

  (
    G167_n_spl_1,
    G167_n_spl_
  );


  buf

  (
    G167_n_spl_10,
    G167_n_spl_1
  );


  buf

  (
    G167_n_spl_11,
    G167_n_spl_1
  );


  buf

  (
    G166_n_spl_,
    G166_n
  );


  buf

  (
    G166_n_spl_0,
    G166_n_spl_
  );


  buf

  (
    G166_n_spl_00,
    G166_n_spl_0
  );


  buf

  (
    G166_n_spl_000,
    G166_n_spl_00
  );


  buf

  (
    G166_n_spl_001,
    G166_n_spl_00
  );


  buf

  (
    G166_n_spl_01,
    G166_n_spl_0
  );


  buf

  (
    G166_n_spl_010,
    G166_n_spl_01
  );


  buf

  (
    G166_n_spl_011,
    G166_n_spl_01
  );


  buf

  (
    G166_n_spl_1,
    G166_n_spl_
  );


  buf

  (
    G166_n_spl_10,
    G166_n_spl_1
  );


  buf

  (
    G166_n_spl_11,
    G166_n_spl_1
  );


  buf

  (
    G150_n_spl_,
    G150_n
  );


  buf

  (
    G150_n_spl_0,
    G150_n_spl_
  );


  buf

  (
    G150_n_spl_00,
    G150_n_spl_0
  );


  buf

  (
    G150_n_spl_1,
    G150_n_spl_
  );


  buf

  (
    G126_p_spl_,
    G126_p
  );


  buf

  (
    G126_p_spl_0,
    G126_p_spl_
  );


  buf

  (
    G126_p_spl_00,
    G126_p_spl_0
  );


  buf

  (
    G126_p_spl_000,
    G126_p_spl_00
  );


  buf

  (
    G126_p_spl_01,
    G126_p_spl_0
  );


  buf

  (
    G126_p_spl_1,
    G126_p_spl_
  );


  buf

  (
    G126_p_spl_10,
    G126_p_spl_1
  );


  buf

  (
    G126_p_spl_11,
    G126_p_spl_1
  );


  buf

  (
    G126_n_spl_,
    G126_n
  );


  buf

  (
    G126_n_spl_0,
    G126_n_spl_
  );


  buf

  (
    G126_n_spl_00,
    G126_n_spl_0
  );


  buf

  (
    G126_n_spl_000,
    G126_n_spl_00
  );


  buf

  (
    G126_n_spl_01,
    G126_n_spl_0
  );


  buf

  (
    G126_n_spl_1,
    G126_n_spl_
  );


  buf

  (
    G126_n_spl_10,
    G126_n_spl_1
  );


  buf

  (
    G126_n_spl_11,
    G126_n_spl_1
  );


  buf

  (
    G149_p_spl_,
    G149_p
  );


  buf

  (
    G149_p_spl_0,
    G149_p_spl_
  );


  buf

  (
    G149_p_spl_00,
    G149_p_spl_0
  );


  buf

  (
    G149_p_spl_1,
    G149_p_spl_
  );


  buf

  (
    G149_n_spl_,
    G149_n
  );


  buf

  (
    G149_n_spl_0,
    G149_n_spl_
  );


  buf

  (
    G149_n_spl_00,
    G149_n_spl_0
  );


  buf

  (
    G149_n_spl_1,
    G149_n_spl_
  );


  buf

  (
    g233_n_spl_,
    g233_n
  );


  buf

  (
    g224_n_spl_,
    g224_n
  );


  buf

  (
    G113_p_spl_,
    G113_p
  );


  buf

  (
    G113_p_spl_0,
    G113_p_spl_
  );


  buf

  (
    G113_p_spl_00,
    G113_p_spl_0
  );


  buf

  (
    G113_p_spl_1,
    G113_p_spl_
  );


  buf

  (
    G102_p_spl_,
    G102_p
  );


  buf

  (
    G102_p_spl_0,
    G102_p_spl_
  );


  buf

  (
    G102_p_spl_00,
    G102_p_spl_0
  );


  buf

  (
    G102_p_spl_000,
    G102_p_spl_00
  );


  buf

  (
    G102_p_spl_001,
    G102_p_spl_00
  );


  buf

  (
    G102_p_spl_01,
    G102_p_spl_0
  );


  buf

  (
    G102_p_spl_010,
    G102_p_spl_01
  );


  buf

  (
    G102_p_spl_011,
    G102_p_spl_01
  );


  buf

  (
    G102_p_spl_1,
    G102_p_spl_
  );


  buf

  (
    G102_p_spl_10,
    G102_p_spl_1
  );


  buf

  (
    G102_p_spl_100,
    G102_p_spl_10
  );


  buf

  (
    G102_p_spl_101,
    G102_p_spl_10
  );


  buf

  (
    G102_p_spl_11,
    G102_p_spl_1
  );


  buf

  (
    G102_p_spl_110,
    G102_p_spl_11
  );


  buf

  (
    G113_n_spl_,
    G113_n
  );


  buf

  (
    G113_n_spl_0,
    G113_n_spl_
  );


  buf

  (
    G113_n_spl_00,
    G113_n_spl_0
  );


  buf

  (
    G113_n_spl_01,
    G113_n_spl_0
  );


  buf

  (
    G113_n_spl_1,
    G113_n_spl_
  );


  buf

  (
    G102_n_spl_,
    G102_n
  );


  buf

  (
    G102_n_spl_0,
    G102_n_spl_
  );


  buf

  (
    G102_n_spl_00,
    G102_n_spl_0
  );


  buf

  (
    G102_n_spl_000,
    G102_n_spl_00
  );


  buf

  (
    G102_n_spl_001,
    G102_n_spl_00
  );


  buf

  (
    G102_n_spl_01,
    G102_n_spl_0
  );


  buf

  (
    G102_n_spl_010,
    G102_n_spl_01
  );


  buf

  (
    G102_n_spl_011,
    G102_n_spl_01
  );


  buf

  (
    G102_n_spl_1,
    G102_n_spl_
  );


  buf

  (
    G102_n_spl_10,
    G102_n_spl_1
  );


  buf

  (
    G102_n_spl_100,
    G102_n_spl_10
  );


  buf

  (
    G102_n_spl_101,
    G102_n_spl_10
  );


  buf

  (
    G102_n_spl_11,
    G102_n_spl_1
  );


  buf

  (
    G102_n_spl_110,
    G102_n_spl_11
  );


  buf

  (
    G98_p_spl_,
    G98_p
  );


  buf

  (
    G98_p_spl_0,
    G98_p_spl_
  );


  buf

  (
    G98_p_spl_00,
    G98_p_spl_0
  );


  buf

  (
    G98_p_spl_000,
    G98_p_spl_00
  );


  buf

  (
    G98_p_spl_001,
    G98_p_spl_00
  );


  buf

  (
    G98_p_spl_01,
    G98_p_spl_0
  );


  buf

  (
    G98_p_spl_010,
    G98_p_spl_01
  );


  buf

  (
    G98_p_spl_011,
    G98_p_spl_01
  );


  buf

  (
    G98_p_spl_1,
    G98_p_spl_
  );


  buf

  (
    G98_p_spl_10,
    G98_p_spl_1
  );


  buf

  (
    G98_p_spl_100,
    G98_p_spl_10
  );


  buf

  (
    G98_p_spl_101,
    G98_p_spl_10
  );


  buf

  (
    G98_p_spl_11,
    G98_p_spl_1
  );


  buf

  (
    G98_p_spl_110,
    G98_p_spl_11
  );


  buf

  (
    G98_p_spl_111,
    G98_p_spl_11
  );


  buf

  (
    G98_n_spl_,
    G98_n
  );


  buf

  (
    G98_n_spl_0,
    G98_n_spl_
  );


  buf

  (
    G98_n_spl_00,
    G98_n_spl_0
  );


  buf

  (
    G98_n_spl_000,
    G98_n_spl_00
  );


  buf

  (
    G98_n_spl_001,
    G98_n_spl_00
  );


  buf

  (
    G98_n_spl_01,
    G98_n_spl_0
  );


  buf

  (
    G98_n_spl_010,
    G98_n_spl_01
  );


  buf

  (
    G98_n_spl_011,
    G98_n_spl_01
  );


  buf

  (
    G98_n_spl_1,
    G98_n_spl_
  );


  buf

  (
    G98_n_spl_10,
    G98_n_spl_1
  );


  buf

  (
    G98_n_spl_100,
    G98_n_spl_10
  );


  buf

  (
    G98_n_spl_101,
    G98_n_spl_10
  );


  buf

  (
    G98_n_spl_11,
    G98_n_spl_1
  );


  buf

  (
    G98_n_spl_110,
    G98_n_spl_11
  );


  buf

  (
    G98_n_spl_111,
    G98_n_spl_11
  );


  buf

  (
    G115_p_spl_,
    G115_p
  );


  buf

  (
    G115_p_spl_0,
    G115_p_spl_
  );


  buf

  (
    G115_p_spl_00,
    G115_p_spl_0
  );


  buf

  (
    G115_p_spl_1,
    G115_p_spl_
  );


  buf

  (
    G101_p_spl_,
    G101_p
  );


  buf

  (
    G101_p_spl_0,
    G101_p_spl_
  );


  buf

  (
    G101_p_spl_00,
    G101_p_spl_0
  );


  buf

  (
    G101_p_spl_000,
    G101_p_spl_00
  );


  buf

  (
    G101_p_spl_001,
    G101_p_spl_00
  );


  buf

  (
    G101_p_spl_01,
    G101_p_spl_0
  );


  buf

  (
    G101_p_spl_010,
    G101_p_spl_01
  );


  buf

  (
    G101_p_spl_011,
    G101_p_spl_01
  );


  buf

  (
    G101_p_spl_1,
    G101_p_spl_
  );


  buf

  (
    G101_p_spl_10,
    G101_p_spl_1
  );


  buf

  (
    G101_p_spl_100,
    G101_p_spl_10
  );


  buf

  (
    G101_p_spl_101,
    G101_p_spl_10
  );


  buf

  (
    G101_p_spl_11,
    G101_p_spl_1
  );


  buf

  (
    G101_p_spl_110,
    G101_p_spl_11
  );


  buf

  (
    G101_p_spl_111,
    G101_p_spl_11
  );


  buf

  (
    G115_n_spl_,
    G115_n
  );


  buf

  (
    G115_n_spl_0,
    G115_n_spl_
  );


  buf

  (
    G115_n_spl_00,
    G115_n_spl_0
  );


  buf

  (
    G115_n_spl_1,
    G115_n_spl_
  );


  buf

  (
    G101_n_spl_,
    G101_n
  );


  buf

  (
    G101_n_spl_0,
    G101_n_spl_
  );


  buf

  (
    G101_n_spl_00,
    G101_n_spl_0
  );


  buf

  (
    G101_n_spl_000,
    G101_n_spl_00
  );


  buf

  (
    G101_n_spl_001,
    G101_n_spl_00
  );


  buf

  (
    G101_n_spl_01,
    G101_n_spl_0
  );


  buf

  (
    G101_n_spl_010,
    G101_n_spl_01
  );


  buf

  (
    G101_n_spl_011,
    G101_n_spl_01
  );


  buf

  (
    G101_n_spl_1,
    G101_n_spl_
  );


  buf

  (
    G101_n_spl_10,
    G101_n_spl_1
  );


  buf

  (
    G101_n_spl_100,
    G101_n_spl_10
  );


  buf

  (
    G101_n_spl_101,
    G101_n_spl_10
  );


  buf

  (
    G101_n_spl_11,
    G101_n_spl_1
  );


  buf

  (
    G101_n_spl_110,
    G101_n_spl_11
  );


  buf

  (
    G101_n_spl_111,
    G101_n_spl_11
  );


  buf

  (
    G100_p_spl_,
    G100_p
  );


  buf

  (
    G100_p_spl_0,
    G100_p_spl_
  );


  buf

  (
    G100_p_spl_00,
    G100_p_spl_0
  );


  buf

  (
    G100_p_spl_000,
    G100_p_spl_00
  );


  buf

  (
    G100_p_spl_0000,
    G100_p_spl_000
  );


  buf

  (
    G100_p_spl_001,
    G100_p_spl_00
  );


  buf

  (
    G100_p_spl_01,
    G100_p_spl_0
  );


  buf

  (
    G100_p_spl_010,
    G100_p_spl_01
  );


  buf

  (
    G100_p_spl_011,
    G100_p_spl_01
  );


  buf

  (
    G100_p_spl_1,
    G100_p_spl_
  );


  buf

  (
    G100_p_spl_10,
    G100_p_spl_1
  );


  buf

  (
    G100_p_spl_100,
    G100_p_spl_10
  );


  buf

  (
    G100_p_spl_101,
    G100_p_spl_10
  );


  buf

  (
    G100_p_spl_11,
    G100_p_spl_1
  );


  buf

  (
    G100_p_spl_110,
    G100_p_spl_11
  );


  buf

  (
    G100_p_spl_111,
    G100_p_spl_11
  );


  buf

  (
    G100_n_spl_,
    G100_n
  );


  buf

  (
    G100_n_spl_0,
    G100_n_spl_
  );


  buf

  (
    G100_n_spl_00,
    G100_n_spl_0
  );


  buf

  (
    G100_n_spl_000,
    G100_n_spl_00
  );


  buf

  (
    G100_n_spl_0000,
    G100_n_spl_000
  );


  buf

  (
    G100_n_spl_001,
    G100_n_spl_00
  );


  buf

  (
    G100_n_spl_01,
    G100_n_spl_0
  );


  buf

  (
    G100_n_spl_010,
    G100_n_spl_01
  );


  buf

  (
    G100_n_spl_011,
    G100_n_spl_01
  );


  buf

  (
    G100_n_spl_1,
    G100_n_spl_
  );


  buf

  (
    G100_n_spl_10,
    G100_n_spl_1
  );


  buf

  (
    G100_n_spl_100,
    G100_n_spl_10
  );


  buf

  (
    G100_n_spl_101,
    G100_n_spl_10
  );


  buf

  (
    G100_n_spl_11,
    G100_n_spl_1
  );


  buf

  (
    G100_n_spl_110,
    G100_n_spl_11
  );


  buf

  (
    G100_n_spl_111,
    G100_n_spl_11
  );


  buf

  (
    g240_p_spl_,
    g240_p
  );


  buf

  (
    g237_n_spl_,
    g237_n
  );


  buf

  (
    g237_n_spl_0,
    g237_n_spl_
  );


  buf

  (
    g237_n_spl_1,
    g237_n_spl_
  );


  buf

  (
    g240_n_spl_,
    g240_n
  );


  buf

  (
    g240_n_spl_0,
    g240_n_spl_
  );


  buf

  (
    g237_p_spl_,
    g237_p
  );


  buf

  (
    g241_n_spl_,
    g241_n
  );


  buf

  (
    G130_p_spl_,
    G130_p
  );


  buf

  (
    G130_p_spl_0,
    G130_p_spl_
  );


  buf

  (
    G130_p_spl_00,
    G130_p_spl_0
  );


  buf

  (
    G130_p_spl_1,
    G130_p_spl_
  );


  buf

  (
    G130_n_spl_,
    G130_n
  );


  buf

  (
    G130_n_spl_0,
    G130_n_spl_
  );


  buf

  (
    G130_n_spl_00,
    G130_n_spl_0
  );


  buf

  (
    G130_n_spl_1,
    G130_n_spl_
  );


  buf

  (
    G148_n_spl_,
    G148_n
  );


  buf

  (
    G148_n_spl_0,
    G148_n_spl_
  );


  buf

  (
    G148_n_spl_00,
    G148_n_spl_0
  );


  buf

  (
    G148_n_spl_1,
    G148_n_spl_
  );


  buf

  (
    G148_p_spl_,
    G148_p
  );


  buf

  (
    G148_p_spl_0,
    G148_p_spl_
  );


  buf

  (
    G148_p_spl_00,
    G148_p_spl_0
  );


  buf

  (
    G148_p_spl_1,
    G148_p_spl_
  );


  buf

  (
    g248_n_spl_,
    g248_n
  );


  buf

  (
    g245_n_spl_,
    g245_n
  );


  buf

  (
    g245_n_spl_0,
    g245_n_spl_
  );


  buf

  (
    g245_n_spl_1,
    g245_n_spl_
  );


  buf

  (
    G119_p_spl_,
    G119_p
  );


  buf

  (
    G119_p_spl_0,
    G119_p_spl_
  );


  buf

  (
    G119_p_spl_00,
    G119_p_spl_0
  );


  buf

  (
    G119_p_spl_01,
    G119_p_spl_0
  );


  buf

  (
    G119_p_spl_1,
    G119_p_spl_
  );


  buf

  (
    G119_p_spl_10,
    G119_p_spl_1
  );


  buf

  (
    G119_n_spl_,
    G119_n
  );


  buf

  (
    G119_n_spl_0,
    G119_n_spl_
  );


  buf

  (
    G119_n_spl_00,
    G119_n_spl_0
  );


  buf

  (
    G119_n_spl_01,
    G119_n_spl_0
  );


  buf

  (
    G119_n_spl_1,
    G119_n_spl_
  );


  buf

  (
    G119_n_spl_10,
    G119_n_spl_1
  );


  buf

  (
    G146_p_spl_,
    G146_p
  );


  buf

  (
    G146_p_spl_0,
    G146_p_spl_
  );


  buf

  (
    G146_p_spl_1,
    G146_p_spl_
  );


  buf

  (
    G146_n_spl_,
    G146_n
  );


  buf

  (
    G146_n_spl_0,
    G146_n_spl_
  );


  buf

  (
    G146_n_spl_1,
    G146_n_spl_
  );


  buf

  (
    G117_p_spl_,
    G117_p
  );


  buf

  (
    G117_p_spl_0,
    G117_p_spl_
  );


  buf

  (
    G117_p_spl_00,
    G117_p_spl_0
  );


  buf

  (
    G117_p_spl_01,
    G117_p_spl_0
  );


  buf

  (
    G117_p_spl_1,
    G117_p_spl_
  );


  buf

  (
    G117_p_spl_10,
    G117_p_spl_1
  );


  buf

  (
    G117_n_spl_,
    G117_n
  );


  buf

  (
    G117_n_spl_0,
    G117_n_spl_
  );


  buf

  (
    G117_n_spl_00,
    G117_n_spl_0
  );


  buf

  (
    G117_n_spl_01,
    G117_n_spl_0
  );


  buf

  (
    G117_n_spl_1,
    G117_n_spl_
  );


  buf

  (
    G117_n_spl_10,
    G117_n_spl_1
  );


  buf

  (
    G145_p_spl_,
    G145_p
  );


  buf

  (
    G145_p_spl_0,
    G145_p_spl_
  );


  buf

  (
    G145_p_spl_1,
    G145_p_spl_
  );


  buf

  (
    G145_n_spl_,
    G145_n
  );


  buf

  (
    G145_n_spl_0,
    G145_n_spl_
  );


  buf

  (
    G145_n_spl_1,
    G145_n_spl_
  );


  buf

  (
    g267_p_spl_,
    g267_p
  );


  buf

  (
    g258_p_spl_,
    g258_p
  );


  buf

  (
    g267_n_spl_,
    g267_n
  );


  buf

  (
    g267_n_spl_0,
    g267_n_spl_
  );


  buf

  (
    g258_n_spl_,
    g258_n
  );


  buf

  (
    g258_n_spl_0,
    g258_n_spl_
  );


  buf

  (
    G121_p_spl_,
    G121_p
  );


  buf

  (
    G121_p_spl_0,
    G121_p_spl_
  );


  buf

  (
    G121_p_spl_00,
    G121_p_spl_0
  );


  buf

  (
    G121_p_spl_000,
    G121_p_spl_00
  );


  buf

  (
    G121_p_spl_01,
    G121_p_spl_0
  );


  buf

  (
    G121_p_spl_1,
    G121_p_spl_
  );


  buf

  (
    G121_p_spl_10,
    G121_p_spl_1
  );


  buf

  (
    G121_p_spl_11,
    G121_p_spl_1
  );


  buf

  (
    G121_n_spl_,
    G121_n
  );


  buf

  (
    G121_n_spl_0,
    G121_n_spl_
  );


  buf

  (
    G121_n_spl_00,
    G121_n_spl_0
  );


  buf

  (
    G121_n_spl_000,
    G121_n_spl_00
  );


  buf

  (
    G121_n_spl_01,
    G121_n_spl_0
  );


  buf

  (
    G121_n_spl_1,
    G121_n_spl_
  );


  buf

  (
    G121_n_spl_10,
    G121_n_spl_1
  );


  buf

  (
    G121_n_spl_11,
    G121_n_spl_1
  );


  buf

  (
    G147_p_spl_,
    G147_p
  );


  buf

  (
    G147_p_spl_0,
    G147_p_spl_
  );


  buf

  (
    G147_p_spl_00,
    G147_p_spl_0
  );


  buf

  (
    G147_p_spl_1,
    G147_p_spl_
  );


  buf

  (
    G147_n_spl_,
    G147_n
  );


  buf

  (
    G147_n_spl_0,
    G147_n_spl_
  );


  buf

  (
    G147_n_spl_00,
    G147_n_spl_0
  );


  buf

  (
    G147_n_spl_1,
    G147_n_spl_
  );


  buf

  (
    g277_n_spl_,
    g277_n
  );


  buf

  (
    g268_n_spl_,
    g268_n
  );


  buf

  (
    G107_p_spl_,
    G107_p
  );


  buf

  (
    G107_p_spl_0,
    G107_p_spl_
  );


  buf

  (
    G107_p_spl_00,
    G107_p_spl_0
  );


  buf

  (
    G107_p_spl_000,
    G107_p_spl_00
  );


  buf

  (
    G107_p_spl_01,
    G107_p_spl_0
  );


  buf

  (
    G107_p_spl_1,
    G107_p_spl_
  );


  buf

  (
    G107_p_spl_10,
    G107_p_spl_1
  );


  buf

  (
    G107_p_spl_11,
    G107_p_spl_1
  );


  buf

  (
    G107_n_spl_,
    G107_n
  );


  buf

  (
    G107_n_spl_0,
    G107_n_spl_
  );


  buf

  (
    G107_n_spl_00,
    G107_n_spl_0
  );


  buf

  (
    G107_n_spl_000,
    G107_n_spl_00
  );


  buf

  (
    G107_n_spl_01,
    G107_n_spl_0
  );


  buf

  (
    G107_n_spl_1,
    G107_n_spl_
  );


  buf

  (
    G107_n_spl_10,
    G107_n_spl_1
  );


  buf

  (
    G107_n_spl_11,
    G107_n_spl_1
  );


  buf

  (
    G139_p_spl_,
    G139_p
  );


  buf

  (
    G139_p_spl_0,
    G139_p_spl_
  );


  buf

  (
    G139_p_spl_00,
    G139_p_spl_0
  );


  buf

  (
    G139_p_spl_1,
    G139_p_spl_
  );


  buf

  (
    G139_n_spl_,
    G139_n
  );


  buf

  (
    G139_n_spl_0,
    G139_n_spl_
  );


  buf

  (
    G139_n_spl_00,
    G139_n_spl_0
  );


  buf

  (
    G139_n_spl_1,
    G139_n_spl_
  );


  buf

  (
    G105_p_spl_,
    G105_p
  );


  buf

  (
    G105_p_spl_0,
    G105_p_spl_
  );


  buf

  (
    G105_p_spl_00,
    G105_p_spl_0
  );


  buf

  (
    G105_p_spl_000,
    G105_p_spl_00
  );


  buf

  (
    G105_p_spl_01,
    G105_p_spl_0
  );


  buf

  (
    G105_p_spl_1,
    G105_p_spl_
  );


  buf

  (
    G105_p_spl_10,
    G105_p_spl_1
  );


  buf

  (
    G105_p_spl_11,
    G105_p_spl_1
  );


  buf

  (
    G105_n_spl_,
    G105_n
  );


  buf

  (
    G105_n_spl_0,
    G105_n_spl_
  );


  buf

  (
    G105_n_spl_00,
    G105_n_spl_0
  );


  buf

  (
    G105_n_spl_000,
    G105_n_spl_00
  );


  buf

  (
    G105_n_spl_01,
    G105_n_spl_0
  );


  buf

  (
    G105_n_spl_1,
    G105_n_spl_
  );


  buf

  (
    G105_n_spl_10,
    G105_n_spl_1
  );


  buf

  (
    G105_n_spl_11,
    G105_n_spl_1
  );


  buf

  (
    G138_p_spl_,
    G138_p
  );


  buf

  (
    G138_p_spl_0,
    G138_p_spl_
  );


  buf

  (
    G138_p_spl_00,
    G138_p_spl_0
  );


  buf

  (
    G138_p_spl_1,
    G138_p_spl_
  );


  buf

  (
    G138_n_spl_,
    G138_n
  );


  buf

  (
    G138_n_spl_0,
    G138_n_spl_
  );


  buf

  (
    G138_n_spl_00,
    G138_n_spl_0
  );


  buf

  (
    G138_n_spl_1,
    G138_n_spl_
  );


  buf

  (
    g298_n_spl_,
    g298_n
  );


  buf

  (
    g289_n_spl_,
    g289_n
  );


  buf

  (
    G109_p_spl_,
    G109_p
  );


  buf

  (
    G109_p_spl_0,
    G109_p_spl_
  );


  buf

  (
    G109_p_spl_00,
    G109_p_spl_0
  );


  buf

  (
    G109_p_spl_000,
    G109_p_spl_00
  );


  buf

  (
    G109_p_spl_01,
    G109_p_spl_0
  );


  buf

  (
    G109_p_spl_1,
    G109_p_spl_
  );


  buf

  (
    G109_p_spl_10,
    G109_p_spl_1
  );


  buf

  (
    G109_p_spl_11,
    G109_p_spl_1
  );


  buf

  (
    G109_n_spl_,
    G109_n
  );


  buf

  (
    G109_n_spl_0,
    G109_n_spl_
  );


  buf

  (
    G109_n_spl_00,
    G109_n_spl_0
  );


  buf

  (
    G109_n_spl_000,
    G109_n_spl_00
  );


  buf

  (
    G109_n_spl_01,
    G109_n_spl_0
  );


  buf

  (
    G109_n_spl_1,
    G109_n_spl_
  );


  buf

  (
    G109_n_spl_10,
    G109_n_spl_1
  );


  buf

  (
    G109_n_spl_11,
    G109_n_spl_1
  );


  buf

  (
    G135_p_spl_,
    G135_p
  );


  buf

  (
    G135_p_spl_0,
    G135_p_spl_
  );


  buf

  (
    G135_p_spl_00,
    G135_p_spl_0
  );


  buf

  (
    G135_p_spl_1,
    G135_p_spl_
  );


  buf

  (
    G135_n_spl_,
    G135_n
  );


  buf

  (
    G135_n_spl_0,
    G135_n_spl_
  );


  buf

  (
    G135_n_spl_00,
    G135_n_spl_0
  );


  buf

  (
    G135_n_spl_1,
    G135_n_spl_
  );


  buf

  (
    G88_p_spl_,
    G88_p
  );


  buf

  (
    G88_p_spl_0,
    G88_p_spl_
  );


  buf

  (
    G88_p_spl_00,
    G88_p_spl_0
  );


  buf

  (
    G88_p_spl_01,
    G88_p_spl_0
  );


  buf

  (
    G88_p_spl_1,
    G88_p_spl_
  );


  buf

  (
    G88_p_spl_10,
    G88_p_spl_1
  );


  buf

  (
    G88_n_spl_,
    G88_n
  );


  buf

  (
    G88_n_spl_0,
    G88_n_spl_
  );


  buf

  (
    G88_n_spl_00,
    G88_n_spl_0
  );


  buf

  (
    G88_n_spl_01,
    G88_n_spl_0
  );


  buf

  (
    G88_n_spl_1,
    G88_n_spl_
  );


  buf

  (
    G88_n_spl_10,
    G88_n_spl_1
  );


  buf

  (
    G142_p_spl_,
    G142_p
  );


  buf

  (
    G142_p_spl_0,
    G142_p_spl_
  );


  buf

  (
    G142_p_spl_1,
    G142_p_spl_
  );


  buf

  (
    G142_n_spl_,
    G142_n
  );


  buf

  (
    G142_n_spl_0,
    G142_n_spl_
  );


  buf

  (
    G142_n_spl_1,
    G142_n_spl_
  );


  buf

  (
    g317_n_spl_,
    g317_n
  );


  buf

  (
    g317_n_spl_0,
    g317_n_spl_
  );


  buf

  (
    g317_n_spl_1,
    g317_n_spl_
  );


  buf

  (
    g308_n_spl_,
    g308_n
  );


  buf

  (
    G90_p_spl_,
    G90_p
  );


  buf

  (
    G90_p_spl_0,
    G90_p_spl_
  );


  buf

  (
    G90_p_spl_00,
    G90_p_spl_0
  );


  buf

  (
    G90_p_spl_000,
    G90_p_spl_00
  );


  buf

  (
    G90_p_spl_01,
    G90_p_spl_0
  );


  buf

  (
    G90_p_spl_1,
    G90_p_spl_
  );


  buf

  (
    G90_p_spl_10,
    G90_p_spl_1
  );


  buf

  (
    G90_p_spl_11,
    G90_p_spl_1
  );


  buf

  (
    G90_n_spl_,
    G90_n
  );


  buf

  (
    G90_n_spl_0,
    G90_n_spl_
  );


  buf

  (
    G90_n_spl_00,
    G90_n_spl_0
  );


  buf

  (
    G90_n_spl_000,
    G90_n_spl_00
  );


  buf

  (
    G90_n_spl_01,
    G90_n_spl_0
  );


  buf

  (
    G90_n_spl_1,
    G90_n_spl_
  );


  buf

  (
    G90_n_spl_10,
    G90_n_spl_1
  );


  buf

  (
    G90_n_spl_11,
    G90_n_spl_1
  );


  buf

  (
    G143_p_spl_,
    G143_p
  );


  buf

  (
    G143_p_spl_0,
    G143_p_spl_
  );


  buf

  (
    G143_p_spl_00,
    G143_p_spl_0
  );


  buf

  (
    G143_p_spl_1,
    G143_p_spl_
  );


  buf

  (
    G143_n_spl_,
    G143_n
  );


  buf

  (
    G143_n_spl_0,
    G143_n_spl_
  );


  buf

  (
    G143_n_spl_00,
    G143_n_spl_0
  );


  buf

  (
    G143_n_spl_1,
    G143_n_spl_
  );


  buf

  (
    G92_p_spl_,
    G92_p
  );


  buf

  (
    G92_p_spl_0,
    G92_p_spl_
  );


  buf

  (
    G92_p_spl_00,
    G92_p_spl_0
  );


  buf

  (
    G92_p_spl_000,
    G92_p_spl_00
  );


  buf

  (
    G92_p_spl_01,
    G92_p_spl_0
  );


  buf

  (
    G92_p_spl_1,
    G92_p_spl_
  );


  buf

  (
    G92_p_spl_10,
    G92_p_spl_1
  );


  buf

  (
    G92_p_spl_11,
    G92_p_spl_1
  );


  buf

  (
    G92_n_spl_,
    G92_n
  );


  buf

  (
    G92_n_spl_0,
    G92_n_spl_
  );


  buf

  (
    G92_n_spl_00,
    G92_n_spl_0
  );


  buf

  (
    G92_n_spl_000,
    G92_n_spl_00
  );


  buf

  (
    G92_n_spl_01,
    G92_n_spl_0
  );


  buf

  (
    G92_n_spl_1,
    G92_n_spl_
  );


  buf

  (
    G92_n_spl_10,
    G92_n_spl_1
  );


  buf

  (
    G92_n_spl_11,
    G92_n_spl_1
  );


  buf

  (
    G144_p_spl_,
    G144_p
  );


  buf

  (
    G144_p_spl_0,
    G144_p_spl_
  );


  buf

  (
    G144_p_spl_00,
    G144_p_spl_0
  );


  buf

  (
    G144_p_spl_1,
    G144_p_spl_
  );


  buf

  (
    G144_n_spl_,
    G144_n
  );


  buf

  (
    G144_n_spl_0,
    G144_n_spl_
  );


  buf

  (
    G144_n_spl_00,
    G144_n_spl_0
  );


  buf

  (
    G144_n_spl_1,
    G144_n_spl_
  );


  buf

  (
    g337_n_spl_,
    g337_n
  );


  buf

  (
    g328_n_spl_,
    g328_n
  );


  buf

  (
    G94_p_spl_,
    G94_p
  );


  buf

  (
    G94_p_spl_0,
    G94_p_spl_
  );


  buf

  (
    G94_p_spl_00,
    G94_p_spl_0
  );


  buf

  (
    G94_p_spl_000,
    G94_p_spl_00
  );


  buf

  (
    G94_p_spl_01,
    G94_p_spl_0
  );


  buf

  (
    G94_p_spl_1,
    G94_p_spl_
  );


  buf

  (
    G94_p_spl_10,
    G94_p_spl_1
  );


  buf

  (
    G94_p_spl_11,
    G94_p_spl_1
  );


  buf

  (
    G94_n_spl_,
    G94_n
  );


  buf

  (
    G94_n_spl_0,
    G94_n_spl_
  );


  buf

  (
    G94_n_spl_00,
    G94_n_spl_0
  );


  buf

  (
    G94_n_spl_000,
    G94_n_spl_00
  );


  buf

  (
    G94_n_spl_01,
    G94_n_spl_0
  );


  buf

  (
    G94_n_spl_1,
    G94_n_spl_
  );


  buf

  (
    G94_n_spl_10,
    G94_n_spl_1
  );


  buf

  (
    G94_n_spl_11,
    G94_n_spl_1
  );


  buf

  (
    G140_p_spl_,
    G140_p
  );


  buf

  (
    G140_p_spl_0,
    G140_p_spl_
  );


  buf

  (
    G140_p_spl_00,
    G140_p_spl_0
  );


  buf

  (
    G140_p_spl_1,
    G140_p_spl_
  );


  buf

  (
    G140_n_spl_,
    G140_n
  );


  buf

  (
    G140_n_spl_0,
    G140_n_spl_
  );


  buf

  (
    G140_n_spl_00,
    G140_n_spl_0
  );


  buf

  (
    G140_n_spl_1,
    G140_n_spl_
  );


  buf

  (
    G96_p_spl_,
    G96_p
  );


  buf

  (
    G96_p_spl_0,
    G96_p_spl_
  );


  buf

  (
    G96_p_spl_00,
    G96_p_spl_0
  );


  buf

  (
    G96_p_spl_000,
    G96_p_spl_00
  );


  buf

  (
    G96_p_spl_01,
    G96_p_spl_0
  );


  buf

  (
    G96_p_spl_1,
    G96_p_spl_
  );


  buf

  (
    G96_p_spl_10,
    G96_p_spl_1
  );


  buf

  (
    G96_p_spl_11,
    G96_p_spl_1
  );


  buf

  (
    G96_n_spl_,
    G96_n
  );


  buf

  (
    G96_n_spl_0,
    G96_n_spl_
  );


  buf

  (
    G96_n_spl_00,
    G96_n_spl_0
  );


  buf

  (
    G96_n_spl_000,
    G96_n_spl_00
  );


  buf

  (
    G96_n_spl_01,
    G96_n_spl_0
  );


  buf

  (
    G96_n_spl_1,
    G96_n_spl_
  );


  buf

  (
    G96_n_spl_10,
    G96_n_spl_1
  );


  buf

  (
    G96_n_spl_11,
    G96_n_spl_1
  );


  buf

  (
    G141_p_spl_,
    G141_p
  );


  buf

  (
    G141_p_spl_0,
    G141_p_spl_
  );


  buf

  (
    G141_p_spl_00,
    G141_p_spl_0
  );


  buf

  (
    G141_p_spl_1,
    G141_p_spl_
  );


  buf

  (
    G141_n_spl_,
    G141_n
  );


  buf

  (
    G141_n_spl_0,
    G141_n_spl_
  );


  buf

  (
    G141_n_spl_00,
    G141_n_spl_0
  );


  buf

  (
    G141_n_spl_1,
    G141_n_spl_
  );


  buf

  (
    G103_p_spl_,
    G103_p
  );


  buf

  (
    G103_p_spl_0,
    G103_p_spl_
  );


  buf

  (
    G103_p_spl_00,
    G103_p_spl_0
  );


  buf

  (
    G103_p_spl_000,
    G103_p_spl_00
  );


  buf

  (
    G103_p_spl_01,
    G103_p_spl_0
  );


  buf

  (
    G103_p_spl_1,
    G103_p_spl_
  );


  buf

  (
    G103_p_spl_10,
    G103_p_spl_1
  );


  buf

  (
    G103_p_spl_11,
    G103_p_spl_1
  );


  buf

  (
    G103_n_spl_,
    G103_n
  );


  buf

  (
    G103_n_spl_0,
    G103_n_spl_
  );


  buf

  (
    G103_n_spl_00,
    G103_n_spl_0
  );


  buf

  (
    G103_n_spl_000,
    G103_n_spl_00
  );


  buf

  (
    G103_n_spl_01,
    G103_n_spl_0
  );


  buf

  (
    G103_n_spl_1,
    G103_n_spl_
  );


  buf

  (
    G103_n_spl_10,
    G103_n_spl_1
  );


  buf

  (
    G103_n_spl_11,
    G103_n_spl_1
  );


  buf

  (
    G137_p_spl_,
    G137_p
  );


  buf

  (
    G137_p_spl_0,
    G137_p_spl_
  );


  buf

  (
    G137_p_spl_00,
    G137_p_spl_0
  );


  buf

  (
    G137_p_spl_1,
    G137_p_spl_
  );


  buf

  (
    G137_n_spl_,
    G137_n
  );


  buf

  (
    G137_n_spl_0,
    G137_n_spl_
  );


  buf

  (
    G137_n_spl_00,
    G137_n_spl_0
  );


  buf

  (
    G137_n_spl_1,
    G137_n_spl_
  );


  buf

  (
    g365_n_spl_,
    g365_n
  );


  buf

  (
    g356_n_spl_,
    g356_n
  );


  buf

  (
    g347_n_spl_,
    g347_n
  );


  buf

  (
    G124_n_spl_,
    G124_n
  );


  buf

  (
    G124_n_spl_0,
    G124_n_spl_
  );


  buf

  (
    G124_n_spl_00,
    G124_n_spl_0
  );


  buf

  (
    G124_n_spl_000,
    G124_n_spl_00
  );


  buf

  (
    G124_n_spl_0000,
    G124_n_spl_000
  );


  buf

  (
    G124_n_spl_0001,
    G124_n_spl_000
  );


  buf

  (
    G124_n_spl_001,
    G124_n_spl_00
  );


  buf

  (
    G124_n_spl_0010,
    G124_n_spl_001
  );


  buf

  (
    G124_n_spl_0011,
    G124_n_spl_001
  );


  buf

  (
    G124_n_spl_01,
    G124_n_spl_0
  );


  buf

  (
    G124_n_spl_010,
    G124_n_spl_01
  );


  buf

  (
    G124_n_spl_011,
    G124_n_spl_01
  );


  buf

  (
    G124_n_spl_1,
    G124_n_spl_
  );


  buf

  (
    G124_n_spl_10,
    G124_n_spl_1
  );


  buf

  (
    G124_n_spl_100,
    G124_n_spl_10
  );


  buf

  (
    G124_n_spl_101,
    G124_n_spl_10
  );


  buf

  (
    G124_n_spl_11,
    G124_n_spl_1
  );


  buf

  (
    G124_n_spl_110,
    G124_n_spl_11
  );


  buf

  (
    G124_n_spl_111,
    G124_n_spl_11
  );


  buf

  (
    G124_p_spl_,
    G124_p
  );


  buf

  (
    G124_p_spl_0,
    G124_p_spl_
  );


  buf

  (
    G124_p_spl_00,
    G124_p_spl_0
  );


  buf

  (
    G124_p_spl_000,
    G124_p_spl_00
  );


  buf

  (
    G124_p_spl_0000,
    G124_p_spl_000
  );


  buf

  (
    G124_p_spl_0001,
    G124_p_spl_000
  );


  buf

  (
    G124_p_spl_001,
    G124_p_spl_00
  );


  buf

  (
    G124_p_spl_0010,
    G124_p_spl_001
  );


  buf

  (
    G124_p_spl_0011,
    G124_p_spl_001
  );


  buf

  (
    G124_p_spl_01,
    G124_p_spl_0
  );


  buf

  (
    G124_p_spl_010,
    G124_p_spl_01
  );


  buf

  (
    G124_p_spl_011,
    G124_p_spl_01
  );


  buf

  (
    G124_p_spl_1,
    G124_p_spl_
  );


  buf

  (
    G124_p_spl_10,
    G124_p_spl_1
  );


  buf

  (
    G124_p_spl_100,
    G124_p_spl_10
  );


  buf

  (
    G124_p_spl_101,
    G124_p_spl_10
  );


  buf

  (
    G124_p_spl_11,
    G124_p_spl_1
  );


  buf

  (
    G124_p_spl_110,
    G124_p_spl_11
  );


  buf

  (
    G124_p_spl_111,
    G124_p_spl_11
  );


  buf

  (
    g372_p_spl_,
    g372_p
  );


  buf

  (
    g372_p_spl_0,
    g372_p_spl_
  );


  buf

  (
    g372_p_spl_1,
    g372_p_spl_
  );


  buf

  (
    g372_n_spl_,
    g372_n
  );


  buf

  (
    g372_n_spl_0,
    g372_n_spl_
  );


  buf

  (
    g372_n_spl_1,
    g372_n_spl_
  );


  buf

  (
    g374_n_spl_,
    g374_n
  );


  buf

  (
    g374_n_spl_0,
    g374_n_spl_
  );


  buf

  (
    g374_n_spl_1,
    g374_n_spl_
  );


  buf

  (
    g373_n_spl_,
    g373_n
  );


  buf

  (
    g373_n_spl_0,
    g373_n_spl_
  );


  buf

  (
    g374_p_spl_,
    g374_p
  );


  buf

  (
    g374_p_spl_0,
    g374_p_spl_
  );


  buf

  (
    g374_p_spl_1,
    g374_p_spl_
  );


  buf

  (
    g373_p_spl_,
    g373_p
  );


  buf

  (
    g373_p_spl_0,
    g373_p_spl_
  );


  buf

  (
    g378_p_spl_,
    g378_p
  );


  buf

  (
    g378_p_spl_0,
    g378_p_spl_
  );


  buf

  (
    g378_p_spl_1,
    g378_p_spl_
  );


  buf

  (
    g378_n_spl_,
    g378_n
  );


  buf

  (
    g378_n_spl_0,
    g378_n_spl_
  );


  buf

  (
    g378_n_spl_1,
    g378_n_spl_
  );


  buf

  (
    g380_n_spl_,
    g380_n
  );


  buf

  (
    g379_n_spl_,
    g379_n
  );


  buf

  (
    g380_p_spl_,
    g380_p
  );


  buf

  (
    g379_p_spl_,
    g379_p
  );


  buf

  (
    g381_p_spl_,
    g381_p
  );


  buf

  (
    g381_p_spl_0,
    g381_p_spl_
  );


  buf

  (
    g381_p_spl_00,
    g381_p_spl_0
  );


  buf

  (
    g381_p_spl_01,
    g381_p_spl_0
  );


  buf

  (
    g381_p_spl_1,
    g381_p_spl_
  );


  buf

  (
    g381_p_spl_10,
    g381_p_spl_1
  );


  buf

  (
    g375_p_spl_,
    g375_p
  );


  buf

  (
    g375_p_spl_0,
    g375_p_spl_
  );


  buf

  (
    g375_p_spl_00,
    g375_p_spl_0
  );


  buf

  (
    g375_p_spl_1,
    g375_p_spl_
  );


  buf

  (
    g381_n_spl_,
    g381_n
  );


  buf

  (
    g381_n_spl_0,
    g381_n_spl_
  );


  buf

  (
    g381_n_spl_00,
    g381_n_spl_0
  );


  buf

  (
    g381_n_spl_01,
    g381_n_spl_0
  );


  buf

  (
    g381_n_spl_1,
    g381_n_spl_
  );


  buf

  (
    g381_n_spl_10,
    g381_n_spl_1
  );


  buf

  (
    g375_n_spl_,
    g375_n
  );


  buf

  (
    g375_n_spl_0,
    g375_n_spl_
  );


  buf

  (
    g375_n_spl_00,
    g375_n_spl_0
  );


  buf

  (
    g375_n_spl_1,
    g375_n_spl_
  );


  buf

  (
    g385_p_spl_,
    g385_p
  );


  buf

  (
    g385_p_spl_0,
    g385_p_spl_
  );


  buf

  (
    g385_p_spl_1,
    g385_p_spl_
  );


  buf

  (
    g385_n_spl_,
    g385_n
  );


  buf

  (
    g385_n_spl_0,
    g385_n_spl_
  );


  buf

  (
    g385_n_spl_1,
    g385_n_spl_
  );


  buf

  (
    g387_n_spl_,
    g387_n
  );


  buf

  (
    g386_n_spl_,
    g386_n
  );


  buf

  (
    g387_p_spl_,
    g387_p
  );


  buf

  (
    g386_p_spl_,
    g386_p
  );


  buf

  (
    g388_p_spl_,
    g388_p
  );


  buf

  (
    g388_p_spl_0,
    g388_p_spl_
  );


  buf

  (
    g388_p_spl_00,
    g388_p_spl_0
  );


  buf

  (
    g388_p_spl_01,
    g388_p_spl_0
  );


  buf

  (
    g388_p_spl_1,
    g388_p_spl_
  );


  buf

  (
    g382_p_spl_,
    g382_p
  );


  buf

  (
    g388_n_spl_,
    g388_n
  );


  buf

  (
    g388_n_spl_0,
    g388_n_spl_
  );


  buf

  (
    g388_n_spl_00,
    g388_n_spl_0
  );


  buf

  (
    g388_n_spl_01,
    g388_n_spl_0
  );


  buf

  (
    g388_n_spl_1,
    g388_n_spl_
  );


  buf

  (
    g382_n_spl_,
    g382_n
  );


  buf

  (
    g392_p_spl_,
    g392_p
  );


  buf

  (
    g392_p_spl_0,
    g392_p_spl_
  );


  buf

  (
    g392_p_spl_1,
    g392_p_spl_
  );


  buf

  (
    g392_n_spl_,
    g392_n
  );


  buf

  (
    g392_n_spl_0,
    g392_n_spl_
  );


  buf

  (
    g392_n_spl_1,
    g392_n_spl_
  );


  buf

  (
    g393_n_spl_,
    g393_n
  );


  buf

  (
    g395_n_spl_,
    g395_n
  );


  buf

  (
    g395_n_spl_0,
    g395_n_spl_
  );


  buf

  (
    g395_n_spl_00,
    g395_n_spl_0
  );


  buf

  (
    g395_n_spl_01,
    g395_n_spl_0
  );


  buf

  (
    g395_n_spl_1,
    g395_n_spl_
  );


  buf

  (
    g395_n_spl_10,
    g395_n_spl_1
  );


  buf

  (
    g389_n_spl_,
    g389_n
  );


  buf

  (
    g389_n_spl_0,
    g389_n_spl_
  );


  buf

  (
    g399_p_spl_,
    g399_p
  );


  buf

  (
    g399_p_spl_0,
    g399_p_spl_
  );


  buf

  (
    g399_p_spl_1,
    g399_p_spl_
  );


  buf

  (
    g399_n_spl_,
    g399_n
  );


  buf

  (
    g399_n_spl_0,
    g399_n_spl_
  );


  buf

  (
    g399_n_spl_1,
    g399_n_spl_
  );


  buf

  (
    g401_n_spl_,
    g401_n
  );


  buf

  (
    g401_n_spl_0,
    g401_n_spl_
  );


  buf

  (
    g400_n_spl_,
    g400_n
  );


  buf

  (
    g400_n_spl_0,
    g400_n_spl_
  );


  buf

  (
    g400_n_spl_00,
    g400_n_spl_0
  );


  buf

  (
    g400_n_spl_1,
    g400_n_spl_
  );


  buf

  (
    g401_p_spl_,
    g401_p
  );


  buf

  (
    g401_p_spl_0,
    g401_p_spl_
  );


  buf

  (
    g400_p_spl_,
    g400_p
  );


  buf

  (
    g400_p_spl_0,
    g400_p_spl_
  );


  buf

  (
    g400_p_spl_00,
    g400_p_spl_0
  );


  buf

  (
    g400_p_spl_1,
    g400_p_spl_
  );


  buf

  (
    g405_p_spl_,
    g405_p
  );


  buf

  (
    g405_p_spl_0,
    g405_p_spl_
  );


  buf

  (
    g405_p_spl_1,
    g405_p_spl_
  );


  buf

  (
    g405_n_spl_,
    g405_n
  );


  buf

  (
    g405_n_spl_0,
    g405_n_spl_
  );


  buf

  (
    g405_n_spl_1,
    g405_n_spl_
  );


  buf

  (
    g406_n_spl_,
    g406_n
  );


  buf

  (
    g406_n_spl_0,
    g406_n_spl_
  );


  buf

  (
    g406_p_spl_,
    g406_p
  );


  buf

  (
    g406_p_spl_0,
    g406_p_spl_
  );


  buf

  (
    g408_p_spl_,
    g408_p
  );


  buf

  (
    g408_p_spl_0,
    g408_p_spl_
  );


  buf

  (
    g408_p_spl_1,
    g408_p_spl_
  );


  buf

  (
    g402_p_spl_,
    g402_p
  );


  buf

  (
    g402_p_spl_0,
    g402_p_spl_
  );


  buf

  (
    g402_p_spl_1,
    g402_p_spl_
  );


  buf

  (
    g408_n_spl_,
    g408_n
  );


  buf

  (
    g408_n_spl_0,
    g408_n_spl_
  );


  buf

  (
    g408_n_spl_00,
    g408_n_spl_0
  );


  buf

  (
    g408_n_spl_1,
    g408_n_spl_
  );


  buf

  (
    g402_n_spl_,
    g402_n
  );


  buf

  (
    g402_n_spl_0,
    g402_n_spl_
  );


  buf

  (
    g412_p_spl_,
    g412_p
  );


  buf

  (
    g412_p_spl_0,
    g412_p_spl_
  );


  buf

  (
    g412_p_spl_1,
    g412_p_spl_
  );


  buf

  (
    g412_n_spl_,
    g412_n
  );


  buf

  (
    g412_n_spl_0,
    g412_n_spl_
  );


  buf

  (
    g412_n_spl_1,
    g412_n_spl_
  );


  buf

  (
    g413_n_spl_,
    g413_n
  );


  buf

  (
    g413_p_spl_,
    g413_p
  );


  buf

  (
    g415_p_spl_,
    g415_p
  );


  buf

  (
    g415_p_spl_0,
    g415_p_spl_
  );


  buf

  (
    g415_p_spl_00,
    g415_p_spl_0
  );


  buf

  (
    g415_p_spl_1,
    g415_p_spl_
  );


  buf

  (
    g409_p_spl_,
    g409_p
  );


  buf

  (
    g409_p_spl_0,
    g409_p_spl_
  );


  buf

  (
    g415_n_spl_,
    g415_n
  );


  buf

  (
    g415_n_spl_0,
    g415_n_spl_
  );


  buf

  (
    g415_n_spl_00,
    g415_n_spl_0
  );


  buf

  (
    g415_n_spl_1,
    g415_n_spl_
  );


  buf

  (
    g409_n_spl_,
    g409_n
  );


  buf

  (
    g409_n_spl_0,
    g409_n_spl_
  );


  buf

  (
    g419_p_spl_,
    g419_p
  );


  buf

  (
    g419_p_spl_0,
    g419_p_spl_
  );


  buf

  (
    g419_p_spl_1,
    g419_p_spl_
  );


  buf

  (
    g419_n_spl_,
    g419_n
  );


  buf

  (
    g419_n_spl_0,
    g419_n_spl_
  );


  buf

  (
    g419_n_spl_1,
    g419_n_spl_
  );


  buf

  (
    g420_n_spl_,
    g420_n
  );


  buf

  (
    g420_n_spl_0,
    g420_n_spl_
  );


  buf

  (
    g420_p_spl_,
    g420_p
  );


  buf

  (
    g420_p_spl_0,
    g420_p_spl_
  );


  buf

  (
    g422_p_spl_,
    g422_p
  );


  buf

  (
    g422_p_spl_0,
    g422_p_spl_
  );


  buf

  (
    g422_p_spl_00,
    g422_p_spl_0
  );


  buf

  (
    g422_p_spl_1,
    g422_p_spl_
  );


  buf

  (
    g416_p_spl_,
    g416_p
  );


  buf

  (
    g416_p_spl_0,
    g416_p_spl_
  );


  buf

  (
    g422_n_spl_,
    g422_n
  );


  buf

  (
    g422_n_spl_0,
    g422_n_spl_
  );


  buf

  (
    g422_n_spl_00,
    g422_n_spl_0
  );


  buf

  (
    g422_n_spl_01,
    g422_n_spl_0
  );


  buf

  (
    g422_n_spl_1,
    g422_n_spl_
  );


  buf

  (
    g416_n_spl_,
    g416_n
  );


  buf

  (
    g416_n_spl_0,
    g416_n_spl_
  );


  buf

  (
    g426_p_spl_,
    g426_p
  );


  buf

  (
    g426_p_spl_0,
    g426_p_spl_
  );


  buf

  (
    g426_p_spl_1,
    g426_p_spl_
  );


  buf

  (
    g426_n_spl_,
    g426_n
  );


  buf

  (
    g426_n_spl_0,
    g426_n_spl_
  );


  buf

  (
    g426_n_spl_1,
    g426_n_spl_
  );


  buf

  (
    g427_n_spl_,
    g427_n
  );


  buf

  (
    g427_p_spl_,
    g427_p
  );


  buf

  (
    g429_p_spl_,
    g429_p
  );


  buf

  (
    g429_p_spl_0,
    g429_p_spl_
  );


  buf

  (
    g429_p_spl_00,
    g429_p_spl_0
  );


  buf

  (
    g429_p_spl_01,
    g429_p_spl_0
  );


  buf

  (
    g429_p_spl_1,
    g429_p_spl_
  );


  buf

  (
    g429_p_spl_10,
    g429_p_spl_1
  );


  buf

  (
    g423_p_spl_,
    g423_p
  );


  buf

  (
    g429_n_spl_,
    g429_n
  );


  buf

  (
    g429_n_spl_0,
    g429_n_spl_
  );


  buf

  (
    g429_n_spl_00,
    g429_n_spl_0
  );


  buf

  (
    g429_n_spl_01,
    g429_n_spl_0
  );


  buf

  (
    g429_n_spl_1,
    g429_n_spl_
  );


  buf

  (
    g429_n_spl_10,
    g429_n_spl_1
  );


  buf

  (
    g423_n_spl_,
    g423_n
  );


  buf

  (
    g430_n_spl_,
    g430_n
  );


  buf

  (
    g430_n_spl_0,
    g430_n_spl_
  );


  buf

  (
    g430_n_spl_1,
    g430_n_spl_
  );


  buf

  (
    g396_n_spl_,
    g396_n
  );


  buf

  (
    G123_n_spl_,
    G123_n
  );


  buf

  (
    G123_n_spl_0,
    G123_n_spl_
  );


  buf

  (
    G123_n_spl_00,
    G123_n_spl_0
  );


  buf

  (
    G123_n_spl_000,
    G123_n_spl_00
  );


  buf

  (
    G123_n_spl_0000,
    G123_n_spl_000
  );


  buf

  (
    G123_n_spl_0001,
    G123_n_spl_000
  );


  buf

  (
    G123_n_spl_001,
    G123_n_spl_00
  );


  buf

  (
    G123_n_spl_0010,
    G123_n_spl_001
  );


  buf

  (
    G123_n_spl_01,
    G123_n_spl_0
  );


  buf

  (
    G123_n_spl_010,
    G123_n_spl_01
  );


  buf

  (
    G123_n_spl_011,
    G123_n_spl_01
  );


  buf

  (
    G123_n_spl_1,
    G123_n_spl_
  );


  buf

  (
    G123_n_spl_10,
    G123_n_spl_1
  );


  buf

  (
    G123_n_spl_100,
    G123_n_spl_10
  );


  buf

  (
    G123_n_spl_101,
    G123_n_spl_10
  );


  buf

  (
    G123_n_spl_11,
    G123_n_spl_1
  );


  buf

  (
    G123_n_spl_110,
    G123_n_spl_11
  );


  buf

  (
    G123_n_spl_111,
    G123_n_spl_11
  );


  buf

  (
    G123_p_spl_,
    G123_p
  );


  buf

  (
    G123_p_spl_0,
    G123_p_spl_
  );


  buf

  (
    G123_p_spl_00,
    G123_p_spl_0
  );


  buf

  (
    G123_p_spl_000,
    G123_p_spl_00
  );


  buf

  (
    G123_p_spl_0000,
    G123_p_spl_000
  );


  buf

  (
    G123_p_spl_0001,
    G123_p_spl_000
  );


  buf

  (
    G123_p_spl_001,
    G123_p_spl_00
  );


  buf

  (
    G123_p_spl_0010,
    G123_p_spl_001
  );


  buf

  (
    G123_p_spl_01,
    G123_p_spl_0
  );


  buf

  (
    G123_p_spl_010,
    G123_p_spl_01
  );


  buf

  (
    G123_p_spl_011,
    G123_p_spl_01
  );


  buf

  (
    G123_p_spl_1,
    G123_p_spl_
  );


  buf

  (
    G123_p_spl_10,
    G123_p_spl_1
  );


  buf

  (
    G123_p_spl_100,
    G123_p_spl_10
  );


  buf

  (
    G123_p_spl_101,
    G123_p_spl_10
  );


  buf

  (
    G123_p_spl_11,
    G123_p_spl_1
  );


  buf

  (
    G123_p_spl_110,
    G123_p_spl_11
  );


  buf

  (
    G123_p_spl_111,
    G123_p_spl_11
  );


  buf

  (
    g434_p_spl_,
    g434_p
  );


  buf

  (
    g434_p_spl_0,
    g434_p_spl_
  );


  buf

  (
    g434_p_spl_1,
    g434_p_spl_
  );


  buf

  (
    g434_n_spl_,
    g434_n
  );


  buf

  (
    g434_n_spl_0,
    g434_n_spl_
  );


  buf

  (
    g434_n_spl_1,
    g434_n_spl_
  );


  buf

  (
    g435_n_spl_,
    g435_n
  );


  buf

  (
    g435_p_spl_,
    g435_p
  );


  buf

  (
    g440_p_spl_,
    g440_p
  );


  buf

  (
    g440_p_spl_0,
    g440_p_spl_
  );


  buf

  (
    g440_p_spl_1,
    g440_p_spl_
  );


  buf

  (
    g440_n_spl_,
    g440_n
  );


  buf

  (
    g440_n_spl_0,
    g440_n_spl_
  );


  buf

  (
    g440_n_spl_1,
    g440_n_spl_
  );


  buf

  (
    g442_n_spl_,
    g442_n
  );


  buf

  (
    g442_n_spl_0,
    g442_n_spl_
  );


  buf

  (
    g442_n_spl_1,
    g442_n_spl_
  );


  buf

  (
    g441_n_spl_,
    g441_n
  );


  buf

  (
    g441_n_spl_0,
    g441_n_spl_
  );


  buf

  (
    g441_n_spl_00,
    g441_n_spl_0
  );


  buf

  (
    g441_n_spl_1,
    g441_n_spl_
  );


  buf

  (
    g442_p_spl_,
    g442_p
  );


  buf

  (
    g442_p_spl_0,
    g442_p_spl_
  );


  buf

  (
    g442_p_spl_1,
    g442_p_spl_
  );


  buf

  (
    g441_p_spl_,
    g441_p
  );


  buf

  (
    g441_p_spl_0,
    g441_p_spl_
  );


  buf

  (
    g441_p_spl_00,
    g441_p_spl_0
  );


  buf

  (
    g441_p_spl_1,
    g441_p_spl_
  );


  buf

  (
    g443_p_spl_,
    g443_p
  );


  buf

  (
    g443_p_spl_0,
    g443_p_spl_
  );


  buf

  (
    g443_p_spl_00,
    g443_p_spl_0
  );


  buf

  (
    g443_p_spl_1,
    g443_p_spl_
  );


  buf

  (
    g437_p_spl_,
    g437_p
  );


  buf

  (
    g437_p_spl_0,
    g437_p_spl_
  );


  buf

  (
    g437_p_spl_00,
    g437_p_spl_0
  );


  buf

  (
    g437_p_spl_01,
    g437_p_spl_0
  );


  buf

  (
    g437_p_spl_1,
    g437_p_spl_
  );


  buf

  (
    g443_n_spl_,
    g443_n
  );


  buf

  (
    g443_n_spl_0,
    g443_n_spl_
  );


  buf

  (
    g443_n_spl_00,
    g443_n_spl_0
  );


  buf

  (
    g443_n_spl_1,
    g443_n_spl_
  );


  buf

  (
    g437_n_spl_,
    g437_n
  );


  buf

  (
    g437_n_spl_0,
    g437_n_spl_
  );


  buf

  (
    g437_n_spl_00,
    g437_n_spl_0
  );


  buf

  (
    g437_n_spl_01,
    g437_n_spl_0
  );


  buf

  (
    g437_n_spl_1,
    g437_n_spl_
  );


  buf

  (
    g447_p_spl_,
    g447_p
  );


  buf

  (
    g447_p_spl_0,
    g447_p_spl_
  );


  buf

  (
    g447_p_spl_1,
    g447_p_spl_
  );


  buf

  (
    g447_n_spl_,
    g447_n
  );


  buf

  (
    g447_n_spl_0,
    g447_n_spl_
  );


  buf

  (
    g447_n_spl_1,
    g447_n_spl_
  );


  buf

  (
    g448_n_spl_,
    g448_n
  );


  buf

  (
    g448_p_spl_,
    g448_p
  );


  buf

  (
    G125_n_spl_,
    G125_n
  );


  buf

  (
    g451_n_spl_,
    g451_n
  );


  buf

  (
    g451_n_spl_0,
    g451_n_spl_
  );


  buf

  (
    g451_n_spl_1,
    g451_n_spl_
  );


  buf

  (
    g451_p_spl_,
    g451_p
  );


  buf

  (
    g451_p_spl_0,
    g451_p_spl_
  );


  buf

  (
    g451_p_spl_1,
    g451_p_spl_
  );


  buf

  (
    g452_n_spl_,
    g452_n
  );


  buf

  (
    g452_n_spl_0,
    g452_n_spl_
  );


  buf

  (
    g452_p_spl_,
    g452_p
  );


  buf

  (
    g452_p_spl_0,
    g452_p_spl_
  );


  buf

  (
    g454_p_spl_,
    g454_p
  );


  buf

  (
    g454_p_spl_0,
    g454_p_spl_
  );


  buf

  (
    g454_p_spl_1,
    g454_p_spl_
  );


  buf

  (
    g450_p_spl_,
    g450_p
  );


  buf

  (
    g450_p_spl_0,
    g450_p_spl_
  );


  buf

  (
    g450_p_spl_1,
    g450_p_spl_
  );


  buf

  (
    g454_n_spl_,
    g454_n
  );


  buf

  (
    g454_n_spl_0,
    g454_n_spl_
  );


  buf

  (
    g454_n_spl_00,
    g454_n_spl_0
  );


  buf

  (
    g454_n_spl_1,
    g454_n_spl_
  );


  buf

  (
    g450_n_spl_,
    g450_n
  );


  buf

  (
    g450_n_spl_0,
    g450_n_spl_
  );


  buf

  (
    g450_n_spl_1,
    g450_n_spl_
  );


  buf

  (
    G129_n_spl_,
    G129_n
  );


  buf

  (
    g458_p_spl_,
    g458_p
  );


  buf

  (
    g458_p_spl_0,
    g458_p_spl_
  );


  buf

  (
    g458_p_spl_1,
    g458_p_spl_
  );


  buf

  (
    g458_n_spl_,
    g458_n
  );


  buf

  (
    g458_n_spl_0,
    g458_n_spl_
  );


  buf

  (
    g458_n_spl_1,
    g458_n_spl_
  );


  buf

  (
    g459_n_spl_,
    g459_n
  );


  buf

  (
    g459_n_spl_0,
    g459_n_spl_
  );


  buf

  (
    g459_p_spl_,
    g459_p
  );


  buf

  (
    g459_p_spl_0,
    g459_p_spl_
  );


  buf

  (
    G131_n_spl_,
    G131_n
  );


  buf

  (
    g464_n_spl_,
    g464_n
  );


  buf

  (
    g464_n_spl_0,
    g464_n_spl_
  );


  buf

  (
    g464_n_spl_00,
    g464_n_spl_0
  );


  buf

  (
    g464_n_spl_01,
    g464_n_spl_0
  );


  buf

  (
    g464_n_spl_1,
    g464_n_spl_
  );


  buf

  (
    g464_n_spl_10,
    g464_n_spl_1
  );


  buf

  (
    g461_p_spl_,
    g461_p
  );


  buf

  (
    g461_p_spl_0,
    g461_p_spl_
  );


  buf

  (
    g464_p_spl_,
    g464_p
  );


  buf

  (
    g464_p_spl_0,
    g464_p_spl_
  );


  buf

  (
    g464_p_spl_00,
    g464_p_spl_0
  );


  buf

  (
    g464_p_spl_01,
    g464_p_spl_0
  );


  buf

  (
    g464_p_spl_1,
    g464_p_spl_
  );


  buf

  (
    g464_p_spl_10,
    g464_p_spl_1
  );


  buf

  (
    g461_n_spl_,
    g461_n
  );


  buf

  (
    g461_n_spl_0,
    g461_n_spl_
  );


  buf

  (
    G127_n_spl_,
    G127_n
  );


  buf

  (
    g468_p_spl_,
    g468_p
  );


  buf

  (
    g468_p_spl_0,
    g468_p_spl_
  );


  buf

  (
    g468_p_spl_1,
    g468_p_spl_
  );


  buf

  (
    g468_n_spl_,
    g468_n
  );


  buf

  (
    g468_n_spl_0,
    g468_n_spl_
  );


  buf

  (
    g468_n_spl_1,
    g468_n_spl_
  );


  buf

  (
    g469_n_spl_,
    g469_n
  );


  buf

  (
    g469_n_spl_0,
    g469_n_spl_
  );


  buf

  (
    g469_p_spl_,
    g469_p
  );


  buf

  (
    g469_p_spl_0,
    g469_p_spl_
  );


  buf

  (
    g471_p_spl_,
    g471_p
  );


  buf

  (
    g471_p_spl_0,
    g471_p_spl_
  );


  buf

  (
    g471_p_spl_1,
    g471_p_spl_
  );


  buf

  (
    g465_p_spl_,
    g465_p
  );


  buf

  (
    g465_p_spl_0,
    g465_p_spl_
  );


  buf

  (
    g471_n_spl_,
    g471_n
  );


  buf

  (
    g471_n_spl_0,
    g471_n_spl_
  );


  buf

  (
    g471_n_spl_00,
    g471_n_spl_0
  );


  buf

  (
    g471_n_spl_1,
    g471_n_spl_
  );


  buf

  (
    g465_n_spl_,
    g465_n
  );


  buf

  (
    g465_n_spl_0,
    g465_n_spl_
  );


  buf

  (
    g472_p_spl_,
    g472_p
  );


  buf

  (
    g455_p_spl_,
    g455_p
  );


  buf

  (
    g472_n_spl_,
    g472_n
  );


  buf

  (
    g455_n_spl_,
    g455_n
  );


  buf

  (
    G114_n_spl_,
    G114_n
  );


  buf

  (
    G114_n_spl_0,
    G114_n_spl_
  );


  buf

  (
    G114_p_spl_,
    G114_p
  );


  buf

  (
    g479_n_spl_,
    g479_n
  );


  buf

  (
    g479_n_spl_0,
    g479_n_spl_
  );


  buf

  (
    g479_n_spl_00,
    g479_n_spl_0
  );


  buf

  (
    g479_n_spl_01,
    g479_n_spl_0
  );


  buf

  (
    g479_n_spl_1,
    g479_n_spl_
  );


  buf

  (
    g479_n_spl_10,
    g479_n_spl_1
  );


  buf

  (
    g476_n_spl_,
    g476_n
  );


  buf

  (
    g476_n_spl_0,
    g476_n_spl_
  );


  buf

  (
    g476_n_spl_1,
    g476_n_spl_
  );


  buf

  (
    g479_p_spl_,
    g479_p
  );


  buf

  (
    g479_p_spl_0,
    g479_p_spl_
  );


  buf

  (
    g479_p_spl_00,
    g479_p_spl_0
  );


  buf

  (
    g479_p_spl_01,
    g479_p_spl_0
  );


  buf

  (
    g479_p_spl_1,
    g479_p_spl_
  );


  buf

  (
    g479_p_spl_10,
    g479_p_spl_1
  );


  buf

  (
    g476_p_spl_,
    g476_p
  );


  buf

  (
    g476_p_spl_0,
    g476_p_spl_
  );


  buf

  (
    g476_p_spl_00,
    g476_p_spl_0
  );


  buf

  (
    g476_p_spl_1,
    g476_p_spl_
  );


  buf

  (
    g480_p_spl_,
    g480_p
  );


  buf

  (
    g480_p_spl_0,
    g480_p_spl_
  );


  buf

  (
    g473_p_spl_,
    g473_p
  );


  buf

  (
    g444_p_spl_,
    g444_p
  );


  buf

  (
    g444_p_spl_0,
    g444_p_spl_
  );


  buf

  (
    g488_n_spl_,
    g488_n
  );


  buf

  (
    g485_p_spl_,
    g485_p
  );


  buf

  (
    g488_p_spl_,
    g488_p
  );


  buf

  (
    g485_n_spl_,
    g485_n
  );


  buf

  (
    G132_n_spl_,
    G132_n
  );


  buf

  (
    G132_n_spl_0,
    G132_n_spl_
  );


  buf

  (
    G132_p_spl_,
    G132_p
  );


  buf

  (
    G132_p_spl_0,
    G132_p_spl_
  );


  buf

  (
    g494_n_spl_,
    g494_n
  );


  buf

  (
    g494_p_spl_,
    g494_p
  );


  buf

  (
    g500_n_spl_,
    g500_n
  );


  buf

  (
    g497_n_spl_,
    g497_n
  );


  buf

  (
    g500_p_spl_,
    g500_p
  );


  buf

  (
    g497_p_spl_,
    g497_p
  );


  buf

  (
    g512_n_spl_,
    g512_n
  );


  buf

  (
    g509_p_spl_,
    g509_p
  );


  buf

  (
    g512_p_spl_,
    g512_p
  );


  buf

  (
    g509_n_spl_,
    g509_n
  );


  buf

  (
    G111_n_spl_,
    G111_n
  );


  buf

  (
    G111_n_spl_0,
    G111_n_spl_
  );


  buf

  (
    G111_p_spl_,
    G111_p
  );


  buf

  (
    G111_p_spl_0,
    G111_p_spl_
  );


  buf

  (
    g521_n_spl_,
    g521_n
  );


  buf

  (
    g518_n_spl_,
    g518_n
  );


  buf

  (
    g521_p_spl_,
    g521_p
  );


  buf

  (
    g518_p_spl_,
    g518_p
  );


  buf

  (
    g527_n_spl_,
    g527_n
  );


  buf

  (
    g524_n_spl_,
    g524_n
  );


  buf

  (
    g527_p_spl_,
    g527_p
  );


  buf

  (
    g524_p_spl_,
    g524_p
  );


  buf

  (
    g535_n_spl_,
    g535_n
  );


  buf

  (
    g535_n_spl_0,
    g535_n_spl_
  );


  buf

  (
    g535_n_spl_1,
    g535_n_spl_
  );


  buf

  (
    g535_p_spl_,
    g535_p
  );


  buf

  (
    g535_p_spl_0,
    g535_p_spl_
  );


  buf

  (
    g535_p_spl_1,
    g535_p_spl_
  );


  buf

  (
    g537_n_spl_,
    g537_n
  );


  buf

  (
    g537_n_spl_0,
    g537_n_spl_
  );


  buf

  (
    g537_n_spl_00,
    g537_n_spl_0
  );


  buf

  (
    g537_n_spl_1,
    g537_n_spl_
  );


  buf

  (
    g537_p_spl_,
    g537_p
  );


  buf

  (
    g537_p_spl_0,
    g537_p_spl_
  );


  buf

  (
    g537_p_spl_00,
    g537_p_spl_0
  );


  buf

  (
    g537_p_spl_1,
    g537_p_spl_
  );


  buf

  (
    g539_n_spl_,
    g539_n
  );


  buf

  (
    g539_n_spl_0,
    g539_n_spl_
  );


  buf

  (
    g539_n_spl_1,
    g539_n_spl_
  );


  buf

  (
    g539_p_spl_,
    g539_p
  );


  buf

  (
    g539_p_spl_0,
    g539_p_spl_
  );


  buf

  (
    g539_p_spl_1,
    g539_p_spl_
  );


  buf

  (
    g541_p_spl_,
    g541_p
  );


  buf

  (
    g541_p_spl_0,
    g541_p_spl_
  );


  buf

  (
    g541_p_spl_00,
    g541_p_spl_0
  );


  buf

  (
    g541_p_spl_1,
    g541_p_spl_
  );


  buf

  (
    g544_n_spl_,
    g544_n
  );


  buf

  (
    g544_n_spl_0,
    g544_n_spl_
  );


  buf

  (
    g544_n_spl_1,
    g544_n_spl_
  );


  buf

  (
    g544_p_spl_,
    g544_p
  );


  buf

  (
    g544_p_spl_0,
    g544_p_spl_
  );


  buf

  (
    g544_p_spl_1,
    g544_p_spl_
  );


  buf

  (
    g545_n_spl_,
    g545_n
  );


  buf

  (
    g545_p_spl_,
    g545_p
  );


  buf

  (
    g546_p_spl_,
    g546_p
  );


  buf

  (
    g546_p_spl_0,
    g546_p_spl_
  );


  buf

  (
    g546_p_spl_1,
    g546_p_spl_
  );


  buf

  (
    g553_p_spl_,
    g553_p
  );


  buf

  (
    G177_p_spl_,
    G177_p
  );


  buf

  (
    G177_p_spl_0,
    G177_p_spl_
  );


  buf

  (
    G177_p_spl_00,
    G177_p_spl_0
  );


  buf

  (
    G177_p_spl_000,
    G177_p_spl_00
  );


  buf

  (
    G177_p_spl_0000,
    G177_p_spl_000
  );


  buf

  (
    G177_p_spl_0001,
    G177_p_spl_000
  );


  buf

  (
    G177_p_spl_001,
    G177_p_spl_00
  );


  buf

  (
    G177_p_spl_0010,
    G177_p_spl_001
  );


  buf

  (
    G177_p_spl_0011,
    G177_p_spl_001
  );


  buf

  (
    G177_p_spl_01,
    G177_p_spl_0
  );


  buf

  (
    G177_p_spl_010,
    G177_p_spl_01
  );


  buf

  (
    G177_p_spl_0100,
    G177_p_spl_010
  );


  buf

  (
    G177_p_spl_0101,
    G177_p_spl_010
  );


  buf

  (
    G177_p_spl_011,
    G177_p_spl_01
  );


  buf

  (
    G177_p_spl_0110,
    G177_p_spl_011
  );


  buf

  (
    G177_p_spl_0111,
    G177_p_spl_011
  );


  buf

  (
    G177_p_spl_1,
    G177_p_spl_
  );


  buf

  (
    G177_p_spl_10,
    G177_p_spl_1
  );


  buf

  (
    G177_p_spl_100,
    G177_p_spl_10
  );


  buf

  (
    G177_p_spl_1000,
    G177_p_spl_100
  );


  buf

  (
    G177_p_spl_1001,
    G177_p_spl_100
  );


  buf

  (
    G177_p_spl_101,
    G177_p_spl_10
  );


  buf

  (
    G177_p_spl_11,
    G177_p_spl_1
  );


  buf

  (
    G177_p_spl_110,
    G177_p_spl_11
  );


  buf

  (
    G177_p_spl_111,
    G177_p_spl_11
  );


  buf

  (
    G176_p_spl_,
    G176_p
  );


  buf

  (
    G176_p_spl_0,
    G176_p_spl_
  );


  buf

  (
    G176_p_spl_00,
    G176_p_spl_0
  );


  buf

  (
    G176_p_spl_000,
    G176_p_spl_00
  );


  buf

  (
    G176_p_spl_0000,
    G176_p_spl_000
  );


  buf

  (
    G176_p_spl_00000,
    G176_p_spl_0000
  );


  buf

  (
    G176_p_spl_00001,
    G176_p_spl_0000
  );


  buf

  (
    G176_p_spl_0001,
    G176_p_spl_000
  );


  buf

  (
    G176_p_spl_001,
    G176_p_spl_00
  );


  buf

  (
    G176_p_spl_0010,
    G176_p_spl_001
  );


  buf

  (
    G176_p_spl_0011,
    G176_p_spl_001
  );


  buf

  (
    G176_p_spl_01,
    G176_p_spl_0
  );


  buf

  (
    G176_p_spl_010,
    G176_p_spl_01
  );


  buf

  (
    G176_p_spl_0100,
    G176_p_spl_010
  );


  buf

  (
    G176_p_spl_0101,
    G176_p_spl_010
  );


  buf

  (
    G176_p_spl_011,
    G176_p_spl_01
  );


  buf

  (
    G176_p_spl_0110,
    G176_p_spl_011
  );


  buf

  (
    G176_p_spl_0111,
    G176_p_spl_011
  );


  buf

  (
    G176_p_spl_1,
    G176_p_spl_
  );


  buf

  (
    G176_p_spl_10,
    G176_p_spl_1
  );


  buf

  (
    G176_p_spl_100,
    G176_p_spl_10
  );


  buf

  (
    G176_p_spl_1000,
    G176_p_spl_100
  );


  buf

  (
    G176_p_spl_1001,
    G176_p_spl_100
  );


  buf

  (
    G176_p_spl_101,
    G176_p_spl_10
  );


  buf

  (
    G176_p_spl_1010,
    G176_p_spl_101
  );


  buf

  (
    G176_p_spl_1011,
    G176_p_spl_101
  );


  buf

  (
    G176_p_spl_11,
    G176_p_spl_1
  );


  buf

  (
    G176_p_spl_110,
    G176_p_spl_11
  );


  buf

  (
    G176_p_spl_1100,
    G176_p_spl_110
  );


  buf

  (
    G176_p_spl_1101,
    G176_p_spl_110
  );


  buf

  (
    G176_p_spl_111,
    G176_p_spl_11
  );


  buf

  (
    G176_p_spl_1110,
    G176_p_spl_111
  );


  buf

  (
    G176_p_spl_1111,
    G176_p_spl_111
  );


  buf

  (
    G177_n_spl_,
    G177_n
  );


  buf

  (
    G177_n_spl_0,
    G177_n_spl_
  );


  buf

  (
    G177_n_spl_00,
    G177_n_spl_0
  );


  buf

  (
    G177_n_spl_000,
    G177_n_spl_00
  );


  buf

  (
    G177_n_spl_0000,
    G177_n_spl_000
  );


  buf

  (
    G177_n_spl_0001,
    G177_n_spl_000
  );


  buf

  (
    G177_n_spl_001,
    G177_n_spl_00
  );


  buf

  (
    G177_n_spl_0010,
    G177_n_spl_001
  );


  buf

  (
    G177_n_spl_0011,
    G177_n_spl_001
  );


  buf

  (
    G177_n_spl_01,
    G177_n_spl_0
  );


  buf

  (
    G177_n_spl_010,
    G177_n_spl_01
  );


  buf

  (
    G177_n_spl_011,
    G177_n_spl_01
  );


  buf

  (
    G177_n_spl_1,
    G177_n_spl_
  );


  buf

  (
    G177_n_spl_10,
    G177_n_spl_1
  );


  buf

  (
    G177_n_spl_100,
    G177_n_spl_10
  );


  buf

  (
    G177_n_spl_101,
    G177_n_spl_10
  );


  buf

  (
    G177_n_spl_11,
    G177_n_spl_1
  );


  buf

  (
    G177_n_spl_110,
    G177_n_spl_11
  );


  buf

  (
    G177_n_spl_111,
    G177_n_spl_11
  );


  buf

  (
    G176_n_spl_,
    G176_n
  );


  buf

  (
    G176_n_spl_0,
    G176_n_spl_
  );


  buf

  (
    G176_n_spl_00,
    G176_n_spl_0
  );


  buf

  (
    G176_n_spl_000,
    G176_n_spl_00
  );


  buf

  (
    G176_n_spl_0000,
    G176_n_spl_000
  );


  buf

  (
    G176_n_spl_0001,
    G176_n_spl_000
  );


  buf

  (
    G176_n_spl_001,
    G176_n_spl_00
  );


  buf

  (
    G176_n_spl_0010,
    G176_n_spl_001
  );


  buf

  (
    G176_n_spl_0011,
    G176_n_spl_001
  );


  buf

  (
    G176_n_spl_01,
    G176_n_spl_0
  );


  buf

  (
    G176_n_spl_010,
    G176_n_spl_01
  );


  buf

  (
    G176_n_spl_0100,
    G176_n_spl_010
  );


  buf

  (
    G176_n_spl_0101,
    G176_n_spl_010
  );


  buf

  (
    G176_n_spl_011,
    G176_n_spl_01
  );


  buf

  (
    G176_n_spl_1,
    G176_n_spl_
  );


  buf

  (
    G176_n_spl_10,
    G176_n_spl_1
  );


  buf

  (
    G176_n_spl_100,
    G176_n_spl_10
  );


  buf

  (
    G176_n_spl_101,
    G176_n_spl_10
  );


  buf

  (
    G176_n_spl_11,
    G176_n_spl_1
  );


  buf

  (
    G176_n_spl_110,
    G176_n_spl_11
  );


  buf

  (
    G176_n_spl_111,
    G176_n_spl_11
  );


  buf

  (
    g562_n_spl_,
    g562_n
  );


  buf

  (
    g562_n_spl_0,
    g562_n_spl_
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G2_p_spl_0,
    G2_p_spl_
  );


  buf

  (
    G2_p_spl_1,
    G2_p_spl_
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G2_n_spl_0,
    G2_n_spl_
  );


  buf

  (
    g570_n_spl_,
    g570_n
  );


  buf

  (
    g572_p_spl_,
    g572_p
  );


  buf

  (
    G173_n_spl_,
    G173_n
  );


  buf

  (
    G173_n_spl_0,
    G173_n_spl_
  );


  buf

  (
    G173_n_spl_00,
    G173_n_spl_0
  );


  buf

  (
    G173_n_spl_000,
    G173_n_spl_00
  );


  buf

  (
    G173_n_spl_0000,
    G173_n_spl_000
  );


  buf

  (
    G173_n_spl_0001,
    G173_n_spl_000
  );


  buf

  (
    G173_n_spl_001,
    G173_n_spl_00
  );


  buf

  (
    G173_n_spl_0010,
    G173_n_spl_001
  );


  buf

  (
    G173_n_spl_0011,
    G173_n_spl_001
  );


  buf

  (
    G173_n_spl_01,
    G173_n_spl_0
  );


  buf

  (
    G173_n_spl_010,
    G173_n_spl_01
  );


  buf

  (
    G173_n_spl_011,
    G173_n_spl_01
  );


  buf

  (
    G173_n_spl_1,
    G173_n_spl_
  );


  buf

  (
    G173_n_spl_10,
    G173_n_spl_1
  );


  buf

  (
    G173_n_spl_100,
    G173_n_spl_10
  );


  buf

  (
    G173_n_spl_101,
    G173_n_spl_10
  );


  buf

  (
    G173_n_spl_11,
    G173_n_spl_1
  );


  buf

  (
    G173_n_spl_110,
    G173_n_spl_11
  );


  buf

  (
    G173_n_spl_111,
    G173_n_spl_11
  );


  buf

  (
    G22_p_spl_,
    G22_p
  );


  buf

  (
    G173_p_spl_,
    G173_p
  );


  buf

  (
    G173_p_spl_0,
    G173_p_spl_
  );


  buf

  (
    G173_p_spl_00,
    G173_p_spl_0
  );


  buf

  (
    G173_p_spl_000,
    G173_p_spl_00
  );


  buf

  (
    G173_p_spl_0000,
    G173_p_spl_000
  );


  buf

  (
    G173_p_spl_0001,
    G173_p_spl_000
  );


  buf

  (
    G173_p_spl_001,
    G173_p_spl_00
  );


  buf

  (
    G173_p_spl_0010,
    G173_p_spl_001
  );


  buf

  (
    G173_p_spl_0011,
    G173_p_spl_001
  );


  buf

  (
    G173_p_spl_01,
    G173_p_spl_0
  );


  buf

  (
    G173_p_spl_010,
    G173_p_spl_01
  );


  buf

  (
    G173_p_spl_011,
    G173_p_spl_01
  );


  buf

  (
    G173_p_spl_1,
    G173_p_spl_
  );


  buf

  (
    G173_p_spl_10,
    G173_p_spl_1
  );


  buf

  (
    G173_p_spl_100,
    G173_p_spl_10
  );


  buf

  (
    G173_p_spl_101,
    G173_p_spl_10
  );


  buf

  (
    G173_p_spl_11,
    G173_p_spl_1
  );


  buf

  (
    G173_p_spl_110,
    G173_p_spl_11
  );


  buf

  (
    G173_p_spl_111,
    G173_p_spl_11
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G172_n_spl_,
    G172_n
  );


  buf

  (
    G172_n_spl_0,
    G172_n_spl_
  );


  buf

  (
    G172_n_spl_00,
    G172_n_spl_0
  );


  buf

  (
    G172_n_spl_000,
    G172_n_spl_00
  );


  buf

  (
    G172_n_spl_001,
    G172_n_spl_00
  );


  buf

  (
    G172_n_spl_01,
    G172_n_spl_0
  );


  buf

  (
    G172_n_spl_1,
    G172_n_spl_
  );


  buf

  (
    G172_n_spl_10,
    G172_n_spl_1
  );


  buf

  (
    G172_n_spl_11,
    G172_n_spl_1
  );


  buf

  (
    g579_p_spl_,
    g579_p
  );


  buf

  (
    g579_p_spl_0,
    g579_p_spl_
  );


  buf

  (
    g579_p_spl_00,
    g579_p_spl_0
  );


  buf

  (
    g579_p_spl_1,
    g579_p_spl_
  );


  buf

  (
    g560_p_spl_,
    g560_p
  );


  buf

  (
    g560_p_spl_0,
    g560_p_spl_
  );


  buf

  (
    g560_p_spl_00,
    g560_p_spl_0
  );


  buf

  (
    g560_p_spl_1,
    g560_p_spl_
  );


  buf

  (
    G172_p_spl_,
    G172_p
  );


  buf

  (
    G172_p_spl_0,
    G172_p_spl_
  );


  buf

  (
    G172_p_spl_00,
    G172_p_spl_0
  );


  buf

  (
    G172_p_spl_000,
    G172_p_spl_00
  );


  buf

  (
    G172_p_spl_001,
    G172_p_spl_00
  );


  buf

  (
    G172_p_spl_01,
    G172_p_spl_0
  );


  buf

  (
    G172_p_spl_1,
    G172_p_spl_
  );


  buf

  (
    G172_p_spl_10,
    G172_p_spl_1
  );


  buf

  (
    G172_p_spl_11,
    G172_p_spl_1
  );


  buf

  (
    g594_n_spl_,
    g594_n
  );


  buf

  (
    g594_p_spl_,
    g594_p
  );


  buf

  (
    g595_n_spl_,
    g595_n
  );


  buf

  (
    g596_n_spl_,
    g596_n
  );


  buf

  (
    g596_n_spl_0,
    g596_n_spl_
  );


  buf

  (
    g596_p_spl_,
    g596_p
  );


  buf

  (
    g596_p_spl_0,
    g596_p_spl_
  );


  buf

  (
    g596_p_spl_1,
    g596_p_spl_
  );


  buf

  (
    g597_p_spl_,
    g597_p
  );


  buf

  (
    g598_p_spl_,
    g598_p
  );


  buf

  (
    g598_p_spl_0,
    g598_p_spl_
  );


  buf

  (
    g598_n_spl_,
    g598_n
  );


  buf

  (
    g598_n_spl_0,
    g598_n_spl_
  );


  buf

  (
    g601_p_spl_,
    g601_p
  );


  buf

  (
    g610_n_spl_,
    g610_n
  );


  buf

  (
    g617_p_spl_,
    g617_p
  );


  buf

  (
    g617_p_spl_0,
    g617_p_spl_
  );


  buf

  (
    g619_n_spl_,
    g619_n
  );


  buf

  (
    G174_n_spl_,
    G174_n
  );


  buf

  (
    G174_n_spl_0,
    G174_n_spl_
  );


  buf

  (
    G174_n_spl_00,
    G174_n_spl_0
  );


  buf

  (
    G174_n_spl_000,
    G174_n_spl_00
  );


  buf

  (
    G174_n_spl_0000,
    G174_n_spl_000
  );


  buf

  (
    G174_n_spl_0001,
    G174_n_spl_000
  );


  buf

  (
    G174_n_spl_001,
    G174_n_spl_00
  );


  buf

  (
    G174_n_spl_0010,
    G174_n_spl_001
  );


  buf

  (
    G174_n_spl_0011,
    G174_n_spl_001
  );


  buf

  (
    G174_n_spl_01,
    G174_n_spl_0
  );


  buf

  (
    G174_n_spl_010,
    G174_n_spl_01
  );


  buf

  (
    G174_n_spl_011,
    G174_n_spl_01
  );


  buf

  (
    G174_n_spl_1,
    G174_n_spl_
  );


  buf

  (
    G174_n_spl_10,
    G174_n_spl_1
  );


  buf

  (
    G174_n_spl_100,
    G174_n_spl_10
  );


  buf

  (
    G174_n_spl_101,
    G174_n_spl_10
  );


  buf

  (
    G174_n_spl_11,
    G174_n_spl_1
  );


  buf

  (
    G174_n_spl_110,
    G174_n_spl_11
  );


  buf

  (
    G174_n_spl_111,
    G174_n_spl_11
  );


  buf

  (
    G174_p_spl_,
    G174_p
  );


  buf

  (
    G174_p_spl_0,
    G174_p_spl_
  );


  buf

  (
    G174_p_spl_00,
    G174_p_spl_0
  );


  buf

  (
    G174_p_spl_000,
    G174_p_spl_00
  );


  buf

  (
    G174_p_spl_0000,
    G174_p_spl_000
  );


  buf

  (
    G174_p_spl_0001,
    G174_p_spl_000
  );


  buf

  (
    G174_p_spl_001,
    G174_p_spl_00
  );


  buf

  (
    G174_p_spl_0010,
    G174_p_spl_001
  );


  buf

  (
    G174_p_spl_0011,
    G174_p_spl_001
  );


  buf

  (
    G174_p_spl_01,
    G174_p_spl_0
  );


  buf

  (
    G174_p_spl_010,
    G174_p_spl_01
  );


  buf

  (
    G174_p_spl_011,
    G174_p_spl_01
  );


  buf

  (
    G174_p_spl_1,
    G174_p_spl_
  );


  buf

  (
    G174_p_spl_10,
    G174_p_spl_1
  );


  buf

  (
    G174_p_spl_100,
    G174_p_spl_10
  );


  buf

  (
    G174_p_spl_101,
    G174_p_spl_10
  );


  buf

  (
    G174_p_spl_11,
    G174_p_spl_1
  );


  buf

  (
    G174_p_spl_110,
    G174_p_spl_11
  );


  buf

  (
    G174_p_spl_111,
    G174_p_spl_11
  );


  buf

  (
    G175_n_spl_,
    G175_n
  );


  buf

  (
    G175_n_spl_0,
    G175_n_spl_
  );


  buf

  (
    G175_n_spl_00,
    G175_n_spl_0
  );


  buf

  (
    G175_n_spl_000,
    G175_n_spl_00
  );


  buf

  (
    G175_n_spl_001,
    G175_n_spl_00
  );


  buf

  (
    G175_n_spl_01,
    G175_n_spl_0
  );


  buf

  (
    G175_n_spl_1,
    G175_n_spl_
  );


  buf

  (
    G175_n_spl_10,
    G175_n_spl_1
  );


  buf

  (
    G175_n_spl_11,
    G175_n_spl_1
  );


  buf

  (
    G175_p_spl_,
    G175_p
  );


  buf

  (
    G175_p_spl_0,
    G175_p_spl_
  );


  buf

  (
    G175_p_spl_00,
    G175_p_spl_0
  );


  buf

  (
    G175_p_spl_000,
    G175_p_spl_00
  );


  buf

  (
    G175_p_spl_001,
    G175_p_spl_00
  );


  buf

  (
    G175_p_spl_01,
    G175_p_spl_0
  );


  buf

  (
    G175_p_spl_1,
    G175_p_spl_
  );


  buf

  (
    G175_p_spl_10,
    G175_p_spl_1
  );


  buf

  (
    G175_p_spl_11,
    G175_p_spl_1
  );


  buf

  (
    g638_p_spl_,
    g638_p
  );


  buf

  (
    g639_p_spl_,
    g639_p
  );


  buf

  (
    g643_n_spl_,
    g643_n
  );


  buf

  (
    g652_n_spl_,
    g652_n
  );


  buf

  (
    g659_p_spl_,
    g659_p
  );


  buf

  (
    g660_p_spl_,
    g660_p
  );


  buf

  (
    g664_n_spl_,
    g664_n
  );


  buf

  (
    g673_n_spl_,
    g673_n
  );


  buf

  (
    g681_p_spl_,
    g681_p
  );


  buf

  (
    g581_n_spl_,
    g581_n
  );


  buf

  (
    g581_n_spl_0,
    g581_n_spl_
  );


  buf

  (
    g581_n_spl_00,
    g581_n_spl_0
  );


  buf

  (
    g581_n_spl_01,
    g581_n_spl_0
  );


  buf

  (
    g581_n_spl_1,
    g581_n_spl_
  );


  buf

  (
    g581_n_spl_10,
    g581_n_spl_1
  );


  buf

  (
    g581_n_spl_11,
    g581_n_spl_1
  );


  buf

  (
    g681_n_spl_,
    g681_n
  );


  buf

  (
    g581_p_spl_,
    g581_p
  );


  buf

  (
    g581_p_spl_0,
    g581_p_spl_
  );


  buf

  (
    g581_p_spl_00,
    g581_p_spl_0
  );


  buf

  (
    g581_p_spl_01,
    g581_p_spl_0
  );


  buf

  (
    g581_p_spl_1,
    g581_p_spl_
  );


  buf

  (
    g687_n_spl_,
    g687_n
  );


  buf

  (
    g687_p_spl_,
    g687_p
  );


  buf

  (
    g696_n_spl_,
    g696_n
  );


  buf

  (
    g693_n_spl_,
    g693_n
  );


  buf

  (
    g696_p_spl_,
    g696_p
  );


  buf

  (
    g693_p_spl_,
    g693_p
  );


  buf

  (
    g699_n_spl_,
    g699_n
  );


  buf

  (
    g690_p_spl_,
    g690_p
  );


  buf

  (
    g699_p_spl_,
    g699_p
  );


  buf

  (
    g690_n_spl_,
    g690_n
  );


  buf

  (
    g711_n_spl_,
    g711_n
  );


  buf

  (
    g708_p_spl_,
    g708_p
  );


  buf

  (
    g711_p_spl_,
    g711_p
  );


  buf

  (
    g708_n_spl_,
    g708_n
  );


  buf

  (
    g717_n_spl_,
    g717_n
  );


  buf

  (
    g717_p_spl_,
    g717_p
  );


  buf

  (
    g723_n_spl_,
    g723_n
  );


  buf

  (
    g720_p_spl_,
    g720_p
  );


  buf

  (
    g723_p_spl_,
    g723_p
  );


  buf

  (
    g720_n_spl_,
    g720_n
  );


  buf

  (
    g729_n_spl_,
    g729_n
  );


  buf

  (
    g726_n_spl_,
    g726_n
  );


  buf

  (
    g729_p_spl_,
    g729_p
  );


  buf

  (
    g726_p_spl_,
    g726_p
  );


  buf

  (
    g430_p_spl_,
    g430_p
  );


  buf

  (
    g430_p_spl_0,
    g430_p_spl_
  );


  buf

  (
    g541_n_spl_,
    g541_n
  );


  buf

  (
    g541_n_spl_0,
    g541_n_spl_
  );


  buf

  (
    g541_n_spl_1,
    g541_n_spl_
  );


  buf

  (
    g737_p_spl_,
    g737_p
  );


  buf

  (
    g737_p_spl_0,
    g737_p_spl_
  );


  buf

  (
    g737_p_spl_00,
    g737_p_spl_0
  );


  buf

  (
    g737_p_spl_1,
    g737_p_spl_
  );


  buf

  (
    g737_n_spl_,
    g737_n
  );


  buf

  (
    g737_n_spl_0,
    g737_n_spl_
  );


  buf

  (
    g737_n_spl_00,
    g737_n_spl_0
  );


  buf

  (
    g737_n_spl_1,
    g737_n_spl_
  );


  buf

  (
    g743_p_spl_,
    g743_p
  );


  buf

  (
    g747_p_spl_,
    g747_p
  );


  buf

  (
    g389_p_spl_,
    g389_p
  );


  buf

  (
    g546_n_spl_,
    g546_n
  );


  buf

  (
    g546_n_spl_0,
    g546_n_spl_
  );


  buf

  (
    g395_p_spl_,
    g395_p
  );


  buf

  (
    g395_p_spl_0,
    g395_p_spl_
  );


  buf

  (
    g395_p_spl_00,
    g395_p_spl_0
  );


  buf

  (
    g395_p_spl_1,
    g395_p_spl_
  );


  buf

  (
    g760_p_spl_,
    g760_p
  );


  buf

  (
    g755_p_spl_,
    g755_p
  );


  buf

  (
    g774_p_spl_,
    g774_p
  );


  buf

  (
    g774_p_spl_0,
    g774_p_spl_
  );


  buf

  (
    g774_p_spl_00,
    g774_p_spl_0
  );


  buf

  (
    g774_p_spl_01,
    g774_p_spl_0
  );


  buf

  (
    g774_p_spl_1,
    g774_p_spl_
  );


  buf

  (
    g774_n_spl_,
    g774_n
  );


  buf

  (
    g774_n_spl_0,
    g774_n_spl_
  );


  buf

  (
    g774_n_spl_00,
    g774_n_spl_0
  );


  buf

  (
    g774_n_spl_01,
    g774_n_spl_0
  );


  buf

  (
    g774_n_spl_1,
    g774_n_spl_
  );


  buf

  (
    g777_p_spl_,
    g777_p
  );


  buf

  (
    g444_n_spl_,
    g444_n
  );


  buf

  (
    g780_p_spl_,
    g780_p
  );


  buf

  (
    g780_p_spl_0,
    g780_p_spl_
  );


  buf

  (
    g780_p_spl_1,
    g780_p_spl_
  );


  buf

  (
    g780_n_spl_,
    g780_n
  );


  buf

  (
    g780_n_spl_0,
    g780_n_spl_
  );


  buf

  (
    g780_n_spl_1,
    g780_n_spl_
  );


  buf

  (
    g791_p_spl_,
    g791_p
  );


  buf

  (
    g785_p_spl_,
    g785_p
  );


  buf

  (
    G158_n_spl_,
    G158_n
  );


  buf

  (
    G158_n_spl_0,
    G158_n_spl_
  );


  buf

  (
    G158_n_spl_00,
    G158_n_spl_0
  );


  buf

  (
    G158_n_spl_000,
    G158_n_spl_00
  );


  buf

  (
    G158_n_spl_0000,
    G158_n_spl_000
  );


  buf

  (
    G158_n_spl_0001,
    G158_n_spl_000
  );


  buf

  (
    G158_n_spl_001,
    G158_n_spl_00
  );


  buf

  (
    G158_n_spl_0010,
    G158_n_spl_001
  );


  buf

  (
    G158_n_spl_0011,
    G158_n_spl_001
  );


  buf

  (
    G158_n_spl_01,
    G158_n_spl_0
  );


  buf

  (
    G158_n_spl_010,
    G158_n_spl_01
  );


  buf

  (
    G158_n_spl_011,
    G158_n_spl_01
  );


  buf

  (
    G158_n_spl_1,
    G158_n_spl_
  );


  buf

  (
    G158_n_spl_10,
    G158_n_spl_1
  );


  buf

  (
    G158_n_spl_100,
    G158_n_spl_10
  );


  buf

  (
    G158_n_spl_101,
    G158_n_spl_10
  );


  buf

  (
    G158_n_spl_11,
    G158_n_spl_1
  );


  buf

  (
    G158_n_spl_110,
    G158_n_spl_11
  );


  buf

  (
    G158_n_spl_111,
    G158_n_spl_11
  );


  buf

  (
    G81_p_spl_,
    G81_p
  );


  buf

  (
    G158_p_spl_,
    G158_p
  );


  buf

  (
    G158_p_spl_0,
    G158_p_spl_
  );


  buf

  (
    G158_p_spl_00,
    G158_p_spl_0
  );


  buf

  (
    G158_p_spl_000,
    G158_p_spl_00
  );


  buf

  (
    G158_p_spl_0000,
    G158_p_spl_000
  );


  buf

  (
    G158_p_spl_0001,
    G158_p_spl_000
  );


  buf

  (
    G158_p_spl_001,
    G158_p_spl_00
  );


  buf

  (
    G158_p_spl_0010,
    G158_p_spl_001
  );


  buf

  (
    G158_p_spl_0011,
    G158_p_spl_001
  );


  buf

  (
    G158_p_spl_01,
    G158_p_spl_0
  );


  buf

  (
    G158_p_spl_010,
    G158_p_spl_01
  );


  buf

  (
    G158_p_spl_011,
    G158_p_spl_01
  );


  buf

  (
    G158_p_spl_1,
    G158_p_spl_
  );


  buf

  (
    G158_p_spl_10,
    G158_p_spl_1
  );


  buf

  (
    G158_p_spl_100,
    G158_p_spl_10
  );


  buf

  (
    G158_p_spl_101,
    G158_p_spl_10
  );


  buf

  (
    G158_p_spl_11,
    G158_p_spl_1
  );


  buf

  (
    G158_p_spl_110,
    G158_p_spl_11
  );


  buf

  (
    G158_p_spl_111,
    G158_p_spl_11
  );


  buf

  (
    G80_p_spl_,
    G80_p
  );


  buf

  (
    G159_n_spl_,
    G159_n
  );


  buf

  (
    G159_n_spl_0,
    G159_n_spl_
  );


  buf

  (
    G159_n_spl_00,
    G159_n_spl_0
  );


  buf

  (
    G159_n_spl_000,
    G159_n_spl_00
  );


  buf

  (
    G159_n_spl_001,
    G159_n_spl_00
  );


  buf

  (
    G159_n_spl_01,
    G159_n_spl_0
  );


  buf

  (
    G159_n_spl_1,
    G159_n_spl_
  );


  buf

  (
    G159_n_spl_10,
    G159_n_spl_1
  );


  buf

  (
    G159_n_spl_11,
    G159_n_spl_1
  );


  buf

  (
    G159_p_spl_,
    G159_p
  );


  buf

  (
    G159_p_spl_0,
    G159_p_spl_
  );


  buf

  (
    G159_p_spl_00,
    G159_p_spl_0
  );


  buf

  (
    G159_p_spl_000,
    G159_p_spl_00
  );


  buf

  (
    G159_p_spl_001,
    G159_p_spl_00
  );


  buf

  (
    G159_p_spl_01,
    G159_p_spl_0
  );


  buf

  (
    G159_p_spl_1,
    G159_p_spl_
  );


  buf

  (
    G159_p_spl_10,
    G159_p_spl_1
  );


  buf

  (
    G159_p_spl_11,
    G159_p_spl_1
  );


  buf

  (
    G64_p_spl_,
    G64_p
  );


  buf

  (
    G64_p_spl_0,
    G64_p_spl_
  );


  buf

  (
    G64_p_spl_00,
    G64_p_spl_0
  );


  buf

  (
    G64_p_spl_000,
    G64_p_spl_00
  );


  buf

  (
    G64_p_spl_0000,
    G64_p_spl_000
  );


  buf

  (
    G64_p_spl_0001,
    G64_p_spl_000
  );


  buf

  (
    G64_p_spl_001,
    G64_p_spl_00
  );


  buf

  (
    G64_p_spl_0010,
    G64_p_spl_001
  );


  buf

  (
    G64_p_spl_01,
    G64_p_spl_0
  );


  buf

  (
    G64_p_spl_010,
    G64_p_spl_01
  );


  buf

  (
    G64_p_spl_011,
    G64_p_spl_01
  );


  buf

  (
    G64_p_spl_1,
    G64_p_spl_
  );


  buf

  (
    G64_p_spl_10,
    G64_p_spl_1
  );


  buf

  (
    G64_p_spl_100,
    G64_p_spl_10
  );


  buf

  (
    G64_p_spl_101,
    G64_p_spl_10
  );


  buf

  (
    G64_p_spl_11,
    G64_p_spl_1
  );


  buf

  (
    G64_p_spl_110,
    G64_p_spl_11
  );


  buf

  (
    G64_p_spl_111,
    G64_p_spl_11
  );


  buf

  (
    G160_n_spl_,
    G160_n
  );


  buf

  (
    G160_n_spl_0,
    G160_n_spl_
  );


  buf

  (
    G160_n_spl_00,
    G160_n_spl_0
  );


  buf

  (
    G160_n_spl_000,
    G160_n_spl_00
  );


  buf

  (
    G160_n_spl_0000,
    G160_n_spl_000
  );


  buf

  (
    G160_n_spl_0001,
    G160_n_spl_000
  );


  buf

  (
    G160_n_spl_001,
    G160_n_spl_00
  );


  buf

  (
    G160_n_spl_0010,
    G160_n_spl_001
  );


  buf

  (
    G160_n_spl_0011,
    G160_n_spl_001
  );


  buf

  (
    G160_n_spl_01,
    G160_n_spl_0
  );


  buf

  (
    G160_n_spl_010,
    G160_n_spl_01
  );


  buf

  (
    G160_n_spl_011,
    G160_n_spl_01
  );


  buf

  (
    G160_n_spl_1,
    G160_n_spl_
  );


  buf

  (
    G160_n_spl_10,
    G160_n_spl_1
  );


  buf

  (
    G160_n_spl_100,
    G160_n_spl_10
  );


  buf

  (
    G160_n_spl_101,
    G160_n_spl_10
  );


  buf

  (
    G160_n_spl_11,
    G160_n_spl_1
  );


  buf

  (
    G160_n_spl_110,
    G160_n_spl_11
  );


  buf

  (
    G160_n_spl_111,
    G160_n_spl_11
  );


  buf

  (
    G160_p_spl_,
    G160_p
  );


  buf

  (
    G160_p_spl_0,
    G160_p_spl_
  );


  buf

  (
    G160_p_spl_00,
    G160_p_spl_0
  );


  buf

  (
    G160_p_spl_000,
    G160_p_spl_00
  );


  buf

  (
    G160_p_spl_0000,
    G160_p_spl_000
  );


  buf

  (
    G160_p_spl_0001,
    G160_p_spl_000
  );


  buf

  (
    G160_p_spl_001,
    G160_p_spl_00
  );


  buf

  (
    G160_p_spl_0010,
    G160_p_spl_001
  );


  buf

  (
    G160_p_spl_0011,
    G160_p_spl_001
  );


  buf

  (
    G160_p_spl_01,
    G160_p_spl_0
  );


  buf

  (
    G160_p_spl_010,
    G160_p_spl_01
  );


  buf

  (
    G160_p_spl_011,
    G160_p_spl_01
  );


  buf

  (
    G160_p_spl_1,
    G160_p_spl_
  );


  buf

  (
    G160_p_spl_10,
    G160_p_spl_1
  );


  buf

  (
    G160_p_spl_100,
    G160_p_spl_10
  );


  buf

  (
    G160_p_spl_101,
    G160_p_spl_10
  );


  buf

  (
    G160_p_spl_11,
    G160_p_spl_1
  );


  buf

  (
    G160_p_spl_110,
    G160_p_spl_11
  );


  buf

  (
    G160_p_spl_111,
    G160_p_spl_11
  );


  buf

  (
    G161_n_spl_,
    G161_n
  );


  buf

  (
    G161_n_spl_0,
    G161_n_spl_
  );


  buf

  (
    G161_n_spl_00,
    G161_n_spl_0
  );


  buf

  (
    G161_n_spl_000,
    G161_n_spl_00
  );


  buf

  (
    G161_n_spl_001,
    G161_n_spl_00
  );


  buf

  (
    G161_n_spl_01,
    G161_n_spl_0
  );


  buf

  (
    G161_n_spl_1,
    G161_n_spl_
  );


  buf

  (
    G161_n_spl_10,
    G161_n_spl_1
  );


  buf

  (
    G161_n_spl_11,
    G161_n_spl_1
  );


  buf

  (
    G161_p_spl_,
    G161_p
  );


  buf

  (
    G161_p_spl_0,
    G161_p_spl_
  );


  buf

  (
    G161_p_spl_00,
    G161_p_spl_0
  );


  buf

  (
    G161_p_spl_000,
    G161_p_spl_00
  );


  buf

  (
    G161_p_spl_001,
    G161_p_spl_00
  );


  buf

  (
    G161_p_spl_01,
    G161_p_spl_0
  );


  buf

  (
    G161_p_spl_1,
    G161_p_spl_
  );


  buf

  (
    G161_p_spl_10,
    G161_p_spl_1
  );


  buf

  (
    G161_p_spl_11,
    G161_p_spl_1
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    g647_n_spl_,
    g647_n
  );


  buf

  (
    g647_n_spl_0,
    g647_n_spl_
  );


  buf

  (
    g647_n_spl_00,
    g647_n_spl_0
  );


  buf

  (
    g647_n_spl_1,
    g647_n_spl_
  );


  buf

  (
    g605_n_spl_,
    g605_n
  );


  buf

  (
    g605_n_spl_0,
    g605_n_spl_
  );


  buf

  (
    g605_n_spl_00,
    g605_n_spl_0
  );


  buf

  (
    g605_n_spl_1,
    g605_n_spl_
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G27_p_spl_,
    G27_p
  );


  buf

  (
    g656_n_spl_,
    g656_n
  );


  buf

  (
    g656_n_spl_0,
    g656_n_spl_
  );


  buf

  (
    g656_n_spl_00,
    g656_n_spl_0
  );


  buf

  (
    g656_n_spl_1,
    g656_n_spl_
  );


  buf

  (
    g614_n_spl_,
    g614_n
  );


  buf

  (
    g614_n_spl_0,
    g614_n_spl_
  );


  buf

  (
    g614_n_spl_00,
    g614_n_spl_0
  );


  buf

  (
    g614_n_spl_1,
    g614_n_spl_
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G26_p_spl_,
    G26_p
  );


  buf

  (
    g669_n_spl_,
    g669_n
  );


  buf

  (
    g669_n_spl_0,
    g669_n_spl_
  );


  buf

  (
    g669_n_spl_00,
    g669_n_spl_0
  );


  buf

  (
    g669_n_spl_1,
    g669_n_spl_
  );


  buf

  (
    g624_n_spl_,
    g624_n
  );


  buf

  (
    g624_n_spl_0,
    g624_n_spl_
  );


  buf

  (
    g624_n_spl_00,
    g624_n_spl_0
  );


  buf

  (
    g624_n_spl_1,
    g624_n_spl_
  );


  buf

  (
    G25_p_spl_,
    G25_p
  );


  buf

  (
    G24_p_spl_,
    G24_p
  );


  buf

  (
    g678_n_spl_,
    g678_n
  );


  buf

  (
    g678_n_spl_0,
    g678_n_spl_
  );


  buf

  (
    g678_n_spl_00,
    g678_n_spl_0
  );


  buf

  (
    g678_n_spl_1,
    g678_n_spl_
  );


  buf

  (
    g569_p_spl_,
    g569_p
  );


  buf

  (
    g569_p_spl_0,
    g569_p_spl_
  );


  buf

  (
    g569_p_spl_00,
    g569_p_spl_0
  );


  buf

  (
    g569_p_spl_1,
    g569_p_spl_
  );


  buf

  (
    G76_p_spl_,
    G76_p
  );


  buf

  (
    G86_p_spl_,
    G86_p
  );


  buf

  (
    G72_p_spl_,
    G72_p
  );


  buf

  (
    G82_p_spl_,
    G82_p
  );


  buf

  (
    G70_p_spl_,
    G70_p
  );


  buf

  (
    G71_p_spl_,
    G71_p
  );


  buf

  (
    G68_p_spl_,
    G68_p
  );


  buf

  (
    G69_p_spl_,
    G69_p
  );


  buf

  (
    G171_p_spl_,
    G171_p
  );


  buf

  (
    G171_n_spl_,
    G171_n
  );


  buf

  (
    G54_p_spl_,
    G54_p
  );


  buf

  (
    G61_n_spl_,
    G61_n
  );


  buf

  (
    G61_p_spl_,
    G61_p
  );


  buf

  (
    g975_p_spl_,
    g975_p
  );


  buf

  (
    g533_n_spl_,
    g533_n
  );


  buf

  (
    G99_n_spl_,
    G99_n
  );


  buf

  (
    g735_n_spl_,
    g735_n
  );


  buf

  (
    g184_n_spl_,
    g184_n
  );


  buf

  (
    G155_n_spl_,
    G155_n
  );


  buf

  (
    g179_n_spl_,
    g179_n
  );


  buf

  (
    g705_n_spl_,
    g705_n
  );


  buf

  (
    g506_n_spl_,
    g506_n
  );


  buf

  (
    g1025_n_spl_,
    g1025_n
  );


  buf

  (
    g1025_n_spl_0,
    g1025_n_spl_
  );


  buf

  (
    g1025_n_spl_00,
    g1025_n_spl_0
  );


  buf

  (
    g1025_n_spl_1,
    g1025_n_spl_
  );


  buf

  (
    g990_p_spl_,
    g990_p
  );


  buf

  (
    g990_p_spl_0,
    g990_p_spl_
  );


  buf

  (
    g990_p_spl_00,
    g990_p_spl_0
  );


  buf

  (
    g990_p_spl_1,
    g990_p_spl_
  );


  buf

  (
    G41_p_spl_,
    G41_p
  );


  buf

  (
    G42_p_spl_,
    G42_p
  );


  buf

  (
    G18_p_spl_,
    G18_p
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    g1032_n_spl_,
    g1032_n
  );


  buf

  (
    g1032_n_spl_0,
    g1032_n_spl_
  );


  buf

  (
    g1032_n_spl_00,
    g1032_n_spl_0
  );


  buf

  (
    g1032_n_spl_1,
    g1032_n_spl_
  );


  buf

  (
    g997_n_spl_,
    g997_n
  );


  buf

  (
    g997_n_spl_0,
    g997_n_spl_
  );


  buf

  (
    g997_n_spl_00,
    g997_n_spl_0
  );


  buf

  (
    g997_n_spl_1,
    g997_n_spl_
  );


  buf

  (
    G40_p_spl_,
    G40_p
  );


  buf

  (
    G39_p_spl_,
    G39_p
  );


  buf

  (
    g1039_n_spl_,
    g1039_n
  );


  buf

  (
    g1039_n_spl_0,
    g1039_n_spl_
  );


  buf

  (
    g1039_n_spl_00,
    g1039_n_spl_0
  );


  buf

  (
    g1039_n_spl_1,
    g1039_n_spl_
  );


  buf

  (
    g1004_n_spl_,
    g1004_n
  );


  buf

  (
    g1004_n_spl_0,
    g1004_n_spl_
  );


  buf

  (
    g1004_n_spl_00,
    g1004_n_spl_0
  );


  buf

  (
    g1004_n_spl_1,
    g1004_n_spl_
  );


  buf

  (
    G15_p_spl_,
    G15_p
  );


  buf

  (
    G36_p_spl_,
    G36_p
  );


  buf

  (
    g1046_n_spl_,
    g1046_n
  );


  buf

  (
    g1046_n_spl_0,
    g1046_n_spl_
  );


  buf

  (
    g1046_n_spl_00,
    g1046_n_spl_0
  );


  buf

  (
    g1046_n_spl_1,
    g1046_n_spl_
  );


  buf

  (
    g1011_n_spl_,
    g1011_n
  );


  buf

  (
    g1011_n_spl_0,
    g1011_n_spl_
  );


  buf

  (
    g1011_n_spl_00,
    g1011_n_spl_0
  );


  buf

  (
    g1011_n_spl_1,
    g1011_n_spl_
  );


  buf

  (
    G77_p_spl_,
    G77_p
  );


  buf

  (
    G87_p_spl_,
    G87_p
  );


  buf

  (
    G75_p_spl_,
    G75_p
  );


  buf

  (
    G85_p_spl_,
    G85_p
  );


  buf

  (
    G74_p_spl_,
    G74_p
  );


  buf

  (
    G84_p_spl_,
    G84_p
  );


  buf

  (
    G73_p_spl_,
    G73_p
  );


  buf

  (
    G83_p_spl_,
    G83_p
  );


  buf

  (
    g1202_n_spl_,
    g1202_n
  );


  buf

  (
    g1200_p_spl_,
    g1200_p
  );


  buf

  (
    g1202_p_spl_,
    g1202_p
  );


  buf

  (
    g1200_n_spl_,
    g1200_n
  );


  buf

  (
    g1223_p_spl_,
    g1223_p
  );


  buf

  (
    g1214_n_spl_,
    g1214_n
  );


  buf

  (
    g1223_n_spl_,
    g1223_n
  );


  buf

  (
    g1214_p_spl_,
    g1214_p
  );


  buf

  (
    g1238_p_spl_,
    g1238_p
  );


  buf

  (
    g1229_n_spl_,
    g1229_n
  );


  buf

  (
    g1238_n_spl_,
    g1238_n
  );


  buf

  (
    g1229_p_spl_,
    g1229_p
  );


  buf

  (
    g1241_p_spl_,
    g1241_p
  );


  buf

  (
    g1241_n_spl_,
    g1241_n
  );


  buf

  (
    g245_p_spl_,
    g245_p
  );


  buf

  (
    g1244_n_spl_,
    g1244_n
  );


  buf

  (
    g1226_p_spl_,
    g1226_p
  );


  buf

  (
    g1244_p_spl_,
    g1244_p
  );


  buf

  (
    g1226_n_spl_,
    g1226_n
  );


  buf

  (
    g1254_n_spl_,
    g1254_n
  );


  buf

  (
    g1254_p_spl_,
    g1254_p
  );


  buf

  (
    g617_n_spl_,
    g617_n
  );


  buf

  (
    g1257_p_spl_,
    g1257_p
  );


  buf

  (
    g1257_n_spl_,
    g1257_n
  );


  buf

  (
    G162_n_spl_,
    G162_n
  );


  buf

  (
    G162_p_spl_,
    G162_p
  );


  buf

  (
    g1263_p_spl_,
    g1263_p
  );


  buf

  (
    g1260_p_spl_,
    g1260_p
  );


  buf

  (
    g1263_n_spl_,
    g1263_n
  );


  buf

  (
    g1260_n_spl_,
    g1260_n
  );


  buf

  (
    g1268_n_spl_,
    g1268_n
  );


  buf

  (
    g1268_p_spl_,
    g1268_p
  );


  buf

  (
    g1271_n_spl_,
    g1271_n
  );


  buf

  (
    g1266_n_spl_,
    g1266_n
  );


  buf

  (
    g1271_p_spl_,
    g1271_p
  );


  buf

  (
    g1266_p_spl_,
    g1266_p
  );


  buf

  (
    g1275_n_spl_,
    g1275_n
  );


  buf

  (
    g1275_p_spl_,
    g1275_p
  );


  buf

  (
    g1278_p_spl_,
    g1278_p
  );


  buf

  (
    g1278_n_spl_,
    g1278_n
  );


  buf

  (
    g1281_p_spl_,
    g1281_p
  );


  buf

  (
    g1281_n_spl_,
    g1281_n
  );


  buf

  (
    g1282_n_spl_,
    g1282_n
  );


  buf

  (
    g1282_p_spl_,
    g1282_p
  );


  buf

  (
    g1284_n_spl_,
    g1284_n
  );


  buf

  (
    g1284_p_spl_,
    g1284_p
  );


  buf

  (
    g1288_n_spl_,
    g1288_n
  );


  buf

  (
    g1288_p_spl_,
    g1288_p
  );


  buf

  (
    g1299_p_spl_,
    g1299_p
  );


  buf

  (
    g1299_n_spl_,
    g1299_n
  );


  buf

  (
    g1308_n_spl_,
    g1308_n
  );


  buf

  (
    g1329_p_spl_,
    g1329_p
  );


  buf

  (
    g1320_n_spl_,
    g1320_n
  );


  buf

  (
    g1329_n_spl_,
    g1329_n
  );


  buf

  (
    g1320_p_spl_,
    g1320_p
  );


  buf

  (
    g1341_n_spl_,
    g1341_n
  );


  buf

  (
    g1341_p_spl_,
    g1341_p
  );


  buf

  (
    g317_p_spl_,
    g317_p
  );


  buf

  (
    g1344_p_spl_,
    g1344_p
  );


  buf

  (
    g1332_n_spl_,
    g1332_n
  );


  buf

  (
    g1344_n_spl_,
    g1344_n
  );


  buf

  (
    g1332_p_spl_,
    g1332_p
  );


  buf

  (
    g1365_p_spl_,
    g1365_p
  );


  buf

  (
    g1356_n_spl_,
    g1356_n
  );


  buf

  (
    g1365_n_spl_,
    g1365_n
  );


  buf

  (
    g1356_p_spl_,
    g1356_p
  );


  buf

  (
    g1386_p_spl_,
    g1386_p
  );


  buf

  (
    g1377_n_spl_,
    g1377_n
  );


  buf

  (
    g1386_n_spl_,
    g1386_n
  );


  buf

  (
    g1377_p_spl_,
    g1377_p
  );


  buf

  (
    g1398_n_spl_,
    g1398_n
  );


  buf

  (
    g1389_p_spl_,
    g1389_p
  );


  buf

  (
    g1398_p_spl_,
    g1398_p
  );


  buf

  (
    g1389_n_spl_,
    g1389_n
  );


  buf

  (
    g1401_n_spl_,
    g1401_n
  );


  buf

  (
    g1368_p_spl_,
    g1368_p
  );


  buf

  (
    g1401_p_spl_,
    g1401_p
  );


  buf

  (
    g1368_n_spl_,
    g1368_n
  );


  buf

  (
    g1412_n_spl_,
    g1412_n
  );


  buf

  (
    g1409_n_spl_,
    g1409_n
  );


  buf

  (
    g1412_p_spl_,
    g1412_p
  );


  buf

  (
    g1409_p_spl_,
    g1409_p
  );


  buf

  (
    g1415_p_spl_,
    g1415_p
  );


  buf

  (
    g1415_n_spl_,
    g1415_n
  );


  buf

  (
    g1416_n_spl_,
    g1416_n
  );


  buf

  (
    g1416_p_spl_,
    g1416_p
  );


  buf

  (
    g1420_p_spl_,
    g1420_p
  );


  buf

  (
    g1420_n_spl_,
    g1420_n
  );


  buf

  (
    g1423_p_spl_,
    g1423_p
  );


  buf

  (
    g1423_n_spl_,
    g1423_n
  );


  buf

  (
    g1426_p_spl_,
    g1426_p
  );


  buf

  (
    g1426_n_spl_,
    g1426_n
  );


  buf

  (
    g1432_p_spl_,
    g1432_p
  );


  buf

  (
    g1432_n_spl_,
    g1432_n
  );


  buf

  (
    g1435_p_spl_,
    g1435_p
  );


  buf

  (
    g1435_n_spl_,
    g1435_n
  );


  buf

  (
    g1438_p_spl_,
    g1438_p
  );


  buf

  (
    g1438_n_spl_,
    g1438_n
  );


  buf

  (
    g1441_n_spl_,
    g1441_n
  );


  buf

  (
    g1441_p_spl_,
    g1441_p
  );


  buf

  (
    g1430_n_spl_,
    g1430_n
  );


  buf

  (
    g1430_p_spl_,
    g1430_p
  );


  buf

  (
    G157_n_spl_,
    G157_n
  );


  buf

  (
    G157_n_spl_0,
    G157_n_spl_
  );


  buf

  (
    G157_n_spl_1,
    G157_n_spl_
  );


  buf

  (
    G157_p_spl_,
    G157_p
  );


  buf

  (
    G157_p_spl_0,
    G157_p_spl_
  );


  buf

  (
    G157_p_spl_1,
    G157_p_spl_
  );


  buf

  (
    g1453_n_spl_,
    g1453_n
  );


  buf

  (
    g1453_p_spl_,
    g1453_p
  );


  buf

  (
    g1458_n_spl_,
    g1458_n
  );


  buf

  (
    g1458_n_spl_0,
    g1458_n_spl_
  );


  buf

  (
    g1458_n_spl_1,
    g1458_n_spl_
  );


  buf

  (
    g1458_p_spl_,
    g1458_p
  );


  buf

  (
    g1458_p_spl_0,
    g1458_p_spl_
  );


  buf

  (
    g1458_p_spl_1,
    g1458_p_spl_
  );


  buf

  (
    g1461_p_spl_,
    g1461_p
  );


  buf

  (
    g1456_n_spl_,
    g1456_n
  );


  buf

  (
    g1461_n_spl_,
    g1461_n
  );


  buf

  (
    g1456_p_spl_,
    g1456_p
  );


  buf

  (
    g1464_n_spl_,
    g1464_n
  );


  buf

  (
    g1464_p_spl_,
    g1464_p
  );


  buf

  (
    g1471_n_spl_,
    g1471_n
  );


  buf

  (
    g1471_p_spl_,
    g1471_p
  );


  buf

  (
    g1474_p_spl_,
    g1474_p
  );


  buf

  (
    g1470_n_spl_,
    g1470_n
  );


  buf

  (
    g1474_n_spl_,
    g1474_n
  );


  buf

  (
    g1470_p_spl_,
    g1470_p
  );


  buf

  (
    g1477_p_spl_,
    g1477_p
  );


  buf

  (
    g1469_n_spl_,
    g1469_n
  );


  buf

  (
    g1477_n_spl_,
    g1477_n
  );


  buf

  (
    g1469_p_spl_,
    g1469_p
  );


  buf

  (
    g1483_p_spl_,
    g1483_p
  );


  buf

  (
    g1480_n_spl_,
    g1480_n
  );


  buf

  (
    g1483_n_spl_,
    g1483_n
  );


  buf

  (
    g1480_p_spl_,
    g1480_p
  );


  buf

  (
    g1488_p_spl_,
    g1488_p
  );


  buf

  (
    g1488_n_spl_,
    g1488_n
  );


  buf

  (
    g1491_n_spl_,
    g1491_n
  );


  buf

  (
    g1491_p_spl_,
    g1491_p
  );


  buf

  (
    g1500_n_spl_,
    g1500_n
  );


  buf

  (
    G23_n_spl_,
    G23_n
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    g1509_p_spl_,
    g1509_p
  );


  buf

  (
    g1509_p_spl_0,
    g1509_p_spl_
  );


  buf

  (
    g1509_p_spl_1,
    g1509_p_spl_
  );


  buf

  (
    g1512_p_spl_,
    g1512_p
  );


  buf

  (
    g1512_p_spl_0,
    g1512_p_spl_
  );


  buf

  (
    g1512_p_spl_1,
    g1512_p_spl_
  );


  buf

  (
    G79_n_spl_,
    G79_n
  );


  buf

  (
    G78_n_spl_,
    G78_n
  );


  buf

  (
    G64_n_spl_,
    G64_n
  );


  buf

  (
    G151_n_spl_,
    G151_n
  );


  buf

  (
    G151_n_spl_0,
    G151_n_spl_
  );


  buf

  (
    G152_p_spl_,
    G152_p
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    G1_n_spl_1,
    G1_n_spl_
  );


  buf

  (
    g194_n_spl_,
    g194_n
  );


  buf

  (
    g431_n_spl_,
    g431_n
  );


  buf

  (
    g482_p_spl_,
    g482_p
  );


  buf

  (
    g549_p_spl_,
    g549_p
  );


  buf

  (
    g550_n_spl_,
    g550_n
  );


endmodule
