// Benchmark "mymod" written by ABC on Sun Oct 29 19:31:51 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41,
    G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
    G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
    G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
    G1354, G1355  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
    G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
    G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
    G1354, G1355;
  reg n630_lo, n642_lo, n654_lo, n666_lo, n678_lo, n690_lo, n702_lo,
    n714_lo, n726_lo, n738_lo, n750_lo, n762_lo, n774_lo, n786_lo, n798_lo,
    n810_lo, n822_lo, n834_lo, n846_lo, n858_lo, n870_lo, n882_lo, n894_lo,
    n906_lo, n918_lo, n930_lo, n942_lo, n954_lo, n966_lo, n978_lo, n990_lo,
    n1002_lo, n1005_lo, n1008_lo, n1017_lo, n1020_lo, n1029_lo, n1032_lo,
    n1041_lo, n1044_lo, n1053_lo, n1056_lo, n1065_lo, n1068_lo, n1077_lo,
    n1080_lo, n1089_lo, n1092_lo, n1101_lo, n1104_lo, n1837_o2, n1838_o2,
    n1839_o2, n1840_o2, n1841_o2, n1842_o2, n1843_o2, n1844_o2, n1845_o2,
    n1846_o2, n1847_o2, n1848_o2, n1849_o2, n1850_o2, n1851_o2, n1852_o2,
    n1853_o2, n1854_o2, n1855_o2, n1856_o2, n1857_o2, n1858_o2, n1859_o2,
    n1860_o2, n1861_o2, n1862_o2, n1863_o2, n1864_o2, n1865_o2, n1866_o2,
    n1867_o2, n1868_o2, G834_o2, G847_o2, G860_o2, G873_o2, G925_o2,
    G886_o2, G912_o2, G899_o2, n2151_o2, n2152_o2, n2153_o2, n2154_o2,
    n2155_o2, n2156_o2, n2157_o2, n2158_o2, n2159_o2, n2160_o2, n2161_o2,
    n2162_o2, n2163_o2, n2164_o2, n2165_o2, n2166_o2, n2167_o2, n2168_o2,
    n2169_o2, n2170_o2, n2171_o2, n2172_o2, n2173_o2, n2174_o2, n2175_o2,
    n2176_o2, n2177_o2, n2178_o2, n2179_o2, n2180_o2, n2181_o2, n2182_o2,
    G974_o2, G976_o2, G970_o2, G972_o2, G973_o2, G977_o2, G971_o2, G975_o2,
    G954_o2, G956_o2, G950_o2, G952_o2, G953_o2, G957_o2, G951_o2, G955_o2,
    G986_o2, G991_o2, G770_o2, G773_o2, G776_o2, G779_o2, G782_o2, G785_o2,
    G788_o2, G791_o2, G642_o2, G645_o2, G648_o2, G651_o2, G654_o2, G657_o2,
    G660_o2, G663_o2, G602_o2, G607_o2, G612_o2, G617_o2, G622_o2, G627_o2,
    G632_o2, G637_o2, n627_lo_buf_o2, n639_lo_buf_o2, n651_lo_buf_o2,
    n663_lo_buf_o2, n675_lo_buf_o2, n687_lo_buf_o2, n699_lo_buf_o2,
    n711_lo_buf_o2, n723_lo_buf_o2, n735_lo_buf_o2, n747_lo_buf_o2,
    n759_lo_buf_o2, n771_lo_buf_o2, n783_lo_buf_o2, n795_lo_buf_o2,
    n807_lo_buf_o2, n819_lo_buf_o2, n831_lo_buf_o2, n843_lo_buf_o2,
    n855_lo_buf_o2, n867_lo_buf_o2, n879_lo_buf_o2, n891_lo_buf_o2,
    n903_lo_buf_o2, n915_lo_buf_o2, n927_lo_buf_o2, n939_lo_buf_o2,
    n951_lo_buf_o2, n963_lo_buf_o2, n975_lo_buf_o2, n987_lo_buf_o2,
    n999_lo_buf_o2;
  wire new_n467_, new_n469_, new_n471_, new_n473_, new_n475_, new_n477_,
    new_n479_, new_n481_, new_n483_, new_n485_, new_n487_, new_n489_,
    new_n491_, new_n493_, new_n495_, new_n497_, new_n499_, new_n501_,
    new_n503_, new_n505_, new_n507_, new_n509_, new_n511_, new_n513_,
    new_n515_, new_n517_, new_n519_, new_n521_, new_n523_, new_n525_,
    new_n527_, new_n529_, new_n531_, new_n533_, new_n535_, new_n537_,
    new_n539_, new_n541_, new_n543_, new_n545_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n629_, new_n630_, new_n631_,
    new_n633_, new_n634_, new_n635_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n651_, new_n653_, new_n655_, new_n657_, new_n659_,
    new_n661_, new_n663_, new_n665_, new_n667_, new_n669_, new_n671_,
    new_n673_, new_n675_, new_n677_, new_n679_, new_n681_, new_n683_,
    new_n685_, new_n687_, new_n689_, new_n691_, new_n693_, new_n695_,
    new_n697_, new_n699_, new_n701_, new_n703_, new_n705_, new_n707_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_,
    new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_,
    new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_,
    new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_,
    new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_,
    new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_,
    new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_,
    new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_,
    new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_,
    new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_,
    new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_,
    new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_,
    new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_,
    new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_,
    new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_,
    new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_,
    new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_,
    new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_,
    new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_,
    new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_,
    new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_,
    new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_,
    new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_,
    new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_,
    new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_,
    new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_,
    new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_,
    new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_,
    new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_,
    new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_,
    new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_,
    new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_,
    new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_,
    new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_,
    new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_,
    new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_,
    new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_,
    new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_,
    new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_,
    new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_,
    new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_,
    new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_,
    new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_,
    new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_,
    new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_,
    new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_,
    new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_,
    new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_,
    new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_,
    new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_,
    new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_,
    new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_,
    new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_,
    new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_,
    new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_,
    new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_,
    new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_,
    new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_,
    new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_,
    new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_,
    new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_,
    new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_,
    new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_,
    new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_,
    new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_,
    new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_,
    new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_,
    new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_,
    new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_,
    new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_,
    new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_,
    new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_,
    new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_,
    new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_,
    new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_,
    new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_,
    new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_,
    new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_,
    new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_,
    new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_,
    new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_,
    new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_,
    new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_,
    new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_,
    new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_,
    new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_,
    new_n1718_, new_n1719_, new_n1948_, new_n1949_, new_n1950_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_,
    new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_,
    new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_,
    new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_,
    new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_,
    new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_,
    new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_,
    new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_,
    new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_,
    new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_,
    new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_,
    new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_,
    new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_,
    new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_,
    new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_,
    new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_,
    new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_,
    new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_,
    new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_,
    new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_,
    new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_,
    new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_,
    new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_,
    new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_,
    new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_,
    new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_,
    new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_,
    new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_,
    new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_,
    new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_,
    new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_,
    new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_,
    new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_,
    new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_,
    new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_,
    new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_,
    new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_,
    new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_,
    new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_,
    new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_,
    new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_,
    new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_,
    new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_,
    new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_,
    new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_,
    new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_,
    new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_,
    new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_,
    new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_,
    new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_,
    new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_,
    new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_,
    new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_,
    new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_,
    new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_,
    new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_,
    new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_,
    new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_,
    new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_,
    new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_,
    new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_,
    new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_,
    new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_,
    new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_,
    new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_,
    new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_,
    new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_,
    new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_,
    new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_,
    new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_,
    new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_,
    new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_,
    new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_,
    new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_,
    new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_,
    new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_,
    new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_,
    new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_,
    new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_,
    new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_,
    new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_,
    new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_,
    new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_,
    new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_,
    new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_,
    new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_,
    new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_,
    new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_,
    new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_,
    new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_,
    new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_,
    new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_,
    new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_,
    new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_,
    new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_,
    new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_,
    new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_,
    n630_li, n642_li, n654_li, n666_li, n678_li, n690_li, n702_li, n714_li,
    n726_li, n738_li, n750_li, n762_li, n774_li, n786_li, n798_li, n810_li,
    n822_li, n834_li, n846_li, n858_li, n870_li, n882_li, n894_li, n906_li,
    n918_li, n930_li, n942_li, n954_li, n966_li, n978_li, n990_li,
    n1002_li, n1005_li, n1008_li, n1017_li, n1020_li, n1029_li, n1032_li,
    n1041_li, n1044_li, n1053_li, n1056_li, n1065_li, n1068_li, n1077_li,
    n1080_li, n1089_li, n1092_li, n1101_li, n1104_li, n1837_i2, n1838_i2,
    n1839_i2, n1840_i2, n1841_i2, n1842_i2, n1843_i2, n1844_i2, n1845_i2,
    n1846_i2, n1847_i2, n1848_i2, n1849_i2, n1850_i2, n1851_i2, n1852_i2,
    n1853_i2, n1854_i2, n1855_i2, n1856_i2, n1857_i2, n1858_i2, n1859_i2,
    n1860_i2, n1861_i2, n1862_i2, n1863_i2, n1864_i2, n1865_i2, n1866_i2,
    n1867_i2, n1868_i2, G834_i2, G847_i2, G860_i2, G873_i2, G925_i2,
    G886_i2, G912_i2, G899_i2, n2151_i2, n2152_i2, n2153_i2, n2154_i2,
    n2155_i2, n2156_i2, n2157_i2, n2158_i2, n2159_i2, n2160_i2, n2161_i2,
    n2162_i2, n2163_i2, n2164_i2, n2165_i2, n2166_i2, n2167_i2, n2168_i2,
    n2169_i2, n2170_i2, n2171_i2, n2172_i2, n2173_i2, n2174_i2, n2175_i2,
    n2176_i2, n2177_i2, n2178_i2, n2179_i2, n2180_i2, n2181_i2, n2182_i2,
    G974_i2, G976_i2, G970_i2, G972_i2, G973_i2, G977_i2, G971_i2, G975_i2,
    G954_i2, G956_i2, G950_i2, G952_i2, G953_i2, G957_i2, G951_i2, G955_i2,
    G986_i2, G991_i2, G770_i2, G773_i2, G776_i2, G779_i2, G782_i2, G785_i2,
    G788_i2, G791_i2, G642_i2, G645_i2, G648_i2, G651_i2, G654_i2, G657_i2,
    G660_i2, G663_i2, G602_i2, G607_i2, G612_i2, G617_i2, G622_i2, G627_i2,
    G632_i2, G637_i2, n627_lo_buf_i2, n639_lo_buf_i2, n651_lo_buf_i2,
    n663_lo_buf_i2, n675_lo_buf_i2, n687_lo_buf_i2, n699_lo_buf_i2,
    n711_lo_buf_i2, n723_lo_buf_i2, n735_lo_buf_i2, n747_lo_buf_i2,
    n759_lo_buf_i2, n771_lo_buf_i2, n783_lo_buf_i2, n795_lo_buf_i2,
    n807_lo_buf_i2, n819_lo_buf_i2, n831_lo_buf_i2, n843_lo_buf_i2,
    n855_lo_buf_i2, n867_lo_buf_i2, n879_lo_buf_i2, n891_lo_buf_i2,
    n903_lo_buf_i2, n915_lo_buf_i2, n927_lo_buf_i2, n939_lo_buf_i2,
    n951_lo_buf_i2, n963_lo_buf_i2, n975_lo_buf_i2, n987_lo_buf_i2,
    n999_lo_buf_i2;
  assign new_n467_ = ~G1;
  assign new_n469_ = ~G2;
  assign new_n471_ = ~G3;
  assign new_n473_ = ~G4;
  assign new_n475_ = ~G5;
  assign new_n477_ = ~G6;
  assign new_n479_ = ~G7;
  assign new_n481_ = ~G8;
  assign new_n483_ = ~G9;
  assign new_n485_ = ~G10;
  assign new_n487_ = ~G11;
  assign new_n489_ = ~G12;
  assign new_n491_ = ~G13;
  assign new_n493_ = ~G14;
  assign new_n495_ = ~G15;
  assign new_n497_ = ~G16;
  assign new_n499_ = ~G17;
  assign new_n501_ = ~G18;
  assign new_n503_ = ~G19;
  assign new_n505_ = ~G20;
  assign new_n507_ = ~G21;
  assign new_n509_ = ~G22;
  assign new_n511_ = ~G23;
  assign new_n513_ = ~G24;
  assign new_n515_ = ~G25;
  assign new_n517_ = ~G26;
  assign new_n519_ = ~G27;
  assign new_n521_ = ~G28;
  assign new_n523_ = ~G29;
  assign new_n525_ = ~G30;
  assign new_n527_ = ~G31;
  assign new_n529_ = ~G32;
  assign new_n531_ = ~G33;
  assign new_n533_ = ~G34;
  assign new_n535_ = ~G35;
  assign new_n537_ = ~G36;
  assign new_n539_ = ~G37;
  assign new_n541_ = ~G38;
  assign new_n543_ = ~G39;
  assign new_n545_ = ~G40;
  assign new_n547_ = ~G41;
  assign new_n548_ = n630_lo;
  assign new_n549_ = ~n630_lo;
  assign new_n550_ = n642_lo;
  assign new_n551_ = ~n642_lo;
  assign new_n552_ = n654_lo;
  assign new_n553_ = ~n654_lo;
  assign new_n554_ = n666_lo;
  assign new_n555_ = ~n666_lo;
  assign new_n556_ = n678_lo;
  assign new_n557_ = ~n678_lo;
  assign new_n558_ = n690_lo;
  assign new_n559_ = ~n690_lo;
  assign new_n560_ = n702_lo;
  assign new_n561_ = ~n702_lo;
  assign new_n562_ = n714_lo;
  assign new_n563_ = ~n714_lo;
  assign new_n564_ = n726_lo;
  assign new_n565_ = ~n726_lo;
  assign new_n566_ = n738_lo;
  assign new_n567_ = ~n738_lo;
  assign new_n568_ = n750_lo;
  assign new_n569_ = ~n750_lo;
  assign new_n570_ = n762_lo;
  assign new_n571_ = ~n762_lo;
  assign new_n572_ = n774_lo;
  assign new_n573_ = ~n774_lo;
  assign new_n574_ = n786_lo;
  assign new_n575_ = ~n786_lo;
  assign new_n576_ = n798_lo;
  assign new_n577_ = ~n798_lo;
  assign new_n578_ = n810_lo;
  assign new_n579_ = ~n810_lo;
  assign new_n580_ = n822_lo;
  assign new_n581_ = ~n822_lo;
  assign new_n582_ = n834_lo;
  assign new_n583_ = ~n834_lo;
  assign new_n584_ = n846_lo;
  assign new_n585_ = ~n846_lo;
  assign new_n586_ = n858_lo;
  assign new_n587_ = ~n858_lo;
  assign new_n588_ = n870_lo;
  assign new_n589_ = ~n870_lo;
  assign new_n590_ = n882_lo;
  assign new_n591_ = ~n882_lo;
  assign new_n592_ = n894_lo;
  assign new_n593_ = ~n894_lo;
  assign new_n594_ = n906_lo;
  assign new_n595_ = ~n906_lo;
  assign new_n596_ = n918_lo;
  assign new_n597_ = ~n918_lo;
  assign new_n598_ = n930_lo;
  assign new_n599_ = ~n930_lo;
  assign new_n600_ = n942_lo;
  assign new_n601_ = ~n942_lo;
  assign new_n602_ = n954_lo;
  assign new_n603_ = ~n954_lo;
  assign new_n604_ = n966_lo;
  assign new_n605_ = ~n966_lo;
  assign new_n606_ = n978_lo;
  assign new_n607_ = ~n978_lo;
  assign new_n608_ = n990_lo;
  assign new_n609_ = ~n990_lo;
  assign new_n610_ = n1002_lo;
  assign new_n611_ = ~n1002_lo;
  assign new_n613_ = ~n1005_lo;
  assign new_n614_ = n1008_lo;
  assign new_n615_ = ~n1008_lo;
  assign new_n617_ = ~n1017_lo;
  assign new_n618_ = n1020_lo;
  assign new_n619_ = ~n1020_lo;
  assign new_n621_ = ~n1029_lo;
  assign new_n622_ = n1032_lo;
  assign new_n623_ = ~n1032_lo;
  assign new_n625_ = ~n1041_lo;
  assign new_n626_ = n1044_lo;
  assign new_n627_ = ~n1044_lo;
  assign new_n629_ = ~n1053_lo;
  assign new_n630_ = n1056_lo;
  assign new_n631_ = ~n1056_lo;
  assign new_n633_ = ~n1065_lo;
  assign new_n634_ = n1068_lo;
  assign new_n635_ = ~n1068_lo;
  assign new_n637_ = ~n1077_lo;
  assign new_n638_ = n1080_lo;
  assign new_n639_ = ~n1080_lo;
  assign new_n641_ = ~n1089_lo;
  assign new_n642_ = n1092_lo;
  assign new_n643_ = ~n1092_lo;
  assign new_n645_ = ~n1101_lo;
  assign new_n646_ = n1104_lo;
  assign new_n647_ = ~n1104_lo;
  assign new_n649_ = ~n1837_o2;
  assign new_n651_ = ~n1838_o2;
  assign new_n653_ = ~n1839_o2;
  assign new_n655_ = ~n1840_o2;
  assign new_n657_ = ~n1841_o2;
  assign new_n659_ = ~n1842_o2;
  assign new_n661_ = ~n1843_o2;
  assign new_n663_ = ~n1844_o2;
  assign new_n665_ = ~n1845_o2;
  assign new_n667_ = ~n1846_o2;
  assign new_n669_ = ~n1847_o2;
  assign new_n671_ = ~n1848_o2;
  assign new_n673_ = ~n1849_o2;
  assign new_n675_ = ~n1850_o2;
  assign new_n677_ = ~n1851_o2;
  assign new_n679_ = ~n1852_o2;
  assign new_n681_ = ~n1853_o2;
  assign new_n683_ = ~n1854_o2;
  assign new_n685_ = ~n1855_o2;
  assign new_n687_ = ~n1856_o2;
  assign new_n689_ = ~n1857_o2;
  assign new_n691_ = ~n1858_o2;
  assign new_n693_ = ~n1859_o2;
  assign new_n695_ = ~n1860_o2;
  assign new_n697_ = ~n1861_o2;
  assign new_n699_ = ~n1862_o2;
  assign new_n701_ = ~n1863_o2;
  assign new_n703_ = ~n1864_o2;
  assign new_n705_ = ~n1865_o2;
  assign new_n707_ = ~n1866_o2;
  assign new_n709_ = ~n1867_o2;
  assign new_n711_ = ~n1868_o2;
  assign new_n712_ = G834_o2;
  assign new_n713_ = ~G834_o2;
  assign new_n714_ = G847_o2;
  assign new_n715_ = ~G847_o2;
  assign new_n716_ = G860_o2;
  assign new_n717_ = ~G860_o2;
  assign new_n718_ = G873_o2;
  assign new_n719_ = ~G873_o2;
  assign new_n720_ = G925_o2;
  assign new_n721_ = ~G925_o2;
  assign new_n722_ = G886_o2;
  assign new_n723_ = ~G886_o2;
  assign new_n724_ = G912_o2;
  assign new_n725_ = ~G912_o2;
  assign new_n726_ = G899_o2;
  assign new_n727_ = ~G899_o2;
  assign new_n728_ = n2151_o2;
  assign new_n729_ = ~n2151_o2;
  assign new_n730_ = n2152_o2;
  assign new_n731_ = ~n2152_o2;
  assign new_n732_ = n2153_o2;
  assign new_n733_ = ~n2153_o2;
  assign new_n734_ = n2154_o2;
  assign new_n735_ = ~n2154_o2;
  assign new_n736_ = n2155_o2;
  assign new_n737_ = ~n2155_o2;
  assign new_n738_ = n2156_o2;
  assign new_n739_ = ~n2156_o2;
  assign new_n740_ = n2157_o2;
  assign new_n741_ = ~n2157_o2;
  assign new_n742_ = n2158_o2;
  assign new_n743_ = ~n2158_o2;
  assign new_n744_ = n2159_o2;
  assign new_n745_ = ~n2159_o2;
  assign new_n746_ = n2160_o2;
  assign new_n747_ = ~n2160_o2;
  assign new_n748_ = n2161_o2;
  assign new_n749_ = ~n2161_o2;
  assign new_n750_ = n2162_o2;
  assign new_n751_ = ~n2162_o2;
  assign new_n752_ = n2163_o2;
  assign new_n753_ = ~n2163_o2;
  assign new_n754_ = n2164_o2;
  assign new_n755_ = ~n2164_o2;
  assign new_n756_ = n2165_o2;
  assign new_n757_ = ~n2165_o2;
  assign new_n758_ = n2166_o2;
  assign new_n759_ = ~n2166_o2;
  assign new_n760_ = n2167_o2;
  assign new_n761_ = ~n2167_o2;
  assign new_n762_ = n2168_o2;
  assign new_n763_ = ~n2168_o2;
  assign new_n764_ = n2169_o2;
  assign new_n765_ = ~n2169_o2;
  assign new_n766_ = n2170_o2;
  assign new_n767_ = ~n2170_o2;
  assign new_n768_ = n2171_o2;
  assign new_n769_ = ~n2171_o2;
  assign new_n770_ = n2172_o2;
  assign new_n771_ = ~n2172_o2;
  assign new_n772_ = n2173_o2;
  assign new_n773_ = ~n2173_o2;
  assign new_n774_ = n2174_o2;
  assign new_n775_ = ~n2174_o2;
  assign new_n776_ = n2175_o2;
  assign new_n777_ = ~n2175_o2;
  assign new_n778_ = n2176_o2;
  assign new_n779_ = ~n2176_o2;
  assign new_n780_ = n2177_o2;
  assign new_n781_ = ~n2177_o2;
  assign new_n782_ = n2178_o2;
  assign new_n783_ = ~n2178_o2;
  assign new_n784_ = n2179_o2;
  assign new_n785_ = ~n2179_o2;
  assign new_n786_ = n2180_o2;
  assign new_n787_ = ~n2180_o2;
  assign new_n788_ = n2181_o2;
  assign new_n789_ = ~n2181_o2;
  assign new_n790_ = n2182_o2;
  assign new_n791_ = ~n2182_o2;
  assign new_n792_ = G974_o2;
  assign new_n793_ = ~G974_o2;
  assign new_n794_ = G976_o2;
  assign new_n795_ = ~G976_o2;
  assign new_n796_ = G970_o2;
  assign new_n797_ = ~G970_o2;
  assign new_n798_ = G972_o2;
  assign new_n799_ = ~G972_o2;
  assign new_n800_ = G973_o2;
  assign new_n801_ = ~G973_o2;
  assign new_n802_ = G977_o2;
  assign new_n803_ = ~G977_o2;
  assign new_n804_ = G971_o2;
  assign new_n805_ = ~G971_o2;
  assign new_n806_ = G975_o2;
  assign new_n807_ = ~G975_o2;
  assign new_n808_ = G954_o2;
  assign new_n809_ = ~G954_o2;
  assign new_n810_ = G956_o2;
  assign new_n811_ = ~G956_o2;
  assign new_n812_ = G950_o2;
  assign new_n813_ = ~G950_o2;
  assign new_n814_ = G952_o2;
  assign new_n815_ = ~G952_o2;
  assign new_n816_ = G953_o2;
  assign new_n817_ = ~G953_o2;
  assign new_n818_ = G957_o2;
  assign new_n819_ = ~G957_o2;
  assign new_n820_ = G951_o2;
  assign new_n821_ = ~G951_o2;
  assign new_n822_ = G955_o2;
  assign new_n823_ = ~G955_o2;
  assign new_n824_ = G986_o2;
  assign new_n825_ = ~G986_o2;
  assign new_n826_ = G991_o2;
  assign new_n827_ = ~G991_o2;
  assign new_n828_ = G770_o2;
  assign new_n829_ = ~G770_o2;
  assign new_n830_ = G773_o2;
  assign new_n831_ = ~G773_o2;
  assign new_n832_ = G776_o2;
  assign new_n833_ = ~G776_o2;
  assign new_n834_ = G779_o2;
  assign new_n835_ = ~G779_o2;
  assign new_n836_ = G782_o2;
  assign new_n837_ = ~G782_o2;
  assign new_n838_ = G785_o2;
  assign new_n839_ = ~G785_o2;
  assign new_n840_ = G788_o2;
  assign new_n841_ = ~G788_o2;
  assign new_n842_ = G791_o2;
  assign new_n843_ = ~G791_o2;
  assign new_n844_ = G642_o2;
  assign new_n845_ = ~G642_o2;
  assign new_n846_ = G645_o2;
  assign new_n847_ = ~G645_o2;
  assign new_n848_ = G648_o2;
  assign new_n849_ = ~G648_o2;
  assign new_n850_ = G651_o2;
  assign new_n851_ = ~G651_o2;
  assign new_n852_ = G654_o2;
  assign new_n853_ = ~G654_o2;
  assign new_n854_ = G657_o2;
  assign new_n855_ = ~G657_o2;
  assign new_n856_ = G660_o2;
  assign new_n857_ = ~G660_o2;
  assign new_n858_ = G663_o2;
  assign new_n859_ = ~G663_o2;
  assign new_n860_ = G602_o2;
  assign new_n861_ = ~G602_o2;
  assign new_n862_ = G607_o2;
  assign new_n863_ = ~G607_o2;
  assign new_n864_ = G612_o2;
  assign new_n865_ = ~G612_o2;
  assign new_n866_ = G617_o2;
  assign new_n867_ = ~G617_o2;
  assign new_n868_ = G622_o2;
  assign new_n869_ = ~G622_o2;
  assign new_n870_ = G627_o2;
  assign new_n871_ = ~G627_o2;
  assign new_n872_ = G632_o2;
  assign new_n873_ = ~G632_o2;
  assign new_n874_ = G637_o2;
  assign new_n875_ = ~G637_o2;
  assign new_n876_ = n627_lo_buf_o2;
  assign new_n877_ = ~n627_lo_buf_o2;
  assign new_n878_ = n639_lo_buf_o2;
  assign new_n879_ = ~n639_lo_buf_o2;
  assign new_n880_ = n651_lo_buf_o2;
  assign new_n881_ = ~n651_lo_buf_o2;
  assign new_n882_ = n663_lo_buf_o2;
  assign new_n883_ = ~n663_lo_buf_o2;
  assign new_n884_ = n675_lo_buf_o2;
  assign new_n885_ = ~n675_lo_buf_o2;
  assign new_n886_ = n687_lo_buf_o2;
  assign new_n887_ = ~n687_lo_buf_o2;
  assign new_n888_ = n699_lo_buf_o2;
  assign new_n889_ = ~n699_lo_buf_o2;
  assign new_n890_ = n711_lo_buf_o2;
  assign new_n891_ = ~n711_lo_buf_o2;
  assign new_n892_ = n723_lo_buf_o2;
  assign new_n893_ = ~n723_lo_buf_o2;
  assign new_n894_ = n735_lo_buf_o2;
  assign new_n895_ = ~n735_lo_buf_o2;
  assign new_n896_ = n747_lo_buf_o2;
  assign new_n897_ = ~n747_lo_buf_o2;
  assign new_n898_ = n759_lo_buf_o2;
  assign new_n899_ = ~n759_lo_buf_o2;
  assign new_n900_ = n771_lo_buf_o2;
  assign new_n901_ = ~n771_lo_buf_o2;
  assign new_n902_ = n783_lo_buf_o2;
  assign new_n903_ = ~n783_lo_buf_o2;
  assign new_n904_ = n795_lo_buf_o2;
  assign new_n905_ = ~n795_lo_buf_o2;
  assign new_n906_ = n807_lo_buf_o2;
  assign new_n907_ = ~n807_lo_buf_o2;
  assign new_n908_ = n819_lo_buf_o2;
  assign new_n909_ = ~n819_lo_buf_o2;
  assign new_n910_ = n831_lo_buf_o2;
  assign new_n911_ = ~n831_lo_buf_o2;
  assign new_n912_ = n843_lo_buf_o2;
  assign new_n913_ = ~n843_lo_buf_o2;
  assign new_n914_ = n855_lo_buf_o2;
  assign new_n915_ = ~n855_lo_buf_o2;
  assign new_n916_ = n867_lo_buf_o2;
  assign new_n917_ = ~n867_lo_buf_o2;
  assign new_n918_ = n879_lo_buf_o2;
  assign new_n919_ = ~n879_lo_buf_o2;
  assign new_n920_ = n891_lo_buf_o2;
  assign new_n921_ = ~n891_lo_buf_o2;
  assign new_n922_ = n903_lo_buf_o2;
  assign new_n923_ = ~n903_lo_buf_o2;
  assign new_n924_ = n915_lo_buf_o2;
  assign new_n925_ = ~n915_lo_buf_o2;
  assign new_n926_ = n927_lo_buf_o2;
  assign new_n927_ = ~n927_lo_buf_o2;
  assign new_n928_ = n939_lo_buf_o2;
  assign new_n929_ = ~n939_lo_buf_o2;
  assign new_n930_ = n951_lo_buf_o2;
  assign new_n931_ = ~n951_lo_buf_o2;
  assign new_n932_ = n963_lo_buf_o2;
  assign new_n933_ = ~n963_lo_buf_o2;
  assign new_n934_ = n975_lo_buf_o2;
  assign new_n935_ = ~n975_lo_buf_o2;
  assign new_n936_ = n987_lo_buf_o2;
  assign new_n937_ = ~n987_lo_buf_o2;
  assign new_n938_ = n999_lo_buf_o2;
  assign new_n939_ = ~n999_lo_buf_o2;
  assign new_n940_ = new_n813_ & new_n1950_;
  assign new_n941_ = new_n812_ | new_n1955_;
  assign new_n942_ = new_n940_ & new_n1960_;
  assign new_n943_ = new_n941_ | new_n1965_;
  assign new_n944_ = new_n942_ & new_n821_;
  assign new_n945_ = new_n943_ | new_n820_;
  assign new_n946_ = new_n944_ & new_n1969_;
  assign new_n947_ = new_n945_ | new_n1972_;
  assign new_n948_ = new_n1975_ & new_n1979_;
  assign new_n949_ = new_n1983_ | new_n1987_;
  assign new_n950_ = new_n949_ | new_n549_;
  assign new_n951_ = new_n1990_ & new_n548_;
  assign new_n952_ = new_n1990_ & new_n948_;
  assign new_n953_ = new_n952_ | new_n951_;
  assign new_n954_ = new_n1975_ & new_n1993_;
  assign new_n955_ = new_n1983_ | new_n1998_;
  assign new_n956_ = new_n955_ | new_n551_;
  assign new_n957_ = new_n2001_ & new_n550_;
  assign new_n958_ = new_n2001_ & new_n954_;
  assign new_n959_ = new_n958_ | new_n957_;
  assign new_n960_ = new_n1976_ & new_n2004_;
  assign new_n961_ = new_n1984_ | new_n2009_;
  assign new_n962_ = new_n961_ | new_n553_;
  assign new_n963_ = new_n2012_ & new_n552_;
  assign new_n964_ = new_n2012_ & new_n960_;
  assign new_n965_ = new_n964_ | new_n963_;
  assign new_n966_ = new_n1976_ & new_n2015_;
  assign new_n967_ = new_n1984_ | new_n2020_;
  assign new_n968_ = new_n967_ | new_n555_;
  assign new_n969_ = new_n2023_ & new_n554_;
  assign new_n970_ = new_n2023_ & new_n966_;
  assign new_n971_ = new_n970_ | new_n969_;
  assign new_n972_ = new_n815_ & new_n1950_;
  assign new_n973_ = new_n814_ | new_n1955_;
  assign new_n974_ = new_n972_ & new_n817_;
  assign new_n975_ = new_n973_ | new_n816_;
  assign new_n976_ = new_n974_ & new_n2026_;
  assign new_n977_ = new_n975_ | new_n2031_;
  assign new_n978_ = new_n976_ & new_n1969_;
  assign new_n979_ = new_n977_ | new_n1972_;
  assign new_n980_ = new_n2035_ & new_n1979_;
  assign new_n981_ = new_n2038_ | new_n1987_;
  assign new_n982_ = new_n981_ | new_n557_;
  assign new_n983_ = new_n2040_ & new_n556_;
  assign new_n984_ = new_n2040_ & new_n980_;
  assign new_n985_ = new_n984_ | new_n983_;
  assign new_n986_ = new_n2035_ & new_n1993_;
  assign new_n987_ = new_n2038_ | new_n1998_;
  assign new_n988_ = new_n987_ | new_n559_;
  assign new_n989_ = new_n2041_ & new_n558_;
  assign new_n990_ = new_n2041_ & new_n986_;
  assign new_n991_ = new_n990_ | new_n989_;
  assign new_n992_ = new_n2036_ & new_n2004_;
  assign new_n993_ = new_n2039_ | new_n2009_;
  assign new_n994_ = new_n993_ | new_n561_;
  assign new_n995_ = new_n2042_ & new_n560_;
  assign new_n996_ = new_n2042_ & new_n992_;
  assign new_n997_ = new_n996_ | new_n995_;
  assign new_n998_ = new_n2036_ & new_n2015_;
  assign new_n999_ = new_n2039_ | new_n2020_;
  assign new_n1000_ = new_n999_ | new_n563_;
  assign new_n1001_ = new_n2043_ & new_n562_;
  assign new_n1002_ = new_n2043_ & new_n998_;
  assign new_n1003_ = new_n1002_ | new_n1001_;
  assign new_n1004_ = new_n809_ & new_n2046_;
  assign new_n1005_ = new_n808_ | new_n2051_;
  assign new_n1006_ = new_n1004_ & new_n1960_;
  assign new_n1007_ = new_n1005_ | new_n1965_;
  assign new_n1008_ = new_n1006_ & new_n823_;
  assign new_n1009_ = new_n1007_ | new_n822_;
  assign new_n1010_ = new_n1008_ & new_n1970_;
  assign new_n1011_ = new_n1009_ | new_n1973_;
  assign new_n1012_ = new_n2055_ & new_n1980_;
  assign new_n1013_ = new_n2058_ | new_n1988_;
  assign new_n1014_ = new_n1013_ | new_n565_;
  assign new_n1015_ = new_n2060_ & new_n564_;
  assign new_n1016_ = new_n2060_ & new_n1012_;
  assign new_n1017_ = new_n1016_ | new_n1015_;
  assign new_n1018_ = new_n2055_ & new_n1994_;
  assign new_n1019_ = new_n2058_ | new_n1999_;
  assign new_n1020_ = new_n1019_ | new_n567_;
  assign new_n1021_ = new_n2061_ & new_n566_;
  assign new_n1022_ = new_n2061_ & new_n1018_;
  assign new_n1023_ = new_n1022_ | new_n1021_;
  assign new_n1024_ = new_n2056_ & new_n2005_;
  assign new_n1025_ = new_n2059_ | new_n2010_;
  assign new_n1026_ = new_n1025_ | new_n569_;
  assign new_n1027_ = new_n2062_ & new_n568_;
  assign new_n1028_ = new_n2062_ & new_n1024_;
  assign new_n1029_ = new_n1028_ | new_n1027_;
  assign new_n1030_ = new_n2056_ & new_n2016_;
  assign new_n1031_ = new_n2059_ | new_n2021_;
  assign new_n1032_ = new_n1031_ | new_n571_;
  assign new_n1033_ = new_n2063_ & new_n570_;
  assign new_n1034_ = new_n2063_ & new_n1030_;
  assign new_n1035_ = new_n1034_ | new_n1033_;
  assign new_n1036_ = new_n811_ & new_n2046_;
  assign new_n1037_ = new_n810_ | new_n2051_;
  assign new_n1038_ = new_n1036_ & new_n819_;
  assign new_n1039_ = new_n1037_ | new_n818_;
  assign new_n1040_ = new_n1038_ & new_n2026_;
  assign new_n1041_ = new_n1039_ | new_n2031_;
  assign new_n1042_ = new_n1040_ & new_n1970_;
  assign new_n1043_ = new_n1041_ | new_n1973_;
  assign new_n1044_ = new_n2065_ & new_n1980_;
  assign new_n1045_ = new_n2068_ | new_n1988_;
  assign new_n1046_ = new_n1045_ | new_n573_;
  assign new_n1047_ = new_n2070_ & new_n572_;
  assign new_n1048_ = new_n2070_ & new_n1044_;
  assign new_n1049_ = new_n1048_ | new_n1047_;
  assign new_n1050_ = new_n2065_ & new_n1994_;
  assign new_n1051_ = new_n2068_ | new_n1999_;
  assign new_n1052_ = new_n1051_ | new_n575_;
  assign new_n1053_ = new_n2071_ & new_n574_;
  assign new_n1054_ = new_n2071_ & new_n1050_;
  assign new_n1055_ = new_n1054_ | new_n1053_;
  assign new_n1056_ = new_n2066_ & new_n2005_;
  assign new_n1057_ = new_n2069_ | new_n2010_;
  assign new_n1058_ = new_n1057_ | new_n577_;
  assign new_n1059_ = new_n2072_ & new_n576_;
  assign new_n1060_ = new_n2072_ & new_n1056_;
  assign new_n1061_ = new_n1060_ | new_n1059_;
  assign new_n1062_ = new_n2066_ & new_n2016_;
  assign new_n1063_ = new_n2069_ | new_n2021_;
  assign new_n1064_ = new_n1063_ | new_n579_;
  assign new_n1065_ = new_n2073_ & new_n578_;
  assign new_n1066_ = new_n2073_ & new_n1062_;
  assign new_n1067_ = new_n1066_ | new_n1065_;
  assign new_n1068_ = new_n797_ & new_n1981_;
  assign new_n1069_ = new_n796_ | new_n1989_;
  assign new_n1070_ = new_n1068_ & new_n2006_;
  assign new_n1071_ = new_n1069_ | new_n2011_;
  assign new_n1072_ = new_n1070_ & new_n805_;
  assign new_n1073_ = new_n1071_ | new_n804_;
  assign new_n1074_ = new_n1072_ & new_n2075_;
  assign new_n1075_ = new_n1073_ | new_n2078_;
  assign new_n1076_ = new_n2081_ & new_n1951_;
  assign new_n1077_ = new_n2084_ | new_n1956_;
  assign new_n1078_ = new_n1077_ | new_n581_;
  assign new_n1079_ = new_n2086_ & new_n580_;
  assign new_n1080_ = new_n2086_ & new_n1076_;
  assign new_n1081_ = new_n1080_ | new_n1079_;
  assign new_n1082_ = new_n2081_ & new_n2047_;
  assign new_n1083_ = new_n2084_ | new_n2052_;
  assign new_n1084_ = new_n1083_ | new_n583_;
  assign new_n1085_ = new_n2087_ & new_n582_;
  assign new_n1086_ = new_n2087_ & new_n1082_;
  assign new_n1087_ = new_n1086_ | new_n1085_;
  assign new_n1088_ = new_n2082_ & new_n1961_;
  assign new_n1089_ = new_n2085_ | new_n1966_;
  assign new_n1090_ = new_n1089_ | new_n585_;
  assign new_n1091_ = new_n2088_ & new_n584_;
  assign new_n1092_ = new_n2088_ & new_n1088_;
  assign new_n1093_ = new_n1092_ | new_n1091_;
  assign new_n1094_ = new_n2082_ & new_n2027_;
  assign new_n1095_ = new_n2085_ | new_n2032_;
  assign new_n1096_ = new_n1095_ | new_n587_;
  assign new_n1097_ = new_n2089_ & new_n586_;
  assign new_n1098_ = new_n2089_ & new_n1094_;
  assign new_n1099_ = new_n1098_ | new_n1097_;
  assign new_n1100_ = new_n799_ & new_n1981_;
  assign new_n1101_ = new_n798_ | new_n1989_;
  assign new_n1102_ = new_n1100_ & new_n801_;
  assign new_n1103_ = new_n1101_ | new_n800_;
  assign new_n1104_ = new_n1102_ & new_n2017_;
  assign new_n1105_ = new_n1103_ | new_n2022_;
  assign new_n1106_ = new_n1104_ & new_n2075_;
  assign new_n1107_ = new_n1105_ | new_n2078_;
  assign new_n1108_ = new_n2091_ & new_n1951_;
  assign new_n1109_ = new_n2094_ | new_n1956_;
  assign new_n1110_ = new_n1109_ | new_n589_;
  assign new_n1111_ = new_n2096_ & new_n588_;
  assign new_n1112_ = new_n2096_ & new_n1108_;
  assign new_n1113_ = new_n1112_ | new_n1111_;
  assign new_n1114_ = new_n2091_ & new_n2047_;
  assign new_n1115_ = new_n2094_ | new_n2052_;
  assign new_n1116_ = new_n1115_ | new_n591_;
  assign new_n1117_ = new_n2097_ & new_n590_;
  assign new_n1118_ = new_n2097_ & new_n1114_;
  assign new_n1119_ = new_n1118_ | new_n1117_;
  assign new_n1120_ = new_n2092_ & new_n1961_;
  assign new_n1121_ = new_n2095_ | new_n1966_;
  assign new_n1122_ = new_n1121_ | new_n593_;
  assign new_n1123_ = new_n2098_ & new_n592_;
  assign new_n1124_ = new_n2098_ & new_n1120_;
  assign new_n1125_ = new_n1124_ | new_n1123_;
  assign new_n1126_ = new_n2092_ & new_n2027_;
  assign new_n1127_ = new_n2095_ | new_n2032_;
  assign new_n1128_ = new_n1127_ | new_n595_;
  assign new_n1129_ = new_n2099_ & new_n594_;
  assign new_n1130_ = new_n2099_ & new_n1126_;
  assign new_n1131_ = new_n1130_ | new_n1129_;
  assign new_n1132_ = new_n793_ & new_n1995_;
  assign new_n1133_ = new_n792_ | new_n2000_;
  assign new_n1134_ = new_n1132_ & new_n2006_;
  assign new_n1135_ = new_n1133_ | new_n2011_;
  assign new_n1136_ = new_n1134_ & new_n807_;
  assign new_n1137_ = new_n1135_ | new_n806_;
  assign new_n1138_ = new_n1136_ & new_n2076_;
  assign new_n1139_ = new_n1137_ | new_n2079_;
  assign new_n1140_ = new_n2101_ & new_n1952_;
  assign new_n1141_ = new_n2104_ | new_n1957_;
  assign new_n1142_ = new_n1141_ | new_n597_;
  assign new_n1143_ = new_n2106_ & new_n596_;
  assign new_n1144_ = new_n2106_ & new_n1140_;
  assign new_n1145_ = new_n1144_ | new_n1143_;
  assign new_n1146_ = new_n2101_ & new_n2048_;
  assign new_n1147_ = new_n2104_ | new_n2053_;
  assign new_n1148_ = new_n1147_ | new_n599_;
  assign new_n1149_ = new_n2107_ & new_n598_;
  assign new_n1150_ = new_n2107_ & new_n1146_;
  assign new_n1151_ = new_n1150_ | new_n1149_;
  assign new_n1152_ = new_n2102_ & new_n1962_;
  assign new_n1153_ = new_n2105_ | new_n1967_;
  assign new_n1154_ = new_n1153_ | new_n601_;
  assign new_n1155_ = new_n2108_ & new_n600_;
  assign new_n1156_ = new_n2108_ & new_n1152_;
  assign new_n1157_ = new_n1156_ | new_n1155_;
  assign new_n1158_ = new_n2102_ & new_n2028_;
  assign new_n1159_ = new_n2105_ | new_n2033_;
  assign new_n1160_ = new_n1159_ | new_n603_;
  assign new_n1161_ = new_n2109_ & new_n602_;
  assign new_n1162_ = new_n2109_ & new_n1158_;
  assign new_n1163_ = new_n1162_ | new_n1161_;
  assign new_n1164_ = new_n795_ & new_n1995_;
  assign new_n1165_ = new_n794_ | new_n2000_;
  assign new_n1166_ = new_n1164_ & new_n803_;
  assign new_n1167_ = new_n1165_ | new_n802_;
  assign new_n1168_ = new_n1166_ & new_n2017_;
  assign new_n1169_ = new_n1167_ | new_n2022_;
  assign new_n1170_ = new_n1168_ & new_n2076_;
  assign new_n1171_ = new_n1169_ | new_n2079_;
  assign new_n1172_ = new_n2111_ & new_n1952_;
  assign new_n1173_ = new_n2114_ | new_n1957_;
  assign new_n1174_ = new_n1173_ | new_n605_;
  assign new_n1175_ = new_n2116_ & new_n604_;
  assign new_n1176_ = new_n2116_ & new_n1172_;
  assign new_n1177_ = new_n1176_ | new_n1175_;
  assign new_n1178_ = new_n2111_ & new_n2048_;
  assign new_n1179_ = new_n2114_ | new_n2053_;
  assign new_n1180_ = new_n1179_ | new_n607_;
  assign new_n1181_ = new_n2117_ & new_n606_;
  assign new_n1182_ = new_n2117_ & new_n1178_;
  assign new_n1183_ = new_n1182_ | new_n1181_;
  assign new_n1184_ = new_n2112_ & new_n1962_;
  assign new_n1185_ = new_n2115_ | new_n1967_;
  assign new_n1186_ = new_n1185_ | new_n609_;
  assign new_n1187_ = new_n2118_ & new_n608_;
  assign new_n1188_ = new_n2118_ & new_n1184_;
  assign new_n1189_ = new_n1188_ | new_n1187_;
  assign new_n1190_ = new_n2112_ & new_n2028_;
  assign new_n1191_ = new_n2115_ | new_n2033_;
  assign new_n1192_ = new_n1191_ | new_n611_;
  assign new_n1193_ = new_n2119_ & new_n610_;
  assign new_n1194_ = new_n2119_ & new_n1190_;
  assign new_n1195_ = new_n1194_ | new_n1193_;
  assign new_n1196_ = new_n2120_ & new_n2121_;
  assign new_n1197_ = new_n2122_ | new_n2123_;
  assign new_n1198_ = new_n2124_ & new_n2120_;
  assign new_n1199_ = new_n2125_ | new_n2122_;
  assign new_n1200_ = new_n2124_ & new_n2121_;
  assign new_n1201_ = new_n2125_ | new_n2123_;
  assign new_n1202_ = new_n1201_ & new_n1199_;
  assign new_n1203_ = new_n1200_ | new_n1198_;
  assign new_n1204_ = new_n2126_ & new_n2127_;
  assign new_n1205_ = new_n2128_ | new_n2129_;
  assign new_n1206_ = new_n2130_ & new_n2126_;
  assign new_n1207_ = new_n2131_ | new_n2128_;
  assign new_n1208_ = new_n2130_ & new_n2127_;
  assign new_n1209_ = new_n2131_ | new_n2129_;
  assign new_n1210_ = new_n1209_ & new_n1207_;
  assign new_n1211_ = new_n1208_ | new_n1206_;
  assign new_n1212_ = new_n2132_ & new_n2133_;
  assign new_n1213_ = new_n2134_ | new_n2135_;
  assign new_n1214_ = new_n2136_ & new_n2132_;
  assign new_n1215_ = new_n2137_ | new_n2134_;
  assign new_n1216_ = new_n2136_ & new_n2133_;
  assign new_n1217_ = new_n2137_ | new_n2135_;
  assign new_n1218_ = new_n1217_ & new_n1215_;
  assign new_n1219_ = new_n1216_ | new_n1214_;
  assign new_n1220_ = new_n2138_ & new_n2139_;
  assign new_n1221_ = new_n2140_ | new_n2141_;
  assign new_n1222_ = new_n2142_ & new_n2138_;
  assign new_n1223_ = new_n2143_ | new_n2140_;
  assign new_n1224_ = new_n2142_ & new_n2139_;
  assign new_n1225_ = new_n2143_ | new_n2141_;
  assign new_n1226_ = new_n1225_ & new_n1223_;
  assign new_n1227_ = new_n1224_ | new_n1222_;
  assign new_n1228_ = new_n2144_ & new_n2145_;
  assign new_n1229_ = new_n2146_ | new_n2147_;
  assign new_n1230_ = new_n2148_ & new_n2144_;
  assign new_n1231_ = new_n2149_ | new_n2146_;
  assign new_n1232_ = new_n2148_ & new_n2145_;
  assign new_n1233_ = new_n2149_ | new_n2147_;
  assign new_n1234_ = new_n1233_ & new_n1231_;
  assign new_n1235_ = new_n1232_ | new_n1230_;
  assign new_n1236_ = new_n2150_ & new_n2151_;
  assign new_n1237_ = new_n2152_ | new_n2153_;
  assign new_n1238_ = new_n2154_ & new_n2150_;
  assign new_n1239_ = new_n2155_ | new_n2152_;
  assign new_n1240_ = new_n2154_ & new_n2151_;
  assign new_n1241_ = new_n2155_ | new_n2153_;
  assign new_n1242_ = new_n1241_ & new_n1239_;
  assign new_n1243_ = new_n1240_ | new_n1238_;
  assign new_n1244_ = new_n2156_ & new_n2157_;
  assign new_n1245_ = new_n2158_ | new_n2159_;
  assign new_n1246_ = new_n2160_ & new_n2156_;
  assign new_n1247_ = new_n2161_ | new_n2158_;
  assign new_n1248_ = new_n2160_ & new_n2157_;
  assign new_n1249_ = new_n2161_ | new_n2159_;
  assign new_n1250_ = new_n1249_ & new_n1247_;
  assign new_n1251_ = new_n1248_ | new_n1246_;
  assign new_n1252_ = new_n2162_ & new_n2163_;
  assign new_n1253_ = new_n2164_ | new_n2165_;
  assign new_n1254_ = new_n2166_ & new_n2162_;
  assign new_n1255_ = new_n2167_ | new_n2164_;
  assign new_n1256_ = new_n2166_ & new_n2163_;
  assign new_n1257_ = new_n2167_ | new_n2165_;
  assign new_n1258_ = new_n1257_ & new_n1255_;
  assign new_n1259_ = new_n1256_ | new_n1254_;
  assign new_n1260_ = new_n2168_ | new_n2169_;
  assign new_n1261_ = new_n2170_ | new_n2172_;
  assign new_n1262_ = new_n1261_ | new_n2174_;
  assign new_n1263_ = new_n2170_ | new_n2177_;
  assign new_n1264_ = new_n1263_ | new_n2180_;
  assign new_n1265_ = new_n2182_ | new_n2169_;
  assign new_n1266_ = new_n1265_ | new_n2172_;
  assign new_n1267_ = new_n1266_ | new_n2180_;
  assign new_n1268_ = new_n2168_ | new_n2185_;
  assign new_n1269_ = new_n1268_ | new_n2171_;
  assign new_n1270_ = new_n1269_ | new_n2179_;
  assign new_n1271_ = new_n1264_ & new_n1262_;
  assign new_n1272_ = new_n1271_ & new_n1267_;
  assign new_n1273_ = new_n1272_ & new_n1270_;
  assign new_n1274_ = new_n2187_ | new_n2188_;
  assign new_n1275_ = new_n2189_ | new_n2191_;
  assign new_n1276_ = new_n1275_ | new_n2193_;
  assign new_n1277_ = new_n2189_ | new_n2196_;
  assign new_n1278_ = new_n1277_ | new_n2199_;
  assign new_n1279_ = new_n2201_ | new_n2188_;
  assign new_n1280_ = new_n1279_ | new_n2191_;
  assign new_n1281_ = new_n1280_ | new_n2199_;
  assign new_n1282_ = new_n2187_ | new_n2204_;
  assign new_n1283_ = new_n1282_ | new_n2190_;
  assign new_n1284_ = new_n1283_ | new_n2198_;
  assign new_n1285_ = new_n1278_ & new_n1276_;
  assign new_n1286_ = new_n1285_ & new_n1281_;
  assign new_n1287_ = new_n1286_ & new_n1284_;
  assign new_n1288_ = new_n2208_ & new_n614_;
  assign new_n1289_ = new_n2215_ | new_n615_;
  assign new_n1290_ = new_n2221_ & new_n2224_;
  assign new_n1291_ = new_n2227_ | new_n2230_;
  assign new_n1292_ = new_n2232_ & new_n2224_;
  assign new_n1293_ = new_n2233_ | new_n2230_;
  assign new_n1294_ = new_n2232_ & new_n2221_;
  assign new_n1295_ = new_n2233_ | new_n2227_;
  assign new_n1296_ = new_n1295_ & new_n1293_;
  assign new_n1297_ = new_n1294_ | new_n1292_;
  assign new_n1298_ = new_n1297_ & new_n1288_;
  assign new_n1299_ = new_n2234_ | new_n1289_;
  assign new_n1300_ = new_n2234_ | new_n1296_;
  assign new_n1301_ = new_n1300_ & new_n1299_;
  assign new_n1302_ = new_n2208_ & new_n618_;
  assign new_n1303_ = new_n2215_ | new_n619_;
  assign new_n1304_ = new_n2236_ & new_n2239_;
  assign new_n1305_ = new_n2242_ | new_n2245_;
  assign new_n1306_ = new_n2247_ & new_n2239_;
  assign new_n1307_ = new_n2248_ | new_n2245_;
  assign new_n1308_ = new_n2247_ & new_n2236_;
  assign new_n1309_ = new_n2248_ | new_n2242_;
  assign new_n1310_ = new_n1309_ & new_n1307_;
  assign new_n1311_ = new_n1308_ | new_n1306_;
  assign new_n1312_ = new_n1311_ & new_n1302_;
  assign new_n1313_ = new_n2249_ | new_n1303_;
  assign new_n1314_ = new_n2249_ | new_n1310_;
  assign new_n1315_ = new_n1314_ & new_n1313_;
  assign new_n1316_ = new_n2209_ & new_n622_;
  assign new_n1317_ = new_n2216_ | new_n623_;
  assign new_n1318_ = new_n2240_ & new_n2225_;
  assign new_n1319_ = new_n2246_ | new_n2231_;
  assign new_n1320_ = new_n2250_ & new_n2225_;
  assign new_n1321_ = new_n2251_ | new_n2231_;
  assign new_n1322_ = new_n2250_ & new_n2240_;
  assign new_n1323_ = new_n2251_ | new_n2246_;
  assign new_n1324_ = new_n1323_ & new_n1321_;
  assign new_n1325_ = new_n1322_ | new_n1320_;
  assign new_n1326_ = new_n1325_ & new_n1316_;
  assign new_n1327_ = new_n2252_ | new_n1317_;
  assign new_n1328_ = new_n2252_ | new_n1324_;
  assign new_n1329_ = new_n1328_ & new_n1327_;
  assign new_n1330_ = new_n2209_ & new_n626_;
  assign new_n1331_ = new_n2216_ | new_n627_;
  assign new_n1332_ = new_n2237_ & new_n2222_;
  assign new_n1333_ = new_n2243_ | new_n2228_;
  assign new_n1334_ = new_n2253_ & new_n2222_;
  assign new_n1335_ = new_n2254_ | new_n2228_;
  assign new_n1336_ = new_n2253_ & new_n2237_;
  assign new_n1337_ = new_n2254_ | new_n2243_;
  assign new_n1338_ = new_n1337_ & new_n1335_;
  assign new_n1339_ = new_n1336_ | new_n1334_;
  assign new_n1340_ = new_n1339_ & new_n1330_;
  assign new_n1341_ = new_n2255_ | new_n1331_;
  assign new_n1342_ = new_n2255_ | new_n1338_;
  assign new_n1343_ = new_n1342_ & new_n1341_;
  assign new_n1344_ = new_n2211_ & new_n630_;
  assign new_n1345_ = new_n2218_ | new_n631_;
  assign new_n1346_ = new_n2257_ & new_n2260_;
  assign new_n1347_ = new_n2263_ | new_n2266_;
  assign new_n1348_ = new_n2268_ & new_n2260_;
  assign new_n1349_ = new_n2269_ | new_n2266_;
  assign new_n1350_ = new_n2268_ & new_n2257_;
  assign new_n1351_ = new_n2269_ | new_n2263_;
  assign new_n1352_ = new_n1351_ & new_n1349_;
  assign new_n1353_ = new_n1350_ | new_n1348_;
  assign new_n1354_ = new_n1353_ & new_n1344_;
  assign new_n1355_ = new_n2270_ | new_n1345_;
  assign new_n1356_ = new_n2270_ | new_n1352_;
  assign new_n1357_ = new_n1356_ & new_n1355_;
  assign new_n1358_ = new_n2211_ & new_n634_;
  assign new_n1359_ = new_n2218_ | new_n635_;
  assign new_n1360_ = new_n2272_ & new_n2275_;
  assign new_n1361_ = new_n2278_ | new_n2281_;
  assign new_n1362_ = new_n2283_ & new_n2275_;
  assign new_n1363_ = new_n2284_ | new_n2281_;
  assign new_n1364_ = new_n2283_ & new_n2272_;
  assign new_n1365_ = new_n2284_ | new_n2278_;
  assign new_n1366_ = new_n1365_ & new_n1363_;
  assign new_n1367_ = new_n1364_ | new_n1362_;
  assign new_n1368_ = new_n1367_ & new_n1358_;
  assign new_n1369_ = new_n2285_ | new_n1359_;
  assign new_n1370_ = new_n2285_ | new_n1366_;
  assign new_n1371_ = new_n1370_ & new_n1369_;
  assign new_n1372_ = new_n2212_ & new_n638_;
  assign new_n1373_ = new_n2219_ | new_n639_;
  assign new_n1374_ = new_n2276_ & new_n2261_;
  assign new_n1375_ = new_n2282_ | new_n2267_;
  assign new_n1376_ = new_n2286_ & new_n2261_;
  assign new_n1377_ = new_n2287_ | new_n2267_;
  assign new_n1378_ = new_n2286_ & new_n2276_;
  assign new_n1379_ = new_n2287_ | new_n2282_;
  assign new_n1380_ = new_n1379_ & new_n1377_;
  assign new_n1381_ = new_n1378_ | new_n1376_;
  assign new_n1382_ = new_n1381_ & new_n1372_;
  assign new_n1383_ = new_n2288_ | new_n1373_;
  assign new_n1384_ = new_n2288_ | new_n1380_;
  assign new_n1385_ = new_n1384_ & new_n1383_;
  assign new_n1386_ = new_n2212_ & new_n642_;
  assign new_n1387_ = new_n2219_ | new_n643_;
  assign new_n1388_ = new_n2273_ & new_n2258_;
  assign new_n1389_ = new_n2279_ | new_n2264_;
  assign new_n1390_ = new_n2289_ & new_n2258_;
  assign new_n1391_ = new_n2290_ | new_n2264_;
  assign new_n1392_ = new_n2289_ & new_n2273_;
  assign new_n1393_ = new_n2290_ | new_n2279_;
  assign new_n1394_ = new_n1393_ & new_n1391_;
  assign new_n1395_ = new_n1392_ | new_n1390_;
  assign new_n1396_ = new_n1395_ & new_n1386_;
  assign new_n1397_ = new_n2291_ | new_n1387_;
  assign new_n1398_ = new_n2291_ | new_n1394_;
  assign new_n1399_ = new_n1398_ & new_n1397_;
  assign new_n1400_ = new_n2292_ & new_n2293_;
  assign new_n1401_ = new_n2295_ | new_n2297_;
  assign new_n1402_ = new_n2298_ & new_n2293_;
  assign new_n1403_ = new_n2299_ | new_n2297_;
  assign new_n1404_ = new_n2298_ & new_n2292_;
  assign new_n1405_ = new_n2299_ | new_n2295_;
  assign new_n1406_ = new_n1405_ & new_n1403_;
  assign new_n1407_ = new_n1404_ | new_n1402_;
  assign new_n1408_ = new_n2300_ & new_n2301_;
  assign new_n1409_ = new_n2303_ | new_n2305_;
  assign new_n1410_ = new_n2306_ & new_n2301_;
  assign new_n1411_ = new_n2307_ | new_n2305_;
  assign new_n1412_ = new_n2306_ & new_n2300_;
  assign new_n1413_ = new_n2307_ | new_n2303_;
  assign new_n1414_ = new_n1413_ & new_n1411_;
  assign new_n1415_ = new_n1412_ | new_n1410_;
  assign new_n1416_ = new_n1415_ & new_n1407_;
  assign new_n1417_ = new_n2308_ | new_n1406_;
  assign new_n1418_ = new_n2308_ | new_n1414_;
  assign new_n1419_ = new_n1418_ & new_n1417_;
  assign new_n1420_ = new_n2309_ & new_n2310_;
  assign new_n1421_ = new_n2312_ | new_n2314_;
  assign new_n1422_ = new_n2315_ & new_n2310_;
  assign new_n1423_ = new_n2316_ | new_n2314_;
  assign new_n1424_ = new_n2315_ & new_n2309_;
  assign new_n1425_ = new_n2316_ | new_n2312_;
  assign new_n1426_ = new_n1425_ & new_n1423_;
  assign new_n1427_ = new_n1424_ | new_n1422_;
  assign new_n1428_ = new_n2317_ & new_n2318_;
  assign new_n1429_ = new_n2320_ | new_n2322_;
  assign new_n1430_ = new_n2323_ & new_n2318_;
  assign new_n1431_ = new_n2324_ | new_n2322_;
  assign new_n1432_ = new_n2323_ & new_n2317_;
  assign new_n1433_ = new_n2324_ | new_n2320_;
  assign new_n1434_ = new_n1433_ & new_n1431_;
  assign new_n1435_ = new_n1432_ | new_n1430_;
  assign new_n1436_ = new_n1435_ & new_n1427_;
  assign new_n1437_ = new_n2325_ | new_n1426_;
  assign new_n1438_ = new_n2325_ | new_n1434_;
  assign new_n1439_ = new_n1438_ & new_n1437_;
  assign new_n1440_ = new_n2326_ & new_n2327_;
  assign new_n1441_ = new_n2329_ | new_n2331_;
  assign new_n1442_ = new_n2332_ & new_n2327_;
  assign new_n1443_ = new_n2333_ | new_n2331_;
  assign new_n1444_ = new_n2332_ & new_n2326_;
  assign new_n1445_ = new_n2333_ | new_n2329_;
  assign new_n1446_ = new_n1445_ & new_n1443_;
  assign new_n1447_ = new_n1444_ | new_n1442_;
  assign new_n1448_ = new_n2334_ & new_n2335_;
  assign new_n1449_ = new_n2337_ | new_n2339_;
  assign new_n1450_ = new_n2340_ & new_n2335_;
  assign new_n1451_ = new_n2341_ | new_n2339_;
  assign new_n1452_ = new_n2340_ & new_n2334_;
  assign new_n1453_ = new_n2341_ | new_n2337_;
  assign new_n1454_ = new_n1453_ & new_n1451_;
  assign new_n1455_ = new_n1452_ | new_n1450_;
  assign new_n1456_ = new_n1455_ & new_n1447_;
  assign new_n1457_ = new_n2342_ | new_n1446_;
  assign new_n1458_ = new_n2342_ | new_n1454_;
  assign new_n1459_ = new_n1458_ & new_n1457_;
  assign new_n1460_ = new_n2343_ & new_n2344_;
  assign new_n1461_ = new_n2346_ | new_n2348_;
  assign new_n1462_ = new_n2349_ & new_n2344_;
  assign new_n1463_ = new_n2350_ | new_n2348_;
  assign new_n1464_ = new_n2349_ & new_n2343_;
  assign new_n1465_ = new_n2350_ | new_n2346_;
  assign new_n1466_ = new_n1465_ & new_n1463_;
  assign new_n1467_ = new_n1464_ | new_n1462_;
  assign new_n1468_ = new_n2351_ & new_n2352_;
  assign new_n1469_ = new_n2354_ | new_n2356_;
  assign new_n1470_ = new_n2357_ & new_n2352_;
  assign new_n1471_ = new_n2358_ | new_n2356_;
  assign new_n1472_ = new_n2357_ & new_n2351_;
  assign new_n1473_ = new_n2358_ | new_n2354_;
  assign new_n1474_ = new_n1473_ & new_n1471_;
  assign new_n1475_ = new_n1472_ | new_n1470_;
  assign new_n1476_ = new_n1475_ & new_n1467_;
  assign new_n1477_ = new_n2359_ | new_n1466_;
  assign new_n1478_ = new_n2359_ | new_n1474_;
  assign new_n1479_ = new_n1478_ & new_n1477_;
  assign new_n1480_ = new_n2360_ & new_n2361_;
  assign new_n1481_ = new_n2363_ | new_n2365_;
  assign new_n1482_ = new_n2366_ & new_n2361_;
  assign new_n1483_ = new_n2367_ | new_n2365_;
  assign new_n1484_ = new_n2366_ & new_n2360_;
  assign new_n1485_ = new_n2367_ | new_n2363_;
  assign new_n1486_ = new_n1485_ & new_n1483_;
  assign new_n1487_ = new_n1484_ | new_n1482_;
  assign new_n1488_ = new_n2368_ & new_n2369_;
  assign new_n1489_ = new_n2371_ | new_n2373_;
  assign new_n1490_ = new_n2374_ & new_n2369_;
  assign new_n1491_ = new_n2375_ | new_n2373_;
  assign new_n1492_ = new_n2374_ & new_n2368_;
  assign new_n1493_ = new_n2375_ | new_n2371_;
  assign new_n1494_ = new_n1493_ & new_n1491_;
  assign new_n1495_ = new_n1492_ | new_n1490_;
  assign new_n1496_ = new_n1495_ & new_n1487_;
  assign new_n1497_ = new_n2376_ | new_n1486_;
  assign new_n1498_ = new_n2376_ | new_n1494_;
  assign new_n1499_ = new_n1498_ & new_n1497_;
  assign new_n1500_ = new_n2377_ & new_n2378_;
  assign new_n1501_ = new_n2380_ | new_n2382_;
  assign new_n1502_ = new_n2383_ & new_n2378_;
  assign new_n1503_ = new_n2384_ | new_n2382_;
  assign new_n1504_ = new_n2383_ & new_n2377_;
  assign new_n1505_ = new_n2384_ | new_n2380_;
  assign new_n1506_ = new_n1505_ & new_n1503_;
  assign new_n1507_ = new_n1504_ | new_n1502_;
  assign new_n1508_ = new_n2385_ & new_n2386_;
  assign new_n1509_ = new_n2388_ | new_n2390_;
  assign new_n1510_ = new_n2391_ & new_n2386_;
  assign new_n1511_ = new_n2392_ | new_n2390_;
  assign new_n1512_ = new_n2391_ & new_n2385_;
  assign new_n1513_ = new_n2392_ | new_n2388_;
  assign new_n1514_ = new_n1513_ & new_n1511_;
  assign new_n1515_ = new_n1512_ | new_n1510_;
  assign new_n1516_ = new_n1515_ & new_n1507_;
  assign new_n1517_ = new_n2393_ | new_n1506_;
  assign new_n1518_ = new_n2393_ | new_n1514_;
  assign new_n1519_ = new_n1518_ & new_n1517_;
  assign new_n1520_ = new_n2394_ & new_n2395_;
  assign new_n1521_ = new_n2397_ | new_n2399_;
  assign new_n1522_ = new_n2400_ & new_n2395_;
  assign new_n1523_ = new_n2401_ | new_n2399_;
  assign new_n1524_ = new_n2400_ & new_n2394_;
  assign new_n1525_ = new_n2401_ | new_n2397_;
  assign new_n1526_ = new_n1525_ & new_n1523_;
  assign new_n1527_ = new_n1524_ | new_n1522_;
  assign new_n1528_ = new_n2402_ & new_n2403_;
  assign new_n1529_ = new_n2405_ | new_n2407_;
  assign new_n1530_ = new_n2408_ & new_n2403_;
  assign new_n1531_ = new_n2409_ | new_n2407_;
  assign new_n1532_ = new_n2408_ & new_n2402_;
  assign new_n1533_ = new_n2409_ | new_n2405_;
  assign new_n1534_ = new_n1533_ & new_n1531_;
  assign new_n1535_ = new_n1532_ | new_n1530_;
  assign new_n1536_ = new_n1535_ & new_n1527_;
  assign new_n1537_ = new_n2410_ | new_n1526_;
  assign new_n1538_ = new_n2410_ | new_n1534_;
  assign new_n1539_ = new_n1538_ & new_n1537_;
  assign new_n1540_ = new_n2411_ & new_n2412_;
  assign new_n1541_ = new_n2414_ | new_n2416_;
  assign new_n1542_ = new_n2417_ & new_n2412_;
  assign new_n1543_ = new_n2418_ | new_n2416_;
  assign new_n1544_ = new_n2417_ & new_n2411_;
  assign new_n1545_ = new_n2418_ | new_n2414_;
  assign new_n1546_ = new_n1545_ & new_n1543_;
  assign new_n1547_ = new_n1544_ | new_n1542_;
  assign new_n1548_ = new_n2419_ & new_n2420_;
  assign new_n1549_ = new_n2422_ | new_n2424_;
  assign new_n1550_ = new_n2425_ & new_n2420_;
  assign new_n1551_ = new_n2426_ | new_n2424_;
  assign new_n1552_ = new_n2425_ & new_n2419_;
  assign new_n1553_ = new_n2426_ | new_n2422_;
  assign new_n1554_ = new_n1553_ & new_n1551_;
  assign new_n1555_ = new_n1552_ | new_n1550_;
  assign new_n1556_ = new_n1555_ & new_n1547_;
  assign new_n1557_ = new_n2427_ | new_n1546_;
  assign new_n1558_ = new_n2427_ | new_n1554_;
  assign new_n1559_ = new_n1558_ & new_n1557_;
  assign new_n1560_ = new_n2428_ & new_n2429_;
  assign new_n1561_ = new_n2431_ | new_n2433_;
  assign new_n1562_ = new_n2434_ & new_n2429_;
  assign new_n1563_ = new_n2435_ | new_n2433_;
  assign new_n1564_ = new_n2434_ & new_n2428_;
  assign new_n1565_ = new_n2435_ | new_n2431_;
  assign new_n1566_ = new_n1565_ & new_n1563_;
  assign new_n1567_ = new_n1564_ | new_n1562_;
  assign new_n1568_ = new_n2436_ & new_n2437_;
  assign new_n1569_ = new_n2439_ | new_n2441_;
  assign new_n1570_ = new_n2442_ & new_n2437_;
  assign new_n1571_ = new_n2443_ | new_n2441_;
  assign new_n1572_ = new_n2442_ & new_n2436_;
  assign new_n1573_ = new_n2443_ | new_n2439_;
  assign new_n1574_ = new_n1573_ & new_n1571_;
  assign new_n1575_ = new_n1572_ | new_n1570_;
  assign new_n1576_ = new_n1575_ & new_n1567_;
  assign new_n1577_ = new_n2444_ | new_n1566_;
  assign new_n1578_ = new_n2444_ | new_n1574_;
  assign new_n1579_ = new_n1578_ & new_n1577_;
  assign new_n1580_ = new_n2445_ & new_n2446_;
  assign new_n1581_ = new_n2448_ | new_n2450_;
  assign new_n1582_ = new_n2451_ & new_n2446_;
  assign new_n1583_ = new_n2452_ | new_n2450_;
  assign new_n1584_ = new_n2451_ & new_n2445_;
  assign new_n1585_ = new_n2452_ | new_n2448_;
  assign new_n1586_ = new_n1585_ & new_n1583_;
  assign new_n1587_ = new_n1584_ | new_n1582_;
  assign new_n1588_ = new_n2453_ & new_n2454_;
  assign new_n1589_ = new_n2456_ | new_n2458_;
  assign new_n1590_ = new_n2459_ & new_n2454_;
  assign new_n1591_ = new_n2460_ | new_n2458_;
  assign new_n1592_ = new_n2459_ & new_n2453_;
  assign new_n1593_ = new_n2460_ | new_n2456_;
  assign new_n1594_ = new_n1593_ & new_n1591_;
  assign new_n1595_ = new_n1592_ | new_n1590_;
  assign new_n1596_ = new_n1595_ & new_n1587_;
  assign new_n1597_ = new_n2461_ | new_n1586_;
  assign new_n1598_ = new_n2461_ | new_n1594_;
  assign new_n1599_ = new_n1598_ & new_n1597_;
  assign new_n1600_ = new_n2462_ & new_n2463_;
  assign new_n1601_ = new_n2465_ | new_n2467_;
  assign new_n1602_ = new_n2468_ & new_n2463_;
  assign new_n1603_ = new_n2469_ | new_n2467_;
  assign new_n1604_ = new_n2468_ & new_n2462_;
  assign new_n1605_ = new_n2469_ | new_n2465_;
  assign new_n1606_ = new_n1605_ & new_n1603_;
  assign new_n1607_ = new_n1604_ | new_n1602_;
  assign new_n1608_ = new_n2470_ & new_n2471_;
  assign new_n1609_ = new_n2473_ | new_n2475_;
  assign new_n1610_ = new_n2476_ & new_n2471_;
  assign new_n1611_ = new_n2477_ | new_n2475_;
  assign new_n1612_ = new_n2476_ & new_n2470_;
  assign new_n1613_ = new_n2477_ | new_n2473_;
  assign new_n1614_ = new_n1613_ & new_n1611_;
  assign new_n1615_ = new_n1612_ | new_n1610_;
  assign new_n1616_ = new_n1615_ & new_n1607_;
  assign new_n1617_ = new_n2478_ | new_n1606_;
  assign new_n1618_ = new_n2478_ | new_n1614_;
  assign new_n1619_ = new_n1618_ & new_n1617_;
  assign new_n1620_ = new_n2479_ & new_n2480_;
  assign new_n1621_ = new_n2482_ | new_n2484_;
  assign new_n1622_ = new_n2485_ & new_n2480_;
  assign new_n1623_ = new_n2486_ | new_n2484_;
  assign new_n1624_ = new_n2485_ & new_n2479_;
  assign new_n1625_ = new_n2486_ | new_n2482_;
  assign new_n1626_ = new_n1625_ & new_n1623_;
  assign new_n1627_ = new_n1624_ | new_n1622_;
  assign new_n1628_ = new_n2487_ & new_n2488_;
  assign new_n1629_ = new_n2490_ | new_n2492_;
  assign new_n1630_ = new_n2493_ & new_n2488_;
  assign new_n1631_ = new_n2494_ | new_n2492_;
  assign new_n1632_ = new_n2493_ & new_n2487_;
  assign new_n1633_ = new_n2494_ | new_n2490_;
  assign new_n1634_ = new_n1633_ & new_n1631_;
  assign new_n1635_ = new_n1632_ | new_n1630_;
  assign new_n1636_ = new_n1635_ & new_n1627_;
  assign new_n1637_ = new_n2495_ | new_n1626_;
  assign new_n1638_ = new_n2495_ | new_n1634_;
  assign new_n1639_ = new_n1638_ & new_n1637_;
  assign new_n1640_ = new_n2496_ & new_n2497_;
  assign new_n1641_ = new_n2499_ | new_n2501_;
  assign new_n1642_ = new_n2502_ & new_n2497_;
  assign new_n1643_ = new_n2503_ | new_n2501_;
  assign new_n1644_ = new_n2502_ & new_n2496_;
  assign new_n1645_ = new_n2503_ | new_n2499_;
  assign new_n1646_ = new_n1645_ & new_n1643_;
  assign new_n1647_ = new_n1644_ | new_n1642_;
  assign new_n1648_ = new_n2504_ & new_n2505_;
  assign new_n1649_ = new_n2507_ | new_n2509_;
  assign new_n1650_ = new_n2510_ & new_n2505_;
  assign new_n1651_ = new_n2511_ | new_n2509_;
  assign new_n1652_ = new_n2510_ & new_n2504_;
  assign new_n1653_ = new_n2511_ | new_n2507_;
  assign new_n1654_ = new_n1653_ & new_n1651_;
  assign new_n1655_ = new_n1652_ | new_n1650_;
  assign new_n1656_ = new_n1655_ & new_n1647_;
  assign new_n1657_ = new_n2512_ | new_n1646_;
  assign new_n1658_ = new_n2512_ | new_n1654_;
  assign new_n1659_ = new_n1658_ & new_n1657_;
  assign new_n1660_ = new_n2513_ & new_n2514_;
  assign new_n1661_ = new_n2516_ | new_n2518_;
  assign new_n1662_ = new_n2519_ & new_n2514_;
  assign new_n1663_ = new_n2520_ | new_n2518_;
  assign new_n1664_ = new_n2519_ & new_n2513_;
  assign new_n1665_ = new_n2520_ | new_n2516_;
  assign new_n1666_ = new_n1665_ & new_n1663_;
  assign new_n1667_ = new_n1664_ | new_n1662_;
  assign new_n1668_ = new_n2521_ & new_n2522_;
  assign new_n1669_ = new_n2524_ | new_n2526_;
  assign new_n1670_ = new_n2527_ & new_n2522_;
  assign new_n1671_ = new_n2528_ | new_n2526_;
  assign new_n1672_ = new_n2527_ & new_n2521_;
  assign new_n1673_ = new_n2528_ | new_n2524_;
  assign new_n1674_ = new_n1673_ & new_n1671_;
  assign new_n1675_ = new_n1672_ | new_n1670_;
  assign new_n1676_ = new_n1675_ & new_n1667_;
  assign new_n1677_ = new_n2529_ | new_n1666_;
  assign new_n1678_ = new_n2529_ | new_n1674_;
  assign new_n1679_ = new_n1678_ & new_n1677_;
  assign new_n1680_ = new_n2530_ & new_n2531_;
  assign new_n1681_ = new_n2533_ | new_n2535_;
  assign new_n1682_ = new_n2536_ & new_n2531_;
  assign new_n1683_ = new_n2537_ | new_n2535_;
  assign new_n1684_ = new_n2536_ & new_n2530_;
  assign new_n1685_ = new_n2537_ | new_n2533_;
  assign new_n1686_ = new_n1685_ & new_n1683_;
  assign new_n1687_ = new_n1684_ | new_n1682_;
  assign new_n1688_ = new_n2538_ & new_n2539_;
  assign new_n1689_ = new_n2541_ | new_n2543_;
  assign new_n1690_ = new_n2544_ & new_n2539_;
  assign new_n1691_ = new_n2545_ | new_n2543_;
  assign new_n1692_ = new_n2544_ & new_n2538_;
  assign new_n1693_ = new_n2545_ | new_n2541_;
  assign new_n1694_ = new_n1693_ & new_n1691_;
  assign new_n1695_ = new_n1692_ | new_n1690_;
  assign new_n1696_ = new_n1695_ & new_n1687_;
  assign new_n1697_ = new_n2546_ | new_n1686_;
  assign new_n1698_ = new_n2546_ | new_n1694_;
  assign new_n1699_ = new_n1698_ & new_n1697_;
  assign new_n1700_ = new_n2547_ & new_n2548_;
  assign new_n1701_ = new_n2550_ | new_n2552_;
  assign new_n1702_ = new_n2553_ & new_n2548_;
  assign new_n1703_ = new_n2554_ | new_n2552_;
  assign new_n1704_ = new_n2553_ & new_n2547_;
  assign new_n1705_ = new_n2554_ | new_n2550_;
  assign new_n1706_ = new_n1705_ & new_n1703_;
  assign new_n1707_ = new_n1704_ | new_n1702_;
  assign new_n1708_ = new_n2555_ & new_n2556_;
  assign new_n1709_ = new_n2558_ | new_n2560_;
  assign new_n1710_ = new_n2561_ & new_n2556_;
  assign new_n1711_ = new_n2562_ | new_n2560_;
  assign new_n1712_ = new_n2561_ & new_n2555_;
  assign new_n1713_ = new_n2562_ | new_n2558_;
  assign new_n1714_ = new_n1713_ & new_n1711_;
  assign new_n1715_ = new_n1712_ | new_n1710_;
  assign new_n1716_ = new_n1715_ & new_n1707_;
  assign new_n1717_ = new_n2563_ | new_n1706_;
  assign new_n1718_ = new_n2563_ | new_n1714_;
  assign new_n1719_ = new_n1718_ & new_n1717_;
  assign G1324 = ~new_n953_;
  assign G1325 = ~new_n959_;
  assign G1326 = ~new_n965_;
  assign G1327 = ~new_n971_;
  assign G1328 = ~new_n985_;
  assign G1329 = ~new_n991_;
  assign G1330 = ~new_n997_;
  assign G1331 = ~new_n1003_;
  assign G1332 = ~new_n1017_;
  assign G1333 = ~new_n1023_;
  assign G1334 = ~new_n1029_;
  assign G1335 = ~new_n1035_;
  assign G1336 = ~new_n1049_;
  assign G1337 = ~new_n1055_;
  assign G1338 = ~new_n1061_;
  assign G1339 = ~new_n1067_;
  assign G1340 = ~new_n1081_;
  assign G1341 = ~new_n1087_;
  assign G1342 = ~new_n1093_;
  assign G1343 = ~new_n1099_;
  assign G1344 = ~new_n1113_;
  assign G1345 = ~new_n1119_;
  assign G1346 = ~new_n1125_;
  assign G1347 = ~new_n1131_;
  assign G1348 = ~new_n1145_;
  assign G1349 = ~new_n1151_;
  assign G1350 = ~new_n1157_;
  assign G1351 = ~new_n1163_;
  assign G1352 = ~new_n1177_;
  assign G1353 = ~new_n1183_;
  assign G1354 = ~new_n1189_;
  assign G1355 = ~new_n1195_;
  assign n630_li = ~new_n649_;
  assign n642_li = ~new_n651_;
  assign n654_li = ~new_n653_;
  assign n666_li = ~new_n655_;
  assign n678_li = ~new_n657_;
  assign n690_li = ~new_n659_;
  assign n702_li = ~new_n661_;
  assign n714_li = ~new_n663_;
  assign n726_li = ~new_n665_;
  assign n738_li = ~new_n667_;
  assign n750_li = ~new_n669_;
  assign n762_li = ~new_n671_;
  assign n774_li = ~new_n673_;
  assign n786_li = ~new_n675_;
  assign n798_li = ~new_n677_;
  assign n810_li = ~new_n679_;
  assign n822_li = ~new_n681_;
  assign n834_li = ~new_n683_;
  assign n846_li = ~new_n685_;
  assign n858_li = ~new_n687_;
  assign n870_li = ~new_n689_;
  assign n882_li = ~new_n691_;
  assign n894_li = ~new_n693_;
  assign n906_li = ~new_n695_;
  assign n918_li = ~new_n697_;
  assign n930_li = ~new_n699_;
  assign n942_li = ~new_n701_;
  assign n954_li = ~new_n703_;
  assign n966_li = ~new_n705_;
  assign n978_li = ~new_n707_;
  assign n990_li = ~new_n709_;
  assign n1002_li = ~new_n711_;
  assign n1005_li = ~new_n531_;
  assign n1008_li = ~new_n613_;
  assign n1017_li = ~new_n533_;
  assign n1020_li = ~new_n617_;
  assign n1029_li = ~new_n535_;
  assign n1032_li = ~new_n621_;
  assign n1041_li = ~new_n537_;
  assign n1044_li = ~new_n625_;
  assign n1053_li = ~new_n539_;
  assign n1056_li = ~new_n629_;
  assign n1065_li = ~new_n541_;
  assign n1068_li = ~new_n633_;
  assign n1077_li = ~new_n543_;
  assign n1080_li = ~new_n637_;
  assign n1089_li = ~new_n545_;
  assign n1092_li = ~new_n641_;
  assign n1101_li = ~new_n547_;
  assign n1104_li = ~new_n645_;
  assign n1837_i2 = ~new_n2296_;
  assign n1838_i2 = ~new_n2313_;
  assign n1839_i2 = ~new_n2330_;
  assign n1840_i2 = ~new_n2347_;
  assign n1841_i2 = ~new_n2294_;
  assign n1842_i2 = ~new_n2311_;
  assign n1843_i2 = ~new_n2328_;
  assign n1844_i2 = ~new_n2345_;
  assign n1845_i2 = ~new_n2304_;
  assign n1846_i2 = ~new_n2321_;
  assign n1847_i2 = ~new_n2338_;
  assign n1848_i2 = ~new_n2355_;
  assign n1849_i2 = ~new_n2302_;
  assign n1850_i2 = ~new_n2319_;
  assign n1851_i2 = ~new_n2336_;
  assign n1852_i2 = ~new_n2353_;
  assign n1853_i2 = ~new_n2364_;
  assign n1854_i2 = ~new_n2381_;
  assign n1855_i2 = ~new_n2398_;
  assign n1856_i2 = ~new_n2415_;
  assign n1857_i2 = ~new_n2362_;
  assign n1858_i2 = ~new_n2379_;
  assign n1859_i2 = ~new_n2396_;
  assign n1860_i2 = ~new_n2413_;
  assign n1861_i2 = ~new_n2372_;
  assign n1862_i2 = ~new_n2389_;
  assign n1863_i2 = ~new_n2406_;
  assign n1864_i2 = ~new_n2423_;
  assign n1865_i2 = ~new_n2370_;
  assign n1866_i2 = ~new_n2387_;
  assign n1867_i2 = ~new_n2404_;
  assign n1868_i2 = ~new_n2421_;
  assign G834_i2 = ~new_n2185_;
  assign G847_i2 = ~new_n2182_;
  assign G860_i2 = ~new_n2177_;
  assign G873_i2 = ~new_n2174_;
  assign G925_i2 = ~new_n2204_;
  assign G886_i2 = ~new_n2201_;
  assign G912_i2 = ~new_n2196_;
  assign G899_i2 = ~new_n2193_;
  assign n2151_i2 = ~new_n2432_;
  assign n2152_i2 = ~new_n2430_;
  assign n2153_i2 = ~new_n2440_;
  assign n2154_i2 = ~new_n2438_;
  assign n2155_i2 = ~new_n2449_;
  assign n2156_i2 = ~new_n2447_;
  assign n2157_i2 = ~new_n2457_;
  assign n2158_i2 = ~new_n2455_;
  assign n2159_i2 = ~new_n2466_;
  assign n2160_i2 = ~new_n2464_;
  assign n2161_i2 = ~new_n2474_;
  assign n2162_i2 = ~new_n2472_;
  assign n2163_i2 = ~new_n2483_;
  assign n2164_i2 = ~new_n2481_;
  assign n2165_i2 = ~new_n2491_;
  assign n2166_i2 = ~new_n2489_;
  assign n2167_i2 = ~new_n2500_;
  assign n2168_i2 = ~new_n2498_;
  assign n2169_i2 = ~new_n2508_;
  assign n2170_i2 = ~new_n2506_;
  assign n2171_i2 = ~new_n2517_;
  assign n2172_i2 = ~new_n2515_;
  assign n2173_i2 = ~new_n2525_;
  assign n2174_i2 = ~new_n2523_;
  assign n2175_i2 = ~new_n2534_;
  assign n2176_i2 = ~new_n2532_;
  assign n2177_i2 = ~new_n2542_;
  assign n2178_i2 = ~new_n2540_;
  assign n2179_i2 = ~new_n2551_;
  assign n2180_i2 = ~new_n2549_;
  assign n2181_i2 = ~new_n2559_;
  assign n2182_i2 = ~new_n2557_;
  assign G974_i2 = ~new_n2186_;
  assign G976_i2 = G974_i2;
  assign G970_i2 = ~new_n2183_;
  assign G972_i2 = G970_i2;
  assign G973_i2 = ~new_n2178_;
  assign G977_i2 = G973_i2;
  assign G971_i2 = ~new_n2175_;
  assign G975_i2 = G971_i2;
  assign G954_i2 = ~new_n2205_;
  assign G956_i2 = G954_i2;
  assign G950_i2 = ~new_n2202_;
  assign G952_i2 = G950_i2;
  assign G953_i2 = ~new_n2197_;
  assign G957_i2 = G953_i2;
  assign G951_i2 = ~new_n2194_;
  assign G955_i2 = G951_i2;
  assign G986_i2 = ~new_n1273_;
  assign G991_i2 = ~new_n1287_;
  assign G770_i2 = ~new_n1301_;
  assign G773_i2 = ~new_n1315_;
  assign G776_i2 = ~new_n1329_;
  assign G779_i2 = ~new_n1343_;
  assign G782_i2 = ~new_n1357_;
  assign G785_i2 = ~new_n1371_;
  assign G788_i2 = ~new_n1385_;
  assign G791_i2 = ~new_n1399_;
  assign G642_i2 = ~new_n1419_;
  assign G645_i2 = ~new_n1439_;
  assign G648_i2 = ~new_n1459_;
  assign G651_i2 = ~new_n1479_;
  assign G654_i2 = ~new_n1499_;
  assign G657_i2 = ~new_n1519_;
  assign G660_i2 = ~new_n1539_;
  assign G663_i2 = ~new_n1559_;
  assign G602_i2 = ~new_n1579_;
  assign G607_i2 = ~new_n1599_;
  assign G612_i2 = ~new_n1619_;
  assign G617_i2 = ~new_n1639_;
  assign G622_i2 = ~new_n1659_;
  assign G627_i2 = ~new_n1679_;
  assign G632_i2 = ~new_n1699_;
  assign G637_i2 = ~new_n1719_;
  assign n627_lo_buf_i2 = ~new_n467_;
  assign n639_lo_buf_i2 = ~new_n469_;
  assign n651_lo_buf_i2 = ~new_n471_;
  assign n663_lo_buf_i2 = ~new_n473_;
  assign n675_lo_buf_i2 = ~new_n475_;
  assign n687_lo_buf_i2 = ~new_n477_;
  assign n699_lo_buf_i2 = ~new_n479_;
  assign n711_lo_buf_i2 = ~new_n481_;
  assign n723_lo_buf_i2 = ~new_n483_;
  assign n735_lo_buf_i2 = ~new_n485_;
  assign n747_lo_buf_i2 = ~new_n487_;
  assign n759_lo_buf_i2 = ~new_n489_;
  assign n771_lo_buf_i2 = ~new_n491_;
  assign n783_lo_buf_i2 = ~new_n493_;
  assign n795_lo_buf_i2 = ~new_n495_;
  assign n807_lo_buf_i2 = ~new_n497_;
  assign n819_lo_buf_i2 = ~new_n499_;
  assign n831_lo_buf_i2 = ~new_n501_;
  assign n843_lo_buf_i2 = ~new_n503_;
  assign n855_lo_buf_i2 = ~new_n505_;
  assign n867_lo_buf_i2 = ~new_n507_;
  assign n879_lo_buf_i2 = ~new_n509_;
  assign n891_lo_buf_i2 = ~new_n511_;
  assign n903_lo_buf_i2 = ~new_n513_;
  assign n915_lo_buf_i2 = ~new_n515_;
  assign n927_lo_buf_i2 = ~new_n517_;
  assign n939_lo_buf_i2 = ~new_n519_;
  assign n951_lo_buf_i2 = ~new_n521_;
  assign n963_lo_buf_i2 = ~new_n523_;
  assign n975_lo_buf_i2 = ~new_n525_;
  assign n987_lo_buf_i2 = ~new_n527_;
  assign n999_lo_buf_i2 = ~new_n529_;
  assign new_n1948_ = new_n720_;
  assign new_n1949_ = new_n1948_;
  assign new_n1950_ = new_n1949_;
  assign new_n1951_ = new_n1949_;
  assign new_n1952_ = new_n1948_;
  assign new_n1953_ = new_n721_;
  assign new_n1954_ = new_n1953_;
  assign new_n1955_ = new_n1954_;
  assign new_n1956_ = new_n1954_;
  assign new_n1957_ = new_n1953_;
  assign new_n1958_ = new_n724_;
  assign new_n1959_ = new_n1958_;
  assign new_n1960_ = new_n1959_;
  assign new_n1961_ = new_n1959_;
  assign new_n1962_ = new_n1958_;
  assign new_n1963_ = new_n725_;
  assign new_n1964_ = new_n1963_;
  assign new_n1965_ = new_n1964_;
  assign new_n1966_ = new_n1964_;
  assign new_n1967_ = new_n1963_;
  assign new_n1968_ = new_n824_;
  assign new_n1969_ = new_n1968_;
  assign new_n1970_ = new_n1968_;
  assign new_n1971_ = new_n825_;
  assign new_n1972_ = new_n1971_;
  assign new_n1973_ = new_n1971_;
  assign new_n1974_ = new_n946_;
  assign new_n1975_ = new_n1974_;
  assign new_n1976_ = new_n1974_;
  assign new_n1977_ = new_n712_;
  assign new_n1978_ = new_n1977_;
  assign new_n1979_ = new_n1978_;
  assign new_n1980_ = new_n1978_;
  assign new_n1981_ = new_n1977_;
  assign new_n1982_ = new_n947_;
  assign new_n1983_ = new_n1982_;
  assign new_n1984_ = new_n1982_;
  assign new_n1985_ = new_n713_;
  assign new_n1986_ = new_n1985_;
  assign new_n1987_ = new_n1986_;
  assign new_n1988_ = new_n1986_;
  assign new_n1989_ = new_n1985_;
  assign new_n1990_ = new_n950_;
  assign new_n1991_ = new_n714_;
  assign new_n1992_ = new_n1991_;
  assign new_n1993_ = new_n1992_;
  assign new_n1994_ = new_n1992_;
  assign new_n1995_ = new_n1991_;
  assign new_n1996_ = new_n715_;
  assign new_n1997_ = new_n1996_;
  assign new_n1998_ = new_n1997_;
  assign new_n1999_ = new_n1997_;
  assign new_n2000_ = new_n1996_;
  assign new_n2001_ = new_n956_;
  assign new_n2002_ = new_n716_;
  assign new_n2003_ = new_n2002_;
  assign new_n2004_ = new_n2003_;
  assign new_n2005_ = new_n2003_;
  assign new_n2006_ = new_n2002_;
  assign new_n2007_ = new_n717_;
  assign new_n2008_ = new_n2007_;
  assign new_n2009_ = new_n2008_;
  assign new_n2010_ = new_n2008_;
  assign new_n2011_ = new_n2007_;
  assign new_n2012_ = new_n962_;
  assign new_n2013_ = new_n718_;
  assign new_n2014_ = new_n2013_;
  assign new_n2015_ = new_n2014_;
  assign new_n2016_ = new_n2014_;
  assign new_n2017_ = new_n2013_;
  assign new_n2018_ = new_n719_;
  assign new_n2019_ = new_n2018_;
  assign new_n2020_ = new_n2019_;
  assign new_n2021_ = new_n2019_;
  assign new_n2022_ = new_n2018_;
  assign new_n2023_ = new_n968_;
  assign new_n2024_ = new_n726_;
  assign new_n2025_ = new_n2024_;
  assign new_n2026_ = new_n2025_;
  assign new_n2027_ = new_n2025_;
  assign new_n2028_ = new_n2024_;
  assign new_n2029_ = new_n727_;
  assign new_n2030_ = new_n2029_;
  assign new_n2031_ = new_n2030_;
  assign new_n2032_ = new_n2030_;
  assign new_n2033_ = new_n2029_;
  assign new_n2034_ = new_n978_;
  assign new_n2035_ = new_n2034_;
  assign new_n2036_ = new_n2034_;
  assign new_n2037_ = new_n979_;
  assign new_n2038_ = new_n2037_;
  assign new_n2039_ = new_n2037_;
  assign new_n2040_ = new_n982_;
  assign new_n2041_ = new_n988_;
  assign new_n2042_ = new_n994_;
  assign new_n2043_ = new_n1000_;
  assign new_n2044_ = new_n722_;
  assign new_n2045_ = new_n2044_;
  assign new_n2046_ = new_n2045_;
  assign new_n2047_ = new_n2045_;
  assign new_n2048_ = new_n2044_;
  assign new_n2049_ = new_n723_;
  assign new_n2050_ = new_n2049_;
  assign new_n2051_ = new_n2050_;
  assign new_n2052_ = new_n2050_;
  assign new_n2053_ = new_n2049_;
  assign new_n2054_ = new_n1010_;
  assign new_n2055_ = new_n2054_;
  assign new_n2056_ = new_n2054_;
  assign new_n2057_ = new_n1011_;
  assign new_n2058_ = new_n2057_;
  assign new_n2059_ = new_n2057_;
  assign new_n2060_ = new_n1014_;
  assign new_n2061_ = new_n1020_;
  assign new_n2062_ = new_n1026_;
  assign new_n2063_ = new_n1032_;
  assign new_n2064_ = new_n1042_;
  assign new_n2065_ = new_n2064_;
  assign new_n2066_ = new_n2064_;
  assign new_n2067_ = new_n1043_;
  assign new_n2068_ = new_n2067_;
  assign new_n2069_ = new_n2067_;
  assign new_n2070_ = new_n1046_;
  assign new_n2071_ = new_n1052_;
  assign new_n2072_ = new_n1058_;
  assign new_n2073_ = new_n1064_;
  assign new_n2074_ = new_n826_;
  assign new_n2075_ = new_n2074_;
  assign new_n2076_ = new_n2074_;
  assign new_n2077_ = new_n827_;
  assign new_n2078_ = new_n2077_;
  assign new_n2079_ = new_n2077_;
  assign new_n2080_ = new_n1074_;
  assign new_n2081_ = new_n2080_;
  assign new_n2082_ = new_n2080_;
  assign new_n2083_ = new_n1075_;
  assign new_n2084_ = new_n2083_;
  assign new_n2085_ = new_n2083_;
  assign new_n2086_ = new_n1078_;
  assign new_n2087_ = new_n1084_;
  assign new_n2088_ = new_n1090_;
  assign new_n2089_ = new_n1096_;
  assign new_n2090_ = new_n1106_;
  assign new_n2091_ = new_n2090_;
  assign new_n2092_ = new_n2090_;
  assign new_n2093_ = new_n1107_;
  assign new_n2094_ = new_n2093_;
  assign new_n2095_ = new_n2093_;
  assign new_n2096_ = new_n1110_;
  assign new_n2097_ = new_n1116_;
  assign new_n2098_ = new_n1122_;
  assign new_n2099_ = new_n1128_;
  assign new_n2100_ = new_n1138_;
  assign new_n2101_ = new_n2100_;
  assign new_n2102_ = new_n2100_;
  assign new_n2103_ = new_n1139_;
  assign new_n2104_ = new_n2103_;
  assign new_n2105_ = new_n2103_;
  assign new_n2106_ = new_n1142_;
  assign new_n2107_ = new_n1148_;
  assign new_n2108_ = new_n1154_;
  assign new_n2109_ = new_n1160_;
  assign new_n2110_ = new_n1170_;
  assign new_n2111_ = new_n2110_;
  assign new_n2112_ = new_n2110_;
  assign new_n2113_ = new_n1171_;
  assign new_n2114_ = new_n2113_;
  assign new_n2115_ = new_n2113_;
  assign new_n2116_ = new_n1174_;
  assign new_n2117_ = new_n1180_;
  assign new_n2118_ = new_n1186_;
  assign new_n2119_ = new_n1192_;
  assign new_n2120_ = new_n844_;
  assign new_n2121_ = new_n828_;
  assign new_n2122_ = new_n845_;
  assign new_n2123_ = new_n829_;
  assign new_n2124_ = new_n1197_;
  assign new_n2125_ = new_n1196_;
  assign new_n2126_ = new_n846_;
  assign new_n2127_ = new_n830_;
  assign new_n2128_ = new_n847_;
  assign new_n2129_ = new_n831_;
  assign new_n2130_ = new_n1205_;
  assign new_n2131_ = new_n1204_;
  assign new_n2132_ = new_n848_;
  assign new_n2133_ = new_n832_;
  assign new_n2134_ = new_n849_;
  assign new_n2135_ = new_n833_;
  assign new_n2136_ = new_n1213_;
  assign new_n2137_ = new_n1212_;
  assign new_n2138_ = new_n850_;
  assign new_n2139_ = new_n834_;
  assign new_n2140_ = new_n851_;
  assign new_n2141_ = new_n835_;
  assign new_n2142_ = new_n1221_;
  assign new_n2143_ = new_n1220_;
  assign new_n2144_ = new_n852_;
  assign new_n2145_ = new_n836_;
  assign new_n2146_ = new_n853_;
  assign new_n2147_ = new_n837_;
  assign new_n2148_ = new_n1229_;
  assign new_n2149_ = new_n1228_;
  assign new_n2150_ = new_n854_;
  assign new_n2151_ = new_n838_;
  assign new_n2152_ = new_n855_;
  assign new_n2153_ = new_n839_;
  assign new_n2154_ = new_n1237_;
  assign new_n2155_ = new_n1236_;
  assign new_n2156_ = new_n856_;
  assign new_n2157_ = new_n840_;
  assign new_n2158_ = new_n857_;
  assign new_n2159_ = new_n841_;
  assign new_n2160_ = new_n1245_;
  assign new_n2161_ = new_n1244_;
  assign new_n2162_ = new_n858_;
  assign new_n2163_ = new_n842_;
  assign new_n2164_ = new_n859_;
  assign new_n2165_ = new_n843_;
  assign new_n2166_ = new_n1253_;
  assign new_n2167_ = new_n1252_;
  assign new_n2168_ = new_n1211_;
  assign new_n2169_ = new_n1203_;
  assign new_n2170_ = new_n1260_;
  assign new_n2171_ = new_n1219_;
  assign new_n2172_ = new_n2171_;
  assign new_n2173_ = new_n1226_;
  assign new_n2174_ = new_n2173_;
  assign new_n2175_ = new_n2173_;
  assign new_n2176_ = new_n1218_;
  assign new_n2177_ = new_n2176_;
  assign new_n2178_ = new_n2176_;
  assign new_n2179_ = new_n1227_;
  assign new_n2180_ = new_n2179_;
  assign new_n2181_ = new_n1210_;
  assign new_n2182_ = new_n2181_;
  assign new_n2183_ = new_n2181_;
  assign new_n2184_ = new_n1202_;
  assign new_n2185_ = new_n2184_;
  assign new_n2186_ = new_n2184_;
  assign new_n2187_ = new_n1243_;
  assign new_n2188_ = new_n1235_;
  assign new_n2189_ = new_n1274_;
  assign new_n2190_ = new_n1251_;
  assign new_n2191_ = new_n2190_;
  assign new_n2192_ = new_n1258_;
  assign new_n2193_ = new_n2192_;
  assign new_n2194_ = new_n2192_;
  assign new_n2195_ = new_n1250_;
  assign new_n2196_ = new_n2195_;
  assign new_n2197_ = new_n2195_;
  assign new_n2198_ = new_n1259_;
  assign new_n2199_ = new_n2198_;
  assign new_n2200_ = new_n1242_;
  assign new_n2201_ = new_n2200_;
  assign new_n2202_ = new_n2200_;
  assign new_n2203_ = new_n1234_;
  assign new_n2204_ = new_n2203_;
  assign new_n2205_ = new_n2203_;
  assign new_n2206_ = new_n646_;
  assign new_n2207_ = new_n2206_;
  assign new_n2208_ = new_n2207_;
  assign new_n2209_ = new_n2207_;
  assign new_n2210_ = new_n2206_;
  assign new_n2211_ = new_n2210_;
  assign new_n2212_ = new_n2210_;
  assign new_n2213_ = new_n647_;
  assign new_n2214_ = new_n2213_;
  assign new_n2215_ = new_n2214_;
  assign new_n2216_ = new_n2214_;
  assign new_n2217_ = new_n2213_;
  assign new_n2218_ = new_n2217_;
  assign new_n2219_ = new_n2217_;
  assign new_n2220_ = new_n870_;
  assign new_n2221_ = new_n2220_;
  assign new_n2222_ = new_n2220_;
  assign new_n2223_ = new_n868_;
  assign new_n2224_ = new_n2223_;
  assign new_n2225_ = new_n2223_;
  assign new_n2226_ = new_n871_;
  assign new_n2227_ = new_n2226_;
  assign new_n2228_ = new_n2226_;
  assign new_n2229_ = new_n869_;
  assign new_n2230_ = new_n2229_;
  assign new_n2231_ = new_n2229_;
  assign new_n2232_ = new_n1291_;
  assign new_n2233_ = new_n1290_;
  assign new_n2234_ = new_n1298_;
  assign new_n2235_ = new_n874_;
  assign new_n2236_ = new_n2235_;
  assign new_n2237_ = new_n2235_;
  assign new_n2238_ = new_n872_;
  assign new_n2239_ = new_n2238_;
  assign new_n2240_ = new_n2238_;
  assign new_n2241_ = new_n875_;
  assign new_n2242_ = new_n2241_;
  assign new_n2243_ = new_n2241_;
  assign new_n2244_ = new_n873_;
  assign new_n2245_ = new_n2244_;
  assign new_n2246_ = new_n2244_;
  assign new_n2247_ = new_n1305_;
  assign new_n2248_ = new_n1304_;
  assign new_n2249_ = new_n1312_;
  assign new_n2250_ = new_n1319_;
  assign new_n2251_ = new_n1318_;
  assign new_n2252_ = new_n1326_;
  assign new_n2253_ = new_n1333_;
  assign new_n2254_ = new_n1332_;
  assign new_n2255_ = new_n1340_;
  assign new_n2256_ = new_n862_;
  assign new_n2257_ = new_n2256_;
  assign new_n2258_ = new_n2256_;
  assign new_n2259_ = new_n860_;
  assign new_n2260_ = new_n2259_;
  assign new_n2261_ = new_n2259_;
  assign new_n2262_ = new_n863_;
  assign new_n2263_ = new_n2262_;
  assign new_n2264_ = new_n2262_;
  assign new_n2265_ = new_n861_;
  assign new_n2266_ = new_n2265_;
  assign new_n2267_ = new_n2265_;
  assign new_n2268_ = new_n1347_;
  assign new_n2269_ = new_n1346_;
  assign new_n2270_ = new_n1354_;
  assign new_n2271_ = new_n866_;
  assign new_n2272_ = new_n2271_;
  assign new_n2273_ = new_n2271_;
  assign new_n2274_ = new_n864_;
  assign new_n2275_ = new_n2274_;
  assign new_n2276_ = new_n2274_;
  assign new_n2277_ = new_n867_;
  assign new_n2278_ = new_n2277_;
  assign new_n2279_ = new_n2277_;
  assign new_n2280_ = new_n865_;
  assign new_n2281_ = new_n2280_;
  assign new_n2282_ = new_n2280_;
  assign new_n2283_ = new_n1361_;
  assign new_n2284_ = new_n1360_;
  assign new_n2285_ = new_n1368_;
  assign new_n2286_ = new_n1375_;
  assign new_n2287_ = new_n1374_;
  assign new_n2288_ = new_n1382_;
  assign new_n2289_ = new_n1389_;
  assign new_n2290_ = new_n1388_;
  assign new_n2291_ = new_n1396_;
  assign new_n2292_ = new_n736_;
  assign new_n2293_ = new_n728_;
  assign new_n2294_ = new_n737_;
  assign new_n2295_ = new_n2294_;
  assign new_n2296_ = new_n729_;
  assign new_n2297_ = new_n2296_;
  assign new_n2298_ = new_n1401_;
  assign new_n2299_ = new_n1400_;
  assign new_n2300_ = new_n752_;
  assign new_n2301_ = new_n744_;
  assign new_n2302_ = new_n753_;
  assign new_n2303_ = new_n2302_;
  assign new_n2304_ = new_n745_;
  assign new_n2305_ = new_n2304_;
  assign new_n2306_ = new_n1409_;
  assign new_n2307_ = new_n1408_;
  assign new_n2308_ = new_n1416_;
  assign new_n2309_ = new_n738_;
  assign new_n2310_ = new_n730_;
  assign new_n2311_ = new_n739_;
  assign new_n2312_ = new_n2311_;
  assign new_n2313_ = new_n731_;
  assign new_n2314_ = new_n2313_;
  assign new_n2315_ = new_n1421_;
  assign new_n2316_ = new_n1420_;
  assign new_n2317_ = new_n754_;
  assign new_n2318_ = new_n746_;
  assign new_n2319_ = new_n755_;
  assign new_n2320_ = new_n2319_;
  assign new_n2321_ = new_n747_;
  assign new_n2322_ = new_n2321_;
  assign new_n2323_ = new_n1429_;
  assign new_n2324_ = new_n1428_;
  assign new_n2325_ = new_n1436_;
  assign new_n2326_ = new_n740_;
  assign new_n2327_ = new_n732_;
  assign new_n2328_ = new_n741_;
  assign new_n2329_ = new_n2328_;
  assign new_n2330_ = new_n733_;
  assign new_n2331_ = new_n2330_;
  assign new_n2332_ = new_n1441_;
  assign new_n2333_ = new_n1440_;
  assign new_n2334_ = new_n756_;
  assign new_n2335_ = new_n748_;
  assign new_n2336_ = new_n757_;
  assign new_n2337_ = new_n2336_;
  assign new_n2338_ = new_n749_;
  assign new_n2339_ = new_n2338_;
  assign new_n2340_ = new_n1449_;
  assign new_n2341_ = new_n1448_;
  assign new_n2342_ = new_n1456_;
  assign new_n2343_ = new_n742_;
  assign new_n2344_ = new_n734_;
  assign new_n2345_ = new_n743_;
  assign new_n2346_ = new_n2345_;
  assign new_n2347_ = new_n735_;
  assign new_n2348_ = new_n2347_;
  assign new_n2349_ = new_n1461_;
  assign new_n2350_ = new_n1460_;
  assign new_n2351_ = new_n758_;
  assign new_n2352_ = new_n750_;
  assign new_n2353_ = new_n759_;
  assign new_n2354_ = new_n2353_;
  assign new_n2355_ = new_n751_;
  assign new_n2356_ = new_n2355_;
  assign new_n2357_ = new_n1469_;
  assign new_n2358_ = new_n1468_;
  assign new_n2359_ = new_n1476_;
  assign new_n2360_ = new_n768_;
  assign new_n2361_ = new_n760_;
  assign new_n2362_ = new_n769_;
  assign new_n2363_ = new_n2362_;
  assign new_n2364_ = new_n761_;
  assign new_n2365_ = new_n2364_;
  assign new_n2366_ = new_n1481_;
  assign new_n2367_ = new_n1480_;
  assign new_n2368_ = new_n784_;
  assign new_n2369_ = new_n776_;
  assign new_n2370_ = new_n785_;
  assign new_n2371_ = new_n2370_;
  assign new_n2372_ = new_n777_;
  assign new_n2373_ = new_n2372_;
  assign new_n2374_ = new_n1489_;
  assign new_n2375_ = new_n1488_;
  assign new_n2376_ = new_n1496_;
  assign new_n2377_ = new_n770_;
  assign new_n2378_ = new_n762_;
  assign new_n2379_ = new_n771_;
  assign new_n2380_ = new_n2379_;
  assign new_n2381_ = new_n763_;
  assign new_n2382_ = new_n2381_;
  assign new_n2383_ = new_n1501_;
  assign new_n2384_ = new_n1500_;
  assign new_n2385_ = new_n786_;
  assign new_n2386_ = new_n778_;
  assign new_n2387_ = new_n787_;
  assign new_n2388_ = new_n2387_;
  assign new_n2389_ = new_n779_;
  assign new_n2390_ = new_n2389_;
  assign new_n2391_ = new_n1509_;
  assign new_n2392_ = new_n1508_;
  assign new_n2393_ = new_n1516_;
  assign new_n2394_ = new_n772_;
  assign new_n2395_ = new_n764_;
  assign new_n2396_ = new_n773_;
  assign new_n2397_ = new_n2396_;
  assign new_n2398_ = new_n765_;
  assign new_n2399_ = new_n2398_;
  assign new_n2400_ = new_n1521_;
  assign new_n2401_ = new_n1520_;
  assign new_n2402_ = new_n788_;
  assign new_n2403_ = new_n780_;
  assign new_n2404_ = new_n789_;
  assign new_n2405_ = new_n2404_;
  assign new_n2406_ = new_n781_;
  assign new_n2407_ = new_n2406_;
  assign new_n2408_ = new_n1529_;
  assign new_n2409_ = new_n1528_;
  assign new_n2410_ = new_n1536_;
  assign new_n2411_ = new_n774_;
  assign new_n2412_ = new_n766_;
  assign new_n2413_ = new_n775_;
  assign new_n2414_ = new_n2413_;
  assign new_n2415_ = new_n767_;
  assign new_n2416_ = new_n2415_;
  assign new_n2417_ = new_n1541_;
  assign new_n2418_ = new_n1540_;
  assign new_n2419_ = new_n790_;
  assign new_n2420_ = new_n782_;
  assign new_n2421_ = new_n791_;
  assign new_n2422_ = new_n2421_;
  assign new_n2423_ = new_n783_;
  assign new_n2424_ = new_n2423_;
  assign new_n2425_ = new_n1549_;
  assign new_n2426_ = new_n1548_;
  assign new_n2427_ = new_n1556_;
  assign new_n2428_ = new_n878_;
  assign new_n2429_ = new_n876_;
  assign new_n2430_ = new_n879_;
  assign new_n2431_ = new_n2430_;
  assign new_n2432_ = new_n877_;
  assign new_n2433_ = new_n2432_;
  assign new_n2434_ = new_n1561_;
  assign new_n2435_ = new_n1560_;
  assign new_n2436_ = new_n882_;
  assign new_n2437_ = new_n880_;
  assign new_n2438_ = new_n883_;
  assign new_n2439_ = new_n2438_;
  assign new_n2440_ = new_n881_;
  assign new_n2441_ = new_n2440_;
  assign new_n2442_ = new_n1569_;
  assign new_n2443_ = new_n1568_;
  assign new_n2444_ = new_n1576_;
  assign new_n2445_ = new_n886_;
  assign new_n2446_ = new_n884_;
  assign new_n2447_ = new_n887_;
  assign new_n2448_ = new_n2447_;
  assign new_n2449_ = new_n885_;
  assign new_n2450_ = new_n2449_;
  assign new_n2451_ = new_n1581_;
  assign new_n2452_ = new_n1580_;
  assign new_n2453_ = new_n890_;
  assign new_n2454_ = new_n888_;
  assign new_n2455_ = new_n891_;
  assign new_n2456_ = new_n2455_;
  assign new_n2457_ = new_n889_;
  assign new_n2458_ = new_n2457_;
  assign new_n2459_ = new_n1589_;
  assign new_n2460_ = new_n1588_;
  assign new_n2461_ = new_n1596_;
  assign new_n2462_ = new_n894_;
  assign new_n2463_ = new_n892_;
  assign new_n2464_ = new_n895_;
  assign new_n2465_ = new_n2464_;
  assign new_n2466_ = new_n893_;
  assign new_n2467_ = new_n2466_;
  assign new_n2468_ = new_n1601_;
  assign new_n2469_ = new_n1600_;
  assign new_n2470_ = new_n898_;
  assign new_n2471_ = new_n896_;
  assign new_n2472_ = new_n899_;
  assign new_n2473_ = new_n2472_;
  assign new_n2474_ = new_n897_;
  assign new_n2475_ = new_n2474_;
  assign new_n2476_ = new_n1609_;
  assign new_n2477_ = new_n1608_;
  assign new_n2478_ = new_n1616_;
  assign new_n2479_ = new_n902_;
  assign new_n2480_ = new_n900_;
  assign new_n2481_ = new_n903_;
  assign new_n2482_ = new_n2481_;
  assign new_n2483_ = new_n901_;
  assign new_n2484_ = new_n2483_;
  assign new_n2485_ = new_n1621_;
  assign new_n2486_ = new_n1620_;
  assign new_n2487_ = new_n906_;
  assign new_n2488_ = new_n904_;
  assign new_n2489_ = new_n907_;
  assign new_n2490_ = new_n2489_;
  assign new_n2491_ = new_n905_;
  assign new_n2492_ = new_n2491_;
  assign new_n2493_ = new_n1629_;
  assign new_n2494_ = new_n1628_;
  assign new_n2495_ = new_n1636_;
  assign new_n2496_ = new_n910_;
  assign new_n2497_ = new_n908_;
  assign new_n2498_ = new_n911_;
  assign new_n2499_ = new_n2498_;
  assign new_n2500_ = new_n909_;
  assign new_n2501_ = new_n2500_;
  assign new_n2502_ = new_n1641_;
  assign new_n2503_ = new_n1640_;
  assign new_n2504_ = new_n914_;
  assign new_n2505_ = new_n912_;
  assign new_n2506_ = new_n915_;
  assign new_n2507_ = new_n2506_;
  assign new_n2508_ = new_n913_;
  assign new_n2509_ = new_n2508_;
  assign new_n2510_ = new_n1649_;
  assign new_n2511_ = new_n1648_;
  assign new_n2512_ = new_n1656_;
  assign new_n2513_ = new_n918_;
  assign new_n2514_ = new_n916_;
  assign new_n2515_ = new_n919_;
  assign new_n2516_ = new_n2515_;
  assign new_n2517_ = new_n917_;
  assign new_n2518_ = new_n2517_;
  assign new_n2519_ = new_n1661_;
  assign new_n2520_ = new_n1660_;
  assign new_n2521_ = new_n922_;
  assign new_n2522_ = new_n920_;
  assign new_n2523_ = new_n923_;
  assign new_n2524_ = new_n2523_;
  assign new_n2525_ = new_n921_;
  assign new_n2526_ = new_n2525_;
  assign new_n2527_ = new_n1669_;
  assign new_n2528_ = new_n1668_;
  assign new_n2529_ = new_n1676_;
  assign new_n2530_ = new_n926_;
  assign new_n2531_ = new_n924_;
  assign new_n2532_ = new_n927_;
  assign new_n2533_ = new_n2532_;
  assign new_n2534_ = new_n925_;
  assign new_n2535_ = new_n2534_;
  assign new_n2536_ = new_n1681_;
  assign new_n2537_ = new_n1680_;
  assign new_n2538_ = new_n930_;
  assign new_n2539_ = new_n928_;
  assign new_n2540_ = new_n931_;
  assign new_n2541_ = new_n2540_;
  assign new_n2542_ = new_n929_;
  assign new_n2543_ = new_n2542_;
  assign new_n2544_ = new_n1689_;
  assign new_n2545_ = new_n1688_;
  assign new_n2546_ = new_n1696_;
  assign new_n2547_ = new_n934_;
  assign new_n2548_ = new_n932_;
  assign new_n2549_ = new_n935_;
  assign new_n2550_ = new_n2549_;
  assign new_n2551_ = new_n933_;
  assign new_n2552_ = new_n2551_;
  assign new_n2553_ = new_n1701_;
  assign new_n2554_ = new_n1700_;
  assign new_n2555_ = new_n938_;
  assign new_n2556_ = new_n936_;
  assign new_n2557_ = new_n939_;
  assign new_n2558_ = new_n2557_;
  assign new_n2559_ = new_n937_;
  assign new_n2560_ = new_n2559_;
  assign new_n2561_ = new_n1709_;
  assign new_n2562_ = new_n1708_;
  assign new_n2563_ = new_n1716_;
  always @ (posedge clock) begin
    n630_lo <= n630_li;
    n642_lo <= n642_li;
    n654_lo <= n654_li;
    n666_lo <= n666_li;
    n678_lo <= n678_li;
    n690_lo <= n690_li;
    n702_lo <= n702_li;
    n714_lo <= n714_li;
    n726_lo <= n726_li;
    n738_lo <= n738_li;
    n750_lo <= n750_li;
    n762_lo <= n762_li;
    n774_lo <= n774_li;
    n786_lo <= n786_li;
    n798_lo <= n798_li;
    n810_lo <= n810_li;
    n822_lo <= n822_li;
    n834_lo <= n834_li;
    n846_lo <= n846_li;
    n858_lo <= n858_li;
    n870_lo <= n870_li;
    n882_lo <= n882_li;
    n894_lo <= n894_li;
    n906_lo <= n906_li;
    n918_lo <= n918_li;
    n930_lo <= n930_li;
    n942_lo <= n942_li;
    n954_lo <= n954_li;
    n966_lo <= n966_li;
    n978_lo <= n978_li;
    n990_lo <= n990_li;
    n1002_lo <= n1002_li;
    n1005_lo <= n1005_li;
    n1008_lo <= n1008_li;
    n1017_lo <= n1017_li;
    n1020_lo <= n1020_li;
    n1029_lo <= n1029_li;
    n1032_lo <= n1032_li;
    n1041_lo <= n1041_li;
    n1044_lo <= n1044_li;
    n1053_lo <= n1053_li;
    n1056_lo <= n1056_li;
    n1065_lo <= n1065_li;
    n1068_lo <= n1068_li;
    n1077_lo <= n1077_li;
    n1080_lo <= n1080_li;
    n1089_lo <= n1089_li;
    n1092_lo <= n1092_li;
    n1101_lo <= n1101_li;
    n1104_lo <= n1104_li;
    n1837_o2 <= n1837_i2;
    n1838_o2 <= n1838_i2;
    n1839_o2 <= n1839_i2;
    n1840_o2 <= n1840_i2;
    n1841_o2 <= n1841_i2;
    n1842_o2 <= n1842_i2;
    n1843_o2 <= n1843_i2;
    n1844_o2 <= n1844_i2;
    n1845_o2 <= n1845_i2;
    n1846_o2 <= n1846_i2;
    n1847_o2 <= n1847_i2;
    n1848_o2 <= n1848_i2;
    n1849_o2 <= n1849_i2;
    n1850_o2 <= n1850_i2;
    n1851_o2 <= n1851_i2;
    n1852_o2 <= n1852_i2;
    n1853_o2 <= n1853_i2;
    n1854_o2 <= n1854_i2;
    n1855_o2 <= n1855_i2;
    n1856_o2 <= n1856_i2;
    n1857_o2 <= n1857_i2;
    n1858_o2 <= n1858_i2;
    n1859_o2 <= n1859_i2;
    n1860_o2 <= n1860_i2;
    n1861_o2 <= n1861_i2;
    n1862_o2 <= n1862_i2;
    n1863_o2 <= n1863_i2;
    n1864_o2 <= n1864_i2;
    n1865_o2 <= n1865_i2;
    n1866_o2 <= n1866_i2;
    n1867_o2 <= n1867_i2;
    n1868_o2 <= n1868_i2;
    G834_o2 <= G834_i2;
    G847_o2 <= G847_i2;
    G860_o2 <= G860_i2;
    G873_o2 <= G873_i2;
    G925_o2 <= G925_i2;
    G886_o2 <= G886_i2;
    G912_o2 <= G912_i2;
    G899_o2 <= G899_i2;
    n2151_o2 <= n2151_i2;
    n2152_o2 <= n2152_i2;
    n2153_o2 <= n2153_i2;
    n2154_o2 <= n2154_i2;
    n2155_o2 <= n2155_i2;
    n2156_o2 <= n2156_i2;
    n2157_o2 <= n2157_i2;
    n2158_o2 <= n2158_i2;
    n2159_o2 <= n2159_i2;
    n2160_o2 <= n2160_i2;
    n2161_o2 <= n2161_i2;
    n2162_o2 <= n2162_i2;
    n2163_o2 <= n2163_i2;
    n2164_o2 <= n2164_i2;
    n2165_o2 <= n2165_i2;
    n2166_o2 <= n2166_i2;
    n2167_o2 <= n2167_i2;
    n2168_o2 <= n2168_i2;
    n2169_o2 <= n2169_i2;
    n2170_o2 <= n2170_i2;
    n2171_o2 <= n2171_i2;
    n2172_o2 <= n2172_i2;
    n2173_o2 <= n2173_i2;
    n2174_o2 <= n2174_i2;
    n2175_o2 <= n2175_i2;
    n2176_o2 <= n2176_i2;
    n2177_o2 <= n2177_i2;
    n2178_o2 <= n2178_i2;
    n2179_o2 <= n2179_i2;
    n2180_o2 <= n2180_i2;
    n2181_o2 <= n2181_i2;
    n2182_o2 <= n2182_i2;
    G974_o2 <= G974_i2;
    G976_o2 <= G976_i2;
    G970_o2 <= G970_i2;
    G972_o2 <= G972_i2;
    G973_o2 <= G973_i2;
    G977_o2 <= G977_i2;
    G971_o2 <= G971_i2;
    G975_o2 <= G975_i2;
    G954_o2 <= G954_i2;
    G956_o2 <= G956_i2;
    G950_o2 <= G950_i2;
    G952_o2 <= G952_i2;
    G953_o2 <= G953_i2;
    G957_o2 <= G957_i2;
    G951_o2 <= G951_i2;
    G955_o2 <= G955_i2;
    G986_o2 <= G986_i2;
    G991_o2 <= G991_i2;
    G770_o2 <= G770_i2;
    G773_o2 <= G773_i2;
    G776_o2 <= G776_i2;
    G779_o2 <= G779_i2;
    G782_o2 <= G782_i2;
    G785_o2 <= G785_i2;
    G788_o2 <= G788_i2;
    G791_o2 <= G791_i2;
    G642_o2 <= G642_i2;
    G645_o2 <= G645_i2;
    G648_o2 <= G648_i2;
    G651_o2 <= G651_i2;
    G654_o2 <= G654_i2;
    G657_o2 <= G657_i2;
    G660_o2 <= G660_i2;
    G663_o2 <= G663_i2;
    G602_o2 <= G602_i2;
    G607_o2 <= G607_i2;
    G612_o2 <= G612_i2;
    G617_o2 <= G617_i2;
    G622_o2 <= G622_i2;
    G627_o2 <= G627_i2;
    G632_o2 <= G632_i2;
    G637_o2 <= G637_i2;
    n627_lo_buf_o2 <= n627_lo_buf_i2;
    n639_lo_buf_o2 <= n639_lo_buf_i2;
    n651_lo_buf_o2 <= n651_lo_buf_i2;
    n663_lo_buf_o2 <= n663_lo_buf_i2;
    n675_lo_buf_o2 <= n675_lo_buf_i2;
    n687_lo_buf_o2 <= n687_lo_buf_i2;
    n699_lo_buf_o2 <= n699_lo_buf_i2;
    n711_lo_buf_o2 <= n711_lo_buf_i2;
    n723_lo_buf_o2 <= n723_lo_buf_i2;
    n735_lo_buf_o2 <= n735_lo_buf_i2;
    n747_lo_buf_o2 <= n747_lo_buf_i2;
    n759_lo_buf_o2 <= n759_lo_buf_i2;
    n771_lo_buf_o2 <= n771_lo_buf_i2;
    n783_lo_buf_o2 <= n783_lo_buf_i2;
    n795_lo_buf_o2 <= n795_lo_buf_i2;
    n807_lo_buf_o2 <= n807_lo_buf_i2;
    n819_lo_buf_o2 <= n819_lo_buf_i2;
    n831_lo_buf_o2 <= n831_lo_buf_i2;
    n843_lo_buf_o2 <= n843_lo_buf_i2;
    n855_lo_buf_o2 <= n855_lo_buf_i2;
    n867_lo_buf_o2 <= n867_lo_buf_i2;
    n879_lo_buf_o2 <= n879_lo_buf_i2;
    n891_lo_buf_o2 <= n891_lo_buf_i2;
    n903_lo_buf_o2 <= n903_lo_buf_i2;
    n915_lo_buf_o2 <= n915_lo_buf_i2;
    n927_lo_buf_o2 <= n927_lo_buf_i2;
    n939_lo_buf_o2 <= n939_lo_buf_i2;
    n951_lo_buf_o2 <= n951_lo_buf_i2;
    n963_lo_buf_o2 <= n963_lo_buf_i2;
    n975_lo_buf_o2 <= n975_lo_buf_i2;
    n987_lo_buf_o2 <= n987_lo_buf_i2;
    n999_lo_buf_o2 <= n999_lo_buf_i2;
  end
  initial begin
    n630_lo <= 1'b0;
    n642_lo <= 1'b0;
    n654_lo <= 1'b0;
    n666_lo <= 1'b0;
    n678_lo <= 1'b0;
    n690_lo <= 1'b0;
    n702_lo <= 1'b0;
    n714_lo <= 1'b0;
    n726_lo <= 1'b0;
    n738_lo <= 1'b0;
    n750_lo <= 1'b0;
    n762_lo <= 1'b0;
    n774_lo <= 1'b0;
    n786_lo <= 1'b0;
    n798_lo <= 1'b0;
    n810_lo <= 1'b0;
    n822_lo <= 1'b0;
    n834_lo <= 1'b0;
    n846_lo <= 1'b0;
    n858_lo <= 1'b0;
    n870_lo <= 1'b0;
    n882_lo <= 1'b0;
    n894_lo <= 1'b0;
    n906_lo <= 1'b0;
    n918_lo <= 1'b0;
    n930_lo <= 1'b0;
    n942_lo <= 1'b0;
    n954_lo <= 1'b0;
    n966_lo <= 1'b0;
    n978_lo <= 1'b0;
    n990_lo <= 1'b0;
    n1002_lo <= 1'b0;
    n1005_lo <= 1'b0;
    n1008_lo <= 1'b0;
    n1017_lo <= 1'b0;
    n1020_lo <= 1'b0;
    n1029_lo <= 1'b0;
    n1032_lo <= 1'b0;
    n1041_lo <= 1'b0;
    n1044_lo <= 1'b0;
    n1053_lo <= 1'b0;
    n1056_lo <= 1'b0;
    n1065_lo <= 1'b0;
    n1068_lo <= 1'b0;
    n1077_lo <= 1'b0;
    n1080_lo <= 1'b0;
    n1089_lo <= 1'b0;
    n1092_lo <= 1'b0;
    n1101_lo <= 1'b0;
    n1104_lo <= 1'b0;
    n1837_o2 <= 1'b0;
    n1838_o2 <= 1'b0;
    n1839_o2 <= 1'b0;
    n1840_o2 <= 1'b0;
    n1841_o2 <= 1'b0;
    n1842_o2 <= 1'b0;
    n1843_o2 <= 1'b0;
    n1844_o2 <= 1'b0;
    n1845_o2 <= 1'b0;
    n1846_o2 <= 1'b0;
    n1847_o2 <= 1'b0;
    n1848_o2 <= 1'b0;
    n1849_o2 <= 1'b0;
    n1850_o2 <= 1'b0;
    n1851_o2 <= 1'b0;
    n1852_o2 <= 1'b0;
    n1853_o2 <= 1'b0;
    n1854_o2 <= 1'b0;
    n1855_o2 <= 1'b0;
    n1856_o2 <= 1'b0;
    n1857_o2 <= 1'b0;
    n1858_o2 <= 1'b0;
    n1859_o2 <= 1'b0;
    n1860_o2 <= 1'b0;
    n1861_o2 <= 1'b0;
    n1862_o2 <= 1'b0;
    n1863_o2 <= 1'b0;
    n1864_o2 <= 1'b0;
    n1865_o2 <= 1'b0;
    n1866_o2 <= 1'b0;
    n1867_o2 <= 1'b0;
    n1868_o2 <= 1'b0;
    G834_o2 <= 1'b0;
    G847_o2 <= 1'b0;
    G860_o2 <= 1'b0;
    G873_o2 <= 1'b0;
    G925_o2 <= 1'b0;
    G886_o2 <= 1'b0;
    G912_o2 <= 1'b0;
    G899_o2 <= 1'b0;
    n2151_o2 <= 1'b0;
    n2152_o2 <= 1'b0;
    n2153_o2 <= 1'b0;
    n2154_o2 <= 1'b0;
    n2155_o2 <= 1'b0;
    n2156_o2 <= 1'b0;
    n2157_o2 <= 1'b0;
    n2158_o2 <= 1'b0;
    n2159_o2 <= 1'b0;
    n2160_o2 <= 1'b0;
    n2161_o2 <= 1'b0;
    n2162_o2 <= 1'b0;
    n2163_o2 <= 1'b0;
    n2164_o2 <= 1'b0;
    n2165_o2 <= 1'b0;
    n2166_o2 <= 1'b0;
    n2167_o2 <= 1'b0;
    n2168_o2 <= 1'b0;
    n2169_o2 <= 1'b0;
    n2170_o2 <= 1'b0;
    n2171_o2 <= 1'b0;
    n2172_o2 <= 1'b0;
    n2173_o2 <= 1'b0;
    n2174_o2 <= 1'b0;
    n2175_o2 <= 1'b0;
    n2176_o2 <= 1'b0;
    n2177_o2 <= 1'b0;
    n2178_o2 <= 1'b0;
    n2179_o2 <= 1'b0;
    n2180_o2 <= 1'b0;
    n2181_o2 <= 1'b0;
    n2182_o2 <= 1'b0;
    G974_o2 <= 1'b0;
    G976_o2 <= 1'b0;
    G970_o2 <= 1'b0;
    G972_o2 <= 1'b0;
    G973_o2 <= 1'b0;
    G977_o2 <= 1'b0;
    G971_o2 <= 1'b0;
    G975_o2 <= 1'b0;
    G954_o2 <= 1'b0;
    G956_o2 <= 1'b0;
    G950_o2 <= 1'b0;
    G952_o2 <= 1'b0;
    G953_o2 <= 1'b0;
    G957_o2 <= 1'b0;
    G951_o2 <= 1'b0;
    G955_o2 <= 1'b0;
    G986_o2 <= 1'b0;
    G991_o2 <= 1'b0;
    G770_o2 <= 1'b0;
    G773_o2 <= 1'b0;
    G776_o2 <= 1'b0;
    G779_o2 <= 1'b0;
    G782_o2 <= 1'b0;
    G785_o2 <= 1'b0;
    G788_o2 <= 1'b0;
    G791_o2 <= 1'b0;
    G642_o2 <= 1'b0;
    G645_o2 <= 1'b0;
    G648_o2 <= 1'b0;
    G651_o2 <= 1'b0;
    G654_o2 <= 1'b0;
    G657_o2 <= 1'b0;
    G660_o2 <= 1'b0;
    G663_o2 <= 1'b0;
    G602_o2 <= 1'b0;
    G607_o2 <= 1'b0;
    G612_o2 <= 1'b0;
    G617_o2 <= 1'b0;
    G622_o2 <= 1'b0;
    G627_o2 <= 1'b0;
    G632_o2 <= 1'b0;
    G637_o2 <= 1'b0;
    n627_lo_buf_o2 <= 1'b0;
    n639_lo_buf_o2 <= 1'b0;
    n651_lo_buf_o2 <= 1'b0;
    n663_lo_buf_o2 <= 1'b0;
    n675_lo_buf_o2 <= 1'b0;
    n687_lo_buf_o2 <= 1'b0;
    n699_lo_buf_o2 <= 1'b0;
    n711_lo_buf_o2 <= 1'b0;
    n723_lo_buf_o2 <= 1'b0;
    n735_lo_buf_o2 <= 1'b0;
    n747_lo_buf_o2 <= 1'b0;
    n759_lo_buf_o2 <= 1'b0;
    n771_lo_buf_o2 <= 1'b0;
    n783_lo_buf_o2 <= 1'b0;
    n795_lo_buf_o2 <= 1'b0;
    n807_lo_buf_o2 <= 1'b0;
    n819_lo_buf_o2 <= 1'b0;
    n831_lo_buf_o2 <= 1'b0;
    n843_lo_buf_o2 <= 1'b0;
    n855_lo_buf_o2 <= 1'b0;
    n867_lo_buf_o2 <= 1'b0;
    n879_lo_buf_o2 <= 1'b0;
    n891_lo_buf_o2 <= 1'b0;
    n903_lo_buf_o2 <= 1'b0;
    n915_lo_buf_o2 <= 1'b0;
    n927_lo_buf_o2 <= 1'b0;
    n939_lo_buf_o2 <= 1'b0;
    n951_lo_buf_o2 <= 1'b0;
    n963_lo_buf_o2 <= 1'b0;
    n975_lo_buf_o2 <= 1'b0;
    n987_lo_buf_o2 <= 1'b0;
    n999_lo_buf_o2 <= 1'b0;
  end
endmodule


