
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  G42,
  G43,
  G44,
  G45,
  G46,
  G47,
  G48,
  G49,
  G50,
  G51,
  G52,
  G53,
  G54,
  G55,
  G56,
  G57,
  G58,
  G59,
  G60,
  G855,
  G856,
  G857,
  G858,
  G859,
  G860,
  G861,
  G862,
  G863,
  G864,
  G865,
  G866,
  G867,
  G868,
  G869,
  G870,
  G871,
  G872,
  G873,
  G874,
  G875,
  G876,
  G877,
  G878,
  G879,
  G880
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input G42;input G43;input G44;input G45;input G46;input G47;input G48;input G49;input G50;input G51;input G52;input G53;input G54;input G55;input G56;input G57;input G58;input G59;input G60;
  output G855;output G856;output G857;output G858;output G859;output G860;output G861;output G862;output G863;output G864;output G865;output G866;output G867;output G868;output G869;output G870;output G871;output G872;output G873;output G874;output G875;output G876;output G877;output G878;output G879;output G880;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire G51_p;
  wire G51_n;
  wire G52_p;
  wire G52_n;
  wire G53_p;
  wire G53_n;
  wire G54_p;
  wire G54_n;
  wire G55_p;
  wire G55_n;
  wire G56_p;
  wire G56_n;
  wire G57_p;
  wire G57_n;
  wire G58_p;
  wire G58_n;
  wire G59_p;
  wire G59_n;
  wire G60_p;
  wire G60_n;
  wire g61_p;
  wire g61_n;
  wire g62_p;
  wire g62_n;
  wire g63_p;
  wire g63_n;
  wire g64_p;
  wire g64_n;
  wire g65_p;
  wire g65_n;
  wire g66_p;
  wire g66_n;
  wire g67_p;
  wire g67_n;
  wire g68_p;
  wire g68_n;
  wire g69_p;
  wire g69_n;
  wire g70_p;
  wire g70_n;
  wire g71_p;
  wire g71_n;
  wire g72_p;
  wire g72_n;
  wire g73_p;
  wire g73_n;
  wire g74_p;
  wire g74_n;
  wire g75_p;
  wire g75_n;
  wire g76_p;
  wire g76_n;
  wire g77_p;
  wire g77_n;
  wire g78_p;
  wire g78_n;
  wire g79_p;
  wire g79_n;
  wire g80_p;
  wire g80_n;
  wire g81_p;
  wire g81_n;
  wire g82_p;
  wire g82_n;
  wire g83_p;
  wire g83_n;
  wire g84_p;
  wire g84_n;
  wire g85_p;
  wire g85_n;
  wire g86_p;
  wire g86_n;
  wire g87_p;
  wire g87_n;
  wire g88_p;
  wire g88_n;
  wire g89_p;
  wire g89_n;
  wire g90_p;
  wire g90_n;
  wire g91_p;
  wire g91_n;
  wire g92_p;
  wire g92_n;
  wire g93_p;
  wire g93_n;
  wire g94_p;
  wire g94_n;
  wire g95_p;
  wire g95_n;
  wire g96_p;
  wire g96_n;
  wire g97_p;
  wire g97_n;
  wire g98_p;
  wire g98_n;
  wire g99_p;
  wire g99_n;
  wire g100_p;
  wire g100_n;
  wire g101_p;
  wire g101_n;
  wire g102_p;
  wire g102_n;
  wire g103_p;
  wire g103_n;
  wire g104_p;
  wire g104_n;
  wire g105_p;
  wire g105_n;
  wire g106_p;
  wire g106_n;
  wire g107_p;
  wire g107_n;
  wire g108_p;
  wire g108_n;
  wire g109_p;
  wire g109_n;
  wire g110_p;
  wire g110_n;
  wire g111_p;
  wire g111_n;
  wire g112_p;
  wire g112_n;
  wire g113_p;
  wire g113_n;
  wire g114_p;
  wire g114_n;
  wire g115_p;
  wire g115_n;
  wire g116_p;
  wire g116_n;
  wire g117_p;
  wire g117_n;
  wire g118_p;
  wire g118_n;
  wire g119_p;
  wire g119_n;
  wire g120_p;
  wire g120_n;
  wire g121_p;
  wire g121_n;
  wire g122_p;
  wire g122_n;
  wire g123_p;
  wire g123_n;
  wire g124_p;
  wire g124_n;
  wire g125_p;
  wire g125_n;
  wire g126_p;
  wire g126_n;
  wire g127_p;
  wire g127_n;
  wire g128_p;
  wire g128_n;
  wire g129_p;
  wire g129_n;
  wire g130_p;
  wire g130_n;
  wire g131_p;
  wire g131_n;
  wire g132_p;
  wire g132_n;
  wire g133_p;
  wire g133_n;
  wire g134_p;
  wire g134_n;
  wire g135_p;
  wire g135_n;
  wire g136_p;
  wire g136_n;
  wire g137_p;
  wire g137_n;
  wire g138_p;
  wire g138_n;
  wire g139_p;
  wire g139_n;
  wire g140_p;
  wire g140_n;
  wire g141_p;
  wire g141_n;
  wire g142_p;
  wire g142_n;
  wire g143_p;
  wire g143_n;
  wire g144_p;
  wire g144_n;
  wire g145_p;
  wire g145_n;
  wire g146_p;
  wire g146_n;
  wire g147_p;
  wire g147_n;
  wire g148_p;
  wire g148_n;
  wire g149_p;
  wire g149_n;
  wire g150_p;
  wire g150_n;
  wire g151_p;
  wire g151_n;
  wire g152_p;
  wire g152_n;
  wire g153_p;
  wire g153_n;
  wire g154_p;
  wire g154_n;
  wire g155_p;
  wire g155_n;
  wire g156_p;
  wire g156_n;
  wire g157_p;
  wire g157_n;
  wire g158_p;
  wire g158_n;
  wire g159_p;
  wire g159_n;
  wire g160_p;
  wire g160_n;
  wire g161_p;
  wire g161_n;
  wire g162_p;
  wire g162_n;
  wire g163_p;
  wire g163_n;
  wire g164_p;
  wire g164_n;
  wire g165_p;
  wire g165_n;
  wire g166_p;
  wire g166_n;
  wire g167_p;
  wire g167_n;
  wire g168_p;
  wire g168_n;
  wire g169_p;
  wire g169_n;
  wire g170_p;
  wire g170_n;
  wire g171_p;
  wire g171_n;
  wire g172_p;
  wire g172_n;
  wire g173_p;
  wire g173_n;
  wire g174_p;
  wire g174_n;
  wire g175_p;
  wire g175_n;
  wire g176_p;
  wire g176_n;
  wire g177_p;
  wire g177_n;
  wire g178_p;
  wire g178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire G16_p_spl_;
  wire G6_n_spl_;
  wire G6_n_spl_0;
  wire G16_n_spl_;
  wire G8_n_spl_;
  wire G8_n_spl_0;
  wire G8_n_spl_00;
  wire G8_n_spl_01;
  wire G8_n_spl_1;
  wire G8_n_spl_10;
  wire g61_n_spl_;
  wire G7_n_spl_;
  wire G17_n_spl_;
  wire G17_n_spl_0;
  wire g63_n_spl_;
  wire G1_p_spl_;
  wire G1_p_spl_0;
  wire G2_p_spl_;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire G2_n_spl_;
  wire G3_n_spl_;
  wire g67_n_spl_;
  wire G4_n_spl_;
  wire G4_n_spl_0;
  wire G4_n_spl_00;
  wire G4_n_spl_01;
  wire G4_n_spl_1;
  wire G4_n_spl_10;
  wire G4_n_spl_11;
  wire g68_n_spl_;
  wire g70_p_spl_;
  wire g70_n_spl_;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_00;
  wire G4_p_spl_01;
  wire G4_p_spl_1;
  wire G4_p_spl_10;
  wire g65_n_spl_;
  wire g65_n_spl_0;
  wire G11_p_spl_;
  wire G11_n_spl_;
  wire G11_n_spl_0;
  wire G11_n_spl_1;
  wire G17_p_spl_;
  wire g74_p_spl_;
  wire g76_n_spl_;
  wire g79_n_spl_;
  wire G9_p_spl_;
  wire G9_p_spl_0;
  wire G9_n_spl_;
  wire G9_n_spl_0;
  wire G10_n_spl_;
  wire G10_n_spl_0;
  wire g83_n_spl_;
  wire g83_n_spl_0;
  wire G12_n_spl_;
  wire g86_n_spl_;
  wire G24_p_spl_;
  wire G24_p_spl_0;
  wire G25_n_spl_;
  wire G25_n_spl_0;
  wire G25_n_spl_1;
  wire G24_n_spl_;
  wire G24_n_spl_0;
  wire G24_n_spl_1;
  wire G25_p_spl_;
  wire G25_p_spl_0;
  wire G26_p_spl_;
  wire G26_p_spl_0;
  wire G27_n_spl_;
  wire G27_n_spl_0;
  wire G27_n_spl_1;
  wire G26_n_spl_;
  wire G26_n_spl_0;
  wire G26_n_spl_1;
  wire G27_p_spl_;
  wire G27_p_spl_0;
  wire g92_p_spl_;
  wire g95_p_spl_;
  wire g92_n_spl_;
  wire g95_n_spl_;
  wire G32_p_spl_;
  wire G32_p_spl_0;
  wire G32_p_spl_1;
  wire g98_p_spl_;
  wire G32_n_spl_;
  wire G32_n_spl_0;
  wire G32_n_spl_1;
  wire g98_n_spl_;
  wire G28_p_spl_;
  wire G28_p_spl_0;
  wire G29_n_spl_;
  wire G29_n_spl_0;
  wire G29_n_spl_1;
  wire G28_n_spl_;
  wire G28_n_spl_0;
  wire G28_n_spl_1;
  wire G29_p_spl_;
  wire G29_p_spl_0;
  wire G30_p_spl_;
  wire G30_p_spl_0;
  wire G31_n_spl_;
  wire G31_n_spl_0;
  wire G30_n_spl_;
  wire G30_n_spl_0;
  wire G30_n_spl_1;
  wire G31_p_spl_;
  wire G31_p_spl_0;
  wire g104_p_spl_;
  wire g107_p_spl_;
  wire g104_n_spl_;
  wire g107_n_spl_;
  wire G33_p_spl_;
  wire g110_p_spl_;
  wire G33_n_spl_;
  wire g110_n_spl_;
  wire G41_p_spl_;
  wire G41_p_spl_0;
  wire G41_p_spl_1;
  wire G42_n_spl_;
  wire G42_n_spl_0;
  wire G42_n_spl_00;
  wire G42_n_spl_1;
  wire G41_n_spl_;
  wire G41_n_spl_0;
  wire G41_n_spl_00;
  wire G41_n_spl_1;
  wire G42_p_spl_;
  wire G42_p_spl_0;
  wire G42_p_spl_1;
  wire G43_p_spl_;
  wire G43_p_spl_0;
  wire G43_p_spl_1;
  wire G44_n_spl_;
  wire G44_n_spl_0;
  wire G44_n_spl_00;
  wire G44_n_spl_1;
  wire G43_n_spl_;
  wire G43_n_spl_0;
  wire G43_n_spl_00;
  wire G43_n_spl_1;
  wire G44_p_spl_;
  wire G44_p_spl_0;
  wire G44_p_spl_1;
  wire g119_p_spl_;
  wire g122_p_spl_;
  wire g119_n_spl_;
  wire g122_n_spl_;
  wire g125_p_spl_;
  wire g125_n_spl_;
  wire G45_p_spl_;
  wire G45_p_spl_0;
  wire G45_p_spl_1;
  wire G46_n_spl_;
  wire G46_n_spl_0;
  wire G46_n_spl_00;
  wire G46_n_spl_1;
  wire G45_n_spl_;
  wire G45_n_spl_0;
  wire G45_n_spl_00;
  wire G45_n_spl_1;
  wire G46_p_spl_;
  wire G46_p_spl_0;
  wire G46_p_spl_1;
  wire G47_p_spl_;
  wire G47_p_spl_0;
  wire G47_p_spl_1;
  wire G48_n_spl_;
  wire G48_n_spl_0;
  wire G48_n_spl_00;
  wire G48_n_spl_1;
  wire G47_n_spl_;
  wire G47_n_spl_0;
  wire G47_n_spl_00;
  wire G47_n_spl_1;
  wire G48_p_spl_;
  wire G48_p_spl_0;
  wire G48_p_spl_1;
  wire g131_p_spl_;
  wire g134_p_spl_;
  wire g131_n_spl_;
  wire g134_n_spl_;
  wire G49_p_spl_;
  wire g137_p_spl_;
  wire G49_n_spl_;
  wire g137_n_spl_;
  wire G55_n_spl_;
  wire G55_n_spl_0;
  wire G50_n_spl_;
  wire G50_n_spl_0;
  wire G50_n_spl_00;
  wire G50_n_spl_01;
  wire G50_n_spl_1;
  wire G50_n_spl_10;
  wire G50_n_spl_11;
  wire g82_p_spl_;
  wire g82_p_spl_0;
  wire g82_n_spl_;
  wire g82_n_spl_0;
  wire g82_n_spl_1;
  wire G10_p_spl_;
  wire g147_p_spl_;
  wire g147_n_spl_;
  wire G60_n_spl_;
  wire G60_n_spl_0;
  wire G60_p_spl_;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire g153_p_spl_;
  wire g153_n_spl_;
  wire g160_n_spl_;
  wire g160_n_spl_0;
  wire g160_n_spl_00;
  wire g160_n_spl_01;
  wire g160_n_spl_1;
  wire g160_n_spl_10;
  wire g160_n_spl_11;
  wire g160_p_spl_;
  wire g160_p_spl_0;
  wire g160_p_spl_00;
  wire g160_p_spl_01;
  wire g160_p_spl_1;
  wire g160_p_spl_10;
  wire g160_p_spl_11;
  wire g162_p_spl_;
  wire g162_n_spl_;
  wire G39_p_spl_;
  wire g164_n_spl_;
  wire g164_n_spl_0;
  wire g164_n_spl_1;
  wire G39_n_spl_;
  wire g164_p_spl_;
  wire g164_p_spl_0;
  wire g164_p_spl_1;
  wire g149_n_spl_;
  wire g149_n_spl_0;
  wire g149_n_spl_1;
  wire g149_p_spl_;
  wire g149_p_spl_0;
  wire g149_p_spl_1;
  wire G54_n_spl_;
  wire G54_n_spl_0;
  wire G54_n_spl_00;
  wire G54_n_spl_01;
  wire G54_n_spl_1;
  wire G54_n_spl_10;
  wire G54_n_spl_11;
  wire g167_p_spl_;
  wire g167_p_spl_0;
  wire g172_n_spl_;
  wire g172_n_spl_0;
  wire g172_n_spl_00;
  wire g172_n_spl_01;
  wire g172_n_spl_1;
  wire g172_n_spl_10;
  wire g172_n_spl_11;
  wire g167_n_spl_;
  wire G53_n_spl_;
  wire G53_n_spl_0;
  wire G53_n_spl_00;
  wire G53_n_spl_01;
  wire G53_n_spl_1;
  wire G53_n_spl_10;
  wire G53_n_spl_11;
  wire g174_p_spl_;
  wire g176_p_spl_;
  wire G51_n_spl_;
  wire G51_n_spl_0;
  wire G51_n_spl_00;
  wire G51_n_spl_000;
  wire G51_n_spl_001;
  wire G51_n_spl_01;
  wire G51_n_spl_010;
  wire G51_n_spl_011;
  wire G51_n_spl_1;
  wire G51_n_spl_10;
  wire G51_n_spl_11;
  wire G58_n_spl_;
  wire g180_p_spl_;
  wire G52_n_spl_;
  wire G52_n_spl_0;
  wire G52_n_spl_00;
  wire G52_n_spl_01;
  wire G52_n_spl_1;
  wire G52_n_spl_10;
  wire G52_n_spl_11;
  wire g174_n_spl_;
  wire G35_p_spl_;
  wire G35_n_spl_;
  wire g194_p_spl_;
  wire g194_p_spl_0;
  wire G36_p_spl_;
  wire G36_n_spl_;
  wire g199_n_spl_;
  wire g199_p_spl_;
  wire g199_p_spl_0;
  wire G37_p_spl_;
  wire G37_n_spl_;
  wire g205_n_spl_;
  wire g205_p_spl_;
  wire g205_p_spl_0;
  wire g207_p_spl_;
  wire g208_p_spl_;
  wire g206_n_spl_;
  wire g206_p_spl_;
  wire g209_p_spl_;
  wire g201_p_spl_;
  wire g210_p_spl_;
  wire g200_n_spl_;
  wire g200_p_spl_;
  wire g211_p_spl_;
  wire g212_p_spl_;
  wire g194_n_spl_;
  wire g214_p_spl_;
  wire g216_p_spl_;
  wire g219_p_spl_;
  wire g214_n_spl_;
  wire g259_p_spl_;
  wire g259_p_spl_0;
  wire g259_p_spl_1;
  wire g259_n_spl_;
  wire g259_n_spl_0;
  wire g259_n_spl_1;
  wire G34_p_spl_;
  wire G34_p_spl_0;
  wire G34_p_spl_1;
  wire G34_n_spl_;
  wire G34_n_spl_0;
  wire G34_n_spl_1;
  wire g265_n_spl_;
  wire g265_n_spl_0;
  wire g265_n_spl_1;
  wire g265_p_spl_;
  wire g265_p_spl_0;
  wire g265_p_spl_1;
  wire g267_n_spl_;
  wire g267_p_spl_;
  wire g267_p_spl_0;
  wire g274_n_spl_;
  wire g274_p_spl_;
  wire g274_p_spl_0;
  wire g282_n_spl_;
  wire g282_p_spl_;
  wire g282_p_spl_0;
  wire g291_p_spl_;
  wire g291_p_spl_0;
  wire g291_n_spl_;
  wire g285_n_spl_;
  wire g292_n_spl_;
  wire g285_p_spl_;
  wire g292_p_spl_;
  wire g294_n_spl_;
  wire g294_n_spl_0;
  wire g294_p_spl_;
  wire g284_n_spl_;
  wire g295_n_spl_;
  wire g284_p_spl_;
  wire g295_p_spl_;
  wire g283_n_spl_;
  wire g283_n_spl_0;
  wire g283_p_spl_;
  wire g276_n_spl_;
  wire g297_n_spl_;
  wire g276_p_spl_;
  wire g297_p_spl_;
  wire g275_n_spl_;
  wire g275_n_spl_0;
  wire g275_p_spl_;
  wire g299_p_spl_;
  wire g300_p_spl_;
  wire g268_n_spl_;
  wire g268_n_spl_0;
  wire g303_n_spl_;
  wire g322_n_spl_;
  wire g337_n_spl_;
  wire g352_n_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  buf

  (
    G42_p,
    G42
  );


  not

  (
    G42_n,
    G42
  );


  buf

  (
    G43_p,
    G43
  );


  not

  (
    G43_n,
    G43
  );


  buf

  (
    G44_p,
    G44
  );


  not

  (
    G44_n,
    G44
  );


  buf

  (
    G45_p,
    G45
  );


  not

  (
    G45_n,
    G45
  );


  buf

  (
    G46_p,
    G46
  );


  not

  (
    G46_n,
    G46
  );


  buf

  (
    G47_p,
    G47
  );


  not

  (
    G47_n,
    G47
  );


  buf

  (
    G48_p,
    G48
  );


  not

  (
    G48_n,
    G48
  );


  buf

  (
    G49_p,
    G49
  );


  not

  (
    G49_n,
    G49
  );


  buf

  (
    G50_p,
    G50
  );


  not

  (
    G50_n,
    G50
  );


  buf

  (
    G51_p,
    G51
  );


  not

  (
    G51_n,
    G51
  );


  buf

  (
    G52_p,
    G52
  );


  not

  (
    G52_n,
    G52
  );


  buf

  (
    G53_p,
    G53
  );


  not

  (
    G53_n,
    G53
  );


  buf

  (
    G54_p,
    G54
  );


  not

  (
    G54_n,
    G54
  );


  buf

  (
    G55_p,
    G55
  );


  not

  (
    G55_n,
    G55
  );


  buf

  (
    G56_p,
    G56
  );


  not

  (
    G56_n,
    G56
  );


  buf

  (
    G57_p,
    G57
  );


  not

  (
    G57_n,
    G57
  );


  buf

  (
    G58_p,
    G58
  );


  not

  (
    G58_n,
    G58
  );


  buf

  (
    G59_p,
    G59
  );


  not

  (
    G59_n,
    G59
  );


  buf

  (
    G60_p,
    G60
  );


  not

  (
    G60_n,
    G60
  );


  and

  (
    g61_p,
    G6_p,
    G16_p_spl_
  );


  or

  (
    g61_n,
    G6_n_spl_0,
    G16_n_spl_
  );


  or

  (
    g62_n,
    G8_n_spl_00,
    g61_n_spl_
  );


  or

  (
    g63_n,
    G6_n_spl_0,
    G7_n_spl_
  );


  or

  (
    g64_n,
    G17_n_spl_0,
    g63_n_spl_
  );


  or

  (
    g65_n,
    G8_n_spl_00,
    g63_n_spl_
  );


  or

  (
    g66_n,
    G18_n,
    G19_n
  );


  and

  (
    g67_p,
    G1_p_spl_0,
    G2_p_spl_
  );


  or

  (
    g67_n,
    G1_n_spl_0,
    G2_n_spl_
  );


  or

  (
    g68_n,
    G3_n_spl_,
    g67_n_spl_
  );


  or

  (
    g69_n,
    G4_n_spl_00,
    g68_n_spl_
  );


  and

  (
    g70_p,
    G1_p_spl_0,
    G5_p
  );


  or

  (
    g70_n,
    G1_n_spl_0,
    G5_n
  );


  and

  (
    g71_p,
    G3_p,
    g70_p_spl_
  );


  or

  (
    g71_n,
    G3_n_spl_,
    g70_n_spl_
  );


  and

  (
    g72_p,
    G4_p_spl_00,
    g71_p
  );


  or

  (
    g72_n,
    G4_n_spl_00,
    g71_n
  );


  and

  (
    g73_p,
    g65_n_spl_0,
    g72_p
  );


  and

  (
    g74_p,
    G11_p_spl_,
    G16_p_spl_
  );


  or

  (
    g74_n,
    G11_n_spl_0,
    G16_n_spl_
  );


  and

  (
    g75_p,
    G17_p_spl_,
    g74_p_spl_
  );


  or

  (
    g76_n,
    G7_n_spl_,
    G11_n_spl_0
  );


  or

  (
    g77_n,
    G17_n_spl_0,
    g76_n_spl_
  );


  or

  (
    g78_n,
    G8_n_spl_01,
    g76_n_spl_
  );


  or

  (
    g79_n,
    G20_p,
    G21_p
  );


  and

  (
    g80_p,
    G23_p,
    g79_n_spl_
  );


  or

  (
    g81_n,
    g65_n_spl_0,
    g72_n
  );


  and

  (
    g82_p,
    G9_p_spl_0,
    g70_p_spl_
  );


  or

  (
    g82_n,
    G9_n_spl_0,
    g70_n_spl_
  );


  or

  (
    g83_n,
    G10_n_spl_0,
    g68_n_spl_
  );


  or

  (
    g84_n,
    G6_n_spl_,
    g83_n_spl_0
  );


  or

  (
    g85_n,
    G12_n_spl_,
    g84_n
  );


  or

  (
    g86_n,
    G11_n_spl_1,
    G12_n_spl_
  );


  or

  (
    g87_n,
    G15_n,
    g83_n_spl_0
  );


  or

  (
    g88_n,
    g86_n_spl_,
    g87_n
  );


  and

  (
    g89_p,
    G22_p,
    g79_n_spl_
  );


  and

  (
    g90_p,
    G24_p_spl_0,
    G25_n_spl_0
  );


  or

  (
    g90_n,
    G24_n_spl_0,
    G25_p_spl_0
  );


  and

  (
    g91_p,
    G24_n_spl_0,
    G25_p_spl_0
  );


  or

  (
    g91_n,
    G24_p_spl_0,
    G25_n_spl_0
  );


  and

  (
    g92_p,
    g90_n,
    g91_n
  );


  or

  (
    g92_n,
    g90_p,
    g91_p
  );


  and

  (
    g93_p,
    G26_p_spl_0,
    G27_n_spl_0
  );


  or

  (
    g93_n,
    G26_n_spl_0,
    G27_p_spl_0
  );


  and

  (
    g94_p,
    G26_n_spl_0,
    G27_p_spl_0
  );


  or

  (
    g94_n,
    G26_p_spl_0,
    G27_n_spl_0
  );


  and

  (
    g95_p,
    g93_n,
    g94_n
  );


  or

  (
    g95_n,
    g93_p,
    g94_p
  );


  and

  (
    g96_p,
    g92_p_spl_,
    g95_p_spl_
  );


  or

  (
    g96_n,
    g92_n_spl_,
    g95_n_spl_
  );


  and

  (
    g97_p,
    g92_n_spl_,
    g95_n_spl_
  );


  or

  (
    g97_n,
    g92_p_spl_,
    g95_p_spl_
  );


  and

  (
    g98_p,
    g96_n,
    g97_n
  );


  or

  (
    g98_n,
    g96_p,
    g97_p
  );


  and

  (
    g99_p,
    G32_p_spl_0,
    g98_p_spl_
  );


  or

  (
    g99_n,
    G32_n_spl_0,
    g98_n_spl_
  );


  and

  (
    g100_p,
    G32_n_spl_0,
    g98_n_spl_
  );


  or

  (
    g100_n,
    G32_p_spl_0,
    g98_p_spl_
  );


  and

  (
    g101_p,
    g99_n,
    g100_n
  );


  or

  (
    g101_n,
    g99_p,
    g100_p
  );


  and

  (
    g102_p,
    G28_p_spl_0,
    G29_n_spl_0
  );


  or

  (
    g102_n,
    G28_n_spl_0,
    G29_p_spl_0
  );


  and

  (
    g103_p,
    G28_n_spl_0,
    G29_p_spl_0
  );


  or

  (
    g103_n,
    G28_p_spl_0,
    G29_n_spl_0
  );


  and

  (
    g104_p,
    g102_n,
    g103_n
  );


  or

  (
    g104_n,
    g102_p,
    g103_p
  );


  and

  (
    g105_p,
    G30_p_spl_0,
    G31_n_spl_0
  );


  or

  (
    g105_n,
    G30_n_spl_0,
    G31_p_spl_0
  );


  and

  (
    g106_p,
    G30_n_spl_0,
    G31_p_spl_0
  );


  or

  (
    g106_n,
    G30_p_spl_0,
    G31_n_spl_0
  );


  and

  (
    g107_p,
    g105_n,
    g106_n
  );


  or

  (
    g107_n,
    g105_p,
    g106_p
  );


  and

  (
    g108_p,
    g104_p_spl_,
    g107_p_spl_
  );


  or

  (
    g108_n,
    g104_n_spl_,
    g107_n_spl_
  );


  and

  (
    g109_p,
    g104_n_spl_,
    g107_n_spl_
  );


  or

  (
    g109_n,
    g104_p_spl_,
    g107_p_spl_
  );


  and

  (
    g110_p,
    g108_n,
    g109_n
  );


  or

  (
    g110_n,
    g108_p,
    g109_p
  );


  and

  (
    g111_p,
    G33_p_spl_,
    g110_p_spl_
  );


  or

  (
    g111_n,
    G33_n_spl_,
    g110_n_spl_
  );


  and

  (
    g112_p,
    G33_n_spl_,
    g110_n_spl_
  );


  or

  (
    g112_n,
    G33_p_spl_,
    g110_p_spl_
  );


  and

  (
    g113_p,
    g111_n,
    g112_n
  );


  or

  (
    g113_n,
    g111_p,
    g112_p
  );


  and

  (
    g114_p,
    g101_n,
    g113_n
  );


  and

  (
    g115_p,
    g101_p,
    g113_p
  );


  or

  (
    g116_n,
    g114_p,
    g115_p
  );


  and

  (
    g117_p,
    G41_p_spl_0,
    G42_n_spl_00
  );


  or

  (
    g117_n,
    G41_n_spl_00,
    G42_p_spl_0
  );


  and

  (
    g118_p,
    G41_n_spl_00,
    G42_p_spl_0
  );


  or

  (
    g118_n,
    G41_p_spl_0,
    G42_n_spl_00
  );


  and

  (
    g119_p,
    g117_n,
    g118_n
  );


  or

  (
    g119_n,
    g117_p,
    g118_p
  );


  and

  (
    g120_p,
    G43_p_spl_0,
    G44_n_spl_00
  );


  or

  (
    g120_n,
    G43_n_spl_00,
    G44_p_spl_0
  );


  and

  (
    g121_p,
    G43_n_spl_00,
    G44_p_spl_0
  );


  or

  (
    g121_n,
    G43_p_spl_0,
    G44_n_spl_00
  );


  and

  (
    g122_p,
    g120_n,
    g121_n
  );


  or

  (
    g122_n,
    g120_p,
    g121_p
  );


  and

  (
    g123_p,
    g119_p_spl_,
    g122_p_spl_
  );


  or

  (
    g123_n,
    g119_n_spl_,
    g122_n_spl_
  );


  and

  (
    g124_p,
    g119_n_spl_,
    g122_n_spl_
  );


  or

  (
    g124_n,
    g119_p_spl_,
    g122_p_spl_
  );


  and

  (
    g125_p,
    g123_n,
    g124_n
  );


  or

  (
    g125_n,
    g123_p,
    g124_p
  );


  and

  (
    g126_p,
    G32_p_spl_1,
    g125_p_spl_
  );


  or

  (
    g126_n,
    G32_n_spl_1,
    g125_n_spl_
  );


  and

  (
    g127_p,
    G32_n_spl_1,
    g125_n_spl_
  );


  or

  (
    g127_n,
    G32_p_spl_1,
    g125_p_spl_
  );


  and

  (
    g128_p,
    g126_n,
    g127_n
  );


  or

  (
    g128_n,
    g126_p,
    g127_p
  );


  and

  (
    g129_p,
    G45_p_spl_0,
    G46_n_spl_00
  );


  or

  (
    g129_n,
    G45_n_spl_00,
    G46_p_spl_0
  );


  and

  (
    g130_p,
    G45_n_spl_00,
    G46_p_spl_0
  );


  or

  (
    g130_n,
    G45_p_spl_0,
    G46_n_spl_00
  );


  and

  (
    g131_p,
    g129_n,
    g130_n
  );


  or

  (
    g131_n,
    g129_p,
    g130_p
  );


  and

  (
    g132_p,
    G47_p_spl_0,
    G48_n_spl_00
  );


  or

  (
    g132_n,
    G47_n_spl_00,
    G48_p_spl_0
  );


  and

  (
    g133_p,
    G47_n_spl_00,
    G48_p_spl_0
  );


  or

  (
    g133_n,
    G47_p_spl_0,
    G48_n_spl_00
  );


  and

  (
    g134_p,
    g132_n,
    g133_n
  );


  or

  (
    g134_n,
    g132_p,
    g133_p
  );


  and

  (
    g135_p,
    g131_p_spl_,
    g134_p_spl_
  );


  or

  (
    g135_n,
    g131_n_spl_,
    g134_n_spl_
  );


  and

  (
    g136_p,
    g131_n_spl_,
    g134_n_spl_
  );


  or

  (
    g136_n,
    g131_p_spl_,
    g134_p_spl_
  );


  and

  (
    g137_p,
    g135_n,
    g136_n
  );


  or

  (
    g137_n,
    g135_p,
    g136_p
  );


  and

  (
    g138_p,
    G49_p_spl_,
    g137_p_spl_
  );


  or

  (
    g138_n,
    G49_n_spl_,
    g137_n_spl_
  );


  and

  (
    g139_p,
    G49_n_spl_,
    g137_n_spl_
  );


  or

  (
    g139_n,
    G49_p_spl_,
    g137_p_spl_
  );


  and

  (
    g140_p,
    g138_n,
    g139_n
  );


  or

  (
    g140_n,
    g138_p,
    g139_p
  );


  and

  (
    g141_p,
    g128_n,
    g140_n
  );


  and

  (
    g142_p,
    g128_p,
    g140_p
  );


  or

  (
    g143_n,
    g141_p,
    g142_p
  );


  or

  (
    g144_n,
    G55_n_spl_0,
    G59_n
  );


  or

  (
    g145_n,
    G30_n_spl_1,
    G50_n_spl_00
  );


  and

  (
    g146_p,
    G17_p_spl_,
    g82_p_spl_0
  );


  or

  (
    g146_n,
    G17_n_spl_,
    g82_n_spl_0
  );


  and

  (
    g147_p,
    g61_p,
    g146_p
  );


  or

  (
    g147_n,
    g61_n_spl_,
    g146_n
  );


  and

  (
    g148_p,
    G10_p_spl_,
    g147_p_spl_
  );


  or

  (
    g148_n,
    G10_n_spl_0,
    g147_n_spl_
  );


  and

  (
    g149_p,
    G60_n_spl_0,
    g148_p
  );


  or

  (
    g149_n,
    G60_p_spl_,
    g148_n
  );


  and

  (
    g150_p,
    G4_n_spl_01,
    G8_n_spl_01
  );


  or

  (
    g150_n,
    G4_p_spl_00,
    G8_p_spl_0
  );


  and

  (
    g151_p,
    G4_p_spl_01,
    G8_p_spl_0
  );


  or

  (
    g151_n,
    G4_n_spl_01,
    G8_n_spl_10
  );


  and

  (
    g152_p,
    g150_n,
    g151_n
  );


  or

  (
    g152_n,
    g150_p,
    g151_p
  );


  and

  (
    g153_p,
    G11_p_spl_,
    G40_p
  );


  or

  (
    g153_n,
    G11_n_spl_1,
    G40_n
  );


  and

  (
    g154_p,
    g82_p_spl_0,
    g153_p_spl_
  );


  or

  (
    g154_n,
    g82_n_spl_0,
    g153_n_spl_
  );


  and

  (
    g155_p,
    g152_p,
    g154_p
  );


  or

  (
    g155_n,
    g152_n,
    g154_n
  );


  and

  (
    g156_p,
    G4_p_spl_01,
    g67_p
  );


  or

  (
    g156_n,
    G4_n_spl_10,
    g67_n_spl_
  );


  and

  (
    g157_p,
    G8_p_spl_,
    g74_p_spl_
  );


  or

  (
    g157_n,
    G8_n_spl_10,
    g74_n
  );


  and

  (
    g158_p,
    G9_p_spl_0,
    g157_n
  );


  or

  (
    g158_n,
    G9_n_spl_0,
    g157_p
  );


  and

  (
    g159_p,
    g156_p,
    g158_p
  );


  or

  (
    g159_n,
    g156_n,
    g158_n
  );


  and

  (
    g160_p,
    g155_n,
    g159_n
  );


  or

  (
    g160_n,
    g155_p,
    g159_p
  );


  and

  (
    g161_p,
    G31_p_spl_,
    g160_n_spl_00
  );


  or

  (
    g161_n,
    G31_n_spl_,
    g160_p_spl_00
  );


  and

  (
    g162_p,
    g82_p_spl_,
    g153_n_spl_
  );


  or

  (
    g162_n,
    g82_n_spl_1,
    g153_p_spl_
  );


  and

  (
    g163_p,
    G4_p_spl_10,
    g162_p_spl_
  );


  or

  (
    g163_n,
    G4_n_spl_10,
    g162_n_spl_
  );


  and

  (
    g164_p,
    G1_p_spl_,
    g163_n
  );


  or

  (
    g164_n,
    G1_n_spl_,
    g163_p
  );


  and

  (
    g165_p,
    G39_p_spl_,
    g164_n_spl_0
  );


  or

  (
    g165_n,
    G39_n_spl_,
    g164_p_spl_0
  );


  and

  (
    g166_p,
    g161_n,
    g165_n
  );


  or

  (
    g166_n,
    g161_p,
    g165_p
  );


  and

  (
    g167_p,
    g149_n_spl_0,
    g166_p
  );


  or

  (
    g167_n,
    g149_p_spl_0,
    g166_n
  );


  or

  (
    g168_n,
    G54_n_spl_00,
    g167_p_spl_0
  );


  or

  (
    g169_n,
    G8_n_spl_1,
    g83_n_spl_
  );


  or

  (
    g170_n,
    G13_n,
    g86_n_spl_
  );


  or

  (
    g171_n,
    G14_n,
    g170_n
  );


  or

  (
    g172_n,
    g169_n,
    g171_n
  );


  or

  (
    g173_n,
    G48_n_spl_0,
    g172_n_spl_00
  );


  and

  (
    g174_p,
    G48_p_spl_1,
    g167_n_spl_
  );


  or

  (
    g174_n,
    G48_n_spl_1,
    g167_p_spl_0
  );


  and

  (
    g175_p,
    G53_n_spl_00,
    g174_p_spl_
  );


  and

  (
    g176_p,
    G48_n_spl_1,
    g167_p_spl_
  );


  or

  (
    g176_n,
    G48_p_spl_1,
    g167_n_spl_
  );


  or

  (
    g177_n,
    g175_p,
    g176_p_spl_
  );


  or

  (
    g178_n,
    G51_n_spl_000,
    G58_n_spl_
  );


  and

  (
    g179_p,
    g177_n,
    g178_n
  );


  and

  (
    g180_p,
    G58_p,
    g176_n
  );


  or

  (
    g180_n,
    G58_n_spl_,
    g176_p_spl_
  );


  or

  (
    g181_n,
    G51_n_spl_000,
    g180_p_spl_
  );


  and

  (
    g182_p,
    G52_n_spl_00,
    g181_n
  );


  and

  (
    g183_p,
    g174_n_spl_,
    g182_p
  );


  or

  (
    g184_n,
    g179_p,
    g183_p
  );


  and

  (
    g185_p,
    g173_n,
    g184_n
  );


  and

  (
    g186_p,
    g168_n,
    g185_p
  );


  and

  (
    g187_p,
    g145_n,
    g186_p
  );


  and

  (
    g188_p,
    g144_n,
    g187_p
  );


  or

  (
    g189_n,
    G27_n_spl_1,
    G50_n_spl_00
  );


  or

  (
    g190_n,
    G45_n_spl_0,
    g172_n_spl_00
  );


  and

  (
    g191_p,
    G28_p_spl_,
    g160_n_spl_00
  );


  or

  (
    g191_n,
    G28_n_spl_1,
    g160_p_spl_00
  );


  and

  (
    g192_p,
    G35_p_spl_,
    g164_n_spl_0
  );


  or

  (
    g192_n,
    G35_n_spl_,
    g164_p_spl_0
  );


  and

  (
    g193_p,
    g191_n,
    g192_n
  );


  or

  (
    g193_n,
    g191_p,
    g192_p
  );


  and

  (
    g194_p,
    g149_n_spl_0,
    g193_p
  );


  or

  (
    g194_n,
    g149_p_spl_0,
    g193_n
  );


  or

  (
    g195_n,
    G54_n_spl_00,
    g194_p_spl_0
  );


  and

  (
    g196_p,
    G29_p_spl_,
    g160_n_spl_01
  );


  or

  (
    g196_n,
    G29_n_spl_1,
    g160_p_spl_01
  );


  and

  (
    g197_p,
    G36_p_spl_,
    g164_n_spl_1
  );


  or

  (
    g197_n,
    G36_n_spl_,
    g164_p_spl_1
  );


  and

  (
    g198_p,
    g196_n,
    g197_n
  );


  or

  (
    g198_n,
    g196_p,
    g197_p
  );


  and

  (
    g199_p,
    g149_n_spl_1,
    g198_p
  );


  or

  (
    g199_n,
    g149_p_spl_1,
    g198_n
  );


  and

  (
    g200_p,
    G46_p_spl_1,
    g199_n_spl_
  );


  or

  (
    g200_n,
    G46_n_spl_0,
    g199_p_spl_0
  );


  and

  (
    g201_p,
    G46_n_spl_1,
    g199_p_spl_0
  );


  or

  (
    g201_n,
    G46_p_spl_1,
    g199_n_spl_
  );


  and

  (
    g202_p,
    G30_p_spl_,
    g160_n_spl_01
  );


  or

  (
    g202_n,
    G30_n_spl_1,
    g160_p_spl_01
  );


  and

  (
    g203_p,
    G37_p_spl_,
    g164_n_spl_1
  );


  or

  (
    g203_n,
    G37_n_spl_,
    g164_p_spl_1
  );


  and

  (
    g204_p,
    g202_n,
    g203_n
  );


  or

  (
    g204_n,
    g202_p,
    g203_p
  );


  and

  (
    g205_p,
    g149_n_spl_1,
    g204_p
  );


  or

  (
    g205_n,
    g149_p_spl_1,
    g204_n
  );


  and

  (
    g206_p,
    G47_p_spl_1,
    g205_n_spl_
  );


  or

  (
    g206_n,
    G47_n_spl_0,
    g205_p_spl_0
  );


  and

  (
    g207_p,
    G47_n_spl_1,
    g205_p_spl_0
  );


  or

  (
    g207_n,
    G47_p_spl_1,
    g205_n_spl_
  );


  and

  (
    g208_p,
    g174_n_spl_,
    g180_n
  );


  or

  (
    g208_n,
    g174_p_spl_,
    g180_p_spl_
  );


  and

  (
    g209_p,
    g207_n,
    g208_n
  );


  or

  (
    g209_n,
    g207_p_spl_,
    g208_p_spl_
  );


  and

  (
    g210_p,
    g206_n_spl_,
    g209_n
  );


  or

  (
    g210_n,
    g206_p_spl_,
    g209_p_spl_
  );


  and

  (
    g211_p,
    g201_n,
    g210_n
  );


  or

  (
    g211_n,
    g201_p_spl_,
    g210_p_spl_
  );


  and

  (
    g212_p,
    g200_n_spl_,
    g211_n
  );


  or

  (
    g212_n,
    g200_p_spl_,
    g211_p_spl_
  );


  or

  (
    g213_n,
    G51_n_spl_001,
    g212_p_spl_
  );


  and

  (
    g214_p,
    G45_p_spl_1,
    g194_n_spl_
  );


  or

  (
    g214_n,
    G45_n_spl_1,
    g194_p_spl_0
  );


  and

  (
    g215_p,
    G53_n_spl_00,
    g214_p_spl_
  );


  and

  (
    g216_p,
    G45_n_spl_1,
    g194_p_spl_
  );


  or

  (
    g216_n,
    G45_p_spl_1,
    g194_n_spl_
  );


  or

  (
    g217_n,
    g215_p,
    g216_p_spl_
  );


  and

  (
    g218_p,
    g213_n,
    g217_n
  );


  and

  (
    g219_p,
    g212_n,
    g216_n
  );


  or

  (
    g219_n,
    g212_p_spl_,
    g216_p_spl_
  );


  or

  (
    g220_n,
    G51_n_spl_001,
    g219_p_spl_
  );


  and

  (
    g221_p,
    G52_n_spl_00,
    g220_n
  );


  and

  (
    g222_p,
    g214_n_spl_,
    g221_p
  );


  or

  (
    g223_n,
    g218_p,
    g222_p
  );


  and

  (
    g224_p,
    g195_n,
    g223_n
  );


  and

  (
    g225_p,
    g190_n,
    g224_p
  );


  and

  (
    g226_p,
    g189_n,
    g225_p
  );


  or

  (
    g227_n,
    G46_n_spl_1,
    g172_n_spl_01
  );


  or

  (
    g228_n,
    G55_n_spl_0,
    G56_n
  );


  or

  (
    g229_n,
    G28_n_spl_1,
    G50_n_spl_01
  );


  or

  (
    g230_n,
    G54_n_spl_01,
    g199_p_spl_
  );


  and

  (
    g231_p,
    G53_n_spl_01,
    g200_p_spl_
  );


  or

  (
    g232_n,
    g201_p_spl_,
    g231_p
  );


  or

  (
    g233_n,
    G51_n_spl_010,
    g210_p_spl_
  );


  and

  (
    g234_p,
    g232_n,
    g233_n
  );


  or

  (
    g235_n,
    G51_n_spl_010,
    g211_p_spl_
  );


  and

  (
    g236_p,
    G52_n_spl_01,
    g235_n
  );


  and

  (
    g237_p,
    g200_n_spl_,
    g236_p
  );


  or

  (
    g238_n,
    g234_p,
    g237_p
  );


  and

  (
    g239_p,
    g230_n,
    g238_n
  );


  and

  (
    g240_p,
    g229_n,
    g239_p
  );


  and

  (
    g241_p,
    g228_n,
    g240_p
  );


  and

  (
    g242_p,
    g227_n,
    g241_p
  );


  or

  (
    g243_n,
    G55_n_spl_,
    G57_n
  );


  or

  (
    g244_n,
    G29_n_spl_1,
    G50_n_spl_01
  );


  or

  (
    g245_n,
    G54_n_spl_01,
    g205_p_spl_
  );


  or

  (
    g246_n,
    G47_n_spl_1,
    g172_n_spl_01
  );


  and

  (
    g247_p,
    G53_n_spl_01,
    g206_p_spl_
  );


  or

  (
    g248_n,
    g207_p_spl_,
    g247_p
  );


  or

  (
    g249_n,
    G51_n_spl_011,
    g208_p_spl_
  );


  and

  (
    g250_p,
    g248_n,
    g249_n
  );


  or

  (
    g251_n,
    G51_n_spl_011,
    g209_p_spl_
  );


  and

  (
    g252_p,
    G52_n_spl_01,
    g251_n
  );


  and

  (
    g253_p,
    g206_n_spl_,
    g252_p
  );


  or

  (
    g254_n,
    g250_p,
    g253_p
  );


  and

  (
    g255_p,
    g246_n,
    g254_n
  );


  and

  (
    g256_p,
    g245_n,
    g255_p
  );


  and

  (
    g257_p,
    g244_n,
    g256_p
  );


  and

  (
    g258_p,
    g243_n,
    g257_p
  );


  and

  (
    g259_p,
    G10_p_spl_,
    g162_p_spl_
  );


  or

  (
    g259_n,
    G10_n_spl_,
    g162_n_spl_
  );


  and

  (
    g260_p,
    G35_p_spl_,
    g259_p_spl_0
  );


  or

  (
    g260_n,
    G35_n_spl_,
    g259_n_spl_0
  );


  and

  (
    g261_p,
    G2_p_spl_,
    G34_p_spl_0
  );


  or

  (
    g261_n,
    G2_n_spl_,
    G34_n_spl_0
  );


  and

  (
    g262_p,
    g260_n,
    g261_n
  );


  or

  (
    g262_n,
    g260_p,
    g261_p
  );


  and

  (
    g263_p,
    G24_p_spl_,
    g160_n_spl_10
  );


  or

  (
    g263_n,
    G24_n_spl_1,
    g160_p_spl_10
  );


  and

  (
    g264_p,
    G4_p_spl_10,
    g147_p_spl_
  );


  or

  (
    g264_n,
    G4_n_spl_11,
    g147_n_spl_
  );


  and

  (
    g265_p,
    G60_n_spl_0,
    g264_p
  );


  or

  (
    g265_n,
    G60_p_spl_,
    g264_n
  );


  and

  (
    g266_p,
    g263_n,
    g265_n_spl_0
  );


  or

  (
    g266_n,
    g263_p,
    g265_p_spl_0
  );


  and

  (
    g267_p,
    g262_p,
    g266_p
  );


  or

  (
    g267_n,
    g262_n,
    g266_n
  );


  and

  (
    g268_p,
    G41_p_spl_1,
    g267_n_spl_
  );


  or

  (
    g268_n,
    G41_n_spl_0,
    g267_p_spl_0
  );


  and

  (
    g269_p,
    G36_p_spl_,
    g259_p_spl_0
  );


  or

  (
    g269_n,
    G36_n_spl_,
    g259_n_spl_0
  );


  and

  (
    g270_p,
    G9_p_spl_,
    G34_p_spl_0
  );


  or

  (
    g270_n,
    G9_n_spl_,
    G34_n_spl_0
  );


  and

  (
    g271_p,
    g269_n,
    g270_n
  );


  or

  (
    g271_n,
    g269_p,
    g270_p
  );


  and

  (
    g272_p,
    G25_p_spl_,
    g160_n_spl_10
  );


  or

  (
    g272_n,
    G25_n_spl_1,
    g160_p_spl_10
  );


  and

  (
    g273_p,
    g265_n_spl_0,
    g272_n
  );


  or

  (
    g273_n,
    g265_p_spl_0,
    g272_p
  );


  and

  (
    g274_p,
    g271_p,
    g273_p
  );


  or

  (
    g274_n,
    g271_n,
    g273_n
  );


  and

  (
    g275_p,
    G42_p_spl_1,
    g274_n_spl_
  );


  or

  (
    g275_n,
    G42_n_spl_0,
    g274_p_spl_0
  );


  and

  (
    g276_p,
    G42_n_spl_1,
    g274_p_spl_0
  );


  or

  (
    g276_n,
    G42_p_spl_1,
    g274_n_spl_
  );


  and

  (
    g277_p,
    G37_p_spl_,
    g259_p_spl_1
  );


  or

  (
    g277_n,
    G37_n_spl_,
    g259_n_spl_1
  );


  and

  (
    g278_p,
    G4_p_spl_1,
    G34_p_spl_1
  );


  or

  (
    g278_n,
    G4_n_spl_11,
    G34_n_spl_1
  );


  and

  (
    g279_p,
    g277_n,
    g278_n
  );


  or

  (
    g279_n,
    g277_p,
    g278_p
  );


  and

  (
    g280_p,
    G26_p_spl_,
    g160_n_spl_11
  );


  or

  (
    g280_n,
    G26_n_spl_1,
    g160_p_spl_11
  );


  and

  (
    g281_p,
    g265_n_spl_1,
    g280_n
  );


  or

  (
    g281_n,
    g265_p_spl_1,
    g280_p
  );


  and

  (
    g282_p,
    g279_p,
    g281_p
  );


  or

  (
    g282_n,
    g279_n,
    g281_n
  );


  and

  (
    g283_p,
    G43_p_spl_1,
    g282_n_spl_
  );


  or

  (
    g283_n,
    G43_n_spl_0,
    g282_p_spl_0
  );


  and

  (
    g284_p,
    G43_n_spl_1,
    g282_p_spl_0
  );


  or

  (
    g284_n,
    G43_p_spl_1,
    g282_n_spl_
  );


  and

  (
    g285_p,
    g214_n_spl_,
    g219_n
  );


  or

  (
    g285_n,
    g214_p_spl_,
    g219_p_spl_
  );


  and

  (
    g286_p,
    G39_p_spl_,
    g259_p_spl_1
  );


  or

  (
    g286_n,
    G39_n_spl_,
    g259_n_spl_1
  );


  and

  (
    g287_p,
    G34_p_spl_1,
    G38_p
  );


  or

  (
    g287_n,
    G34_n_spl_1,
    G38_n
  );


  and

  (
    g288_p,
    g286_n,
    g287_n
  );


  or

  (
    g288_n,
    g286_p,
    g287_p
  );


  and

  (
    g289_p,
    G27_p_spl_,
    g160_n_spl_11
  );


  or

  (
    g289_n,
    G27_n_spl_1,
    g160_p_spl_11
  );


  and

  (
    g290_p,
    g265_n_spl_1,
    g289_n
  );


  or

  (
    g290_n,
    g265_p_spl_1,
    g289_p
  );


  and

  (
    g291_p,
    g288_p,
    g290_p
  );


  or

  (
    g291_n,
    g288_n,
    g290_n
  );


  and

  (
    g292_p,
    G44_n_spl_0,
    g291_p_spl_0
  );


  or

  (
    g292_n,
    G44_p_spl_1,
    g291_n_spl_
  );


  and

  (
    g293_p,
    g285_n_spl_,
    g292_n_spl_
  );


  or

  (
    g293_n,
    g285_p_spl_,
    g292_p_spl_
  );


  and

  (
    g294_p,
    G44_p_spl_1,
    g291_n_spl_
  );


  or

  (
    g294_n,
    G44_n_spl_1,
    g291_p_spl_0
  );


  and

  (
    g295_p,
    g293_n,
    g294_n_spl_0
  );


  or

  (
    g295_n,
    g293_p,
    g294_p_spl_
  );


  and

  (
    g296_p,
    g284_n_spl_,
    g295_n_spl_
  );


  or

  (
    g296_n,
    g284_p_spl_,
    g295_p_spl_
  );


  and

  (
    g297_p,
    g283_n_spl_0,
    g296_n
  );


  or

  (
    g297_n,
    g283_p_spl_,
    g296_p
  );


  and

  (
    g298_p,
    g276_n_spl_,
    g297_n_spl_
  );


  or

  (
    g298_n,
    g276_p_spl_,
    g297_p_spl_
  );


  and

  (
    g299_p,
    g275_n_spl_0,
    g298_n
  );


  or

  (
    g299_n,
    g275_p_spl_,
    g298_p
  );


  and

  (
    g300_p,
    G41_n_spl_1,
    g267_p_spl_0
  );


  or

  (
    g300_n,
    G41_p_spl_1,
    g267_n_spl_
  );


  or

  (
    g301_n,
    g299_p_spl_,
    g300_p_spl_
  );


  and

  (
    g302_p,
    g268_n_spl_0,
    g301_n
  );


  and

  (
    g303_p,
    g292_n_spl_,
    g294_n_spl_0
  );


  or

  (
    g303_n,
    g292_p_spl_,
    g294_p_spl_
  );


  or

  (
    g304_n,
    g285_p_spl_,
    g303_p
  );


  or

  (
    g305_n,
    g285_n_spl_,
    g303_n_spl_
  );


  and

  (
    g306_p,
    g304_n,
    g305_n
  );


  or

  (
    g307_n,
    G51_n_spl_10,
    g306_p
  );


  or

  (
    g308_n,
    G52_n_spl_10,
    g303_n_spl_
  );


  or

  (
    g309_n,
    G54_n_spl_10,
    g291_p_spl_
  );


  and

  (
    g310_p,
    g308_n,
    g309_n
  );


  or

  (
    g311_n,
    G44_n_spl_1,
    g172_n_spl_10
  );


  or

  (
    g312_n,
    G53_n_spl_10,
    g294_n_spl_
  );


  or

  (
    g313_n,
    G26_n_spl_1,
    G50_n_spl_10
  );


  and

  (
    g314_p,
    g312_n,
    g313_n
  );


  and

  (
    g315_p,
    g311_n,
    g314_p
  );


  and

  (
    g316_p,
    g310_p,
    g315_p
  );


  and

  (
    g317_p,
    g307_n,
    g316_p
  );


  or

  (
    g318_n,
    G53_n_spl_10,
    g268_n_spl_0
  );


  or

  (
    g319_n,
    G50_n_spl_10,
    G60_n_spl_
  );


  and

  (
    g320_p,
    g318_n,
    g319_n
  );


  or

  (
    g321_n,
    G41_n_spl_1,
    g172_n_spl_10
  );


  and

  (
    g322_p,
    g268_n_spl_,
    g300_n
  );


  or

  (
    g322_n,
    g268_p,
    g300_p_spl_
  );


  or

  (
    g323_n,
    G52_n_spl_10,
    g322_n_spl_
  );


  or

  (
    g324_n,
    G54_n_spl_10,
    g267_p_spl_
  );


  and

  (
    g325_p,
    g323_n,
    g324_n
  );


  and

  (
    g326_p,
    g321_n,
    g325_p
  );


  and

  (
    g327_p,
    g320_p,
    g326_p
  );


  and

  (
    g328_p,
    g299_p_spl_,
    g322_n_spl_
  );


  and

  (
    g329_p,
    g299_n,
    g322_p
  );


  or

  (
    g330_n,
    G51_n_spl_10,
    g329_p
  );


  or

  (
    g331_n,
    g328_p,
    g330_n
  );


  and

  (
    g332_p,
    g327_p,
    g331_n
  );


  or

  (
    g333_n,
    G53_n_spl_11,
    g275_n_spl_0
  );


  or

  (
    g334_n,
    G24_n_spl_1,
    G50_n_spl_11
  );


  and

  (
    g335_p,
    g333_n,
    g334_n
  );


  or

  (
    g336_n,
    G42_n_spl_1,
    g172_n_spl_11
  );


  and

  (
    g337_p,
    g275_n_spl_,
    g276_n_spl_
  );


  or

  (
    g337_n,
    g275_p_spl_,
    g276_p_spl_
  );


  or

  (
    g338_n,
    G52_n_spl_11,
    g337_n_spl_
  );


  or

  (
    g339_n,
    G54_n_spl_11,
    g274_p_spl_
  );


  and

  (
    g340_p,
    g338_n,
    g339_n
  );


  and

  (
    g341_p,
    g336_n,
    g340_p
  );


  and

  (
    g342_p,
    g335_p,
    g341_p
  );


  and

  (
    g343_p,
    g297_p_spl_,
    g337_n_spl_
  );


  and

  (
    g344_p,
    g297_n_spl_,
    g337_p
  );


  or

  (
    g345_n,
    G51_n_spl_11,
    g344_p
  );


  or

  (
    g346_n,
    g343_p,
    g345_n
  );


  and

  (
    g347_p,
    g342_p,
    g346_n
  );


  or

  (
    g348_n,
    G53_n_spl_11,
    g283_n_spl_0
  );


  or

  (
    g349_n,
    G25_n_spl_1,
    G50_n_spl_11
  );


  and

  (
    g350_p,
    g348_n,
    g349_n
  );


  or

  (
    g351_n,
    G43_n_spl_1,
    g172_n_spl_11
  );


  and

  (
    g352_p,
    g283_n_spl_,
    g284_n_spl_
  );


  or

  (
    g352_n,
    g283_p_spl_,
    g284_p_spl_
  );


  or

  (
    g353_n,
    G52_n_spl_11,
    g352_n_spl_
  );


  or

  (
    g354_n,
    G54_n_spl_11,
    g282_p_spl_
  );


  and

  (
    g355_p,
    g353_n,
    g354_n
  );


  and

  (
    g356_p,
    g351_n,
    g355_p
  );


  and

  (
    g357_p,
    g295_p_spl_,
    g352_n_spl_
  );


  and

  (
    g358_p,
    g295_n_spl_,
    g352_p
  );


  or

  (
    g359_n,
    G51_n_spl_11,
    g358_p
  );


  or

  (
    g360_n,
    g357_p,
    g359_n
  );


  and

  (
    g361_p,
    g356_p,
    g360_n
  );


  and

  (
    g362_p,
    g350_p,
    g361_p
  );


  buf

  (
    G855,
    g62_n
  );


  buf

  (
    G856,
    g64_n
  );


  buf

  (
    G857,
    g65_n_spl_
  );


  buf

  (
    G858,
    g66_n
  );


  buf

  (
    G859,
    g69_n
  );


  buf

  (
    G860,
    g73_p
  );


  buf

  (
    G861,
    g75_p
  );


  not

  (
    G862,
    g77_n
  );


  not

  (
    G863,
    g78_n
  );


  not

  (
    G864,
    g80_p
  );


  not

  (
    G865,
    g81_n
  );


  buf

  (
    G866,
    g82_n_spl_1
  );


  buf

  (
    G867,
    g85_n
  );


  buf

  (
    G868,
    g88_n
  );


  not

  (
    G869,
    g89_p
  );


  buf

  (
    G870,
    g116_n
  );


  buf

  (
    G871,
    g143_n
  );


  buf

  (
    G872,
    g188_p
  );


  buf

  (
    G873,
    g226_p
  );


  buf

  (
    G874,
    g242_p
  );


  buf

  (
    G875,
    g258_p
  );


  buf

  (
    G876,
    g302_p
  );


  buf

  (
    G877,
    g317_p
  );


  buf

  (
    G878,
    g332_p
  );


  buf

  (
    G879,
    g347_p
  );


  buf

  (
    G880,
    g362_p
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    G6_n_spl_,
    G6_n
  );


  buf

  (
    G6_n_spl_0,
    G6_n_spl_
  );


  buf

  (
    G16_n_spl_,
    G16_n
  );


  buf

  (
    G8_n_spl_,
    G8_n
  );


  buf

  (
    G8_n_spl_0,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_00,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_01,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_1,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_10,
    G8_n_spl_1
  );


  buf

  (
    g61_n_spl_,
    g61_n
  );


  buf

  (
    G7_n_spl_,
    G7_n
  );


  buf

  (
    G17_n_spl_,
    G17_n
  );


  buf

  (
    G17_n_spl_0,
    G17_n_spl_
  );


  buf

  (
    g63_n_spl_,
    g63_n
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G1_p_spl_0,
    G1_p_spl_
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G3_n_spl_,
    G3_n
  );


  buf

  (
    g67_n_spl_,
    g67_n
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    G4_n_spl_0,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_00,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_01,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_1,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_10,
    G4_n_spl_1
  );


  buf

  (
    G4_n_spl_11,
    G4_n_spl_1
  );


  buf

  (
    g68_n_spl_,
    g68_n
  );


  buf

  (
    g70_p_spl_,
    g70_p
  );


  buf

  (
    g70_n_spl_,
    g70_n
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_00,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_01,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_10,
    G4_p_spl_1
  );


  buf

  (
    g65_n_spl_,
    g65_n
  );


  buf

  (
    g65_n_spl_0,
    g65_n_spl_
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    G11_n_spl_0,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_1,
    G11_n_spl_
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    g74_p_spl_,
    g74_p
  );


  buf

  (
    g76_n_spl_,
    g76_n
  );


  buf

  (
    g79_n_spl_,
    g79_n
  );


  buf

  (
    G9_p_spl_,
    G9_p
  );


  buf

  (
    G9_p_spl_0,
    G9_p_spl_
  );


  buf

  (
    G9_n_spl_,
    G9_n
  );


  buf

  (
    G9_n_spl_0,
    G9_n_spl_
  );


  buf

  (
    G10_n_spl_,
    G10_n
  );


  buf

  (
    G10_n_spl_0,
    G10_n_spl_
  );


  buf

  (
    g83_n_spl_,
    g83_n
  );


  buf

  (
    g83_n_spl_0,
    g83_n_spl_
  );


  buf

  (
    G12_n_spl_,
    G12_n
  );


  buf

  (
    g86_n_spl_,
    g86_n
  );


  buf

  (
    G24_p_spl_,
    G24_p
  );


  buf

  (
    G24_p_spl_0,
    G24_p_spl_
  );


  buf

  (
    G25_n_spl_,
    G25_n
  );


  buf

  (
    G25_n_spl_0,
    G25_n_spl_
  );


  buf

  (
    G25_n_spl_1,
    G25_n_spl_
  );


  buf

  (
    G24_n_spl_,
    G24_n
  );


  buf

  (
    G24_n_spl_0,
    G24_n_spl_
  );


  buf

  (
    G24_n_spl_1,
    G24_n_spl_
  );


  buf

  (
    G25_p_spl_,
    G25_p
  );


  buf

  (
    G25_p_spl_0,
    G25_p_spl_
  );


  buf

  (
    G26_p_spl_,
    G26_p
  );


  buf

  (
    G26_p_spl_0,
    G26_p_spl_
  );


  buf

  (
    G27_n_spl_,
    G27_n
  );


  buf

  (
    G27_n_spl_0,
    G27_n_spl_
  );


  buf

  (
    G27_n_spl_1,
    G27_n_spl_
  );


  buf

  (
    G26_n_spl_,
    G26_n
  );


  buf

  (
    G26_n_spl_0,
    G26_n_spl_
  );


  buf

  (
    G26_n_spl_1,
    G26_n_spl_
  );


  buf

  (
    G27_p_spl_,
    G27_p
  );


  buf

  (
    G27_p_spl_0,
    G27_p_spl_
  );


  buf

  (
    g92_p_spl_,
    g92_p
  );


  buf

  (
    g95_p_spl_,
    g95_p
  );


  buf

  (
    g92_n_spl_,
    g92_n
  );


  buf

  (
    g95_n_spl_,
    g95_n
  );


  buf

  (
    G32_p_spl_,
    G32_p
  );


  buf

  (
    G32_p_spl_0,
    G32_p_spl_
  );


  buf

  (
    G32_p_spl_1,
    G32_p_spl_
  );


  buf

  (
    g98_p_spl_,
    g98_p
  );


  buf

  (
    G32_n_spl_,
    G32_n
  );


  buf

  (
    G32_n_spl_0,
    G32_n_spl_
  );


  buf

  (
    G32_n_spl_1,
    G32_n_spl_
  );


  buf

  (
    g98_n_spl_,
    g98_n
  );


  buf

  (
    G28_p_spl_,
    G28_p
  );


  buf

  (
    G28_p_spl_0,
    G28_p_spl_
  );


  buf

  (
    G29_n_spl_,
    G29_n
  );


  buf

  (
    G29_n_spl_0,
    G29_n_spl_
  );


  buf

  (
    G29_n_spl_1,
    G29_n_spl_
  );


  buf

  (
    G28_n_spl_,
    G28_n
  );


  buf

  (
    G28_n_spl_0,
    G28_n_spl_
  );


  buf

  (
    G28_n_spl_1,
    G28_n_spl_
  );


  buf

  (
    G29_p_spl_,
    G29_p
  );


  buf

  (
    G29_p_spl_0,
    G29_p_spl_
  );


  buf

  (
    G30_p_spl_,
    G30_p
  );


  buf

  (
    G30_p_spl_0,
    G30_p_spl_
  );


  buf

  (
    G31_n_spl_,
    G31_n
  );


  buf

  (
    G31_n_spl_0,
    G31_n_spl_
  );


  buf

  (
    G30_n_spl_,
    G30_n
  );


  buf

  (
    G30_n_spl_0,
    G30_n_spl_
  );


  buf

  (
    G30_n_spl_1,
    G30_n_spl_
  );


  buf

  (
    G31_p_spl_,
    G31_p
  );


  buf

  (
    G31_p_spl_0,
    G31_p_spl_
  );


  buf

  (
    g104_p_spl_,
    g104_p
  );


  buf

  (
    g107_p_spl_,
    g107_p
  );


  buf

  (
    g104_n_spl_,
    g104_n
  );


  buf

  (
    g107_n_spl_,
    g107_n
  );


  buf

  (
    G33_p_spl_,
    G33_p
  );


  buf

  (
    g110_p_spl_,
    g110_p
  );


  buf

  (
    G33_n_spl_,
    G33_n
  );


  buf

  (
    g110_n_spl_,
    g110_n
  );


  buf

  (
    G41_p_spl_,
    G41_p
  );


  buf

  (
    G41_p_spl_0,
    G41_p_spl_
  );


  buf

  (
    G41_p_spl_1,
    G41_p_spl_
  );


  buf

  (
    G42_n_spl_,
    G42_n
  );


  buf

  (
    G42_n_spl_0,
    G42_n_spl_
  );


  buf

  (
    G42_n_spl_00,
    G42_n_spl_0
  );


  buf

  (
    G42_n_spl_1,
    G42_n_spl_
  );


  buf

  (
    G41_n_spl_,
    G41_n
  );


  buf

  (
    G41_n_spl_0,
    G41_n_spl_
  );


  buf

  (
    G41_n_spl_00,
    G41_n_spl_0
  );


  buf

  (
    G41_n_spl_1,
    G41_n_spl_
  );


  buf

  (
    G42_p_spl_,
    G42_p
  );


  buf

  (
    G42_p_spl_0,
    G42_p_spl_
  );


  buf

  (
    G42_p_spl_1,
    G42_p_spl_
  );


  buf

  (
    G43_p_spl_,
    G43_p
  );


  buf

  (
    G43_p_spl_0,
    G43_p_spl_
  );


  buf

  (
    G43_p_spl_1,
    G43_p_spl_
  );


  buf

  (
    G44_n_spl_,
    G44_n
  );


  buf

  (
    G44_n_spl_0,
    G44_n_spl_
  );


  buf

  (
    G44_n_spl_00,
    G44_n_spl_0
  );


  buf

  (
    G44_n_spl_1,
    G44_n_spl_
  );


  buf

  (
    G43_n_spl_,
    G43_n
  );


  buf

  (
    G43_n_spl_0,
    G43_n_spl_
  );


  buf

  (
    G43_n_spl_00,
    G43_n_spl_0
  );


  buf

  (
    G43_n_spl_1,
    G43_n_spl_
  );


  buf

  (
    G44_p_spl_,
    G44_p
  );


  buf

  (
    G44_p_spl_0,
    G44_p_spl_
  );


  buf

  (
    G44_p_spl_1,
    G44_p_spl_
  );


  buf

  (
    g119_p_spl_,
    g119_p
  );


  buf

  (
    g122_p_spl_,
    g122_p
  );


  buf

  (
    g119_n_spl_,
    g119_n
  );


  buf

  (
    g122_n_spl_,
    g122_n
  );


  buf

  (
    g125_p_spl_,
    g125_p
  );


  buf

  (
    g125_n_spl_,
    g125_n
  );


  buf

  (
    G45_p_spl_,
    G45_p
  );


  buf

  (
    G45_p_spl_0,
    G45_p_spl_
  );


  buf

  (
    G45_p_spl_1,
    G45_p_spl_
  );


  buf

  (
    G46_n_spl_,
    G46_n
  );


  buf

  (
    G46_n_spl_0,
    G46_n_spl_
  );


  buf

  (
    G46_n_spl_00,
    G46_n_spl_0
  );


  buf

  (
    G46_n_spl_1,
    G46_n_spl_
  );


  buf

  (
    G45_n_spl_,
    G45_n
  );


  buf

  (
    G45_n_spl_0,
    G45_n_spl_
  );


  buf

  (
    G45_n_spl_00,
    G45_n_spl_0
  );


  buf

  (
    G45_n_spl_1,
    G45_n_spl_
  );


  buf

  (
    G46_p_spl_,
    G46_p
  );


  buf

  (
    G46_p_spl_0,
    G46_p_spl_
  );


  buf

  (
    G46_p_spl_1,
    G46_p_spl_
  );


  buf

  (
    G47_p_spl_,
    G47_p
  );


  buf

  (
    G47_p_spl_0,
    G47_p_spl_
  );


  buf

  (
    G47_p_spl_1,
    G47_p_spl_
  );


  buf

  (
    G48_n_spl_,
    G48_n
  );


  buf

  (
    G48_n_spl_0,
    G48_n_spl_
  );


  buf

  (
    G48_n_spl_00,
    G48_n_spl_0
  );


  buf

  (
    G48_n_spl_1,
    G48_n_spl_
  );


  buf

  (
    G47_n_spl_,
    G47_n
  );


  buf

  (
    G47_n_spl_0,
    G47_n_spl_
  );


  buf

  (
    G47_n_spl_00,
    G47_n_spl_0
  );


  buf

  (
    G47_n_spl_1,
    G47_n_spl_
  );


  buf

  (
    G48_p_spl_,
    G48_p
  );


  buf

  (
    G48_p_spl_0,
    G48_p_spl_
  );


  buf

  (
    G48_p_spl_1,
    G48_p_spl_
  );


  buf

  (
    g131_p_spl_,
    g131_p
  );


  buf

  (
    g134_p_spl_,
    g134_p
  );


  buf

  (
    g131_n_spl_,
    g131_n
  );


  buf

  (
    g134_n_spl_,
    g134_n
  );


  buf

  (
    G49_p_spl_,
    G49_p
  );


  buf

  (
    g137_p_spl_,
    g137_p
  );


  buf

  (
    G49_n_spl_,
    G49_n
  );


  buf

  (
    g137_n_spl_,
    g137_n
  );


  buf

  (
    G55_n_spl_,
    G55_n
  );


  buf

  (
    G55_n_spl_0,
    G55_n_spl_
  );


  buf

  (
    G50_n_spl_,
    G50_n
  );


  buf

  (
    G50_n_spl_0,
    G50_n_spl_
  );


  buf

  (
    G50_n_spl_00,
    G50_n_spl_0
  );


  buf

  (
    G50_n_spl_01,
    G50_n_spl_0
  );


  buf

  (
    G50_n_spl_1,
    G50_n_spl_
  );


  buf

  (
    G50_n_spl_10,
    G50_n_spl_1
  );


  buf

  (
    G50_n_spl_11,
    G50_n_spl_1
  );


  buf

  (
    g82_p_spl_,
    g82_p
  );


  buf

  (
    g82_p_spl_0,
    g82_p_spl_
  );


  buf

  (
    g82_n_spl_,
    g82_n
  );


  buf

  (
    g82_n_spl_0,
    g82_n_spl_
  );


  buf

  (
    g82_n_spl_1,
    g82_n_spl_
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


  buf

  (
    g147_p_spl_,
    g147_p
  );


  buf

  (
    g147_n_spl_,
    g147_n
  );


  buf

  (
    G60_n_spl_,
    G60_n
  );


  buf

  (
    G60_n_spl_0,
    G60_n_spl_
  );


  buf

  (
    G60_p_spl_,
    G60_p
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    g153_p_spl_,
    g153_p
  );


  buf

  (
    g153_n_spl_,
    g153_n
  );


  buf

  (
    g160_n_spl_,
    g160_n
  );


  buf

  (
    g160_n_spl_0,
    g160_n_spl_
  );


  buf

  (
    g160_n_spl_00,
    g160_n_spl_0
  );


  buf

  (
    g160_n_spl_01,
    g160_n_spl_0
  );


  buf

  (
    g160_n_spl_1,
    g160_n_spl_
  );


  buf

  (
    g160_n_spl_10,
    g160_n_spl_1
  );


  buf

  (
    g160_n_spl_11,
    g160_n_spl_1
  );


  buf

  (
    g160_p_spl_,
    g160_p
  );


  buf

  (
    g160_p_spl_0,
    g160_p_spl_
  );


  buf

  (
    g160_p_spl_00,
    g160_p_spl_0
  );


  buf

  (
    g160_p_spl_01,
    g160_p_spl_0
  );


  buf

  (
    g160_p_spl_1,
    g160_p_spl_
  );


  buf

  (
    g160_p_spl_10,
    g160_p_spl_1
  );


  buf

  (
    g160_p_spl_11,
    g160_p_spl_1
  );


  buf

  (
    g162_p_spl_,
    g162_p
  );


  buf

  (
    g162_n_spl_,
    g162_n
  );


  buf

  (
    G39_p_spl_,
    G39_p
  );


  buf

  (
    g164_n_spl_,
    g164_n
  );


  buf

  (
    g164_n_spl_0,
    g164_n_spl_
  );


  buf

  (
    g164_n_spl_1,
    g164_n_spl_
  );


  buf

  (
    G39_n_spl_,
    G39_n
  );


  buf

  (
    g164_p_spl_,
    g164_p
  );


  buf

  (
    g164_p_spl_0,
    g164_p_spl_
  );


  buf

  (
    g164_p_spl_1,
    g164_p_spl_
  );


  buf

  (
    g149_n_spl_,
    g149_n
  );


  buf

  (
    g149_n_spl_0,
    g149_n_spl_
  );


  buf

  (
    g149_n_spl_1,
    g149_n_spl_
  );


  buf

  (
    g149_p_spl_,
    g149_p
  );


  buf

  (
    g149_p_spl_0,
    g149_p_spl_
  );


  buf

  (
    g149_p_spl_1,
    g149_p_spl_
  );


  buf

  (
    G54_n_spl_,
    G54_n
  );


  buf

  (
    G54_n_spl_0,
    G54_n_spl_
  );


  buf

  (
    G54_n_spl_00,
    G54_n_spl_0
  );


  buf

  (
    G54_n_spl_01,
    G54_n_spl_0
  );


  buf

  (
    G54_n_spl_1,
    G54_n_spl_
  );


  buf

  (
    G54_n_spl_10,
    G54_n_spl_1
  );


  buf

  (
    G54_n_spl_11,
    G54_n_spl_1
  );


  buf

  (
    g167_p_spl_,
    g167_p
  );


  buf

  (
    g167_p_spl_0,
    g167_p_spl_
  );


  buf

  (
    g172_n_spl_,
    g172_n
  );


  buf

  (
    g172_n_spl_0,
    g172_n_spl_
  );


  buf

  (
    g172_n_spl_00,
    g172_n_spl_0
  );


  buf

  (
    g172_n_spl_01,
    g172_n_spl_0
  );


  buf

  (
    g172_n_spl_1,
    g172_n_spl_
  );


  buf

  (
    g172_n_spl_10,
    g172_n_spl_1
  );


  buf

  (
    g172_n_spl_11,
    g172_n_spl_1
  );


  buf

  (
    g167_n_spl_,
    g167_n
  );


  buf

  (
    G53_n_spl_,
    G53_n
  );


  buf

  (
    G53_n_spl_0,
    G53_n_spl_
  );


  buf

  (
    G53_n_spl_00,
    G53_n_spl_0
  );


  buf

  (
    G53_n_spl_01,
    G53_n_spl_0
  );


  buf

  (
    G53_n_spl_1,
    G53_n_spl_
  );


  buf

  (
    G53_n_spl_10,
    G53_n_spl_1
  );


  buf

  (
    G53_n_spl_11,
    G53_n_spl_1
  );


  buf

  (
    g174_p_spl_,
    g174_p
  );


  buf

  (
    g176_p_spl_,
    g176_p
  );


  buf

  (
    G51_n_spl_,
    G51_n
  );


  buf

  (
    G51_n_spl_0,
    G51_n_spl_
  );


  buf

  (
    G51_n_spl_00,
    G51_n_spl_0
  );


  buf

  (
    G51_n_spl_000,
    G51_n_spl_00
  );


  buf

  (
    G51_n_spl_001,
    G51_n_spl_00
  );


  buf

  (
    G51_n_spl_01,
    G51_n_spl_0
  );


  buf

  (
    G51_n_spl_010,
    G51_n_spl_01
  );


  buf

  (
    G51_n_spl_011,
    G51_n_spl_01
  );


  buf

  (
    G51_n_spl_1,
    G51_n_spl_
  );


  buf

  (
    G51_n_spl_10,
    G51_n_spl_1
  );


  buf

  (
    G51_n_spl_11,
    G51_n_spl_1
  );


  buf

  (
    G58_n_spl_,
    G58_n
  );


  buf

  (
    g180_p_spl_,
    g180_p
  );


  buf

  (
    G52_n_spl_,
    G52_n
  );


  buf

  (
    G52_n_spl_0,
    G52_n_spl_
  );


  buf

  (
    G52_n_spl_00,
    G52_n_spl_0
  );


  buf

  (
    G52_n_spl_01,
    G52_n_spl_0
  );


  buf

  (
    G52_n_spl_1,
    G52_n_spl_
  );


  buf

  (
    G52_n_spl_10,
    G52_n_spl_1
  );


  buf

  (
    G52_n_spl_11,
    G52_n_spl_1
  );


  buf

  (
    g174_n_spl_,
    g174_n
  );


  buf

  (
    G35_p_spl_,
    G35_p
  );


  buf

  (
    G35_n_spl_,
    G35_n
  );


  buf

  (
    g194_p_spl_,
    g194_p
  );


  buf

  (
    g194_p_spl_0,
    g194_p_spl_
  );


  buf

  (
    G36_p_spl_,
    G36_p
  );


  buf

  (
    G36_n_spl_,
    G36_n
  );


  buf

  (
    g199_n_spl_,
    g199_n
  );


  buf

  (
    g199_p_spl_,
    g199_p
  );


  buf

  (
    g199_p_spl_0,
    g199_p_spl_
  );


  buf

  (
    G37_p_spl_,
    G37_p
  );


  buf

  (
    G37_n_spl_,
    G37_n
  );


  buf

  (
    g205_n_spl_,
    g205_n
  );


  buf

  (
    g205_p_spl_,
    g205_p
  );


  buf

  (
    g205_p_spl_0,
    g205_p_spl_
  );


  buf

  (
    g207_p_spl_,
    g207_p
  );


  buf

  (
    g208_p_spl_,
    g208_p
  );


  buf

  (
    g206_n_spl_,
    g206_n
  );


  buf

  (
    g206_p_spl_,
    g206_p
  );


  buf

  (
    g209_p_spl_,
    g209_p
  );


  buf

  (
    g201_p_spl_,
    g201_p
  );


  buf

  (
    g210_p_spl_,
    g210_p
  );


  buf

  (
    g200_n_spl_,
    g200_n
  );


  buf

  (
    g200_p_spl_,
    g200_p
  );


  buf

  (
    g211_p_spl_,
    g211_p
  );


  buf

  (
    g212_p_spl_,
    g212_p
  );


  buf

  (
    g194_n_spl_,
    g194_n
  );


  buf

  (
    g214_p_spl_,
    g214_p
  );


  buf

  (
    g216_p_spl_,
    g216_p
  );


  buf

  (
    g219_p_spl_,
    g219_p
  );


  buf

  (
    g214_n_spl_,
    g214_n
  );


  buf

  (
    g259_p_spl_,
    g259_p
  );


  buf

  (
    g259_p_spl_0,
    g259_p_spl_
  );


  buf

  (
    g259_p_spl_1,
    g259_p_spl_
  );


  buf

  (
    g259_n_spl_,
    g259_n
  );


  buf

  (
    g259_n_spl_0,
    g259_n_spl_
  );


  buf

  (
    g259_n_spl_1,
    g259_n_spl_
  );


  buf

  (
    G34_p_spl_,
    G34_p
  );


  buf

  (
    G34_p_spl_0,
    G34_p_spl_
  );


  buf

  (
    G34_p_spl_1,
    G34_p_spl_
  );


  buf

  (
    G34_n_spl_,
    G34_n
  );


  buf

  (
    G34_n_spl_0,
    G34_n_spl_
  );


  buf

  (
    G34_n_spl_1,
    G34_n_spl_
  );


  buf

  (
    g265_n_spl_,
    g265_n
  );


  buf

  (
    g265_n_spl_0,
    g265_n_spl_
  );


  buf

  (
    g265_n_spl_1,
    g265_n_spl_
  );


  buf

  (
    g265_p_spl_,
    g265_p
  );


  buf

  (
    g265_p_spl_0,
    g265_p_spl_
  );


  buf

  (
    g265_p_spl_1,
    g265_p_spl_
  );


  buf

  (
    g267_n_spl_,
    g267_n
  );


  buf

  (
    g267_p_spl_,
    g267_p
  );


  buf

  (
    g267_p_spl_0,
    g267_p_spl_
  );


  buf

  (
    g274_n_spl_,
    g274_n
  );


  buf

  (
    g274_p_spl_,
    g274_p
  );


  buf

  (
    g274_p_spl_0,
    g274_p_spl_
  );


  buf

  (
    g282_n_spl_,
    g282_n
  );


  buf

  (
    g282_p_spl_,
    g282_p
  );


  buf

  (
    g282_p_spl_0,
    g282_p_spl_
  );


  buf

  (
    g291_p_spl_,
    g291_p
  );


  buf

  (
    g291_p_spl_0,
    g291_p_spl_
  );


  buf

  (
    g291_n_spl_,
    g291_n
  );


  buf

  (
    g285_n_spl_,
    g285_n
  );


  buf

  (
    g292_n_spl_,
    g292_n
  );


  buf

  (
    g285_p_spl_,
    g285_p
  );


  buf

  (
    g292_p_spl_,
    g292_p
  );


  buf

  (
    g294_n_spl_,
    g294_n
  );


  buf

  (
    g294_n_spl_0,
    g294_n_spl_
  );


  buf

  (
    g294_p_spl_,
    g294_p
  );


  buf

  (
    g284_n_spl_,
    g284_n
  );


  buf

  (
    g295_n_spl_,
    g295_n
  );


  buf

  (
    g284_p_spl_,
    g284_p
  );


  buf

  (
    g295_p_spl_,
    g295_p
  );


  buf

  (
    g283_n_spl_,
    g283_n
  );


  buf

  (
    g283_n_spl_0,
    g283_n_spl_
  );


  buf

  (
    g283_p_spl_,
    g283_p
  );


  buf

  (
    g276_n_spl_,
    g276_n
  );


  buf

  (
    g297_n_spl_,
    g297_n
  );


  buf

  (
    g276_p_spl_,
    g276_p
  );


  buf

  (
    g297_p_spl_,
    g297_p
  );


  buf

  (
    g275_n_spl_,
    g275_n
  );


  buf

  (
    g275_n_spl_0,
    g275_n_spl_
  );


  buf

  (
    g275_p_spl_,
    g275_p
  );


  buf

  (
    g299_p_spl_,
    g299_p
  );


  buf

  (
    g300_p_spl_,
    g300_p
  );


  buf

  (
    g268_n_spl_,
    g268_n
  );


  buf

  (
    g268_n_spl_0,
    g268_n_spl_
  );


  buf

  (
    g303_n_spl_,
    g303_n
  );


  buf

  (
    g322_n_spl_,
    g322_n
  );


  buf

  (
    g337_n_spl_,
    g337_n
  );


  buf

  (
    g352_n_spl_,
    g352_n
  );


endmodule
