
module mymod
(
  G1_p,
  G1_n,
  G2_p,
  G2_n,
  G3_p,
  G3_n,
  G4_p,
  G4_n,
  G5_p,
  G5_n,
  G6_p,
  G6_n,
  G7_p,
  G7_n,
  G8_p,
  G8_n,
  G9_p,
  G9_n,
  G10_p,
  G10_n,
  G11_p,
  G11_n,
  G12_p,
  G12_n,
  G13_p,
  G13_n,
  G14_p,
  G14_n,
  G15_p,
  G15_n,
  G16_p,
  G16_n,
  G17_p,
  G17_n,
  G18_p,
  G18_n,
  G19_p,
  G19_n,
  G20_p,
  G20_n,
  G21_p,
  G21_n,
  G22_p,
  G22_n,
  G23_p,
  G23_n,
  G24_p,
  G24_n,
  G25_p,
  G25_n,
  G26_p,
  G26_n,
  G27_p,
  G27_n,
  G28_p,
  G28_n,
  G29_p,
  G29_n,
  G30_p,
  G30_n,
  G31_p,
  G31_n,
  G32_p,
  G32_n,
  G33_p,
  G33_n,
  G34_p,
  G34_n,
  G35_p,
  G35_n,
  G36_p,
  G36_n,
  G37_p,
  G37_n,
  G38_p,
  G38_n,
  G39_p,
  G39_n,
  G40_p,
  G40_n,
  G41_p,
  G41_n,
  G42_p,
  G42_n,
  G43_p,
  G43_n,
  G44_p,
  G44_n,
  G45_p,
  G45_n,
  G46_p,
  G46_n,
  G47_p,
  G47_n,
  G48_p,
  G48_n,
  G49_p,
  G49_n,
  G50_p,
  G50_n,
  G51_p,
  G51_n,
  G52_p,
  G52_n,
  G53_p,
  G53_n,
  G54_p,
  G54_n,
  G55_p,
  G55_n,
  G56_p,
  G56_n,
  G57_p,
  G57_n,
  G58_p,
  G58_n,
  G59_p,
  G59_n,
  G60_p,
  G60_n,
  G61_p,
  G61_n,
  G62_p,
  G62_n,
  G63_p,
  G63_n,
  G64_p,
  G64_n,
  G65_p,
  G65_n,
  G66_p,
  G66_n,
  G67_p,
  G67_n,
  G68_p,
  G68_n,
  G69_p,
  G69_n,
  G70_p,
  G70_n,
  G71_p,
  G71_n,
  G72_p,
  G72_n,
  G73_p,
  G73_n,
  G74_p,
  G74_n,
  G75_p,
  G75_n,
  G76_p,
  G76_n,
  G77_p,
  G77_n,
  G78_p,
  G78_n,
  G79_p,
  G79_n,
  G80_p,
  G80_n,
  G81_p,
  G81_n,
  G82_p,
  G82_n,
  G83_p,
  G83_n,
  G84_p,
  G84_n,
  G85_p,
  G85_n,
  G86_p,
  G86_n,
  G87_p,
  G87_n,
  G88_p,
  G88_n,
  G89_p,
  G89_n,
  G90_p,
  G90_n,
  G91_p,
  G91_n,
  G92_p,
  G92_n,
  G93_p,
  G93_n,
  G94_p,
  G94_n,
  G95_p,
  G95_n,
  G96_p,
  G96_n,
  G97_p,
  G97_n,
  G98_p,
  G98_n,
  G99_p,
  G99_n,
  G100_p,
  G100_n,
  G101_p,
  G101_n,
  G102_p,
  G102_n,
  G103_p,
  G103_n,
  G104_p,
  G104_n,
  G105_p,
  G105_n,
  G106_p,
  G106_n,
  G107_p,
  G107_n,
  G108_p,
  G108_n,
  G109_p,
  G109_n,
  G110_p,
  G110_n,
  G111_p,
  G111_n,
  G112_p,
  G112_n,
  G113_p,
  G113_n,
  G114_p,
  G114_n,
  G115_p,
  G115_n,
  G116_p,
  G116_n,
  G117_p,
  G117_n,
  G118_p,
  G118_n,
  G119_p,
  G119_n,
  G120_p,
  G120_n,
  G121_p,
  G121_n,
  G122_p,
  G122_n,
  G123_p,
  G123_n,
  G124_p,
  G124_n,
  G125_p,
  G125_n,
  G126_p,
  G126_n,
  G127_p,
  G127_n,
  G128_p,
  G128_n,
  G129_p,
  G129_n,
  G130_p,
  G130_n,
  G131_p,
  G131_n,
  G132_p,
  G132_n,
  G133_p,
  G133_n,
  G134_p,
  G134_n,
  G135_p,
  G135_n,
  G136_p,
  G136_n,
  G137_p,
  G137_n,
  G138_p,
  G138_n,
  G139_p,
  G139_n,
  G140_p,
  G140_n,
  G141_p,
  G141_n,
  G142_p,
  G142_n,
  G143_p,
  G143_n,
  G144_p,
  G144_n,
  G145_p,
  G145_n,
  G146_p,
  G146_n,
  G147_p,
  G147_n,
  G148_p,
  G148_n,
  G149_p,
  G149_n,
  G150_p,
  G150_n,
  G151_p,
  G151_n,
  G152_p,
  G152_n,
  G153_p,
  G153_n,
  G154_p,
  G154_n,
  G155_p,
  G155_n,
  G156_p,
  G156_n,
  G157_p,
  G157_n,
  G2531_p,
  G2532_p,
  G2533_p,
  G2534_p,
  G2535_p,
  G2536_p,
  G2537_p,
  G2538_p,
  G2539_p,
  G2540_p,
  G2541_p,
  G2542_p,
  G2543_p,
  G2544_p,
  G2545_p,
  G2546_p,
  G2547_p,
  G2548_p,
  G2549_p,
  G2550_p,
  G2551_p,
  G2552_p,
  G2553_p,
  G2554_p,
  G2555_p,
  G2556_p,
  G2557_p,
  G2558_p,
  G2559_p,
  G2560_p,
  G2561_p,
  G2562_p,
  G2563_p,
  G2564_p,
  G2565_p,
  G2566_p,
  G2567_p,
  G2568_p,
  G2569_p,
  G2570_p,
  G2571_p,
  G2572_p,
  G2573_p,
  G2574_p,
  G2575_p,
  G2576_p,
  G2577_p,
  G2578_p,
  G2579_p,
  G2580_p,
  G2581_n,
  G2582_p,
  G2583_p,
  G2584_p,
  G2585_p,
  G2586_p,
  G2587_n,
  G2588_p,
  G2589_p,
  G2590_n,
  G2591_p,
  G2592_p,
  G2593_p,
  G2594_p
);

  input G1_p;input G1_n;input G2_p;input G2_n;input G3_p;input G3_n;input G4_p;input G4_n;input G5_p;input G5_n;input G6_p;input G6_n;input G7_p;input G7_n;input G8_p;input G8_n;input G9_p;input G9_n;input G10_p;input G10_n;input G11_p;input G11_n;input G12_p;input G12_n;input G13_p;input G13_n;input G14_p;input G14_n;input G15_p;input G15_n;input G16_p;input G16_n;input G17_p;input G17_n;input G18_p;input G18_n;input G19_p;input G19_n;input G20_p;input G20_n;input G21_p;input G21_n;input G22_p;input G22_n;input G23_p;input G23_n;input G24_p;input G24_n;input G25_p;input G25_n;input G26_p;input G26_n;input G27_p;input G27_n;input G28_p;input G28_n;input G29_p;input G29_n;input G30_p;input G30_n;input G31_p;input G31_n;input G32_p;input G32_n;input G33_p;input G33_n;input G34_p;input G34_n;input G35_p;input G35_n;input G36_p;input G36_n;input G37_p;input G37_n;input G38_p;input G38_n;input G39_p;input G39_n;input G40_p;input G40_n;input G41_p;input G41_n;input G42_p;input G42_n;input G43_p;input G43_n;input G44_p;input G44_n;input G45_p;input G45_n;input G46_p;input G46_n;input G47_p;input G47_n;input G48_p;input G48_n;input G49_p;input G49_n;input G50_p;input G50_n;input G51_p;input G51_n;input G52_p;input G52_n;input G53_p;input G53_n;input G54_p;input G54_n;input G55_p;input G55_n;input G56_p;input G56_n;input G57_p;input G57_n;input G58_p;input G58_n;input G59_p;input G59_n;input G60_p;input G60_n;input G61_p;input G61_n;input G62_p;input G62_n;input G63_p;input G63_n;input G64_p;input G64_n;input G65_p;input G65_n;input G66_p;input G66_n;input G67_p;input G67_n;input G68_p;input G68_n;input G69_p;input G69_n;input G70_p;input G70_n;input G71_p;input G71_n;input G72_p;input G72_n;input G73_p;input G73_n;input G74_p;input G74_n;input G75_p;input G75_n;input G76_p;input G76_n;input G77_p;input G77_n;input G78_p;input G78_n;input G79_p;input G79_n;input G80_p;input G80_n;input G81_p;input G81_n;input G82_p;input G82_n;input G83_p;input G83_n;input G84_p;input G84_n;input G85_p;input G85_n;input G86_p;input G86_n;input G87_p;input G87_n;input G88_p;input G88_n;input G89_p;input G89_n;input G90_p;input G90_n;input G91_p;input G91_n;input G92_p;input G92_n;input G93_p;input G93_n;input G94_p;input G94_n;input G95_p;input G95_n;input G96_p;input G96_n;input G97_p;input G97_n;input G98_p;input G98_n;input G99_p;input G99_n;input G100_p;input G100_n;input G101_p;input G101_n;input G102_p;input G102_n;input G103_p;input G103_n;input G104_p;input G104_n;input G105_p;input G105_n;input G106_p;input G106_n;input G107_p;input G107_n;input G108_p;input G108_n;input G109_p;input G109_n;input G110_p;input G110_n;input G111_p;input G111_n;input G112_p;input G112_n;input G113_p;input G113_n;input G114_p;input G114_n;input G115_p;input G115_n;input G116_p;input G116_n;input G117_p;input G117_n;input G118_p;input G118_n;input G119_p;input G119_n;input G120_p;input G120_n;input G121_p;input G121_n;input G122_p;input G122_n;input G123_p;input G123_n;input G124_p;input G124_n;input G125_p;input G125_n;input G126_p;input G126_n;input G127_p;input G127_n;input G128_p;input G128_n;input G129_p;input G129_n;input G130_p;input G130_n;input G131_p;input G131_n;input G132_p;input G132_n;input G133_p;input G133_n;input G134_p;input G134_n;input G135_p;input G135_n;input G136_p;input G136_n;input G137_p;input G137_n;input G138_p;input G138_n;input G139_p;input G139_n;input G140_p;input G140_n;input G141_p;input G141_n;input G142_p;input G142_n;input G143_p;input G143_n;input G144_p;input G144_n;input G145_p;input G145_n;input G146_p;input G146_n;input G147_p;input G147_n;input G148_p;input G148_n;input G149_p;input G149_n;input G150_p;input G150_n;input G151_p;input G151_n;input G152_p;input G152_n;input G153_p;input G153_n;input G154_p;input G154_n;input G155_p;input G155_n;input G156_p;input G156_n;input G157_p;input G157_n;
  output G2531_p;output G2532_p;output G2533_p;output G2534_p;output G2535_p;output G2536_p;output G2537_p;output G2538_p;output G2539_p;output G2540_p;output G2541_p;output G2542_p;output G2543_p;output G2544_p;output G2545_p;output G2546_p;output G2547_p;output G2548_p;output G2549_p;output G2550_p;output G2551_p;output G2552_p;output G2553_p;output G2554_p;output G2555_p;output G2556_p;output G2557_p;output G2558_p;output G2559_p;output G2560_p;output G2561_p;output G2562_p;output G2563_p;output G2564_p;output G2565_p;output G2566_p;output G2567_p;output G2568_p;output G2569_p;output G2570_p;output G2571_p;output G2572_p;output G2573_p;output G2574_p;output G2575_p;output G2576_p;output G2577_p;output G2578_p;output G2579_p;output G2580_p;output G2581_n;output G2582_p;output G2583_p;output G2584_p;output G2585_p;output G2586_p;output G2587_n;output G2588_p;output G2589_p;output G2590_n;output G2591_p;output G2592_p;output G2593_p;output G2594_p;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire G51_p;
  wire G51_n;
  wire G52_p;
  wire G52_n;
  wire G53_p;
  wire G53_n;
  wire G54_p;
  wire G54_n;
  wire G55_p;
  wire G55_n;
  wire G56_p;
  wire G56_n;
  wire G57_p;
  wire G57_n;
  wire G58_p;
  wire G58_n;
  wire G59_p;
  wire G59_n;
  wire G60_p;
  wire G60_n;
  wire G61_p;
  wire G61_n;
  wire G62_p;
  wire G62_n;
  wire G63_p;
  wire G63_n;
  wire G64_p;
  wire G64_n;
  wire G65_p;
  wire G65_n;
  wire G66_p;
  wire G66_n;
  wire G67_p;
  wire G67_n;
  wire G68_p;
  wire G68_n;
  wire G69_p;
  wire G69_n;
  wire G70_p;
  wire G70_n;
  wire G71_p;
  wire G71_n;
  wire G72_p;
  wire G72_n;
  wire G73_p;
  wire G73_n;
  wire G74_p;
  wire G74_n;
  wire G75_p;
  wire G75_n;
  wire G76_p;
  wire G76_n;
  wire G77_p;
  wire G77_n;
  wire G78_p;
  wire G78_n;
  wire G79_p;
  wire G79_n;
  wire G80_p;
  wire G80_n;
  wire G81_p;
  wire G81_n;
  wire G82_p;
  wire G82_n;
  wire G83_p;
  wire G83_n;
  wire G84_p;
  wire G84_n;
  wire G85_p;
  wire G85_n;
  wire G86_p;
  wire G86_n;
  wire G87_p;
  wire G87_n;
  wire G88_p;
  wire G88_n;
  wire G89_p;
  wire G89_n;
  wire G90_p;
  wire G90_n;
  wire G91_p;
  wire G91_n;
  wire G92_p;
  wire G92_n;
  wire G93_p;
  wire G93_n;
  wire G94_p;
  wire G94_n;
  wire G95_p;
  wire G95_n;
  wire G96_p;
  wire G96_n;
  wire G97_p;
  wire G97_n;
  wire G98_p;
  wire G98_n;
  wire G99_p;
  wire G99_n;
  wire G100_p;
  wire G100_n;
  wire G101_p;
  wire G101_n;
  wire G102_p;
  wire G102_n;
  wire G103_p;
  wire G103_n;
  wire G104_p;
  wire G104_n;
  wire G105_p;
  wire G105_n;
  wire G106_p;
  wire G106_n;
  wire G107_p;
  wire G107_n;
  wire G108_p;
  wire G108_n;
  wire G109_p;
  wire G109_n;
  wire G110_p;
  wire G110_n;
  wire G111_p;
  wire G111_n;
  wire G112_p;
  wire G112_n;
  wire G113_p;
  wire G113_n;
  wire G114_p;
  wire G114_n;
  wire G115_p;
  wire G115_n;
  wire G116_p;
  wire G116_n;
  wire G117_p;
  wire G117_n;
  wire G118_p;
  wire G118_n;
  wire G119_p;
  wire G119_n;
  wire G120_p;
  wire G120_n;
  wire G121_p;
  wire G121_n;
  wire G122_p;
  wire G122_n;
  wire G123_p;
  wire G123_n;
  wire G124_p;
  wire G124_n;
  wire G125_p;
  wire G125_n;
  wire G126_p;
  wire G126_n;
  wire G127_p;
  wire G127_n;
  wire G128_p;
  wire G128_n;
  wire G129_p;
  wire G129_n;
  wire G130_p;
  wire G130_n;
  wire G131_p;
  wire G131_n;
  wire G132_p;
  wire G132_n;
  wire G133_p;
  wire G133_n;
  wire G134_p;
  wire G134_n;
  wire G135_p;
  wire G135_n;
  wire G136_p;
  wire G136_n;
  wire G137_p;
  wire G137_n;
  wire G138_p;
  wire G138_n;
  wire G139_p;
  wire G139_n;
  wire G140_p;
  wire G140_n;
  wire G141_p;
  wire G141_n;
  wire G142_p;
  wire G142_n;
  wire G143_p;
  wire G143_n;
  wire G144_p;
  wire G144_n;
  wire G145_p;
  wire G145_n;
  wire G146_p;
  wire G146_n;
  wire G147_p;
  wire G147_n;
  wire G148_p;
  wire G148_n;
  wire G149_p;
  wire G149_n;
  wire G150_p;
  wire G150_n;
  wire G151_p;
  wire G151_n;
  wire G152_p;
  wire G152_n;
  wire G153_p;
  wire G153_n;
  wire G154_p;
  wire G154_n;
  wire G155_p;
  wire G155_n;
  wire G156_p;
  wire G156_n;
  wire G157_p;
  wire G157_n;
  wire g158_p;
  wire g158_n;
  wire g159_p;
  wire g159_n;
  wire g160_p;
  wire g160_n;
  wire g161_p;
  wire g161_n;
  wire g162_p;
  wire g162_n;
  wire g163_p;
  wire g163_n;
  wire g164_p;
  wire g164_n;
  wire g165_p;
  wire g165_n;
  wire g166_p;
  wire g166_n;
  wire g167_p;
  wire g167_n;
  wire g168_p;
  wire g168_n;
  wire g169_p;
  wire g169_n;
  wire g170_p;
  wire g170_n;
  wire g171_p;
  wire g171_n;
  wire g172_p;
  wire g172_n;
  wire g173_p;
  wire g173_n;
  wire g174_p;
  wire g174_n;
  wire g175_p;
  wire g175_n;
  wire g176_p;
  wire g176_n;
  wire g177_p;
  wire g177_n;
  wire g178_p;
  wire g178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire g693_p;
  wire g693_n;
  wire g694_p;
  wire g694_n;
  wire g695_p;
  wire g695_n;
  wire g696_p;
  wire g696_n;
  wire g697_p;
  wire g697_n;
  wire g698_p;
  wire g698_n;
  wire g699_p;
  wire g699_n;
  wire g700_p;
  wire g700_n;
  wire g701_p;
  wire g701_n;
  wire g702_p;
  wire g702_n;
  wire g703_p;
  wire g703_n;
  wire g704_p;
  wire g704_n;
  wire g705_p;
  wire g705_n;
  wire g706_p;
  wire g706_n;
  wire g707_p;
  wire g707_n;
  wire g708_p;
  wire g708_n;
  wire g709_p;
  wire g709_n;
  wire g710_p;
  wire g710_n;
  wire g711_p;
  wire g711_n;
  wire g712_p;
  wire g712_n;
  wire g713_p;
  wire g713_n;
  wire g714_p;
  wire g714_n;
  wire g715_p;
  wire g715_n;
  wire g716_p;
  wire g716_n;
  wire g717_p;
  wire g717_n;
  wire g718_p;
  wire g718_n;
  wire G141_p_spl_;
  wire G141_p_spl_0;
  wire G141_p_spl_1;
  wire G142_p_spl_;
  wire G142_p_spl_0;
  wire G142_p_spl_1;
  wire G141_n_spl_;
  wire G141_n_spl_0;
  wire G142_n_spl_;
  wire G142_n_spl_0;
  wire G139_p_spl_;
  wire G139_p_spl_0;
  wire G139_p_spl_1;
  wire G140_p_spl_;
  wire G140_p_spl_0;
  wire G140_p_spl_1;
  wire G139_n_spl_;
  wire G139_n_spl_0;
  wire G140_n_spl_;
  wire G140_n_spl_0;
  wire g158_n_spl_;
  wire g159_n_spl_;
  wire G121_n_spl_;
  wire G115_n_spl_;
  wire G115_n_spl_0;
  wire G115_n_spl_1;
  wire g164_n_spl_;
  wire g164_n_spl_0;
  wire G43_n_spl_;
  wire G53_n_spl_;
  wire G86_n_spl_;
  wire G96_n_spl_;
  wire G32_n_spl_;
  wire G64_n_spl_;
  wire G76_n_spl_;
  wire G106_n_spl_;
  wire g169_n_spl_;
  wire g172_n_spl_;
  wire G145_n_spl_;
  wire G145_n_spl_0;
  wire G145_n_spl_00;
  wire G145_n_spl_000;
  wire G145_n_spl_0000;
  wire G145_n_spl_00000;
  wire G145_n_spl_00001;
  wire G145_n_spl_0001;
  wire G145_n_spl_00010;
  wire G145_n_spl_00011;
  wire G145_n_spl_001;
  wire G145_n_spl_0010;
  wire G145_n_spl_0011;
  wire G145_n_spl_01;
  wire G145_n_spl_010;
  wire G145_n_spl_0100;
  wire G145_n_spl_0101;
  wire G145_n_spl_011;
  wire G145_n_spl_0110;
  wire G145_n_spl_0111;
  wire G145_n_spl_1;
  wire G145_n_spl_10;
  wire G145_n_spl_100;
  wire G145_n_spl_1000;
  wire G145_n_spl_1001;
  wire G145_n_spl_101;
  wire G145_n_spl_1010;
  wire G145_n_spl_1011;
  wire G145_n_spl_11;
  wire G145_n_spl_110;
  wire G145_n_spl_1100;
  wire G145_n_spl_1101;
  wire G145_n_spl_111;
  wire G145_n_spl_1110;
  wire G145_n_spl_1111;
  wire G145_p_spl_;
  wire G145_p_spl_0;
  wire G145_p_spl_00;
  wire G145_p_spl_000;
  wire G145_p_spl_0000;
  wire G145_p_spl_00000;
  wire G145_p_spl_00001;
  wire G145_p_spl_0001;
  wire G145_p_spl_00010;
  wire G145_p_spl_00011;
  wire G145_p_spl_001;
  wire G145_p_spl_0010;
  wire G145_p_spl_0011;
  wire G145_p_spl_01;
  wire G145_p_spl_010;
  wire G145_p_spl_0100;
  wire G145_p_spl_0101;
  wire G145_p_spl_011;
  wire G145_p_spl_0110;
  wire G145_p_spl_0111;
  wire G145_p_spl_1;
  wire G145_p_spl_10;
  wire G145_p_spl_100;
  wire G145_p_spl_1000;
  wire G145_p_spl_1001;
  wire G145_p_spl_101;
  wire G145_p_spl_1010;
  wire G145_p_spl_1011;
  wire G145_p_spl_11;
  wire G145_p_spl_110;
  wire G145_p_spl_1100;
  wire G145_p_spl_1101;
  wire G145_p_spl_111;
  wire G145_p_spl_1110;
  wire G145_p_spl_1111;
  wire G146_p_spl_;
  wire G146_p_spl_0;
  wire G146_p_spl_00;
  wire G146_p_spl_000;
  wire G146_p_spl_0000;
  wire G146_p_spl_0001;
  wire G146_p_spl_001;
  wire G146_p_spl_01;
  wire G146_p_spl_010;
  wire G146_p_spl_011;
  wire G146_p_spl_1;
  wire G146_p_spl_10;
  wire G146_p_spl_100;
  wire G146_p_spl_101;
  wire G146_p_spl_11;
  wire G146_p_spl_110;
  wire G146_p_spl_111;
  wire G146_n_spl_;
  wire G146_n_spl_0;
  wire G146_n_spl_00;
  wire G146_n_spl_000;
  wire G146_n_spl_0000;
  wire G146_n_spl_0001;
  wire G146_n_spl_001;
  wire G146_n_spl_01;
  wire G146_n_spl_010;
  wire G146_n_spl_011;
  wire G146_n_spl_1;
  wire G146_n_spl_10;
  wire G146_n_spl_100;
  wire G146_n_spl_101;
  wire G146_n_spl_11;
  wire G146_n_spl_110;
  wire G146_n_spl_111;
  wire G117_p_spl_;
  wire G117_p_spl_0;
  wire G117_p_spl_00;
  wire G117_p_spl_000;
  wire G117_p_spl_0000;
  wire G117_p_spl_0001;
  wire G117_p_spl_001;
  wire G117_p_spl_0010;
  wire G117_p_spl_0011;
  wire G117_p_spl_01;
  wire G117_p_spl_010;
  wire G117_p_spl_0100;
  wire G117_p_spl_0101;
  wire G117_p_spl_011;
  wire G117_p_spl_0110;
  wire G117_p_spl_0111;
  wire G117_p_spl_1;
  wire G117_p_spl_10;
  wire G117_p_spl_100;
  wire G117_p_spl_1000;
  wire G117_p_spl_1001;
  wire G117_p_spl_101;
  wire G117_p_spl_1010;
  wire G117_p_spl_1011;
  wire G117_p_spl_11;
  wire G117_p_spl_110;
  wire G117_p_spl_1100;
  wire G117_p_spl_1101;
  wire G117_p_spl_111;
  wire G117_p_spl_1110;
  wire G120_n_spl_;
  wire G120_n_spl_0;
  wire G120_n_spl_00;
  wire G120_n_spl_000;
  wire G120_n_spl_0000;
  wire G120_n_spl_0001;
  wire G120_n_spl_001;
  wire G120_n_spl_0010;
  wire G120_n_spl_0011;
  wire G120_n_spl_01;
  wire G120_n_spl_010;
  wire G120_n_spl_0100;
  wire G120_n_spl_011;
  wire G120_n_spl_1;
  wire G120_n_spl_10;
  wire G120_n_spl_100;
  wire G120_n_spl_101;
  wire G120_n_spl_11;
  wire G120_n_spl_110;
  wire G120_n_spl_111;
  wire G117_n_spl_;
  wire G117_n_spl_0;
  wire G117_n_spl_00;
  wire G117_n_spl_000;
  wire G117_n_spl_0000;
  wire G117_n_spl_0001;
  wire G117_n_spl_001;
  wire G117_n_spl_0010;
  wire G117_n_spl_0011;
  wire G117_n_spl_01;
  wire G117_n_spl_010;
  wire G117_n_spl_0100;
  wire G117_n_spl_0101;
  wire G117_n_spl_011;
  wire G117_n_spl_0110;
  wire G117_n_spl_0111;
  wire G117_n_spl_1;
  wire G117_n_spl_10;
  wire G117_n_spl_100;
  wire G117_n_spl_1000;
  wire G117_n_spl_1001;
  wire G117_n_spl_101;
  wire G117_n_spl_1010;
  wire G117_n_spl_1011;
  wire G117_n_spl_11;
  wire G117_n_spl_110;
  wire G117_n_spl_1100;
  wire G117_n_spl_1101;
  wire G117_n_spl_111;
  wire G117_n_spl_1110;
  wire G120_p_spl_;
  wire G120_p_spl_0;
  wire G120_p_spl_00;
  wire G120_p_spl_000;
  wire G120_p_spl_0000;
  wire G120_p_spl_0001;
  wire G120_p_spl_001;
  wire G120_p_spl_0010;
  wire G120_p_spl_0011;
  wire G120_p_spl_01;
  wire G120_p_spl_010;
  wire G120_p_spl_0100;
  wire G120_p_spl_011;
  wire G120_p_spl_1;
  wire G120_p_spl_10;
  wire G120_p_spl_100;
  wire G120_p_spl_101;
  wire G120_p_spl_11;
  wire G120_p_spl_110;
  wire G120_p_spl_111;
  wire g204_p_spl_;
  wire g204_p_spl_0;
  wire g204_p_spl_00;
  wire g204_p_spl_000;
  wire g204_p_spl_01;
  wire g204_p_spl_1;
  wire g204_p_spl_10;
  wire g204_p_spl_11;
  wire g204_n_spl_;
  wire g204_n_spl_0;
  wire g204_n_spl_00;
  wire g204_n_spl_000;
  wire g204_n_spl_01;
  wire g204_n_spl_1;
  wire g204_n_spl_10;
  wire g204_n_spl_11;
  wire G122_n_spl_;
  wire G122_n_spl_0;
  wire g240_n_spl_;
  wire g240_n_spl_0;
  wire g240_n_spl_00;
  wire g240_n_spl_1;
  wire g176_n_spl_;
  wire g176_n_spl_0;
  wire g243_n_spl_;
  wire G123_p_spl_;
  wire G123_p_spl_0;
  wire G123_p_spl_1;
  wire g231_n_spl_;
  wire g231_n_spl_0;
  wire g231_n_spl_00;
  wire g231_n_spl_1;
  wire G123_n_spl_;
  wire G123_n_spl_0;
  wire G123_n_spl_1;
  wire g290_p_spl_;
  wire g290_p_spl_0;
  wire g290_p_spl_00;
  wire g290_p_spl_01;
  wire g290_p_spl_1;
  wire g222_p_spl_;
  wire g222_p_spl_0;
  wire g222_p_spl_00;
  wire g222_p_spl_01;
  wire g222_p_spl_1;
  wire g255_n_spl_;
  wire g255_n_spl_0;
  wire g255_n_spl_00;
  wire g255_n_spl_1;
  wire G118_p_spl_;
  wire G118_p_spl_0;
  wire g290_n_spl_;
  wire g290_n_spl_0;
  wire g290_n_spl_00;
  wire g290_n_spl_01;
  wire g290_n_spl_1;
  wire g290_n_spl_10;
  wire g290_n_spl_11;
  wire G118_n_spl_;
  wire g298_p_spl_;
  wire g298_p_spl_0;
  wire g240_p_spl_;
  wire g240_p_spl_0;
  wire g240_p_spl_1;
  wire G143_n_spl_;
  wire G143_n_spl_0;
  wire g310_p_spl_;
  wire g310_p_spl_0;
  wire G143_p_spl_;
  wire G143_p_spl_0;
  wire g310_n_spl_;
  wire g310_n_spl_0;
  wire g310_n_spl_1;
  wire G144_p_spl_;
  wire G144_p_spl_0;
  wire G154_n_spl_;
  wire G155_n_spl_;
  wire G154_p_spl_;
  wire G155_p_spl_;
  wire G125_n_spl_;
  wire G125_n_spl_0;
  wire G126_n_spl_;
  wire G126_n_spl_0;
  wire G125_p_spl_;
  wire G125_p_spl_0;
  wire G125_p_spl_1;
  wire G126_p_spl_;
  wire G126_p_spl_0;
  wire G126_p_spl_1;
  wire g317_p_spl_;
  wire g320_n_spl_;
  wire g317_n_spl_;
  wire g320_p_spl_;
  wire G152_n_spl_;
  wire G153_n_spl_;
  wire G152_p_spl_;
  wire G153_p_spl_;
  wire G148_n_spl_;
  wire G149_n_spl_;
  wire G148_p_spl_;
  wire G149_p_spl_;
  wire g326_n_spl_;
  wire g329_n_spl_;
  wire g326_p_spl_;
  wire g329_p_spl_;
  wire G150_n_spl_;
  wire G151_n_spl_;
  wire G150_p_spl_;
  wire G151_p_spl_;
  wire g332_n_spl_;
  wire g335_n_spl_;
  wire g332_p_spl_;
  wire g335_p_spl_;
  wire G138_p_spl_;
  wire G138_p_spl_0;
  wire G138_p_spl_00;
  wire G138_p_spl_1;
  wire G157_n_spl_;
  wire G138_n_spl_;
  wire G138_n_spl_0;
  wire G138_n_spl_1;
  wire G157_p_spl_;
  wire g346_n_spl_;
  wire g349_n_spl_;
  wire g346_p_spl_;
  wire g349_p_spl_;
  wire g344_n_spl_;
  wire g352_n_spl_;
  wire g344_p_spl_;
  wire g352_p_spl_;
  wire G144_n_spl_;
  wire G133_n_spl_;
  wire G133_n_spl_0;
  wire G134_n_spl_;
  wire G134_n_spl_0;
  wire G134_n_spl_1;
  wire G133_p_spl_;
  wire G133_p_spl_0;
  wire G133_p_spl_1;
  wire G134_p_spl_;
  wire G134_p_spl_0;
  wire G134_p_spl_1;
  wire G135_n_spl_;
  wire G135_n_spl_0;
  wire G135_n_spl_1;
  wire G136_n_spl_;
  wire G136_n_spl_0;
  wire G136_n_spl_1;
  wire G135_p_spl_;
  wire G135_p_spl_0;
  wire G135_p_spl_1;
  wire G136_p_spl_;
  wire G136_p_spl_0;
  wire G136_p_spl_00;
  wire G136_p_spl_1;
  wire g364_p_spl_;
  wire g367_n_spl_;
  wire g364_n_spl_;
  wire g367_p_spl_;
  wire G131_n_spl_;
  wire G131_n_spl_0;
  wire G132_n_spl_;
  wire G132_n_spl_0;
  wire G131_p_spl_;
  wire G131_p_spl_0;
  wire G131_p_spl_1;
  wire G132_p_spl_;
  wire G132_p_spl_0;
  wire G132_p_spl_1;
  wire G128_p_spl_;
  wire G128_p_spl_0;
  wire G128_p_spl_1;
  wire G156_n_spl_;
  wire G128_n_spl_;
  wire G128_n_spl_0;
  wire G156_p_spl_;
  wire g373_n_spl_;
  wire g376_n_spl_;
  wire g373_p_spl_;
  wire g376_p_spl_;
  wire G129_n_spl_;
  wire G129_n_spl_0;
  wire G130_n_spl_;
  wire G130_n_spl_0;
  wire G129_p_spl_;
  wire G129_p_spl_0;
  wire G129_p_spl_1;
  wire G130_p_spl_;
  wire G130_p_spl_0;
  wire G130_p_spl_1;
  wire g379_n_spl_;
  wire g382_n_spl_;
  wire g379_p_spl_;
  wire g382_p_spl_;
  wire G12_n_spl_;
  wire G12_n_spl_0;
  wire G12_n_spl_00;
  wire G12_n_spl_000;
  wire G12_n_spl_0000;
  wire G12_n_spl_0001;
  wire G12_n_spl_001;
  wire G12_n_spl_01;
  wire G12_n_spl_010;
  wire G12_n_spl_011;
  wire G12_n_spl_1;
  wire G12_n_spl_10;
  wire G12_n_spl_100;
  wire G12_n_spl_101;
  wire G12_n_spl_11;
  wire G12_n_spl_110;
  wire G12_n_spl_111;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire G12_p_spl_00;
  wire G12_p_spl_000;
  wire G12_p_spl_0000;
  wire G12_p_spl_0001;
  wire G12_p_spl_001;
  wire G12_p_spl_01;
  wire G12_p_spl_010;
  wire G12_p_spl_011;
  wire G12_p_spl_1;
  wire G12_p_spl_10;
  wire G12_p_spl_100;
  wire G12_p_spl_101;
  wire G12_p_spl_11;
  wire G12_p_spl_110;
  wire G12_p_spl_111;
  wire g222_n_spl_;
  wire g222_n_spl_0;
  wire g222_n_spl_1;
  wire g231_p_spl_;
  wire g231_p_spl_0;
  wire g231_p_spl_00;
  wire g231_p_spl_01;
  wire g231_p_spl_1;
  wire g213_p_spl_;
  wire g213_p_spl_0;
  wire g213_p_spl_00;
  wire g213_p_spl_1;
  wire g213_n_spl_;
  wire g213_n_spl_0;
  wire g213_n_spl_1;
  wire G23_n_spl_;
  wire G23_n_spl_0;
  wire G23_n_spl_00;
  wire G23_n_spl_000;
  wire G23_n_spl_001;
  wire G23_n_spl_01;
  wire G23_n_spl_010;
  wire G23_n_spl_011;
  wire G23_n_spl_1;
  wire G23_n_spl_10;
  wire G23_n_spl_100;
  wire G23_n_spl_101;
  wire G23_n_spl_11;
  wire G23_n_spl_110;
  wire G23_p_spl_;
  wire G23_p_spl_0;
  wire G23_p_spl_00;
  wire G23_p_spl_000;
  wire G23_p_spl_001;
  wire G23_p_spl_01;
  wire G23_p_spl_010;
  wire G23_p_spl_011;
  wire G23_p_spl_1;
  wire G23_p_spl_10;
  wire G23_p_spl_100;
  wire G23_p_spl_101;
  wire G23_p_spl_11;
  wire G23_p_spl_110;
  wire g185_n_spl_;
  wire g185_n_spl_0;
  wire g185_n_spl_00;
  wire g185_n_spl_1;
  wire g185_p_spl_;
  wire g185_p_spl_0;
  wire g185_p_spl_1;
  wire g203_n_spl_;
  wire g203_n_spl_0;
  wire g203_n_spl_00;
  wire g203_n_spl_1;
  wire g203_p_spl_;
  wire g203_p_spl_0;
  wire g203_p_spl_1;
  wire g427_n_spl_;
  wire g427_n_spl_0;
  wire g427_n_spl_1;
  wire g427_p_spl_;
  wire g427_p_spl_0;
  wire g427_p_spl_1;
  wire g255_p_spl_;
  wire g255_p_spl_0;
  wire g255_p_spl_00;
  wire g255_p_spl_1;
  wire g262_n_spl_;
  wire g262_n_spl_0;
  wire g262_n_spl_1;
  wire g262_p_spl_;
  wire g262_p_spl_0;
  wire g262_p_spl_1;
  wire g271_p_spl_;
  wire g271_p_spl_0;
  wire g271_p_spl_1;
  wire g271_n_spl_;
  wire g271_n_spl_0;
  wire g271_n_spl_1;
  wire g280_p_spl_;
  wire g280_p_spl_0;
  wire g280_p_spl_1;
  wire g280_n_spl_;
  wire g280_n_spl_0;
  wire g280_n_spl_00;
  wire g280_n_spl_1;
  wire g484_n_spl_;
  wire g484_n_spl_0;
  wire g484_n_spl_1;
  wire g484_p_spl_;
  wire g484_p_spl_0;
  wire g484_p_spl_1;
  wire g503_n_spl_;
  wire g503_n_spl_0;
  wire g503_p_spl_;
  wire g503_p_spl_0;
  wire g194_n_spl_;
  wire g194_n_spl_0;
  wire g194_n_spl_1;
  wire g194_p_spl_;
  wire g194_p_spl_0;
  wire g522_n_spl_;
  wire g522_n_spl_0;
  wire g522_n_spl_1;
  wire g522_p_spl_;
  wire g522_p_spl_0;
  wire g522_p_spl_1;
  wire g550_n_spl_;
  wire g550_n_spl_0;
  wire g550_n_spl_1;
  wire g550_p_spl_;
  wire g553_n_spl_;
  wire g553_n_spl_0;
  wire g553_p_spl_;
  wire g553_p_spl_0;
  wire g562_p_spl_;
  wire g562_n_spl_;
  wire g574_p_spl_;
  wire g574_n_spl_;
  wire g577_p_spl_;
  wire g580_n_spl_;
  wire g577_n_spl_;
  wire g580_p_spl_;
  wire g583_n_spl_;
  wire g586_n_spl_;
  wire g583_p_spl_;
  wire g586_p_spl_;
  wire G29_n_spl_;
  wire g597_p_spl_;
  wire g600_n_spl_;
  wire g597_n_spl_;
  wire g600_p_spl_;
  wire g606_n_spl_;
  wire g606_p_spl_;
  wire g609_n_spl_;
  wire g609_n_spl_0;
  wire g609_n_spl_1;
  wire g298_n_spl_;
  wire g609_p_spl_;
  wire g609_p_spl_0;
  wire g609_p_spl_1;
  wire g603_p_spl_;
  wire g603_n_spl_;
  wire g620_p_spl_;
  wire g620_n_spl_;
  wire g628_p_spl_;
  wire g629_p_spl_;
  wire g628_n_spl_;
  wire g629_n_spl_;
  wire G8_n_spl_;
  wire g630_p_spl_;
  wire g630_p_spl_0;
  wire g630_p_spl_00;
  wire g630_p_spl_01;
  wire g630_p_spl_1;
  wire g631_n_spl_;
  wire g631_n_spl_0;
  wire g631_n_spl_1;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire g630_n_spl_;
  wire g630_n_spl_0;
  wire g630_n_spl_00;
  wire g630_n_spl_1;
  wire g633_p_spl_;
  wire g633_n_spl_;
  wire g637_p_spl_;
  wire g640_p_spl_;
  wire g643_p_spl_;
  wire g646_p_spl_;
  wire g651_n_spl_;
  wire g656_n_spl_;
  wire g661_n_spl_;
  wire g682_p_spl_;
  wire g682_p_spl_0;
  wire g682_p_spl_00;
  wire g682_p_spl_01;
  wire g682_p_spl_1;
  wire g682_p_spl_10;
  wire g682_p_spl_11;
  wire g682_n_spl_;
  wire g682_n_spl_0;
  wire g682_n_spl_00;
  wire g682_n_spl_01;
  wire g682_n_spl_1;
  wire g682_n_spl_10;
  wire g682_n_spl_11;
  wire g683_n_spl_;
  wire g684_p_spl_;
  wire g686_n_spl_;
  wire g687_p_spl_;
  wire g690_n_spl_;
  wire g694_n_spl_;
  wire g695_p_spl_;
  wire g699_p_spl_;
  wire g700_n_spl_;
  wire g698_n_spl_;
  wire g693_n_spl_;
  wire g342_p_spl_;
  wire g361_p_spl_;
  wire g388_p_spl_;
  wire g593_p_spl_;
  wire g627_p_spl_;
  wire G124_n_spl_;
  wire G137_n_spl_;
  wire G137_n_spl_0;
  wire g173_n_spl_;
  wire g292_n_spl_;
  wire g295_n_spl_;
  wire g301_n_spl_;
  wire g540_n_spl_;
  wire g617_p_spl_;
  wire g718_n_spl_;

  LA
  g_g158_p
  (
    .dout(g158_p),
    .din1(G141_p_spl_0),
    .din2(G142_p_spl_0)
  );


  FA
  g_g158_n
  (
    .dout(g158_n),
    .din1(G141_n_spl_0),
    .din2(G142_n_spl_0)
  );


  LA
  g_g159_p
  (
    .dout(g159_p),
    .din1(G139_p_spl_0),
    .din2(G140_p_spl_0)
  );


  FA
  g_g159_n
  (
    .dout(g159_n),
    .din1(G139_n_spl_0),
    .din2(G140_n_spl_0)
  );


  FA
  g_g160_n
  (
    .dout(g160_n),
    .din1(g158_n_spl_),
    .din2(g159_n_spl_)
  );


  FA
  g_g161_n
  (
    .dout(g161_n),
    .din1(G2_n),
    .din2(G121_n_spl_)
  );


  FA
  g_g162_n
  (
    .dout(g162_n),
    .din1(G11_n),
    .din2(g161_n)
  );


  LA
  g_g163_p
  (
    .dout(g163_p),
    .din1(G74_p),
    .din2(G115_n_spl_0)
  );


  FA
  g_g164_n
  (
    .dout(g164_n),
    .din1(G7_n),
    .din2(G121_n_spl_)
  );


  FA
  g_g165_n
  (
    .dout(g165_n),
    .din1(G119_n),
    .din2(g164_n_spl_0)
  );


  FA
  g_g166_n
  (
    .dout(g166_n),
    .din1(G147_n),
    .din2(g164_n_spl_0)
  );


  FA
  g_g167_n
  (
    .dout(g167_n),
    .din1(G43_n_spl_),
    .din2(G53_n_spl_)
  );


  FA
  g_g168_n
  (
    .dout(g168_n),
    .din1(G86_n_spl_),
    .din2(G96_n_spl_)
  );


  FA
  g_g169_n
  (
    .dout(g169_n),
    .din1(g167_n),
    .din2(g168_n)
  );


  FA
  g_g170_n
  (
    .dout(g170_n),
    .din1(G32_n_spl_),
    .din2(G64_n_spl_)
  );


  FA
  g_g171_n
  (
    .dout(g171_n),
    .din1(G76_n_spl_),
    .din2(G106_n_spl_)
  );


  FA
  g_g172_n
  (
    .dout(g172_n),
    .din1(g170_n),
    .din2(g171_n)
  );


  FA
  g_g173_n
  (
    .dout(g173_n),
    .din1(g169_n_spl_),
    .din2(g172_n_spl_)
  );


  LA
  g_g174_p
  (
    .dout(g174_p),
    .din1(G147_p),
    .din2(g172_n_spl_)
  );


  LA
  g_g175_p
  (
    .dout(g175_p),
    .din1(G119_p),
    .din2(g169_n_spl_)
  );


  FA
  g_g176_n
  (
    .dout(g176_n),
    .din1(g174_p),
    .din2(g175_p)
  );


  LA
  g_g177_p
  (
    .dout(g177_p),
    .din1(G79_n),
    .din2(G145_n_spl_00000)
  );


  FA
  g_g177_n
  (
    .dout(g177_n),
    .din1(G79_p),
    .din2(G145_p_spl_00000)
  );


  LA
  g_g178_p
  (
    .dout(g178_p),
    .din1(G109_n),
    .din2(G145_p_spl_00000)
  );


  FA
  g_g178_n
  (
    .dout(g178_n),
    .din1(G109_p),
    .din2(G145_n_spl_00000)
  );


  LA
  g_g179_p
  (
    .dout(g179_p),
    .din1(g177_n),
    .din2(g178_n)
  );


  FA
  g_g179_n
  (
    .dout(g179_n),
    .din1(g177_p),
    .din2(g178_p)
  );


  LA
  g_g180_p
  (
    .dout(g180_p),
    .din1(G146_p_spl_0000),
    .din2(g179_n)
  );


  FA
  g_g180_n
  (
    .dout(g180_n),
    .din1(G146_n_spl_0000),
    .din2(g179_p)
  );


  LA
  g_g181_p
  (
    .dout(g181_p),
    .din1(G99_n),
    .din2(G145_p_spl_00001)
  );


  FA
  g_g181_n
  (
    .dout(g181_n),
    .din1(G99_p),
    .din2(G145_n_spl_00001)
  );


  LA
  g_g182_p
  (
    .dout(g182_p),
    .din1(G89_n),
    .din2(G145_n_spl_00001)
  );


  FA
  g_g182_n
  (
    .dout(g182_n),
    .din1(G89_p),
    .din2(G145_p_spl_00001)
  );


  LA
  g_g183_p
  (
    .dout(g183_p),
    .din1(g181_n),
    .din2(g182_n)
  );


  FA
  g_g183_n
  (
    .dout(g183_n),
    .din1(g181_p),
    .din2(g182_p)
  );


  LA
  g_g184_p
  (
    .dout(g184_p),
    .din1(G146_n_spl_0000),
    .din2(g183_n)
  );


  FA
  g_g184_n
  (
    .dout(g184_n),
    .din1(G146_p_spl_0000),
    .din2(g183_p)
  );


  LA
  g_g185_p
  (
    .dout(g185_p),
    .din1(g180_n),
    .din2(g184_n)
  );


  FA
  g_g185_n
  (
    .dout(g185_n),
    .din1(g180_p),
    .din2(g184_p)
  );


  LA
  g_g186_p
  (
    .dout(g186_p),
    .din1(G78_n),
    .din2(G145_n_spl_00010)
  );


  FA
  g_g186_n
  (
    .dout(g186_n),
    .din1(G78_p),
    .din2(G145_p_spl_00010)
  );


  LA
  g_g187_p
  (
    .dout(g187_p),
    .din1(G108_n),
    .din2(G145_p_spl_00010)
  );


  FA
  g_g187_n
  (
    .dout(g187_n),
    .din1(G108_p),
    .din2(G145_n_spl_00010)
  );


  LA
  g_g188_p
  (
    .dout(g188_p),
    .din1(g186_n),
    .din2(g187_n)
  );


  FA
  g_g188_n
  (
    .dout(g188_n),
    .din1(g186_p),
    .din2(g187_p)
  );


  LA
  g_g189_p
  (
    .dout(g189_p),
    .din1(G146_p_spl_0001),
    .din2(g188_n)
  );


  FA
  g_g189_n
  (
    .dout(g189_n),
    .din1(G146_n_spl_0001),
    .din2(g188_p)
  );


  LA
  g_g190_p
  (
    .dout(g190_p),
    .din1(G98_n),
    .din2(G145_p_spl_00011)
  );


  FA
  g_g190_n
  (
    .dout(g190_n),
    .din1(G98_p),
    .din2(G145_n_spl_00011)
  );


  LA
  g_g191_p
  (
    .dout(g191_p),
    .din1(G88_n),
    .din2(G145_n_spl_00011)
  );


  FA
  g_g191_n
  (
    .dout(g191_n),
    .din1(G88_p),
    .din2(G145_p_spl_00011)
  );


  LA
  g_g192_p
  (
    .dout(g192_p),
    .din1(g190_n),
    .din2(g191_n)
  );


  FA
  g_g192_n
  (
    .dout(g192_n),
    .din1(g190_p),
    .din2(g191_p)
  );


  LA
  g_g193_p
  (
    .dout(g193_p),
    .din1(G146_n_spl_0001),
    .din2(g192_n)
  );


  FA
  g_g193_n
  (
    .dout(g193_n),
    .din1(G146_p_spl_0001),
    .din2(g192_p)
  );


  LA
  g_g194_p
  (
    .dout(g194_p),
    .din1(g189_n),
    .din2(g193_n)
  );


  FA
  g_g194_n
  (
    .dout(g194_n),
    .din1(g189_p),
    .din2(g193_p)
  );


  LA
  g_g195_p
  (
    .dout(g195_p),
    .din1(G80_n),
    .din2(G145_n_spl_0010)
  );


  FA
  g_g195_n
  (
    .dout(g195_n),
    .din1(G80_p),
    .din2(G145_p_spl_0010)
  );


  LA
  g_g196_p
  (
    .dout(g196_p),
    .din1(G110_n),
    .din2(G145_p_spl_0010)
  );


  FA
  g_g196_n
  (
    .dout(g196_n),
    .din1(G110_p),
    .din2(G145_n_spl_0010)
  );


  LA
  g_g197_p
  (
    .dout(g197_p),
    .din1(g195_n),
    .din2(g196_n)
  );


  FA
  g_g197_n
  (
    .dout(g197_n),
    .din1(g195_p),
    .din2(g196_p)
  );


  LA
  g_g198_p
  (
    .dout(g198_p),
    .din1(G146_p_spl_001),
    .din2(g197_n)
  );


  FA
  g_g198_n
  (
    .dout(g198_n),
    .din1(G146_n_spl_001),
    .din2(g197_p)
  );


  LA
  g_g199_p
  (
    .dout(g199_p),
    .din1(G100_n),
    .din2(G145_p_spl_0011)
  );


  FA
  g_g199_n
  (
    .dout(g199_n),
    .din1(G100_p),
    .din2(G145_n_spl_0011)
  );


  LA
  g_g200_p
  (
    .dout(g200_p),
    .din1(G90_n),
    .din2(G145_n_spl_0011)
  );


  FA
  g_g200_n
  (
    .dout(g200_n),
    .din1(G90_p),
    .din2(G145_p_spl_0011)
  );


  LA
  g_g201_p
  (
    .dout(g201_p),
    .din1(g199_n),
    .din2(g200_n)
  );


  FA
  g_g201_n
  (
    .dout(g201_n),
    .din1(g199_p),
    .din2(g200_p)
  );


  LA
  g_g202_p
  (
    .dout(g202_p),
    .din1(G146_n_spl_001),
    .din2(g201_n)
  );


  FA
  g_g202_n
  (
    .dout(g202_n),
    .din1(G146_p_spl_001),
    .din2(g201_p)
  );


  LA
  g_g203_p
  (
    .dout(g203_p),
    .din1(g198_n),
    .din2(g202_n)
  );


  FA
  g_g203_n
  (
    .dout(g203_n),
    .din1(g198_p),
    .din2(g202_p)
  );


  LA
  g_g204_p
  (
    .dout(g204_p),
    .din1(G117_p_spl_0000),
    .din2(G120_n_spl_0000)
  );


  FA
  g_g204_n
  (
    .dout(g204_n),
    .din1(G117_n_spl_0000),
    .din2(G120_p_spl_0000)
  );


  LA
  g_g205_p
  (
    .dout(g205_p),
    .din1(G46_p),
    .din2(g204_p_spl_000)
  );


  FA
  g_g205_n
  (
    .dout(g205_n),
    .din1(G46_n),
    .din2(g204_n_spl_000)
  );


  LA
  g_g206_p
  (
    .dout(g206_p),
    .din1(G57_p),
    .din2(G117_n_spl_0000)
  );


  FA
  g_g206_n
  (
    .dout(g206_n),
    .din1(G57_n),
    .din2(G117_p_spl_0000)
  );


  LA
  g_g207_p
  (
    .dout(g207_p),
    .din1(G120_n_spl_0000),
    .din2(g206_n)
  );


  FA
  g_g207_n
  (
    .dout(g207_n),
    .din1(G120_p_spl_0000),
    .din2(g206_p)
  );


  LA
  g_g208_p
  (
    .dout(g208_p),
    .din1(G36_n),
    .din2(G117_n_spl_0001)
  );


  FA
  g_g208_n
  (
    .dout(g208_n),
    .din1(G36_p),
    .din2(G117_p_spl_0001)
  );


  LA
  g_g209_p
  (
    .dout(g209_p),
    .din1(G120_p_spl_0001),
    .din2(g208_p)
  );


  FA
  g_g209_n
  (
    .dout(g209_n),
    .din1(G120_n_spl_0001),
    .din2(g208_n)
  );


  LA
  g_g210_p
  (
    .dout(g210_p),
    .din1(G68_n),
    .din2(G117_p_spl_0001)
  );


  FA
  g_g210_n
  (
    .dout(g210_n),
    .din1(G68_p),
    .din2(G117_n_spl_0001)
  );


  LA
  g_g211_p
  (
    .dout(g211_p),
    .din1(g209_n),
    .din2(g210_n)
  );


  FA
  g_g211_n
  (
    .dout(g211_n),
    .din1(g209_p),
    .din2(g210_p)
  );


  LA
  g_g212_p
  (
    .dout(g212_p),
    .din1(g207_n),
    .din2(g211_p)
  );


  FA
  g_g212_n
  (
    .dout(g212_n),
    .din1(g207_p),
    .din2(g211_n)
  );


  LA
  g_g213_p
  (
    .dout(g213_p),
    .din1(g205_n),
    .din2(g212_n)
  );


  FA
  g_g213_n
  (
    .dout(g213_n),
    .din1(g205_p),
    .din2(g212_p)
  );


  LA
  g_g214_p
  (
    .dout(g214_p),
    .din1(G47_p),
    .din2(g204_p_spl_000)
  );


  FA
  g_g214_n
  (
    .dout(g214_n),
    .din1(G47_n),
    .din2(g204_n_spl_000)
  );


  LA
  g_g215_p
  (
    .dout(g215_p),
    .din1(G58_p),
    .din2(G117_n_spl_0010)
  );


  FA
  g_g215_n
  (
    .dout(g215_n),
    .din1(G58_n),
    .din2(G117_p_spl_0010)
  );


  LA
  g_g216_p
  (
    .dout(g216_p),
    .din1(G120_n_spl_0001),
    .din2(g215_n)
  );


  FA
  g_g216_n
  (
    .dout(g216_n),
    .din1(G120_p_spl_0001),
    .din2(g215_p)
  );


  LA
  g_g217_p
  (
    .dout(g217_p),
    .din1(G37_n),
    .din2(G117_n_spl_0010)
  );


  FA
  g_g217_n
  (
    .dout(g217_n),
    .din1(G37_p),
    .din2(G117_p_spl_0010)
  );


  LA
  g_g218_p
  (
    .dout(g218_p),
    .din1(G120_p_spl_0010),
    .din2(g217_p)
  );


  FA
  g_g218_n
  (
    .dout(g218_n),
    .din1(G120_n_spl_0010),
    .din2(g217_n)
  );


  LA
  g_g219_p
  (
    .dout(g219_p),
    .din1(G69_n),
    .din2(G117_p_spl_0011)
  );


  FA
  g_g219_n
  (
    .dout(g219_n),
    .din1(G69_p),
    .din2(G117_n_spl_0011)
  );


  LA
  g_g220_p
  (
    .dout(g220_p),
    .din1(g218_n),
    .din2(g219_n)
  );


  FA
  g_g220_n
  (
    .dout(g220_n),
    .din1(g218_p),
    .din2(g219_p)
  );


  LA
  g_g221_p
  (
    .dout(g221_p),
    .din1(g216_n),
    .din2(g220_p)
  );


  FA
  g_g221_n
  (
    .dout(g221_n),
    .din1(g216_p),
    .din2(g220_n)
  );


  LA
  g_g222_p
  (
    .dout(g222_p),
    .din1(g214_n),
    .din2(g221_n)
  );


  FA
  g_g222_n
  (
    .dout(g222_n),
    .din1(g214_p),
    .din2(g221_p)
  );


  LA
  g_g223_p
  (
    .dout(g223_p),
    .din1(G48_p),
    .din2(g204_p_spl_00)
  );


  FA
  g_g223_n
  (
    .dout(g223_n),
    .din1(G48_n),
    .din2(g204_n_spl_00)
  );


  LA
  g_g224_p
  (
    .dout(g224_p),
    .din1(G59_p),
    .din2(G117_n_spl_0011)
  );


  FA
  g_g224_n
  (
    .dout(g224_n),
    .din1(G59_n),
    .din2(G117_p_spl_0011)
  );


  LA
  g_g225_p
  (
    .dout(g225_p),
    .din1(G120_n_spl_0010),
    .din2(g224_n)
  );


  FA
  g_g225_n
  (
    .dout(g225_n),
    .din1(G120_p_spl_0010),
    .din2(g224_p)
  );


  LA
  g_g226_p
  (
    .dout(g226_p),
    .din1(G38_n),
    .din2(G117_n_spl_0100)
  );


  FA
  g_g226_n
  (
    .dout(g226_n),
    .din1(G38_p),
    .din2(G117_p_spl_0100)
  );


  LA
  g_g227_p
  (
    .dout(g227_p),
    .din1(G120_p_spl_0011),
    .din2(g226_p)
  );


  FA
  g_g227_n
  (
    .dout(g227_n),
    .din1(G120_n_spl_0011),
    .din2(g226_n)
  );


  LA
  g_g228_p
  (
    .dout(g228_p),
    .din1(G70_n),
    .din2(G117_p_spl_0100)
  );


  FA
  g_g228_n
  (
    .dout(g228_n),
    .din1(G70_p),
    .din2(G117_n_spl_0100)
  );


  LA
  g_g229_p
  (
    .dout(g229_p),
    .din1(g227_n),
    .din2(g228_n)
  );


  FA
  g_g229_n
  (
    .dout(g229_n),
    .din1(g227_p),
    .din2(g228_p)
  );


  LA
  g_g230_p
  (
    .dout(g230_p),
    .din1(g225_n),
    .din2(g229_p)
  );


  FA
  g_g230_n
  (
    .dout(g230_n),
    .din1(g225_p),
    .din2(g229_n)
  );


  LA
  g_g231_p
  (
    .dout(g231_p),
    .din1(g223_n),
    .din2(g230_n)
  );


  FA
  g_g231_n
  (
    .dout(g231_n),
    .din1(g223_p),
    .din2(g230_p)
  );


  LA
  g_g232_p
  (
    .dout(g232_p),
    .din1(G42_p),
    .din2(g204_p_spl_01)
  );


  FA
  g_g232_n
  (
    .dout(g232_n),
    .din1(G42_n),
    .din2(g204_n_spl_01)
  );


  LA
  g_g233_p
  (
    .dout(g233_p),
    .din1(G52_p),
    .din2(G117_n_spl_0101)
  );


  FA
  g_g233_n
  (
    .dout(g233_n),
    .din1(G52_n),
    .din2(G117_p_spl_0101)
  );


  LA
  g_g234_p
  (
    .dout(g234_p),
    .din1(G120_n_spl_0011),
    .din2(g233_n)
  );


  FA
  g_g234_n
  (
    .dout(g234_n),
    .din1(G120_p_spl_0011),
    .din2(g233_p)
  );


  LA
  g_g235_p
  (
    .dout(g235_p),
    .din1(G31_n),
    .din2(G117_n_spl_0101)
  );


  FA
  g_g235_n
  (
    .dout(g235_n),
    .din1(G31_p),
    .din2(G117_p_spl_0101)
  );


  LA
  g_g236_p
  (
    .dout(g236_p),
    .din1(G120_p_spl_0100),
    .din2(g235_p)
  );


  FA
  g_g236_n
  (
    .dout(g236_n),
    .din1(G120_n_spl_0100),
    .din2(g235_n)
  );


  LA
  g_g237_p
  (
    .dout(g237_p),
    .din1(G63_n),
    .din2(G117_p_spl_0110)
  );


  FA
  g_g237_n
  (
    .dout(g237_n),
    .din1(G63_p),
    .din2(G117_n_spl_0110)
  );


  LA
  g_g238_p
  (
    .dout(g238_p),
    .din1(g236_n),
    .din2(g237_n)
  );


  FA
  g_g238_n
  (
    .dout(g238_n),
    .din1(g236_p),
    .din2(g237_p)
  );


  LA
  g_g239_p
  (
    .dout(g239_p),
    .din1(g234_n),
    .din2(g238_p)
  );


  FA
  g_g239_n
  (
    .dout(g239_n),
    .din1(g234_p),
    .din2(g238_n)
  );


  LA
  g_g240_p
  (
    .dout(g240_p),
    .din1(g232_n),
    .din2(g239_n)
  );


  FA
  g_g240_n
  (
    .dout(g240_n),
    .din1(g232_p),
    .din2(g239_p)
  );


  FA
  g_g241_n
  (
    .dout(g241_n),
    .din1(G122_n_spl_0),
    .din2(g240_n_spl_00)
  );


  FA
  g_g242_n
  (
    .dout(g242_n),
    .din1(G116_n),
    .din2(g176_n_spl_0)
  );


  FA
  g_g243_n
  (
    .dout(g243_n),
    .din1(G121_p),
    .din2(g242_n)
  );


  FA
  g_g244_n
  (
    .dout(g244_n),
    .din1(G28_n),
    .din2(g243_n_spl_)
  );


  LA
  g_g245_p
  (
    .dout(g245_p),
    .din1(G1_p),
    .din2(G3_p)
  );


  FA
  g_g246_n
  (
    .dout(g246_n),
    .din1(g243_n_spl_),
    .din2(g245_p)
  );


  LA
  g_g247_p
  (
    .dout(g247_p),
    .din1(G49_p),
    .din2(g204_p_spl_01)
  );


  FA
  g_g247_n
  (
    .dout(g247_n),
    .din1(G49_n),
    .din2(g204_n_spl_01)
  );


  LA
  g_g248_p
  (
    .dout(g248_p),
    .din1(G60_p),
    .din2(G117_n_spl_0110)
  );


  FA
  g_g248_n
  (
    .dout(g248_n),
    .din1(G60_n),
    .din2(G117_p_spl_0110)
  );


  LA
  g_g249_p
  (
    .dout(g249_p),
    .din1(G120_n_spl_0100),
    .din2(g248_n)
  );


  FA
  g_g249_n
  (
    .dout(g249_n),
    .din1(G120_p_spl_0100),
    .din2(g248_p)
  );


  LA
  g_g250_p
  (
    .dout(g250_p),
    .din1(G39_n),
    .din2(G117_n_spl_0111)
  );


  FA
  g_g250_n
  (
    .dout(g250_n),
    .din1(G39_p),
    .din2(G117_p_spl_0111)
  );


  LA
  g_g251_p
  (
    .dout(g251_p),
    .din1(G120_p_spl_010),
    .din2(g250_p)
  );


  FA
  g_g251_n
  (
    .dout(g251_n),
    .din1(G120_n_spl_010),
    .din2(g250_n)
  );


  LA
  g_g252_p
  (
    .dout(g252_p),
    .din1(G71_n),
    .din2(G117_p_spl_0111)
  );


  FA
  g_g252_n
  (
    .dout(g252_n),
    .din1(G71_p),
    .din2(G117_n_spl_0111)
  );


  LA
  g_g253_p
  (
    .dout(g253_p),
    .din1(g251_n),
    .din2(g252_n)
  );


  FA
  g_g253_n
  (
    .dout(g253_n),
    .din1(g251_p),
    .din2(g252_p)
  );


  LA
  g_g254_p
  (
    .dout(g254_p),
    .din1(g249_n),
    .din2(g253_p)
  );


  FA
  g_g254_n
  (
    .dout(g254_n),
    .din1(g249_p),
    .din2(g253_n)
  );


  LA
  g_g255_p
  (
    .dout(g255_p),
    .din1(g247_n),
    .din2(g254_n)
  );


  FA
  g_g255_n
  (
    .dout(g255_n),
    .din1(g247_p),
    .din2(g254_p)
  );


  LA
  g_g256_p
  (
    .dout(g256_p),
    .din1(G35_n),
    .din2(G117_n_spl_1000)
  );


  FA
  g_g256_n
  (
    .dout(g256_n),
    .din1(G35_p),
    .din2(G117_p_spl_1000)
  );


  LA
  g_g257_p
  (
    .dout(g257_p),
    .din1(G67_n),
    .din2(G117_p_spl_1000)
  );


  FA
  g_g257_n
  (
    .dout(g257_n),
    .din1(G67_p),
    .din2(G117_n_spl_1000)
  );


  LA
  g_g258_p
  (
    .dout(g258_p),
    .din1(g256_n),
    .din2(g257_n)
  );


  FA
  g_g258_n
  (
    .dout(g258_n),
    .din1(g256_p),
    .din2(g257_p)
  );


  LA
  g_g259_p
  (
    .dout(g259_p),
    .din1(G120_p_spl_011),
    .din2(g258_n)
  );


  FA
  g_g259_n
  (
    .dout(g259_n),
    .din1(G120_n_spl_011),
    .din2(g258_p)
  );


  LA
  g_g260_p
  (
    .dout(g260_p),
    .din1(G56_n),
    .din2(G117_n_spl_1001)
  );


  FA
  g_g260_n
  (
    .dout(g260_n),
    .din1(G56_p),
    .din2(G117_p_spl_1001)
  );


  LA
  g_g261_p
  (
    .dout(g261_p),
    .din1(G120_n_spl_011),
    .din2(g260_p)
  );


  FA
  g_g261_n
  (
    .dout(g261_n),
    .din1(G120_p_spl_011),
    .din2(g260_n)
  );


  LA
  g_g262_p
  (
    .dout(g262_p),
    .din1(g259_n),
    .din2(g261_n)
  );


  FA
  g_g262_n
  (
    .dout(g262_n),
    .din1(g259_p),
    .din2(g261_p)
  );


  LA
  g_g263_p
  (
    .dout(g263_p),
    .din1(G45_p),
    .din2(g204_p_spl_10)
  );


  FA
  g_g263_n
  (
    .dout(g263_n),
    .din1(G45_n),
    .din2(g204_n_spl_10)
  );


  LA
  g_g264_p
  (
    .dout(g264_p),
    .din1(G55_p),
    .din2(G117_n_spl_1001)
  );


  FA
  g_g264_n
  (
    .dout(g264_n),
    .din1(G55_n),
    .din2(G117_p_spl_1001)
  );


  LA
  g_g265_p
  (
    .dout(g265_p),
    .din1(G120_n_spl_100),
    .din2(g264_n)
  );


  FA
  g_g265_n
  (
    .dout(g265_n),
    .din1(G120_p_spl_100),
    .din2(g264_p)
  );


  LA
  g_g266_p
  (
    .dout(g266_p),
    .din1(G34_n),
    .din2(G117_n_spl_1010)
  );


  FA
  g_g266_n
  (
    .dout(g266_n),
    .din1(G34_p),
    .din2(G117_p_spl_1010)
  );


  LA
  g_g267_p
  (
    .dout(g267_p),
    .din1(G120_p_spl_100),
    .din2(g266_p)
  );


  FA
  g_g267_n
  (
    .dout(g267_n),
    .din1(G120_n_spl_100),
    .din2(g266_n)
  );


  LA
  g_g268_p
  (
    .dout(g268_p),
    .din1(G66_n),
    .din2(G117_p_spl_1010)
  );


  FA
  g_g268_n
  (
    .dout(g268_n),
    .din1(G66_p),
    .din2(G117_n_spl_1010)
  );


  LA
  g_g269_p
  (
    .dout(g269_p),
    .din1(g267_n),
    .din2(g268_n)
  );


  FA
  g_g269_n
  (
    .dout(g269_n),
    .din1(g267_p),
    .din2(g268_p)
  );


  LA
  g_g270_p
  (
    .dout(g270_p),
    .din1(g265_n),
    .din2(g269_p)
  );


  FA
  g_g270_n
  (
    .dout(g270_n),
    .din1(g265_p),
    .din2(g269_n)
  );


  LA
  g_g271_p
  (
    .dout(g271_p),
    .din1(g263_n),
    .din2(g270_n)
  );


  FA
  g_g271_n
  (
    .dout(g271_n),
    .din1(g263_p),
    .din2(g270_p)
  );


  LA
  g_g272_p
  (
    .dout(g272_p),
    .din1(G44_p),
    .din2(g204_p_spl_10)
  );


  FA
  g_g272_n
  (
    .dout(g272_n),
    .din1(G44_n),
    .din2(g204_n_spl_10)
  );


  LA
  g_g273_p
  (
    .dout(g273_p),
    .din1(G54_p),
    .din2(G117_n_spl_1011)
  );


  FA
  g_g273_n
  (
    .dout(g273_n),
    .din1(G54_n),
    .din2(G117_p_spl_1011)
  );


  LA
  g_g274_p
  (
    .dout(g274_p),
    .din1(G120_n_spl_101),
    .din2(g273_n)
  );


  FA
  g_g274_n
  (
    .dout(g274_n),
    .din1(G120_p_spl_101),
    .din2(g273_p)
  );


  LA
  g_g275_p
  (
    .dout(g275_p),
    .din1(G33_n),
    .din2(G117_n_spl_1011)
  );


  FA
  g_g275_n
  (
    .dout(g275_n),
    .din1(G33_p),
    .din2(G117_p_spl_1011)
  );


  LA
  g_g276_p
  (
    .dout(g276_p),
    .din1(G120_p_spl_101),
    .din2(g275_p)
  );


  FA
  g_g276_n
  (
    .dout(g276_n),
    .din1(G120_n_spl_101),
    .din2(g275_n)
  );


  LA
  g_g277_p
  (
    .dout(g277_p),
    .din1(G65_n),
    .din2(G117_p_spl_1100)
  );


  FA
  g_g277_n
  (
    .dout(g277_n),
    .din1(G65_p),
    .din2(G117_n_spl_1100)
  );


  LA
  g_g278_p
  (
    .dout(g278_p),
    .din1(g276_n),
    .din2(g277_n)
  );


  FA
  g_g278_n
  (
    .dout(g278_n),
    .din1(g276_p),
    .din2(g277_p)
  );


  LA
  g_g279_p
  (
    .dout(g279_p),
    .din1(g274_n),
    .din2(g278_p)
  );


  FA
  g_g279_n
  (
    .dout(g279_n),
    .din1(g274_p),
    .din2(g278_n)
  );


  LA
  g_g280_p
  (
    .dout(g280_p),
    .din1(g272_n),
    .din2(g279_n)
  );


  FA
  g_g280_n
  (
    .dout(g280_n),
    .din1(g272_p),
    .din2(g279_p)
  );


  LA
  g_g281_p
  (
    .dout(g281_p),
    .din1(G123_p_spl_0),
    .din2(g231_n_spl_00)
  );


  LA
  g_g282_p
  (
    .dout(g282_p),
    .din1(G50_p),
    .din2(g204_p_spl_11)
  );


  FA
  g_g282_n
  (
    .dout(g282_n),
    .din1(G50_n),
    .din2(g204_n_spl_11)
  );


  LA
  g_g283_p
  (
    .dout(g283_p),
    .din1(G61_p),
    .din2(G117_n_spl_1100)
  );


  FA
  g_g283_n
  (
    .dout(g283_n),
    .din1(G61_n),
    .din2(G117_p_spl_1100)
  );


  LA
  g_g284_p
  (
    .dout(g284_p),
    .din1(G120_n_spl_110),
    .din2(g283_n)
  );


  FA
  g_g284_n
  (
    .dout(g284_n),
    .din1(G120_p_spl_110),
    .din2(g283_p)
  );


  LA
  g_g285_p
  (
    .dout(g285_p),
    .din1(G40_n),
    .din2(G117_n_spl_1101)
  );


  FA
  g_g285_n
  (
    .dout(g285_n),
    .din1(G40_p),
    .din2(G117_p_spl_1101)
  );


  LA
  g_g286_p
  (
    .dout(g286_p),
    .din1(G120_p_spl_110),
    .din2(g285_p)
  );


  FA
  g_g286_n
  (
    .dout(g286_n),
    .din1(G120_n_spl_110),
    .din2(g285_n)
  );


  LA
  g_g287_p
  (
    .dout(g287_p),
    .din1(G72_n),
    .din2(G117_p_spl_1101)
  );


  FA
  g_g287_n
  (
    .dout(g287_n),
    .din1(G72_p),
    .din2(G117_n_spl_1101)
  );


  LA
  g_g288_p
  (
    .dout(g288_p),
    .din1(g286_n),
    .din2(g287_n)
  );


  FA
  g_g288_n
  (
    .dout(g288_n),
    .din1(g286_p),
    .din2(g287_p)
  );


  LA
  g_g289_p
  (
    .dout(g289_p),
    .din1(g284_n),
    .din2(g288_p)
  );


  FA
  g_g289_n
  (
    .dout(g289_n),
    .din1(g284_p),
    .din2(g288_n)
  );


  LA
  g_g290_p
  (
    .dout(g290_p),
    .din1(g282_n),
    .din2(g289_n)
  );


  FA
  g_g290_n
  (
    .dout(g290_n),
    .din1(g282_p),
    .din2(g289_p)
  );


  LA
  g_g291_p
  (
    .dout(g291_p),
    .din1(G123_n_spl_0),
    .din2(g290_p_spl_00)
  );


  FA
  g_g292_n
  (
    .dout(g292_n),
    .din1(g281_p),
    .din2(g291_p)
  );


  LA
  g_g293_p
  (
    .dout(g293_p),
    .din1(G123_p_spl_0),
    .din2(g222_p_spl_00)
  );


  LA
  g_g294_p
  (
    .dout(g294_p),
    .din1(G123_n_spl_0),
    .din2(g255_n_spl_00)
  );


  FA
  g_g295_n
  (
    .dout(g295_n),
    .din1(g293_p),
    .din2(g294_p)
  );


  LA
  g_g296_p
  (
    .dout(g296_p),
    .din1(G118_p_spl_0),
    .din2(G122_n_spl_0)
  );


  FA
  g_g297_n
  (
    .dout(g297_n),
    .din1(g290_n_spl_00),
    .din2(g296_p)
  );


  LA
  g_g298_p
  (
    .dout(g298_p),
    .din1(G118_n_spl_),
    .din2(g290_p_spl_00)
  );


  FA
  g_g298_n
  (
    .dout(g298_n),
    .din1(G118_p_spl_0),
    .din2(g290_n_spl_00)
  );


  LA
  g_g299_p
  (
    .dout(g299_p),
    .din1(G123_p_spl_1),
    .din2(g298_p_spl_0)
  );


  LA
  g_g300_p
  (
    .dout(g300_p),
    .din1(G123_n_spl_1),
    .din2(g240_p_spl_0)
  );


  FA
  g_g301_n
  (
    .dout(g301_n),
    .din1(g299_p),
    .din2(g300_p)
  );


  LA
  g_g302_p
  (
    .dout(g302_p),
    .din1(G77_n),
    .din2(G145_n_spl_0100)
  );


  FA
  g_g302_n
  (
    .dout(g302_n),
    .din1(G77_p),
    .din2(G145_p_spl_0100)
  );


  LA
  g_g303_p
  (
    .dout(g303_p),
    .din1(G107_n),
    .din2(G145_p_spl_0100)
  );


  FA
  g_g303_n
  (
    .dout(g303_n),
    .din1(G107_p),
    .din2(G145_n_spl_0100)
  );


  LA
  g_g304_p
  (
    .dout(g304_p),
    .din1(g302_n),
    .din2(g303_n)
  );


  FA
  g_g304_n
  (
    .dout(g304_n),
    .din1(g302_p),
    .din2(g303_p)
  );


  LA
  g_g305_p
  (
    .dout(g305_p),
    .din1(G146_p_spl_010),
    .din2(g304_n)
  );


  FA
  g_g305_n
  (
    .dout(g305_n),
    .din1(G146_n_spl_010),
    .din2(g304_p)
  );


  LA
  g_g306_p
  (
    .dout(g306_p),
    .din1(G97_n),
    .din2(G145_p_spl_0101)
  );


  FA
  g_g306_n
  (
    .dout(g306_n),
    .din1(G97_p),
    .din2(G145_n_spl_0101)
  );


  LA
  g_g307_p
  (
    .dout(g307_p),
    .din1(G87_n),
    .din2(G145_n_spl_0101)
  );


  FA
  g_g307_n
  (
    .dout(g307_n),
    .din1(G87_p),
    .din2(G145_p_spl_0101)
  );


  LA
  g_g308_p
  (
    .dout(g308_p),
    .din1(g306_n),
    .din2(g307_n)
  );


  FA
  g_g308_n
  (
    .dout(g308_n),
    .din1(g306_p),
    .din2(g307_p)
  );


  LA
  g_g309_p
  (
    .dout(g309_p),
    .din1(G146_n_spl_010),
    .din2(g308_n)
  );


  FA
  g_g309_n
  (
    .dout(g309_n),
    .din1(G146_p_spl_010),
    .din2(g308_p)
  );


  LA
  g_g310_p
  (
    .dout(g310_p),
    .din1(g305_n),
    .din2(g309_n)
  );


  FA
  g_g310_n
  (
    .dout(g310_n),
    .din1(g305_p),
    .din2(g309_p)
  );


  FA
  g_g311_n
  (
    .dout(g311_n),
    .din1(G143_n_spl_0),
    .din2(g310_p_spl_0)
  );


  FA
  g_g312_n
  (
    .dout(g312_n),
    .din1(G143_p_spl_0),
    .din2(g310_n_spl_0)
  );


  LA
  g_g313_p
  (
    .dout(g313_p),
    .din1(g311_n),
    .din2(g312_n)
  );


  FA
  g_g314_n
  (
    .dout(g314_n),
    .din1(G144_p_spl_0),
    .din2(g313_p)
  );


  LA
  g_g315_p
  (
    .dout(g315_p),
    .din1(G154_n_spl_),
    .din2(G155_n_spl_)
  );


  FA
  g_g315_n
  (
    .dout(g315_n),
    .din1(G154_p_spl_),
    .din2(G155_p_spl_)
  );


  LA
  g_g316_p
  (
    .dout(g316_p),
    .din1(G154_p_spl_),
    .din2(G155_p_spl_)
  );


  FA
  g_g316_n
  (
    .dout(g316_n),
    .din1(G154_n_spl_),
    .din2(G155_n_spl_)
  );


  LA
  g_g317_p
  (
    .dout(g317_p),
    .din1(g315_n),
    .din2(g316_n)
  );


  FA
  g_g317_n
  (
    .dout(g317_n),
    .din1(g315_p),
    .din2(g316_p)
  );


  LA
  g_g318_p
  (
    .dout(g318_p),
    .din1(G125_n_spl_0),
    .din2(G126_n_spl_0)
  );


  FA
  g_g318_n
  (
    .dout(g318_n),
    .din1(G125_p_spl_0),
    .din2(G126_p_spl_0)
  );


  LA
  g_g319_p
  (
    .dout(g319_p),
    .din1(G125_p_spl_0),
    .din2(G126_p_spl_0)
  );


  FA
  g_g319_n
  (
    .dout(g319_n),
    .din1(G125_n_spl_0),
    .din2(G126_n_spl_0)
  );


  LA
  g_g320_p
  (
    .dout(g320_p),
    .din1(g318_n),
    .din2(g319_n)
  );


  FA
  g_g320_n
  (
    .dout(g320_n),
    .din1(g318_p),
    .din2(g319_p)
  );


  LA
  g_g321_p
  (
    .dout(g321_p),
    .din1(g317_p_spl_),
    .din2(g320_n_spl_)
  );


  FA
  g_g321_n
  (
    .dout(g321_n),
    .din1(g317_n_spl_),
    .din2(g320_p_spl_)
  );


  LA
  g_g322_p
  (
    .dout(g322_p),
    .din1(g317_n_spl_),
    .din2(g320_p_spl_)
  );


  FA
  g_g322_n
  (
    .dout(g322_n),
    .din1(g317_p_spl_),
    .din2(g320_n_spl_)
  );


  LA
  g_g323_p
  (
    .dout(g323_p),
    .din1(g321_n),
    .din2(g322_n)
  );


  FA
  g_g323_n
  (
    .dout(g323_n),
    .din1(g321_p),
    .din2(g322_p)
  );


  LA
  g_g324_p
  (
    .dout(g324_p),
    .din1(G152_n_spl_),
    .din2(G153_n_spl_)
  );


  FA
  g_g324_n
  (
    .dout(g324_n),
    .din1(G152_p_spl_),
    .din2(G153_p_spl_)
  );


  LA
  g_g325_p
  (
    .dout(g325_p),
    .din1(G152_p_spl_),
    .din2(G153_p_spl_)
  );


  FA
  g_g325_n
  (
    .dout(g325_n),
    .din1(G152_n_spl_),
    .din2(G153_n_spl_)
  );


  LA
  g_g326_p
  (
    .dout(g326_p),
    .din1(g324_n),
    .din2(g325_n)
  );


  FA
  g_g326_n
  (
    .dout(g326_n),
    .din1(g324_p),
    .din2(g325_p)
  );


  LA
  g_g327_p
  (
    .dout(g327_p),
    .din1(G148_n_spl_),
    .din2(G149_n_spl_)
  );


  FA
  g_g327_n
  (
    .dout(g327_n),
    .din1(G148_p_spl_),
    .din2(G149_p_spl_)
  );


  LA
  g_g328_p
  (
    .dout(g328_p),
    .din1(G148_p_spl_),
    .din2(G149_p_spl_)
  );


  FA
  g_g328_n
  (
    .dout(g328_n),
    .din1(G148_n_spl_),
    .din2(G149_n_spl_)
  );


  LA
  g_g329_p
  (
    .dout(g329_p),
    .din1(g327_n),
    .din2(g328_n)
  );


  FA
  g_g329_n
  (
    .dout(g329_n),
    .din1(g327_p),
    .din2(g328_p)
  );


  LA
  g_g330_p
  (
    .dout(g330_p),
    .din1(g326_n_spl_),
    .din2(g329_n_spl_)
  );


  FA
  g_g330_n
  (
    .dout(g330_n),
    .din1(g326_p_spl_),
    .din2(g329_p_spl_)
  );


  LA
  g_g331_p
  (
    .dout(g331_p),
    .din1(g326_p_spl_),
    .din2(g329_p_spl_)
  );


  FA
  g_g331_n
  (
    .dout(g331_n),
    .din1(g326_n_spl_),
    .din2(g329_n_spl_)
  );


  LA
  g_g332_p
  (
    .dout(g332_p),
    .din1(g330_n),
    .din2(g331_n)
  );


  FA
  g_g332_n
  (
    .dout(g332_n),
    .din1(g330_p),
    .din2(g331_p)
  );


  LA
  g_g333_p
  (
    .dout(g333_p),
    .din1(G150_n_spl_),
    .din2(G151_n_spl_)
  );


  FA
  g_g333_n
  (
    .dout(g333_n),
    .din1(G150_p_spl_),
    .din2(G151_p_spl_)
  );


  LA
  g_g334_p
  (
    .dout(g334_p),
    .din1(G150_p_spl_),
    .din2(G151_p_spl_)
  );


  FA
  g_g334_n
  (
    .dout(g334_n),
    .din1(G150_n_spl_),
    .din2(G151_n_spl_)
  );


  LA
  g_g335_p
  (
    .dout(g335_p),
    .din1(g333_n),
    .din2(g334_n)
  );


  FA
  g_g335_n
  (
    .dout(g335_n),
    .din1(g333_p),
    .din2(g334_p)
  );


  LA
  g_g336_p
  (
    .dout(g336_p),
    .din1(g332_n_spl_),
    .din2(g335_n_spl_)
  );


  FA
  g_g336_n
  (
    .dout(g336_n),
    .din1(g332_p_spl_),
    .din2(g335_p_spl_)
  );


  LA
  g_g337_p
  (
    .dout(g337_p),
    .din1(g332_p_spl_),
    .din2(g335_p_spl_)
  );


  FA
  g_g337_n
  (
    .dout(g337_n),
    .din1(g332_n_spl_),
    .din2(g335_n_spl_)
  );


  LA
  g_g338_p
  (
    .dout(g338_p),
    .din1(g336_n),
    .din2(g337_n)
  );


  FA
  g_g338_n
  (
    .dout(g338_n),
    .din1(g336_p),
    .din2(g337_p)
  );


  FA
  g_g339_n
  (
    .dout(g339_n),
    .din1(g323_n),
    .din2(g338_p)
  );


  FA
  g_g340_n
  (
    .dout(g340_n),
    .din1(g323_p),
    .din2(g338_n)
  );


  LA
  g_g341_p
  (
    .dout(g341_p),
    .din1(G10_p),
    .din2(g340_n)
  );


  LA
  g_g342_p
  (
    .dout(g342_p),
    .din1(g339_n),
    .din2(g341_p)
  );


  LA
  g_g343_p
  (
    .dout(g343_p),
    .din1(G141_n_spl_0),
    .din2(G142_n_spl_0)
  );


  FA
  g_g343_n
  (
    .dout(g343_n),
    .din1(G141_p_spl_0),
    .din2(G142_p_spl_0)
  );


  LA
  g_g344_p
  (
    .dout(g344_p),
    .din1(g158_n_spl_),
    .din2(g343_n)
  );


  FA
  g_g344_n
  (
    .dout(g344_n),
    .din1(g158_p),
    .din2(g343_p)
  );


  LA
  g_g345_p
  (
    .dout(g345_p),
    .din1(G139_n_spl_0),
    .din2(G140_n_spl_0)
  );


  FA
  g_g345_n
  (
    .dout(g345_n),
    .din1(G139_p_spl_0),
    .din2(G140_p_spl_0)
  );


  LA
  g_g346_p
  (
    .dout(g346_p),
    .din1(g159_n_spl_),
    .din2(g345_n)
  );


  FA
  g_g346_n
  (
    .dout(g346_n),
    .din1(g159_p),
    .din2(g345_p)
  );


  LA
  g_g347_p
  (
    .dout(g347_p),
    .din1(G138_p_spl_00),
    .din2(G157_n_spl_)
  );


  FA
  g_g347_n
  (
    .dout(g347_n),
    .din1(G138_n_spl_0),
    .din2(G157_p_spl_)
  );


  LA
  g_g348_p
  (
    .dout(g348_p),
    .din1(G138_n_spl_0),
    .din2(G157_p_spl_)
  );


  FA
  g_g348_n
  (
    .dout(g348_n),
    .din1(G138_p_spl_00),
    .din2(G157_n_spl_)
  );


  LA
  g_g349_p
  (
    .dout(g349_p),
    .din1(g347_n),
    .din2(g348_n)
  );


  FA
  g_g349_n
  (
    .dout(g349_n),
    .din1(g347_p),
    .din2(g348_p)
  );


  LA
  g_g350_p
  (
    .dout(g350_p),
    .din1(g346_n_spl_),
    .din2(g349_n_spl_)
  );


  FA
  g_g350_n
  (
    .dout(g350_n),
    .din1(g346_p_spl_),
    .din2(g349_p_spl_)
  );


  LA
  g_g351_p
  (
    .dout(g351_p),
    .din1(g346_p_spl_),
    .din2(g349_p_spl_)
  );


  FA
  g_g351_n
  (
    .dout(g351_n),
    .din1(g346_n_spl_),
    .din2(g349_n_spl_)
  );


  LA
  g_g352_p
  (
    .dout(g352_p),
    .din1(g350_n),
    .din2(g351_n)
  );


  FA
  g_g352_n
  (
    .dout(g352_n),
    .din1(g350_p),
    .din2(g351_p)
  );


  LA
  g_g353_p
  (
    .dout(g353_p),
    .din1(g344_n_spl_),
    .din2(g352_n_spl_)
  );


  FA
  g_g353_n
  (
    .dout(g353_n),
    .din1(g344_p_spl_),
    .din2(g352_p_spl_)
  );


  LA
  g_g354_p
  (
    .dout(g354_p),
    .din1(g344_p_spl_),
    .din2(g352_p_spl_)
  );


  FA
  g_g354_n
  (
    .dout(g354_n),
    .din1(g344_n_spl_),
    .din2(g352_n_spl_)
  );


  LA
  g_g355_p
  (
    .dout(g355_p),
    .din1(g353_n),
    .din2(g354_n)
  );


  FA
  g_g355_n
  (
    .dout(g355_n),
    .din1(g353_p),
    .din2(g354_p)
  );


  LA
  g_g356_p
  (
    .dout(g356_p),
    .din1(G143_n_spl_0),
    .din2(G144_n_spl_)
  );


  FA
  g_g356_n
  (
    .dout(g356_n),
    .din1(G143_p_spl_0),
    .din2(G144_p_spl_0)
  );


  LA
  g_g357_p
  (
    .dout(g357_p),
    .din1(G143_p_spl_),
    .din2(G144_p_spl_)
  );


  FA
  g_g357_n
  (
    .dout(g357_n),
    .din1(G143_n_spl_),
    .din2(G144_n_spl_)
  );


  LA
  g_g358_p
  (
    .dout(g358_p),
    .din1(g356_n),
    .din2(g357_n)
  );


  FA
  g_g358_n
  (
    .dout(g358_n),
    .din1(g356_p),
    .din2(g357_p)
  );


  FA
  g_g359_n
  (
    .dout(g359_n),
    .din1(g355_n),
    .din2(g358_n)
  );


  FA
  g_g360_n
  (
    .dout(g360_n),
    .din1(g355_p),
    .din2(g358_p)
  );


  LA
  g_g361_p
  (
    .dout(g361_p),
    .din1(g359_n),
    .din2(g360_n)
  );


  LA
  g_g362_p
  (
    .dout(g362_p),
    .din1(G133_n_spl_0),
    .din2(G134_n_spl_0)
  );


  FA
  g_g362_n
  (
    .dout(g362_n),
    .din1(G133_p_spl_0),
    .din2(G134_p_spl_0)
  );


  LA
  g_g363_p
  (
    .dout(g363_p),
    .din1(G133_p_spl_0),
    .din2(G134_p_spl_0)
  );


  FA
  g_g363_n
  (
    .dout(g363_n),
    .din1(G133_n_spl_0),
    .din2(G134_n_spl_0)
  );


  LA
  g_g364_p
  (
    .dout(g364_p),
    .din1(g362_n),
    .din2(g363_n)
  );


  FA
  g_g364_n
  (
    .dout(g364_n),
    .din1(g362_p),
    .din2(g363_p)
  );


  LA
  g_g365_p
  (
    .dout(g365_p),
    .din1(G135_n_spl_0),
    .din2(G136_n_spl_0)
  );


  FA
  g_g365_n
  (
    .dout(g365_n),
    .din1(G135_p_spl_0),
    .din2(G136_p_spl_00)
  );


  LA
  g_g366_p
  (
    .dout(g366_p),
    .din1(G135_p_spl_0),
    .din2(G136_p_spl_00)
  );


  FA
  g_g366_n
  (
    .dout(g366_n),
    .din1(G135_n_spl_0),
    .din2(G136_n_spl_0)
  );


  LA
  g_g367_p
  (
    .dout(g367_p),
    .din1(g365_n),
    .din2(g366_n)
  );


  FA
  g_g367_n
  (
    .dout(g367_n),
    .din1(g365_p),
    .din2(g366_p)
  );


  LA
  g_g368_p
  (
    .dout(g368_p),
    .din1(g364_p_spl_),
    .din2(g367_n_spl_)
  );


  FA
  g_g368_n
  (
    .dout(g368_n),
    .din1(g364_n_spl_),
    .din2(g367_p_spl_)
  );


  LA
  g_g369_p
  (
    .dout(g369_p),
    .din1(g364_n_spl_),
    .din2(g367_p_spl_)
  );


  FA
  g_g369_n
  (
    .dout(g369_n),
    .din1(g364_p_spl_),
    .din2(g367_n_spl_)
  );


  LA
  g_g370_p
  (
    .dout(g370_p),
    .din1(g368_n),
    .din2(g369_n)
  );


  FA
  g_g370_n
  (
    .dout(g370_n),
    .din1(g368_p),
    .din2(g369_p)
  );


  LA
  g_g371_p
  (
    .dout(g371_p),
    .din1(G131_n_spl_0),
    .din2(G132_n_spl_0)
  );


  FA
  g_g371_n
  (
    .dout(g371_n),
    .din1(G131_p_spl_0),
    .din2(G132_p_spl_0)
  );


  LA
  g_g372_p
  (
    .dout(g372_p),
    .din1(G131_p_spl_0),
    .din2(G132_p_spl_0)
  );


  FA
  g_g372_n
  (
    .dout(g372_n),
    .din1(G131_n_spl_0),
    .din2(G132_n_spl_0)
  );


  LA
  g_g373_p
  (
    .dout(g373_p),
    .din1(g371_n),
    .din2(g372_n)
  );


  FA
  g_g373_n
  (
    .dout(g373_n),
    .din1(g371_p),
    .din2(g372_p)
  );


  LA
  g_g374_p
  (
    .dout(g374_p),
    .din1(G128_p_spl_0),
    .din2(G156_n_spl_)
  );


  FA
  g_g374_n
  (
    .dout(g374_n),
    .din1(G128_n_spl_0),
    .din2(G156_p_spl_)
  );


  LA
  g_g375_p
  (
    .dout(g375_p),
    .din1(G128_n_spl_0),
    .din2(G156_p_spl_)
  );


  FA
  g_g375_n
  (
    .dout(g375_n),
    .din1(G128_p_spl_0),
    .din2(G156_n_spl_)
  );


  LA
  g_g376_p
  (
    .dout(g376_p),
    .din1(g374_n),
    .din2(g375_n)
  );


  FA
  g_g376_n
  (
    .dout(g376_n),
    .din1(g374_p),
    .din2(g375_p)
  );


  LA
  g_g377_p
  (
    .dout(g377_p),
    .din1(g373_n_spl_),
    .din2(g376_n_spl_)
  );


  FA
  g_g377_n
  (
    .dout(g377_n),
    .din1(g373_p_spl_),
    .din2(g376_p_spl_)
  );


  LA
  g_g378_p
  (
    .dout(g378_p),
    .din1(g373_p_spl_),
    .din2(g376_p_spl_)
  );


  FA
  g_g378_n
  (
    .dout(g378_n),
    .din1(g373_n_spl_),
    .din2(g376_n_spl_)
  );


  LA
  g_g379_p
  (
    .dout(g379_p),
    .din1(g377_n),
    .din2(g378_n)
  );


  FA
  g_g379_n
  (
    .dout(g379_n),
    .din1(g377_p),
    .din2(g378_p)
  );


  LA
  g_g380_p
  (
    .dout(g380_p),
    .din1(G129_n_spl_0),
    .din2(G130_n_spl_0)
  );


  FA
  g_g380_n
  (
    .dout(g380_n),
    .din1(G129_p_spl_0),
    .din2(G130_p_spl_0)
  );


  LA
  g_g381_p
  (
    .dout(g381_p),
    .din1(G129_p_spl_0),
    .din2(G130_p_spl_0)
  );


  FA
  g_g381_n
  (
    .dout(g381_n),
    .din1(G129_n_spl_0),
    .din2(G130_n_spl_0)
  );


  LA
  g_g382_p
  (
    .dout(g382_p),
    .din1(g380_n),
    .din2(g381_n)
  );


  FA
  g_g382_n
  (
    .dout(g382_n),
    .din1(g380_p),
    .din2(g381_p)
  );


  LA
  g_g383_p
  (
    .dout(g383_p),
    .din1(g379_n_spl_),
    .din2(g382_n_spl_)
  );


  FA
  g_g383_n
  (
    .dout(g383_n),
    .din1(g379_p_spl_),
    .din2(g382_p_spl_)
  );


  LA
  g_g384_p
  (
    .dout(g384_p),
    .din1(g379_p_spl_),
    .din2(g382_p_spl_)
  );


  FA
  g_g384_n
  (
    .dout(g384_n),
    .din1(g379_n_spl_),
    .din2(g382_n_spl_)
  );


  LA
  g_g385_p
  (
    .dout(g385_p),
    .din1(g383_n),
    .din2(g384_n)
  );


  FA
  g_g385_n
  (
    .dout(g385_n),
    .din1(g383_p),
    .din2(g384_p)
  );


  FA
  g_g386_n
  (
    .dout(g386_n),
    .din1(g370_p),
    .din2(g385_n)
  );


  FA
  g_g387_n
  (
    .dout(g387_n),
    .din1(g370_n),
    .din2(g385_p)
  );


  LA
  g_g388_p
  (
    .dout(g388_p),
    .din1(g386_n),
    .din2(g387_n)
  );


  LA
  g_g389_p
  (
    .dout(g389_p),
    .din1(G12_n_spl_0000),
    .din2(g222_p_spl_00)
  );


  FA
  g_g389_n
  (
    .dout(g389_n),
    .din1(G12_p_spl_0000),
    .din2(g222_n_spl_0)
  );


  LA
  g_g390_p
  (
    .dout(g390_p),
    .din1(G12_p_spl_0000),
    .din2(G15_n)
  );


  FA
  g_g390_n
  (
    .dout(g390_n),
    .din1(G12_n_spl_0000),
    .din2(G15_p)
  );


  LA
  g_g391_p
  (
    .dout(g391_p),
    .din1(g389_n),
    .din2(g390_n)
  );


  FA
  g_g391_n
  (
    .dout(g391_n),
    .din1(g389_p),
    .din2(g390_p)
  );


  LA
  g_g392_p
  (
    .dout(g392_p),
    .din1(G130_p_spl_1),
    .din2(g391_n)
  );


  LA
  g_g393_p
  (
    .dout(g393_p),
    .din1(G12_n_spl_0001),
    .din2(g231_p_spl_00)
  );


  FA
  g_g393_n
  (
    .dout(g393_n),
    .din1(G12_p_spl_0001),
    .din2(g231_n_spl_00)
  );


  LA
  g_g394_p
  (
    .dout(g394_p),
    .din1(G5_n),
    .din2(G12_p_spl_0001)
  );


  FA
  g_g394_n
  (
    .dout(g394_n),
    .din1(G5_p),
    .din2(G12_n_spl_0001)
  );


  LA
  g_g395_p
  (
    .dout(g395_p),
    .din1(g393_n),
    .din2(g394_n)
  );


  FA
  g_g395_n
  (
    .dout(g395_n),
    .din1(g393_p),
    .din2(g394_p)
  );


  LA
  g_g396_p
  (
    .dout(g396_p),
    .din1(G129_n_spl_),
    .din2(g395_p)
  );


  FA
  g_g397_n
  (
    .dout(g397_n),
    .din1(g392_p),
    .din2(g396_p)
  );


  LA
  g_g398_p
  (
    .dout(g398_p),
    .din1(G12_n_spl_001),
    .din2(g213_p_spl_00)
  );


  FA
  g_g398_n
  (
    .dout(g398_n),
    .din1(G12_p_spl_001),
    .din2(g213_n_spl_0)
  );


  LA
  g_g399_p
  (
    .dout(g399_p),
    .din1(G12_p_spl_001),
    .din2(G16_n)
  );


  FA
  g_g399_n
  (
    .dout(g399_n),
    .din1(G12_n_spl_001),
    .din2(G16_p)
  );


  LA
  g_g400_p
  (
    .dout(g400_p),
    .din1(g398_n),
    .din2(g399_n)
  );


  FA
  g_g400_n
  (
    .dout(g400_n),
    .din1(g398_p),
    .din2(g399_p)
  );


  LA
  g_g401_p
  (
    .dout(g401_p),
    .din1(G131_n_spl_),
    .din2(g400_p)
  );


  FA
  g_g402_n
  (
    .dout(g402_n),
    .din1(G22_n),
    .din2(G23_n_spl_000)
  );


  FA
  g_g403_n
  (
    .dout(g403_n),
    .din1(G23_p_spl_000),
    .din2(g310_n_spl_0)
  );


  LA
  g_g404_p
  (
    .dout(g404_p),
    .din1(g402_n),
    .din2(g403_n)
  );


  FA
  g_g405_n
  (
    .dout(g405_n),
    .din1(g401_p),
    .din2(g404_p)
  );


  FA
  g_g406_n
  (
    .dout(g406_n),
    .din1(G9_n),
    .din2(g405_n)
  );


  LA
  g_g407_p
  (
    .dout(g407_p),
    .din1(G23_n_spl_000),
    .din2(g185_n_spl_00)
  );


  FA
  g_g407_n
  (
    .dout(g407_n),
    .din1(G23_p_spl_000),
    .din2(g185_p_spl_0)
  );


  LA
  g_g408_p
  (
    .dout(g408_p),
    .din1(G23_p_spl_001),
    .din2(G26_n)
  );


  FA
  g_g408_n
  (
    .dout(g408_n),
    .din1(G23_n_spl_001),
    .din2(G26_p)
  );


  LA
  g_g409_p
  (
    .dout(g409_p),
    .din1(g407_n),
    .din2(g408_n)
  );


  FA
  g_g409_n
  (
    .dout(g409_n),
    .din1(g407_p),
    .din2(g408_p)
  );


  LA
  g_g410_p
  (
    .dout(g410_p),
    .din1(G141_p_spl_1),
    .din2(g409_n)
  );


  LA
  g_g411_p
  (
    .dout(g411_p),
    .din1(G23_n_spl_001),
    .din2(g203_n_spl_00)
  );


  FA
  g_g411_n
  (
    .dout(g411_n),
    .din1(G23_p_spl_001),
    .din2(g203_p_spl_0)
  );


  LA
  g_g412_p
  (
    .dout(g412_p),
    .din1(G21_n),
    .din2(G23_p_spl_010)
  );


  FA
  g_g412_n
  (
    .dout(g412_n),
    .din1(G21_p),
    .din2(G23_n_spl_010)
  );


  LA
  g_g413_p
  (
    .dout(g413_p),
    .din1(g411_n),
    .din2(g412_n)
  );


  FA
  g_g413_n
  (
    .dout(g413_n),
    .din1(g411_p),
    .din2(g412_p)
  );


  LA
  g_g414_p
  (
    .dout(g414_p),
    .din1(G140_p_spl_1),
    .din2(g413_n)
  );


  LA
  g_g415_p
  (
    .dout(g415_p),
    .din1(G141_n_spl_),
    .din2(g409_p)
  );


  FA
  g_g416_n
  (
    .dout(g416_n),
    .din1(g414_p),
    .din2(g415_p)
  );


  FA
  g_g417_n
  (
    .dout(g417_n),
    .din1(g410_p),
    .din2(g416_n)
  );


  LA
  g_g418_p
  (
    .dout(g418_p),
    .din1(G140_n_spl_),
    .din2(g413_p)
  );


  LA
  g_g419_p
  (
    .dout(g419_p),
    .din1(G83_n),
    .din2(G145_n_spl_0110)
  );


  FA
  g_g419_n
  (
    .dout(g419_n),
    .din1(G83_p),
    .din2(G145_p_spl_0110)
  );


  LA
  g_g420_p
  (
    .dout(g420_p),
    .din1(G113_n),
    .din2(G145_p_spl_0110)
  );


  FA
  g_g420_n
  (
    .dout(g420_n),
    .din1(G113_p),
    .din2(G145_n_spl_0110)
  );


  LA
  g_g421_p
  (
    .dout(g421_p),
    .din1(g419_n),
    .din2(g420_n)
  );


  FA
  g_g421_n
  (
    .dout(g421_n),
    .din1(g419_p),
    .din2(g420_p)
  );


  LA
  g_g422_p
  (
    .dout(g422_p),
    .din1(G146_p_spl_011),
    .din2(g421_n)
  );


  FA
  g_g422_n
  (
    .dout(g422_n),
    .din1(G146_n_spl_011),
    .din2(g421_p)
  );


  LA
  g_g423_p
  (
    .dout(g423_p),
    .din1(G103_n),
    .din2(G145_p_spl_0111)
  );


  FA
  g_g423_n
  (
    .dout(g423_n),
    .din1(G103_p),
    .din2(G145_n_spl_0111)
  );


  LA
  g_g424_p
  (
    .dout(g424_p),
    .din1(G93_n),
    .din2(G145_n_spl_0111)
  );


  FA
  g_g424_n
  (
    .dout(g424_n),
    .din1(G93_p),
    .din2(G145_p_spl_0111)
  );


  LA
  g_g425_p
  (
    .dout(g425_p),
    .din1(g423_n),
    .din2(g424_n)
  );


  FA
  g_g425_n
  (
    .dout(g425_n),
    .din1(g423_p),
    .din2(g424_p)
  );


  LA
  g_g426_p
  (
    .dout(g426_p),
    .din1(G146_n_spl_011),
    .din2(g425_n)
  );


  FA
  g_g426_n
  (
    .dout(g426_n),
    .din1(G146_p_spl_011),
    .din2(g425_p)
  );


  LA
  g_g427_p
  (
    .dout(g427_p),
    .din1(g422_n),
    .din2(g426_n)
  );


  FA
  g_g427_n
  (
    .dout(g427_n),
    .din1(g422_p),
    .din2(g426_p)
  );


  LA
  g_g428_p
  (
    .dout(g428_p),
    .din1(G23_n_spl_010),
    .din2(g427_n_spl_0)
  );


  FA
  g_g428_n
  (
    .dout(g428_n),
    .din1(G23_p_spl_010),
    .din2(g427_p_spl_0)
  );


  LA
  g_g429_p
  (
    .dout(g429_p),
    .din1(G23_p_spl_011),
    .din2(G24_n)
  );


  FA
  g_g429_n
  (
    .dout(g429_n),
    .din1(G23_n_spl_011),
    .din2(G24_p)
  );


  LA
  g_g430_p
  (
    .dout(g430_p),
    .din1(g428_n),
    .din2(g429_n)
  );


  FA
  g_g430_n
  (
    .dout(g430_n),
    .din1(g428_p),
    .din2(g429_p)
  );


  LA
  g_g431_p
  (
    .dout(g431_p),
    .din1(G136_n_spl_1),
    .din2(g430_p)
  );


  LA
  g_g432_p
  (
    .dout(g432_p),
    .din1(G136_p_spl_0),
    .din2(g430_n)
  );


  FA
  g_g433_n
  (
    .dout(g433_n),
    .din1(g431_p),
    .din2(g432_p)
  );


  FA
  g_g434_n
  (
    .dout(g434_n),
    .din1(g418_p),
    .din2(g433_n)
  );


  FA
  g_g435_n
  (
    .dout(g435_n),
    .din1(g417_n),
    .din2(g434_n)
  );


  FA
  g_g436_n
  (
    .dout(g436_n),
    .din1(g406_n),
    .din2(g435_n)
  );


  FA
  g_g437_n
  (
    .dout(g437_n),
    .din1(g397_n),
    .din2(g436_n)
  );


  LA
  g_g438_p
  (
    .dout(g438_p),
    .din1(G12_n_spl_010),
    .din2(g255_p_spl_00)
  );


  FA
  g_g438_n
  (
    .dout(g438_n),
    .din1(G12_p_spl_010),
    .din2(g255_n_spl_00)
  );


  LA
  g_g439_p
  (
    .dout(g439_p),
    .din1(G12_p_spl_010),
    .din2(G14_n)
  );


  FA
  g_g439_n
  (
    .dout(g439_n),
    .din1(G12_n_spl_010),
    .din2(G14_p)
  );


  LA
  g_g440_p
  (
    .dout(g440_p),
    .din1(g438_n),
    .din2(g439_n)
  );


  FA
  g_g440_n
  (
    .dout(g440_n),
    .din1(g438_p),
    .din2(g439_p)
  );


  LA
  g_g441_p
  (
    .dout(g441_p),
    .din1(G128_p_spl_1),
    .din2(g440_n)
  );


  LA
  g_g442_p
  (
    .dout(g442_p),
    .din1(G130_n_spl_),
    .din2(g391_p)
  );


  FA
  g_g443_n
  (
    .dout(g443_n),
    .din1(g441_p),
    .din2(g442_p)
  );


  LA
  g_g444_p
  (
    .dout(g444_p),
    .din1(G131_p_spl_1),
    .din2(g400_n)
  );


  LA
  g_g445_p
  (
    .dout(g445_p),
    .din1(G12_n_spl_011),
    .din2(g262_n_spl_0)
  );


  FA
  g_g445_n
  (
    .dout(g445_n),
    .din1(G12_p_spl_011),
    .din2(g262_p_spl_0)
  );


  LA
  g_g446_p
  (
    .dout(g446_p),
    .din1(G12_p_spl_011),
    .din2(G17_n)
  );


  FA
  g_g446_n
  (
    .dout(g446_n),
    .din1(G12_n_spl_011),
    .din2(G17_p)
  );


  LA
  g_g447_p
  (
    .dout(g447_p),
    .din1(g445_n),
    .din2(g446_n)
  );


  FA
  g_g447_n
  (
    .dout(g447_n),
    .din1(g445_p),
    .din2(g446_p)
  );


  LA
  g_g448_p
  (
    .dout(g448_p),
    .din1(G132_n_spl_),
    .din2(g447_p)
  );


  FA
  g_g449_n
  (
    .dout(g449_n),
    .din1(g444_p),
    .din2(g448_p)
  );


  LA
  g_g450_p
  (
    .dout(g450_p),
    .din1(G132_p_spl_1),
    .din2(g447_n)
  );


  LA
  g_g451_p
  (
    .dout(g451_p),
    .din1(G12_n_spl_100),
    .din2(g271_p_spl_0)
  );


  FA
  g_g451_n
  (
    .dout(g451_n),
    .din1(G12_p_spl_100),
    .din2(g271_n_spl_0)
  );


  LA
  g_g452_p
  (
    .dout(g452_p),
    .din1(G6_n),
    .din2(G12_p_spl_100)
  );


  FA
  g_g452_n
  (
    .dout(g452_n),
    .din1(G6_p),
    .din2(G12_n_spl_100)
  );


  LA
  g_g453_p
  (
    .dout(g453_p),
    .din1(g451_n),
    .din2(g452_n)
  );


  FA
  g_g453_n
  (
    .dout(g453_n),
    .din1(g451_p),
    .din2(g452_p)
  );


  LA
  g_g454_p
  (
    .dout(g454_p),
    .din1(G133_n_spl_),
    .din2(g453_p)
  );


  FA
  g_g455_n
  (
    .dout(g455_n),
    .din1(g450_p),
    .din2(g454_p)
  );


  LA
  g_g456_p
  (
    .dout(g456_p),
    .din1(G12_n_spl_101),
    .din2(g240_p_spl_0)
  );


  FA
  g_g456_n
  (
    .dout(g456_n),
    .din1(G12_p_spl_101),
    .din2(g240_n_spl_00)
  );


  LA
  g_g457_p
  (
    .dout(g457_p),
    .din1(G12_p_spl_101),
    .din2(G13_n)
  );


  FA
  g_g457_n
  (
    .dout(g457_n),
    .din1(G12_n_spl_101),
    .din2(G13_p)
  );


  LA
  g_g458_p
  (
    .dout(g458_p),
    .din1(g456_n),
    .din2(g457_n)
  );


  FA
  g_g458_n
  (
    .dout(g458_n),
    .din1(g456_p),
    .din2(g457_p)
  );


  LA
  g_g459_p
  (
    .dout(g459_p),
    .din1(G125_p_spl_1),
    .din2(g458_n)
  );


  FA
  g_g460_n
  (
    .dout(g460_n),
    .din1(g455_n),
    .din2(g459_p)
  );


  FA
  g_g461_n
  (
    .dout(g461_n),
    .din1(g449_n),
    .din2(g460_n)
  );


  FA
  g_g462_n
  (
    .dout(g462_n),
    .din1(g443_n),
    .din2(g461_n)
  );


  FA
  g_g463_n
  (
    .dout(g463_n),
    .din1(g437_n),
    .din2(g462_n)
  );


  LA
  g_g464_p
  (
    .dout(g464_p),
    .din1(G12_n_spl_110),
    .din2(g290_p_spl_01)
  );


  FA
  g_g464_n
  (
    .dout(g464_n),
    .din1(G12_p_spl_110),
    .din2(g290_n_spl_01)
  );


  LA
  g_g465_p
  (
    .dout(g465_p),
    .din1(G4_n),
    .din2(G12_p_spl_110)
  );


  FA
  g_g465_n
  (
    .dout(g465_n),
    .din1(G4_p),
    .din2(G12_n_spl_110)
  );


  LA
  g_g466_p
  (
    .dout(g466_p),
    .din1(g464_n),
    .din2(g465_n)
  );


  FA
  g_g466_n
  (
    .dout(g466_n),
    .din1(g464_p),
    .din2(g465_p)
  );


  LA
  g_g467_p
  (
    .dout(g467_p),
    .din1(G126_n_spl_),
    .din2(g466_p)
  );


  LA
  g_g468_p
  (
    .dout(g468_p),
    .din1(G133_p_spl_1),
    .din2(g453_n)
  );


  FA
  g_g469_n
  (
    .dout(g469_n),
    .din1(g467_p),
    .din2(g468_p)
  );


  LA
  g_g470_p
  (
    .dout(g470_p),
    .din1(G12_n_spl_111),
    .din2(g280_p_spl_0)
  );


  FA
  g_g470_n
  (
    .dout(g470_n),
    .din1(G12_p_spl_111),
    .din2(g280_n_spl_00)
  );


  LA
  g_g471_p
  (
    .dout(g471_p),
    .din1(G12_p_spl_111),
    .din2(G18_n)
  );


  FA
  g_g471_n
  (
    .dout(g471_n),
    .din1(G12_n_spl_111),
    .din2(G18_p)
  );


  LA
  g_g472_p
  (
    .dout(g472_p),
    .din1(g470_n),
    .din2(g471_n)
  );


  FA
  g_g472_n
  (
    .dout(g472_n),
    .din1(g470_p),
    .din2(g471_p)
  );


  LA
  g_g473_p
  (
    .dout(g473_p),
    .din1(G134_p_spl_1),
    .din2(g472_n)
  );


  LA
  g_g474_p
  (
    .dout(g474_p),
    .din1(G125_n_spl_),
    .din2(g458_p)
  );


  FA
  g_g475_n
  (
    .dout(g475_n),
    .din1(g473_p),
    .din2(g474_p)
  );


  LA
  g_g476_p
  (
    .dout(g476_p),
    .din1(G75_n),
    .din2(G145_n_spl_1000)
  );


  FA
  g_g476_n
  (
    .dout(g476_n),
    .din1(G75_p),
    .din2(G145_p_spl_1000)
  );


  LA
  g_g477_p
  (
    .dout(g477_p),
    .din1(G105_n),
    .din2(G145_p_spl_1000)
  );


  FA
  g_g477_n
  (
    .dout(g477_n),
    .din1(G105_p),
    .din2(G145_n_spl_1000)
  );


  LA
  g_g478_p
  (
    .dout(g478_p),
    .din1(g476_n),
    .din2(g477_n)
  );


  FA
  g_g478_n
  (
    .dout(g478_n),
    .din1(g476_p),
    .din2(g477_p)
  );


  LA
  g_g479_p
  (
    .dout(g479_p),
    .din1(G146_p_spl_100),
    .din2(g478_n)
  );


  FA
  g_g479_n
  (
    .dout(g479_n),
    .din1(G146_n_spl_100),
    .din2(g478_p)
  );


  LA
  g_g480_p
  (
    .dout(g480_p),
    .din1(G95_n),
    .din2(G145_p_spl_1001)
  );


  FA
  g_g480_n
  (
    .dout(g480_n),
    .din1(G95_p),
    .din2(G145_n_spl_1001)
  );


  LA
  g_g481_p
  (
    .dout(g481_p),
    .din1(G85_n),
    .din2(G145_n_spl_1001)
  );


  FA
  g_g481_n
  (
    .dout(g481_n),
    .din1(G85_p),
    .din2(G145_p_spl_1001)
  );


  LA
  g_g482_p
  (
    .dout(g482_p),
    .din1(g480_n),
    .din2(g481_n)
  );


  FA
  g_g482_n
  (
    .dout(g482_n),
    .din1(g480_p),
    .din2(g481_p)
  );


  LA
  g_g483_p
  (
    .dout(g483_p),
    .din1(G146_n_spl_100),
    .din2(g482_n)
  );


  FA
  g_g483_n
  (
    .dout(g483_n),
    .din1(G146_p_spl_100),
    .din2(g482_p)
  );


  LA
  g_g484_p
  (
    .dout(g484_p),
    .din1(g479_n),
    .din2(g483_n)
  );


  FA
  g_g484_n
  (
    .dout(g484_n),
    .din1(g479_p),
    .din2(g483_p)
  );


  LA
  g_g485_p
  (
    .dout(g485_p),
    .din1(G23_n_spl_011),
    .din2(g484_n_spl_0)
  );


  FA
  g_g485_n
  (
    .dout(g485_n),
    .din1(G23_p_spl_011),
    .din2(g484_p_spl_0)
  );


  LA
  g_g486_p
  (
    .dout(g486_p),
    .din1(G19_n),
    .din2(G23_p_spl_100)
  );


  FA
  g_g486_n
  (
    .dout(g486_n),
    .din1(G19_p),
    .din2(G23_n_spl_100)
  );


  LA
  g_g487_p
  (
    .dout(g487_p),
    .din1(g485_n),
    .din2(g486_n)
  );


  FA
  g_g487_n
  (
    .dout(g487_n),
    .din1(g485_p),
    .din2(g486_p)
  );


  LA
  g_g488_p
  (
    .dout(g488_p),
    .din1(G135_n_spl_1),
    .din2(g487_p)
  );


  LA
  g_g489_p
  (
    .dout(g489_p),
    .din1(G135_p_spl_1),
    .din2(g487_n)
  );


  LA
  g_g490_p
  (
    .dout(g490_p),
    .din1(G134_n_spl_1),
    .din2(g472_p)
  );


  FA
  g_g491_n
  (
    .dout(g491_n),
    .din1(g489_p),
    .din2(g490_p)
  );


  FA
  g_g492_n
  (
    .dout(g492_n),
    .din1(g488_p),
    .din2(g491_n)
  );


  FA
  g_g493_n
  (
    .dout(g493_n),
    .din1(g475_n),
    .din2(g492_n)
  );


  FA
  g_g494_n
  (
    .dout(g494_n),
    .din1(g469_n),
    .din2(g493_n)
  );


  LA
  g_g495_p
  (
    .dout(g495_p),
    .din1(G81_n),
    .din2(G145_n_spl_1010)
  );


  FA
  g_g495_n
  (
    .dout(g495_n),
    .din1(G81_p),
    .din2(G145_p_spl_1010)
  );


  LA
  g_g496_p
  (
    .dout(g496_p),
    .din1(G111_n),
    .din2(G145_p_spl_1010)
  );


  FA
  g_g496_n
  (
    .dout(g496_n),
    .din1(G111_p),
    .din2(G145_n_spl_1010)
  );


  LA
  g_g497_p
  (
    .dout(g497_p),
    .din1(g495_n),
    .din2(g496_n)
  );


  FA
  g_g497_n
  (
    .dout(g497_n),
    .din1(g495_p),
    .din2(g496_p)
  );


  LA
  g_g498_p
  (
    .dout(g498_p),
    .din1(G146_p_spl_101),
    .din2(g497_n)
  );


  FA
  g_g498_n
  (
    .dout(g498_n),
    .din1(G146_n_spl_101),
    .din2(g497_p)
  );


  LA
  g_g499_p
  (
    .dout(g499_p),
    .din1(G101_n),
    .din2(G145_p_spl_1011)
  );


  FA
  g_g499_n
  (
    .dout(g499_n),
    .din1(G101_p),
    .din2(G145_n_spl_1011)
  );


  LA
  g_g500_p
  (
    .dout(g500_p),
    .din1(G91_n),
    .din2(G145_n_spl_1011)
  );


  FA
  g_g500_n
  (
    .dout(g500_n),
    .din1(G91_p),
    .din2(G145_p_spl_1011)
  );


  LA
  g_g501_p
  (
    .dout(g501_p),
    .din1(g499_n),
    .din2(g500_n)
  );


  FA
  g_g501_n
  (
    .dout(g501_n),
    .din1(g499_p),
    .din2(g500_p)
  );


  LA
  g_g502_p
  (
    .dout(g502_p),
    .din1(G146_n_spl_101),
    .din2(g501_n)
  );


  FA
  g_g502_n
  (
    .dout(g502_n),
    .din1(G146_p_spl_101),
    .din2(g501_p)
  );


  LA
  g_g503_p
  (
    .dout(g503_p),
    .din1(g498_n),
    .din2(g502_n)
  );


  FA
  g_g503_n
  (
    .dout(g503_n),
    .din1(g498_p),
    .din2(g502_p)
  );


  LA
  g_g504_p
  (
    .dout(g504_p),
    .din1(G23_n_spl_100),
    .din2(g503_n_spl_0)
  );


  FA
  g_g504_n
  (
    .dout(g504_n),
    .din1(G23_p_spl_100),
    .din2(g503_p_spl_0)
  );


  LA
  g_g505_p
  (
    .dout(g505_p),
    .din1(G23_p_spl_101),
    .din2(G25_n)
  );


  FA
  g_g505_n
  (
    .dout(g505_n),
    .din1(G23_n_spl_101),
    .din2(G25_p)
  );


  LA
  g_g506_p
  (
    .dout(g506_p),
    .din1(g504_n),
    .din2(g505_n)
  );


  FA
  g_g506_n
  (
    .dout(g506_n),
    .din1(g504_p),
    .din2(g505_p)
  );


  LA
  g_g507_p
  (
    .dout(g507_p),
    .din1(G139_p_spl_1),
    .din2(g506_n)
  );


  LA
  g_g508_p
  (
    .dout(g508_p),
    .din1(G23_n_spl_101),
    .din2(g194_n_spl_0)
  );


  FA
  g_g508_n
  (
    .dout(g508_n),
    .din1(G23_p_spl_101),
    .din2(g194_p_spl_0)
  );


  LA
  g_g509_p
  (
    .dout(g509_p),
    .din1(G23_p_spl_110),
    .din2(G27_n)
  );


  FA
  g_g509_n
  (
    .dout(g509_n),
    .din1(G23_n_spl_110),
    .din2(G27_p)
  );


  LA
  g_g510_p
  (
    .dout(g510_p),
    .din1(g508_n),
    .din2(g509_n)
  );


  FA
  g_g510_n
  (
    .dout(g510_n),
    .din1(g508_p),
    .din2(g509_p)
  );


  LA
  g_g511_p
  (
    .dout(g511_p),
    .din1(G142_p_spl_1),
    .din2(g510_n)
  );


  FA
  g_g512_n
  (
    .dout(g512_n),
    .din1(g507_p),
    .din2(g511_p)
  );


  LA
  g_g513_p
  (
    .dout(g513_p),
    .din1(G139_n_spl_),
    .din2(g506_p)
  );


  LA
  g_g514_p
  (
    .dout(g514_p),
    .din1(G82_n),
    .din2(G145_n_spl_1100)
  );


  FA
  g_g514_n
  (
    .dout(g514_n),
    .din1(G82_p),
    .din2(G145_p_spl_1100)
  );


  LA
  g_g515_p
  (
    .dout(g515_p),
    .din1(G112_n),
    .din2(G145_p_spl_1100)
  );


  FA
  g_g515_n
  (
    .dout(g515_n),
    .din1(G112_p),
    .din2(G145_n_spl_1100)
  );


  LA
  g_g516_p
  (
    .dout(g516_p),
    .din1(g514_n),
    .din2(g515_n)
  );


  FA
  g_g516_n
  (
    .dout(g516_n),
    .din1(g514_p),
    .din2(g515_p)
  );


  LA
  g_g517_p
  (
    .dout(g517_p),
    .din1(G146_p_spl_110),
    .din2(g516_n)
  );


  FA
  g_g517_n
  (
    .dout(g517_n),
    .din1(G146_n_spl_110),
    .din2(g516_p)
  );


  LA
  g_g518_p
  (
    .dout(g518_p),
    .din1(G102_n),
    .din2(G145_p_spl_1101)
  );


  FA
  g_g518_n
  (
    .dout(g518_n),
    .din1(G102_p),
    .din2(G145_n_spl_1101)
  );


  LA
  g_g519_p
  (
    .dout(g519_p),
    .din1(G92_n),
    .din2(G145_n_spl_1101)
  );


  FA
  g_g519_n
  (
    .dout(g519_n),
    .din1(G92_p),
    .din2(G145_p_spl_1101)
  );


  LA
  g_g520_p
  (
    .dout(g520_p),
    .din1(g518_n),
    .din2(g519_n)
  );


  FA
  g_g520_n
  (
    .dout(g520_n),
    .din1(g518_p),
    .din2(g519_p)
  );


  LA
  g_g521_p
  (
    .dout(g521_p),
    .din1(G146_n_spl_110),
    .din2(g520_n)
  );


  FA
  g_g521_n
  (
    .dout(g521_n),
    .din1(G146_p_spl_110),
    .din2(g520_p)
  );


  LA
  g_g522_p
  (
    .dout(g522_p),
    .din1(g517_n),
    .din2(g521_n)
  );


  FA
  g_g522_n
  (
    .dout(g522_n),
    .din1(g517_p),
    .din2(g521_p)
  );


  LA
  g_g523_p
  (
    .dout(g523_p),
    .din1(G23_n_spl_110),
    .din2(g522_n_spl_0)
  );


  FA
  g_g523_n
  (
    .dout(g523_n),
    .din1(G23_p_spl_110),
    .din2(g522_p_spl_0)
  );


  LA
  g_g524_p
  (
    .dout(g524_p),
    .din1(G20_n),
    .din2(G23_p_spl_11)
  );


  FA
  g_g524_n
  (
    .dout(g524_n),
    .din1(G20_p),
    .din2(G23_n_spl_11)
  );


  LA
  g_g525_p
  (
    .dout(g525_p),
    .din1(g523_n),
    .din2(g524_n)
  );


  FA
  g_g525_n
  (
    .dout(g525_n),
    .din1(g523_p),
    .din2(g524_p)
  );


  LA
  g_g526_p
  (
    .dout(g526_p),
    .din1(G138_p_spl_0),
    .din2(g525_n)
  );


  LA
  g_g527_p
  (
    .dout(g527_p),
    .din1(G138_n_spl_1),
    .din2(g525_p)
  );


  FA
  g_g528_n
  (
    .dout(g528_n),
    .din1(g526_p),
    .din2(g527_p)
  );


  FA
  g_g529_n
  (
    .dout(g529_n),
    .din1(g513_p),
    .din2(g528_n)
  );


  FA
  g_g530_n
  (
    .dout(g530_n),
    .din1(g512_n),
    .din2(g529_n)
  );


  LA
  g_g531_p
  (
    .dout(g531_p),
    .din1(G129_p_spl_1),
    .din2(g395_n)
  );


  LA
  g_g532_p
  (
    .dout(g532_p),
    .din1(G142_n_spl_),
    .din2(g510_p)
  );


  FA
  g_g533_n
  (
    .dout(g533_n),
    .din1(g531_p),
    .din2(g532_p)
  );


  LA
  g_g534_p
  (
    .dout(g534_p),
    .din1(G126_p_spl_1),
    .din2(g466_n)
  );


  LA
  g_g535_p
  (
    .dout(g535_p),
    .din1(G128_n_spl_),
    .din2(g440_p)
  );


  FA
  g_g536_n
  (
    .dout(g536_n),
    .din1(g534_p),
    .din2(g535_p)
  );


  FA
  g_g537_n
  (
    .dout(g537_n),
    .din1(g533_n),
    .din2(g536_n)
  );


  FA
  g_g538_n
  (
    .dout(g538_n),
    .din1(g530_n),
    .din2(g537_n)
  );


  FA
  g_g539_n
  (
    .dout(g539_n),
    .din1(g494_n),
    .din2(g538_n)
  );


  FA
  g_g540_n
  (
    .dout(g540_n),
    .din1(g463_n),
    .din2(g539_n)
  );


  LA
  g_g541_p
  (
    .dout(g541_p),
    .din1(G118_p_spl_),
    .din2(g290_p_spl_01)
  );


  FA
  g_g541_n
  (
    .dout(g541_n),
    .din1(G118_n_spl_),
    .din2(g290_n_spl_01)
  );


  LA
  g_g542_p
  (
    .dout(g542_p),
    .din1(G51_p),
    .din2(g204_p_spl_11)
  );


  FA
  g_g542_n
  (
    .dout(g542_n),
    .din1(G51_n),
    .din2(g204_n_spl_11)
  );


  LA
  g_g543_p
  (
    .dout(g543_p),
    .din1(G62_p),
    .din2(G117_n_spl_1110)
  );


  FA
  g_g543_n
  (
    .dout(g543_n),
    .din1(G62_n),
    .din2(G117_p_spl_1110)
  );


  LA
  g_g544_p
  (
    .dout(g544_p),
    .din1(G120_n_spl_111),
    .din2(g543_n)
  );


  FA
  g_g544_n
  (
    .dout(g544_n),
    .din1(G120_p_spl_111),
    .din2(g543_p)
  );


  LA
  g_g545_p
  (
    .dout(g545_p),
    .din1(G41_n),
    .din2(G117_n_spl_1110)
  );


  FA
  g_g545_n
  (
    .dout(g545_n),
    .din1(G41_p),
    .din2(G117_p_spl_1110)
  );


  LA
  g_g546_p
  (
    .dout(g546_p),
    .din1(G120_p_spl_111),
    .din2(g545_p)
  );


  FA
  g_g546_n
  (
    .dout(g546_n),
    .din1(G120_n_spl_111),
    .din2(g545_n)
  );


  LA
  g_g547_p
  (
    .dout(g547_p),
    .din1(G73_n),
    .din2(G117_p_spl_111)
  );


  FA
  g_g547_n
  (
    .dout(g547_n),
    .din1(G73_p),
    .din2(G117_n_spl_111)
  );


  LA
  g_g548_p
  (
    .dout(g548_p),
    .din1(g546_n),
    .din2(g547_n)
  );


  FA
  g_g548_n
  (
    .dout(g548_n),
    .din1(g546_p),
    .din2(g547_p)
  );


  LA
  g_g549_p
  (
    .dout(g549_p),
    .din1(g544_n),
    .din2(g548_p)
  );


  FA
  g_g549_n
  (
    .dout(g549_n),
    .din1(g544_p),
    .din2(g548_n)
  );


  LA
  g_g550_p
  (
    .dout(g550_p),
    .din1(g542_n),
    .din2(g549_n)
  );


  FA
  g_g550_n
  (
    .dout(g550_n),
    .din1(g542_p),
    .din2(g549_p)
  );


  LA
  g_g551_p
  (
    .dout(g551_p),
    .din1(g240_n_spl_0),
    .din2(g550_n_spl_0)
  );


  FA
  g_g551_n
  (
    .dout(g551_n),
    .din1(g240_p_spl_1),
    .din2(g550_p_spl_)
  );


  LA
  g_g552_p
  (
    .dout(g552_p),
    .din1(g240_p_spl_1),
    .din2(g550_p_spl_)
  );


  FA
  g_g552_n
  (
    .dout(g552_n),
    .din1(g240_n_spl_1),
    .din2(g550_n_spl_0)
  );


  LA
  g_g553_p
  (
    .dout(g553_p),
    .din1(g551_n),
    .din2(g552_n)
  );


  FA
  g_g553_n
  (
    .dout(g553_n),
    .din1(g551_p),
    .din2(g552_p)
  );


  LA
  g_g554_p
  (
    .dout(g554_p),
    .din1(g541_p),
    .din2(g553_n_spl_0)
  );


  LA
  g_g555_p
  (
    .dout(g555_p),
    .din1(g541_n),
    .din2(g553_p_spl_0)
  );


  FA
  g_g556_n
  (
    .dout(g556_n),
    .din1(g554_p),
    .din2(g555_p)
  );


  LA
  g_g557_p
  (
    .dout(g557_p),
    .din1(G122_n_spl_),
    .din2(g556_n)
  );


  LA
  g_g558_p
  (
    .dout(g558_p),
    .din1(G122_p),
    .din2(g550_n_spl_1)
  );


  FA
  g_g559_n
  (
    .dout(g559_n),
    .din1(g557_p),
    .din2(g558_p)
  );


  LA
  g_g560_p
  (
    .dout(g560_p),
    .din1(g185_n_spl_00),
    .din2(g194_n_spl_0)
  );


  FA
  g_g560_n
  (
    .dout(g560_n),
    .din1(g185_p_spl_0),
    .din2(g194_p_spl_0)
  );


  LA
  g_g561_p
  (
    .dout(g561_p),
    .din1(g185_p_spl_1),
    .din2(g194_p_spl_)
  );


  FA
  g_g561_n
  (
    .dout(g561_n),
    .din1(g185_n_spl_0),
    .din2(g194_n_spl_1)
  );


  LA
  g_g562_p
  (
    .dout(g562_p),
    .din1(g560_n),
    .din2(g561_n)
  );


  FA
  g_g562_n
  (
    .dout(g562_n),
    .din1(g560_p),
    .din2(g561_p)
  );


  LA
  g_g563_p
  (
    .dout(g563_p),
    .din1(g310_p_spl_0),
    .din2(g562_p_spl_)
  );


  FA
  g_g563_n
  (
    .dout(g563_n),
    .din1(g310_n_spl_1),
    .din2(g562_n_spl_)
  );


  LA
  g_g564_p
  (
    .dout(g564_p),
    .din1(g310_n_spl_1),
    .din2(g562_n_spl_)
  );


  FA
  g_g564_n
  (
    .dout(g564_n),
    .din1(g310_p_spl_),
    .din2(g562_p_spl_)
  );


  LA
  g_g565_p
  (
    .dout(g565_p),
    .din1(g563_n),
    .din2(g564_n)
  );


  FA
  g_g565_n
  (
    .dout(g565_n),
    .din1(g563_p),
    .din2(g564_p)
  );


  LA
  g_g566_p
  (
    .dout(g566_p),
    .din1(G84_n),
    .din2(G145_n_spl_1110)
  );


  FA
  g_g566_n
  (
    .dout(g566_n),
    .din1(G84_p),
    .din2(G145_p_spl_1110)
  );


  LA
  g_g567_p
  (
    .dout(g567_p),
    .din1(G114_n),
    .din2(G145_p_spl_1110)
  );


  FA
  g_g567_n
  (
    .dout(g567_n),
    .din1(G114_p),
    .din2(G145_n_spl_1110)
  );


  LA
  g_g568_p
  (
    .dout(g568_p),
    .din1(g566_n),
    .din2(g567_n)
  );


  FA
  g_g568_n
  (
    .dout(g568_n),
    .din1(g566_p),
    .din2(g567_p)
  );


  LA
  g_g569_p
  (
    .dout(g569_p),
    .din1(G146_p_spl_111),
    .din2(g568_n)
  );


  FA
  g_g569_n
  (
    .dout(g569_n),
    .din1(G146_n_spl_111),
    .din2(g568_p)
  );


  LA
  g_g570_p
  (
    .dout(g570_p),
    .din1(G104_n),
    .din2(G145_p_spl_1111)
  );


  FA
  g_g570_n
  (
    .dout(g570_n),
    .din1(G104_p),
    .din2(G145_n_spl_1111)
  );


  LA
  g_g571_p
  (
    .dout(g571_p),
    .din1(G94_n),
    .din2(G145_n_spl_1111)
  );


  FA
  g_g571_n
  (
    .dout(g571_n),
    .din1(G94_p),
    .din2(G145_p_spl_1111)
  );


  LA
  g_g572_p
  (
    .dout(g572_p),
    .din1(g570_n),
    .din2(g571_n)
  );


  FA
  g_g572_n
  (
    .dout(g572_n),
    .din1(g570_p),
    .din2(g571_p)
  );


  LA
  g_g573_p
  (
    .dout(g573_p),
    .din1(G146_n_spl_111),
    .din2(g572_n)
  );


  FA
  g_g573_n
  (
    .dout(g573_n),
    .din1(G146_p_spl_111),
    .din2(g572_p)
  );


  LA
  g_g574_p
  (
    .dout(g574_p),
    .din1(g569_n),
    .din2(g573_n)
  );


  FA
  g_g574_n
  (
    .dout(g574_n),
    .din1(g569_p),
    .din2(g573_p)
  );


  LA
  g_g575_p
  (
    .dout(g575_p),
    .din1(g484_p_spl_0),
    .din2(g574_p_spl_)
  );


  FA
  g_g575_n
  (
    .dout(g575_n),
    .din1(g484_n_spl_0),
    .din2(g574_n_spl_)
  );


  LA
  g_g576_p
  (
    .dout(g576_p),
    .din1(g484_n_spl_1),
    .din2(g574_n_spl_)
  );


  FA
  g_g576_n
  (
    .dout(g576_n),
    .din1(g484_p_spl_1),
    .din2(g574_p_spl_)
  );


  LA
  g_g577_p
  (
    .dout(g577_p),
    .din1(g575_n),
    .din2(g576_n)
  );


  FA
  g_g577_n
  (
    .dout(g577_n),
    .din1(g575_p),
    .din2(g576_p)
  );


  LA
  g_g578_p
  (
    .dout(g578_p),
    .din1(g203_n_spl_00),
    .din2(g503_n_spl_0)
  );


  FA
  g_g578_n
  (
    .dout(g578_n),
    .din1(g203_p_spl_0),
    .din2(g503_p_spl_0)
  );


  LA
  g_g579_p
  (
    .dout(g579_p),
    .din1(g203_p_spl_1),
    .din2(g503_p_spl_)
  );


  FA
  g_g579_n
  (
    .dout(g579_n),
    .din1(g203_n_spl_0),
    .din2(g503_n_spl_)
  );


  LA
  g_g580_p
  (
    .dout(g580_p),
    .din1(g578_n),
    .din2(g579_n)
  );


  FA
  g_g580_n
  (
    .dout(g580_n),
    .din1(g578_p),
    .din2(g579_p)
  );


  LA
  g_g581_p
  (
    .dout(g581_p),
    .din1(g577_p_spl_),
    .din2(g580_n_spl_)
  );


  FA
  g_g581_n
  (
    .dout(g581_n),
    .din1(g577_n_spl_),
    .din2(g580_p_spl_)
  );


  LA
  g_g582_p
  (
    .dout(g582_p),
    .din1(g577_n_spl_),
    .din2(g580_p_spl_)
  );


  FA
  g_g582_n
  (
    .dout(g582_n),
    .din1(g577_p_spl_),
    .din2(g580_n_spl_)
  );


  LA
  g_g583_p
  (
    .dout(g583_p),
    .din1(g581_n),
    .din2(g582_n)
  );


  FA
  g_g583_n
  (
    .dout(g583_n),
    .din1(g581_p),
    .din2(g582_p)
  );


  LA
  g_g584_p
  (
    .dout(g584_p),
    .din1(g427_n_spl_0),
    .din2(g522_n_spl_0)
  );


  FA
  g_g584_n
  (
    .dout(g584_n),
    .din1(g427_p_spl_0),
    .din2(g522_p_spl_0)
  );


  LA
  g_g585_p
  (
    .dout(g585_p),
    .din1(g427_p_spl_1),
    .din2(g522_p_spl_1)
  );


  FA
  g_g585_n
  (
    .dout(g585_n),
    .din1(g427_n_spl_1),
    .din2(g522_n_spl_1)
  );


  LA
  g_g586_p
  (
    .dout(g586_p),
    .din1(g584_n),
    .din2(g585_n)
  );


  FA
  g_g586_n
  (
    .dout(g586_n),
    .din1(g584_p),
    .din2(g585_p)
  );


  LA
  g_g587_p
  (
    .dout(g587_p),
    .din1(g583_n_spl_),
    .din2(g586_n_spl_)
  );


  FA
  g_g587_n
  (
    .dout(g587_n),
    .din1(g583_p_spl_),
    .din2(g586_p_spl_)
  );


  LA
  g_g588_p
  (
    .dout(g588_p),
    .din1(g583_p_spl_),
    .din2(g586_p_spl_)
  );


  FA
  g_g588_n
  (
    .dout(g588_n),
    .din1(g583_n_spl_),
    .din2(g586_n_spl_)
  );


  LA
  g_g589_p
  (
    .dout(g589_p),
    .din1(g587_n),
    .din2(g588_n)
  );


  FA
  g_g589_n
  (
    .dout(g589_n),
    .din1(g587_p),
    .din2(g588_p)
  );


  FA
  g_g590_n
  (
    .dout(g590_n),
    .din1(g565_n),
    .din2(g589_p)
  );


  FA
  g_g591_n
  (
    .dout(g591_n),
    .din1(g565_p),
    .din2(g589_n)
  );


  LA
  g_g592_p
  (
    .dout(g592_p),
    .din1(G29_n_spl_),
    .din2(g591_n)
  );


  LA
  g_g593_p
  (
    .dout(g593_p),
    .din1(g590_n),
    .din2(g592_p)
  );


  FA
  g_g594_n
  (
    .dout(g594_n),
    .din1(G123_p_spl_1),
    .din2(g550_n_spl_1)
  );


  LA
  g_g595_p
  (
    .dout(g595_p),
    .din1(g213_p_spl_00),
    .din2(g262_n_spl_0)
  );


  FA
  g_g595_n
  (
    .dout(g595_n),
    .din1(g213_n_spl_0),
    .din2(g262_p_spl_0)
  );


  LA
  g_g596_p
  (
    .dout(g596_p),
    .din1(g213_n_spl_1),
    .din2(g262_p_spl_1)
  );


  FA
  g_g596_n
  (
    .dout(g596_n),
    .din1(g213_p_spl_0),
    .din2(g262_n_spl_1)
  );


  LA
  g_g597_p
  (
    .dout(g597_p),
    .din1(g595_n),
    .din2(g596_n)
  );


  FA
  g_g597_n
  (
    .dout(g597_n),
    .din1(g595_p),
    .din2(g596_p)
  );


  LA
  g_g598_p
  (
    .dout(g598_p),
    .din1(g271_n_spl_0),
    .din2(g280_n_spl_00)
  );


  FA
  g_g598_n
  (
    .dout(g598_n),
    .din1(g271_p_spl_0),
    .din2(g280_p_spl_0)
  );


  LA
  g_g599_p
  (
    .dout(g599_p),
    .din1(g271_p_spl_1),
    .din2(g280_p_spl_1)
  );


  FA
  g_g599_n
  (
    .dout(g599_n),
    .din1(g271_n_spl_1),
    .din2(g280_n_spl_0)
  );


  LA
  g_g600_p
  (
    .dout(g600_p),
    .din1(g598_n),
    .din2(g599_n)
  );


  FA
  g_g600_n
  (
    .dout(g600_n),
    .din1(g598_p),
    .din2(g599_p)
  );


  LA
  g_g601_p
  (
    .dout(g601_p),
    .din1(g597_p_spl_),
    .din2(g600_n_spl_)
  );


  FA
  g_g601_n
  (
    .dout(g601_n),
    .din1(g597_n_spl_),
    .din2(g600_p_spl_)
  );


  LA
  g_g602_p
  (
    .dout(g602_p),
    .din1(g597_n_spl_),
    .din2(g600_p_spl_)
  );


  FA
  g_g602_n
  (
    .dout(g602_n),
    .din1(g597_p_spl_),
    .din2(g600_n_spl_)
  );


  LA
  g_g603_p
  (
    .dout(g603_p),
    .din1(g601_n),
    .din2(g602_n)
  );


  FA
  g_g603_n
  (
    .dout(g603_n),
    .din1(g601_p),
    .din2(g602_p)
  );


  LA
  g_g604_p
  (
    .dout(g604_p),
    .din1(g255_p_spl_00),
    .din2(g290_n_spl_10)
  );


  FA
  g_g604_n
  (
    .dout(g604_n),
    .din1(g255_n_spl_0),
    .din2(g290_p_spl_1)
  );


  LA
  g_g605_p
  (
    .dout(g605_p),
    .din1(g255_n_spl_1),
    .din2(g290_p_spl_1)
  );


  FA
  g_g605_n
  (
    .dout(g605_n),
    .din1(g255_p_spl_0),
    .din2(g290_n_spl_10)
  );


  LA
  g_g606_p
  (
    .dout(g606_p),
    .din1(g604_n),
    .din2(g605_n)
  );


  FA
  g_g606_n
  (
    .dout(g606_n),
    .din1(g604_p),
    .din2(g605_p)
  );


  LA
  g_g607_p
  (
    .dout(g607_p),
    .din1(g553_p_spl_0),
    .din2(g606_n_spl_)
  );


  FA
  g_g607_n
  (
    .dout(g607_n),
    .din1(g553_n_spl_0),
    .din2(g606_p_spl_)
  );


  LA
  g_g608_p
  (
    .dout(g608_p),
    .din1(g553_n_spl_),
    .din2(g606_p_spl_)
  );


  FA
  g_g608_n
  (
    .dout(g608_n),
    .din1(g553_p_spl_),
    .din2(g606_n_spl_)
  );


  LA
  g_g609_p
  (
    .dout(g609_p),
    .din1(g607_n),
    .din2(g608_n)
  );


  FA
  g_g609_n
  (
    .dout(g609_n),
    .din1(g607_p),
    .din2(g608_p)
  );


  LA
  g_g610_p
  (
    .dout(g610_p),
    .din1(g298_p_spl_0),
    .din2(g609_n_spl_0)
  );


  FA
  g_g610_n
  (
    .dout(g610_n),
    .din1(g298_n_spl_),
    .din2(g609_p_spl_0)
  );


  LA
  g_g611_p
  (
    .dout(g611_p),
    .din1(g298_n_spl_),
    .din2(g609_p_spl_0)
  );


  FA
  g_g611_n
  (
    .dout(g611_n),
    .din1(g298_p_spl_),
    .din2(g609_n_spl_0)
  );


  LA
  g_g612_p
  (
    .dout(g612_p),
    .din1(g610_n),
    .din2(g611_n)
  );


  FA
  g_g612_n
  (
    .dout(g612_n),
    .din1(g610_p),
    .din2(g611_p)
  );


  FA
  g_g613_n
  (
    .dout(g613_n),
    .din1(g603_p_spl_),
    .din2(g612_n)
  );


  FA
  g_g614_n
  (
    .dout(g614_n),
    .din1(g603_n_spl_),
    .din2(g612_p)
  );


  LA
  g_g615_p
  (
    .dout(g615_p),
    .din1(g613_n),
    .din2(g614_n)
  );


  FA
  g_g616_n
  (
    .dout(g616_n),
    .din1(G123_n_spl_1),
    .din2(g615_p)
  );


  LA
  g_g617_p
  (
    .dout(g617_p),
    .din1(g594_n),
    .din2(g616_n)
  );


  LA
  g_g618_p
  (
    .dout(g618_p),
    .din1(g222_p_spl_01),
    .din2(g231_n_spl_0)
  );


  FA
  g_g618_n
  (
    .dout(g618_n),
    .din1(g222_n_spl_0),
    .din2(g231_p_spl_00)
  );


  LA
  g_g619_p
  (
    .dout(g619_p),
    .din1(g222_n_spl_1),
    .din2(g231_p_spl_01)
  );


  FA
  g_g619_n
  (
    .dout(g619_n),
    .din1(g222_p_spl_01),
    .din2(g231_n_spl_1)
  );


  LA
  g_g620_p
  (
    .dout(g620_p),
    .din1(g618_n),
    .din2(g619_n)
  );


  FA
  g_g620_n
  (
    .dout(g620_n),
    .din1(g618_p),
    .din2(g619_p)
  );


  LA
  g_g621_p
  (
    .dout(g621_p),
    .din1(g609_n_spl_1),
    .din2(g620_p_spl_)
  );


  FA
  g_g621_n
  (
    .dout(g621_n),
    .din1(g609_p_spl_1),
    .din2(g620_n_spl_)
  );


  LA
  g_g622_p
  (
    .dout(g622_p),
    .din1(g609_p_spl_1),
    .din2(g620_n_spl_)
  );


  FA
  g_g622_n
  (
    .dout(g622_n),
    .din1(g609_n_spl_1),
    .din2(g620_p_spl_)
  );


  LA
  g_g623_p
  (
    .dout(g623_p),
    .din1(g621_n),
    .din2(g622_n)
  );


  FA
  g_g623_n
  (
    .dout(g623_n),
    .din1(g621_p),
    .din2(g622_p)
  );


  FA
  g_g624_n
  (
    .dout(g624_n),
    .din1(g603_n_spl_),
    .din2(g623_p)
  );


  FA
  g_g625_n
  (
    .dout(g625_n),
    .din1(g603_p_spl_),
    .din2(g623_n)
  );


  LA
  g_g626_p
  (
    .dout(g626_p),
    .din1(G29_n_spl_),
    .din2(g625_n)
  );


  LA
  g_g627_p
  (
    .dout(g627_p),
    .din1(g624_n),
    .din2(g626_p)
  );


  LA
  g_g628_p
  (
    .dout(g628_p),
    .din1(G127_n),
    .din2(g203_p_spl_1)
  );


  FA
  g_g628_n
  (
    .dout(g628_n),
    .din1(G127_p),
    .din2(g203_n_spl_1)
  );


  LA
  g_g629_p
  (
    .dout(g629_p),
    .din1(G30_p),
    .din2(g185_n_spl_1)
  );


  FA
  g_g629_n
  (
    .dout(g629_n),
    .din1(G30_n),
    .din2(g185_p_spl_1)
  );


  LA
  g_g630_p
  (
    .dout(g630_p),
    .din1(g628_p_spl_),
    .din2(g629_p_spl_)
  );


  FA
  g_g630_n
  (
    .dout(g630_n),
    .din1(g628_n_spl_),
    .din2(g629_n_spl_)
  );


  FA
  g_g631_n
  (
    .dout(g631_n),
    .din1(G8_n_spl_),
    .din2(g630_p_spl_00)
  );


  FA
  g_g632_n
  (
    .dout(g632_n),
    .din1(G133_p_spl_1),
    .din2(g631_n_spl_0)
  );


  LA
  g_g633_p
  (
    .dout(g633_p),
    .din1(G8_p_spl_0),
    .din2(g630_p_spl_00)
  );


  FA
  g_g633_n
  (
    .dout(g633_n),
    .din1(G8_n_spl_),
    .din2(g630_n_spl_00)
  );


  LA
  g_g634_p
  (
    .dout(g634_p),
    .din1(g271_p_spl_1),
    .din2(g633_p_spl_)
  );


  FA
  g_g635_n
  (
    .dout(g635_n),
    .din1(G132_p_spl_1),
    .din2(g631_n_spl_0)
  );


  LA
  g_g636_p
  (
    .dout(g636_p),
    .din1(g262_n_spl_1),
    .din2(g633_p_spl_)
  );


  LA
  g_g637_p
  (
    .dout(g637_p),
    .din1(G8_p_spl_0),
    .din2(g213_p_spl_1)
  );


  FA
  g_g638_n
  (
    .dout(g638_n),
    .din1(G131_p_spl_1),
    .din2(g631_n_spl_1)
  );


  FA
  g_g639_n
  (
    .dout(g639_n),
    .din1(G142_p_spl_1),
    .din2(g633_n_spl_)
  );


  LA
  g_g640_p
  (
    .dout(g640_p),
    .din1(g638_n),
    .din2(g639_n)
  );


  FA
  g_g641_n
  (
    .dout(g641_n),
    .din1(g637_p_spl_),
    .din2(g640_p_spl_)
  );


  LA
  g_g642_p
  (
    .dout(g642_p),
    .din1(g637_p_spl_),
    .din2(g640_p_spl_)
  );


  LA
  g_g643_p
  (
    .dout(g643_p),
    .din1(G8_p_spl_),
    .din2(g222_p_spl_1)
  );


  FA
  g_g644_n
  (
    .dout(g644_n),
    .din1(G130_p_spl_1),
    .din2(g631_n_spl_1)
  );


  FA
  g_g645_n
  (
    .dout(g645_n),
    .din1(G141_p_spl_1),
    .din2(g633_n_spl_)
  );


  LA
  g_g646_p
  (
    .dout(g646_p),
    .din1(g644_n),
    .din2(g645_n)
  );


  FA
  g_g647_n
  (
    .dout(g647_n),
    .din1(g643_p_spl_),
    .din2(g646_p_spl_)
  );


  LA
  g_g648_p
  (
    .dout(g648_p),
    .din1(g643_p_spl_),
    .din2(g646_p_spl_)
  );


  LA
  g_g649_p
  (
    .dout(g649_p),
    .din1(G129_p_spl_1),
    .din2(g630_n_spl_00)
  );


  LA
  g_g650_p
  (
    .dout(g650_p),
    .din1(G140_p_spl_1),
    .din2(g630_p_spl_01)
  );


  FA
  g_g651_n
  (
    .dout(g651_n),
    .din1(g649_p),
    .din2(g650_p)
  );


  FA
  g_g652_n
  (
    .dout(g652_n),
    .din1(g231_p_spl_01),
    .din2(g651_n_spl_)
  );


  LA
  g_g653_p
  (
    .dout(g653_p),
    .din1(g231_p_spl_1),
    .din2(g651_n_spl_)
  );


  LA
  g_g654_p
  (
    .dout(g654_p),
    .din1(G128_p_spl_1),
    .din2(g630_n_spl_0)
  );


  LA
  g_g655_p
  (
    .dout(g655_p),
    .din1(G139_p_spl_1),
    .din2(g630_p_spl_01)
  );


  FA
  g_g656_n
  (
    .dout(g656_n),
    .din1(g654_p),
    .din2(g655_p)
  );


  LA
  g_g657_p
  (
    .dout(g657_p),
    .din1(g255_p_spl_1),
    .din2(g656_n_spl_)
  );


  FA
  g_g658_n
  (
    .dout(g658_n),
    .din1(g653_p),
    .din2(g657_p)
  );


  LA
  g_g659_p
  (
    .dout(g659_p),
    .din1(G126_p_spl_1),
    .din2(g630_n_spl_1)
  );


  LA
  g_g660_p
  (
    .dout(g660_p),
    .din1(G138_p_spl_1),
    .din2(g630_p_spl_1)
  );


  FA
  g_g661_n
  (
    .dout(g661_n),
    .din1(g659_p),
    .din2(g660_p)
  );


  LA
  g_g662_p
  (
    .dout(g662_p),
    .din1(g290_n_spl_11),
    .din2(g661_n_spl_)
  );


  FA
  g_g663_n
  (
    .dout(g663_n),
    .din1(G136_p_spl_1),
    .din2(g630_n_spl_1)
  );


  FA
  g_g664_n
  (
    .dout(g664_n),
    .din1(G125_p_spl_1),
    .din2(g630_p_spl_1)
  );


  LA
  g_g665_p
  (
    .dout(g665_p),
    .din1(g663_n),
    .din2(g664_n)
  );


  FA
  g_g666_n
  (
    .dout(g666_n),
    .din1(g662_p),
    .din2(g665_p)
  );


  FA
  g_g667_n
  (
    .dout(g667_n),
    .din1(g240_n_spl_1),
    .din2(g666_n)
  );


  FA
  g_g668_n
  (
    .dout(g668_n),
    .din1(g290_n_spl_11),
    .din2(g661_n_spl_)
  );


  FA
  g_g669_n
  (
    .dout(g669_n),
    .din1(g255_p_spl_1),
    .din2(g656_n_spl_)
  );


  LA
  g_g670_p
  (
    .dout(g670_p),
    .din1(g668_n),
    .din2(g669_n)
  );


  LA
  g_g671_p
  (
    .dout(g671_p),
    .din1(g667_n),
    .din2(g670_p)
  );


  FA
  g_g672_n
  (
    .dout(g672_n),
    .din1(g658_n),
    .din2(g671_p)
  );


  LA
  g_g673_p
  (
    .dout(g673_p),
    .din1(g652_n),
    .din2(g672_n)
  );


  FA
  g_g674_n
  (
    .dout(g674_n),
    .din1(g648_p),
    .din2(g673_p)
  );


  LA
  g_g675_p
  (
    .dout(g675_p),
    .din1(g647_n),
    .din2(g674_n)
  );


  FA
  g_g676_n
  (
    .dout(g676_n),
    .din1(g642_p),
    .din2(g675_p)
  );


  LA
  g_g677_p
  (
    .dout(g677_p),
    .din1(g641_n),
    .din2(g676_n)
  );


  FA
  g_g678_n
  (
    .dout(g678_n),
    .din1(g636_p),
    .din2(g677_p)
  );


  LA
  g_g679_p
  (
    .dout(g679_p),
    .din1(g635_n),
    .din2(g678_n)
  );


  FA
  g_g680_n
  (
    .dout(g680_n),
    .din1(g634_p),
    .din2(g679_p)
  );


  LA
  g_g681_p
  (
    .dout(g681_p),
    .din1(g632_n),
    .din2(g680_n)
  );


  LA
  g_g682_p
  (
    .dout(g682_p),
    .din1(g628_n_spl_),
    .din2(g629_p_spl_)
  );


  FA
  g_g682_n
  (
    .dout(g682_n),
    .din1(g628_p_spl_),
    .din2(g629_n_spl_)
  );


  LA
  g_g683_p
  (
    .dout(g683_p),
    .din1(G136_n_spl_1),
    .din2(g682_p_spl_00)
  );


  FA
  g_g683_n
  (
    .dout(g683_n),
    .din1(G136_p_spl_1),
    .din2(g682_n_spl_00)
  );


  LA
  g_g684_p
  (
    .dout(g684_p),
    .din1(g427_p_spl_1),
    .din2(g682_p_spl_00)
  );


  FA
  g_g684_n
  (
    .dout(g684_n),
    .din1(g427_n_spl_1),
    .din2(g682_n_spl_00)
  );


  LA
  g_g685_p
  (
    .dout(g685_p),
    .din1(g683_n_spl_),
    .din2(g684_p_spl_)
  );


  LA
  g_g686_p
  (
    .dout(g686_p),
    .din1(G138_n_spl_1),
    .din2(g682_p_spl_01)
  );


  FA
  g_g686_n
  (
    .dout(g686_n),
    .din1(G138_p_spl_1),
    .din2(g682_n_spl_01)
  );


  LA
  g_g687_p
  (
    .dout(g687_p),
    .din1(g522_n_spl_1),
    .din2(g682_p_spl_01)
  );


  FA
  g_g687_n
  (
    .dout(g687_n),
    .din1(g522_p_spl_1),
    .din2(g682_n_spl_01)
  );


  LA
  g_g688_p
  (
    .dout(g688_p),
    .din1(g686_p),
    .din2(g687_n)
  );


  FA
  g_g688_n
  (
    .dout(g688_n),
    .din1(g686_n_spl_),
    .din2(g687_p_spl_)
  );


  LA
  g_g689_p
  (
    .dout(g689_p),
    .din1(g686_n_spl_),
    .din2(g687_p_spl_)
  );


  FA
  g_g690_n
  (
    .dout(g690_n),
    .din1(g688_p),
    .din2(g689_p)
  );


  LA
  g_g691_p
  (
    .dout(g691_p),
    .din1(g683_p),
    .din2(g684_n)
  );


  FA
  g_g691_n
  (
    .dout(g691_n),
    .din1(g683_n_spl_),
    .din2(g684_p_spl_)
  );


  FA
  g_g692_n
  (
    .dout(g692_n),
    .din1(g690_n_spl_),
    .din2(g691_p)
  );


  FA
  g_g693_n
  (
    .dout(g693_n),
    .din1(g685_p),
    .din2(g692_n)
  );


  LA
  g_g694_p
  (
    .dout(g694_p),
    .din1(G135_n_spl_1),
    .din2(g682_p_spl_10)
  );


  FA
  g_g694_n
  (
    .dout(g694_n),
    .din1(G135_p_spl_1),
    .din2(g682_n_spl_10)
  );


  LA
  g_g695_p
  (
    .dout(g695_p),
    .din1(g484_p_spl_1),
    .din2(g682_p_spl_10)
  );


  FA
  g_g695_n
  (
    .dout(g695_n),
    .din1(g484_n_spl_1),
    .din2(g682_n_spl_10)
  );


  LA
  g_g696_p
  (
    .dout(g696_p),
    .din1(g694_p),
    .din2(g695_n)
  );


  FA
  g_g696_n
  (
    .dout(g696_n),
    .din1(g694_n_spl_),
    .din2(g695_p_spl_)
  );


  LA
  g_g697_p
  (
    .dout(g697_p),
    .din1(g694_n_spl_),
    .din2(g695_p_spl_)
  );


  FA
  g_g698_n
  (
    .dout(g698_n),
    .din1(g696_p),
    .din2(g697_p)
  );


  LA
  g_g699_p
  (
    .dout(g699_p),
    .din1(g280_p_spl_1),
    .din2(g682_p_spl_11)
  );


  FA
  g_g699_n
  (
    .dout(g699_n),
    .din1(g280_n_spl_1),
    .din2(g682_n_spl_11)
  );


  LA
  g_g700_p
  (
    .dout(g700_p),
    .din1(G134_n_spl_1),
    .din2(g682_p_spl_11)
  );


  FA
  g_g700_n
  (
    .dout(g700_n),
    .din1(G134_p_spl_1),
    .din2(g682_n_spl_11)
  );


  LA
  g_g701_p
  (
    .dout(g701_p),
    .din1(g699_n),
    .din2(g700_p)
  );


  FA
  g_g701_n
  (
    .dout(g701_n),
    .din1(g699_p_spl_),
    .din2(g700_n_spl_)
  );


  LA
  g_g702_p
  (
    .dout(g702_p),
    .din1(g699_p_spl_),
    .din2(g700_n_spl_)
  );


  FA
  g_g703_n
  (
    .dout(g703_n),
    .din1(g701_p),
    .din2(g702_p)
  );


  FA
  g_g704_n
  (
    .dout(g704_n),
    .din1(g698_n_spl_),
    .din2(g703_n)
  );


  FA
  g_g705_n
  (
    .dout(g705_n),
    .din1(g693_n_spl_),
    .din2(g704_n)
  );


  FA
  g_g706_n
  (
    .dout(g706_n),
    .din1(g681_p),
    .din2(g705_n)
  );


  FA
  g_g707_n
  (
    .dout(g707_n),
    .din1(g698_n_spl_),
    .din2(g701_n)
  );


  LA
  g_g708_p
  (
    .dout(g708_p),
    .din1(g696_n),
    .din2(g707_n)
  );


  FA
  g_g709_n
  (
    .dout(g709_n),
    .din1(g693_n_spl_),
    .din2(g708_p)
  );


  FA
  g_g710_n
  (
    .dout(g710_n),
    .din1(g690_n_spl_),
    .din2(g691_n)
  );


  LA
  g_g711_p
  (
    .dout(g711_p),
    .din1(g709_n),
    .din2(g710_n)
  );


  LA
  g_g712_p
  (
    .dout(g712_p),
    .din1(g688_n),
    .din2(g711_p)
  );


  LA
  g_g713_p
  (
    .dout(g713_p),
    .din1(g706_n),
    .din2(g712_p)
  );


  FA
  g_g714_n
  (
    .dout(g714_n),
    .din1(g342_p_spl_),
    .din2(g361_p_spl_)
  );


  FA
  g_g715_n
  (
    .dout(g715_n),
    .din1(g388_p_spl_),
    .din2(g714_n)
  );


  FA
  g_g716_n
  (
    .dout(g716_n),
    .din1(g176_n_spl_0),
    .din2(g593_p_spl_)
  );


  FA
  g_g717_n
  (
    .dout(g717_n),
    .din1(g627_p_spl_),
    .din2(g716_n)
  );


  FA
  g_g718_n
  (
    .dout(g718_n),
    .din1(g715_n),
    .din2(g717_n)
  );


  buf

  (
    G2531_p,
    G115_n_spl_0
  );


  buf

  (
    G2532_p,
    G115_n_spl_1
  );


  buf

  (
    G2533_p,
    G115_n_spl_1
  );


  buf

  (
    G2534_p,
    G124_n_spl_
  );


  buf

  (
    G2535_p,
    G124_n_spl_
  );


  buf

  (
    G2536_p,
    G137_n_spl_0
  );


  buf

  (
    G2537_p,
    G137_n_spl_0
  );


  buf

  (
    G2538_p,
    G137_n_spl_
  );


  buf

  (
    G2539_p,
    G32_n_spl_
  );


  buf

  (
    G2540_p,
    G106_n_spl_
  );


  buf

  (
    G2541_p,
    G64_n_spl_
  );


  buf

  (
    G2542_p,
    G76_n_spl_
  );


  buf

  (
    G2543_p,
    G53_n_spl_
  );


  buf

  (
    G2544_p,
    G96_n_spl_
  );


  buf

  (
    G2545_p,
    G43_n_spl_
  );


  buf

  (
    G2546_p,
    G86_n_spl_
  );


  buf

  (
    G2547_p,
    g160_n
  );


  buf

  (
    G2548_p,
    g162_n
  );


  buf

  (
    G2549_p,
    G115_p
  );


  buf

  (
    G2550_p,
    g163_p
  );


  buf

  (
    G2551_p,
    g164_n_spl_
  );


  buf

  (
    G2552_p,
    g165_n
  );


  buf

  (
    G2553_p,
    g166_n
  );


  buf

  (
    G2554_p,
    g173_n_spl_
  );


  buf

  (
    G2555_p,
    g173_n_spl_
  );


  buf

  (
    G2556_p,
    g176_n_spl_
  );


  buf

  (
    G2557_p,
    g185_n_spl_1
  );


  buf

  (
    G2558_p,
    g194_n_spl_1
  );


  buf

  (
    G2559_p,
    g203_n_spl_1
  );


  buf

  (
    G2560_p,
    g213_p_spl_1
  );


  buf

  (
    G2561_p,
    g222_p_spl_1
  );


  buf

  (
    G2562_p,
    g231_p_spl_1
  );


  buf

  (
    G2563_p,
    g241_n
  );


  buf

  (
    G2564_p,
    g244_n
  );


  buf

  (
    G2565_p,
    g246_n
  );


  buf

  (
    G2566_p,
    g255_n_spl_1
  );


  buf

  (
    G2567_p,
    g231_n_spl_1
  );


  buf

  (
    G2568_p,
    g222_n_spl_1
  );


  buf

  (
    G2569_p,
    g213_n_spl_1
  );


  buf

  (
    G2570_p,
    g262_p_spl_1
  );


  buf

  (
    G2571_p,
    g271_n_spl_1
  );


  buf

  (
    G2572_p,
    g280_n_spl_1
  );


  buf

  (
    G2573_p,
    g292_n_spl_
  );


  buf

  (
    G2574_p,
    g292_n_spl_
  );


  buf

  (
    G2575_p,
    g295_n_spl_
  );


  buf

  (
    G2576_p,
    g295_n_spl_
  );


  buf

  (
    G2577_p,
    g297_n
  );


  buf

  (
    G2578_p,
    g301_n_spl_
  );


  buf

  (
    G2579_p,
    g301_n_spl_
  );


  buf

  (
    G2580_p,
    g314_n
  );


  buf

  (
    G2581_n,
    g342_p_spl_
  );


  buf

  (
    G2582_p,
    g361_p_spl_
  );


  buf

  (
    G2583_p,
    g388_p_spl_
  );


  buf

  (
    G2584_p,
    g540_n_spl_
  );


  buf

  (
    G2585_p,
    g540_n_spl_
  );


  buf

  (
    G2586_p,
    g559_n
  );


  buf

  (
    G2587_n,
    g593_p_spl_
  );


  buf

  (
    G2588_p,
    g617_p_spl_
  );


  buf

  (
    G2589_p,
    g617_p_spl_
  );


  buf

  (
    G2590_n,
    g627_p_spl_
  );


  buf

  (
    G2591_p,
    g713_p
  );


  buf

  (
    G2592_p,
    1'b0
  );


  buf

  (
    G2593_p,
    g718_n_spl_
  );


  buf

  (
    G2594_p,
    g718_n_spl_
  );


  buf

  (
    G141_p_spl_,
    G141_p
  );


  buf

  (
    G141_p_spl_0,
    G141_p_spl_
  );


  buf

  (
    G141_p_spl_1,
    G141_p_spl_
  );


  buf

  (
    G142_p_spl_,
    G142_p
  );


  buf

  (
    G142_p_spl_0,
    G142_p_spl_
  );


  buf

  (
    G142_p_spl_1,
    G142_p_spl_
  );


  buf

  (
    G141_n_spl_,
    G141_n
  );


  buf

  (
    G141_n_spl_0,
    G141_n_spl_
  );


  buf

  (
    G142_n_spl_,
    G142_n
  );


  buf

  (
    G142_n_spl_0,
    G142_n_spl_
  );


  buf

  (
    G139_p_spl_,
    G139_p
  );


  buf

  (
    G139_p_spl_0,
    G139_p_spl_
  );


  buf

  (
    G139_p_spl_1,
    G139_p_spl_
  );


  buf

  (
    G140_p_spl_,
    G140_p
  );


  buf

  (
    G140_p_spl_0,
    G140_p_spl_
  );


  buf

  (
    G140_p_spl_1,
    G140_p_spl_
  );


  buf

  (
    G139_n_spl_,
    G139_n
  );


  buf

  (
    G139_n_spl_0,
    G139_n_spl_
  );


  buf

  (
    G140_n_spl_,
    G140_n
  );


  buf

  (
    G140_n_spl_0,
    G140_n_spl_
  );


  buf

  (
    g158_n_spl_,
    g158_n
  );


  buf

  (
    g159_n_spl_,
    g159_n
  );


  buf

  (
    G121_n_spl_,
    G121_n
  );


  buf

  (
    G115_n_spl_,
    G115_n
  );


  buf

  (
    G115_n_spl_0,
    G115_n_spl_
  );


  buf

  (
    G115_n_spl_1,
    G115_n_spl_
  );


  buf

  (
    g164_n_spl_,
    g164_n
  );


  buf

  (
    g164_n_spl_0,
    g164_n_spl_
  );


  buf

  (
    G43_n_spl_,
    G43_n
  );


  buf

  (
    G53_n_spl_,
    G53_n
  );


  buf

  (
    G86_n_spl_,
    G86_n
  );


  buf

  (
    G96_n_spl_,
    G96_n
  );


  buf

  (
    G32_n_spl_,
    G32_n
  );


  buf

  (
    G64_n_spl_,
    G64_n
  );


  buf

  (
    G76_n_spl_,
    G76_n
  );


  buf

  (
    G106_n_spl_,
    G106_n
  );


  buf

  (
    g169_n_spl_,
    g169_n
  );


  buf

  (
    g172_n_spl_,
    g172_n
  );


  buf

  (
    G145_n_spl_,
    G145_n
  );


  buf

  (
    G145_n_spl_0,
    G145_n_spl_
  );


  buf

  (
    G145_n_spl_00,
    G145_n_spl_0
  );


  buf

  (
    G145_n_spl_000,
    G145_n_spl_00
  );


  buf

  (
    G145_n_spl_0000,
    G145_n_spl_000
  );


  buf

  (
    G145_n_spl_00000,
    G145_n_spl_0000
  );


  buf

  (
    G145_n_spl_00001,
    G145_n_spl_0000
  );


  buf

  (
    G145_n_spl_0001,
    G145_n_spl_000
  );


  buf

  (
    G145_n_spl_00010,
    G145_n_spl_0001
  );


  buf

  (
    G145_n_spl_00011,
    G145_n_spl_0001
  );


  buf

  (
    G145_n_spl_001,
    G145_n_spl_00
  );


  buf

  (
    G145_n_spl_0010,
    G145_n_spl_001
  );


  buf

  (
    G145_n_spl_0011,
    G145_n_spl_001
  );


  buf

  (
    G145_n_spl_01,
    G145_n_spl_0
  );


  buf

  (
    G145_n_spl_010,
    G145_n_spl_01
  );


  buf

  (
    G145_n_spl_0100,
    G145_n_spl_010
  );


  buf

  (
    G145_n_spl_0101,
    G145_n_spl_010
  );


  buf

  (
    G145_n_spl_011,
    G145_n_spl_01
  );


  buf

  (
    G145_n_spl_0110,
    G145_n_spl_011
  );


  buf

  (
    G145_n_spl_0111,
    G145_n_spl_011
  );


  buf

  (
    G145_n_spl_1,
    G145_n_spl_
  );


  buf

  (
    G145_n_spl_10,
    G145_n_spl_1
  );


  buf

  (
    G145_n_spl_100,
    G145_n_spl_10
  );


  buf

  (
    G145_n_spl_1000,
    G145_n_spl_100
  );


  buf

  (
    G145_n_spl_1001,
    G145_n_spl_100
  );


  buf

  (
    G145_n_spl_101,
    G145_n_spl_10
  );


  buf

  (
    G145_n_spl_1010,
    G145_n_spl_101
  );


  buf

  (
    G145_n_spl_1011,
    G145_n_spl_101
  );


  buf

  (
    G145_n_spl_11,
    G145_n_spl_1
  );


  buf

  (
    G145_n_spl_110,
    G145_n_spl_11
  );


  buf

  (
    G145_n_spl_1100,
    G145_n_spl_110
  );


  buf

  (
    G145_n_spl_1101,
    G145_n_spl_110
  );


  buf

  (
    G145_n_spl_111,
    G145_n_spl_11
  );


  buf

  (
    G145_n_spl_1110,
    G145_n_spl_111
  );


  buf

  (
    G145_n_spl_1111,
    G145_n_spl_111
  );


  buf

  (
    G145_p_spl_,
    G145_p
  );


  buf

  (
    G145_p_spl_0,
    G145_p_spl_
  );


  buf

  (
    G145_p_spl_00,
    G145_p_spl_0
  );


  buf

  (
    G145_p_spl_000,
    G145_p_spl_00
  );


  buf

  (
    G145_p_spl_0000,
    G145_p_spl_000
  );


  buf

  (
    G145_p_spl_00000,
    G145_p_spl_0000
  );


  buf

  (
    G145_p_spl_00001,
    G145_p_spl_0000
  );


  buf

  (
    G145_p_spl_0001,
    G145_p_spl_000
  );


  buf

  (
    G145_p_spl_00010,
    G145_p_spl_0001
  );


  buf

  (
    G145_p_spl_00011,
    G145_p_spl_0001
  );


  buf

  (
    G145_p_spl_001,
    G145_p_spl_00
  );


  buf

  (
    G145_p_spl_0010,
    G145_p_spl_001
  );


  buf

  (
    G145_p_spl_0011,
    G145_p_spl_001
  );


  buf

  (
    G145_p_spl_01,
    G145_p_spl_0
  );


  buf

  (
    G145_p_spl_010,
    G145_p_spl_01
  );


  buf

  (
    G145_p_spl_0100,
    G145_p_spl_010
  );


  buf

  (
    G145_p_spl_0101,
    G145_p_spl_010
  );


  buf

  (
    G145_p_spl_011,
    G145_p_spl_01
  );


  buf

  (
    G145_p_spl_0110,
    G145_p_spl_011
  );


  buf

  (
    G145_p_spl_0111,
    G145_p_spl_011
  );


  buf

  (
    G145_p_spl_1,
    G145_p_spl_
  );


  buf

  (
    G145_p_spl_10,
    G145_p_spl_1
  );


  buf

  (
    G145_p_spl_100,
    G145_p_spl_10
  );


  buf

  (
    G145_p_spl_1000,
    G145_p_spl_100
  );


  buf

  (
    G145_p_spl_1001,
    G145_p_spl_100
  );


  buf

  (
    G145_p_spl_101,
    G145_p_spl_10
  );


  buf

  (
    G145_p_spl_1010,
    G145_p_spl_101
  );


  buf

  (
    G145_p_spl_1011,
    G145_p_spl_101
  );


  buf

  (
    G145_p_spl_11,
    G145_p_spl_1
  );


  buf

  (
    G145_p_spl_110,
    G145_p_spl_11
  );


  buf

  (
    G145_p_spl_1100,
    G145_p_spl_110
  );


  buf

  (
    G145_p_spl_1101,
    G145_p_spl_110
  );


  buf

  (
    G145_p_spl_111,
    G145_p_spl_11
  );


  buf

  (
    G145_p_spl_1110,
    G145_p_spl_111
  );


  buf

  (
    G145_p_spl_1111,
    G145_p_spl_111
  );


  buf

  (
    G146_p_spl_,
    G146_p
  );


  buf

  (
    G146_p_spl_0,
    G146_p_spl_
  );


  buf

  (
    G146_p_spl_00,
    G146_p_spl_0
  );


  buf

  (
    G146_p_spl_000,
    G146_p_spl_00
  );


  buf

  (
    G146_p_spl_0000,
    G146_p_spl_000
  );


  buf

  (
    G146_p_spl_0001,
    G146_p_spl_000
  );


  buf

  (
    G146_p_spl_001,
    G146_p_spl_00
  );


  buf

  (
    G146_p_spl_01,
    G146_p_spl_0
  );


  buf

  (
    G146_p_spl_010,
    G146_p_spl_01
  );


  buf

  (
    G146_p_spl_011,
    G146_p_spl_01
  );


  buf

  (
    G146_p_spl_1,
    G146_p_spl_
  );


  buf

  (
    G146_p_spl_10,
    G146_p_spl_1
  );


  buf

  (
    G146_p_spl_100,
    G146_p_spl_10
  );


  buf

  (
    G146_p_spl_101,
    G146_p_spl_10
  );


  buf

  (
    G146_p_spl_11,
    G146_p_spl_1
  );


  buf

  (
    G146_p_spl_110,
    G146_p_spl_11
  );


  buf

  (
    G146_p_spl_111,
    G146_p_spl_11
  );


  buf

  (
    G146_n_spl_,
    G146_n
  );


  buf

  (
    G146_n_spl_0,
    G146_n_spl_
  );


  buf

  (
    G146_n_spl_00,
    G146_n_spl_0
  );


  buf

  (
    G146_n_spl_000,
    G146_n_spl_00
  );


  buf

  (
    G146_n_spl_0000,
    G146_n_spl_000
  );


  buf

  (
    G146_n_spl_0001,
    G146_n_spl_000
  );


  buf

  (
    G146_n_spl_001,
    G146_n_spl_00
  );


  buf

  (
    G146_n_spl_01,
    G146_n_spl_0
  );


  buf

  (
    G146_n_spl_010,
    G146_n_spl_01
  );


  buf

  (
    G146_n_spl_011,
    G146_n_spl_01
  );


  buf

  (
    G146_n_spl_1,
    G146_n_spl_
  );


  buf

  (
    G146_n_spl_10,
    G146_n_spl_1
  );


  buf

  (
    G146_n_spl_100,
    G146_n_spl_10
  );


  buf

  (
    G146_n_spl_101,
    G146_n_spl_10
  );


  buf

  (
    G146_n_spl_11,
    G146_n_spl_1
  );


  buf

  (
    G146_n_spl_110,
    G146_n_spl_11
  );


  buf

  (
    G146_n_spl_111,
    G146_n_spl_11
  );


  buf

  (
    G117_p_spl_,
    G117_p
  );


  buf

  (
    G117_p_spl_0,
    G117_p_spl_
  );


  buf

  (
    G117_p_spl_00,
    G117_p_spl_0
  );


  buf

  (
    G117_p_spl_000,
    G117_p_spl_00
  );


  buf

  (
    G117_p_spl_0000,
    G117_p_spl_000
  );


  buf

  (
    G117_p_spl_0001,
    G117_p_spl_000
  );


  buf

  (
    G117_p_spl_001,
    G117_p_spl_00
  );


  buf

  (
    G117_p_spl_0010,
    G117_p_spl_001
  );


  buf

  (
    G117_p_spl_0011,
    G117_p_spl_001
  );


  buf

  (
    G117_p_spl_01,
    G117_p_spl_0
  );


  buf

  (
    G117_p_spl_010,
    G117_p_spl_01
  );


  buf

  (
    G117_p_spl_0100,
    G117_p_spl_010
  );


  buf

  (
    G117_p_spl_0101,
    G117_p_spl_010
  );


  buf

  (
    G117_p_spl_011,
    G117_p_spl_01
  );


  buf

  (
    G117_p_spl_0110,
    G117_p_spl_011
  );


  buf

  (
    G117_p_spl_0111,
    G117_p_spl_011
  );


  buf

  (
    G117_p_spl_1,
    G117_p_spl_
  );


  buf

  (
    G117_p_spl_10,
    G117_p_spl_1
  );


  buf

  (
    G117_p_spl_100,
    G117_p_spl_10
  );


  buf

  (
    G117_p_spl_1000,
    G117_p_spl_100
  );


  buf

  (
    G117_p_spl_1001,
    G117_p_spl_100
  );


  buf

  (
    G117_p_spl_101,
    G117_p_spl_10
  );


  buf

  (
    G117_p_spl_1010,
    G117_p_spl_101
  );


  buf

  (
    G117_p_spl_1011,
    G117_p_spl_101
  );


  buf

  (
    G117_p_spl_11,
    G117_p_spl_1
  );


  buf

  (
    G117_p_spl_110,
    G117_p_spl_11
  );


  buf

  (
    G117_p_spl_1100,
    G117_p_spl_110
  );


  buf

  (
    G117_p_spl_1101,
    G117_p_spl_110
  );


  buf

  (
    G117_p_spl_111,
    G117_p_spl_11
  );


  buf

  (
    G117_p_spl_1110,
    G117_p_spl_111
  );


  buf

  (
    G120_n_spl_,
    G120_n
  );


  buf

  (
    G120_n_spl_0,
    G120_n_spl_
  );


  buf

  (
    G120_n_spl_00,
    G120_n_spl_0
  );


  buf

  (
    G120_n_spl_000,
    G120_n_spl_00
  );


  buf

  (
    G120_n_spl_0000,
    G120_n_spl_000
  );


  buf

  (
    G120_n_spl_0001,
    G120_n_spl_000
  );


  buf

  (
    G120_n_spl_001,
    G120_n_spl_00
  );


  buf

  (
    G120_n_spl_0010,
    G120_n_spl_001
  );


  buf

  (
    G120_n_spl_0011,
    G120_n_spl_001
  );


  buf

  (
    G120_n_spl_01,
    G120_n_spl_0
  );


  buf

  (
    G120_n_spl_010,
    G120_n_spl_01
  );


  buf

  (
    G120_n_spl_0100,
    G120_n_spl_010
  );


  buf

  (
    G120_n_spl_011,
    G120_n_spl_01
  );


  buf

  (
    G120_n_spl_1,
    G120_n_spl_
  );


  buf

  (
    G120_n_spl_10,
    G120_n_spl_1
  );


  buf

  (
    G120_n_spl_100,
    G120_n_spl_10
  );


  buf

  (
    G120_n_spl_101,
    G120_n_spl_10
  );


  buf

  (
    G120_n_spl_11,
    G120_n_spl_1
  );


  buf

  (
    G120_n_spl_110,
    G120_n_spl_11
  );


  buf

  (
    G120_n_spl_111,
    G120_n_spl_11
  );


  buf

  (
    G117_n_spl_,
    G117_n
  );


  buf

  (
    G117_n_spl_0,
    G117_n_spl_
  );


  buf

  (
    G117_n_spl_00,
    G117_n_spl_0
  );


  buf

  (
    G117_n_spl_000,
    G117_n_spl_00
  );


  buf

  (
    G117_n_spl_0000,
    G117_n_spl_000
  );


  buf

  (
    G117_n_spl_0001,
    G117_n_spl_000
  );


  buf

  (
    G117_n_spl_001,
    G117_n_spl_00
  );


  buf

  (
    G117_n_spl_0010,
    G117_n_spl_001
  );


  buf

  (
    G117_n_spl_0011,
    G117_n_spl_001
  );


  buf

  (
    G117_n_spl_01,
    G117_n_spl_0
  );


  buf

  (
    G117_n_spl_010,
    G117_n_spl_01
  );


  buf

  (
    G117_n_spl_0100,
    G117_n_spl_010
  );


  buf

  (
    G117_n_spl_0101,
    G117_n_spl_010
  );


  buf

  (
    G117_n_spl_011,
    G117_n_spl_01
  );


  buf

  (
    G117_n_spl_0110,
    G117_n_spl_011
  );


  buf

  (
    G117_n_spl_0111,
    G117_n_spl_011
  );


  buf

  (
    G117_n_spl_1,
    G117_n_spl_
  );


  buf

  (
    G117_n_spl_10,
    G117_n_spl_1
  );


  buf

  (
    G117_n_spl_100,
    G117_n_spl_10
  );


  buf

  (
    G117_n_spl_1000,
    G117_n_spl_100
  );


  buf

  (
    G117_n_spl_1001,
    G117_n_spl_100
  );


  buf

  (
    G117_n_spl_101,
    G117_n_spl_10
  );


  buf

  (
    G117_n_spl_1010,
    G117_n_spl_101
  );


  buf

  (
    G117_n_spl_1011,
    G117_n_spl_101
  );


  buf

  (
    G117_n_spl_11,
    G117_n_spl_1
  );


  buf

  (
    G117_n_spl_110,
    G117_n_spl_11
  );


  buf

  (
    G117_n_spl_1100,
    G117_n_spl_110
  );


  buf

  (
    G117_n_spl_1101,
    G117_n_spl_110
  );


  buf

  (
    G117_n_spl_111,
    G117_n_spl_11
  );


  buf

  (
    G117_n_spl_1110,
    G117_n_spl_111
  );


  buf

  (
    G120_p_spl_,
    G120_p
  );


  buf

  (
    G120_p_spl_0,
    G120_p_spl_
  );


  buf

  (
    G120_p_spl_00,
    G120_p_spl_0
  );


  buf

  (
    G120_p_spl_000,
    G120_p_spl_00
  );


  buf

  (
    G120_p_spl_0000,
    G120_p_spl_000
  );


  buf

  (
    G120_p_spl_0001,
    G120_p_spl_000
  );


  buf

  (
    G120_p_spl_001,
    G120_p_spl_00
  );


  buf

  (
    G120_p_spl_0010,
    G120_p_spl_001
  );


  buf

  (
    G120_p_spl_0011,
    G120_p_spl_001
  );


  buf

  (
    G120_p_spl_01,
    G120_p_spl_0
  );


  buf

  (
    G120_p_spl_010,
    G120_p_spl_01
  );


  buf

  (
    G120_p_spl_0100,
    G120_p_spl_010
  );


  buf

  (
    G120_p_spl_011,
    G120_p_spl_01
  );


  buf

  (
    G120_p_spl_1,
    G120_p_spl_
  );


  buf

  (
    G120_p_spl_10,
    G120_p_spl_1
  );


  buf

  (
    G120_p_spl_100,
    G120_p_spl_10
  );


  buf

  (
    G120_p_spl_101,
    G120_p_spl_10
  );


  buf

  (
    G120_p_spl_11,
    G120_p_spl_1
  );


  buf

  (
    G120_p_spl_110,
    G120_p_spl_11
  );


  buf

  (
    G120_p_spl_111,
    G120_p_spl_11
  );


  buf

  (
    g204_p_spl_,
    g204_p
  );


  buf

  (
    g204_p_spl_0,
    g204_p_spl_
  );


  buf

  (
    g204_p_spl_00,
    g204_p_spl_0
  );


  buf

  (
    g204_p_spl_000,
    g204_p_spl_00
  );


  buf

  (
    g204_p_spl_01,
    g204_p_spl_0
  );


  buf

  (
    g204_p_spl_1,
    g204_p_spl_
  );


  buf

  (
    g204_p_spl_10,
    g204_p_spl_1
  );


  buf

  (
    g204_p_spl_11,
    g204_p_spl_1
  );


  buf

  (
    g204_n_spl_,
    g204_n
  );


  buf

  (
    g204_n_spl_0,
    g204_n_spl_
  );


  buf

  (
    g204_n_spl_00,
    g204_n_spl_0
  );


  buf

  (
    g204_n_spl_000,
    g204_n_spl_00
  );


  buf

  (
    g204_n_spl_01,
    g204_n_spl_0
  );


  buf

  (
    g204_n_spl_1,
    g204_n_spl_
  );


  buf

  (
    g204_n_spl_10,
    g204_n_spl_1
  );


  buf

  (
    g204_n_spl_11,
    g204_n_spl_1
  );


  buf

  (
    G122_n_spl_,
    G122_n
  );


  buf

  (
    G122_n_spl_0,
    G122_n_spl_
  );


  buf

  (
    g240_n_spl_,
    g240_n
  );


  buf

  (
    g240_n_spl_0,
    g240_n_spl_
  );


  buf

  (
    g240_n_spl_00,
    g240_n_spl_0
  );


  buf

  (
    g240_n_spl_1,
    g240_n_spl_
  );


  buf

  (
    g176_n_spl_,
    g176_n
  );


  buf

  (
    g176_n_spl_0,
    g176_n_spl_
  );


  buf

  (
    g243_n_spl_,
    g243_n
  );


  buf

  (
    G123_p_spl_,
    G123_p
  );


  buf

  (
    G123_p_spl_0,
    G123_p_spl_
  );


  buf

  (
    G123_p_spl_1,
    G123_p_spl_
  );


  buf

  (
    g231_n_spl_,
    g231_n
  );


  buf

  (
    g231_n_spl_0,
    g231_n_spl_
  );


  buf

  (
    g231_n_spl_00,
    g231_n_spl_0
  );


  buf

  (
    g231_n_spl_1,
    g231_n_spl_
  );


  buf

  (
    G123_n_spl_,
    G123_n
  );


  buf

  (
    G123_n_spl_0,
    G123_n_spl_
  );


  buf

  (
    G123_n_spl_1,
    G123_n_spl_
  );


  buf

  (
    g290_p_spl_,
    g290_p
  );


  buf

  (
    g290_p_spl_0,
    g290_p_spl_
  );


  buf

  (
    g290_p_spl_00,
    g290_p_spl_0
  );


  buf

  (
    g290_p_spl_01,
    g290_p_spl_0
  );


  buf

  (
    g290_p_spl_1,
    g290_p_spl_
  );


  buf

  (
    g222_p_spl_,
    g222_p
  );


  buf

  (
    g222_p_spl_0,
    g222_p_spl_
  );


  buf

  (
    g222_p_spl_00,
    g222_p_spl_0
  );


  buf

  (
    g222_p_spl_01,
    g222_p_spl_0
  );


  buf

  (
    g222_p_spl_1,
    g222_p_spl_
  );


  buf

  (
    g255_n_spl_,
    g255_n
  );


  buf

  (
    g255_n_spl_0,
    g255_n_spl_
  );


  buf

  (
    g255_n_spl_00,
    g255_n_spl_0
  );


  buf

  (
    g255_n_spl_1,
    g255_n_spl_
  );


  buf

  (
    G118_p_spl_,
    G118_p
  );


  buf

  (
    G118_p_spl_0,
    G118_p_spl_
  );


  buf

  (
    g290_n_spl_,
    g290_n
  );


  buf

  (
    g290_n_spl_0,
    g290_n_spl_
  );


  buf

  (
    g290_n_spl_00,
    g290_n_spl_0
  );


  buf

  (
    g290_n_spl_01,
    g290_n_spl_0
  );


  buf

  (
    g290_n_spl_1,
    g290_n_spl_
  );


  buf

  (
    g290_n_spl_10,
    g290_n_spl_1
  );


  buf

  (
    g290_n_spl_11,
    g290_n_spl_1
  );


  buf

  (
    G118_n_spl_,
    G118_n
  );


  buf

  (
    g298_p_spl_,
    g298_p
  );


  buf

  (
    g298_p_spl_0,
    g298_p_spl_
  );


  buf

  (
    g240_p_spl_,
    g240_p
  );


  buf

  (
    g240_p_spl_0,
    g240_p_spl_
  );


  buf

  (
    g240_p_spl_1,
    g240_p_spl_
  );


  buf

  (
    G143_n_spl_,
    G143_n
  );


  buf

  (
    G143_n_spl_0,
    G143_n_spl_
  );


  buf

  (
    g310_p_spl_,
    g310_p
  );


  buf

  (
    g310_p_spl_0,
    g310_p_spl_
  );


  buf

  (
    G143_p_spl_,
    G143_p
  );


  buf

  (
    G143_p_spl_0,
    G143_p_spl_
  );


  buf

  (
    g310_n_spl_,
    g310_n
  );


  buf

  (
    g310_n_spl_0,
    g310_n_spl_
  );


  buf

  (
    g310_n_spl_1,
    g310_n_spl_
  );


  buf

  (
    G144_p_spl_,
    G144_p
  );


  buf

  (
    G144_p_spl_0,
    G144_p_spl_
  );


  buf

  (
    G154_n_spl_,
    G154_n
  );


  buf

  (
    G155_n_spl_,
    G155_n
  );


  buf

  (
    G154_p_spl_,
    G154_p
  );


  buf

  (
    G155_p_spl_,
    G155_p
  );


  buf

  (
    G125_n_spl_,
    G125_n
  );


  buf

  (
    G125_n_spl_0,
    G125_n_spl_
  );


  buf

  (
    G126_n_spl_,
    G126_n
  );


  buf

  (
    G126_n_spl_0,
    G126_n_spl_
  );


  buf

  (
    G125_p_spl_,
    G125_p
  );


  buf

  (
    G125_p_spl_0,
    G125_p_spl_
  );


  buf

  (
    G125_p_spl_1,
    G125_p_spl_
  );


  buf

  (
    G126_p_spl_,
    G126_p
  );


  buf

  (
    G126_p_spl_0,
    G126_p_spl_
  );


  buf

  (
    G126_p_spl_1,
    G126_p_spl_
  );


  buf

  (
    g317_p_spl_,
    g317_p
  );


  buf

  (
    g320_n_spl_,
    g320_n
  );


  buf

  (
    g317_n_spl_,
    g317_n
  );


  buf

  (
    g320_p_spl_,
    g320_p
  );


  buf

  (
    G152_n_spl_,
    G152_n
  );


  buf

  (
    G153_n_spl_,
    G153_n
  );


  buf

  (
    G152_p_spl_,
    G152_p
  );


  buf

  (
    G153_p_spl_,
    G153_p
  );


  buf

  (
    G148_n_spl_,
    G148_n
  );


  buf

  (
    G149_n_spl_,
    G149_n
  );


  buf

  (
    G148_p_spl_,
    G148_p
  );


  buf

  (
    G149_p_spl_,
    G149_p
  );


  buf

  (
    g326_n_spl_,
    g326_n
  );


  buf

  (
    g329_n_spl_,
    g329_n
  );


  buf

  (
    g326_p_spl_,
    g326_p
  );


  buf

  (
    g329_p_spl_,
    g329_p
  );


  buf

  (
    G150_n_spl_,
    G150_n
  );


  buf

  (
    G151_n_spl_,
    G151_n
  );


  buf

  (
    G150_p_spl_,
    G150_p
  );


  buf

  (
    G151_p_spl_,
    G151_p
  );


  buf

  (
    g332_n_spl_,
    g332_n
  );


  buf

  (
    g335_n_spl_,
    g335_n
  );


  buf

  (
    g332_p_spl_,
    g332_p
  );


  buf

  (
    g335_p_spl_,
    g335_p
  );


  buf

  (
    G138_p_spl_,
    G138_p
  );


  buf

  (
    G138_p_spl_0,
    G138_p_spl_
  );


  buf

  (
    G138_p_spl_00,
    G138_p_spl_0
  );


  buf

  (
    G138_p_spl_1,
    G138_p_spl_
  );


  buf

  (
    G157_n_spl_,
    G157_n
  );


  buf

  (
    G138_n_spl_,
    G138_n
  );


  buf

  (
    G138_n_spl_0,
    G138_n_spl_
  );


  buf

  (
    G138_n_spl_1,
    G138_n_spl_
  );


  buf

  (
    G157_p_spl_,
    G157_p
  );


  buf

  (
    g346_n_spl_,
    g346_n
  );


  buf

  (
    g349_n_spl_,
    g349_n
  );


  buf

  (
    g346_p_spl_,
    g346_p
  );


  buf

  (
    g349_p_spl_,
    g349_p
  );


  buf

  (
    g344_n_spl_,
    g344_n
  );


  buf

  (
    g352_n_spl_,
    g352_n
  );


  buf

  (
    g344_p_spl_,
    g344_p
  );


  buf

  (
    g352_p_spl_,
    g352_p
  );


  buf

  (
    G144_n_spl_,
    G144_n
  );


  buf

  (
    G133_n_spl_,
    G133_n
  );


  buf

  (
    G133_n_spl_0,
    G133_n_spl_
  );


  buf

  (
    G134_n_spl_,
    G134_n
  );


  buf

  (
    G134_n_spl_0,
    G134_n_spl_
  );


  buf

  (
    G134_n_spl_1,
    G134_n_spl_
  );


  buf

  (
    G133_p_spl_,
    G133_p
  );


  buf

  (
    G133_p_spl_0,
    G133_p_spl_
  );


  buf

  (
    G133_p_spl_1,
    G133_p_spl_
  );


  buf

  (
    G134_p_spl_,
    G134_p
  );


  buf

  (
    G134_p_spl_0,
    G134_p_spl_
  );


  buf

  (
    G134_p_spl_1,
    G134_p_spl_
  );


  buf

  (
    G135_n_spl_,
    G135_n
  );


  buf

  (
    G135_n_spl_0,
    G135_n_spl_
  );


  buf

  (
    G135_n_spl_1,
    G135_n_spl_
  );


  buf

  (
    G136_n_spl_,
    G136_n
  );


  buf

  (
    G136_n_spl_0,
    G136_n_spl_
  );


  buf

  (
    G136_n_spl_1,
    G136_n_spl_
  );


  buf

  (
    G135_p_spl_,
    G135_p
  );


  buf

  (
    G135_p_spl_0,
    G135_p_spl_
  );


  buf

  (
    G135_p_spl_1,
    G135_p_spl_
  );


  buf

  (
    G136_p_spl_,
    G136_p
  );


  buf

  (
    G136_p_spl_0,
    G136_p_spl_
  );


  buf

  (
    G136_p_spl_00,
    G136_p_spl_0
  );


  buf

  (
    G136_p_spl_1,
    G136_p_spl_
  );


  buf

  (
    g364_p_spl_,
    g364_p
  );


  buf

  (
    g367_n_spl_,
    g367_n
  );


  buf

  (
    g364_n_spl_,
    g364_n
  );


  buf

  (
    g367_p_spl_,
    g367_p
  );


  buf

  (
    G131_n_spl_,
    G131_n
  );


  buf

  (
    G131_n_spl_0,
    G131_n_spl_
  );


  buf

  (
    G132_n_spl_,
    G132_n
  );


  buf

  (
    G132_n_spl_0,
    G132_n_spl_
  );


  buf

  (
    G131_p_spl_,
    G131_p
  );


  buf

  (
    G131_p_spl_0,
    G131_p_spl_
  );


  buf

  (
    G131_p_spl_1,
    G131_p_spl_
  );


  buf

  (
    G132_p_spl_,
    G132_p
  );


  buf

  (
    G132_p_spl_0,
    G132_p_spl_
  );


  buf

  (
    G132_p_spl_1,
    G132_p_spl_
  );


  buf

  (
    G128_p_spl_,
    G128_p
  );


  buf

  (
    G128_p_spl_0,
    G128_p_spl_
  );


  buf

  (
    G128_p_spl_1,
    G128_p_spl_
  );


  buf

  (
    G156_n_spl_,
    G156_n
  );


  buf

  (
    G128_n_spl_,
    G128_n
  );


  buf

  (
    G128_n_spl_0,
    G128_n_spl_
  );


  buf

  (
    G156_p_spl_,
    G156_p
  );


  buf

  (
    g373_n_spl_,
    g373_n
  );


  buf

  (
    g376_n_spl_,
    g376_n
  );


  buf

  (
    g373_p_spl_,
    g373_p
  );


  buf

  (
    g376_p_spl_,
    g376_p
  );


  buf

  (
    G129_n_spl_,
    G129_n
  );


  buf

  (
    G129_n_spl_0,
    G129_n_spl_
  );


  buf

  (
    G130_n_spl_,
    G130_n
  );


  buf

  (
    G130_n_spl_0,
    G130_n_spl_
  );


  buf

  (
    G129_p_spl_,
    G129_p
  );


  buf

  (
    G129_p_spl_0,
    G129_p_spl_
  );


  buf

  (
    G129_p_spl_1,
    G129_p_spl_
  );


  buf

  (
    G130_p_spl_,
    G130_p
  );


  buf

  (
    G130_p_spl_0,
    G130_p_spl_
  );


  buf

  (
    G130_p_spl_1,
    G130_p_spl_
  );


  buf

  (
    g379_n_spl_,
    g379_n
  );


  buf

  (
    g382_n_spl_,
    g382_n
  );


  buf

  (
    g379_p_spl_,
    g379_p
  );


  buf

  (
    g382_p_spl_,
    g382_p
  );


  buf

  (
    G12_n_spl_,
    G12_n
  );


  buf

  (
    G12_n_spl_0,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_00,
    G12_n_spl_0
  );


  buf

  (
    G12_n_spl_000,
    G12_n_spl_00
  );


  buf

  (
    G12_n_spl_0000,
    G12_n_spl_000
  );


  buf

  (
    G12_n_spl_0001,
    G12_n_spl_000
  );


  buf

  (
    G12_n_spl_001,
    G12_n_spl_00
  );


  buf

  (
    G12_n_spl_01,
    G12_n_spl_0
  );


  buf

  (
    G12_n_spl_010,
    G12_n_spl_01
  );


  buf

  (
    G12_n_spl_011,
    G12_n_spl_01
  );


  buf

  (
    G12_n_spl_1,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_10,
    G12_n_spl_1
  );


  buf

  (
    G12_n_spl_100,
    G12_n_spl_10
  );


  buf

  (
    G12_n_spl_101,
    G12_n_spl_10
  );


  buf

  (
    G12_n_spl_11,
    G12_n_spl_1
  );


  buf

  (
    G12_n_spl_110,
    G12_n_spl_11
  );


  buf

  (
    G12_n_spl_111,
    G12_n_spl_11
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_00,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_000,
    G12_p_spl_00
  );


  buf

  (
    G12_p_spl_0000,
    G12_p_spl_000
  );


  buf

  (
    G12_p_spl_0001,
    G12_p_spl_000
  );


  buf

  (
    G12_p_spl_001,
    G12_p_spl_00
  );


  buf

  (
    G12_p_spl_01,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_010,
    G12_p_spl_01
  );


  buf

  (
    G12_p_spl_011,
    G12_p_spl_01
  );


  buf

  (
    G12_p_spl_1,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_10,
    G12_p_spl_1
  );


  buf

  (
    G12_p_spl_100,
    G12_p_spl_10
  );


  buf

  (
    G12_p_spl_101,
    G12_p_spl_10
  );


  buf

  (
    G12_p_spl_11,
    G12_p_spl_1
  );


  buf

  (
    G12_p_spl_110,
    G12_p_spl_11
  );


  buf

  (
    G12_p_spl_111,
    G12_p_spl_11
  );


  buf

  (
    g222_n_spl_,
    g222_n
  );


  buf

  (
    g222_n_spl_0,
    g222_n_spl_
  );


  buf

  (
    g222_n_spl_1,
    g222_n_spl_
  );


  buf

  (
    g231_p_spl_,
    g231_p
  );


  buf

  (
    g231_p_spl_0,
    g231_p_spl_
  );


  buf

  (
    g231_p_spl_00,
    g231_p_spl_0
  );


  buf

  (
    g231_p_spl_01,
    g231_p_spl_0
  );


  buf

  (
    g231_p_spl_1,
    g231_p_spl_
  );


  buf

  (
    g213_p_spl_,
    g213_p
  );


  buf

  (
    g213_p_spl_0,
    g213_p_spl_
  );


  buf

  (
    g213_p_spl_00,
    g213_p_spl_0
  );


  buf

  (
    g213_p_spl_1,
    g213_p_spl_
  );


  buf

  (
    g213_n_spl_,
    g213_n
  );


  buf

  (
    g213_n_spl_0,
    g213_n_spl_
  );


  buf

  (
    g213_n_spl_1,
    g213_n_spl_
  );


  buf

  (
    G23_n_spl_,
    G23_n
  );


  buf

  (
    G23_n_spl_0,
    G23_n_spl_
  );


  buf

  (
    G23_n_spl_00,
    G23_n_spl_0
  );


  buf

  (
    G23_n_spl_000,
    G23_n_spl_00
  );


  buf

  (
    G23_n_spl_001,
    G23_n_spl_00
  );


  buf

  (
    G23_n_spl_01,
    G23_n_spl_0
  );


  buf

  (
    G23_n_spl_010,
    G23_n_spl_01
  );


  buf

  (
    G23_n_spl_011,
    G23_n_spl_01
  );


  buf

  (
    G23_n_spl_1,
    G23_n_spl_
  );


  buf

  (
    G23_n_spl_10,
    G23_n_spl_1
  );


  buf

  (
    G23_n_spl_100,
    G23_n_spl_10
  );


  buf

  (
    G23_n_spl_101,
    G23_n_spl_10
  );


  buf

  (
    G23_n_spl_11,
    G23_n_spl_1
  );


  buf

  (
    G23_n_spl_110,
    G23_n_spl_11
  );


  buf

  (
    G23_p_spl_,
    G23_p
  );


  buf

  (
    G23_p_spl_0,
    G23_p_spl_
  );


  buf

  (
    G23_p_spl_00,
    G23_p_spl_0
  );


  buf

  (
    G23_p_spl_000,
    G23_p_spl_00
  );


  buf

  (
    G23_p_spl_001,
    G23_p_spl_00
  );


  buf

  (
    G23_p_spl_01,
    G23_p_spl_0
  );


  buf

  (
    G23_p_spl_010,
    G23_p_spl_01
  );


  buf

  (
    G23_p_spl_011,
    G23_p_spl_01
  );


  buf

  (
    G23_p_spl_1,
    G23_p_spl_
  );


  buf

  (
    G23_p_spl_10,
    G23_p_spl_1
  );


  buf

  (
    G23_p_spl_100,
    G23_p_spl_10
  );


  buf

  (
    G23_p_spl_101,
    G23_p_spl_10
  );


  buf

  (
    G23_p_spl_11,
    G23_p_spl_1
  );


  buf

  (
    G23_p_spl_110,
    G23_p_spl_11
  );


  buf

  (
    g185_n_spl_,
    g185_n
  );


  buf

  (
    g185_n_spl_0,
    g185_n_spl_
  );


  buf

  (
    g185_n_spl_00,
    g185_n_spl_0
  );


  buf

  (
    g185_n_spl_1,
    g185_n_spl_
  );


  buf

  (
    g185_p_spl_,
    g185_p
  );


  buf

  (
    g185_p_spl_0,
    g185_p_spl_
  );


  buf

  (
    g185_p_spl_1,
    g185_p_spl_
  );


  buf

  (
    g203_n_spl_,
    g203_n
  );


  buf

  (
    g203_n_spl_0,
    g203_n_spl_
  );


  buf

  (
    g203_n_spl_00,
    g203_n_spl_0
  );


  buf

  (
    g203_n_spl_1,
    g203_n_spl_
  );


  buf

  (
    g203_p_spl_,
    g203_p
  );


  buf

  (
    g203_p_spl_0,
    g203_p_spl_
  );


  buf

  (
    g203_p_spl_1,
    g203_p_spl_
  );


  buf

  (
    g427_n_spl_,
    g427_n
  );


  buf

  (
    g427_n_spl_0,
    g427_n_spl_
  );


  buf

  (
    g427_n_spl_1,
    g427_n_spl_
  );


  buf

  (
    g427_p_spl_,
    g427_p
  );


  buf

  (
    g427_p_spl_0,
    g427_p_spl_
  );


  buf

  (
    g427_p_spl_1,
    g427_p_spl_
  );


  buf

  (
    g255_p_spl_,
    g255_p
  );


  buf

  (
    g255_p_spl_0,
    g255_p_spl_
  );


  buf

  (
    g255_p_spl_00,
    g255_p_spl_0
  );


  buf

  (
    g255_p_spl_1,
    g255_p_spl_
  );


  buf

  (
    g262_n_spl_,
    g262_n
  );


  buf

  (
    g262_n_spl_0,
    g262_n_spl_
  );


  buf

  (
    g262_n_spl_1,
    g262_n_spl_
  );


  buf

  (
    g262_p_spl_,
    g262_p
  );


  buf

  (
    g262_p_spl_0,
    g262_p_spl_
  );


  buf

  (
    g262_p_spl_1,
    g262_p_spl_
  );


  buf

  (
    g271_p_spl_,
    g271_p
  );


  buf

  (
    g271_p_spl_0,
    g271_p_spl_
  );


  buf

  (
    g271_p_spl_1,
    g271_p_spl_
  );


  buf

  (
    g271_n_spl_,
    g271_n
  );


  buf

  (
    g271_n_spl_0,
    g271_n_spl_
  );


  buf

  (
    g271_n_spl_1,
    g271_n_spl_
  );


  buf

  (
    g280_p_spl_,
    g280_p
  );


  buf

  (
    g280_p_spl_0,
    g280_p_spl_
  );


  buf

  (
    g280_p_spl_1,
    g280_p_spl_
  );


  buf

  (
    g280_n_spl_,
    g280_n
  );


  buf

  (
    g280_n_spl_0,
    g280_n_spl_
  );


  buf

  (
    g280_n_spl_00,
    g280_n_spl_0
  );


  buf

  (
    g280_n_spl_1,
    g280_n_spl_
  );


  buf

  (
    g484_n_spl_,
    g484_n
  );


  buf

  (
    g484_n_spl_0,
    g484_n_spl_
  );


  buf

  (
    g484_n_spl_1,
    g484_n_spl_
  );


  buf

  (
    g484_p_spl_,
    g484_p
  );


  buf

  (
    g484_p_spl_0,
    g484_p_spl_
  );


  buf

  (
    g484_p_spl_1,
    g484_p_spl_
  );


  buf

  (
    g503_n_spl_,
    g503_n
  );


  buf

  (
    g503_n_spl_0,
    g503_n_spl_
  );


  buf

  (
    g503_p_spl_,
    g503_p
  );


  buf

  (
    g503_p_spl_0,
    g503_p_spl_
  );


  buf

  (
    g194_n_spl_,
    g194_n
  );


  buf

  (
    g194_n_spl_0,
    g194_n_spl_
  );


  buf

  (
    g194_n_spl_1,
    g194_n_spl_
  );


  buf

  (
    g194_p_spl_,
    g194_p
  );


  buf

  (
    g194_p_spl_0,
    g194_p_spl_
  );


  buf

  (
    g522_n_spl_,
    g522_n
  );


  buf

  (
    g522_n_spl_0,
    g522_n_spl_
  );


  buf

  (
    g522_n_spl_1,
    g522_n_spl_
  );


  buf

  (
    g522_p_spl_,
    g522_p
  );


  buf

  (
    g522_p_spl_0,
    g522_p_spl_
  );


  buf

  (
    g522_p_spl_1,
    g522_p_spl_
  );


  buf

  (
    g550_n_spl_,
    g550_n
  );


  buf

  (
    g550_n_spl_0,
    g550_n_spl_
  );


  buf

  (
    g550_n_spl_1,
    g550_n_spl_
  );


  buf

  (
    g550_p_spl_,
    g550_p
  );


  buf

  (
    g553_n_spl_,
    g553_n
  );


  buf

  (
    g553_n_spl_0,
    g553_n_spl_
  );


  buf

  (
    g553_p_spl_,
    g553_p
  );


  buf

  (
    g553_p_spl_0,
    g553_p_spl_
  );


  buf

  (
    g562_p_spl_,
    g562_p
  );


  buf

  (
    g562_n_spl_,
    g562_n
  );


  buf

  (
    g574_p_spl_,
    g574_p
  );


  buf

  (
    g574_n_spl_,
    g574_n
  );


  buf

  (
    g577_p_spl_,
    g577_p
  );


  buf

  (
    g580_n_spl_,
    g580_n
  );


  buf

  (
    g577_n_spl_,
    g577_n
  );


  buf

  (
    g580_p_spl_,
    g580_p
  );


  buf

  (
    g583_n_spl_,
    g583_n
  );


  buf

  (
    g586_n_spl_,
    g586_n
  );


  buf

  (
    g583_p_spl_,
    g583_p
  );


  buf

  (
    g586_p_spl_,
    g586_p
  );


  buf

  (
    G29_n_spl_,
    G29_n
  );


  buf

  (
    g597_p_spl_,
    g597_p
  );


  buf

  (
    g600_n_spl_,
    g600_n
  );


  buf

  (
    g597_n_spl_,
    g597_n
  );


  buf

  (
    g600_p_spl_,
    g600_p
  );


  buf

  (
    g606_n_spl_,
    g606_n
  );


  buf

  (
    g606_p_spl_,
    g606_p
  );


  buf

  (
    g609_n_spl_,
    g609_n
  );


  buf

  (
    g609_n_spl_0,
    g609_n_spl_
  );


  buf

  (
    g609_n_spl_1,
    g609_n_spl_
  );


  buf

  (
    g298_n_spl_,
    g298_n
  );


  buf

  (
    g609_p_spl_,
    g609_p
  );


  buf

  (
    g609_p_spl_0,
    g609_p_spl_
  );


  buf

  (
    g609_p_spl_1,
    g609_p_spl_
  );


  buf

  (
    g603_p_spl_,
    g603_p
  );


  buf

  (
    g603_n_spl_,
    g603_n
  );


  buf

  (
    g620_p_spl_,
    g620_p
  );


  buf

  (
    g620_n_spl_,
    g620_n
  );


  buf

  (
    g628_p_spl_,
    g628_p
  );


  buf

  (
    g629_p_spl_,
    g629_p
  );


  buf

  (
    g628_n_spl_,
    g628_n
  );


  buf

  (
    g629_n_spl_,
    g629_n
  );


  buf

  (
    G8_n_spl_,
    G8_n
  );


  buf

  (
    g630_p_spl_,
    g630_p
  );


  buf

  (
    g630_p_spl_0,
    g630_p_spl_
  );


  buf

  (
    g630_p_spl_00,
    g630_p_spl_0
  );


  buf

  (
    g630_p_spl_01,
    g630_p_spl_0
  );


  buf

  (
    g630_p_spl_1,
    g630_p_spl_
  );


  buf

  (
    g631_n_spl_,
    g631_n
  );


  buf

  (
    g631_n_spl_0,
    g631_n_spl_
  );


  buf

  (
    g631_n_spl_1,
    g631_n_spl_
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    g630_n_spl_,
    g630_n
  );


  buf

  (
    g630_n_spl_0,
    g630_n_spl_
  );


  buf

  (
    g630_n_spl_00,
    g630_n_spl_0
  );


  buf

  (
    g630_n_spl_1,
    g630_n_spl_
  );


  buf

  (
    g633_p_spl_,
    g633_p
  );


  buf

  (
    g633_n_spl_,
    g633_n
  );


  buf

  (
    g637_p_spl_,
    g637_p
  );


  buf

  (
    g640_p_spl_,
    g640_p
  );


  buf

  (
    g643_p_spl_,
    g643_p
  );


  buf

  (
    g646_p_spl_,
    g646_p
  );


  buf

  (
    g651_n_spl_,
    g651_n
  );


  buf

  (
    g656_n_spl_,
    g656_n
  );


  buf

  (
    g661_n_spl_,
    g661_n
  );


  buf

  (
    g682_p_spl_,
    g682_p
  );


  buf

  (
    g682_p_spl_0,
    g682_p_spl_
  );


  buf

  (
    g682_p_spl_00,
    g682_p_spl_0
  );


  buf

  (
    g682_p_spl_01,
    g682_p_spl_0
  );


  buf

  (
    g682_p_spl_1,
    g682_p_spl_
  );


  buf

  (
    g682_p_spl_10,
    g682_p_spl_1
  );


  buf

  (
    g682_p_spl_11,
    g682_p_spl_1
  );


  buf

  (
    g682_n_spl_,
    g682_n
  );


  buf

  (
    g682_n_spl_0,
    g682_n_spl_
  );


  buf

  (
    g682_n_spl_00,
    g682_n_spl_0
  );


  buf

  (
    g682_n_spl_01,
    g682_n_spl_0
  );


  buf

  (
    g682_n_spl_1,
    g682_n_spl_
  );


  buf

  (
    g682_n_spl_10,
    g682_n_spl_1
  );


  buf

  (
    g682_n_spl_11,
    g682_n_spl_1
  );


  buf

  (
    g683_n_spl_,
    g683_n
  );


  buf

  (
    g684_p_spl_,
    g684_p
  );


  buf

  (
    g686_n_spl_,
    g686_n
  );


  buf

  (
    g687_p_spl_,
    g687_p
  );


  buf

  (
    g690_n_spl_,
    g690_n
  );


  buf

  (
    g694_n_spl_,
    g694_n
  );


  buf

  (
    g695_p_spl_,
    g695_p
  );


  buf

  (
    g699_p_spl_,
    g699_p
  );


  buf

  (
    g700_n_spl_,
    g700_n
  );


  buf

  (
    g698_n_spl_,
    g698_n
  );


  buf

  (
    g693_n_spl_,
    g693_n
  );


  buf

  (
    g342_p_spl_,
    g342_p
  );


  buf

  (
    g361_p_spl_,
    g361_p
  );


  buf

  (
    g388_p_spl_,
    g388_p
  );


  buf

  (
    g593_p_spl_,
    g593_p
  );


  buf

  (
    g627_p_spl_,
    g627_p
  );


  buf

  (
    G124_n_spl_,
    G124_n
  );


  buf

  (
    G137_n_spl_,
    G137_n
  );


  buf

  (
    G137_n_spl_0,
    G137_n_spl_
  );


  buf

  (
    g173_n_spl_,
    g173_n
  );


  buf

  (
    g292_n_spl_,
    g292_n
  );


  buf

  (
    g295_n_spl_,
    g295_n
  );


  buf

  (
    g301_n_spl_,
    g301_n
  );


  buf

  (
    g540_n_spl_,
    g540_n
  );


  buf

  (
    g617_p_spl_,
    g617_p
  );


  buf

  (
    g718_n_spl_,
    g718_n
  );


endmodule
