
module mymod
(
  G1_p,
  G1_n,
  G2_p,
  G2_n,
  G3_p,
  G3_n,
  G4_p,
  G4_n,
  G5_p,
  G5_n,
  G6_p,
  G6_n,
  G7_p,
  G7_n,
  G8_p,
  G8_n,
  G9_p,
  G9_n,
  G10_p,
  G10_n,
  G11_p,
  G11_n,
  G12_p,
  G12_n,
  G13_p,
  G13_n,
  G14_p,
  G14_n,
  G15_p,
  G15_n,
  G16_p,
  G16_n,
  G17_p,
  G17_n,
  G18_p,
  G18_n,
  G19_p,
  G19_n,
  G20_p,
  G20_n,
  G21_p,
  G21_n,
  G22_p,
  G22_n,
  G23_p,
  G23_n,
  G24_p,
  G24_n,
  G25_p,
  G25_n,
  G26_p,
  G26_n,
  G27_p,
  G27_n,
  G28_p,
  G28_n,
  G29_p,
  G29_n,
  G30_p,
  G30_n,
  G31_p,
  G31_n,
  G32_p,
  G32_n,
  G33_p,
  G33_n,
  G34_p,
  G34_n,
  G35_p,
  G35_n,
  G36_p,
  G36_n,
  G37_p,
  G37_n,
  G38_p,
  G38_n,
  G39_p,
  G39_n,
  G40_p,
  G40_n,
  G41_p,
  G41_n,
  G42_p,
  G42_n,
  G43_p,
  G43_n,
  G44_p,
  G44_n,
  G45_p,
  G45_n,
  G46_p,
  G46_n,
  G47_p,
  G47_n,
  G48_p,
  G48_n,
  G49_p,
  G49_n,
  G50_p,
  G50_n,
  G51_p,
  G51_n,
  G52_p,
  G52_n,
  G53_p,
  G53_n,
  G54_p,
  G54_n,
  G55_p,
  G55_n,
  G56_p,
  G56_n,
  G57_p,
  G57_n,
  G58_p,
  G58_n,
  G59_p,
  G59_n,
  G60_p,
  G60_n,
  G855_p,
  G856_p,
  G857_p,
  G858_p,
  G859_p,
  G860_n,
  G861_n,
  G862_n,
  G863_p,
  G864_n,
  G865_n,
  G866_p,
  G867_p,
  G868_p,
  G869_n,
  G870_p,
  G871_p,
  G872_p,
  G873_p,
  G874_p,
  G875_p,
  G876_p,
  G877_p,
  G878_p,
  G879_p,
  G880_p
);

  input G1_p;input G1_n;input G2_p;input G2_n;input G3_p;input G3_n;input G4_p;input G4_n;input G5_p;input G5_n;input G6_p;input G6_n;input G7_p;input G7_n;input G8_p;input G8_n;input G9_p;input G9_n;input G10_p;input G10_n;input G11_p;input G11_n;input G12_p;input G12_n;input G13_p;input G13_n;input G14_p;input G14_n;input G15_p;input G15_n;input G16_p;input G16_n;input G17_p;input G17_n;input G18_p;input G18_n;input G19_p;input G19_n;input G20_p;input G20_n;input G21_p;input G21_n;input G22_p;input G22_n;input G23_p;input G23_n;input G24_p;input G24_n;input G25_p;input G25_n;input G26_p;input G26_n;input G27_p;input G27_n;input G28_p;input G28_n;input G29_p;input G29_n;input G30_p;input G30_n;input G31_p;input G31_n;input G32_p;input G32_n;input G33_p;input G33_n;input G34_p;input G34_n;input G35_p;input G35_n;input G36_p;input G36_n;input G37_p;input G37_n;input G38_p;input G38_n;input G39_p;input G39_n;input G40_p;input G40_n;input G41_p;input G41_n;input G42_p;input G42_n;input G43_p;input G43_n;input G44_p;input G44_n;input G45_p;input G45_n;input G46_p;input G46_n;input G47_p;input G47_n;input G48_p;input G48_n;input G49_p;input G49_n;input G50_p;input G50_n;input G51_p;input G51_n;input G52_p;input G52_n;input G53_p;input G53_n;input G54_p;input G54_n;input G55_p;input G55_n;input G56_p;input G56_n;input G57_p;input G57_n;input G58_p;input G58_n;input G59_p;input G59_n;input G60_p;input G60_n;
  output G855_p;output G856_p;output G857_p;output G858_p;output G859_p;output G860_n;output G861_n;output G862_n;output G863_p;output G864_n;output G865_n;output G866_p;output G867_p;output G868_p;output G869_n;output G870_p;output G871_p;output G872_p;output G873_p;output G874_p;output G875_p;output G876_p;output G877_p;output G878_p;output G879_p;output G880_p;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire G51_p;
  wire G51_n;
  wire G52_p;
  wire G52_n;
  wire G53_p;
  wire G53_n;
  wire G54_p;
  wire G54_n;
  wire G55_p;
  wire G55_n;
  wire G56_p;
  wire G56_n;
  wire G57_p;
  wire G57_n;
  wire G58_p;
  wire G58_n;
  wire G59_p;
  wire G59_n;
  wire G60_p;
  wire G60_n;
  wire ffc_0_p;
  wire ffc_0_n;
  wire ffc_1_p;
  wire ffc_1_n;
  wire ffc_2_p;
  wire ffc_2_n;
  wire ffc_3_p;
  wire ffc_3_n;
  wire ffc_4_p;
  wire ffc_4_n;
  wire ffc_5_p;
  wire ffc_5_n;
  wire ffc_6_p;
  wire ffc_6_n;
  wire ffc_7_p;
  wire ffc_7_n;
  wire ffc_8_p;
  wire ffc_8_n;
  wire ffc_9_p;
  wire ffc_9_n;
  wire ffc_10_p;
  wire ffc_10_n;
  wire ffc_11_p;
  wire ffc_11_n;
  wire ffc_12_p;
  wire ffc_12_n;
  wire ffc_13_p;
  wire ffc_13_n;
  wire ffc_14_p;
  wire ffc_14_n;
  wire ffc_15_p;
  wire ffc_15_n;
  wire ffc_16_p;
  wire ffc_16_n;
  wire ffc_17_p;
  wire ffc_17_n;
  wire ffc_18_p;
  wire ffc_18_n;
  wire ffc_19_p;
  wire ffc_19_n;
  wire ffc_20_p;
  wire ffc_20_n;
  wire ffc_21_p;
  wire ffc_21_n;
  wire ffc_22_p;
  wire ffc_22_n;
  wire ffc_23_p;
  wire ffc_23_n;
  wire ffc_24_p;
  wire ffc_24_n;
  wire ffc_25_p;
  wire ffc_25_n;
  wire ffc_26_p;
  wire ffc_26_n;
  wire ffc_27_p;
  wire ffc_27_n;
  wire ffc_28_p;
  wire ffc_28_n;
  wire ffc_29_p;
  wire ffc_29_n;
  wire ffc_30_p;
  wire ffc_30_n;
  wire ffc_31_p;
  wire ffc_31_n;
  wire ffc_32_p;
  wire ffc_32_n;
  wire ffc_33_p;
  wire ffc_33_n;
  wire ffc_34_p;
  wire ffc_34_n;
  wire ffc_35_p;
  wire ffc_35_n;
  wire ffc_36_p;
  wire ffc_36_n;
  wire ffc_37_p;
  wire ffc_37_n;
  wire ffc_38_p;
  wire ffc_38_n;
  wire ffc_39_p;
  wire ffc_39_n;
  wire ffc_40_p;
  wire ffc_40_n;
  wire ffc_41_p;
  wire ffc_41_n;
  wire ffc_42_p;
  wire ffc_42_n;
  wire ffc_43_p;
  wire ffc_43_n;
  wire ffc_44_p;
  wire ffc_44_n;
  wire ffc_45_p;
  wire ffc_45_n;
  wire ffc_46_p;
  wire ffc_46_n;
  wire ffc_47_p;
  wire ffc_47_n;
  wire ffc_48_p;
  wire ffc_48_n;
  wire ffc_49_p;
  wire ffc_49_n;
  wire ffc_50_p;
  wire ffc_50_n;
  wire ffc_51_p;
  wire ffc_51_n;
  wire ffc_52_p;
  wire ffc_52_n;
  wire ffc_53_p;
  wire ffc_53_n;
  wire ffc_54_p;
  wire ffc_54_n;
  wire ffc_55_p;
  wire ffc_55_n;
  wire ffc_56_p;
  wire ffc_56_n;
  wire ffc_57_p;
  wire ffc_57_n;
  wire ffc_58_p;
  wire ffc_58_n;
  wire ffc_59_p;
  wire ffc_59_n;
  wire ffc_60_p;
  wire ffc_60_n;
  wire ffc_61_p;
  wire ffc_61_n;
  wire ffc_62_p;
  wire ffc_62_n;
  wire ffc_63_p;
  wire ffc_63_n;
  wire ffc_64_p;
  wire ffc_64_n;
  wire ffc_65_p;
  wire ffc_65_n;
  wire ffc_66_p;
  wire ffc_66_n;
  wire ffc_67_p;
  wire ffc_67_n;
  wire ffc_68_p;
  wire ffc_68_n;
  wire ffc_69_p;
  wire ffc_69_n;
  wire ffc_70_p;
  wire ffc_70_n;
  wire ffc_71_p;
  wire ffc_71_n;
  wire ffc_72_p;
  wire ffc_72_n;
  wire ffc_73_p;
  wire ffc_73_n;
  wire ffc_74_p;
  wire ffc_74_n;
  wire ffc_75_p;
  wire ffc_75_n;
  wire ffc_76_p;
  wire ffc_76_n;
  wire ffc_77_p;
  wire ffc_77_n;
  wire ffc_78_p;
  wire ffc_78_n;
  wire ffc_79_p;
  wire ffc_79_n;
  wire ffc_80_p;
  wire ffc_80_n;
  wire ffc_81_p;
  wire ffc_81_n;
  wire ffc_82_p;
  wire ffc_82_n;
  wire ffc_83_p;
  wire ffc_83_n;
  wire ffc_84_p;
  wire ffc_84_n;
  wire ffc_85_p;
  wire ffc_85_n;
  wire ffc_86_p;
  wire ffc_86_n;
  wire ffc_87_p;
  wire ffc_87_n;
  wire ffc_88_p;
  wire ffc_88_n;
  wire ffc_89_p;
  wire ffc_89_n;
  wire ffc_90_p;
  wire ffc_90_n;
  wire ffc_91_p;
  wire ffc_91_n;
  wire ffc_92_p;
  wire ffc_92_n;
  wire ffc_93_p;
  wire ffc_93_n;
  wire ffc_94_p;
  wire ffc_94_n;
  wire ffc_95_p;
  wire ffc_95_n;
  wire ffc_96_p;
  wire ffc_96_n;
  wire ffc_97_p;
  wire ffc_97_n;
  wire ffc_98_p;
  wire ffc_98_n;
  wire ffc_99_p;
  wire ffc_99_n;
  wire ffc_100_p;
  wire ffc_100_n;
  wire ffc_101_p;
  wire ffc_101_n;
  wire ffc_102_p;
  wire ffc_102_n;
  wire ffc_103_p;
  wire ffc_103_n;
  wire ffc_104_p;
  wire ffc_104_n;
  wire ffc_105_p;
  wire ffc_105_n;
  wire ffc_106_p;
  wire ffc_106_n;
  wire ffc_107_p;
  wire ffc_107_n;
  wire ffc_108_p;
  wire ffc_108_n;
  wire ffc_109_p;
  wire ffc_109_n;
  wire ffc_110_p;
  wire ffc_110_n;
  wire ffc_111_p;
  wire ffc_111_n;
  wire ffc_112_p;
  wire ffc_112_n;
  wire ffc_113_p;
  wire ffc_113_n;
  wire ffc_114_p;
  wire ffc_114_n;
  wire ffc_115_p;
  wire ffc_115_n;
  wire ffc_116_p;
  wire ffc_116_n;
  wire ffc_117_p;
  wire ffc_117_n;
  wire ffc_118_p;
  wire ffc_118_n;
  wire ffc_119_p;
  wire ffc_119_n;
  wire ffc_120_p;
  wire ffc_120_n;
  wire ffc_121_p;
  wire ffc_121_n;
  wire ffc_122_p;
  wire ffc_122_n;
  wire ffc_123_p;
  wire ffc_123_n;
  wire ffc_124_p;
  wire ffc_124_n;
  wire ffc_125_p;
  wire ffc_125_n;
  wire ffc_126_p;
  wire ffc_126_n;
  wire ffc_127_p;
  wire ffc_127_n;
  wire ffc_128_p;
  wire ffc_128_n;
  wire ffc_129_p;
  wire ffc_129_n;
  wire ffc_130_p;
  wire ffc_130_n;
  wire ffc_131_p;
  wire ffc_131_n;
  wire ffc_132_p;
  wire ffc_132_n;
  wire ffc_133_p;
  wire ffc_133_n;
  wire ffc_134_p;
  wire ffc_134_n;
  wire ffc_135_p;
  wire ffc_135_n;
  wire ffc_136_p;
  wire ffc_136_n;
  wire ffc_137_p;
  wire ffc_137_n;
  wire ffc_138_p;
  wire ffc_138_n;
  wire ffc_139_p;
  wire ffc_139_n;
  wire ffc_140_p;
  wire ffc_140_n;
  wire ffc_141_p;
  wire ffc_141_n;
  wire ffc_142_p;
  wire ffc_142_n;
  wire ffc_143_p;
  wire ffc_143_n;
  wire ffc_144_p;
  wire ffc_144_n;
  wire ffc_145_p;
  wire ffc_145_n;
  wire ffc_146_p;
  wire ffc_146_n;
  wire ffc_147_p;
  wire ffc_147_n;
  wire ffc_148_p;
  wire ffc_148_n;
  wire ffc_149_p;
  wire ffc_149_n;
  wire ffc_150_p;
  wire ffc_150_n;
  wire ffc_151_p;
  wire ffc_151_n;
  wire ffc_152_p;
  wire ffc_152_n;
  wire ffc_153_p;
  wire ffc_153_n;
  wire ffc_154_p;
  wire ffc_154_n;
  wire ffc_155_p;
  wire ffc_155_n;
  wire ffc_156_p;
  wire ffc_156_n;
  wire ffc_157_p;
  wire ffc_157_n;
  wire ffc_158_p;
  wire ffc_158_n;
  wire ffc_159_p;
  wire ffc_159_n;
  wire ffc_160_p;
  wire ffc_160_n;
  wire ffc_161_p;
  wire ffc_161_n;
  wire ffc_162_p;
  wire ffc_162_n;
  wire ffc_163_p;
  wire ffc_163_n;
  wire ffc_164_p;
  wire ffc_164_n;
  wire ffc_165_p;
  wire ffc_165_n;
  wire ffc_166_p;
  wire ffc_166_n;
  wire ffc_167_p;
  wire ffc_167_n;
  wire ffc_168_p;
  wire ffc_168_n;
  wire ffc_169_p;
  wire ffc_169_n;
  wire ffc_170_p;
  wire ffc_170_n;
  wire ffc_171_p;
  wire ffc_171_n;
  wire ffc_172_p;
  wire ffc_172_n;
  wire ffc_173_p;
  wire ffc_173_n;
  wire ffc_174_p;
  wire ffc_174_n;
  wire ffc_175_p;
  wire ffc_175_n;
  wire ffc_176_p;
  wire ffc_176_n;
  wire ffc_177_p;
  wire ffc_177_n;
  wire ffc_178_p;
  wire ffc_178_n;
  wire ffc_179_p;
  wire ffc_179_n;
  wire ffc_180_p;
  wire ffc_180_n;
  wire ffc_181_p;
  wire ffc_181_n;
  wire ffc_182_p;
  wire ffc_182_n;
  wire ffc_183_p;
  wire ffc_183_n;
  wire ffc_184_p;
  wire ffc_184_n;
  wire ffc_185_p;
  wire ffc_185_n;
  wire ffc_186_p;
  wire ffc_186_n;
  wire ffc_187_p;
  wire ffc_187_n;
  wire ffc_188_p;
  wire ffc_188_n;
  wire ffc_189_p;
  wire ffc_189_n;
  wire ffc_190_p;
  wire ffc_190_n;
  wire ffc_191_p;
  wire ffc_191_n;
  wire ffc_192_p;
  wire ffc_192_n;
  wire ffc_193_p;
  wire ffc_193_n;
  wire ffc_194_p;
  wire ffc_194_n;
  wire ffc_195_p;
  wire ffc_195_n;
  wire ffc_196_p;
  wire ffc_196_n;
  wire ffc_197_p;
  wire ffc_197_n;
  wire ffc_198_p;
  wire ffc_198_n;
  wire ffc_199_p;
  wire ffc_199_n;
  wire ffc_200_p;
  wire ffc_200_n;
  wire ffc_201_p;
  wire ffc_201_n;
  wire ffc_202_p;
  wire ffc_202_n;
  wire ffc_203_p;
  wire ffc_203_n;
  wire ffc_204_p;
  wire ffc_204_n;
  wire ffc_205_p;
  wire ffc_205_n;
  wire ffc_206_p;
  wire ffc_206_n;
  wire ffc_207_p;
  wire ffc_207_n;
  wire ffc_208_p;
  wire ffc_208_n;
  wire ffc_209_p;
  wire ffc_209_n;
  wire ffc_210_p;
  wire ffc_210_n;
  wire ffc_211_p;
  wire ffc_211_n;
  wire ffc_212_p;
  wire ffc_212_n;
  wire ffc_213_p;
  wire ffc_213_n;
  wire ffc_214_p;
  wire ffc_214_n;
  wire ffc_215_p;
  wire ffc_215_n;
  wire ffc_216_p;
  wire ffc_216_n;
  wire ffc_217_p;
  wire ffc_217_n;
  wire ffc_218_p;
  wire ffc_218_n;
  wire ffc_219_p;
  wire ffc_219_n;
  wire ffc_220_p;
  wire ffc_220_n;
  wire ffc_221_p;
  wire ffc_221_n;
  wire ffc_222_p;
  wire ffc_222_n;
  wire ffc_223_p;
  wire ffc_223_n;
  wire ffc_224_p;
  wire ffc_224_n;
  wire ffc_225_p;
  wire ffc_225_n;
  wire ffc_226_p;
  wire ffc_226_n;
  wire ffc_227_p;
  wire ffc_227_n;
  wire ffc_228_p;
  wire ffc_228_n;
  wire ffc_229_p;
  wire ffc_229_n;
  wire ffc_230_p;
  wire ffc_230_n;
  wire ffc_231_p;
  wire ffc_231_n;
  wire ffc_232_p;
  wire ffc_232_n;
  wire ffc_233_p;
  wire ffc_233_n;
  wire ffc_234_p;
  wire ffc_234_n;
  wire ffc_235_p;
  wire ffc_235_n;
  wire ffc_236_p;
  wire ffc_236_n;
  wire ffc_237_p;
  wire ffc_237_n;
  wire ffc_238_p;
  wire ffc_238_n;
  wire ffc_239_p;
  wire ffc_239_n;
  wire ffc_240_p;
  wire ffc_240_n;
  wire ffc_241_p;
  wire ffc_241_n;
  wire ffc_242_p;
  wire ffc_242_n;
  wire ffc_243_p;
  wire ffc_243_n;
  wire ffc_244_p;
  wire ffc_244_n;
  wire ffc_245_p;
  wire ffc_245_n;
  wire ffc_246_p;
  wire ffc_246_n;
  wire ffc_247_p;
  wire ffc_247_n;
  wire ffc_248_p;
  wire ffc_248_n;
  wire ffc_249_p;
  wire ffc_249_n;
  wire ffc_250_p;
  wire ffc_250_n;
  wire ffc_251_p;
  wire ffc_251_n;
  wire ffc_252_p;
  wire ffc_252_n;
  wire ffc_253_p;
  wire ffc_253_n;
  wire ffc_254_p;
  wire ffc_254_n;
  wire ffc_255_p;
  wire ffc_255_n;
  wire ffc_256_p;
  wire ffc_256_n;
  wire ffc_257_p;
  wire ffc_257_n;
  wire ffc_258_p;
  wire ffc_258_n;
  wire ffc_259_p;
  wire ffc_259_n;
  wire ffc_260_p;
  wire ffc_260_n;
  wire ffc_261_p;
  wire ffc_261_n;
  wire ffc_262_p;
  wire ffc_262_n;
  wire ffc_263_p;
  wire ffc_263_n;
  wire ffc_264_p;
  wire ffc_264_n;
  wire ffc_265_p;
  wire ffc_265_n;
  wire ffc_266_p;
  wire ffc_266_n;
  wire ffc_267_p;
  wire ffc_267_n;
  wire ffc_268_p;
  wire ffc_268_n;
  wire ffc_269_p;
  wire ffc_269_n;
  wire ffc_270_p;
  wire ffc_270_n;
  wire ffc_271_p;
  wire ffc_271_n;
  wire ffc_272_p;
  wire ffc_272_n;
  wire ffc_273_p;
  wire ffc_273_n;
  wire ffc_274_p;
  wire ffc_274_n;
  wire ffc_275_p;
  wire ffc_275_n;
  wire ffc_276_p;
  wire ffc_276_n;
  wire ffc_277_p;
  wire ffc_277_n;
  wire ffc_278_p;
  wire ffc_278_n;
  wire ffc_279_p;
  wire ffc_279_n;
  wire ffc_280_p;
  wire ffc_280_n;
  wire ffc_281_p;
  wire ffc_281_n;
  wire ffc_282_p;
  wire ffc_282_n;
  wire ffc_283_p;
  wire ffc_283_n;
  wire ffc_284_p;
  wire ffc_284_n;
  wire ffc_285_p;
  wire ffc_285_n;
  wire ffc_286_p;
  wire ffc_286_n;
  wire ffc_287_p;
  wire ffc_287_n;
  wire ffc_288_p;
  wire ffc_288_n;
  wire ffc_289_p;
  wire ffc_289_n;
  wire ffc_290_p;
  wire ffc_290_n;
  wire ffc_291_p;
  wire ffc_291_n;
  wire ffc_292_p;
  wire ffc_292_n;
  wire ffc_293_p;
  wire ffc_293_n;
  wire ffc_294_p;
  wire ffc_294_n;
  wire ffc_295_p;
  wire ffc_295_n;
  wire ffc_296_p;
  wire ffc_296_n;
  wire ffc_297_p;
  wire ffc_297_n;
  wire ffc_298_p;
  wire ffc_298_n;
  wire ffc_299_p;
  wire ffc_299_n;
  wire ffc_300_p;
  wire ffc_300_n;
  wire ffc_301_p;
  wire ffc_301_n;
  wire ffc_302_p;
  wire ffc_302_n;
  wire ffc_303_p;
  wire ffc_303_n;
  wire ffc_304_p;
  wire ffc_304_n;
  wire ffc_305_p;
  wire ffc_305_n;
  wire ffc_306_p;
  wire ffc_306_n;
  wire ffc_307_p;
  wire ffc_307_n;
  wire ffc_308_p;
  wire ffc_308_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire ffc_6_n_spl_;
  wire ffc_26_n_spl_;
  wire g370_n_spl_;
  wire ffc_10_n_spl_;
  wire ffc_10_n_spl_0;
  wire ffc_10_p_spl_;
  wire g375_n_spl_;
  wire g377_n_spl_;
  wire ffc_12_n_spl_;
  wire g379_n_spl_;
  wire g383_n_spl_;
  wire g373_n_spl_;
  wire ffc_237_n_spl_;
  wire ffc_259_n_spl_;
  wire ffc_261_n_spl_;
  wire ffc_259_p_spl_;
  wire ffc_261_p_spl_;
  wire ffc_77_p_spl_;
  wire ffc_77_p_spl_0;
  wire ffc_77_p_spl_1;
  wire g392_p_spl_;
  wire ffc_77_n_spl_;
  wire ffc_77_n_spl_0;
  wire ffc_77_n_spl_1;
  wire g392_n_spl_;
  wire ffc_262_n_spl_;
  wire ffc_263_n_spl_;
  wire ffc_262_p_spl_;
  wire ffc_263_p_spl_;
  wire ffc_81_p_spl_;
  wire g398_p_spl_;
  wire ffc_81_n_spl_;
  wire g398_n_spl_;
  wire ffc_264_n_spl_;
  wire ffc_265_n_spl_;
  wire ffc_264_p_spl_;
  wire ffc_265_p_spl_;
  wire g407_p_spl_;
  wire g407_n_spl_;
  wire ffc_267_n_spl_;
  wire ffc_269_n_spl_;
  wire ffc_267_p_spl_;
  wire ffc_269_p_spl_;
  wire ffc_119_p_spl_;
  wire g413_p_spl_;
  wire ffc_119_n_spl_;
  wire g413_n_spl_;
  wire ffc_135_n_spl_;
  wire ffc_135_n_spl_0;
  wire ffc_135_n_spl_00;
  wire ffc_135_n_spl_01;
  wire ffc_135_n_spl_1;
  wire ffc_135_n_spl_10;
  wire ffc_135_n_spl_11;
  wire ffc_127_n_spl_;
  wire ffc_127_n_spl_0;
  wire ffc_127_n_spl_00;
  wire ffc_127_n_spl_000;
  wire ffc_127_n_spl_001;
  wire ffc_127_n_spl_01;
  wire ffc_127_n_spl_010;
  wire ffc_127_n_spl_1;
  wire ffc_127_n_spl_10;
  wire ffc_127_n_spl_11;
  wire ffc_131_n_spl_;
  wire ffc_131_n_spl_0;
  wire ffc_131_n_spl_00;
  wire ffc_131_n_spl_01;
  wire ffc_131_n_spl_1;
  wire ffc_131_n_spl_10;
  wire ffc_131_n_spl_11;
  wire ffc_139_n_spl_;
  wire ffc_139_n_spl_0;
  wire ffc_139_n_spl_00;
  wire ffc_139_n_spl_01;
  wire ffc_139_n_spl_1;
  wire ffc_139_n_spl_10;
  wire ffc_139_n_spl_11;
  wire ffc_270_n_spl_;
  wire ffc_270_n_spl_0;
  wire ffc_270_n_spl_00;
  wire ffc_270_n_spl_01;
  wire ffc_270_n_spl_1;
  wire ffc_270_n_spl_10;
  wire ffc_270_n_spl_11;
  wire ffc_123_n_spl_;
  wire ffc_123_n_spl_0;
  wire ffc_123_n_spl_00;
  wire ffc_123_n_spl_01;
  wire ffc_123_n_spl_1;
  wire ffc_123_n_spl_10;
  wire ffc_143_n_spl_;
  wire ffc_171_n_spl_;
  wire g450_n_spl_;
  wire ffc_93_p_spl_;
  wire ffc_260_p_spl_;
  wire ffc_93_n_spl_;
  wire ffc_93_n_spl_0;
  wire ffc_260_n_spl_;
  wire ffc_260_n_spl_0;
  wire ffc_97_n_spl_;
  wire ffc_238_n_spl_;
  wire ffc_256_n_spl_;
  wire ffc_256_n_spl_0;
  wire ffc_266_n_spl_;
  wire ffc_256_p_spl_;
  wire ffc_266_p_spl_;
  wire g483_n_spl_;
  wire g483_p_spl_;
  wire g482_p_spl_;
  wire g485_n_spl_;
  wire g481_n_spl_;
  wire g481_n_spl_0;
  wire ffc_201_n_spl_;
  wire g488_n_spl_;
  wire g503_n_spl_;
  wire g518_n_spl_;
  wire ffc_235_n_spl_;
  wire g533_n_spl_;
  wire ffc_257_n_spl_;
  wire ffc_104_n_spl_;
  wire ffc_104_n_spl_0;
  wire g549_p_spl_;
  wire g549_p_spl_0;
  wire g548_n_spl_;
  wire g550_n_spl_;
  wire ffc_62_n_spl_;
  wire ffc_100_n_spl_;
  wire ffc_100_n_spl_0;
  wire g558_p_spl_;
  wire g558_p_spl_0;
  wire g551_p_spl_;
  wire g552_p_spl_;
  wire g553_n_spl_;
  wire ffc_287_n_spl_;
  wire g565_p_spl_;
  wire g565_p_spl_0;
  wire g563_n_spl_;
  wire g564_n_spl_;
  wire g559_n_spl_;
  wire ffc_58_p_spl_;
  wire ffc_58_p_spl_0;
  wire ffc_198_p_spl_;
  wire ffc_244_p_spl_;
  wire ffc_234_p_spl_;
  wire ffc_245_p_spl_;
  wire g566_p_spl_;
  wire g567_p_spl_;
  wire ffc_243_p_spl_;
  wire ffc_306_p_spl_;
  wire ffc_306_p_spl_0;
  wire ffc_306_p_spl_1;
  wire ffc_305_p_spl_;
  wire ffc_307_p_spl_;
  wire ffc_110_n_spl_;
  wire g582_p_spl_;
  wire g582_p_spl_0;
  wire g578_n_spl_;
  wire g583_n_spl_;
  wire ffc_298_p_spl_;
  wire ffc_303_p_spl_;
  wire g591_p_spl_;
  wire ffc_122_p_spl_;
  wire ffc_233_p_spl_;
  wire ffc_96_p_spl_;
  wire ffc_96_p_spl_0;
  wire g577_n_spl_;
  wire ffc_142_p_spl_;
  wire ffc_54_p_spl_;
  wire ffc_54_p_spl_0;
  wire ffc_180_p_spl_;
  wire ffc_62_p_spl_;
  wire ffc_254_p_spl_;
  wire ffc_209_p_spl_;
  wire ffc_200_p_spl_;
  wire ffc_92_p_spl_;
  wire ffc_100_p_spl_;
  wire ffc_104_p_spl_;
  wire g560_p_spl_;
  wire g562_p_spl_;
  wire g568_n_spl_;
  wire ffc_236_p_spl_;
  wire ffc_257_p_spl_;
  wire ffc_202_p_spl_;
  wire ffc_211_p_spl_;
  wire g571_n_spl_;
  wire ffc_68_p_spl_;
  wire ffc_252_p_spl_;
  wire ffc_252_p_spl_0;
  wire ffc_85_p_spl_;
  wire ffc_83_p_spl_;
  wire ffc_217_p_spl_;
  wire ffc_65_p_spl_;
  wire ffc_107_p_spl_;
  wire g644_n_spl_;
  wire g585_n_spl_;
  wire g587_n_spl_;
  wire g592_n_spl_;
  wire g593_p_spl_;
  wire g634_p_spl_;
  wire ffc_73_p_spl_;
  wire g599_n_spl_;
  wire g599_n_spl_0;
  wire ffc_299_p_spl_;
  wire g589_n_spl_;
  wire g589_n_spl_0;
  wire g601_p_spl_;
  wire g601_p_spl_0;
  wire ffc_71_p_spl_;
  wire ffc_87_p_spl_;
  wire ffc_114_p_spl_;
  wire g657_n_spl_;
  wire G2_p_spl_;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_1;
  wire g663_n_spl_;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire G11_p_spl_;
  wire g662_n_spl_;
  wire G6_p_spl_;
  wire G17_p_spl_;

  andX
  g_g370_p
  (
    .dout(g370_p),
    .din1(ffc_6_p),
    .din2(ffc_11_p)
  );


  orX
  g_g370_n
  (
    .dout(g370_n),
    .din1(ffc_6_n_spl_),
    .din2(ffc_11_n)
  );


  orX
  g_g371_n
  (
    .dout(g371_n),
    .din1(ffc_26_n_spl_),
    .din2(g370_n_spl_)
  );


  orX
  g_g372_n
  (
    .dout(g372_n),
    .din1(ffc_10_n_spl_0),
    .din2(ffc_159_n)
  );


  andX
  g_g373_p
  (
    .dout(g373_p),
    .din1(ffc_10_p_spl_),
    .din2(g370_p)
  );


  orX
  g_g373_n
  (
    .dout(g373_n),
    .din1(ffc_10_n_spl_0),
    .din2(g370_n_spl_)
  );


  orX
  g_g374_n
  (
    .dout(g374_n),
    .din1(ffc_31_n),
    .din2(ffc_35_n)
  );


  orX
  g_g375_n
  (
    .dout(g375_n),
    .din1(ffc_4_n),
    .din2(ffc_208_n)
  );


  orX
  g_g376_n
  (
    .dout(g376_n),
    .din1(ffc_0_n),
    .din2(g375_n_spl_)
  );


  orX
  g_g377_n
  (
    .dout(g377_n),
    .din1(ffc_5_n),
    .din2(g375_n_spl_)
  );


  orX
  g_g378_n
  (
    .dout(g378_n),
    .din1(g373_p),
    .din2(g377_n_spl_)
  );


  orX
  g_g379_n
  (
    .dout(g379_n),
    .din1(ffc_12_n_spl_),
    .din2(ffc_27_n)
  );


  orX
  g_g380_n
  (
    .dout(g380_n),
    .din1(ffc_26_n_spl_),
    .din2(g379_n_spl_)
  );


  orX
  g_g381_n
  (
    .dout(g381_n),
    .din1(ffc_10_n_spl_),
    .din2(g379_n_spl_)
  );


  andX
  g_g382_p
  (
    .dout(g382_p),
    .din1(ffc_10_p_spl_),
    .din2(ffc_160_p)
  );


  orX
  g_g383_n
  (
    .dout(g383_n),
    .din1(ffc_39_p),
    .din2(ffc_43_p)
  );


  andX
  g_g384_p
  (
    .dout(g384_p),
    .din1(ffc_51_p),
    .din2(g383_n_spl_)
  );


  orX
  g_g385_n
  (
    .dout(g385_n),
    .din1(g373_n_spl_),
    .din2(g377_n_spl_)
  );


  orX
  g_g386_n
  (
    .dout(g386_n),
    .din1(ffc_6_n_spl_),
    .din2(ffc_237_n_spl_)
  );


  orX
  g_g387_n
  (
    .dout(g387_n),
    .din1(ffc_12_n_spl_),
    .din2(ffc_25_n)
  );


  orX
  g_g388_n
  (
    .dout(g388_n),
    .din1(ffc_237_n_spl_),
    .din2(g387_n)
  );


  andX
  g_g389_p
  (
    .dout(g389_p),
    .din1(ffc_47_p),
    .din2(g383_n_spl_)
  );


  andX
  g_g390_p
  (
    .dout(g390_p),
    .din1(ffc_259_n_spl_),
    .din2(ffc_261_n_spl_)
  );


  orX
  g_g390_n
  (
    .dout(g390_n),
    .din1(ffc_259_p_spl_),
    .din2(ffc_261_p_spl_)
  );


  andX
  g_g391_p
  (
    .dout(g391_p),
    .din1(ffc_259_p_spl_),
    .din2(ffc_261_p_spl_)
  );


  orX
  g_g391_n
  (
    .dout(g391_n),
    .din1(ffc_259_n_spl_),
    .din2(ffc_261_n_spl_)
  );


  andX
  g_g392_p
  (
    .dout(g392_p),
    .din1(g390_n),
    .din2(g391_n)
  );


  orX
  g_g392_n
  (
    .dout(g392_n),
    .din1(g390_p),
    .din2(g391_p)
  );


  andX
  g_g393_p
  (
    .dout(g393_p),
    .din1(ffc_77_p_spl_0),
    .din2(g392_p_spl_)
  );


  orX
  g_g393_n
  (
    .dout(g393_n),
    .din1(ffc_77_n_spl_0),
    .din2(g392_n_spl_)
  );


  andX
  g_g394_p
  (
    .dout(g394_p),
    .din1(ffc_77_n_spl_0),
    .din2(g392_n_spl_)
  );


  orX
  g_g394_n
  (
    .dout(g394_n),
    .din1(ffc_77_p_spl_0),
    .din2(g392_p_spl_)
  );


  andX
  g_g395_p
  (
    .dout(g395_p),
    .din1(g393_n),
    .din2(g394_n)
  );


  orX
  g_g395_n
  (
    .dout(g395_n),
    .din1(g393_p),
    .din2(g394_p)
  );


  andX
  g_g396_p
  (
    .dout(g396_p),
    .din1(ffc_262_n_spl_),
    .din2(ffc_263_n_spl_)
  );


  orX
  g_g396_n
  (
    .dout(g396_n),
    .din1(ffc_262_p_spl_),
    .din2(ffc_263_p_spl_)
  );


  andX
  g_g397_p
  (
    .dout(g397_p),
    .din1(ffc_262_p_spl_),
    .din2(ffc_263_p_spl_)
  );


  orX
  g_g397_n
  (
    .dout(g397_n),
    .din1(ffc_262_n_spl_),
    .din2(ffc_263_n_spl_)
  );


  andX
  g_g398_p
  (
    .dout(g398_p),
    .din1(g396_n),
    .din2(g397_n)
  );


  orX
  g_g398_n
  (
    .dout(g398_n),
    .din1(g396_p),
    .din2(g397_p)
  );


  andX
  g_g399_p
  (
    .dout(g399_p),
    .din1(ffc_81_p_spl_),
    .din2(g398_p_spl_)
  );


  orX
  g_g399_n
  (
    .dout(g399_n),
    .din1(ffc_81_n_spl_),
    .din2(g398_n_spl_)
  );


  andX
  g_g400_p
  (
    .dout(g400_p),
    .din1(ffc_81_n_spl_),
    .din2(g398_n_spl_)
  );


  orX
  g_g400_n
  (
    .dout(g400_n),
    .din1(ffc_81_p_spl_),
    .din2(g398_p_spl_)
  );


  andX
  g_g401_p
  (
    .dout(g401_p),
    .din1(g399_n),
    .din2(g400_n)
  );


  orX
  g_g401_n
  (
    .dout(g401_n),
    .din1(g399_p),
    .din2(g400_p)
  );


  andX
  g_g402_p
  (
    .dout(g402_p),
    .din1(g395_n),
    .din2(g401_n)
  );


  andX
  g_g403_p
  (
    .dout(g403_p),
    .din1(g395_p),
    .din2(g401_p)
  );


  orX
  g_g404_n
  (
    .dout(g404_n),
    .din1(g402_p),
    .din2(g403_p)
  );


  andX
  g_g405_p
  (
    .dout(g405_p),
    .din1(ffc_264_n_spl_),
    .din2(ffc_265_n_spl_)
  );


  orX
  g_g405_n
  (
    .dout(g405_n),
    .din1(ffc_264_p_spl_),
    .din2(ffc_265_p_spl_)
  );


  andX
  g_g406_p
  (
    .dout(g406_p),
    .din1(ffc_264_p_spl_),
    .din2(ffc_265_p_spl_)
  );


  orX
  g_g406_n
  (
    .dout(g406_n),
    .din1(ffc_264_n_spl_),
    .din2(ffc_265_n_spl_)
  );


  andX
  g_g407_p
  (
    .dout(g407_p),
    .din1(g405_n),
    .din2(g406_n)
  );


  orX
  g_g407_n
  (
    .dout(g407_n),
    .din1(g405_p),
    .din2(g406_p)
  );


  andX
  g_g408_p
  (
    .dout(g408_p),
    .din1(ffc_77_p_spl_1),
    .din2(g407_p_spl_)
  );


  orX
  g_g408_n
  (
    .dout(g408_n),
    .din1(ffc_77_n_spl_1),
    .din2(g407_n_spl_)
  );


  andX
  g_g409_p
  (
    .dout(g409_p),
    .din1(ffc_77_n_spl_1),
    .din2(g407_n_spl_)
  );


  orX
  g_g409_n
  (
    .dout(g409_n),
    .din1(ffc_77_p_spl_1),
    .din2(g407_p_spl_)
  );


  andX
  g_g410_p
  (
    .dout(g410_p),
    .din1(g408_n),
    .din2(g409_n)
  );


  orX
  g_g410_n
  (
    .dout(g410_n),
    .din1(g408_p),
    .din2(g409_p)
  );


  andX
  g_g411_p
  (
    .dout(g411_p),
    .din1(ffc_267_n_spl_),
    .din2(ffc_269_n_spl_)
  );


  orX
  g_g411_n
  (
    .dout(g411_n),
    .din1(ffc_267_p_spl_),
    .din2(ffc_269_p_spl_)
  );


  andX
  g_g412_p
  (
    .dout(g412_p),
    .din1(ffc_267_p_spl_),
    .din2(ffc_269_p_spl_)
  );


  orX
  g_g412_n
  (
    .dout(g412_n),
    .din1(ffc_267_n_spl_),
    .din2(ffc_269_n_spl_)
  );


  andX
  g_g413_p
  (
    .dout(g413_p),
    .din1(g411_n),
    .din2(g412_n)
  );


  orX
  g_g413_n
  (
    .dout(g413_n),
    .din1(g411_p),
    .din2(g412_p)
  );


  andX
  g_g414_p
  (
    .dout(g414_p),
    .din1(ffc_119_p_spl_),
    .din2(g413_p_spl_)
  );


  orX
  g_g414_n
  (
    .dout(g414_n),
    .din1(ffc_119_n_spl_),
    .din2(g413_n_spl_)
  );


  andX
  g_g415_p
  (
    .dout(g415_p),
    .din1(ffc_119_n_spl_),
    .din2(g413_n_spl_)
  );


  orX
  g_g415_n
  (
    .dout(g415_n),
    .din1(ffc_119_p_spl_),
    .din2(g413_p_spl_)
  );


  andX
  g_g416_p
  (
    .dout(g416_p),
    .din1(g414_n),
    .din2(g415_n)
  );


  orX
  g_g416_n
  (
    .dout(g416_n),
    .din1(g414_p),
    .din2(g415_p)
  );


  andX
  g_g417_p
  (
    .dout(g417_p),
    .din1(g410_n),
    .din2(g416_n)
  );


  andX
  g_g418_p
  (
    .dout(g418_p),
    .din1(g410_p),
    .din2(g416_p)
  );


  orX
  g_g419_n
  (
    .dout(g419_n),
    .din1(g417_p),
    .din2(g418_p)
  );


  andX
  g_g420_p
  (
    .dout(g420_p),
    .din1(ffc_135_n_spl_00),
    .din2(ffc_163_p)
  );


  orX
  g_g421_n
  (
    .dout(g421_n),
    .din1(ffc_162_n),
    .din2(g420_p)
  );


  orX
  g_g422_n
  (
    .dout(g422_n),
    .din1(ffc_127_n_spl_000),
    .din2(ffc_152_n)
  );


  andX
  g_g423_p
  (
    .dout(g423_p),
    .din1(g421_n),
    .din2(g422_n)
  );


  orX
  g_g424_n
  (
    .dout(g424_n),
    .din1(ffc_127_n_spl_000),
    .din2(ffc_164_p)
  );


  andX
  g_g425_p
  (
    .dout(g425_p),
    .din1(ffc_131_n_spl_00),
    .din2(ffc_163_n)
  );


  andX
  g_g426_p
  (
    .dout(g426_p),
    .din1(g424_n),
    .din2(g425_p)
  );


  orX
  g_g427_n
  (
    .dout(g427_n),
    .din1(g423_p),
    .din2(g426_p)
  );


  orX
  g_g428_n
  (
    .dout(g428_n),
    .din1(ffc_139_n_spl_00),
    .din2(ffc_161_n)
  );


  orX
  g_g429_n
  (
    .dout(g429_n),
    .din1(ffc_115_n),
    .din2(ffc_270_n_spl_00)
  );


  orX
  g_g430_n
  (
    .dout(g430_n),
    .din1(ffc_72_n),
    .din2(ffc_123_n_spl_00)
  );


  orX
  g_g431_n
  (
    .dout(g431_n),
    .din1(ffc_143_n_spl_),
    .din2(ffc_156_n)
  );


  andX
  g_g432_p
  (
    .dout(g432_p),
    .din1(g430_n),
    .din2(g431_n)
  );


  andX
  g_g433_p
  (
    .dout(g433_p),
    .din1(g429_n),
    .din2(g432_p)
  );


  andX
  g_g434_p
  (
    .dout(g434_p),
    .din1(g428_n),
    .din2(g433_p)
  );


  andX
  g_g435_p
  (
    .dout(g435_p),
    .din1(g427_n),
    .din2(g434_p)
  );


  orX
  g_g436_n
  (
    .dout(g436_n),
    .din1(ffc_127_n_spl_001),
    .din2(ffc_185_n)
  );


  andX
  g_g437_p
  (
    .dout(g437_p),
    .din1(ffc_135_n_spl_00),
    .din2(ffc_191_p)
  );


  orX
  g_g438_n
  (
    .dout(g438_n),
    .din1(ffc_184_n),
    .din2(g437_p)
  );


  andX
  g_g439_p
  (
    .dout(g439_p),
    .din1(g436_n),
    .din2(g438_n)
  );


  orX
  g_g440_n
  (
    .dout(g440_n),
    .din1(ffc_127_n_spl_001),
    .din2(ffc_194_p)
  );


  andX
  g_g441_p
  (
    .dout(g441_p),
    .din1(ffc_131_n_spl_00),
    .din2(ffc_191_n)
  );


  andX
  g_g442_p
  (
    .dout(g442_p),
    .din1(g440_n),
    .din2(g441_p)
  );


  orX
  g_g443_n
  (
    .dout(g443_n),
    .din1(g439_p),
    .din2(g442_p)
  );


  orX
  g_g444_n
  (
    .dout(g444_n),
    .din1(ffc_139_n_spl_00),
    .din2(ffc_174_n)
  );


  orX
  g_g445_n
  (
    .dout(g445_n),
    .din1(ffc_66_n),
    .din2(ffc_123_n_spl_00)
  );


  orX
  g_g446_n
  (
    .dout(g446_n),
    .din1(ffc_108_n),
    .din2(ffc_270_n_spl_00)
  );


  andX
  g_g447_p
  (
    .dout(g447_p),
    .din1(g445_n),
    .din2(g446_n)
  );


  andX
  g_g448_p
  (
    .dout(g448_p),
    .din1(g444_n),
    .din2(g447_p)
  );


  andX
  g_g449_p
  (
    .dout(g449_p),
    .din1(g443_n),
    .din2(g448_p)
  );


  andX
  g_g450_p
  (
    .dout(g450_p),
    .din1(ffc_171_n_spl_),
    .din2(ffc_173_p)
  );


  orX
  g_g450_n
  (
    .dout(g450_n),
    .din1(ffc_171_p),
    .din2(ffc_173_n)
  );


  orX
  g_g451_n
  (
    .dout(g451_n),
    .din1(ffc_172_n),
    .din2(g450_p)
  );


  orX
  g_g452_n
  (
    .dout(g452_n),
    .din1(ffc_172_p),
    .din2(g450_n_spl_)
  );


  andX
  g_g453_p
  (
    .dout(g453_p),
    .din1(g451_n),
    .din2(g452_n)
  );


  orX
  g_g454_n
  (
    .dout(g454_n),
    .din1(ffc_127_n_spl_010),
    .din2(g453_p)
  );


  orX
  g_g455_n
  (
    .dout(g455_n),
    .din1(ffc_131_n_spl_01),
    .din2(g450_n_spl_)
  );


  orX
  g_g456_n
  (
    .dout(g456_n),
    .din1(ffc_135_n_spl_01),
    .din2(ffc_171_n_spl_)
  );


  orX
  g_g457_n
  (
    .dout(g457_n),
    .din1(ffc_139_n_spl_01),
    .din2(ffc_169_n)
  );


  orX
  g_g458_n
  (
    .dout(g458_n),
    .din1(ffc_111_n),
    .din2(ffc_270_n_spl_01)
  );


  andX
  g_g459_p
  (
    .dout(g459_p),
    .din1(ffc_255_n),
    .din2(ffc_258_n)
  );


  andX
  g_g460_p
  (
    .dout(g460_p),
    .din1(g458_n),
    .din2(g459_p)
  );


  andX
  g_g461_p
  (
    .dout(g461_p),
    .din1(g457_n),
    .din2(g460_p)
  );


  andX
  g_g462_p
  (
    .dout(g462_p),
    .din1(g456_n),
    .din2(g461_p)
  );


  andX
  g_g463_p
  (
    .dout(g463_p),
    .din1(g455_n),
    .din2(g462_p)
  );


  andX
  g_g464_p
  (
    .dout(g464_p),
    .din1(g454_n),
    .din2(g463_p)
  );


  andX
  g_g465_p
  (
    .dout(g465_p),
    .din1(ffc_135_n_spl_01),
    .din2(ffc_168_p)
  );


  orX
  g_g466_n
  (
    .dout(g466_n),
    .din1(ffc_166_n),
    .din2(g465_p)
  );


  orX
  g_g467_n
  (
    .dout(g467_n),
    .din1(ffc_127_n_spl_010),
    .din2(ffc_167_n)
  );


  andX
  g_g468_p
  (
    .dout(g468_p),
    .din1(g466_n),
    .din2(g467_n)
  );


  orX
  g_g469_n
  (
    .dout(g469_n),
    .din1(ffc_127_n_spl_01),
    .din2(ffc_170_p)
  );


  andX
  g_g470_p
  (
    .dout(g470_p),
    .din1(ffc_131_n_spl_01),
    .din2(ffc_168_n)
  );


  andX
  g_g471_p
  (
    .dout(g471_p),
    .din1(g469_n),
    .din2(g470_p)
  );


  orX
  g_g472_n
  (
    .dout(g472_n),
    .din1(g468_p),
    .din2(g471_p)
  );


  orX
  g_g473_n
  (
    .dout(g473_n),
    .din1(ffc_139_n_spl_01),
    .din2(ffc_165_n)
  );


  orX
  g_g474_n
  (
    .dout(g474_n),
    .din1(ffc_113_n),
    .din2(ffc_270_n_spl_01)
  );


  orX
  g_g475_n
  (
    .dout(g475_n),
    .din1(ffc_70_n),
    .din2(ffc_123_n_spl_01)
  );


  orX
  g_g476_n
  (
    .dout(g476_n),
    .din1(ffc_143_n_spl_),
    .din2(ffc_150_n)
  );


  andX
  g_g477_p
  (
    .dout(g477_p),
    .din1(g475_n),
    .din2(g476_n)
  );


  andX
  g_g478_p
  (
    .dout(g478_p),
    .din1(g474_n),
    .din2(g477_p)
  );


  andX
  g_g479_p
  (
    .dout(g479_p),
    .din1(g473_n),
    .din2(g478_p)
  );


  andX
  g_g480_p
  (
    .dout(g480_p),
    .din1(g472_n),
    .din2(g479_p)
  );


  andX
  g_g481_p
  (
    .dout(g481_p),
    .din1(ffc_93_p_spl_),
    .din2(ffc_260_p_spl_)
  );


  orX
  g_g481_n
  (
    .dout(g481_n),
    .din1(ffc_93_n_spl_0),
    .din2(ffc_260_n_spl_0)
  );


  andX
  g_g482_p
  (
    .dout(g482_p),
    .din1(ffc_93_n_spl_0),
    .din2(ffc_260_n_spl_0)
  );


  orX
  g_g482_n
  (
    .dout(g482_n),
    .din1(ffc_93_p_spl_),
    .din2(ffc_260_p_spl_)
  );


  andX
  g_g483_p
  (
    .dout(g483_p),
    .din1(ffc_97_n_spl_),
    .din2(ffc_238_n_spl_)
  );


  orX
  g_g483_n
  (
    .dout(g483_n),
    .din1(ffc_97_p),
    .din2(ffc_238_p)
  );


  andX
  g_g484_p
  (
    .dout(g484_p),
    .din1(ffc_256_n_spl_0),
    .din2(ffc_266_n_spl_)
  );


  orX
  g_g484_n
  (
    .dout(g484_n),
    .din1(ffc_256_p_spl_),
    .din2(ffc_266_p_spl_)
  );


  andX
  g_g485_p
  (
    .dout(g485_p),
    .din1(g483_n_spl_),
    .din2(g484_n)
  );


  orX
  g_g485_n
  (
    .dout(g485_n),
    .din1(g483_p_spl_),
    .din2(g484_p)
  );


  orX
  g_g486_n
  (
    .dout(g486_n),
    .din1(g482_p_spl_),
    .din2(g485_n_spl_)
  );


  andX
  g_g487_p
  (
    .dout(g487_p),
    .din1(g481_n_spl_0),
    .din2(g486_n)
  );


  andX
  g_g488_p
  (
    .dout(g488_p),
    .din1(ffc_196_p),
    .din2(ffc_201_n_spl_)
  );


  orX
  g_g488_n
  (
    .dout(g488_n),
    .din1(ffc_196_n),
    .din2(ffc_201_p)
  );


  orX
  g_g489_n
  (
    .dout(g489_n),
    .din1(ffc_197_n),
    .din2(g488_p)
  );


  orX
  g_g490_n
  (
    .dout(g490_n),
    .din1(ffc_197_p),
    .din2(g488_n_spl_)
  );


  andX
  g_g491_p
  (
    .dout(g491_p),
    .din1(g489_n),
    .din2(g490_n)
  );


  orX
  g_g492_n
  (
    .dout(g492_n),
    .din1(ffc_127_n_spl_10),
    .din2(g491_p)
  );


  orX
  g_g493_n
  (
    .dout(g493_n),
    .din1(ffc_131_n_spl_10),
    .din2(g488_n_spl_)
  );


  orX
  g_g494_n
  (
    .dout(g494_n),
    .din1(ffc_135_n_spl_10),
    .din2(ffc_201_n_spl_)
  );


  orX
  g_g495_n
  (
    .dout(g495_n),
    .din1(ffc_139_n_spl_10),
    .din2(ffc_193_n)
  );


  orX
  g_g496_n
  (
    .dout(g496_n),
    .din1(ffc_105_n),
    .din2(ffc_270_n_spl_10)
  );


  orX
  g_g497_n
  (
    .dout(g497_n),
    .din1(ffc_63_n),
    .din2(ffc_123_n_spl_01)
  );


  andX
  g_g498_p
  (
    .dout(g498_p),
    .din1(g496_n),
    .din2(g497_n)
  );


  andX
  g_g499_p
  (
    .dout(g499_p),
    .din1(g495_n),
    .din2(g498_p)
  );


  andX
  g_g500_p
  (
    .dout(g500_p),
    .din1(g494_n),
    .din2(g499_p)
  );


  andX
  g_g501_p
  (
    .dout(g501_p),
    .din1(g493_n),
    .din2(g500_p)
  );


  andX
  g_g502_p
  (
    .dout(g502_p),
    .din1(g492_n),
    .din2(g501_p)
  );


  andX
  g_g503_p
  (
    .dout(g503_p),
    .din1(g481_n_spl_0),
    .din2(g482_n)
  );


  orX
  g_g503_n
  (
    .dout(g503_n),
    .din1(g481_p),
    .din2(g482_p_spl_)
  );


  andX
  g_g504_p
  (
    .dout(g504_p),
    .din1(g485_p),
    .din2(g503_p)
  );


  andX
  g_g505_p
  (
    .dout(g505_p),
    .din1(g485_n_spl_),
    .din2(g503_n_spl_)
  );


  orX
  g_g506_n
  (
    .dout(g506_n),
    .din1(ffc_127_n_spl_10),
    .din2(g505_p)
  );


  orX
  g_g507_n
  (
    .dout(g507_n),
    .din1(g504_p),
    .din2(g506_n)
  );


  orX
  g_g508_n
  (
    .dout(g508_n),
    .din1(ffc_131_n_spl_10),
    .din2(g503_n_spl_)
  );


  orX
  g_g509_n
  (
    .dout(g509_n),
    .din1(ffc_135_n_spl_10),
    .din2(g481_n_spl_)
  );


  orX
  g_g510_n
  (
    .dout(g510_n),
    .din1(ffc_139_n_spl_10),
    .din2(ffc_260_n_spl_)
  );


  orX
  g_g511_n
  (
    .dout(g511_n),
    .din1(ffc_123_n_spl_10),
    .din2(ffc_157_n)
  );


  orX
  g_g512_n
  (
    .dout(g512_n),
    .din1(ffc_93_n_spl_),
    .din2(ffc_270_n_spl_10)
  );


  andX
  g_g513_p
  (
    .dout(g513_p),
    .din1(g511_n),
    .din2(g512_n)
  );


  andX
  g_g514_p
  (
    .dout(g514_p),
    .din1(g510_n),
    .din2(g513_p)
  );


  andX
  g_g515_p
  (
    .dout(g515_p),
    .din1(g509_n),
    .din2(g514_p)
  );


  andX
  g_g516_p
  (
    .dout(g516_p),
    .din1(g508_n),
    .din2(g515_p)
  );


  andX
  g_g517_p
  (
    .dout(g517_p),
    .din1(g507_n),
    .din2(g516_p)
  );


  andX
  g_g518_p
  (
    .dout(g518_p),
    .din1(ffc_256_n_spl_0),
    .din2(g483_n_spl_)
  );


  orX
  g_g518_n
  (
    .dout(g518_n),
    .din1(ffc_256_p_spl_),
    .din2(g483_p_spl_)
  );


  andX
  g_g519_p
  (
    .dout(g519_p),
    .din1(ffc_266_p_spl_),
    .din2(g518_p)
  );


  andX
  g_g520_p
  (
    .dout(g520_p),
    .din1(ffc_266_n_spl_),
    .din2(g518_n_spl_)
  );


  orX
  g_g521_n
  (
    .dout(g521_n),
    .din1(ffc_127_n_spl_11),
    .din2(g520_p)
  );


  orX
  g_g522_n
  (
    .dout(g522_n),
    .din1(g519_p),
    .din2(g521_n)
  );


  orX
  g_g523_n
  (
    .dout(g523_n),
    .din1(ffc_131_n_spl_11),
    .din2(g518_n_spl_)
  );


  orX
  g_g524_n
  (
    .dout(g524_n),
    .din1(ffc_135_n_spl_11),
    .din2(ffc_256_n_spl_)
  );


  orX
  g_g525_n
  (
    .dout(g525_n),
    .din1(ffc_139_n_spl_11),
    .din2(ffc_238_n_spl_)
  );


  orX
  g_g526_n
  (
    .dout(g526_n),
    .din1(ffc_55_n),
    .din2(ffc_123_n_spl_10)
  );


  orX
  g_g527_n
  (
    .dout(g527_n),
    .din1(ffc_97_n_spl_),
    .din2(ffc_270_n_spl_11)
  );


  andX
  g_g528_p
  (
    .dout(g528_p),
    .din1(g526_n),
    .din2(g527_n)
  );


  andX
  g_g529_p
  (
    .dout(g529_p),
    .din1(g525_n),
    .din2(g528_p)
  );


  andX
  g_g530_p
  (
    .dout(g530_p),
    .din1(g524_n),
    .din2(g529_p)
  );


  andX
  g_g531_p
  (
    .dout(g531_p),
    .din1(g523_n),
    .din2(g530_p)
  );


  andX
  g_g532_p
  (
    .dout(g532_p),
    .din1(g522_n),
    .din2(g531_p)
  );


  andX
  g_g533_p
  (
    .dout(g533_p),
    .din1(ffc_210_p),
    .din2(ffc_235_n_spl_)
  );


  orX
  g_g533_n
  (
    .dout(g533_n),
    .din1(ffc_210_n),
    .din2(ffc_235_p)
  );


  andX
  g_g534_p
  (
    .dout(g534_p),
    .din1(ffc_212_n),
    .din2(g533_n_spl_)
  );


  andX
  g_g535_p
  (
    .dout(g535_p),
    .din1(ffc_212_p),
    .din2(g533_p)
  );


  orX
  g_g536_n
  (
    .dout(g536_n),
    .din1(ffc_127_n_spl_11),
    .din2(g535_p)
  );


  orX
  g_g537_n
  (
    .dout(g537_n),
    .din1(g534_p),
    .din2(g536_n)
  );


  orX
  g_g538_n
  (
    .dout(g538_n),
    .din1(ffc_131_n_spl_11),
    .din2(g533_n_spl_)
  );


  orX
  g_g539_n
  (
    .dout(g539_n),
    .din1(ffc_135_n_spl_11),
    .din2(ffc_235_n_spl_)
  );


  orX
  g_g540_n
  (
    .dout(g540_n),
    .din1(ffc_139_n_spl_11),
    .din2(ffc_203_n)
  );


  orX
  g_g541_n
  (
    .dout(g541_n),
    .din1(ffc_59_n),
    .din2(ffc_123_n_spl_1)
  );


  orX
  g_g542_n
  (
    .dout(g542_n),
    .din1(ffc_101_n),
    .din2(ffc_270_n_spl_11)
  );


  andX
  g_g543_p
  (
    .dout(g543_p),
    .din1(g541_n),
    .din2(g542_n)
  );


  andX
  g_g544_p
  (
    .dout(g544_p),
    .din1(g540_n),
    .din2(g543_p)
  );


  andX
  g_g545_p
  (
    .dout(g545_p),
    .din1(g539_n),
    .din2(g544_p)
  );


  andX
  g_g546_p
  (
    .dout(g546_p),
    .din1(g538_n),
    .din2(g545_p)
  );


  andX
  g_g547_p
  (
    .dout(g547_p),
    .din1(g537_n),
    .din2(g546_p)
  );


  orX
  g_g548_n
  (
    .dout(g548_n),
    .din1(ffc_257_n_spl_),
    .din2(ffc_271_n)
  );


  andX
  g_g549_p
  (
    .dout(g549_p),
    .din1(ffc_274_n),
    .din2(ffc_278_n)
  );


  orX
  g_g550_n
  (
    .dout(g550_n),
    .din1(ffc_276_n),
    .din2(ffc_279_n)
  );


  andX
  g_g551_p
  (
    .dout(g551_p),
    .din1(ffc_104_n_spl_0),
    .din2(g549_p_spl_0)
  );


  andX
  g_g552_p
  (
    .dout(g552_p),
    .din1(g548_n_spl_),
    .din2(g550_n_spl_)
  );


  orX
  g_g553_n
  (
    .dout(g553_n),
    .din1(ffc_104_n_spl_0),
    .din2(g549_p_spl_0)
  );


  orX
  g_g554_n
  (
    .dout(g554_n),
    .din1(ffc_62_n_spl_),
    .din2(ffc_198_n)
  );


  orX
  g_g555_n
  (
    .dout(g555_n),
    .din1(ffc_199_n),
    .din2(ffc_244_n)
  );


  andX
  g_g556_p
  (
    .dout(g556_p),
    .din1(ffc_245_n),
    .din2(ffc_273_n)
  );


  andX
  g_g557_p
  (
    .dout(g557_p),
    .din1(g555_n),
    .din2(g556_p)
  );


  andX
  g_g558_p
  (
    .dout(g558_p),
    .din1(g554_n),
    .din2(g557_p)
  );


  orX
  g_g559_n
  (
    .dout(g559_n),
    .din1(ffc_3_n),
    .din2(ffc_175_n)
  );


  andX
  g_g560_p
  (
    .dout(g560_p),
    .din1(ffc_100_n_spl_0),
    .din2(g558_p_spl_0)
  );


  orX
  g_g561_n
  (
    .dout(g561_n),
    .din1(g551_p_spl_),
    .din2(g552_p_spl_)
  );


  andX
  g_g562_p
  (
    .dout(g562_p),
    .din1(g553_n_spl_),
    .din2(g561_n)
  );


  orX
  g_g563_n
  (
    .dout(g563_n),
    .din1(ffc_277_n),
    .din2(ffc_280_n)
  );


  orX
  g_g564_n
  (
    .dout(g564_n),
    .din1(ffc_291_n),
    .din2(ffc_296_n)
  );


  andX
  g_g565_p
  (
    .dout(g565_p),
    .din1(ffc_288_n),
    .din2(ffc_289_n)
  );


  andX
  g_g566_p
  (
    .dout(g566_p),
    .din1(ffc_287_n_spl_),
    .din2(g565_p_spl_0)
  );


  andX
  g_g567_p
  (
    .dout(g567_p),
    .din1(g563_n_spl_),
    .din2(g564_n_spl_)
  );


  orX
  g_g568_n
  (
    .dout(g568_n),
    .din1(ffc_100_n_spl_0),
    .din2(g558_p_spl_0)
  );


  orX
  g_g569_n
  (
    .dout(g569_n),
    .din1(ffc_180_n),
    .din2(ffc_190_n)
  );


  orX
  g_g570_n
  (
    .dout(g570_n),
    .din1(ffc_15_n),
    .din2(g569_n)
  );


  orX
  g_g571_n
  (
    .dout(g571_n),
    .din1(g559_n_spl_),
    .din2(g570_n)
  );


  andX
  g_g572_p
  (
    .dout(g572_p),
    .din1(ffc_58_p_spl_0),
    .din2(ffc_198_p_spl_)
  );


  andX
  g_g573_p
  (
    .dout(g573_p),
    .din1(ffc_205_p),
    .din2(ffc_244_p_spl_)
  );


  andX
  g_g574_p
  (
    .dout(g574_p),
    .din1(ffc_178_p),
    .din2(ffc_234_p_spl_)
  );


  orX
  g_g575_n
  (
    .dout(g575_n),
    .din1(ffc_245_p_spl_),
    .din2(g574_p)
  );


  orX
  g_g576_n
  (
    .dout(g576_n),
    .din1(g573_p),
    .din2(g575_n)
  );


  orX
  g_g577_n
  (
    .dout(g577_n),
    .din1(g572_p),
    .din2(g576_n)
  );


  orX
  g_g578_n
  (
    .dout(g578_n),
    .din1(ffc_287_n_spl_),
    .din2(g565_p_spl_0)
  );


  orX
  g_g579_n
  (
    .dout(g579_n),
    .din1(ffc_252_n),
    .din2(ffc_286_n)
  );


  orX
  g_g580_n
  (
    .dout(g580_n),
    .din1(ffc_246_p),
    .din2(ffc_290_n)
  );


  andX
  g_g581_p
  (
    .dout(g581_p),
    .din1(ffc_253_n),
    .din2(g580_n)
  );


  andX
  g_g582_p
  (
    .dout(g582_p),
    .din1(g579_n),
    .din2(g581_p)
  );


  orX
  g_g583_n
  (
    .dout(g583_n),
    .din1(g566_p_spl_),
    .din2(g567_p_spl_)
  );


  orX
  g_g584_n
  (
    .dout(g584_n),
    .din1(ffc_228_p),
    .din2(ffc_242_n)
  );


  orX
  g_g585_n
  (
    .dout(g585_n),
    .din1(ffc_231_n),
    .din2(g584_n)
  );


  orX
  g_g586_n
  (
    .dout(g586_n),
    .din1(ffc_217_n),
    .din2(ffc_243_p_spl_)
  );


  orX
  g_g587_n
  (
    .dout(g587_n),
    .din1(ffc_247_n),
    .din2(g586_n)
  );


  andX
  g_g588_p
  (
    .dout(g588_p),
    .din1(ffc_301_p),
    .din2(ffc_306_p_spl_0)
  );


  orX
  g_g589_n
  (
    .dout(g589_n),
    .din1(ffc_281_n),
    .din2(g588_p)
  );


  andX
  g_g590_p
  (
    .dout(g590_p),
    .din1(ffc_305_p_spl_),
    .din2(ffc_307_p_spl_)
  );


  andX
  g_g591_p
  (
    .dout(g591_p),
    .din1(ffc_306_p_spl_0),
    .din2(g590_p)
  );


  orX
  g_g592_n
  (
    .dout(g592_n),
    .din1(ffc_110_n_spl_),
    .din2(g582_p_spl_0)
  );


  andX
  g_g593_p
  (
    .dout(g593_p),
    .din1(g578_n_spl_),
    .din2(g583_n_spl_)
  );


  andX
  g_g594_p
  (
    .dout(g594_p),
    .din1(ffc_298_p_spl_),
    .din2(ffc_308_p)
  );


  andX
  g_g595_p
  (
    .dout(g595_p),
    .din1(ffc_306_p_spl_1),
    .din2(g594_p)
  );


  orX
  g_g596_n
  (
    .dout(g596_n),
    .din1(ffc_302_n),
    .din2(ffc_305_n)
  );


  andX
  g_g597_p
  (
    .dout(g597_p),
    .din1(ffc_297_p),
    .din2(ffc_300_p)
  );


  andX
  g_g598_p
  (
    .dout(g598_p),
    .din1(g596_n),
    .din2(g597_p)
  );


  orX
  g_g599_n
  (
    .dout(g599_n),
    .din1(g595_p),
    .din2(g598_p)
  );


  andX
  g_g600_p
  (
    .dout(g600_p),
    .din1(ffc_303_p_spl_),
    .din2(ffc_304_n)
  );


  andX
  g_g601_p
  (
    .dout(g601_p),
    .din1(g591_p_spl_),
    .din2(g600_p)
  );


  andX
  g_g602_p
  (
    .dout(g602_p),
    .din1(ffc_122_p_spl_),
    .din2(ffc_233_p_spl_)
  );


  andX
  g_g603_p
  (
    .dout(g603_p),
    .din1(ffc_96_p_spl_0),
    .din2(g577_n_spl_)
  );


  andX
  g_g604_p
  (
    .dout(g604_p),
    .din1(ffc_142_p_spl_),
    .din2(ffc_146_p)
  );


  orX
  g_g605_n
  (
    .dout(g605_n),
    .din1(ffc_54_p_spl_0),
    .din2(ffc_58_p_spl_0)
  );


  orX
  g_g606_n
  (
    .dout(g606_n),
    .din1(ffc_54_n),
    .din2(ffc_58_n)
  );


  andX
  g_g607_p
  (
    .dout(g607_p),
    .din1(g605_n),
    .din2(g606_n)
  );


  andX
  g_g608_p
  (
    .dout(g608_p),
    .din1(ffc_54_p_spl_0),
    .din2(ffc_198_p_spl_)
  );


  andX
  g_g609_p
  (
    .dout(g609_p),
    .din1(ffc_180_p_spl_),
    .din2(ffc_234_p_spl_)
  );


  orX
  g_g610_n
  (
    .dout(g610_n),
    .din1(ffc_245_p_spl_),
    .din2(g609_p)
  );


  andX
  g_g611_p
  (
    .dout(g611_p),
    .din1(ffc_221_p),
    .din2(ffc_244_p_spl_)
  );


  orX
  g_g612_n
  (
    .dout(g612_n),
    .din1(g610_n),
    .din2(g611_p)
  );


  orX
  g_g613_n
  (
    .dout(g613_n),
    .din1(g608_p),
    .din2(g612_n)
  );


  orX
  g_g614_n
  (
    .dout(g614_n),
    .din1(ffc_62_p_spl_),
    .din2(ffc_254_p_spl_)
  );


  orX
  g_g615_n
  (
    .dout(g615_n),
    .din1(ffc_62_n_spl_),
    .din2(ffc_254_n)
  );


  andX
  g_g616_p
  (
    .dout(g616_p),
    .din1(g614_n),
    .din2(g615_n)
  );


  orX
  g_g617_n
  (
    .dout(g617_n),
    .din1(ffc_209_p_spl_),
    .din2(ffc_233_p_spl_)
  );


  orX
  g_g618_n
  (
    .dout(g618_n),
    .din1(ffc_209_n),
    .din2(ffc_233_n)
  );


  andX
  g_g619_p
  (
    .dout(g619_p),
    .din1(g617_n),
    .din2(g618_n)
  );


  orX
  g_g620_n
  (
    .dout(g620_n),
    .din1(ffc_195_p),
    .din2(ffc_200_p_spl_)
  );


  orX
  g_g621_n
  (
    .dout(g621_n),
    .din1(ffc_195_n),
    .din2(ffc_200_n)
  );


  andX
  g_g622_p
  (
    .dout(g622_p),
    .din1(g620_n),
    .din2(g621_n)
  );


  orX
  g_g623_n
  (
    .dout(g623_n),
    .din1(ffc_92_p_spl_),
    .din2(ffc_96_p_spl_0)
  );


  orX
  g_g624_n
  (
    .dout(g624_n),
    .din1(ffc_92_n),
    .din2(ffc_96_n)
  );


  andX
  g_g625_p
  (
    .dout(g625_p),
    .din1(g623_n),
    .din2(g624_n)
  );


  orX
  g_g626_n
  (
    .dout(g626_n),
    .din1(ffc_100_p_spl_),
    .din2(ffc_104_p_spl_)
  );


  orX
  g_g627_n
  (
    .dout(g627_n),
    .din1(ffc_100_n_spl_),
    .din2(ffc_104_n_spl_)
  );


  andX
  g_g628_p
  (
    .dout(g628_p),
    .din1(g626_n),
    .din2(g627_n)
  );


  orX
  g_g629_n
  (
    .dout(g629_n),
    .din1(g560_p_spl_),
    .din2(g562_p_spl_)
  );


  andX
  g_g630_p
  (
    .dout(g630_p),
    .din1(g568_n_spl_),
    .din2(g629_n)
  );


  orX
  g_g631_n
  (
    .dout(g631_n),
    .din1(ffc_236_p_spl_),
    .din2(ffc_257_p_spl_)
  );


  orX
  g_g632_n
  (
    .dout(g632_n),
    .din1(ffc_236_n),
    .din2(ffc_257_n_spl_)
  );


  andX
  g_g633_p
  (
    .dout(g633_p),
    .din1(g631_n),
    .din2(g632_n)
  );


  andX
  g_g634_p
  (
    .dout(g634_p),
    .din1(ffc_110_n_spl_),
    .din2(g582_p_spl_0)
  );


  orX
  g_g635_n
  (
    .dout(g635_n),
    .din1(ffc_202_p_spl_),
    .din2(ffc_211_p_spl_)
  );


  orX
  g_g636_n
  (
    .dout(g636_n),
    .din1(ffc_202_n),
    .din2(ffc_211_n)
  );


  andX
  g_g637_p
  (
    .dout(g637_p),
    .din1(g635_n),
    .din2(g636_n)
  );


  orX
  g_g638_n
  (
    .dout(g638_n),
    .din1(ffc_18_n),
    .din2(ffc_21_n)
  );


  orX
  g_g639_n
  (
    .dout(g639_n),
    .din1(ffc_187_n),
    .din2(g638_n)
  );


  orX
  g_g640_n
  (
    .dout(g640_n),
    .din1(g571_n_spl_),
    .din2(g639_n)
  );


  andX
  g_g641_p
  (
    .dout(g641_p),
    .din1(ffc_68_p_spl_),
    .din2(ffc_252_p_spl_0)
  );


  andX
  g_g642_p
  (
    .dout(g642_p),
    .din1(ffc_85_p_spl_),
    .din2(ffc_246_n)
  );


  orX
  g_g643_n
  (
    .dout(g643_n),
    .din1(ffc_253_p),
    .din2(g642_p)
  );


  orX
  g_g644_n
  (
    .dout(g644_n),
    .din1(g641_p),
    .din2(g643_n)
  );


  andX
  g_g645_p
  (
    .dout(g645_p),
    .din1(ffc_83_p_spl_),
    .din2(ffc_217_p_spl_)
  );


  andX
  g_g646_p
  (
    .dout(g646_p),
    .din1(ffc_65_p_spl_),
    .din2(ffc_252_p_spl_0)
  );


  orX
  g_g647_n
  (
    .dout(g647_n),
    .din1(ffc_107_p_spl_),
    .din2(g644_n_spl_)
  );


  orX
  g_g648_n
  (
    .dout(g648_n),
    .din1(ffc_248_n),
    .din2(g585_n_spl_)
  );


  orX
  g_g649_n
  (
    .dout(g649_n),
    .din1(ffc_83_n),
    .din2(ffc_89_n)
  );


  andX
  g_g650_p
  (
    .dout(g650_p),
    .din1(g587_n_spl_),
    .din2(g649_n)
  );


  andX
  g_g651_p
  (
    .dout(g651_p),
    .din1(g648_n),
    .din2(g650_p)
  );


  andX
  g_g652_p
  (
    .dout(g652_p),
    .din1(g592_n_spl_),
    .din2(g593_p_spl_)
  );


  orX
  g_g653_n
  (
    .dout(g653_n),
    .din1(g634_p_spl_),
    .din2(g652_p)
  );


  andX
  g_g654_p
  (
    .dout(g654_p),
    .din1(ffc_73_p_spl_),
    .din2(g599_n_spl_0)
  );


  andX
  g_g655_p
  (
    .dout(g655_p),
    .din1(ffc_299_p_spl_),
    .din2(g589_n_spl_0)
  );


  orX
  g_g656_n
  (
    .dout(g656_n),
    .din1(g601_p_spl_0),
    .din2(g655_p)
  );


  orX
  g_g657_n
  (
    .dout(g657_n),
    .din1(g654_p),
    .din2(g656_n)
  );


  andX
  g_g658_p
  (
    .dout(g658_p),
    .din1(ffc_71_p_spl_),
    .din2(g599_n_spl_0)
  );


  andX
  g_g659_p
  (
    .dout(g659_p),
    .din1(ffc_87_p_spl_),
    .din2(g589_n_spl_0)
  );


  orX
  g_g660_n
  (
    .dout(g660_n),
    .din1(g601_p_spl_0),
    .din2(g659_p)
  );


  orX
  g_g661_n
  (
    .dout(g661_n),
    .din1(ffc_114_p_spl_),
    .din2(g657_n_spl_)
  );


  orX
  g_g662_n
  (
    .dout(g662_n),
    .din1(G1_n),
    .din2(G9_n)
  );


  orX
  g_g663_n
  (
    .dout(g663_n),
    .din1(G11_n),
    .din2(G40_n)
  );


  andX
  g_g664_p
  (
    .dout(g664_p),
    .din1(G2_p_spl_),
    .din2(G4_p_spl_0)
  );


  andX
  g_g665_p
  (
    .dout(g665_p),
    .din1(G4_p_spl_0),
    .din2(g663_n_spl_)
  );


  andX
  g_g666_p
  (
    .dout(g666_p),
    .din1(G8_p_spl_0),
    .din2(G11_p_spl_)
  );


  orX
  g_g667_n
  (
    .dout(g667_n),
    .din1(G5_n),
    .din2(g662_n_spl_)
  );


  andX
  g_g668_p
  (
    .dout(g668_p),
    .din1(G6_p_spl_),
    .din2(G17_p_spl_)
  );


  andX
  g_g669_p
  (
    .dout(g669_p),
    .din1(G4_p_spl_1),
    .din2(G8_n)
  );


  andX
  g_g670_p
  (
    .dout(g670_p),
    .din1(G4_n),
    .din2(G8_p_spl_0)
  );


  orX
  g_g671_n
  (
    .dout(g671_n),
    .din1(g669_p),
    .din2(g670_p)
  );


  buf

  (
    G855_p,
    g371_n
  );


  buf

  (
    G856_p,
    g372_n
  );


  buf

  (
    G857_p,
    g373_n_spl_
  );


  buf

  (
    G858_p,
    g374_n
  );


  buf

  (
    G859_p,
    g376_n
  );


  buf

  (
    G860_n,
    g378_n
  );


  buf

  (
    G861_n,
    g380_n
  );


  buf

  (
    G862_n,
    g381_n
  );


  buf

  (
    G863_p,
    g382_p
  );


  buf

  (
    G864_n,
    g384_p
  );


  buf

  (
    G865_n,
    g385_n
  );


  buf

  (
    G866_p,
    ffc_158_n
  );


  buf

  (
    G867_p,
    g386_n
  );


  buf

  (
    G868_p,
    g388_n
  );


  buf

  (
    G869_n,
    g389_p
  );


  buf

  (
    G870_p,
    g404_n
  );


  buf

  (
    G871_p,
    g419_n
  );


  buf

  (
    G872_p,
    g435_p
  );


  buf

  (
    G873_p,
    g449_p
  );


  buf

  (
    G874_p,
    g464_p
  );


  buf

  (
    G875_p,
    g480_p
  );


  buf

  (
    G876_p,
    g487_p
  );


  buf

  (
    G877_p,
    g502_p
  );


  buf

  (
    G878_p,
    g517_p
  );


  buf

  (
    G879_p,
    g532_p
  );


  buf

  (
    G880_p,
    g547_p
  );


  DROC
  ffc_0
  (
    .doutp(ffc_0_p),
    .doutn(ffc_0_n),
    .din(ffc_180_p_spl_)
  );


  DROC
  ffc_1
  (
    .doutp(ffc_1_p),
    .doutn(ffc_1_n),
    .din(G3_p)
  );


  DROC
  ffc_2
  (
    .doutp(ffc_2_p),
    .doutn(ffc_2_n),
    .din(ffc_1_p)
  );


  DROC
  ffc_3
  (
    .doutp(ffc_3_p),
    .doutn(ffc_3_n),
    .din(ffc_2_p)
  );


  DROC
  ffc_4
  (
    .doutp(ffc_4_p),
    .doutn(ffc_4_n),
    .din(ffc_176_p)
  );


  DROC
  ffc_5
  (
    .doutp(ffc_5_p),
    .doutn(ffc_5_n),
    .din(ffc_181_p)
  );


  DROC
  ffc_6
  (
    .doutp(ffc_6_p),
    .doutn(ffc_6_n),
    .din(ffc_182_p)
  );


  DROC
  ffc_7
  (
    .doutp(ffc_7_p),
    .doutn(ffc_7_n),
    .din(G7_p)
  );


  DROC
  ffc_8
  (
    .doutp(ffc_8_p),
    .doutn(ffc_8_n),
    .din(ffc_7_p)
  );


  DROC
  ffc_9
  (
    .doutp(ffc_9_p),
    .doutn(ffc_9_n),
    .din(ffc_8_p)
  );


  DROC
  ffc_10
  (
    .doutp(ffc_10_p),
    .doutn(ffc_10_n),
    .din(ffc_9_p)
  );


  DROC
  ffc_11
  (
    .doutp(ffc_11_p),
    .doutn(ffc_11_n),
    .din(ffc_177_p)
  );


  DROC
  ffc_12
  (
    .doutp(ffc_12_p),
    .doutn(ffc_12_n),
    .din(ffc_179_p)
  );


  DROC
  ffc_13
  (
    .doutp(ffc_13_p),
    .doutn(ffc_13_n),
    .din(G12_p)
  );


  DROC
  ffc_14
  (
    .doutp(ffc_14_p),
    .doutn(ffc_14_n),
    .din(ffc_13_p)
  );


  DROC
  ffc_15
  (
    .doutp(ffc_15_p),
    .doutn(ffc_15_n),
    .din(ffc_14_p)
  );


  DROC
  ffc_16
  (
    .doutp(ffc_16_p),
    .doutn(ffc_16_n),
    .din(G13_p)
  );


  DROC
  ffc_17
  (
    .doutp(ffc_17_p),
    .doutn(ffc_17_n),
    .din(ffc_16_p)
  );


  DROC
  ffc_18
  (
    .doutp(ffc_18_p),
    .doutn(ffc_18_n),
    .din(ffc_17_p)
  );


  DROC
  ffc_19
  (
    .doutp(ffc_19_p),
    .doutn(ffc_19_n),
    .din(G14_p)
  );


  DROC
  ffc_20
  (
    .doutp(ffc_20_p),
    .doutn(ffc_20_n),
    .din(ffc_19_p)
  );


  DROC
  ffc_21
  (
    .doutp(ffc_21_p),
    .doutn(ffc_21_n),
    .din(ffc_20_p)
  );


  DROC
  ffc_22
  (
    .doutp(ffc_22_p),
    .doutn(ffc_22_n),
    .din(G15_p)
  );


  DROC
  ffc_23
  (
    .doutp(ffc_23_p),
    .doutn(ffc_23_n),
    .din(ffc_22_p)
  );


  DROC
  ffc_24
  (
    .doutp(ffc_24_p),
    .doutn(ffc_24_n),
    .din(ffc_23_p)
  );


  DROC
  ffc_25
  (
    .doutp(ffc_25_p),
    .doutn(ffc_25_n),
    .din(ffc_24_p)
  );


  DROC
  ffc_26
  (
    .doutp(ffc_26_p),
    .doutn(ffc_26_n),
    .din(ffc_186_p)
  );


  DROC
  ffc_27
  (
    .doutp(ffc_27_p),
    .doutn(ffc_27_n),
    .din(ffc_183_p)
  );


  DROC
  ffc_28
  (
    .doutp(ffc_28_p),
    .doutn(ffc_28_n),
    .din(G18_p)
  );


  DROC
  ffc_29
  (
    .doutp(ffc_29_p),
    .doutn(ffc_29_n),
    .din(ffc_28_p)
  );


  DROC
  ffc_30
  (
    .doutp(ffc_30_p),
    .doutn(ffc_30_n),
    .din(ffc_29_p)
  );


  DROC
  ffc_31
  (
    .doutp(ffc_31_p),
    .doutn(ffc_31_n),
    .din(ffc_30_p)
  );


  DROC
  ffc_32
  (
    .doutp(ffc_32_p),
    .doutn(ffc_32_n),
    .din(G19_p)
  );


  DROC
  ffc_33
  (
    .doutp(ffc_33_p),
    .doutn(ffc_33_n),
    .din(ffc_32_p)
  );


  DROC
  ffc_34
  (
    .doutp(ffc_34_p),
    .doutn(ffc_34_n),
    .din(ffc_33_p)
  );


  DROC
  ffc_35
  (
    .doutp(ffc_35_p),
    .doutn(ffc_35_n),
    .din(ffc_34_p)
  );


  DROC
  ffc_36
  (
    .doutp(ffc_36_p),
    .doutn(ffc_36_n),
    .din(G20_p)
  );


  DROC
  ffc_37
  (
    .doutp(ffc_37_p),
    .doutn(ffc_37_n),
    .din(ffc_36_p)
  );


  DROC
  ffc_38
  (
    .doutp(ffc_38_p),
    .doutn(ffc_38_n),
    .din(ffc_37_p)
  );


  DROC
  ffc_39
  (
    .doutp(ffc_39_p),
    .doutn(ffc_39_n),
    .din(ffc_38_p)
  );


  DROC
  ffc_40
  (
    .doutp(ffc_40_p),
    .doutn(ffc_40_n),
    .din(G21_p)
  );


  DROC
  ffc_41
  (
    .doutp(ffc_41_p),
    .doutn(ffc_41_n),
    .din(ffc_40_p)
  );


  DROC
  ffc_42
  (
    .doutp(ffc_42_p),
    .doutn(ffc_42_n),
    .din(ffc_41_p)
  );


  DROC
  ffc_43
  (
    .doutp(ffc_43_p),
    .doutn(ffc_43_n),
    .din(ffc_42_p)
  );


  DROC
  ffc_44
  (
    .doutp(ffc_44_p),
    .doutn(ffc_44_n),
    .din(G22_p)
  );


  DROC
  ffc_45
  (
    .doutp(ffc_45_p),
    .doutn(ffc_45_n),
    .din(ffc_44_p)
  );


  DROC
  ffc_46
  (
    .doutp(ffc_46_p),
    .doutn(ffc_46_n),
    .din(ffc_45_p)
  );


  DROC
  ffc_47
  (
    .doutp(ffc_47_p),
    .doutn(ffc_47_n),
    .din(ffc_46_p)
  );


  DROC
  ffc_48
  (
    .doutp(ffc_48_p),
    .doutn(ffc_48_n),
    .din(G23_p)
  );


  DROC
  ffc_49
  (
    .doutp(ffc_49_p),
    .doutn(ffc_49_n),
    .din(ffc_48_p)
  );


  DROC
  ffc_50
  (
    .doutp(ffc_50_p),
    .doutn(ffc_50_n),
    .din(ffc_49_p)
  );


  DROC
  ffc_51
  (
    .doutp(ffc_51_p),
    .doutn(ffc_51_n),
    .din(ffc_50_p)
  );


  DROC
  ffc_52
  (
    .doutp(ffc_52_p),
    .doutn(ffc_52_n),
    .din(G24_p)
  );


  DROC
  ffc_53
  (
    .doutp(ffc_53_p),
    .doutn(ffc_53_n),
    .din(ffc_52_p)
  );


  DROC
  ffc_54
  (
    .doutp(ffc_54_p),
    .doutn(ffc_54_n),
    .din(ffc_53_p)
  );


  DROC
  ffc_55
  (
    .doutp(ffc_55_p),
    .doutn(ffc_55_n),
    .din(ffc_54_p_spl_)
  );


  DROC
  ffc_56
  (
    .doutp(ffc_56_p),
    .doutn(ffc_56_n),
    .din(G25_p)
  );


  DROC
  ffc_57
  (
    .doutp(ffc_57_p),
    .doutn(ffc_57_n),
    .din(ffc_56_p)
  );


  DROC
  ffc_58
  (
    .doutp(ffc_58_p),
    .doutn(ffc_58_n),
    .din(ffc_57_p)
  );


  DROC
  ffc_59
  (
    .doutp(ffc_59_p),
    .doutn(ffc_59_n),
    .din(ffc_58_p_spl_)
  );


  DROC
  ffc_60
  (
    .doutp(ffc_60_p),
    .doutn(ffc_60_n),
    .din(G26_p)
  );


  DROC
  ffc_61
  (
    .doutp(ffc_61_p),
    .doutn(ffc_61_n),
    .din(ffc_60_p)
  );


  DROC
  ffc_62
  (
    .doutp(ffc_62_p),
    .doutn(ffc_62_n),
    .din(ffc_61_p)
  );


  DROC
  ffc_63
  (
    .doutp(ffc_63_p),
    .doutn(ffc_63_n),
    .din(ffc_62_p_spl_)
  );


  DROC
  ffc_64
  (
    .doutp(ffc_64_p),
    .doutn(ffc_64_n),
    .din(G27_p)
  );


  DROC
  ffc_65
  (
    .doutp(ffc_65_p),
    .doutn(ffc_65_n),
    .din(ffc_64_p)
  );


  DROC
  ffc_66
  (
    .doutp(ffc_66_p),
    .doutn(ffc_66_n),
    .din(ffc_254_p_spl_)
  );


  DROC
  ffc_67
  (
    .doutp(ffc_67_p),
    .doutn(ffc_67_n),
    .din(G28_p)
  );


  DROC
  ffc_68
  (
    .doutp(ffc_68_p),
    .doutn(ffc_68_n),
    .din(ffc_67_p)
  );


  DROC
  ffc_69
  (
    .doutp(ffc_69_p),
    .doutn(ffc_69_n),
    .din(G29_p)
  );


  DROC
  ffc_70
  (
    .doutp(ffc_70_p),
    .doutn(ffc_70_n),
    .din(ffc_209_p_spl_)
  );


  DROC
  ffc_71
  (
    .doutp(ffc_71_p),
    .doutn(ffc_71_n),
    .din(G30_p)
  );


  DROC
  ffc_72
  (
    .doutp(ffc_72_p),
    .doutn(ffc_72_n),
    .din(ffc_200_p_spl_)
  );


  DROC
  ffc_73
  (
    .doutp(ffc_73_p),
    .doutn(ffc_73_n),
    .din(G31_p)
  );


  DROC
  ffc_74
  (
    .doutp(ffc_74_p),
    .doutn(ffc_74_n),
    .din(G32_p)
  );


  DROC
  ffc_75
  (
    .doutp(ffc_75_p),
    .doutn(ffc_75_n),
    .din(ffc_74_p)
  );


  DROC
  ffc_76
  (
    .doutp(ffc_76_p),
    .doutn(ffc_76_n),
    .din(ffc_75_p)
  );


  DROC
  ffc_77
  (
    .doutp(ffc_77_p),
    .doutn(ffc_77_n),
    .din(ffc_76_p)
  );


  DROC
  ffc_78
  (
    .doutp(ffc_78_p),
    .doutn(ffc_78_n),
    .din(G33_p)
  );


  DROC
  ffc_79
  (
    .doutp(ffc_79_p),
    .doutn(ffc_79_n),
    .din(ffc_78_p)
  );


  DROC
  ffc_80
  (
    .doutp(ffc_80_p),
    .doutn(ffc_80_n),
    .din(ffc_79_p)
  );


  DROC
  ffc_81
  (
    .doutp(ffc_81_p),
    .doutn(ffc_81_n),
    .din(ffc_80_p)
  );


  DROC
  ffc_82
  (
    .doutp(ffc_82_p),
    .doutn(ffc_82_n),
    .din(G34_p)
  );


  DROC
  ffc_83
  (
    .doutp(ffc_83_p),
    .doutn(ffc_83_n),
    .din(ffc_82_p)
  );


  DROC
  ffc_84
  (
    .doutp(ffc_84_p),
    .doutn(ffc_84_n),
    .din(G35_p)
  );


  DROC
  ffc_85
  (
    .doutp(ffc_85_p),
    .doutn(ffc_85_n),
    .din(ffc_84_p)
  );


  DROC
  ffc_86
  (
    .doutp(ffc_86_p),
    .doutn(ffc_86_n),
    .din(G36_p)
  );


  DROC
  ffc_87
  (
    .doutp(ffc_87_p),
    .doutn(ffc_87_n),
    .din(G37_p)
  );


  DROC
  ffc_88
  (
    .doutp(ffc_88_p),
    .doutn(ffc_88_n),
    .din(G38_p)
  );


  DROC
  ffc_89
  (
    .doutp(ffc_89_p),
    .doutn(ffc_89_n),
    .din(ffc_88_p)
  );


  DROC
  ffc_90
  (
    .doutp(ffc_90_p),
    .doutn(ffc_90_n),
    .din(G41_p)
  );


  DROC
  ffc_91
  (
    .doutp(ffc_91_p),
    .doutn(ffc_91_n),
    .din(ffc_90_p)
  );


  DROC
  ffc_92
  (
    .doutp(ffc_92_p),
    .doutn(ffc_92_n),
    .din(ffc_91_p)
  );


  DROC
  ffc_93
  (
    .doutp(ffc_93_p),
    .doutn(ffc_93_n),
    .din(ffc_92_p_spl_)
  );


  DROC
  ffc_94
  (
    .doutp(ffc_94_p),
    .doutn(ffc_94_n),
    .din(G42_p)
  );


  DROC
  ffc_95
  (
    .doutp(ffc_95_p),
    .doutn(ffc_95_n),
    .din(ffc_94_p)
  );


  DROC
  ffc_96
  (
    .doutp(ffc_96_p),
    .doutn(ffc_96_n),
    .din(ffc_95_p)
  );


  DROC
  ffc_97
  (
    .doutp(ffc_97_p),
    .doutn(ffc_97_n),
    .din(ffc_96_p_spl_)
  );


  DROC
  ffc_98
  (
    .doutp(ffc_98_p),
    .doutn(ffc_98_n),
    .din(G43_p)
  );


  DROC
  ffc_99
  (
    .doutp(ffc_99_p),
    .doutn(ffc_99_n),
    .din(ffc_98_p)
  );


  DROC
  ffc_100
  (
    .doutp(ffc_100_p),
    .doutn(ffc_100_n),
    .din(ffc_99_p)
  );


  DROC
  ffc_101
  (
    .doutp(ffc_101_p),
    .doutn(ffc_101_n),
    .din(ffc_100_p_spl_)
  );


  DROC
  ffc_102
  (
    .doutp(ffc_102_p),
    .doutn(ffc_102_n),
    .din(G44_p)
  );


  DROC
  ffc_103
  (
    .doutp(ffc_103_p),
    .doutn(ffc_103_n),
    .din(ffc_102_p)
  );


  DROC
  ffc_104
  (
    .doutp(ffc_104_p),
    .doutn(ffc_104_n),
    .din(ffc_103_p)
  );


  DROC
  ffc_105
  (
    .doutp(ffc_105_p),
    .doutn(ffc_105_n),
    .din(ffc_104_p_spl_)
  );


  DROC
  ffc_106
  (
    .doutp(ffc_106_p),
    .doutn(ffc_106_n),
    .din(G45_p)
  );


  DROC
  ffc_107
  (
    .doutp(ffc_107_p),
    .doutn(ffc_107_n),
    .din(ffc_106_p)
  );


  DROC
  ffc_108
  (
    .doutp(ffc_108_p),
    .doutn(ffc_108_n),
    .din(ffc_257_p_spl_)
  );


  DROC
  ffc_109
  (
    .doutp(ffc_109_p),
    .doutn(ffc_109_n),
    .din(G46_p)
  );


  DROC
  ffc_110
  (
    .doutp(ffc_110_p),
    .doutn(ffc_110_n),
    .din(ffc_109_p)
  );


  DROC
  ffc_111
  (
    .doutp(ffc_111_p),
    .doutn(ffc_111_n),
    .din(ffc_236_p_spl_)
  );


  DROC
  ffc_112
  (
    .doutp(ffc_112_p),
    .doutn(ffc_112_n),
    .din(G47_p)
  );


  DROC
  ffc_113
  (
    .doutp(ffc_113_p),
    .doutn(ffc_113_n),
    .din(ffc_211_p_spl_)
  );


  DROC
  ffc_114
  (
    .doutp(ffc_114_p),
    .doutn(ffc_114_n),
    .din(G48_p)
  );


  DROC
  ffc_115
  (
    .doutp(ffc_115_p),
    .doutn(ffc_115_n),
    .din(ffc_202_p_spl_)
  );


  DROC
  ffc_116
  (
    .doutp(ffc_116_p),
    .doutn(ffc_116_n),
    .din(G49_p)
  );


  DROC
  ffc_117
  (
    .doutp(ffc_117_p),
    .doutn(ffc_117_n),
    .din(ffc_116_p)
  );


  DROC
  ffc_118
  (
    .doutp(ffc_118_p),
    .doutn(ffc_118_n),
    .din(ffc_117_p)
  );


  DROC
  ffc_119
  (
    .doutp(ffc_119_p),
    .doutn(ffc_119_n),
    .din(ffc_118_p)
  );


  DROC
  ffc_120
  (
    .doutp(ffc_120_p),
    .doutn(ffc_120_n),
    .din(G50_p)
  );


  DROC
  ffc_121
  (
    .doutp(ffc_121_p),
    .doutn(ffc_121_n),
    .din(ffc_120_p)
  );


  DROC
  ffc_122
  (
    .doutp(ffc_122_p),
    .doutn(ffc_122_n),
    .din(ffc_121_p)
  );


  DROC
  ffc_123
  (
    .doutp(ffc_123_p),
    .doutn(ffc_123_n),
    .din(ffc_122_p_spl_)
  );


  DROC
  ffc_124
  (
    .doutp(ffc_124_p),
    .doutn(ffc_124_n),
    .din(G51_p)
  );


  DROC
  ffc_125
  (
    .doutp(ffc_125_p),
    .doutn(ffc_125_n),
    .din(ffc_124_p)
  );


  DROC
  ffc_126
  (
    .doutp(ffc_126_p),
    .doutn(ffc_126_n),
    .din(ffc_125_p)
  );


  DROC
  ffc_127
  (
    .doutp(ffc_127_p),
    .doutn(ffc_127_n),
    .din(ffc_126_p)
  );


  DROC
  ffc_128
  (
    .doutp(ffc_128_p),
    .doutn(ffc_128_n),
    .din(G52_p)
  );


  DROC
  ffc_129
  (
    .doutp(ffc_129_p),
    .doutn(ffc_129_n),
    .din(ffc_128_p)
  );


  DROC
  ffc_130
  (
    .doutp(ffc_130_p),
    .doutn(ffc_130_n),
    .din(ffc_129_p)
  );


  DROC
  ffc_131
  (
    .doutp(ffc_131_p),
    .doutn(ffc_131_n),
    .din(ffc_130_p)
  );


  DROC
  ffc_132
  (
    .doutp(ffc_132_p),
    .doutn(ffc_132_n),
    .din(G53_p)
  );


  DROC
  ffc_133
  (
    .doutp(ffc_133_p),
    .doutn(ffc_133_n),
    .din(ffc_132_p)
  );


  DROC
  ffc_134
  (
    .doutp(ffc_134_p),
    .doutn(ffc_134_n),
    .din(ffc_133_p)
  );


  DROC
  ffc_135
  (
    .doutp(ffc_135_p),
    .doutn(ffc_135_n),
    .din(ffc_134_p)
  );


  DROC
  ffc_136
  (
    .doutp(ffc_136_p),
    .doutn(ffc_136_n),
    .din(G54_p)
  );


  DROC
  ffc_137
  (
    .doutp(ffc_137_p),
    .doutn(ffc_137_n),
    .din(ffc_136_p)
  );


  DROC
  ffc_138
  (
    .doutp(ffc_138_p),
    .doutn(ffc_138_n),
    .din(ffc_137_p)
  );


  DROC
  ffc_139
  (
    .doutp(ffc_139_p),
    .doutn(ffc_139_n),
    .din(ffc_138_p)
  );


  DROC
  ffc_140
  (
    .doutp(ffc_140_p),
    .doutn(ffc_140_n),
    .din(G55_p)
  );


  DROC
  ffc_141
  (
    .doutp(ffc_141_p),
    .doutn(ffc_141_n),
    .din(ffc_140_p)
  );


  DROC
  ffc_142
  (
    .doutp(ffc_142_p),
    .doutn(ffc_142_n),
    .din(ffc_141_p)
  );


  DROC
  ffc_143
  (
    .doutp(ffc_143_p),
    .doutn(ffc_143_n),
    .din(ffc_142_p_spl_)
  );


  DROC
  ffc_144
  (
    .doutp(ffc_144_p),
    .doutn(ffc_144_n),
    .din(G56_p)
  );


  DROC
  ffc_145
  (
    .doutp(ffc_145_p),
    .doutn(ffc_145_n),
    .din(ffc_144_p)
  );


  DROC
  ffc_146
  (
    .doutp(ffc_146_p),
    .doutn(ffc_146_n),
    .din(ffc_145_p)
  );


  DROC
  ffc_147
  (
    .doutp(ffc_147_p),
    .doutn(ffc_147_n),
    .din(G57_p)
  );


  DROC
  ffc_148
  (
    .doutp(ffc_148_p),
    .doutn(ffc_148_n),
    .din(ffc_147_p)
  );


  DROC
  ffc_149
  (
    .doutp(ffc_149_p),
    .doutn(ffc_149_n),
    .din(ffc_148_p)
  );


  DROC
  ffc_150
  (
    .doutp(ffc_150_p),
    .doutn(ffc_150_n),
    .din(ffc_149_p)
  );


  DROC
  ffc_151
  (
    .doutp(ffc_151_p),
    .doutn(ffc_151_n),
    .din(G58_p)
  );


  DROC
  ffc_152
  (
    .doutp(ffc_152_p),
    .doutn(ffc_152_n),
    .din(ffc_206_p)
  );


  DROC
  ffc_153
  (
    .doutp(ffc_153_p),
    .doutn(ffc_153_n),
    .din(G59_p)
  );


  DROC
  ffc_154
  (
    .doutp(ffc_154_p),
    .doutn(ffc_154_n),
    .din(ffc_153_p)
  );


  DROC
  ffc_155
  (
    .doutp(ffc_155_p),
    .doutn(ffc_155_n),
    .din(ffc_154_p)
  );


  DROC
  ffc_156
  (
    .doutp(ffc_156_p),
    .doutn(ffc_156_n),
    .din(ffc_155_p)
  );


  DROC
  ffc_157
  (
    .doutp(ffc_157_p),
    .doutn(ffc_157_n),
    .din(ffc_192_p)
  );


  DROC
  ffc_158
  (
    .doutp(ffc_158_p),
    .doutn(ffc_158_n),
    .din(ffc_188_p)
  );


  DROC
  ffc_159
  (
    .doutp(ffc_159_p),
    .doutn(ffc_159_n),
    .din(ffc_189_p)
  );


  DROC
  ffc_160
  (
    .doutp(ffc_160_p),
    .doutn(ffc_160_n),
    .din(ffc_187_p)
  );


  DROC
  ffc_161
  (
    .doutp(ffc_161_p),
    .doutn(ffc_161_n),
    .din(ffc_204_p)
  );


  DROC
  ffc_162
  (
    .doutp(ffc_162_p),
    .doutn(ffc_162_n),
    .din(ffc_207_p)
  );


  DROC
  ffc_163
  (
    .doutp(ffc_163_p),
    .doutn(ffc_163_n),
    .din(ffc_213_p)
  );


  DROC
  ffc_164
  (
    .doutp(ffc_164_p),
    .doutn(ffc_164_n),
    .din(ffc_214_p)
  );


  DROC
  ffc_165
  (
    .doutp(ffc_165_p),
    .doutn(ffc_165_n),
    .din(ffc_215_p)
  );


  DROC
  ffc_166
  (
    .doutp(ffc_166_p),
    .doutn(ffc_166_n),
    .din(ffc_226_p)
  );


  DROC
  ffc_167
  (
    .doutp(ffc_167_p),
    .doutn(ffc_167_n),
    .din(ffc_227_p)
  );


  DROC
  ffc_168
  (
    .doutp(ffc_168_p),
    .doutn(ffc_168_n),
    .din(ffc_239_p)
  );


  DROC
  ffc_169
  (
    .doutp(ffc_169_p),
    .doutn(ffc_169_n),
    .din(ffc_240_p)
  );


  DROC
  ffc_170
  (
    .doutp(ffc_170_p),
    .doutn(ffc_170_n),
    .din(ffc_241_p)
  );


  DROC
  ffc_171
  (
    .doutp(ffc_171_p),
    .doutn(ffc_171_n),
    .din(ffc_249_p)
  );


  DROC
  ffc_172
  (
    .doutp(ffc_172_p),
    .doutn(ffc_172_n),
    .din(ffc_250_p)
  );


  DROC
  ffc_173
  (
    .doutp(ffc_173_p),
    .doutn(ffc_173_n),
    .din(ffc_268_p)
  );


  DROC
  ffc_174
  (
    .doutp(ffc_174_p),
    .doutn(ffc_174_n),
    .din(ffc_271_p)
  );


  DROC
  ffc_175
  (
    .doutp(ffc_175_p),
    .doutn(ffc_175_n),
    .din(ffc_216_p)
  );


  DROC
  ffc_176
  (
    .doutp(ffc_176_p),
    .doutn(ffc_176_n),
    .din(ffc_217_p_spl_)
  );


  DROC
  ffc_177
  (
    .doutp(ffc_177_p),
    .doutn(ffc_177_n),
    .din(ffc_218_p)
  );


  DROC
  ffc_178
  (
    .doutp(ffc_178_p),
    .doutn(ffc_178_n),
    .din(ffc_219_p)
  );


  DROC
  ffc_179
  (
    .doutp(ffc_179_p),
    .doutn(ffc_179_n),
    .din(ffc_220_p)
  );


  DROC
  ffc_180
  (
    .doutp(ffc_180_p),
    .doutn(ffc_180_n),
    .din(ffc_222_p)
  );


  DROC
  ffc_181
  (
    .doutp(ffc_181_p),
    .doutn(ffc_181_n),
    .din(ffc_223_p)
  );


  DROC
  ffc_182
  (
    .doutp(ffc_182_p),
    .doutn(ffc_182_n),
    .din(ffc_224_p)
  );


  DROC
  ffc_183
  (
    .doutp(ffc_183_p),
    .doutn(ffc_183_n),
    .din(ffc_225_p)
  );


  DROC
  ffc_184
  (
    .doutp(ffc_184_p),
    .doutn(ffc_184_n),
    .din(ffc_276_p)
  );


  DROC
  ffc_185
  (
    .doutp(ffc_185_p),
    .doutn(ffc_185_n),
    .din(ffc_279_p)
  );


  DROC
  ffc_186
  (
    .doutp(ffc_186_p),
    .doutn(ffc_186_n),
    .din(ffc_230_p)
  );


  DROC
  ffc_187
  (
    .doutp(ffc_187_p),
    .doutn(ffc_187_n),
    .din(ffc_229_p)
  );


  DROC
  ffc_188
  (
    .doutp(ffc_188_p),
    .doutn(ffc_188_n),
    .din(ffc_231_p)
  );


  DROC
  ffc_189
  (
    .doutp(ffc_189_p),
    .doutn(ffc_189_n),
    .din(ffc_232_p)
  );


  DROC
  ffc_190
  (
    .doutp(ffc_190_p),
    .doutn(ffc_190_n),
    .din(ffc_242_p)
  );


  DROC
  ffc_191
  (
    .doutp(ffc_191_n),
    .doutn(ffc_191_p),
    .din(g548_n_spl_)
  );


  DROC
  ffc_192
  (
    .doutp(ffc_192_p),
    .doutn(ffc_192_n),
    .din(ffc_243_p_spl_)
  );


  DROC
  ffc_193
  (
    .doutp(ffc_193_n),
    .doutn(ffc_193_p),
    .din(g549_p_spl_)
  );


  DROC
  ffc_194
  (
    .doutp(ffc_194_n),
    .doutn(ffc_194_p),
    .din(g550_n_spl_)
  );


  DROC
  ffc_195
  (
    .doutp(ffc_195_p),
    .doutn(ffc_195_n),
    .din(ffc_251_p)
  );


  DROC
  ffc_196
  (
    .doutp(ffc_196_n),
    .doutn(ffc_196_p),
    .din(g551_p_spl_)
  );


  DROC
  ffc_197
  (
    .doutp(ffc_197_n),
    .doutn(ffc_197_p),
    .din(g552_p_spl_)
  );


  DROC
  ffc_198
  (
    .doutp(ffc_198_p),
    .doutn(ffc_198_n),
    .din(ffc_252_p_spl_)
  );


  DROC
  ffc_199
  (
    .doutp(ffc_199_p),
    .doutn(ffc_199_n),
    .din(ffc_272_p)
  );


  DROC
  ffc_200
  (
    .doutp(ffc_200_p),
    .doutn(ffc_200_n),
    .din(ffc_275_p)
  );


  DROC
  ffc_201
  (
    .doutp(ffc_201_n),
    .doutn(ffc_201_p),
    .din(g553_n_spl_)
  );


  DROC
  ffc_202
  (
    .doutp(ffc_202_p),
    .doutn(ffc_202_n),
    .din(ffc_277_p)
  );


  DROC
  ffc_203
  (
    .doutp(ffc_203_n),
    .doutn(ffc_203_p),
    .din(g558_p_spl_)
  );


  DROC
  ffc_204
  (
    .doutp(ffc_204_p),
    .doutn(ffc_204_n),
    .din(ffc_280_p)
  );


  DROC
  ffc_205
  (
    .doutp(ffc_205_p),
    .doutn(ffc_205_n),
    .din(ffc_290_p)
  );


  DROC
  ffc_206
  (
    .doutp(ffc_206_p),
    .doutn(ffc_206_n),
    .din(ffc_291_p)
  );


  DROC
  ffc_207
  (
    .doutp(ffc_207_p),
    .doutn(ffc_207_n),
    .din(ffc_296_p)
  );


  DROC
  ffc_208
  (
    .doutp(ffc_208_n),
    .doutn(ffc_208_p),
    .din(g559_n_spl_)
  );


  DROC
  ffc_209
  (
    .doutp(ffc_209_p),
    .doutn(ffc_209_n),
    .din(ffc_286_p)
  );


  DROC
  ffc_210
  (
    .doutp(ffc_210_n),
    .doutn(ffc_210_p),
    .din(g560_p_spl_)
  );


  DROC
  ffc_211
  (
    .doutp(ffc_211_p),
    .doutn(ffc_211_n),
    .din(ffc_287_p)
  );


  DROC
  ffc_212
  (
    .doutp(ffc_212_n),
    .doutn(ffc_212_p),
    .din(g562_p_spl_)
  );


  DROC
  ffc_213
  (
    .doutp(ffc_213_n),
    .doutn(ffc_213_p),
    .din(g563_n_spl_)
  );


  DROC
  ffc_214
  (
    .doutp(ffc_214_n),
    .doutn(ffc_214_p),
    .din(g564_n_spl_)
  );


  DROC
  ffc_215
  (
    .doutp(ffc_215_n),
    .doutn(ffc_215_p),
    .din(g565_p_spl_)
  );


  DROC
  ffc_216
  (
    .doutp(ffc_216_p),
    .doutn(ffc_216_n),
    .din(ffc_281_p)
  );


  DROC
  ffc_217
  (
    .doutp(ffc_217_p),
    .doutn(ffc_217_n),
    .din(ffc_282_p)
  );


  DROC
  ffc_218
  (
    .doutp(ffc_218_p),
    .doutn(ffc_218_n),
    .din(ffc_283_p)
  );


  DROC
  ffc_219
  (
    .doutp(ffc_219_p),
    .doutn(ffc_219_n),
    .din(ffc_284_p)
  );


  DROC
  ffc_220
  (
    .doutp(ffc_220_p),
    .doutn(ffc_220_n),
    .din(ffc_285_p)
  );


  DROC
  ffc_221
  (
    .doutp(ffc_221_p),
    .doutn(ffc_221_n),
    .din(ffc_85_p_spl_)
  );


  DROC
  ffc_222
  (
    .doutp(ffc_222_p),
    .doutn(ffc_222_n),
    .din(ffc_292_p)
  );


  DROC
  ffc_223
  (
    .doutp(ffc_223_p),
    .doutn(ffc_223_n),
    .din(ffc_293_p)
  );


  DROC
  ffc_224
  (
    .doutp(ffc_224_p),
    .doutn(ffc_224_n),
    .din(ffc_294_p)
  );


  DROC
  ffc_225
  (
    .doutp(ffc_225_p),
    .doutn(ffc_225_n),
    .din(ffc_295_p)
  );


  DROC
  ffc_226
  (
    .doutp(ffc_226_n),
    .doutn(ffc_226_p),
    .din(g566_p_spl_)
  );


  DROC
  ffc_227
  (
    .doutp(ffc_227_n),
    .doutn(ffc_227_p),
    .din(g567_p_spl_)
  );


  DROC
  ffc_228
  (
    .doutp(ffc_228_p),
    .doutn(ffc_228_n),
    .din(ffc_298_p_spl_)
  );


  DROC
  ffc_229
  (
    .doutp(ffc_229_p),
    .doutn(ffc_229_n),
    .din(ffc_302_p)
  );


  DROC
  ffc_230
  (
    .doutp(ffc_230_p),
    .doutn(ffc_230_n),
    .din(ffc_305_p_spl_)
  );


  DROC
  ffc_231
  (
    .doutp(ffc_231_p),
    .doutn(ffc_231_n),
    .din(ffc_306_p_spl_1)
  );


  DROC
  ffc_232
  (
    .doutp(ffc_232_p),
    .doutn(ffc_232_n),
    .din(ffc_307_p_spl_)
  );


  DROC
  ffc_233
  (
    .doutp(ffc_233_p),
    .doutn(ffc_233_n),
    .din(ffc_68_p_spl_)
  );


  DROC
  ffc_234
  (
    .doutp(ffc_234_p),
    .doutn(ffc_234_n),
    .din(ffc_83_p_spl_)
  );


  DROC
  ffc_235
  (
    .doutp(ffc_235_n),
    .doutn(ffc_235_p),
    .din(g568_n_spl_)
  );


  DROC
  ffc_236
  (
    .doutp(ffc_236_p),
    .doutn(ffc_236_n),
    .din(ffc_110_p)
  );


  DROC
  ffc_237
  (
    .doutp(ffc_237_n),
    .doutn(ffc_237_p),
    .din(g571_n_spl_)
  );


  DROC
  ffc_238
  (
    .doutp(ffc_238_p),
    .doutn(ffc_238_n),
    .din(g577_n_spl_)
  );


  DROC
  ffc_239
  (
    .doutp(ffc_239_n),
    .doutn(ffc_239_p),
    .din(g578_n_spl_)
  );


  DROC
  ffc_240
  (
    .doutp(ffc_240_n),
    .doutn(ffc_240_p),
    .din(g582_p_spl_)
  );


  DROC
  ffc_241
  (
    .doutp(ffc_241_n),
    .doutn(ffc_241_p),
    .din(g583_n_spl_)
  );


  DROC
  ffc_242
  (
    .doutp(ffc_242_p),
    .doutn(ffc_242_n),
    .din(ffc_303_p_spl_)
  );


  DROC
  ffc_243
  (
    .doutp(ffc_243_p),
    .doutn(ffc_243_n),
    .din(ffc_304_p)
  );


  DROC
  ffc_244
  (
    .doutp(ffc_244_n),
    .doutn(ffc_244_p),
    .din(g585_n_spl_)
  );


  DROC
  ffc_245
  (
    .doutp(ffc_245_n),
    .doutn(ffc_245_p),
    .din(g587_n_spl_)
  );


  DROC
  ffc_246
  (
    .doutp(ffc_246_n),
    .doutn(ffc_246_p),
    .din(g589_n_spl_)
  );


  DROC
  ffc_247
  (
    .doutp(ffc_247_p),
    .doutn(ffc_247_n),
    .din(g591_p_spl_)
  );


  DROC
  ffc_248
  (
    .doutp(ffc_248_p),
    .doutn(ffc_248_n),
    .din(ffc_299_p_spl_)
  );


  DROC
  ffc_249
  (
    .doutp(ffc_249_n),
    .doutn(ffc_249_p),
    .din(g592_n_spl_)
  );


  DROC
  ffc_250
  (
    .doutp(ffc_250_n),
    .doutn(ffc_250_p),
    .din(g593_p_spl_)
  );


  DROC
  ffc_251
  (
    .doutp(ffc_251_p),
    .doutn(ffc_251_n),
    .din(ffc_73_p_spl_)
  );


  DROC
  ffc_252
  (
    .doutp(ffc_252_p),
    .doutn(ffc_252_n),
    .din(g599_n_spl_)
  );


  DROC
  ffc_253
  (
    .doutp(ffc_253_p),
    .doutn(ffc_253_n),
    .din(g601_p_spl_)
  );


  DROC
  ffc_254
  (
    .doutp(ffc_254_p),
    .doutn(ffc_254_n),
    .din(ffc_65_p_spl_)
  );


  DROC
  ffc_255
  (
    .doutp(ffc_255_p),
    .doutn(ffc_255_n),
    .din(g602_p)
  );


  DROC
  ffc_256
  (
    .doutp(ffc_256_p),
    .doutn(ffc_256_n),
    .din(g603_p)
  );


  DROC
  ffc_257
  (
    .doutp(ffc_257_p),
    .doutn(ffc_257_n),
    .din(ffc_107_p_spl_)
  );


  DROC
  ffc_258
  (
    .doutp(ffc_258_p),
    .doutn(ffc_258_n),
    .din(g604_p)
  );


  DROC
  ffc_259
  (
    .doutp(ffc_259_p),
    .doutn(ffc_259_n),
    .din(g607_p)
  );


  DROC
  ffc_260
  (
    .doutp(ffc_260_p),
    .doutn(ffc_260_n),
    .din(g613_n)
  );


  DROC
  ffc_261
  (
    .doutp(ffc_261_p),
    .doutn(ffc_261_n),
    .din(g616_p)
  );


  DROC
  ffc_262
  (
    .doutp(ffc_262_p),
    .doutn(ffc_262_n),
    .din(g619_p)
  );


  DROC
  ffc_263
  (
    .doutp(ffc_263_p),
    .doutn(ffc_263_n),
    .din(g622_p)
  );


  DROC
  ffc_264
  (
    .doutp(ffc_264_p),
    .doutn(ffc_264_n),
    .din(g625_p)
  );


  DROC
  ffc_265
  (
    .doutp(ffc_265_p),
    .doutn(ffc_265_n),
    .din(g628_p)
  );


  DROC
  ffc_266
  (
    .doutp(ffc_266_n),
    .doutn(ffc_266_p),
    .din(g630_p)
  );


  DROC
  ffc_267
  (
    .doutp(ffc_267_p),
    .doutn(ffc_267_n),
    .din(g633_p)
  );


  DROC
  ffc_268
  (
    .doutp(ffc_268_n),
    .doutn(ffc_268_p),
    .din(g634_p_spl_)
  );


  DROC
  ffc_269
  (
    .doutp(ffc_269_p),
    .doutn(ffc_269_n),
    .din(g637_p)
  );


  DROC
  ffc_270
  (
    .doutp(ffc_270_n),
    .doutn(ffc_270_p),
    .din(g640_n)
  );


  DROC
  ffc_271
  (
    .doutp(ffc_271_p),
    .doutn(ffc_271_n),
    .din(g644_n_spl_)
  );


  DROC
  ffc_272
  (
    .doutp(ffc_272_p),
    .doutn(ffc_272_n),
    .din(ffc_87_p_spl_)
  );


  DROC
  ffc_273
  (
    .doutp(ffc_273_p),
    .doutn(ffc_273_n),
    .din(g645_p)
  );


  DROC
  ffc_274
  (
    .doutp(ffc_274_p),
    .doutn(ffc_274_n),
    .din(g646_p)
  );


  DROC
  ffc_275
  (
    .doutp(ffc_275_p),
    .doutn(ffc_275_n),
    .din(ffc_71_p_spl_)
  );


  DROC
  ffc_276
  (
    .doutp(ffc_276_p),
    .doutn(ffc_276_n),
    .din(g647_n)
  );


  DROC
  ffc_277
  (
    .doutp(ffc_277_p),
    .doutn(ffc_277_n),
    .din(ffc_114_p_spl_)
  );


  DROC
  ffc_278
  (
    .doutp(ffc_278_n),
    .doutn(ffc_278_p),
    .din(g651_p)
  );


  DROC
  ffc_279
  (
    .doutp(ffc_279_n),
    .doutn(ffc_279_p),
    .din(g653_n)
  );


  DROC
  ffc_280
  (
    .doutp(ffc_280_p),
    .doutn(ffc_280_n),
    .din(g657_n_spl_)
  );


  DROC
  ffc_281
  (
    .doutp(ffc_281_p),
    .doutn(ffc_281_n),
    .din(G1_p)
  );


  DROC
  ffc_282
  (
    .doutp(ffc_282_p),
    .doutn(ffc_282_n),
    .din(G4_p_spl_1)
  );


  DROC
  ffc_283
  (
    .doutp(ffc_283_p),
    .doutn(ffc_283_n),
    .din(G8_p_spl_)
  );


  DROC
  ffc_284
  (
    .doutp(ffc_284_p),
    .doutn(ffc_284_n),
    .din(G9_p)
  );


  DROC
  ffc_285
  (
    .doutp(ffc_285_p),
    .doutn(ffc_285_n),
    .din(G11_p_spl_)
  );


  DROC
  ffc_286
  (
    .doutp(ffc_286_p),
    .doutn(ffc_286_n),
    .din(ffc_69_p)
  );


  DROC
  ffc_287
  (
    .doutp(ffc_287_p),
    .doutn(ffc_287_n),
    .din(ffc_112_p)
  );


  DROC
  ffc_288
  (
    .doutp(ffc_288_p),
    .doutn(ffc_288_n),
    .din(g658_p)
  );


  DROC
  ffc_289
  (
    .doutp(ffc_289_p),
    .doutn(ffc_289_n),
    .din(g660_n)
  );


  DROC
  ffc_290
  (
    .doutp(ffc_290_p),
    .doutn(ffc_290_n),
    .din(ffc_86_p)
  );


  DROC
  ffc_291
  (
    .doutp(ffc_291_p),
    .doutn(ffc_291_n),
    .din(ffc_151_p)
  );


  DROC
  ffc_292
  (
    .doutp(ffc_292_p),
    .doutn(ffc_292_n),
    .din(G2_p_spl_)
  );


  DROC
  ffc_293
  (
    .doutp(ffc_293_p),
    .doutn(ffc_293_n),
    .din(G5_p)
  );


  DROC
  ffc_294
  (
    .doutp(ffc_294_p),
    .doutn(ffc_294_n),
    .din(G6_p_spl_)
  );


  DROC
  ffc_295
  (
    .doutp(ffc_295_p),
    .doutn(ffc_295_n),
    .din(G17_p_spl_)
  );


  DROC
  ffc_296
  (
    .doutp(ffc_296_p),
    .doutn(ffc_296_n),
    .din(g661_n)
  );


  DROC
  ffc_297
  (
    .doutp(ffc_297_n),
    .doutn(ffc_297_p),
    .din(g662_n_spl_)
  );


  DROC
  ffc_298
  (
    .doutp(ffc_298_n),
    .doutn(ffc_298_p),
    .din(g663_n_spl_)
  );


  DROC
  ffc_299
  (
    .doutp(ffc_299_p),
    .doutn(ffc_299_n),
    .din(G39_p)
  );


  DROC
  ffc_300
  (
    .doutp(ffc_300_p),
    .doutn(ffc_300_n),
    .din(g664_p)
  );


  DROC
  ffc_301
  (
    .doutp(ffc_301_p),
    .doutn(ffc_301_n),
    .din(g665_p)
  );


  DROC
  ffc_302
  (
    .doutp(ffc_302_p),
    .doutn(ffc_302_n),
    .din(g666_p)
  );


  DROC
  ffc_303
  (
    .doutp(ffc_303_p),
    .doutn(ffc_303_n),
    .din(G10_p)
  );


  DROC
  ffc_304
  (
    .doutp(ffc_304_p),
    .doutn(ffc_304_n),
    .din(G60_p)
  );


  DROC
  ffc_305
  (
    .doutp(ffc_305_p),
    .doutn(ffc_305_n),
    .din(G16_p)
  );


  DROC
  ffc_306
  (
    .doutp(ffc_306_n),
    .doutn(ffc_306_p),
    .din(g667_n)
  );


  DROC
  ffc_307
  (
    .doutp(ffc_307_p),
    .doutn(ffc_307_n),
    .din(g668_p)
  );


  DROC
  ffc_308
  (
    .doutp(ffc_308_p),
    .doutn(ffc_308_n),
    .din(g671_n)
  );


  buf

  (
    ffc_6_n_spl_,
    ffc_6_n
  );


  buf

  (
    ffc_26_n_spl_,
    ffc_26_n
  );


  buf

  (
    g370_n_spl_,
    g370_n
  );


  buf

  (
    ffc_10_n_spl_,
    ffc_10_n
  );


  buf

  (
    ffc_10_n_spl_0,
    ffc_10_n_spl_
  );


  buf

  (
    ffc_10_p_spl_,
    ffc_10_p
  );


  buf

  (
    g375_n_spl_,
    g375_n
  );


  buf

  (
    g377_n_spl_,
    g377_n
  );


  buf

  (
    ffc_12_n_spl_,
    ffc_12_n
  );


  buf

  (
    g379_n_spl_,
    g379_n
  );


  buf

  (
    g383_n_spl_,
    g383_n
  );


  buf

  (
    g373_n_spl_,
    g373_n
  );


  buf

  (
    ffc_237_n_spl_,
    ffc_237_n
  );


  buf

  (
    ffc_259_n_spl_,
    ffc_259_n
  );


  buf

  (
    ffc_261_n_spl_,
    ffc_261_n
  );


  buf

  (
    ffc_259_p_spl_,
    ffc_259_p
  );


  buf

  (
    ffc_261_p_spl_,
    ffc_261_p
  );


  buf

  (
    ffc_77_p_spl_,
    ffc_77_p
  );


  buf

  (
    ffc_77_p_spl_0,
    ffc_77_p_spl_
  );


  buf

  (
    ffc_77_p_spl_1,
    ffc_77_p_spl_
  );


  buf

  (
    g392_p_spl_,
    g392_p
  );


  buf

  (
    ffc_77_n_spl_,
    ffc_77_n
  );


  buf

  (
    ffc_77_n_spl_0,
    ffc_77_n_spl_
  );


  buf

  (
    ffc_77_n_spl_1,
    ffc_77_n_spl_
  );


  buf

  (
    g392_n_spl_,
    g392_n
  );


  buf

  (
    ffc_262_n_spl_,
    ffc_262_n
  );


  buf

  (
    ffc_263_n_spl_,
    ffc_263_n
  );


  buf

  (
    ffc_262_p_spl_,
    ffc_262_p
  );


  buf

  (
    ffc_263_p_spl_,
    ffc_263_p
  );


  buf

  (
    ffc_81_p_spl_,
    ffc_81_p
  );


  buf

  (
    g398_p_spl_,
    g398_p
  );


  buf

  (
    ffc_81_n_spl_,
    ffc_81_n
  );


  buf

  (
    g398_n_spl_,
    g398_n
  );


  buf

  (
    ffc_264_n_spl_,
    ffc_264_n
  );


  buf

  (
    ffc_265_n_spl_,
    ffc_265_n
  );


  buf

  (
    ffc_264_p_spl_,
    ffc_264_p
  );


  buf

  (
    ffc_265_p_spl_,
    ffc_265_p
  );


  buf

  (
    g407_p_spl_,
    g407_p
  );


  buf

  (
    g407_n_spl_,
    g407_n
  );


  buf

  (
    ffc_267_n_spl_,
    ffc_267_n
  );


  buf

  (
    ffc_269_n_spl_,
    ffc_269_n
  );


  buf

  (
    ffc_267_p_spl_,
    ffc_267_p
  );


  buf

  (
    ffc_269_p_spl_,
    ffc_269_p
  );


  buf

  (
    ffc_119_p_spl_,
    ffc_119_p
  );


  buf

  (
    g413_p_spl_,
    g413_p
  );


  buf

  (
    ffc_119_n_spl_,
    ffc_119_n
  );


  buf

  (
    g413_n_spl_,
    g413_n
  );


  buf

  (
    ffc_135_n_spl_,
    ffc_135_n
  );


  buf

  (
    ffc_135_n_spl_0,
    ffc_135_n_spl_
  );


  buf

  (
    ffc_135_n_spl_00,
    ffc_135_n_spl_0
  );


  buf

  (
    ffc_135_n_spl_01,
    ffc_135_n_spl_0
  );


  buf

  (
    ffc_135_n_spl_1,
    ffc_135_n_spl_
  );


  buf

  (
    ffc_135_n_spl_10,
    ffc_135_n_spl_1
  );


  buf

  (
    ffc_135_n_spl_11,
    ffc_135_n_spl_1
  );


  buf

  (
    ffc_127_n_spl_,
    ffc_127_n
  );


  buf

  (
    ffc_127_n_spl_0,
    ffc_127_n_spl_
  );


  buf

  (
    ffc_127_n_spl_00,
    ffc_127_n_spl_0
  );


  buf

  (
    ffc_127_n_spl_000,
    ffc_127_n_spl_00
  );


  buf

  (
    ffc_127_n_spl_001,
    ffc_127_n_spl_00
  );


  buf

  (
    ffc_127_n_spl_01,
    ffc_127_n_spl_0
  );


  buf

  (
    ffc_127_n_spl_010,
    ffc_127_n_spl_01
  );


  buf

  (
    ffc_127_n_spl_1,
    ffc_127_n_spl_
  );


  buf

  (
    ffc_127_n_spl_10,
    ffc_127_n_spl_1
  );


  buf

  (
    ffc_127_n_spl_11,
    ffc_127_n_spl_1
  );


  buf

  (
    ffc_131_n_spl_,
    ffc_131_n
  );


  buf

  (
    ffc_131_n_spl_0,
    ffc_131_n_spl_
  );


  buf

  (
    ffc_131_n_spl_00,
    ffc_131_n_spl_0
  );


  buf

  (
    ffc_131_n_spl_01,
    ffc_131_n_spl_0
  );


  buf

  (
    ffc_131_n_spl_1,
    ffc_131_n_spl_
  );


  buf

  (
    ffc_131_n_spl_10,
    ffc_131_n_spl_1
  );


  buf

  (
    ffc_131_n_spl_11,
    ffc_131_n_spl_1
  );


  buf

  (
    ffc_139_n_spl_,
    ffc_139_n
  );


  buf

  (
    ffc_139_n_spl_0,
    ffc_139_n_spl_
  );


  buf

  (
    ffc_139_n_spl_00,
    ffc_139_n_spl_0
  );


  buf

  (
    ffc_139_n_spl_01,
    ffc_139_n_spl_0
  );


  buf

  (
    ffc_139_n_spl_1,
    ffc_139_n_spl_
  );


  buf

  (
    ffc_139_n_spl_10,
    ffc_139_n_spl_1
  );


  buf

  (
    ffc_139_n_spl_11,
    ffc_139_n_spl_1
  );


  buf

  (
    ffc_270_n_spl_,
    ffc_270_n
  );


  buf

  (
    ffc_270_n_spl_0,
    ffc_270_n_spl_
  );


  buf

  (
    ffc_270_n_spl_00,
    ffc_270_n_spl_0
  );


  buf

  (
    ffc_270_n_spl_01,
    ffc_270_n_spl_0
  );


  buf

  (
    ffc_270_n_spl_1,
    ffc_270_n_spl_
  );


  buf

  (
    ffc_270_n_spl_10,
    ffc_270_n_spl_1
  );


  buf

  (
    ffc_270_n_spl_11,
    ffc_270_n_spl_1
  );


  buf

  (
    ffc_123_n_spl_,
    ffc_123_n
  );


  buf

  (
    ffc_123_n_spl_0,
    ffc_123_n_spl_
  );


  buf

  (
    ffc_123_n_spl_00,
    ffc_123_n_spl_0
  );


  buf

  (
    ffc_123_n_spl_01,
    ffc_123_n_spl_0
  );


  buf

  (
    ffc_123_n_spl_1,
    ffc_123_n_spl_
  );


  buf

  (
    ffc_123_n_spl_10,
    ffc_123_n_spl_1
  );


  buf

  (
    ffc_143_n_spl_,
    ffc_143_n
  );


  buf

  (
    ffc_171_n_spl_,
    ffc_171_n
  );


  buf

  (
    g450_n_spl_,
    g450_n
  );


  buf

  (
    ffc_93_p_spl_,
    ffc_93_p
  );


  buf

  (
    ffc_260_p_spl_,
    ffc_260_p
  );


  buf

  (
    ffc_93_n_spl_,
    ffc_93_n
  );


  buf

  (
    ffc_93_n_spl_0,
    ffc_93_n_spl_
  );


  buf

  (
    ffc_260_n_spl_,
    ffc_260_n
  );


  buf

  (
    ffc_260_n_spl_0,
    ffc_260_n_spl_
  );


  buf

  (
    ffc_97_n_spl_,
    ffc_97_n
  );


  buf

  (
    ffc_238_n_spl_,
    ffc_238_n
  );


  buf

  (
    ffc_256_n_spl_,
    ffc_256_n
  );


  buf

  (
    ffc_256_n_spl_0,
    ffc_256_n_spl_
  );


  buf

  (
    ffc_266_n_spl_,
    ffc_266_n
  );


  buf

  (
    ffc_256_p_spl_,
    ffc_256_p
  );


  buf

  (
    ffc_266_p_spl_,
    ffc_266_p
  );


  buf

  (
    g483_n_spl_,
    g483_n
  );


  buf

  (
    g483_p_spl_,
    g483_p
  );


  buf

  (
    g482_p_spl_,
    g482_p
  );


  buf

  (
    g485_n_spl_,
    g485_n
  );


  buf

  (
    g481_n_spl_,
    g481_n
  );


  buf

  (
    g481_n_spl_0,
    g481_n_spl_
  );


  buf

  (
    ffc_201_n_spl_,
    ffc_201_n
  );


  buf

  (
    g488_n_spl_,
    g488_n
  );


  buf

  (
    g503_n_spl_,
    g503_n
  );


  buf

  (
    g518_n_spl_,
    g518_n
  );


  buf

  (
    ffc_235_n_spl_,
    ffc_235_n
  );


  buf

  (
    g533_n_spl_,
    g533_n
  );


  buf

  (
    ffc_257_n_spl_,
    ffc_257_n
  );


  buf

  (
    ffc_104_n_spl_,
    ffc_104_n
  );


  buf

  (
    ffc_104_n_spl_0,
    ffc_104_n_spl_
  );


  buf

  (
    g549_p_spl_,
    g549_p
  );


  buf

  (
    g549_p_spl_0,
    g549_p_spl_
  );


  buf

  (
    g548_n_spl_,
    g548_n
  );


  buf

  (
    g550_n_spl_,
    g550_n
  );


  buf

  (
    ffc_62_n_spl_,
    ffc_62_n
  );


  buf

  (
    ffc_100_n_spl_,
    ffc_100_n
  );


  buf

  (
    ffc_100_n_spl_0,
    ffc_100_n_spl_
  );


  buf

  (
    g558_p_spl_,
    g558_p
  );


  buf

  (
    g558_p_spl_0,
    g558_p_spl_
  );


  buf

  (
    g551_p_spl_,
    g551_p
  );


  buf

  (
    g552_p_spl_,
    g552_p
  );


  buf

  (
    g553_n_spl_,
    g553_n
  );


  buf

  (
    ffc_287_n_spl_,
    ffc_287_n
  );


  buf

  (
    g565_p_spl_,
    g565_p
  );


  buf

  (
    g565_p_spl_0,
    g565_p_spl_
  );


  buf

  (
    g563_n_spl_,
    g563_n
  );


  buf

  (
    g564_n_spl_,
    g564_n
  );


  buf

  (
    g559_n_spl_,
    g559_n
  );


  buf

  (
    ffc_58_p_spl_,
    ffc_58_p
  );


  buf

  (
    ffc_58_p_spl_0,
    ffc_58_p_spl_
  );


  buf

  (
    ffc_198_p_spl_,
    ffc_198_p
  );


  buf

  (
    ffc_244_p_spl_,
    ffc_244_p
  );


  buf

  (
    ffc_234_p_spl_,
    ffc_234_p
  );


  buf

  (
    ffc_245_p_spl_,
    ffc_245_p
  );


  buf

  (
    g566_p_spl_,
    g566_p
  );


  buf

  (
    g567_p_spl_,
    g567_p
  );


  buf

  (
    ffc_243_p_spl_,
    ffc_243_p
  );


  buf

  (
    ffc_306_p_spl_,
    ffc_306_p
  );


  buf

  (
    ffc_306_p_spl_0,
    ffc_306_p_spl_
  );


  buf

  (
    ffc_306_p_spl_1,
    ffc_306_p_spl_
  );


  buf

  (
    ffc_305_p_spl_,
    ffc_305_p
  );


  buf

  (
    ffc_307_p_spl_,
    ffc_307_p
  );


  buf

  (
    ffc_110_n_spl_,
    ffc_110_n
  );


  buf

  (
    g582_p_spl_,
    g582_p
  );


  buf

  (
    g582_p_spl_0,
    g582_p_spl_
  );


  buf

  (
    g578_n_spl_,
    g578_n
  );


  buf

  (
    g583_n_spl_,
    g583_n
  );


  buf

  (
    ffc_298_p_spl_,
    ffc_298_p
  );


  buf

  (
    ffc_303_p_spl_,
    ffc_303_p
  );


  buf

  (
    g591_p_spl_,
    g591_p
  );


  buf

  (
    ffc_122_p_spl_,
    ffc_122_p
  );


  buf

  (
    ffc_233_p_spl_,
    ffc_233_p
  );


  buf

  (
    ffc_96_p_spl_,
    ffc_96_p
  );


  buf

  (
    ffc_96_p_spl_0,
    ffc_96_p_spl_
  );


  buf

  (
    g577_n_spl_,
    g577_n
  );


  buf

  (
    ffc_142_p_spl_,
    ffc_142_p
  );


  buf

  (
    ffc_54_p_spl_,
    ffc_54_p
  );


  buf

  (
    ffc_54_p_spl_0,
    ffc_54_p_spl_
  );


  buf

  (
    ffc_180_p_spl_,
    ffc_180_p
  );


  buf

  (
    ffc_62_p_spl_,
    ffc_62_p
  );


  buf

  (
    ffc_254_p_spl_,
    ffc_254_p
  );


  buf

  (
    ffc_209_p_spl_,
    ffc_209_p
  );


  buf

  (
    ffc_200_p_spl_,
    ffc_200_p
  );


  buf

  (
    ffc_92_p_spl_,
    ffc_92_p
  );


  buf

  (
    ffc_100_p_spl_,
    ffc_100_p
  );


  buf

  (
    ffc_104_p_spl_,
    ffc_104_p
  );


  buf

  (
    g560_p_spl_,
    g560_p
  );


  buf

  (
    g562_p_spl_,
    g562_p
  );


  buf

  (
    g568_n_spl_,
    g568_n
  );


  buf

  (
    ffc_236_p_spl_,
    ffc_236_p
  );


  buf

  (
    ffc_257_p_spl_,
    ffc_257_p
  );


  buf

  (
    ffc_202_p_spl_,
    ffc_202_p
  );


  buf

  (
    ffc_211_p_spl_,
    ffc_211_p
  );


  buf

  (
    g571_n_spl_,
    g571_n
  );


  buf

  (
    ffc_68_p_spl_,
    ffc_68_p
  );


  buf

  (
    ffc_252_p_spl_,
    ffc_252_p
  );


  buf

  (
    ffc_252_p_spl_0,
    ffc_252_p_spl_
  );


  buf

  (
    ffc_85_p_spl_,
    ffc_85_p
  );


  buf

  (
    ffc_83_p_spl_,
    ffc_83_p
  );


  buf

  (
    ffc_217_p_spl_,
    ffc_217_p
  );


  buf

  (
    ffc_65_p_spl_,
    ffc_65_p
  );


  buf

  (
    ffc_107_p_spl_,
    ffc_107_p
  );


  buf

  (
    g644_n_spl_,
    g644_n
  );


  buf

  (
    g585_n_spl_,
    g585_n
  );


  buf

  (
    g587_n_spl_,
    g587_n
  );


  buf

  (
    g592_n_spl_,
    g592_n
  );


  buf

  (
    g593_p_spl_,
    g593_p
  );


  buf

  (
    g634_p_spl_,
    g634_p
  );


  buf

  (
    ffc_73_p_spl_,
    ffc_73_p
  );


  buf

  (
    g599_n_spl_,
    g599_n
  );


  buf

  (
    g599_n_spl_0,
    g599_n_spl_
  );


  buf

  (
    ffc_299_p_spl_,
    ffc_299_p
  );


  buf

  (
    g589_n_spl_,
    g589_n
  );


  buf

  (
    g589_n_spl_0,
    g589_n_spl_
  );


  buf

  (
    g601_p_spl_,
    g601_p
  );


  buf

  (
    g601_p_spl_0,
    g601_p_spl_
  );


  buf

  (
    ffc_71_p_spl_,
    ffc_71_p
  );


  buf

  (
    ffc_87_p_spl_,
    ffc_87_p
  );


  buf

  (
    ffc_114_p_spl_,
    ffc_114_p
  );


  buf

  (
    g657_n_spl_,
    g657_n
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    g663_n_spl_,
    g663_n
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    g662_n_spl_,
    g662_n
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


endmodule
