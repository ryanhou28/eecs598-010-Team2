// Benchmark "c2670" written by ABC on Sun Oct 29 19:31:53 2023

module c2670 (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58,
    G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70, G71, G72,
    G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86,
    G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G109, G110, G111, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G124,
    G125, G126, G127, G128, G129, G130, G131, G132, G133, G134, G135, G136,
    G137, G138, G139, G140, G141, G142, G143, G144, G145, G146, G147, G148,
    G149, G150, G151, G152, G153, G154, G155, G156, G157,
    G2531, G2532, G2533, G2534, G2535, G2536, G2537, G2538, G2539, G2540,
    G2541, G2542, G2543, G2544, G2545, G2546, G2547, G2548, G2549, G2550,
    G2551, G2552, G2553, G2554, G2555, G2556, G2557, G2558, G2559, G2560,
    G2561, G2562, G2563, G2564, G2565, G2566, G2567, G2568, G2569, G2570,
    G2571, G2572, G2573, G2574, G2575, G2576, G2577, G2578, G2579, G2580,
    G2581, G2582, G2583, G2584, G2585, G2586, G2587, G2588, G2589, G2590,
    G2591, G2592, G2593, G2594  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70,
    G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98,
    G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G110,
    G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G133, G134,
    G135, G136, G137, G138, G139, G140, G141, G142, G143, G144, G145, G146,
    G147, G148, G149, G150, G151, G152, G153, G154, G155, G156, G157;
  output G2531, G2532, G2533, G2534, G2535, G2536, G2537, G2538, G2539, G2540,
    G2541, G2542, G2543, G2544, G2545, G2546, G2547, G2548, G2549, G2550,
    G2551, G2552, G2553, G2554, G2555, G2556, G2557, G2558, G2559, G2560,
    G2561, G2562, G2563, G2564, G2565, G2566, G2567, G2568, G2569, G2570,
    G2571, G2572, G2573, G2574, G2575, G2576, G2577, G2578, G2579, G2580,
    G2581, G2582, G2583, G2584, G2585, G2586, G2587, G2588, G2589, G2590,
    G2591, G2592, G2593, G2594;
  reg n1416_lo, n1419_lo, n1422_lo, n1425_lo, n1428_lo, n1431_lo, n1434_lo,
    n1437_lo, n1440_lo, n1443_lo, n1446_lo, n1449_lo, n1452_lo, n1455_lo,
    n1458_lo, n1461_lo, n1464_lo, n1467_lo, n1470_lo, n1473_lo, n1476_lo,
    n1479_lo, n1482_lo, n1485_lo, n1488_lo, n1491_lo, n1494_lo, n1497_lo,
    n1500_lo, n1503_lo, n1506_lo, n1509_lo, n1512_lo, n1515_lo, n1518_lo,
    n1521_lo, n1524_lo, n1527_lo, n1530_lo, n1533_lo, n1536_lo, n1539_lo,
    n1542_lo, n1545_lo, n1548_lo, n1551_lo, n1554_lo, n1557_lo, n1560_lo,
    n1563_lo, n1566_lo, n1569_lo, n1572_lo, n1575_lo, n1578_lo, n1581_lo,
    n1584_lo, n1587_lo, n1590_lo, n1593_lo, n1596_lo, n1599_lo, n1602_lo,
    n1605_lo, n1608_lo, n1611_lo, n1614_lo, n1617_lo, n1620_lo, n1623_lo,
    n1626_lo, n1629_lo, n1632_lo, n1635_lo, n1638_lo, n1641_lo, n1644_lo,
    n1647_lo, n1650_lo, n1653_lo, n1656_lo, n1659_lo, n1662_lo, n1665_lo,
    n1668_lo, n1671_lo, n1674_lo, n1677_lo, n1680_lo, n1683_lo, n1686_lo,
    n1689_lo, n1692_lo, n1695_lo, n1698_lo, n1701_lo, n1704_lo, n1707_lo,
    n1710_lo, n1713_lo, n1716_lo, n1719_lo, n1722_lo, n1725_lo, n1728_lo,
    n1731_lo, n1734_lo, n1737_lo, n1740_lo, n1743_lo, n1746_lo, n1749_lo,
    n1752_lo, n1755_lo, n1758_lo, n1761_lo, n1764_lo, n1767_lo, n1770_lo,
    n1773_lo, n1776_lo, n1779_lo, n1782_lo, n1785_lo, n1788_lo, n1791_lo,
    n1794_lo, n1797_lo, n1800_lo, n1803_lo, n1806_lo, n1809_lo, n1812_lo,
    n1815_lo, n1818_lo, n1821_lo, n1824_lo, n1827_lo, n1830_lo, n1833_lo,
    n1836_lo, n1839_lo, n1842_lo, n1845_lo, n1848_lo, n1851_lo, n1854_lo,
    n1857_lo, n1860_lo, n1863_lo, n1866_lo, n1869_lo, n1872_lo, n1875_lo,
    n1878_lo, n1881_lo, n1884_lo, n1887_lo, n1890_lo, n1893_lo, n1896_lo,
    n1899_lo, n1902_lo, n1905_lo, n1908_lo, n1911_lo, n1914_lo, n1917_lo,
    n1920_lo, n1923_lo, n1926_lo, n1929_lo, n1932_lo, n1935_lo, n1938_lo,
    n1941_lo, n1944_lo, n1947_lo, n1950_lo, n1953_lo, n1956_lo, n1959_lo,
    n1962_lo, n1965_lo, n1968_lo, n1971_lo, n1974_lo, n1977_lo, n1980_lo,
    n1983_lo, n1986_lo, n1989_lo, n1992_lo, n1995_lo, n1998_lo, n2001_lo,
    n2004_lo, n2007_lo, n2010_lo, n2013_lo, n2016_lo, n2019_lo, n2022_lo,
    n2025_lo, n2028_lo, n2031_lo, n2034_lo, n2037_lo, n2040_lo, n2043_lo,
    n2046_lo, n2049_lo, n2052_lo, n2055_lo, n2058_lo, n2061_lo, n2064_lo,
    n2067_lo, n2070_lo, n2073_lo, n2076_lo, n2079_lo, n2082_lo, n2085_lo,
    n2088_lo, n2091_lo, n2094_lo, n2097_lo, n2100_lo, n2103_lo, n2106_lo,
    n2109_lo, n2112_lo, n2115_lo, n2118_lo, n2121_lo, n2124_lo, n2127_lo,
    n2130_lo, n2133_lo, n2136_lo, n2139_lo, n2142_lo, n2145_lo, n2148_lo,
    n2151_lo, n2154_lo, n2157_lo, n2160_lo, n2163_lo, n2166_lo, n2169_lo,
    n2172_lo, n2175_lo, n2178_lo, n2181_lo, n2184_lo, n2187_lo, n2190_lo,
    n2193_lo, n2196_lo, n2199_lo, n2202_lo, n2205_lo, n2208_lo, n2211_lo,
    n2214_lo, n2217_lo, n2220_lo, n2223_lo, n2226_lo, n2229_lo, n2232_lo,
    n2235_lo, n2238_lo, n2241_lo, n2244_lo, n2247_lo, n2250_lo, n2253_lo,
    n2256_lo, n2259_lo, n2262_lo, n2265_lo, n2268_lo, n2271_lo, n2274_lo,
    n2277_lo, n2280_lo, n2283_lo, n2286_lo, n2289_lo, n2292_lo, n2295_lo,
    n2298_lo, n2301_lo, n2304_lo, n2307_lo, n2310_lo, n2313_lo, n2316_lo,
    n2319_lo, n2322_lo, n2325_lo, n2328_lo, n2331_lo, n2334_lo, n2337_lo,
    n2340_lo, n2343_lo, n2346_lo, n2349_lo, n2352_lo, n2355_lo, n2358_lo,
    n2361_lo, n2364_lo, n2367_lo, n2370_lo, n2373_lo, n2376_lo, n2379_lo,
    n2382_lo, n2385_lo, n2388_lo, n2391_lo, n2394_lo, n2397_lo, n2400_lo,
    n2403_lo, n2406_lo, n2409_lo, n2412_lo, n2415_lo, n2418_lo, n2421_lo,
    n2424_lo, n2427_lo, n2430_lo, n2433_lo, n2436_lo, n2439_lo, n2442_lo,
    n2445_lo, n2448_lo, n2451_lo, n2454_lo, n2457_lo, n2460_lo, n2463_lo,
    n2466_lo, n2469_lo, n2472_lo, n2475_lo, n2478_lo, n2481_lo, n2484_lo,
    n2487_lo, n2490_lo, n2493_lo, n2496_lo, n2499_lo, n2502_lo, n2505_lo,
    n2508_lo, n2511_lo, n2514_lo, n2517_lo, n2520_lo, n2523_lo, n2526_lo,
    n2529_lo, n2532_lo, n2535_lo, n2538_lo, n2541_lo, n2544_lo, n2547_lo,
    n2550_lo, n2553_lo, n2556_lo, n2559_lo, n2562_lo, n2565_lo, n2568_lo,
    n2571_lo, n2574_lo, n2577_lo, n2580_lo, n2583_lo, n2586_lo, n2589_lo,
    n2592_lo, n2595_lo, n2598_lo, n2601_lo, n2604_lo, n2607_lo, n2610_lo,
    n2613_lo, n2616_lo, n2619_lo, n2622_lo, n2625_lo, n2628_lo, n2631_lo,
    n2634_lo, n2637_lo, n2640_lo, n2643_lo, n2646_lo, n2649_lo, n2652_lo,
    n2655_lo, n2658_lo, n2661_lo, n2664_lo, n2667_lo, n2670_lo, n2673_lo,
    n2676_lo, n2679_lo, n2682_lo, n2685_lo, n2688_lo, n2691_lo, n2694_lo,
    n2697_lo, n2700_lo, n2703_lo, n2706_lo, n2709_lo, n2712_lo, n2715_lo,
    n2718_lo, n2721_lo, n2724_lo, n2727_lo, n2730_lo, n2733_lo, n2736_lo,
    n2739_lo, n2742_lo, n2745_lo, n2748_lo, n2751_lo, n2754_lo, n2757_lo,
    n2760_lo, n2763_lo, n2766_lo, n2769_lo, n2772_lo, n2775_lo, n2778_lo,
    n2781_lo, n2784_lo, n2787_lo, n2790_lo, n2793_lo, n2796_lo, n2799_lo,
    n2802_lo, n2805_lo, n2808_lo, n2811_lo, n2814_lo, n2817_lo, n2820_lo,
    n2823_lo, n2826_lo, n2829_lo, n2832_lo, n2835_lo, n2838_lo, n2841_lo,
    n2844_lo, n2847_lo, n2850_lo, n2853_lo, n2856_lo, n2859_lo, n2862_lo,
    n2865_lo, n2868_lo, n2871_lo, n2874_lo, n2877_lo, n2880_lo, n2883_lo,
    n2886_lo, n2889_lo, n2892_lo, n2895_lo, n2898_lo, n2901_lo, n2904_lo,
    n2907_lo, n2910_lo, n2913_lo, n2916_lo, n2919_lo, n2922_lo, n2925_lo,
    n2928_lo, n2931_lo, n2934_lo, n2937_lo, n2940_lo, n2943_lo, n2946_lo,
    n2949_lo, n2952_lo, n2955_lo, n2958_lo, n2961_lo, n2964_lo, n2967_lo,
    n2970_lo, n2973_lo, n2976_lo, n2979_lo, n2982_lo, n2985_lo, n2988_lo,
    n2991_lo, n2994_lo, n2997_lo, n3000_lo, n3003_lo, n3006_lo, n3009_lo,
    n3012_lo, n3015_lo, n3018_lo, n3021_lo, n3024_lo, n3027_lo, n3030_lo,
    n3033_lo, n3036_lo, n3039_lo, n3042_lo, n3045_lo, n3048_lo, n3051_lo,
    n3054_lo, n3057_lo, n3060_lo, n3063_lo, n3066_lo, n3069_lo, n3072_lo,
    n3075_lo, n3078_lo, n3081_lo, n3084_lo, n3087_lo, n3090_lo, n3093_lo,
    n3096_lo, n3099_lo, n3102_lo, n3105_lo, n3108_lo, n3111_lo, n3114_lo,
    n3117_lo, n3120_lo, n3123_lo, n3126_lo, n3129_lo, n3132_lo, n3135_lo,
    n3138_lo, n3141_lo, n3144_lo, n3147_lo, n3150_lo, n3153_lo, n3156_lo,
    n3159_lo, n3162_lo, n3165_lo, n3168_lo, n3171_lo, n3174_lo, n3177_lo,
    n3180_lo, n3183_lo, n3186_lo, n3189_lo, n3192_lo, n3195_lo, n3198_lo,
    n3201_lo, n3204_lo, n3207_lo, n3210_lo, n3213_lo, n3216_lo, n3219_lo,
    n3222_lo, n3225_lo, n3228_lo, n3231_lo, n3234_lo, n3237_lo, n3240_lo,
    n3243_lo, n3246_lo, n3249_lo, n3252_lo, n3255_lo, n3258_lo, n3261_lo,
    n3264_lo, n3267_lo, n3270_lo, n3273_lo, n3276_lo, n3279_lo, n3282_lo,
    n3285_lo, n3288_lo, n3291_lo, n3294_lo, n3297_lo;
  wire new_G282_, new_G283_, new_G284_, new_G285_, new_G286_, new_G287_,
    new_G288_, new_G291_, new_G292_, new_G295_, new_G298_, new_G301_,
    new_G313_, new_G325_, new_G329_, new_G335_, new_G336_, new_G339_,
    new_G342_, new_G354_, new_G366_, new_G370_, new_G374_, new_G386_,
    new_G398_, new_G399_, new_G400_, new_G401_, new_G402_, new_G403_,
    new_G404_, new_G405_, new_G417_, new_G429_, new_G435_, new_G442_,
    new_G443_, new_G447_, new_G451_, new_G455_, new_G459_, new_G463_,
    new_G467_, new_G471_, new_G475_, new_G479_, new_G485_, new_G491_,
    new_G497_, new_G503_, new_G507_, new_G511_, new_G515_, new_G519_,
    new_G522_, new_G525_, new_G526_, new_G527_, new_G530_, new_G533_,
    new_G536_, new_G539_, new_G542_, new_G545_, new_G548_, new_G551_,
    new_G554_, new_G557_, new_G560_, new_G563_, new_G566_, new_G569_,
    new_G572_, new_G575_, new_G578_, new_G581_, new_G584_, new_G585_,
    new_G586_, new_G587_, new_G588_, new_G589_, new_G590_, new_G591_,
    new_G592_, new_G593_, new_G594_, new_G595_, new_G598_, new_G603_,
    new_G614_, new_G625_, new_G626_, new_G627_, new_G628_, new_G629_,
    new_G630_, new_G631_, new_G636_, new_G647_, new_G658_, new_G659_,
    new_G660_, new_G661_, new_G662_, new_G663_, new_G674_, new_G685_,
    new_G686_, new_G687_, new_G688_, new_G689_, new_G690_, new_G694_,
    new_G698_, new_G701_, new_G702_, new_G703_, new_G704_, new_G705_,
    new_G706_, new_G707_, new_G718_, new_G729_, new_G730_, new_G731_,
    new_G732_, new_G733_, new_G734_, new_G739_, new_G745_, new_G746_,
    new_G747_, new_G748_, new_G749_, new_G750_, new_G751_, new_G756_,
    new_G761_, new_G766_, new_G771_, new_G772_, new_G773_, new_G774_,
    new_G775_, new_G776_, new_G777_, new_G780_, new_G783_, new_G786_,
    new_G789_, new_G792_, new_G795_, new_G798_, new_G801_, new_G804_,
    new_G807_, new_G810_, new_G811_, new_G812_, new_G815_, new_G818_,
    new_G821_, new_G824_, new_G827_, new_G830_, new_G831_, new_G832_,
    new_G833_, new_G834_, new_G835_, new_G836_, new_G837_, new_G838_,
    new_G839_, new_G840_, new_G841_, new_G842_, new_G843_, new_G844_,
    new_G845_, new_G846_, new_G847_, new_G848_, new_G849_, new_G850_,
    new_G851_, new_G852_, new_G853_, new_G854_, new_G855_, new_G856_,
    new_G857_, new_G858_, new_G859_, new_G860_, new_G861_, new_G862_,
    new_G863_, new_G864_, new_G865_, new_G866_, new_G867_, new_G868_,
    new_G869_, new_G870_, new_G871_, new_G872_, new_G873_, new_G874_,
    new_G875_, new_G876_, new_G877_, new_G878_, new_G879_, new_G880_,
    new_G881_, new_G882_, new_G883_, new_G884_, new_G885_, new_G886_,
    new_G887_, new_G888_, new_G889_, new_G890_, new_G891_, new_G892_,
    new_G893_, new_G894_, new_G895_, new_G896_, new_G897_, new_G898_,
    new_G901_, new_G904_, new_G908_, new_G912_, new_G915_, new_G918_,
    new_G921_, new_G922_, new_G923_, new_G924_, new_G925_, new_G926_,
    new_G927_, new_G928_, new_G929_, new_G930_, new_G931_, new_G932_,
    new_G933_, new_G934_, new_G935_, new_G936_, new_G937_, new_G938_,
    new_G939_, new_G940_, new_G941_, new_G942_, new_G943_, new_G944_,
    new_G945_, new_G946_, new_G947_, new_G948_, new_G949_, new_G950_,
    new_G951_, new_G952_, new_G953_, new_G954_, new_G955_, new_G959_,
    new_G963_, new_G966_, new_G967_, new_G968_, new_G969_, new_G970_,
    new_G971_, new_G972_, new_G973_, new_G974_, new_G975_, new_G976_,
    new_G977_, new_G978_, new_G979_, new_G980_, new_G983_, new_G984_,
    new_G987_, new_G990_, new_G993_, new_G998_, new_G1002_, new_G1008_,
    new_G1014_, new_G1017_, new_G1021_, new_G1026_, new_G1030_, new_G1033_,
    new_G1036_, new_G1039_, new_G1044_, new_G1049_, new_G1053_, new_G1058_,
    new_G1062_, new_G1067_, new_G1072_, new_G1076_, new_G1079_, new_G1082_,
    new_G1085_, new_G1088_, new_G1089_, new_G1090_, new_G1093_, new_G1096_,
    new_G1097_, new_G1098_, new_G1101_, new_G1104_, new_G1107_, new_G1110_,
    new_G1111_, new_G1112_, new_G1113_, new_G1114_, new_G1115_, new_G1116_,
    new_G1117_, new_G1118_, new_G1119_, new_G1120_, new_G1123_, new_G1126_,
    new_G1127_, new_G1128_, new_G1129_, new_G1132_, new_G1137_, new_G1144_,
    new_G1148_, new_G1152_, new_G1159_, new_G1166_, new_G1171_, new_G1176_,
    new_G1181_, new_G1184_, new_G1187_, new_G1190_, new_G1193_, new_G1196_,
    new_G1197_, new_G1198_, new_G1199_, new_G1200_, new_G1201_, new_G1202_,
    new_G1203_, new_G1204_, new_G1205_, new_G1206_, new_G1207_, new_G1208_,
    new_G1209_, new_G1210_, new_G1211_, new_G1212_, new_G1213_, new_G1214_,
    new_G1215_, new_G1216_, new_G1219_, new_G1220_, new_G1221_, new_G1222_,
    new_G1225_, new_G1228_, new_G1231_, new_G1234_, new_G1237_, new_G1240_,
    new_G1243_, new_G1246_, new_G1249_, new_G1250_, new_G1251_, new_G1252_,
    new_G1253_, new_G1254_, new_G1255_, new_G1256_, new_G1257_, new_G1258_,
    new_G1259_, new_G1260_, new_G1263_, new_G1266_, new_G1269_, new_G1272_,
    new_G1275_, new_G1278_, new_G1281_, new_G1284_, new_G1287_, new_G1290_,
    new_G1293_, new_G1296_, new_G1299_, new_G1302_, new_G1305_, new_G1308_,
    new_G1311_, new_G1314_, new_G1320_, new_G1321_, new_G1326_, new_G1327_,
    new_G1328_, new_G1329_, new_G1336_, new_G1342_, new_G1345_, new_G1348_,
    new_G1351_, new_G1354_, new_G1355_, new_G1356_, new_G1357_, new_G1358_,
    new_G1359_, new_G1360_, new_G1361_, new_G1362_, new_G1363_, new_G1364_,
    new_G1365_, new_G1366_, new_G1367_, new_G1368_, new_G1371_, new_G1374_,
    new_G1377_, new_G1380_, new_G1383_, new_G1384_, new_G1387_, new_G1390_,
    new_G1393_, new_G1396_, new_G1399_, new_G1402_, new_G1405_, new_G1406_,
    new_G1407_, new_G1408_, new_G1409_, new_G1412_, new_G1415_, new_G1418_,
    new_G1421_, new_G1424_, new_G1425_, new_G1426_, new_G1427_, new_G1428_,
    new_G1429_, new_G1430_, new_G1431_, new_G1432_, new_G1433_, new_G1434_,
    new_G1435_, new_G1436_, new_G1437_, new_G1438_, new_G1439_, new_G1440_,
    new_G1441_, new_G1442_, new_G1443_, new_G1444_, new_G1445_, new_G1446_,
    new_G1447_, new_G1448_, new_G1449_, new_G1450_, new_G1451_, new_G1452_,
    new_G1453_, new_G1454_, new_G1455_, new_G1456_, new_G1457_, new_G1458_,
    new_G1459_, new_G1460_, new_G1461_, new_G1462_, new_G1463_, new_G1464_,
    new_G1465_, new_G1466_, new_G1467_, new_G1468_, new_G1469_, new_G1470_,
    new_G1471_, new_G1472_, new_G1475_, new_G1476_, new_G1477_, new_G1478_,
    new_G1479_, new_G1483_, new_G1484_, new_G1485_, new_G1486_, new_G1487_,
    new_G1488_, new_G1493_, new_G1497_, new_G1498_, new_G1502_, new_G1507_,
    new_G1508_, new_G1509_, new_G1510_, new_G1511_, new_G1512_, new_G1513_,
    new_G1514_, new_G1515_, new_G1516_, new_G1517_, new_G1518_, new_G1519_,
    new_G1520_, new_G1524_, new_G1528_, new_G1531_, new_G1532_, new_G1533_,
    new_G1534_, new_G1535_, new_G1536_, new_G1537_, new_G1540_, new_G1543_,
    new_G1546_, new_G1549_, new_G1552_, new_G1555_, new_G1556_, new_G1557_,
    new_G1560_, new_G1563_, new_G1566_, new_G1569_, new_G1572_, new_G1575_,
    new_G1578_, new_G1581_, new_G1584_, new_G1587_, new_G1590_, new_G1593_,
    new_G1596_, new_G1599_, new_G1600_, new_G1601_, new_G1602_, new_G1603_,
    new_G1606_, new_G1607_, new_G1610_, new_G1613_, new_G1616_, new_G1619_,
    new_G1620_, new_G1621_, new_G1622_, new_G1623_, new_G1624_, new_G1625_,
    new_G1626_, new_G1627_, new_G1628_, new_G1629_, new_G1630_, new_G1631_,
    new_G1632_, new_G1633_, new_G1634_, new_G1635_, new_G1636_, new_G1640_,
    new_G1641_, new_G1642_, new_G1643_, new_G1644_, new_G1645_, new_G1646_,
    new_G1650_, new_G1651_, new_G1652_, new_G1653_, new_G1654_, new_G1657_,
    new_G1661_, new_G1662_, new_G1663_, new_G1664_, new_G1665_, new_G1666_,
    new_G1667_, new_G1668_, new_G1669_, new_G1670_, new_G1675_, new_G1676_,
    new_G1681_, new_G1682_, new_G1683_, new_G1684_, new_G1688_, new_G1689_,
    new_G1690_, new_G1691_, new_G1692_, new_G1693_, new_G1694_, new_G1695_,
    new_G1696_, new_G1697_, new_G1698_, new_G1699_, new_G1700_, new_G1701_,
    new_G1702_, new_G1703_, new_G1704_, new_G1705_, new_G1706_, new_G1709_,
    new_G1712_, new_G1715_, new_G1718_, new_G1719_, new_G1720_, new_G1721_,
    new_G1722_, new_G1723_, new_G1724_, new_G1725_, new_G1726_, new_G1727_,
    new_G1728_, new_G1731_, new_G1732_, new_G1733_, new_G1734_, new_G1735_,
    new_G1736_, new_G1737_, new_G1738_, new_G1739_, new_G1744_, new_G1749_,
    new_G1750_, new_G1751_, new_G1752_, new_G1753_, new_G1754_, new_G1755_,
    new_G1756_, new_G1761_, new_G1766_, new_G1767_, new_G1768_, new_G1769_,
    new_G1770_, new_G1771_, new_G1772_, new_G1773_, new_G1774_, new_G1775_,
    new_G1776_, new_G1777_, new_G1778_, new_G1779_, new_G1780_, new_G1781_,
    new_G1782_, new_G1785_, new_G1789_, new_G1792_, new_G1795_, new_G1798_,
    new_G1799_, new_G1800_, new_G1801_, new_G1802_, new_G1805_, new_G1811_,
    new_G1814_, new_G1815_, new_G1816_, new_G1822_, new_G1823_, new_G1824_,
    new_G1825_, new_G1826_, new_G1829_, new_G1835_, new_G1840_, new_G1846_,
    new_G1851_, new_G1854_, new_G1857_, new_G1858_, new_G1859_, new_G1862_,
    new_G1865_, new_G1868_, new_G1869_, new_G1870_, new_G1871_, new_G1872_,
    new_G1873_, new_G1874_, new_G1875_, new_G1876_, new_G1877_, new_G1878_,
    new_G1879_, new_G1880_, new_G1881_, new_G1882_, new_G1883_, new_G1884_,
    new_G1887_, new_G1888_, new_G1889_, new_G1890_, new_G1893_, new_G1896_,
    new_G1899_, new_G1902_, new_G1903_, new_G1904_, new_G1907_, new_G1910_,
    new_G1913_, new_G1916_, new_G1919_, new_G1922_, new_G1925_, new_G1926_,
    new_G1927_, new_G1928_, new_G1931_, new_G1934_, new_G1937_, new_G1940_,
    new_G1943_, new_G1946_, new_G1947_, new_G1948_, new_G1953_, new_G1954_,
    new_G1955_, new_G1956_, new_G1961_, new_G1962_, new_G1963_, new_G1964_,
    new_G1965_, new_G1966_, new_G1967_, new_G1970_, new_G1971_, new_G1972_,
    new_G1973_, new_G1974_, new_G1975_, new_G1976_, new_G1977_, new_G1978_,
    new_G1981_, new_G1982_, new_G1983_, new_G1984_, new_G1985_, new_G1986_,
    new_G1987_, new_G1988_, new_G1989_, new_G1990_, new_G1991_, new_G1992_,
    new_G1993_, new_G1996_, new_G1999_, new_G2002_, new_G2005_, new_G2008_,
    new_G2011_, new_G2014_, new_G2017_, new_G2020_, new_G2023_, new_G2026_,
    new_G2029_, new_G2032_, new_G2035_, new_G2038_, new_G2041_, new_G2044_,
    new_G2045_, new_G2046_, new_G2047_, new_G2048_, new_G2051_, new_G2052_,
    new_G2053_, new_G2054_, new_G2055_, new_G2056_, new_G2057_, new_G2058_,
    new_G2059_, new_G2060_, new_G2061_, new_G2062_, new_G2063_, new_G2064_,
    new_G2065_, new_G2066_, new_G2067_, new_G2068_, new_G2069_, new_G2070_,
    new_G2071_, new_G2072_, new_G2073_, new_G2076_, new_G2079_, new_G2082_,
    new_G2085_, new_G2088_, new_G2091_, new_G2094_, new_G2097_, new_G2100_,
    new_G2103_, new_G2106_, new_G2109_, new_G2112_, new_G2115_, new_G2116_,
    new_G2117_, new_G2118_, new_G2119_, new_G2120_, new_G2121_, new_G2122_,
    new_G2123_, new_G2124_, new_G2125_, new_G2126_, new_G2127_, new_G2128_,
    new_G2129_, new_G2130_, new_G2131_, new_G2132_, new_G2133_, new_G2134_,
    new_G2135_, new_G2138_, new_G2141_, new_G2144_, new_G2147_, new_G2150_,
    new_G2153_, new_G2154_, new_G2155_, new_G2156_, new_G2157_, new_G2158_,
    new_G2161_, new_G2164_, new_G2167_, new_G2170_, new_G2173_, new_G2176_,
    new_G2179_, new_G2182_, new_G2185_, new_G2188_, new_G2191_, new_G2194_,
    new_G2197_, new_G2200_, new_G2203_, new_G2206_, new_G2207_, new_G2208_,
    new_G2209_, new_G2210_, new_G2211_, new_G2212_, new_G2213_, new_G2214_,
    new_G2215_, new_G2216_, new_G2217_, new_G2218_, new_G2219_, new_G2220_,
    new_G2221_, new_G2222_, new_G2223_, new_G2224_, new_G2225_, new_G2226_,
    new_G2227_, new_G2228_, new_G2231_, new_G2234_, new_G2237_, new_G2240_,
    new_G2241_, new_G2242_, new_G2243_, new_G2244_, new_G2245_, new_G2246_,
    new_G2247_, new_G2248_, new_G2249_, new_G2250_, new_G2251_, new_G2252_,
    new_G2253_, new_G2254_, new_G2255_, new_G2256_, new_G2257_, new_G2258_,
    new_G2259_, new_G2260_, new_G2261_, new_G2262_, new_G2263_, new_G2264_,
    new_G2265_, new_G2266_, new_G2267_, new_G2268_, new_G2269_, new_G2270_,
    new_G2271_, new_G2272_, new_G2273_, new_G2274_, new_G2275_, new_G2276_,
    new_G2279_, new_G2282_, new_G2285_, new_G2288_, new_G2291_, new_G2294_,
    new_G2297_, new_G2300_, new_G2301_, new_G2302_, new_G2303_, new_G2304_,
    new_G2305_, new_G2306_, new_G2307_, new_G2308_, new_G2309_, new_G2310_,
    new_G2311_, new_G2312_, new_G2313_, new_G2314_, new_G2315_, new_G2316_,
    new_G2317_, new_G2320_, new_G2323_, new_G2326_, new_G2329_, new_G2330_,
    new_G2331_, new_G2332_, new_G2333_, new_G2334_, new_G2335_, new_G2336_,
    new_G2337_, new_G2340_, new_G2345_, new_G2349_, new_G2352_, new_G2353_,
    new_G2359_, new_G2364_, new_G2365_, new_G2366_, new_G2367_, new_G2368_,
    new_G2369_, new_G2370_, new_G2375_, new_G2379_, new_G2382_, new_G2383_,
    new_G2389_, new_G2394_, new_G2395_, new_G2396_, new_G2397_, new_G2398_,
    new_G2399_, new_G2400_, new_G2401_, new_G2402_, new_G2403_, new_G2404_,
    new_G2405_, new_G2406_, new_G2407_, new_G2408_, new_G2409_, new_G2410_,
    new_G2411_, new_G2412_, new_G2413_, new_G2414_, new_G2417_, new_G2418_,
    new_G2419_, new_G2420_, new_G2421_, new_G2422_, new_G2423_, new_G2424_,
    new_G2425_, new_G2426_, new_G2427_, new_G2428_, new_G2431_, new_G2432_,
    new_G2433_, new_G2434_, new_G2435_, new_G2436_, new_G2437_, new_G2438_,
    new_G2439_, new_G2440_, new_G2441_, new_G2442_, new_G2443_, new_G2447_,
    new_G2450_, new_G2451_, new_G2454_, new_G2458_, new_G2461_, new_G2462_,
    new_G2465_, new_G2466_, new_G2467_, new_G2470_, new_G2473_, new_G2474_,
    new_G2475_, new_G2476_, new_G2477_, new_G2478_, new_G2479_, new_G2480_,
    new_G2481_, new_G2482_, new_G2483_, new_G2484_, new_G2485_, new_G2486_,
    new_G2487_, new_G2488_, new_G2489_, new_G2490_, new_G2491_, new_G2492_,
    new_G2495_, new_G2496_, new_G2499_, new_G2500_, new_G2501_, new_G2502_,
    new_G2503_, new_G2504_, new_G2505_, new_G2508_, new_G2512_, new_G2515_,
    new_G2516_, new_G2517_, new_G2520_, new_G2523_, new_G2524_, new_G2527_,
    new_G2528_, n1416_li, n1419_li, n1422_li, n1425_li, n1428_li, n1431_li,
    n1434_li, n1437_li, n1440_li, n1443_li, n1446_li, n1449_li, n1452_li,
    n1455_li, n1458_li, n1461_li, n1464_li, n1467_li, n1470_li, n1473_li,
    n1476_li, n1479_li, n1482_li, n1485_li, n1488_li, n1491_li, n1494_li,
    n1497_li, n1500_li, n1503_li, n1506_li, n1509_li, n1512_li, n1515_li,
    n1518_li, n1521_li, n1524_li, n1527_li, n1530_li, n1533_li, n1536_li,
    n1539_li, n1542_li, n1545_li, n1548_li, n1551_li, n1554_li, n1557_li,
    n1560_li, n1563_li, n1566_li, n1569_li, n1572_li, n1575_li, n1578_li,
    n1581_li, n1584_li, n1587_li, n1590_li, n1593_li, n1596_li, n1599_li,
    n1602_li, n1605_li, n1608_li, n1611_li, n1614_li, n1617_li, n1620_li,
    n1623_li, n1626_li, n1629_li, n1632_li, n1635_li, n1638_li, n1641_li,
    n1644_li, n1647_li, n1650_li, n1653_li, n1656_li, n1659_li, n1662_li,
    n1665_li, n1668_li, n1671_li, n1674_li, n1677_li, n1680_li, n1683_li,
    n1686_li, n1689_li, n1692_li, n1695_li, n1698_li, n1701_li, n1704_li,
    n1707_li, n1710_li, n1713_li, n1716_li, n1719_li, n1722_li, n1725_li,
    n1728_li, n1731_li, n1734_li, n1737_li, n1740_li, n1743_li, n1746_li,
    n1749_li, n1752_li, n1755_li, n1758_li, n1761_li, n1764_li, n1767_li,
    n1770_li, n1773_li, n1776_li, n1779_li, n1782_li, n1785_li, n1788_li,
    n1791_li, n1794_li, n1797_li, n1800_li, n1803_li, n1806_li, n1809_li,
    n1812_li, n1815_li, n1818_li, n1821_li, n1824_li, n1827_li, n1830_li,
    n1833_li, n1836_li, n1839_li, n1842_li, n1845_li, n1848_li, n1851_li,
    n1854_li, n1857_li, n1860_li, n1863_li, n1866_li, n1869_li, n1872_li,
    n1875_li, n1878_li, n1881_li, n1884_li, n1887_li, n1890_li, n1893_li,
    n1896_li, n1899_li, n1902_li, n1905_li, n1908_li, n1911_li, n1914_li,
    n1917_li, n1920_li, n1923_li, n1926_li, n1929_li, n1932_li, n1935_li,
    n1938_li, n1941_li, n1944_li, n1947_li, n1950_li, n1953_li, n1956_li,
    n1959_li, n1962_li, n1965_li, n1968_li, n1971_li, n1974_li, n1977_li,
    n1980_li, n1983_li, n1986_li, n1989_li, n1992_li, n1995_li, n1998_li,
    n2001_li, n2004_li, n2007_li, n2010_li, n2013_li, n2016_li, n2019_li,
    n2022_li, n2025_li, n2028_li, n2031_li, n2034_li, n2037_li, n2040_li,
    n2043_li, n2046_li, n2049_li, n2052_li, n2055_li, n2058_li, n2061_li,
    n2064_li, n2067_li, n2070_li, n2073_li, n2076_li, n2079_li, n2082_li,
    n2085_li, n2088_li, n2091_li, n2094_li, n2097_li, n2100_li, n2103_li,
    n2106_li, n2109_li, n2112_li, n2115_li, n2118_li, n2121_li, n2124_li,
    n2127_li, n2130_li, n2133_li, n2136_li, n2139_li, n2142_li, n2145_li,
    n2148_li, n2151_li, n2154_li, n2157_li, n2160_li, n2163_li, n2166_li,
    n2169_li, n2172_li, n2175_li, n2178_li, n2181_li, n2184_li, n2187_li,
    n2190_li, n2193_li, n2196_li, n2199_li, n2202_li, n2205_li, n2208_li,
    n2211_li, n2214_li, n2217_li, n2220_li, n2223_li, n2226_li, n2229_li,
    n2232_li, n2235_li, n2238_li, n2241_li, n2244_li, n2247_li, n2250_li,
    n2253_li, n2256_li, n2259_li, n2262_li, n2265_li, n2268_li, n2271_li,
    n2274_li, n2277_li, n2280_li, n2283_li, n2286_li, n2289_li, n2292_li,
    n2295_li, n2298_li, n2301_li, n2304_li, n2307_li, n2310_li, n2313_li,
    n2316_li, n2319_li, n2322_li, n2325_li, n2328_li, n2331_li, n2334_li,
    n2337_li, n2340_li, n2343_li, n2346_li, n2349_li, n2352_li, n2355_li,
    n2358_li, n2361_li, n2364_li, n2367_li, n2370_li, n2373_li, n2376_li,
    n2379_li, n2382_li, n2385_li, n2388_li, n2391_li, n2394_li, n2397_li,
    n2400_li, n2403_li, n2406_li, n2409_li, n2412_li, n2415_li, n2418_li,
    n2421_li, n2424_li, n2427_li, n2430_li, n2433_li, n2436_li, n2439_li,
    n2442_li, n2445_li, n2448_li, n2451_li, n2454_li, n2457_li, n2460_li,
    n2463_li, n2466_li, n2469_li, n2472_li, n2475_li, n2478_li, n2481_li,
    n2484_li, n2487_li, n2490_li, n2493_li, n2496_li, n2499_li, n2502_li,
    n2505_li, n2508_li, n2511_li, n2514_li, n2517_li, n2520_li, n2523_li,
    n2526_li, n2529_li, n2532_li, n2535_li, n2538_li, n2541_li, n2544_li,
    n2547_li, n2550_li, n2553_li, n2556_li, n2559_li, n2562_li, n2565_li,
    n2568_li, n2571_li, n2574_li, n2577_li, n2580_li, n2583_li, n2586_li,
    n2589_li, n2592_li, n2595_li, n2598_li, n2601_li, n2604_li, n2607_li,
    n2610_li, n2613_li, n2616_li, n2619_li, n2622_li, n2625_li, n2628_li,
    n2631_li, n2634_li, n2637_li, n2640_li, n2643_li, n2646_li, n2649_li,
    n2652_li, n2655_li, n2658_li, n2661_li, n2664_li, n2667_li, n2670_li,
    n2673_li, n2676_li, n2679_li, n2682_li, n2685_li, n2688_li, n2691_li,
    n2694_li, n2697_li, n2700_li, n2703_li, n2706_li, n2709_li, n2712_li,
    n2715_li, n2718_li, n2721_li, n2724_li, n2727_li, n2730_li, n2733_li,
    n2736_li, n2739_li, n2742_li, n2745_li, n2748_li, n2751_li, n2754_li,
    n2757_li, n2760_li, n2763_li, n2766_li, n2769_li, n2772_li, n2775_li,
    n2778_li, n2781_li, n2784_li, n2787_li, n2790_li, n2793_li, n2796_li,
    n2799_li, n2802_li, n2805_li, n2808_li, n2811_li, n2814_li, n2817_li,
    n2820_li, n2823_li, n2826_li, n2829_li, n2832_li, n2835_li, n2838_li,
    n2841_li, n2844_li, n2847_li, n2850_li, n2853_li, n2856_li, n2859_li,
    n2862_li, n2865_li, n2868_li, n2871_li, n2874_li, n2877_li, n2880_li,
    n2883_li, n2886_li, n2889_li, n2892_li, n2895_li, n2898_li, n2901_li,
    n2904_li, n2907_li, n2910_li, n2913_li, n2916_li, n2919_li, n2922_li,
    n2925_li, n2928_li, n2931_li, n2934_li, n2937_li, n2940_li, n2943_li,
    n2946_li, n2949_li, n2952_li, n2955_li, n2958_li, n2961_li, n2964_li,
    n2967_li, n2970_li, n2973_li, n2976_li, n2979_li, n2982_li, n2985_li,
    n2988_li, n2991_li, n2994_li, n2997_li, n3000_li, n3003_li, n3006_li,
    n3009_li, n3012_li, n3015_li, n3018_li, n3021_li, n3024_li, n3027_li,
    n3030_li, n3033_li, n3036_li, n3039_li, n3042_li, n3045_li, n3048_li,
    n3051_li, n3054_li, n3057_li, n3060_li, n3063_li, n3066_li, n3069_li,
    n3072_li, n3075_li, n3078_li, n3081_li, n3084_li, n3087_li, n3090_li,
    n3093_li, n3096_li, n3099_li, n3102_li, n3105_li, n3108_li, n3111_li,
    n3114_li, n3117_li, n3120_li, n3123_li, n3126_li, n3129_li, n3132_li,
    n3135_li, n3138_li, n3141_li, n3144_li, n3147_li, n3150_li, n3153_li,
    n3156_li, n3159_li, n3162_li, n3165_li, n3168_li, n3171_li, n3174_li,
    n3177_li, n3180_li, n3183_li, n3186_li, n3189_li, n3192_li, n3195_li,
    n3198_li, n3201_li, n3204_li, n3207_li, n3210_li, n3213_li, n3216_li,
    n3219_li, n3222_li, n3225_li, n3228_li, n3231_li, n3234_li, n3237_li,
    n3240_li, n3243_li, n3246_li, n3249_li, n3252_li, n3255_li, n3258_li,
    n3261_li, n3264_li, n3267_li, n3270_li, n3273_li, n3276_li, n3279_li,
    n3282_li, n3285_li, n3288_li, n3291_li, n3294_li, n3297_li;
  assign new_G282_ = n1425_lo & n1449_lo;
  assign new_G283_ = ~n2829_lo;
  assign new_G284_ = ~n2937_lo;
  assign new_G285_ = n3081_lo & n3117_lo & n3105_lo & n3093_lo;
  assign new_G286_ = ~new_G282_;
  assign new_G287_ = n1437_lo & n1545_lo & n2865_lo;
  assign new_G288_ = ~n2865_lo;
  assign new_G291_ = n1761_lo & n1761_lo;
  assign new_G292_ = ~n2793_lo;
  assign new_G295_ = ~n1509_lo;
  assign new_G298_ = ~n1509_lo;
  assign new_G301_ = ~n2817_lo;
  assign new_G313_ = ~n2853_lo;
  assign new_G325_ = ~n2877_lo;
  assign new_G329_ = ~n2889_lo;
  assign new_G335_ = n1521_lo & n2889_lo;
  assign new_G336_ = n1797_lo & n2685_lo & n2181_lo & n2325_lo;
  assign new_G339_ = n2049_lo & n2565_lo & n1929_lo & n2445_lo;
  assign new_G342_ = ~n2817_lo;
  assign new_G354_ = ~n2853_lo;
  assign new_G366_ = ~n2913_lo;
  assign new_G370_ = ~n2925_lo;
  assign new_G374_ = ~n3153_lo;
  assign new_G386_ = ~n3165_lo;
  assign new_G398_ = ~n3189_lo;
  assign new_G399_ = ~n3201_lo;
  assign new_G400_ = ~n3213_lo;
  assign new_G401_ = ~n3225_lo;
  assign new_G402_ = ~n3237_lo;
  assign new_G403_ = ~n3249_lo;
  assign new_G404_ = ~n3285_lo;
  assign new_G405_ = ~n3153_lo;
  assign new_G417_ = ~n3165_lo;
  assign new_G429_ = ~n1557_lo;
  assign new_G435_ = ~n1557_lo;
  assign new_G442_ = ~n3297_lo;
  assign new_G443_ = n1497_lo & n2865_lo;
  assign new_G447_ = ~n2949_lo;
  assign new_G451_ = ~n2961_lo;
  assign new_G455_ = ~n2973_lo;
  assign new_G459_ = ~n2985_lo;
  assign new_G463_ = ~n2997_lo;
  assign new_G467_ = ~n3009_lo;
  assign new_G471_ = ~n3021_lo;
  assign new_G475_ = ~n3033_lo;
  assign new_G479_ = ~n3045_lo;
  assign new_G485_ = ~n1689_lo;
  assign new_G491_ = ~n1689_lo;
  assign new_G497_ = ~n3069_lo;
  assign new_G503_ = ~n3081_lo;
  assign new_G507_ = ~n3093_lo;
  assign new_G511_ = ~n3105_lo;
  assign new_G515_ = ~n3117_lo;
  assign new_G519_ = ~n3129_lo;
  assign new_G522_ = ~n3141_lo;
  assign new_G525_ = ~n3261_lo;
  assign new_G526_ = ~n3273_lo;
  assign new_G527_ = ~n2925_lo;
  assign new_G530_ = ~n2913_lo;
  assign new_G533_ = ~n2949_lo;
  assign new_G536_ = ~n2973_lo;
  assign new_G539_ = ~n2961_lo;
  assign new_G542_ = ~n2997_lo;
  assign new_G545_ = ~n2985_lo;
  assign new_G548_ = ~n3021_lo;
  assign new_G551_ = ~n3009_lo;
  assign new_G554_ = ~n3045_lo;
  assign new_G557_ = ~n3033_lo;
  assign new_G560_ = ~n3069_lo;
  assign new_G563_ = ~n3093_lo;
  assign new_G566_ = ~n3081_lo;
  assign new_G569_ = ~n3117_lo;
  assign new_G572_ = ~n3105_lo;
  assign new_G575_ = ~n3141_lo;
  assign new_G578_ = ~n3129_lo;
  assign new_G581_ = ~new_G291_;
  assign new_G584_ = ~n3201_lo | ~new_G398_;
  assign new_G585_ = ~n3189_lo | ~new_G399_;
  assign new_G586_ = ~n3225_lo | ~new_G400_;
  assign new_G587_ = ~n3213_lo | ~new_G401_;
  assign new_G588_ = ~n3249_lo | ~new_G402_;
  assign new_G589_ = ~n3237_lo | ~new_G403_;
  assign new_G590_ = ~n3273_lo | ~new_G525_;
  assign new_G591_ = ~n3261_lo | ~new_G526_;
  assign new_G592_ = n3177_lo & new_G443_;
  assign new_G593_ = ~new_G336_;
  assign new_G594_ = ~new_G339_;
  assign new_G595_ = new_G339_ & new_G336_;
  assign new_G598_ = ~new_G295_;
  assign new_G603_ = ~new_G301_;
  assign new_G614_ = ~new_G313_;
  assign new_G625_ = n2157_lo & new_G301_ & new_G313_;
  assign new_G626_ = n2037_lo & new_G301_ & new_G313_;
  assign new_G627_ = n2145_lo & new_G301_ & new_G313_;
  assign new_G628_ = n2133_lo & new_G301_ & new_G313_;
  assign new_G629_ = n2121_lo & new_G301_ & new_G313_;
  assign new_G630_ = n1521_lo & new_G329_;
  assign new_G631_ = ~new_G295_;
  assign new_G636_ = ~new_G342_;
  assign new_G647_ = ~new_G354_;
  assign new_G658_ = n2109_lo & new_G342_ & new_G354_;
  assign new_G659_ = n2097_lo & new_G342_ & new_G354_;
  assign new_G660_ = n2085_lo & new_G342_ & new_G354_;
  assign new_G661_ = n2073_lo & new_G342_ & new_G354_;
  assign new_G662_ = n2061_lo & new_G342_ & new_G354_;
  assign new_G663_ = ~new_G374_;
  assign new_G674_ = ~new_G386_;
  assign new_G685_ = n2493_lo & new_G374_ & new_G386_;
  assign new_G686_ = n2481_lo & new_G374_ & new_G386_;
  assign new_G687_ = n2469_lo & new_G374_ & new_G386_;
  assign new_G688_ = n2457_lo & new_G374_ & new_G386_;
  assign new_G689_ = new_G374_ & new_G386_;
  assign new_G690_ = ~new_G584_ | ~new_G585_;
  assign new_G694_ = ~new_G586_ | ~new_G587_;
  assign new_G698_ = ~new_G588_ | ~new_G589_;
  assign new_G701_ = ~new_G533_;
  assign new_G702_ = ~new_G533_ | ~new_G404_;
  assign new_G703_ = ~new_G536_;
  assign new_G704_ = ~new_G539_;
  assign new_G705_ = ~new_G542_;
  assign new_G706_ = ~new_G545_;
  assign new_G707_ = ~new_G405_;
  assign new_G718_ = ~new_G417_;
  assign new_G729_ = n2541_lo & new_G405_ & new_G417_;
  assign new_G730_ = n2433_lo & new_G405_ & new_G417_;
  assign new_G731_ = n2529_lo & new_G405_ & new_G417_;
  assign new_G732_ = n2517_lo & new_G405_ & new_G417_;
  assign new_G733_ = n2505_lo & new_G405_ & new_G417_;
  assign new_G734_ = ~new_G429_;
  assign new_G739_ = ~new_G435_;
  assign new_G745_ = ~new_G560_;
  assign new_G746_ = ~new_G560_ | ~new_G442_;
  assign new_G747_ = ~new_G563_;
  assign new_G748_ = ~new_G566_;
  assign new_G749_ = ~new_G569_;
  assign new_G750_ = ~new_G572_;
  assign new_G751_ = ~new_G298_;
  assign new_G756_ = ~new_G298_;
  assign new_G761_ = ~new_G485_;
  assign new_G766_ = ~new_G491_;
  assign new_G771_ = ~new_G527_;
  assign new_G772_ = ~new_G530_;
  assign new_G773_ = ~new_G548_;
  assign new_G774_ = ~new_G551_;
  assign new_G775_ = ~new_G554_;
  assign new_G776_ = ~new_G557_;
  assign new_G777_ = ~new_G590_ | ~new_G591_;
  assign new_G780_ = ~new_G366_;
  assign new_G783_ = ~new_G370_;
  assign new_G786_ = ~new_G447_;
  assign new_G789_ = ~new_G451_;
  assign new_G792_ = ~new_G455_;
  assign new_G795_ = ~new_G459_;
  assign new_G798_ = ~new_G463_;
  assign new_G801_ = ~new_G467_;
  assign new_G804_ = ~new_G471_;
  assign new_G807_ = ~new_G475_;
  assign new_G810_ = ~new_G575_;
  assign new_G811_ = ~new_G578_;
  assign new_G812_ = ~new_G479_;
  assign new_G815_ = ~new_G497_;
  assign new_G818_ = ~new_G503_;
  assign new_G821_ = ~new_G507_;
  assign new_G824_ = ~new_G511_;
  assign new_G827_ = ~new_G515_;
  assign new_G830_ = n3177_lo & new_G593_;
  assign new_G831_ = n2841_lo & new_G594_;
  assign new_G832_ = new_G630_ | new_G335_;
  assign new_G833_ = ~n3285_lo | ~new_G701_;
  assign new_G834_ = ~new_G539_ | ~new_G703_;
  assign new_G835_ = ~new_G536_ | ~new_G704_;
  assign new_G836_ = ~new_G545_ | ~new_G705_;
  assign new_G837_ = ~new_G542_ | ~new_G706_;
  assign new_G838_ = ~n3297_lo | ~new_G745_;
  assign new_G839_ = ~new_G566_ | ~new_G747_;
  assign new_G840_ = ~new_G563_ | ~new_G748_;
  assign new_G841_ = ~new_G572_ | ~new_G749_;
  assign new_G842_ = ~new_G569_ | ~new_G750_;
  assign new_G843_ = ~new_G530_ | ~new_G771_;
  assign new_G844_ = ~new_G527_ | ~new_G772_;
  assign new_G845_ = ~new_G551_ | ~new_G773_;
  assign new_G846_ = ~new_G548_ | ~new_G774_;
  assign new_G847_ = ~new_G557_ | ~new_G775_;
  assign new_G848_ = ~new_G554_ | ~new_G776_;
  assign new_G849_ = ~new_G578_ | ~new_G810_;
  assign new_G850_ = ~new_G575_ | ~new_G811_;
  assign new_G851_ = ~new_G830_;
  assign new_G852_ = ~new_G831_;
  assign new_G853_ = n2289_lo & new_G603_ & new_G614_;
  assign new_G854_ = n1905_lo & new_G301_ & new_G614_;
  assign new_G855_ = n2025_lo & new_G603_ & new_G313_;
  assign new_G856_ = n2169_lo & new_G603_ & new_G614_;
  assign new_G857_ = n1785_lo & new_G301_ & new_G614_;
  assign new_G858_ = n1917_lo & new_G603_ & new_G313_;
  assign new_G859_ = n2277_lo & new_G603_ & new_G614_;
  assign new_G860_ = n1893_lo & new_G301_ & new_G614_;
  assign new_G861_ = n2013_lo & new_G603_ & new_G313_;
  assign new_G862_ = n2265_lo & new_G603_ & new_G614_;
  assign new_G863_ = n1881_lo & new_G301_ & new_G614_;
  assign new_G864_ = n2001_lo & new_G603_ & new_G313_;
  assign new_G865_ = n2253_lo & new_G603_ & new_G614_;
  assign new_G866_ = n1869_lo & new_G301_ & new_G614_;
  assign new_G867_ = n1989_lo & new_G603_ & new_G313_;
  assign new_G868_ = n2241_lo & new_G636_ & new_G647_;
  assign new_G869_ = n1857_lo & new_G342_ & new_G647_;
  assign new_G870_ = n1977_lo & new_G636_ & new_G354_;
  assign new_G871_ = n2229_lo & new_G636_ & new_G647_;
  assign new_G872_ = n1845_lo & new_G342_ & new_G647_;
  assign new_G873_ = n1965_lo & new_G636_ & new_G354_;
  assign new_G874_ = n2217_lo & new_G636_ & new_G647_;
  assign new_G875_ = n1833_lo & new_G342_ & new_G647_;
  assign new_G876_ = new_G636_ & new_G354_;
  assign new_G877_ = n2205_lo & new_G636_ & new_G647_;
  assign new_G878_ = n1821_lo & new_G342_ & new_G647_;
  assign new_G879_ = n1953_lo & new_G636_ & new_G354_;
  assign new_G880_ = n2193_lo & new_G636_ & new_G647_;
  assign new_G881_ = n1809_lo & new_G342_ & new_G647_;
  assign new_G882_ = n1941_lo & new_G636_ & new_G354_;
  assign new_G883_ = n2733_lo & new_G663_ & new_G674_;
  assign new_G884_ = n2373_lo & new_G374_ & new_G674_;
  assign new_G885_ = n2613_lo & new_G663_ & new_G386_;
  assign new_G886_ = n2721_lo & new_G663_ & new_G674_;
  assign new_G887_ = n2361_lo & new_G374_ & new_G674_;
  assign new_G888_ = n2601_lo & new_G663_ & new_G386_;
  assign new_G889_ = n2709_lo & new_G663_ & new_G674_;
  assign new_G890_ = n2349_lo & new_G374_ & new_G674_;
  assign new_G891_ = n2589_lo & new_G663_ & new_G386_;
  assign new_G892_ = n2697_lo & new_G663_ & new_G674_;
  assign new_G893_ = n2337_lo & new_G374_ & new_G674_;
  assign new_G894_ = n2577_lo & new_G663_ & new_G386_;
  assign new_G895_ = new_G663_ & new_G674_;
  assign new_G896_ = new_G374_ & new_G674_;
  assign new_G897_ = new_G663_ & new_G386_;
  assign new_G898_ = ~new_G690_;
  assign new_G901_ = ~new_G694_;
  assign new_G904_ = ~new_G833_ | ~new_G702_;
  assign new_G908_ = ~new_G834_ | ~new_G835_;
  assign new_G912_ = ~new_G836_ | ~new_G837_;
  assign new_G915_ = ~new_G698_;
  assign new_G918_ = ~new_G698_;
  assign new_G921_ = ~new_G780_;
  assign new_G922_ = ~new_G783_;
  assign new_G923_ = ~new_G786_;
  assign new_G924_ = ~new_G789_;
  assign new_G925_ = ~new_G792_;
  assign new_G926_ = ~new_G795_;
  assign new_G927_ = ~new_G798_;
  assign new_G928_ = ~new_G801_;
  assign new_G929_ = ~new_G804_;
  assign new_G930_ = ~new_G807_;
  assign new_G931_ = n2781_lo & new_G707_ & new_G718_;
  assign new_G932_ = n2421_lo & new_G405_ & new_G718_;
  assign new_G933_ = n2661_lo & new_G707_ & new_G417_;
  assign new_G934_ = n2673_lo & new_G707_ & new_G718_;
  assign new_G935_ = n2313_lo & new_G405_ & new_G718_;
  assign new_G936_ = n2553_lo & new_G707_ & new_G417_;
  assign new_G937_ = n2769_lo & new_G707_ & new_G718_;
  assign new_G938_ = n2409_lo & new_G405_ & new_G718_;
  assign new_G939_ = n2649_lo & new_G707_ & new_G417_;
  assign new_G940_ = n2757_lo & new_G707_ & new_G718_;
  assign new_G941_ = n2397_lo & new_G405_ & new_G718_;
  assign new_G942_ = n2637_lo & new_G707_ & new_G417_;
  assign new_G943_ = n2745_lo & new_G707_ & new_G718_;
  assign new_G944_ = n2385_lo & new_G405_ & new_G718_;
  assign new_G945_ = n2625_lo & new_G707_ & new_G417_;
  assign new_G946_ = n1569_lo & new_G734_;
  assign new_G947_ = n1461_lo & new_G734_;
  assign new_G948_ = n1581_lo & new_G734_;
  assign new_G949_ = n1473_lo & new_G734_;
  assign new_G950_ = n1593_lo & new_G739_;
  assign new_G951_ = n1605_lo & new_G739_;
  assign new_G952_ = n1617_lo & new_G739_;
  assign new_G953_ = n1485_lo & new_G739_;
  assign new_G954_ = n1629_lo & new_G739_;
  assign new_G955_ = ~new_G838_ | ~new_G746_;
  assign new_G959_ = ~new_G839_ | ~new_G840_;
  assign new_G963_ = ~new_G841_ | ~new_G842_;
  assign new_G966_ = n1641_lo & new_G761_;
  assign new_G967_ = n1701_lo & new_G761_;
  assign new_G968_ = n1653_lo & new_G761_;
  assign new_G969_ = n1713_lo & new_G761_;
  assign new_G970_ = n1665_lo & new_G766_;
  assign new_G971_ = n1725_lo & new_G766_;
  assign new_G972_ = n1737_lo & new_G766_;
  assign new_G973_ = n1677_lo & new_G766_;
  assign new_G974_ = ~new_G812_;
  assign new_G975_ = ~new_G815_;
  assign new_G976_ = ~new_G818_;
  assign new_G977_ = ~new_G821_;
  assign new_G978_ = ~new_G824_;
  assign new_G979_ = ~new_G827_;
  assign new_G980_ = ~new_G843_ | ~new_G844_;
  assign new_G983_ = ~new_G777_;
  assign new_G984_ = ~new_G847_ | ~new_G848_;
  assign new_G987_ = ~new_G845_ | ~new_G846_;
  assign new_G990_ = ~new_G849_ | ~new_G850_;
  assign new_G993_ = new_G851_ & new_G852_;
  assign new_G998_ = new_G625_ | new_G855_ | new_G853_ | new_G854_;
  assign new_G1002_ = new_G626_ | new_G858_ | new_G856_ | new_G857_;
  assign new_G1008_ = new_G627_ | new_G861_ | new_G859_ | new_G860_;
  assign new_G1014_ = new_G628_ | new_G864_ | new_G862_ | new_G863_;
  assign new_G1017_ = new_G629_ | new_G867_ | new_G865_ | new_G866_;
  assign new_G1021_ = new_G658_ | new_G870_ | new_G868_ | new_G869_;
  assign new_G1026_ = new_G659_ | new_G873_ | new_G871_ | new_G872_;
  assign new_G1030_ = new_G660_ | new_G876_ | new_G874_ | new_G875_;
  assign new_G1033_ = new_G661_ | new_G879_ | new_G877_ | new_G878_;
  assign new_G1036_ = new_G662_ | new_G882_ | new_G880_ | new_G881_;
  assign new_G1039_ = new_G685_ | new_G885_ | new_G883_ | new_G884_;
  assign new_G1044_ = new_G686_ | new_G888_ | new_G886_ | new_G887_;
  assign new_G1049_ = new_G687_ | new_G891_ | new_G889_ | new_G890_;
  assign new_G1053_ = new_G688_ | new_G894_ | new_G892_ | new_G893_;
  assign new_G1058_ = new_G689_ | new_G897_ | new_G895_ | new_G896_;
  assign new_G1062_ = new_G730_ | new_G936_ | new_G934_ | new_G935_;
  assign new_G1067_ = new_G731_ | new_G939_ | new_G937_ | new_G938_;
  assign new_G1072_ = new_G732_ | new_G942_ | new_G940_ | new_G941_;
  assign new_G1076_ = new_G733_ | new_G945_ | new_G943_ | new_G944_;
  assign new_G1079_ = new_G729_ | new_G933_ | new_G931_ | new_G932_;
  assign new_G1082_ = ~new_G904_;
  assign new_G1085_ = ~new_G908_;
  assign new_G1088_ = ~new_G915_;
  assign new_G1089_ = ~new_G918_;
  assign new_G1090_ = ~new_G912_;
  assign new_G1093_ = ~new_G912_;
  assign new_G1096_ = new_G694_ & new_G690_ & new_G915_;
  assign new_G1097_ = new_G901_ & new_G898_ & new_G918_;
  assign new_G1098_ = ~new_G955_;
  assign new_G1101_ = ~new_G959_;
  assign new_G1104_ = ~new_G963_;
  assign new_G1107_ = ~new_G963_;
  assign new_G1110_ = ~new_G990_;
  assign new_G1111_ = ~new_G980_;
  assign new_G1112_ = ~new_G980_ | ~new_G983_;
  assign new_G1113_ = ~new_G984_;
  assign new_G1114_ = ~new_G987_;
  assign new_G1115_ = new_G998_ & n2877_lo;
  assign new_G1116_ = new_G1008_ & n2877_lo;
  assign new_G1117_ = new_G1002_ & n2877_lo;
  assign new_G1118_ = new_G993_ & new_G288_ & n2805_lo & n1749_lo;
  assign new_G1119_ = new_G286_ & new_G288_ & n2805_lo & new_G993_;
  assign new_G1120_ = ~new_G998_;
  assign new_G1123_ = ~new_G1008_;
  assign new_G1126_ = new_G1002_ & new_G329_;
  assign new_G1127_ = new_G1008_ & new_G329_;
  assign new_G1128_ = new_G1021_ & n2889_lo;
  assign new_G1129_ = ~new_G998_;
  assign new_G1132_ = ~new_G1002_;
  assign new_G1137_ = ~new_G1008_;
  assign new_G1144_ = ~new_G1014_;
  assign new_G1148_ = ~new_G1017_;
  assign new_G1152_ = ~new_G1021_;
  assign new_G1159_ = ~new_G1026_;
  assign new_G1166_ = ~new_G1030_;
  assign new_G1171_ = ~new_G1033_;
  assign new_G1176_ = ~new_G1036_;
  assign new_G1181_ = ~new_G519_ | ~new_G1053_;
  assign new_G1184_ = ~new_G522_ | ~new_G1058_;
  assign new_G1187_ = ~new_G1072_;
  assign new_G1190_ = new_G1039_ & new_G284_;
  assign new_G1193_ = ~new_G1044_;
  assign new_G1196_ = new_G898_ & new_G694_ & new_G1088_;
  assign new_G1197_ = new_G690_ & new_G901_ & new_G1089_;
  assign new_G1198_ = new_G1002_ & new_G429_;
  assign new_G1199_ = new_G1008_ & new_G429_;
  assign new_G1200_ = new_G1014_ & new_G429_;
  assign new_G1201_ = new_G1017_ & new_G429_;
  assign new_G1202_ = new_G1021_ & new_G435_;
  assign new_G1203_ = new_G1026_ & new_G435_;
  assign new_G1204_ = new_G1030_ & new_G435_;
  assign new_G1205_ = new_G1033_ & new_G435_;
  assign new_G1206_ = new_G1036_ & new_G435_;
  assign new_G1207_ = ~new_G1079_;
  assign new_G1208_ = new_G1062_ & new_G485_;
  assign new_G1209_ = new_G1067_ & new_G485_;
  assign new_G1210_ = new_G1072_ & new_G485_;
  assign new_G1211_ = new_G1076_ & new_G485_;
  assign new_G1212_ = new_G1039_ & new_G491_;
  assign new_G1213_ = new_G1044_ & new_G491_;
  assign new_G1214_ = new_G1049_ & new_G491_;
  assign new_G1215_ = new_G1053_ & new_G491_;
  assign new_G1216_ = ~new_G1002_;
  assign new_G1219_ = ~new_G777_ | ~new_G1111_;
  assign new_G1220_ = ~new_G987_ | ~new_G1113_;
  assign new_G1221_ = ~new_G984_ | ~new_G1114_;
  assign new_G1222_ = ~new_G1062_;
  assign new_G1225_ = ~new_G1072_;
  assign new_G1228_ = ~new_G1067_;
  assign new_G1231_ = ~new_G1039_;
  assign new_G1234_ = ~new_G1076_;
  assign new_G1237_ = ~new_G1049_;
  assign new_G1240_ = ~new_G1044_;
  assign new_G1243_ = ~new_G1058_;
  assign new_G1246_ = ~new_G1053_;
  assign new_G1249_ = ~new_G1090_;
  assign new_G1250_ = ~new_G1093_;
  assign new_G1251_ = ~new_G1196_ & ~new_G1096_;
  assign new_G1252_ = ~new_G1197_ & ~new_G1097_;
  assign new_G1253_ = new_G908_ & new_G904_ & new_G1090_;
  assign new_G1254_ = new_G1085_ & new_G1082_ & new_G1093_;
  assign new_G1255_ = new_G973_ | new_G1215_;
  assign new_G1256_ = ~new_G1104_;
  assign new_G1257_ = ~new_G1107_;
  assign new_G1258_ = new_G959_ & new_G955_ & new_G1104_;
  assign new_G1259_ = new_G1101_ & new_G1098_ & new_G1107_;
  assign new_G1260_ = ~new_G1219_ | ~new_G1112_;
  assign new_G1263_ = ~new_G1220_ | ~new_G1221_;
  assign new_G1266_ = new_G946_ | new_G1198_;
  assign new_G1269_ = new_G947_ | new_G1199_;
  assign new_G1272_ = new_G948_ | new_G1200_;
  assign new_G1275_ = new_G949_ | new_G1201_;
  assign new_G1278_ = new_G950_ | new_G1202_;
  assign new_G1281_ = new_G951_ | new_G1203_;
  assign new_G1284_ = new_G952_ | new_G1204_;
  assign new_G1287_ = new_G953_ | new_G1205_;
  assign new_G1290_ = new_G954_ | new_G1206_;
  assign new_G1293_ = new_G966_ | new_G1208_;
  assign new_G1296_ = new_G967_ | new_G1209_;
  assign new_G1299_ = new_G968_ | new_G1210_;
  assign new_G1302_ = new_G969_ | new_G1211_;
  assign new_G1305_ = new_G970_ | new_G1212_;
  assign new_G1308_ = new_G971_ | new_G1213_;
  assign new_G1311_ = new_G972_ | new_G1214_;
  assign new_G1314_ = new_G1193_ & new_G1190_ & n1773_lo;
  assign new_G1320_ = ~new_G1190_;
  assign new_G1321_ = ~new_G283_ | ~new_G1123_;
  assign new_G1326_ = new_G1120_ & new_G329_;
  assign new_G1327_ = new_G1148_ & n2889_lo;
  assign new_G1328_ = new_G1144_ & new_G329_;
  assign new_G1329_ = ~new_G1144_;
  assign new_G1336_ = ~new_G1148_;
  assign new_G1342_ = ~new_G1159_;
  assign new_G1345_ = ~new_G1166_;
  assign new_G1348_ = ~new_G1171_;
  assign new_G1351_ = ~new_G1176_;
  assign new_G1354_ = new_G519_ & new_G1181_;
  assign new_G1355_ = new_G1181_ & new_G1053_;
  assign new_G1356_ = new_G522_ & new_G1184_;
  assign new_G1357_ = new_G1184_ & new_G1058_;
  assign new_G1358_ = new_G1082_ & new_G908_ & new_G1249_;
  assign new_G1359_ = new_G904_ & new_G1085_ & new_G1250_;
  assign new_G1360_ = ~new_G1222_;
  assign new_G1361_ = ~new_G1222_ | ~new_G1207_;
  assign new_G1362_ = ~new_G1225_;
  assign new_G1363_ = ~new_G1228_;
  assign new_G1364_ = ~new_G1231_;
  assign new_G1365_ = ~new_G1234_;
  assign new_G1366_ = new_G1098_ & new_G959_ & new_G1256_;
  assign new_G1367_ = new_G955_ & new_G1101_ & new_G1257_;
  assign new_G1368_ = ~new_G1132_;
  assign new_G1371_ = ~new_G1129_;
  assign new_G1374_ = ~new_G1137_;
  assign new_G1377_ = ~new_G1152_;
  assign new_G1380_ = ~new_G1123_;
  assign new_G1383_ = ~new_G1216_;
  assign new_G1384_ = ~new_G1132_;
  assign new_G1387_ = ~new_G1129_;
  assign new_G1390_ = ~new_G1137_;
  assign new_G1393_ = ~new_G1120_;
  assign new_G1396_ = ~new_G1137_;
  assign new_G1399_ = ~new_G1137_;
  assign new_G1402_ = ~new_G1252_ | ~new_G1251_;
  assign new_G1405_ = ~new_G1237_;
  assign new_G1406_ = ~new_G1240_;
  assign new_G1407_ = ~new_G1243_;
  assign new_G1408_ = ~new_G1246_;
  assign new_G1409_ = n1773_lo & new_G1193_ & new_G1320_;
  assign new_G1412_ = new_G1127_ | new_G1327_;
  assign new_G1415_ = new_G1328_ | new_G1128_;
  assign new_G1418_ = new_G1354_ | new_G1355_;
  assign new_G1421_ = new_G1356_ | new_G1357_;
  assign new_G1424_ = ~new_G1358_ & ~new_G1253_;
  assign new_G1425_ = ~new_G1359_ & ~new_G1254_;
  assign new_G1426_ = ~new_G1260_;
  assign new_G1427_ = ~new_G1263_;
  assign new_G1428_ = ~new_G1266_ | ~new_G921_;
  assign new_G1429_ = ~new_G1266_;
  assign new_G1430_ = ~new_G1269_ | ~new_G922_;
  assign new_G1431_ = ~new_G1269_;
  assign new_G1432_ = ~new_G1272_ | ~new_G923_;
  assign new_G1433_ = ~new_G1272_;
  assign new_G1434_ = ~new_G1275_ | ~new_G924_;
  assign new_G1435_ = ~new_G1275_;
  assign new_G1436_ = ~new_G1278_ | ~new_G925_;
  assign new_G1437_ = ~new_G1278_;
  assign new_G1438_ = ~new_G1281_ | ~new_G926_;
  assign new_G1439_ = ~new_G1281_;
  assign new_G1440_ = ~new_G1284_ | ~new_G927_;
  assign new_G1441_ = ~new_G1284_;
  assign new_G1442_ = ~new_G1287_ | ~new_G928_;
  assign new_G1443_ = ~new_G1287_;
  assign new_G1444_ = ~new_G1290_ | ~new_G929_;
  assign new_G1445_ = ~new_G1290_;
  assign new_G1446_ = ~new_G1293_ | ~new_G930_;
  assign new_G1447_ = ~new_G1293_;
  assign new_G1448_ = ~new_G1079_ | ~new_G1360_;
  assign new_G1449_ = ~new_G1228_ | ~new_G1362_;
  assign new_G1450_ = ~new_G1225_ | ~new_G1363_;
  assign new_G1451_ = ~new_G1234_ | ~new_G1364_;
  assign new_G1452_ = ~new_G1231_ | ~new_G1365_;
  assign new_G1453_ = ~new_G1366_ & ~new_G1258_;
  assign new_G1454_ = ~new_G1367_ & ~new_G1259_;
  assign new_G1455_ = ~new_G1296_ | ~new_G974_;
  assign new_G1456_ = ~new_G1296_;
  assign new_G1457_ = ~new_G1299_ | ~new_G975_;
  assign new_G1458_ = ~new_G1299_;
  assign new_G1459_ = ~new_G1302_ | ~new_G976_;
  assign new_G1460_ = ~new_G1302_;
  assign new_G1461_ = ~new_G1305_ | ~new_G977_;
  assign new_G1462_ = ~new_G1305_;
  assign new_G1463_ = ~new_G1308_ | ~new_G978_;
  assign new_G1464_ = ~new_G1308_;
  assign new_G1465_ = ~new_G1311_ | ~new_G979_;
  assign new_G1466_ = ~new_G1311_;
  assign new_G1467_ = ~new_G1240_ | ~new_G1405_;
  assign new_G1468_ = ~new_G1237_ | ~new_G1406_;
  assign new_G1469_ = ~new_G1246_ | ~new_G1407_;
  assign new_G1470_ = ~new_G1243_ | ~new_G1408_;
  assign new_G1471_ = new_G1321_ & new_G325_;
  assign new_G1472_ = ~new_G1314_;
  assign new_G1475_ = ~new_G1368_;
  assign new_G1476_ = ~new_G1371_;
  assign new_G1477_ = ~new_G1374_;
  assign new_G1478_ = ~new_G1377_;
  assign new_G1479_ = ~new_G1321_;
  assign new_G1483_ = ~new_G1384_;
  assign new_G1484_ = ~new_G1387_;
  assign new_G1485_ = ~new_G1390_;
  assign new_G1486_ = ~new_G1393_;
  assign new_G1487_ = ~new_G1396_;
  assign new_G1488_ = ~new_G1314_;
  assign new_G1493_ = ~new_G1314_;
  assign new_G1497_ = new_G1321_ & n2889_lo;
  assign new_G1498_ = ~new_G1314_;
  assign new_G1502_ = ~new_G1314_;
  assign new_G1507_ = ~new_G1402_ | ~new_G1426_;
  assign new_G1508_ = ~new_G1399_;
  assign new_G1509_ = ~new_G1402_;
  assign new_G1510_ = ~new_G780_ | ~new_G1429_;
  assign new_G1511_ = ~new_G783_ | ~new_G1431_;
  assign new_G1512_ = ~new_G786_ | ~new_G1433_;
  assign new_G1513_ = ~new_G789_ | ~new_G1435_;
  assign new_G1514_ = ~new_G792_ | ~new_G1437_;
  assign new_G1515_ = ~new_G795_ | ~new_G1439_;
  assign new_G1516_ = ~new_G798_ | ~new_G1441_;
  assign new_G1517_ = ~new_G801_ | ~new_G1443_;
  assign new_G1518_ = ~new_G804_ | ~new_G1445_;
  assign new_G1519_ = ~new_G807_ | ~new_G1447_;
  assign new_G1520_ = ~new_G1448_ | ~new_G1361_;
  assign new_G1524_ = ~new_G1449_ | ~new_G1450_;
  assign new_G1528_ = ~new_G1451_ | ~new_G1452_;
  assign new_G1531_ = ~new_G812_ | ~new_G1456_;
  assign new_G1532_ = ~new_G815_ | ~new_G1458_;
  assign new_G1533_ = ~new_G818_ | ~new_G1460_;
  assign new_G1534_ = ~new_G821_ | ~new_G1462_;
  assign new_G1535_ = ~new_G824_ | ~new_G1464_;
  assign new_G1536_ = ~new_G827_ | ~new_G1466_;
  assign new_G1537_ = ~new_G1329_;
  assign new_G1540_ = ~new_G1336_;
  assign new_G1543_ = ~new_G1345_;
  assign new_G1546_ = ~new_G1342_;
  assign new_G1549_ = ~new_G1351_;
  assign new_G1552_ = ~new_G1348_;
  assign new_G1555_ = ~new_G1380_;
  assign new_G1556_ = ~new_G1380_ | ~new_G1383_;
  assign new_G1557_ = ~new_G1329_;
  assign new_G1560_ = ~new_G1345_;
  assign new_G1563_ = ~new_G1342_;
  assign new_G1566_ = ~new_G1351_;
  assign new_G1569_ = ~new_G1348_;
  assign new_G1572_ = ~new_G1321_;
  assign new_G1575_ = ~new_G1329_;
  assign new_G1578_ = ~new_G1336_;
  assign new_G1581_ = ~new_G1329_;
  assign new_G1584_ = ~new_G1336_;
  assign new_G1587_ = ~new_G1425_ | ~new_G1424_;
  assign new_G1590_ = ~new_G1469_ | ~new_G1470_;
  assign new_G1593_ = ~new_G1467_ | ~new_G1468_;
  assign new_G1596_ = ~new_G1454_ | ~new_G1453_;
  assign new_G1599_ = ~new_G1371_ | ~new_G1475_;
  assign new_G1600_ = ~new_G1368_ | ~new_G1476_;
  assign new_G1601_ = ~new_G1387_ | ~new_G1483_;
  assign new_G1602_ = ~new_G1384_ | ~new_G1484_;
  assign new_G1603_ = new_G1126_ | new_G1497_;
  assign new_G1606_ = ~new_G1260_ | ~new_G1509_;
  assign new_G1607_ = ~new_G1418_;
  assign new_G1610_ = ~new_G1421_;
  assign new_G1613_ = ~new_G1409_;
  assign new_G1616_ = ~new_G1409_;
  assign new_G1619_ = ~new_G1428_ | ~new_G1510_;
  assign new_G1620_ = ~new_G1430_ | ~new_G1511_;
  assign new_G1621_ = ~new_G1432_ | ~new_G1512_;
  assign new_G1622_ = ~new_G1434_ | ~new_G1513_;
  assign new_G1623_ = ~new_G1436_ | ~new_G1514_;
  assign new_G1624_ = ~new_G1438_ | ~new_G1515_;
  assign new_G1625_ = ~new_G1440_ | ~new_G1516_;
  assign new_G1626_ = ~new_G1442_ | ~new_G1517_;
  assign new_G1627_ = ~new_G1444_ | ~new_G1518_;
  assign new_G1628_ = ~new_G1446_ | ~new_G1519_;
  assign new_G1629_ = ~new_G1455_ | ~new_G1531_;
  assign new_G1630_ = ~new_G1457_ | ~new_G1532_;
  assign new_G1631_ = ~new_G1459_ | ~new_G1533_;
  assign new_G1632_ = ~new_G1461_ | ~new_G1534_;
  assign new_G1633_ = ~new_G1463_ | ~new_G1535_;
  assign new_G1634_ = ~new_G1465_ | ~new_G1536_;
  assign new_G1635_ = ~new_G1216_ | ~new_G1555_;
  assign new_G1636_ = ~new_G1472_;
  assign new_G1640_ = new_G1176_ & new_G1488_;
  assign new_G1641_ = new_G1062_ & new_G1488_;
  assign new_G1642_ = new_G1067_ & new_G1488_;
  assign new_G1643_ = new_G1187_ & new_G1488_;
  assign new_G1644_ = new_G1152_ & new_G1493_;
  assign new_G1645_ = new_G1159_ & new_G1493_;
  assign new_G1646_ = ~new_G1599_ | ~new_G1600_;
  assign new_G1650_ = ~new_G1537_;
  assign new_G1651_ = ~new_G1537_ | ~new_G1477_;
  assign new_G1652_ = ~new_G1540_ | ~new_G1478_;
  assign new_G1653_ = ~new_G1540_;
  assign new_G1654_ = ~new_G1479_;
  assign new_G1657_ = ~new_G1601_ | ~new_G1602_;
  assign new_G1661_ = ~new_G1557_;
  assign new_G1662_ = ~new_G1557_ | ~new_G1485_;
  assign new_G1663_ = ~new_G1575_;
  assign new_G1664_ = new_G1152_ & new_G1498_;
  assign new_G1665_ = new_G1159_ & new_G1498_;
  assign new_G1666_ = new_G1176_ & new_G1502_;
  assign new_G1667_ = new_G1062_ & new_G1502_;
  assign new_G1668_ = new_G1067_ & new_G1502_;
  assign new_G1669_ = new_G1187_ & new_G1502_;
  assign new_G1670_ = ~new_G1493_;
  assign new_G1675_ = ~new_G1578_;
  assign new_G1676_ = ~new_G1498_;
  assign new_G1681_ = ~new_G1606_ | ~new_G1507_;
  assign new_G1682_ = ~new_G1581_;
  assign new_G1683_ = ~new_G1584_;
  assign new_G1684_ = ~new_G1472_;
  assign new_G1688_ = ~new_G1587_;
  assign new_G1689_ = ~new_G1587_ | ~new_G1427_;
  assign new_G1690_ = ~new_G1628_;
  assign new_G1691_ = ~new_G1627_;
  assign new_G1692_ = ~new_G1626_;
  assign new_G1693_ = ~new_G1625_;
  assign new_G1694_ = ~new_G1624_;
  assign new_G1695_ = ~new_G1623_;
  assign new_G1696_ = ~new_G1622_;
  assign new_G1697_ = ~new_G1621_;
  assign new_G1698_ = ~new_G1620_;
  assign new_G1699_ = ~new_G1619_;
  assign new_G1700_ = ~new_G1634_;
  assign new_G1701_ = ~new_G1633_;
  assign new_G1702_ = ~new_G1632_;
  assign new_G1703_ = ~new_G1631_;
  assign new_G1704_ = ~new_G1630_;
  assign new_G1705_ = ~new_G1629_;
  assign new_G1706_ = ~new_G1520_;
  assign new_G1709_ = ~new_G1524_;
  assign new_G1712_ = ~new_G1528_;
  assign new_G1715_ = ~new_G1528_;
  assign new_G1718_ = ~new_G1596_;
  assign new_G1719_ = ~new_G1596_ | ~new_G1110_;
  assign new_G1720_ = ~new_G1543_;
  assign new_G1721_ = ~new_G1546_;
  assign new_G1722_ = ~new_G1549_;
  assign new_G1723_ = ~new_G1552_;
  assign new_G1724_ = ~new_G1560_;
  assign new_G1725_ = ~new_G1563_;
  assign new_G1726_ = ~new_G1566_;
  assign new_G1727_ = ~new_G1569_;
  assign new_G1728_ = ~new_G1635_ | ~new_G1556_;
  assign new_G1731_ = ~new_G1572_;
  assign new_G1732_ = ~new_G1590_;
  assign new_G1733_ = ~new_G1593_;
  assign new_G1734_ = new_G1421_ & new_G1610_;
  assign new_G1735_ = new_G1418_ & new_G1607_;
  assign new_G1736_ = ~new_G1374_ | ~new_G1650_;
  assign new_G1737_ = ~new_G1377_ | ~new_G1653_;
  assign new_G1738_ = ~new_G1390_ | ~new_G1661_;
  assign new_G1739_ = ~new_G1613_;
  assign new_G1744_ = ~new_G1613_;
  assign new_G1749_ = ~new_G1681_;
  assign new_G1750_ = ~new_G1263_ | ~new_G1688_;
  assign new_G1751_ = new_G1693_ & new_G1690_ & new_G1691_ & new_G1692_ & new_G1694_;
  assign new_G1752_ = new_G1698_ & new_G1695_ & new_G1696_ & new_G1697_ & new_G1699_;
  assign new_G1753_ = new_G1255_ & new_G1700_;
  assign new_G1754_ = new_G1704_ & new_G1701_ & new_G1702_ & new_G1703_ & new_G1705_;
  assign new_G1755_ = ~new_G990_ | ~new_G1718_;
  assign new_G1756_ = ~new_G1616_;
  assign new_G1761_ = ~new_G1616_;
  assign new_G1766_ = ~new_G1546_ | ~new_G1720_;
  assign new_G1767_ = ~new_G1543_ | ~new_G1721_;
  assign new_G1768_ = ~new_G1552_ | ~new_G1722_;
  assign new_G1769_ = ~new_G1549_ | ~new_G1723_;
  assign new_G1770_ = ~new_G1563_ | ~new_G1724_;
  assign new_G1771_ = ~new_G1560_ | ~new_G1725_;
  assign new_G1772_ = ~new_G1569_ | ~new_G1726_;
  assign new_G1773_ = ~new_G1566_ | ~new_G1727_;
  assign new_G1774_ = ~new_G1593_ | ~new_G1732_;
  assign new_G1775_ = ~new_G1590_ | ~new_G1733_;
  assign new_G1776_ = new_G1734_ | new_G1610_;
  assign new_G1777_ = new_G1735_ | new_G1607_;
  assign new_G1778_ = new_G1152_ & new_G1670_;
  assign new_G1779_ = new_G1159_ & new_G1670_;
  assign new_G1780_ = new_G1166_ & new_G1670_;
  assign new_G1781_ = new_G1171_ & new_G1670_;
  assign new_G1782_ = ~new_G1646_;
  assign new_G1785_ = ~new_G1736_ | ~new_G1651_;
  assign new_G1789_ = ~new_G1652_ | ~new_G1737_;
  assign new_G1792_ = ~new_G1657_;
  assign new_G1795_ = ~new_G1738_ | ~new_G1662_;
  assign new_G1798_ = new_G1152_ & new_G1676_;
  assign new_G1799_ = new_G1159_ & new_G1676_;
  assign new_G1800_ = new_G1166_ & new_G1676_;
  assign new_G1801_ = new_G1171_ & new_G1676_;
  assign new_G1802_ = new_G1749_ & n1533_lo;
  assign new_G1805_ = ~new_G1636_;
  assign new_G1811_ = ~new_G1750_ | ~new_G1689_;
  assign new_G1814_ = new_G1751_ & new_G1752_;
  assign new_G1815_ = new_G1753_ & new_G1754_;
  assign new_G1816_ = ~new_G1684_;
  assign new_G1822_ = ~new_G1712_;
  assign new_G1823_ = ~new_G1715_;
  assign new_G1824_ = new_G1524_ & new_G1520_ & new_G1712_;
  assign new_G1825_ = new_G1709_ & new_G1706_ & new_G1715_;
  assign new_G1826_ = ~new_G1755_ | ~new_G1719_;
  assign new_G1829_ = ~new_G1636_;
  assign new_G1835_ = ~new_G1636_;
  assign new_G1840_ = ~new_G1684_;
  assign new_G1846_ = ~new_G1684_;
  assign new_G1851_ = ~new_G1768_ | ~new_G1769_;
  assign new_G1854_ = ~new_G1766_ | ~new_G1767_;
  assign new_G1857_ = ~new_G1728_;
  assign new_G1858_ = ~new_G1728_ | ~new_G1731_;
  assign new_G1859_ = ~new_G1772_ | ~new_G1773_;
  assign new_G1862_ = ~new_G1770_ | ~new_G1771_;
  assign new_G1865_ = ~new_G1774_ | ~new_G1775_;
  assign new_G1868_ = new_G1640_ & new_G1739_;
  assign new_G1869_ = new_G1641_ & new_G1739_;
  assign new_G1870_ = new_G1642_ & new_G1739_;
  assign new_G1871_ = new_G1643_ & new_G1739_;
  assign new_G1872_ = new_G1778_ | new_G1644_;
  assign new_G1873_ = new_G1779_ | new_G1645_;
  assign new_G1874_ = new_G1780_ & new_G598_;
  assign new_G1875_ = new_G1781_ & new_G598_;
  assign new_G1876_ = new_G1798_ | new_G1664_;
  assign new_G1877_ = new_G1799_ | new_G1665_;
  assign new_G1878_ = new_G1800_ & new_G631_;
  assign new_G1879_ = new_G1801_ & new_G631_;
  assign new_G1880_ = new_G1666_ & new_G1744_;
  assign new_G1881_ = new_G1667_ & new_G1744_;
  assign new_G1882_ = new_G1668_ & new_G1744_;
  assign new_G1883_ = new_G1669_ & new_G1744_;
  assign new_G1884_ = new_G1814_ & new_G1815_ & new_G832_;
  assign new_G1887_ = new_G1706_ & new_G1524_ & new_G1822_;
  assign new_G1888_ = new_G1520_ & new_G1709_ & new_G1823_;
  assign new_G1889_ = ~new_G1572_ | ~new_G1857_;
  assign new_G1890_ = ~new_G1868_;
  assign new_G1893_ = ~new_G1869_;
  assign new_G1896_ = ~new_G1870_;
  assign new_G1899_ = ~new_G1871_;
  assign new_G1902_ = new_G1872_ & new_G598_;
  assign new_G1903_ = new_G1873_ & new_G598_;
  assign new_G1904_ = ~new_G1874_;
  assign new_G1907_ = ~new_G1875_;
  assign new_G1910_ = ~new_G1785_;
  assign new_G1913_ = ~new_G1789_;
  assign new_G1916_ = ~new_G1789_;
  assign new_G1919_ = ~new_G1795_;
  assign new_G1922_ = ~new_G1795_;
  assign new_G1925_ = new_G366_ & new_G1805_;
  assign new_G1926_ = new_G1876_ & new_G631_;
  assign new_G1927_ = new_G1877_ & new_G631_;
  assign new_G1928_ = ~new_G1878_;
  assign new_G1931_ = ~new_G1879_;
  assign new_G1934_ = ~new_G1880_;
  assign new_G1937_ = ~new_G1881_;
  assign new_G1940_ = ~new_G1882_;
  assign new_G1943_ = ~new_G1883_;
  assign new_G1946_ = ~new_G1802_;
  assign new_G1947_ = new_G366_ & new_G1816_;
  assign new_G1948_ = ~new_G1805_;
  assign new_G1953_ = new_G370_ & new_G1805_;
  assign new_G1954_ = new_G447_ & new_G1805_;
  assign new_G1955_ = new_G451_ & new_G1805_;
  assign new_G1956_ = ~new_G1816_;
  assign new_G1961_ = new_G370_ & new_G1816_;
  assign new_G1962_ = new_G447_ & new_G1816_;
  assign new_G1963_ = new_G451_ & new_G1816_;
  assign new_G1964_ = ~new_G1887_ & ~new_G1824_;
  assign new_G1965_ = ~new_G1888_ & ~new_G1825_;
  assign new_G1966_ = ~new_G1865_;
  assign new_G1967_ = ~new_G1829_;
  assign new_G1970_ = new_G455_ & new_G1829_;
  assign new_G1971_ = new_G459_ & new_G1829_;
  assign new_G1972_ = new_G463_ & new_G1829_;
  assign new_G1973_ = new_G467_ & new_G1829_;
  assign new_G1974_ = new_G471_ & new_G1835_;
  assign new_G1975_ = new_G475_ & new_G1835_;
  assign new_G1976_ = new_G479_ & new_G1835_;
  assign new_G1977_ = new_G497_ & new_G1835_;
  assign new_G1978_ = ~new_G1840_;
  assign new_G1981_ = new_G455_ & new_G1840_;
  assign new_G1982_ = new_G459_ & new_G1840_;
  assign new_G1983_ = new_G463_ & new_G1840_;
  assign new_G1984_ = new_G467_ & new_G1840_;
  assign new_G1985_ = new_G471_ & new_G1846_;
  assign new_G1986_ = new_G475_ & new_G1846_;
  assign new_G1987_ = new_G479_ & new_G1846_;
  assign new_G1988_ = new_G497_ & new_G1846_;
  assign new_G1989_ = ~new_G1851_;
  assign new_G1990_ = ~new_G1854_;
  assign new_G1991_ = ~new_G1859_;
  assign new_G1992_ = ~new_G1862_;
  assign new_G1993_ = ~new_G1858_ | ~new_G1889_;
  assign new_G1996_ = ~new_G1902_;
  assign new_G1999_ = ~new_G1903_;
  assign new_G2002_ = ~new_G1926_;
  assign new_G2005_ = ~new_G1927_;
  assign new_G2008_ = new_G1972_ & new_G751_;
  assign new_G2011_ = new_G1973_ & new_G751_;
  assign new_G2014_ = new_G1974_ & new_G1756_;
  assign new_G2017_ = new_G1975_ & new_G1756_;
  assign new_G2020_ = new_G1976_ & new_G1756_;
  assign new_G2023_ = new_G1977_ & new_G1756_;
  assign new_G2026_ = new_G1983_ & new_G756_;
  assign new_G2029_ = new_G1984_ & new_G756_;
  assign new_G2032_ = new_G1985_ & new_G1761_;
  assign new_G2035_ = new_G1986_ & new_G1761_;
  assign new_G2038_ = new_G1987_ & new_G1761_;
  assign new_G2041_ = new_G1988_ & new_G1761_;
  assign new_G2044_ = ~new_G1854_ | ~new_G1989_;
  assign new_G2045_ = ~new_G1851_ | ~new_G1990_;
  assign new_G2046_ = ~new_G1862_ | ~new_G1991_;
  assign new_G2047_ = ~new_G1859_ | ~new_G1992_;
  assign new_G2048_ = ~new_G1965_ | ~new_G1964_;
  assign new_G2051_ = ~new_G1913_;
  assign new_G2052_ = ~new_G1916_;
  assign new_G2053_ = ~new_G1919_;
  assign new_G2054_ = ~new_G1922_;
  assign new_G2055_ = new_G1785_ & new_G1646_ & new_G1913_;
  assign new_G2056_ = new_G1910_ & new_G1782_ & new_G1916_;
  assign new_G2057_ = new_G1657_ & new_G1479_ & new_G1919_;
  assign new_G2058_ = new_G1792_ & new_G1654_ & new_G1922_;
  assign new_G2059_ = ~new_G1993_ | ~new_G1486_;
  assign new_G2060_ = ~new_G1993_;
  assign new_G2061_ = new_G479_ & new_G1948_;
  assign new_G2062_ = new_G479_ & new_G1956_;
  assign new_G2063_ = new_G497_ & new_G1948_;
  assign new_G2064_ = new_G503_ & new_G1948_;
  assign new_G2065_ = new_G507_ & new_G1948_;
  assign new_G2066_ = new_G497_ & new_G1956_;
  assign new_G2067_ = new_G503_ & new_G1956_;
  assign new_G2068_ = new_G507_ & new_G1956_;
  assign new_G2069_ = new_G511_ & new_G1967_;
  assign new_G2070_ = new_G515_ & new_G1967_;
  assign new_G2071_ = new_G511_ & new_G1978_;
  assign new_G2072_ = new_G515_ & new_G1978_;
  assign new_G2073_ = ~new_G2044_ | ~new_G2045_;
  assign new_G2076_ = ~new_G2046_ | ~new_G2047_;
  assign new_G2079_ = ~new_G1899_;
  assign new_G2082_ = ~new_G1896_;
  assign new_G2085_ = ~new_G1893_;
  assign new_G2088_ = ~new_G1890_;
  assign new_G2091_ = ~new_G1907_;
  assign new_G2094_ = ~new_G1904_;
  assign new_G2097_ = ~new_G1943_;
  assign new_G2100_ = ~new_G1940_;
  assign new_G2103_ = ~new_G1937_;
  assign new_G2106_ = ~new_G1934_;
  assign new_G2109_ = ~new_G1931_;
  assign new_G2112_ = ~new_G1928_;
  assign new_G2115_ = new_G1782_ & new_G1785_ & new_G2051_;
  assign new_G2116_ = new_G1646_ & new_G1910_ & new_G2052_;
  assign new_G2117_ = new_G1654_ & new_G1657_ & new_G2053_;
  assign new_G2118_ = new_G1479_ & new_G1792_ & new_G2054_;
  assign new_G2119_ = ~new_G1393_ | ~new_G2060_;
  assign new_G2120_ = new_G2061_ | new_G1925_;
  assign new_G2121_ = ~new_G2048_ | ~new_G1966_;
  assign new_G2122_ = new_G2023_ & new_G1899_;
  assign new_G2123_ = new_G2020_ & new_G1896_;
  assign new_G2124_ = new_G2017_ & new_G1893_;
  assign new_G2125_ = new_G1890_ & new_G2014_;
  assign new_G2126_ = new_G2011_ & new_G1907_;
  assign new_G2127_ = new_G2008_ & new_G1904_;
  assign new_G2128_ = new_G2062_ | new_G1947_;
  assign new_G2129_ = new_G2041_ & new_G1943_;
  assign new_G2130_ = new_G2038_ & new_G1940_;
  assign new_G2131_ = new_G2035_ & new_G1937_;
  assign new_G2132_ = new_G1934_ & new_G2032_;
  assign new_G2133_ = new_G2029_ & new_G1931_;
  assign new_G2134_ = new_G2026_ & new_G1928_;
  assign new_G2135_ = new_G2063_ | new_G1953_;
  assign new_G2138_ = new_G2064_ | new_G1954_;
  assign new_G2141_ = new_G2065_ | new_G1955_;
  assign new_G2144_ = new_G2066_ | new_G1961_;
  assign new_G2147_ = new_G2067_ | new_G1962_;
  assign new_G2150_ = new_G2068_ | new_G1963_;
  assign new_G2153_ = ~new_G2048_;
  assign new_G2154_ = new_G2069_ | new_G1970_;
  assign new_G2155_ = new_G2070_ | new_G1971_;
  assign new_G2156_ = new_G2071_ | new_G1981_;
  assign new_G2157_ = new_G2072_ | new_G1982_;
  assign new_G2158_ = ~new_G2023_;
  assign new_G2161_ = ~new_G2020_;
  assign new_G2164_ = ~new_G2017_;
  assign new_G2167_ = ~new_G2014_;
  assign new_G2170_ = ~new_G2011_;
  assign new_G2173_ = ~new_G2008_;
  assign new_G2176_ = ~new_G1999_;
  assign new_G2179_ = ~new_G1996_;
  assign new_G2182_ = ~new_G2041_;
  assign new_G2185_ = ~new_G2038_;
  assign new_G2188_ = ~new_G2035_;
  assign new_G2191_ = ~new_G2032_;
  assign new_G2194_ = ~new_G2029_;
  assign new_G2197_ = ~new_G2026_;
  assign new_G2200_ = ~new_G2005_;
  assign new_G2203_ = ~new_G2002_;
  assign new_G2206_ = ~new_G2059_ | ~new_G2119_;
  assign new_G2207_ = ~new_G2115_ & ~new_G2055_;
  assign new_G2208_ = ~new_G2116_ & ~new_G2056_;
  assign new_G2209_ = ~new_G2117_ & ~new_G2057_;
  assign new_G2210_ = ~new_G2118_ & ~new_G2058_;
  assign new_G2211_ = ~new_G2073_;
  assign new_G2212_ = ~new_G2076_;
  assign new_G2213_ = new_G2120_ & new_G1132_;
  assign new_G2214_ = ~new_G1865_ | ~new_G2153_;
  assign new_G2215_ = ~new_G2079_;
  assign new_G2216_ = ~new_G2082_;
  assign new_G2217_ = ~new_G2085_;
  assign new_G2218_ = ~new_G2088_;
  assign new_G2219_ = ~new_G2091_;
  assign new_G2220_ = ~new_G2094_;
  assign new_G2221_ = new_G2128_ & new_G1132_;
  assign new_G2222_ = ~new_G2097_;
  assign new_G2223_ = ~new_G2100_;
  assign new_G2224_ = ~new_G2103_;
  assign new_G2225_ = ~new_G2106_;
  assign new_G2226_ = ~new_G2109_;
  assign new_G2227_ = ~new_G2112_;
  assign new_G2228_ = new_G2154_ & new_G751_;
  assign new_G2231_ = new_G2155_ & new_G751_;
  assign new_G2234_ = new_G2156_ & new_G756_;
  assign new_G2237_ = new_G2157_ & new_G756_;
  assign new_G2240_ = new_G2206_ & new_G325_;
  assign new_G2241_ = new_G2138_ & new_G1329_;
  assign new_G2242_ = new_G2135_ & new_G1137_;
  assign new_G2243_ = ~new_G2214_ | ~new_G2121_;
  assign new_G2244_ = ~new_G2158_;
  assign new_G2245_ = ~new_G2158_ | ~new_G2215_;
  assign new_G2246_ = ~new_G2161_;
  assign new_G2247_ = ~new_G2161_ | ~new_G2216_;
  assign new_G2248_ = ~new_G2164_;
  assign new_G2249_ = ~new_G2164_ | ~new_G2217_;
  assign new_G2250_ = ~new_G2167_;
  assign new_G2251_ = ~new_G2167_ | ~new_G2218_;
  assign new_G2252_ = ~new_G2170_;
  assign new_G2253_ = ~new_G2170_ | ~new_G2219_;
  assign new_G2254_ = ~new_G2173_;
  assign new_G2255_ = ~new_G2173_ | ~new_G2220_;
  assign new_G2256_ = ~new_G2176_;
  assign new_G2257_ = ~new_G2179_;
  assign new_G2258_ = new_G2141_ & new_G1336_;
  assign new_G2259_ = new_G2147_ & new_G1329_;
  assign new_G2260_ = new_G2144_ & new_G1137_;
  assign new_G2261_ = ~new_G2182_;
  assign new_G2262_ = ~new_G2182_ | ~new_G2222_;
  assign new_G2263_ = ~new_G2185_;
  assign new_G2264_ = ~new_G2185_ | ~new_G2223_;
  assign new_G2265_ = ~new_G2188_;
  assign new_G2266_ = ~new_G2188_ | ~new_G2224_;
  assign new_G2267_ = ~new_G2191_;
  assign new_G2268_ = ~new_G2191_ | ~new_G2225_;
  assign new_G2269_ = ~new_G2194_;
  assign new_G2270_ = ~new_G2194_ | ~new_G2226_;
  assign new_G2271_ = ~new_G2197_;
  assign new_G2272_ = ~new_G2197_ | ~new_G2227_;
  assign new_G2273_ = ~new_G2200_;
  assign new_G2274_ = ~new_G2203_;
  assign new_G2275_ = new_G2150_ & new_G1336_;
  assign new_G2276_ = ~new_G2208_ | ~new_G2207_;
  assign new_G2279_ = ~new_G2210_ | ~new_G2209_;
  assign new_G2282_ = ~new_G2138_;
  assign new_G2285_ = ~new_G2135_;
  assign new_G2288_ = ~new_G2141_;
  assign new_G2291_ = ~new_G2147_;
  assign new_G2294_ = ~new_G2144_;
  assign new_G2297_ = ~new_G2150_;
  assign new_G2300_ = ~new_G2243_;
  assign new_G2301_ = ~new_G2079_ | ~new_G2244_;
  assign new_G2302_ = ~new_G2082_ | ~new_G2246_;
  assign new_G2303_ = ~new_G2085_ | ~new_G2248_;
  assign new_G2304_ = ~new_G2088_ | ~new_G2250_;
  assign new_G2305_ = ~new_G2091_ | ~new_G2252_;
  assign new_G2306_ = ~new_G2094_ | ~new_G2254_;
  assign new_G2307_ = new_G2231_ & new_G1999_;
  assign new_G2308_ = new_G2228_ & new_G1996_;
  assign new_G2309_ = ~new_G2097_ | ~new_G2261_;
  assign new_G2310_ = ~new_G2100_ | ~new_G2263_;
  assign new_G2311_ = ~new_G2103_ | ~new_G2265_;
  assign new_G2312_ = ~new_G2106_ | ~new_G2267_;
  assign new_G2313_ = ~new_G2109_ | ~new_G2269_;
  assign new_G2314_ = ~new_G2112_ | ~new_G2271_;
  assign new_G2315_ = new_G2237_ & new_G2005_;
  assign new_G2316_ = new_G2234_ & new_G2002_;
  assign new_G2317_ = ~new_G2231_;
  assign new_G2320_ = ~new_G2228_;
  assign new_G2323_ = ~new_G2237_;
  assign new_G2326_ = ~new_G2234_;
  assign new_G2329_ = ~new_G2276_;
  assign new_G2330_ = ~new_G2276_ | ~new_G2211_;
  assign new_G2331_ = ~new_G2279_;
  assign new_G2332_ = ~new_G2279_ | ~new_G2212_;
  assign new_G2333_ = ~new_G2282_;
  assign new_G2334_ = ~new_G2282_ | ~new_G1663_;
  assign new_G2335_ = ~new_G2285_ | ~new_G1487_;
  assign new_G2336_ = ~new_G2285_;
  assign new_G2337_ = new_G2300_ & new_G581_;
  assign new_G2340_ = ~new_G2301_ | ~new_G2245_;
  assign new_G2345_ = ~new_G2302_ | ~new_G2247_;
  assign new_G2349_ = ~new_G2303_ | ~new_G2249_;
  assign new_G2352_ = ~new_G2304_ | ~new_G2251_;
  assign new_G2353_ = ~new_G2305_ | ~new_G2253_;
  assign new_G2359_ = ~new_G2306_ | ~new_G2255_;
  assign new_G2364_ = ~new_G2288_;
  assign new_G2365_ = ~new_G2288_ | ~new_G1675_;
  assign new_G2366_ = ~new_G2291_;
  assign new_G2367_ = ~new_G2291_ | ~new_G1682_;
  assign new_G2368_ = ~new_G2294_ | ~new_G1508_;
  assign new_G2369_ = ~new_G2294_;
  assign new_G2370_ = ~new_G2309_ | ~new_G2262_;
  assign new_G2375_ = ~new_G2310_ | ~new_G2264_;
  assign new_G2379_ = ~new_G2311_ | ~new_G2266_;
  assign new_G2382_ = ~new_G2312_ | ~new_G2268_;
  assign new_G2383_ = ~new_G2313_ | ~new_G2270_;
  assign new_G2389_ = ~new_G2314_ | ~new_G2272_;
  assign new_G2394_ = ~new_G2297_;
  assign new_G2395_ = ~new_G2297_ | ~new_G1683_;
  assign new_G2396_ = ~new_G2073_ | ~new_G2329_;
  assign new_G2397_ = ~new_G2076_ | ~new_G2331_;
  assign new_G2398_ = ~new_G1575_ | ~new_G2333_;
  assign new_G2399_ = ~new_G1396_ | ~new_G2336_;
  assign new_G2400_ = ~new_G2317_;
  assign new_G2401_ = ~new_G2317_ | ~new_G2256_;
  assign new_G2402_ = ~new_G2320_;
  assign new_G2403_ = ~new_G2320_ | ~new_G2257_;
  assign new_G2404_ = ~new_G1578_ | ~new_G2364_;
  assign new_G2405_ = ~new_G1581_ | ~new_G2366_;
  assign new_G2406_ = ~new_G1399_ | ~new_G2369_;
  assign new_G2407_ = ~new_G2323_;
  assign new_G2408_ = ~new_G2323_ | ~new_G2273_;
  assign new_G2409_ = ~new_G2326_;
  assign new_G2410_ = ~new_G2326_ | ~new_G2274_;
  assign new_G2411_ = ~new_G1584_ | ~new_G2394_;
  assign new_G2412_ = ~new_G2396_ | ~new_G2330_;
  assign new_G2413_ = ~new_G2397_ | ~new_G2332_;
  assign new_G2414_ = ~new_G2398_ | ~new_G2334_;
  assign new_G2417_ = ~new_G2399_ | ~new_G2335_;
  assign new_G2418_ = ~new_G2337_;
  assign new_G2419_ = ~new_G2176_ | ~new_G2400_;
  assign new_G2420_ = ~new_G2179_ | ~new_G2402_;
  assign new_G2421_ = ~new_G2404_ | ~new_G2365_;
  assign new_G2422_ = new_G2340_ & new_G2345_ & new_G2352_ & new_G2349_;
  assign new_G2423_ = new_G2340_ & new_G2123_;
  assign new_G2424_ = new_G2345_ & new_G2340_ & new_G2124_;
  assign new_G2425_ = new_G2345_ & new_G2349_ & new_G2340_ & new_G2125_;
  assign new_G2426_ = new_G2353_ & new_G2127_;
  assign new_G2427_ = new_G2359_ & new_G2353_ & new_G2307_;
  assign new_G2428_ = ~new_G2405_ | ~new_G2367_;
  assign new_G2431_ = ~new_G2406_ | ~new_G2368_;
  assign new_G2432_ = ~new_G2200_ | ~new_G2407_;
  assign new_G2433_ = ~new_G2203_ | ~new_G2409_;
  assign new_G2434_ = ~new_G2411_ | ~new_G2395_;
  assign new_G2435_ = new_G2370_ & new_G2375_ & new_G2382_ & new_G2379_;
  assign new_G2436_ = new_G2370_ & new_G2130_;
  assign new_G2437_ = new_G2375_ & new_G2370_ & new_G2131_;
  assign new_G2438_ = new_G2375_ & new_G2379_ & new_G2370_ & new_G2132_;
  assign new_G2439_ = new_G2383_ & new_G2134_;
  assign new_G2440_ = new_G2389_ & new_G2383_ & new_G2315_;
  assign new_G2441_ = ~new_G2412_;
  assign new_G2442_ = new_G2413_ & n2889_lo;
  assign new_G2443_ = ~new_G2419_ | ~new_G2401_;
  assign new_G2447_ = ~new_G2420_ | ~new_G2403_;
  assign new_G2450_ = ~new_G2422_;
  assign new_G2451_ = new_G2425_ | new_G2424_ | new_G2122_ | new_G2423_;
  assign new_G2454_ = ~new_G2432_ | ~new_G2408_;
  assign new_G2458_ = ~new_G2433_ | ~new_G2410_;
  assign new_G2461_ = ~new_G2435_;
  assign new_G2462_ = new_G2438_ | new_G2437_ | new_G2129_ | new_G2436_;
  assign new_G2465_ = new_G2414_ & new_G2242_;
  assign new_G2466_ = new_G2417_ & new_G2414_ & new_G2213_;
  assign new_G2467_ = new_G1326_ | new_G2442_;
  assign new_G2470_ = new_G2441_ & new_G581_;
  assign new_G2473_ = new_G2428_ & new_G2260_;
  assign new_G2474_ = new_G2431_ & new_G2428_ & new_G2221_;
  assign new_G2475_ = new_G2466_ | new_G2241_ | new_G2465_;
  assign new_G2476_ = ~new_G2451_;
  assign new_G2477_ = new_G2353_ & new_G2359_ & new_G2421_ & new_G2443_ & new_G2447_;
  assign new_G2478_ = new_G2359_ & new_G2443_ & new_G2353_ & new_G2308_;
  assign new_G2479_ = new_G2258_ & new_G2447_ & new_G2443_ & new_G2353_ & new_G2359_;
  assign new_G2480_ = new_G2474_ | new_G2259_ | new_G2473_;
  assign new_G2481_ = ~new_G2462_;
  assign new_G2482_ = new_G2383_ & new_G2389_ & new_G2434_ & new_G2454_ & new_G2458_;
  assign new_G2483_ = new_G2389_ & new_G2454_ & new_G2383_ & new_G2316_;
  assign new_G2484_ = new_G2275_ & new_G2458_ & new_G2454_ & new_G2383_ & new_G2389_;
  assign new_G2485_ = new_G2478_ | new_G2427_ | new_G2126_ | new_G2426_ | new_G2479_;
  assign new_G2486_ = new_G2477_ & new_G2475_;
  assign new_G2487_ = ~new_G2476_ | ~new_G2450_;
  assign new_G2488_ = ~new_G2470_;
  assign new_G2489_ = new_G2483_ | new_G2440_ | new_G2133_ | new_G2439_ | new_G2484_;
  assign new_G2490_ = new_G2482_ & new_G2480_;
  assign new_G2491_ = ~new_G2481_ | ~new_G2461_;
  assign new_G2492_ = new_G2485_ | new_G2486_;
  assign new_G2495_ = new_G2418_ & new_G2488_ & new_G1826_;
  assign new_G2496_ = new_G2489_ | new_G2490_;
  assign new_G2499_ = ~new_G2492_;
  assign new_G2500_ = new_G2487_ & new_G2492_;
  assign new_G2501_ = ~new_G2496_;
  assign new_G2502_ = new_G2491_ & new_G2496_;
  assign new_G2503_ = new_G2451_ & new_G2499_;
  assign new_G2504_ = new_G2462_ & new_G2501_;
  assign new_G2505_ = new_G2503_ | new_G2500_;
  assign new_G2508_ = new_G2504_ | new_G2502_;
  assign new_G2512_ = ~new_G2508_ | ~new_G2505_;
  assign new_G2515_ = new_G2508_ & new_G2512_;
  assign new_G2516_ = new_G2512_ & new_G2505_;
  assign new_G2517_ = new_G2515_ | new_G2516_;
  assign new_G2520_ = ~new_G2517_;
  assign new_G2523_ = new_G2517_ & new_G2520_;
  assign new_G2524_ = new_G2523_ | new_G2520_;
  assign new_G2527_ = new_G1811_ & new_G1946_ & new_G2524_;
  assign new_G2528_ = new_G2495_ & new_G2527_ & new_G993_;
  assign G2531 = ~n2793_lo;
  assign G2532 = G2531;
  assign G2533 = G2531;
  assign G2534 = ~n2901_lo;
  assign G2535 = G2534;
  assign G2536 = ~n3057_lo;
  assign G2537 = G2536;
  assign G2538 = G2536;
  assign G2539 = ~n1797_lo;
  assign G2540 = ~n2685_lo;
  assign G2541 = ~n2181_lo;
  assign G2542 = ~n2325_lo;
  assign G2543 = ~n2049_lo;
  assign G2544 = ~n2565_lo;
  assign G2545 = ~n1929_lo;
  assign G2546 = ~n2445_lo;
  assign G2547 = ~new_G285_;
  assign G2548 = ~new_G287_;
  assign G2549 = ~new_G292_;
  assign G2550 = n2301_lo & new_G292_;
  assign G2551 = ~new_G443_;
  assign G2552 = ~n2841_lo | ~new_G443_;
  assign G2553 = ~new_G592_;
  assign G2554 = ~new_G595_;
  assign G2555 = G2554;
  assign G2556 = ~new_G993_;
  assign G2557 = ~new_G1044_;
  assign G2558 = ~new_G1049_;
  assign G2559 = ~new_G1039_;
  assign G2560 = ~new_G1026_;
  assign G2561 = ~new_G1021_;
  assign G2562 = ~new_G1017_;
  assign G2563 = new_G325_ | new_G1117_;
  assign G2564 = ~new_G1118_;
  assign G2565 = ~new_G1119_;
  assign G2566 = ~new_G1144_;
  assign G2567 = ~new_G1148_;
  assign G2568 = ~new_G1152_;
  assign G2569 = ~new_G1159_;
  assign G2570 = ~new_G1166_;
  assign G2571 = ~new_G1171_;
  assign G2572 = ~new_G1176_;
  assign G2573 = ~new_G1412_;
  assign G2574 = G2573;
  assign G2575 = ~new_G1415_;
  assign G2576 = G2575;
  assign G2577 = new_G1471_ | new_G1116_;
  assign G2578 = ~new_G1603_;
  assign G2579 = G2578;
  assign G2580 = ~new_G1776_ | ~new_G1777_;
  assign G2581 = ~new_G1802_;
  assign G2582 = ~new_G1826_;
  assign G2583 = ~new_G1811_;
  assign G2584 = ~new_G1884_;
  assign G2585 = G2584;
  assign G2586 = new_G2240_ | new_G1115_;
  assign G2587 = ~new_G2337_;
  assign G2588 = ~new_G2467_;
  assign G2589 = G2588;
  assign G2590 = ~new_G2470_;
  assign G2591 = ~new_G2508_;
  assign G2592 = ~new_G2524_;
  assign G2593 = ~new_G2528_;
  assign G2594 = G2593;
  assign n1416_li = G1;
  assign n1419_li = n1416_lo;
  assign n1422_li = n1419_lo;
  assign n1425_li = n1422_lo;
  assign n1428_li = G2;
  assign n1431_li = n1428_lo;
  assign n1434_li = n1431_lo;
  assign n1437_li = n1434_lo;
  assign n1440_li = G3;
  assign n1443_li = n1440_lo;
  assign n1446_li = n1443_lo;
  assign n1449_li = n1446_lo;
  assign n1452_li = G4;
  assign n1455_li = n1452_lo;
  assign n1458_li = n1455_lo;
  assign n1461_li = n1458_lo;
  assign n1464_li = G5;
  assign n1467_li = n1464_lo;
  assign n1470_li = n1467_lo;
  assign n1473_li = n1470_lo;
  assign n1476_li = G6;
  assign n1479_li = n1476_lo;
  assign n1482_li = n1479_lo;
  assign n1485_li = n1482_lo;
  assign n1488_li = G7;
  assign n1491_li = n1488_lo;
  assign n1494_li = n1491_lo;
  assign n1497_li = n1494_lo;
  assign n1500_li = G8;
  assign n1503_li = n1500_lo;
  assign n1506_li = n1503_lo;
  assign n1509_li = n1506_lo;
  assign n1512_li = G9;
  assign n1515_li = n1512_lo;
  assign n1518_li = n1515_lo;
  assign n1521_li = n1518_lo;
  assign n1524_li = G10;
  assign n1527_li = n1524_lo;
  assign n1530_li = n1527_lo;
  assign n1533_li = n1530_lo;
  assign n1536_li = G11;
  assign n1539_li = n1536_lo;
  assign n1542_li = n1539_lo;
  assign n1545_li = n1542_lo;
  assign n1548_li = G12;
  assign n1551_li = n1548_lo;
  assign n1554_li = n1551_lo;
  assign n1557_li = n1554_lo;
  assign n1560_li = G13;
  assign n1563_li = n1560_lo;
  assign n1566_li = n1563_lo;
  assign n1569_li = n1566_lo;
  assign n1572_li = G14;
  assign n1575_li = n1572_lo;
  assign n1578_li = n1575_lo;
  assign n1581_li = n1578_lo;
  assign n1584_li = G15;
  assign n1587_li = n1584_lo;
  assign n1590_li = n1587_lo;
  assign n1593_li = n1590_lo;
  assign n1596_li = G16;
  assign n1599_li = n1596_lo;
  assign n1602_li = n1599_lo;
  assign n1605_li = n1602_lo;
  assign n1608_li = G17;
  assign n1611_li = n1608_lo;
  assign n1614_li = n1611_lo;
  assign n1617_li = n1614_lo;
  assign n1620_li = G18;
  assign n1623_li = n1620_lo;
  assign n1626_li = n1623_lo;
  assign n1629_li = n1626_lo;
  assign n1632_li = G19;
  assign n1635_li = n1632_lo;
  assign n1638_li = n1635_lo;
  assign n1641_li = n1638_lo;
  assign n1644_li = G20;
  assign n1647_li = n1644_lo;
  assign n1650_li = n1647_lo;
  assign n1653_li = n1650_lo;
  assign n1656_li = G21;
  assign n1659_li = n1656_lo;
  assign n1662_li = n1659_lo;
  assign n1665_li = n1662_lo;
  assign n1668_li = G22;
  assign n1671_li = n1668_lo;
  assign n1674_li = n1671_lo;
  assign n1677_li = n1674_lo;
  assign n1680_li = G23;
  assign n1683_li = n1680_lo;
  assign n1686_li = n1683_lo;
  assign n1689_li = n1686_lo;
  assign n1692_li = G24;
  assign n1695_li = n1692_lo;
  assign n1698_li = n1695_lo;
  assign n1701_li = n1698_lo;
  assign n1704_li = G25;
  assign n1707_li = n1704_lo;
  assign n1710_li = n1707_lo;
  assign n1713_li = n1710_lo;
  assign n1716_li = G26;
  assign n1719_li = n1716_lo;
  assign n1722_li = n1719_lo;
  assign n1725_li = n1722_lo;
  assign n1728_li = G27;
  assign n1731_li = n1728_lo;
  assign n1734_li = n1731_lo;
  assign n1737_li = n1734_lo;
  assign n1740_li = G28;
  assign n1743_li = n1740_lo;
  assign n1746_li = n1743_lo;
  assign n1749_li = n1746_lo;
  assign n1752_li = G29;
  assign n1755_li = n1752_lo;
  assign n1758_li = n1755_lo;
  assign n1761_li = n1758_lo;
  assign n1764_li = G30;
  assign n1767_li = n1764_lo;
  assign n1770_li = n1767_lo;
  assign n1773_li = n1770_lo;
  assign n1776_li = G31;
  assign n1779_li = n1776_lo;
  assign n1782_li = n1779_lo;
  assign n1785_li = n1782_lo;
  assign n1788_li = G32;
  assign n1791_li = n1788_lo;
  assign n1794_li = n1791_lo;
  assign n1797_li = n1794_lo;
  assign n1800_li = G33;
  assign n1803_li = n1800_lo;
  assign n1806_li = n1803_lo;
  assign n1809_li = n1806_lo;
  assign n1812_li = G34;
  assign n1815_li = n1812_lo;
  assign n1818_li = n1815_lo;
  assign n1821_li = n1818_lo;
  assign n1824_li = G35;
  assign n1827_li = n1824_lo;
  assign n1830_li = n1827_lo;
  assign n1833_li = n1830_lo;
  assign n1836_li = G36;
  assign n1839_li = n1836_lo;
  assign n1842_li = n1839_lo;
  assign n1845_li = n1842_lo;
  assign n1848_li = G37;
  assign n1851_li = n1848_lo;
  assign n1854_li = n1851_lo;
  assign n1857_li = n1854_lo;
  assign n1860_li = G38;
  assign n1863_li = n1860_lo;
  assign n1866_li = n1863_lo;
  assign n1869_li = n1866_lo;
  assign n1872_li = G39;
  assign n1875_li = n1872_lo;
  assign n1878_li = n1875_lo;
  assign n1881_li = n1878_lo;
  assign n1884_li = G40;
  assign n1887_li = n1884_lo;
  assign n1890_li = n1887_lo;
  assign n1893_li = n1890_lo;
  assign n1896_li = G41;
  assign n1899_li = n1896_lo;
  assign n1902_li = n1899_lo;
  assign n1905_li = n1902_lo;
  assign n1908_li = G42;
  assign n1911_li = n1908_lo;
  assign n1914_li = n1911_lo;
  assign n1917_li = n1914_lo;
  assign n1920_li = G43;
  assign n1923_li = n1920_lo;
  assign n1926_li = n1923_lo;
  assign n1929_li = n1926_lo;
  assign n1932_li = G44;
  assign n1935_li = n1932_lo;
  assign n1938_li = n1935_lo;
  assign n1941_li = n1938_lo;
  assign n1944_li = G45;
  assign n1947_li = n1944_lo;
  assign n1950_li = n1947_lo;
  assign n1953_li = n1950_lo;
  assign n1956_li = G46;
  assign n1959_li = n1956_lo;
  assign n1962_li = n1959_lo;
  assign n1965_li = n1962_lo;
  assign n1968_li = G47;
  assign n1971_li = n1968_lo;
  assign n1974_li = n1971_lo;
  assign n1977_li = n1974_lo;
  assign n1980_li = G48;
  assign n1983_li = n1980_lo;
  assign n1986_li = n1983_lo;
  assign n1989_li = n1986_lo;
  assign n1992_li = G49;
  assign n1995_li = n1992_lo;
  assign n1998_li = n1995_lo;
  assign n2001_li = n1998_lo;
  assign n2004_li = G50;
  assign n2007_li = n2004_lo;
  assign n2010_li = n2007_lo;
  assign n2013_li = n2010_lo;
  assign n2016_li = G51;
  assign n2019_li = n2016_lo;
  assign n2022_li = n2019_lo;
  assign n2025_li = n2022_lo;
  assign n2028_li = G52;
  assign n2031_li = n2028_lo;
  assign n2034_li = n2031_lo;
  assign n2037_li = n2034_lo;
  assign n2040_li = G53;
  assign n2043_li = n2040_lo;
  assign n2046_li = n2043_lo;
  assign n2049_li = n2046_lo;
  assign n2052_li = G54;
  assign n2055_li = n2052_lo;
  assign n2058_li = n2055_lo;
  assign n2061_li = n2058_lo;
  assign n2064_li = G55;
  assign n2067_li = n2064_lo;
  assign n2070_li = n2067_lo;
  assign n2073_li = n2070_lo;
  assign n2076_li = G56;
  assign n2079_li = n2076_lo;
  assign n2082_li = n2079_lo;
  assign n2085_li = n2082_lo;
  assign n2088_li = G57;
  assign n2091_li = n2088_lo;
  assign n2094_li = n2091_lo;
  assign n2097_li = n2094_lo;
  assign n2100_li = G58;
  assign n2103_li = n2100_lo;
  assign n2106_li = n2103_lo;
  assign n2109_li = n2106_lo;
  assign n2112_li = G59;
  assign n2115_li = n2112_lo;
  assign n2118_li = n2115_lo;
  assign n2121_li = n2118_lo;
  assign n2124_li = G60;
  assign n2127_li = n2124_lo;
  assign n2130_li = n2127_lo;
  assign n2133_li = n2130_lo;
  assign n2136_li = G61;
  assign n2139_li = n2136_lo;
  assign n2142_li = n2139_lo;
  assign n2145_li = n2142_lo;
  assign n2148_li = G62;
  assign n2151_li = n2148_lo;
  assign n2154_li = n2151_lo;
  assign n2157_li = n2154_lo;
  assign n2160_li = G63;
  assign n2163_li = n2160_lo;
  assign n2166_li = n2163_lo;
  assign n2169_li = n2166_lo;
  assign n2172_li = G64;
  assign n2175_li = n2172_lo;
  assign n2178_li = n2175_lo;
  assign n2181_li = n2178_lo;
  assign n2184_li = G65;
  assign n2187_li = n2184_lo;
  assign n2190_li = n2187_lo;
  assign n2193_li = n2190_lo;
  assign n2196_li = G66;
  assign n2199_li = n2196_lo;
  assign n2202_li = n2199_lo;
  assign n2205_li = n2202_lo;
  assign n2208_li = G67;
  assign n2211_li = n2208_lo;
  assign n2214_li = n2211_lo;
  assign n2217_li = n2214_lo;
  assign n2220_li = G68;
  assign n2223_li = n2220_lo;
  assign n2226_li = n2223_lo;
  assign n2229_li = n2226_lo;
  assign n2232_li = G69;
  assign n2235_li = n2232_lo;
  assign n2238_li = n2235_lo;
  assign n2241_li = n2238_lo;
  assign n2244_li = G70;
  assign n2247_li = n2244_lo;
  assign n2250_li = n2247_lo;
  assign n2253_li = n2250_lo;
  assign n2256_li = G71;
  assign n2259_li = n2256_lo;
  assign n2262_li = n2259_lo;
  assign n2265_li = n2262_lo;
  assign n2268_li = G72;
  assign n2271_li = n2268_lo;
  assign n2274_li = n2271_lo;
  assign n2277_li = n2274_lo;
  assign n2280_li = G73;
  assign n2283_li = n2280_lo;
  assign n2286_li = n2283_lo;
  assign n2289_li = n2286_lo;
  assign n2292_li = G74;
  assign n2295_li = n2292_lo;
  assign n2298_li = n2295_lo;
  assign n2301_li = n2298_lo;
  assign n2304_li = G75;
  assign n2307_li = n2304_lo;
  assign n2310_li = n2307_lo;
  assign n2313_li = n2310_lo;
  assign n2316_li = G76;
  assign n2319_li = n2316_lo;
  assign n2322_li = n2319_lo;
  assign n2325_li = n2322_lo;
  assign n2328_li = G77;
  assign n2331_li = n2328_lo;
  assign n2334_li = n2331_lo;
  assign n2337_li = n2334_lo;
  assign n2340_li = G78;
  assign n2343_li = n2340_lo;
  assign n2346_li = n2343_lo;
  assign n2349_li = n2346_lo;
  assign n2352_li = G79;
  assign n2355_li = n2352_lo;
  assign n2358_li = n2355_lo;
  assign n2361_li = n2358_lo;
  assign n2364_li = G80;
  assign n2367_li = n2364_lo;
  assign n2370_li = n2367_lo;
  assign n2373_li = n2370_lo;
  assign n2376_li = G81;
  assign n2379_li = n2376_lo;
  assign n2382_li = n2379_lo;
  assign n2385_li = n2382_lo;
  assign n2388_li = G82;
  assign n2391_li = n2388_lo;
  assign n2394_li = n2391_lo;
  assign n2397_li = n2394_lo;
  assign n2400_li = G83;
  assign n2403_li = n2400_lo;
  assign n2406_li = n2403_lo;
  assign n2409_li = n2406_lo;
  assign n2412_li = G84;
  assign n2415_li = n2412_lo;
  assign n2418_li = n2415_lo;
  assign n2421_li = n2418_lo;
  assign n2424_li = G85;
  assign n2427_li = n2424_lo;
  assign n2430_li = n2427_lo;
  assign n2433_li = n2430_lo;
  assign n2436_li = G86;
  assign n2439_li = n2436_lo;
  assign n2442_li = n2439_lo;
  assign n2445_li = n2442_lo;
  assign n2448_li = G87;
  assign n2451_li = n2448_lo;
  assign n2454_li = n2451_lo;
  assign n2457_li = n2454_lo;
  assign n2460_li = G88;
  assign n2463_li = n2460_lo;
  assign n2466_li = n2463_lo;
  assign n2469_li = n2466_lo;
  assign n2472_li = G89;
  assign n2475_li = n2472_lo;
  assign n2478_li = n2475_lo;
  assign n2481_li = n2478_lo;
  assign n2484_li = G90;
  assign n2487_li = n2484_lo;
  assign n2490_li = n2487_lo;
  assign n2493_li = n2490_lo;
  assign n2496_li = G91;
  assign n2499_li = n2496_lo;
  assign n2502_li = n2499_lo;
  assign n2505_li = n2502_lo;
  assign n2508_li = G92;
  assign n2511_li = n2508_lo;
  assign n2514_li = n2511_lo;
  assign n2517_li = n2514_lo;
  assign n2520_li = G93;
  assign n2523_li = n2520_lo;
  assign n2526_li = n2523_lo;
  assign n2529_li = n2526_lo;
  assign n2532_li = G94;
  assign n2535_li = n2532_lo;
  assign n2538_li = n2535_lo;
  assign n2541_li = n2538_lo;
  assign n2544_li = G95;
  assign n2547_li = n2544_lo;
  assign n2550_li = n2547_lo;
  assign n2553_li = n2550_lo;
  assign n2556_li = G96;
  assign n2559_li = n2556_lo;
  assign n2562_li = n2559_lo;
  assign n2565_li = n2562_lo;
  assign n2568_li = G97;
  assign n2571_li = n2568_lo;
  assign n2574_li = n2571_lo;
  assign n2577_li = n2574_lo;
  assign n2580_li = G98;
  assign n2583_li = n2580_lo;
  assign n2586_li = n2583_lo;
  assign n2589_li = n2586_lo;
  assign n2592_li = G99;
  assign n2595_li = n2592_lo;
  assign n2598_li = n2595_lo;
  assign n2601_li = n2598_lo;
  assign n2604_li = G100;
  assign n2607_li = n2604_lo;
  assign n2610_li = n2607_lo;
  assign n2613_li = n2610_lo;
  assign n2616_li = G101;
  assign n2619_li = n2616_lo;
  assign n2622_li = n2619_lo;
  assign n2625_li = n2622_lo;
  assign n2628_li = G102;
  assign n2631_li = n2628_lo;
  assign n2634_li = n2631_lo;
  assign n2637_li = n2634_lo;
  assign n2640_li = G103;
  assign n2643_li = n2640_lo;
  assign n2646_li = n2643_lo;
  assign n2649_li = n2646_lo;
  assign n2652_li = G104;
  assign n2655_li = n2652_lo;
  assign n2658_li = n2655_lo;
  assign n2661_li = n2658_lo;
  assign n2664_li = G105;
  assign n2667_li = n2664_lo;
  assign n2670_li = n2667_lo;
  assign n2673_li = n2670_lo;
  assign n2676_li = G106;
  assign n2679_li = n2676_lo;
  assign n2682_li = n2679_lo;
  assign n2685_li = n2682_lo;
  assign n2688_li = G107;
  assign n2691_li = n2688_lo;
  assign n2694_li = n2691_lo;
  assign n2697_li = n2694_lo;
  assign n2700_li = G108;
  assign n2703_li = n2700_lo;
  assign n2706_li = n2703_lo;
  assign n2709_li = n2706_lo;
  assign n2712_li = G109;
  assign n2715_li = n2712_lo;
  assign n2718_li = n2715_lo;
  assign n2721_li = n2718_lo;
  assign n2724_li = G110;
  assign n2727_li = n2724_lo;
  assign n2730_li = n2727_lo;
  assign n2733_li = n2730_lo;
  assign n2736_li = G111;
  assign n2739_li = n2736_lo;
  assign n2742_li = n2739_lo;
  assign n2745_li = n2742_lo;
  assign n2748_li = G112;
  assign n2751_li = n2748_lo;
  assign n2754_li = n2751_lo;
  assign n2757_li = n2754_lo;
  assign n2760_li = G113;
  assign n2763_li = n2760_lo;
  assign n2766_li = n2763_lo;
  assign n2769_li = n2766_lo;
  assign n2772_li = G114;
  assign n2775_li = n2772_lo;
  assign n2778_li = n2775_lo;
  assign n2781_li = n2778_lo;
  assign n2784_li = G115;
  assign n2787_li = n2784_lo;
  assign n2790_li = n2787_lo;
  assign n2793_li = n2790_lo;
  assign n2796_li = G116;
  assign n2799_li = n2796_lo;
  assign n2802_li = n2799_lo;
  assign n2805_li = n2802_lo;
  assign n2808_li = G117;
  assign n2811_li = n2808_lo;
  assign n2814_li = n2811_lo;
  assign n2817_li = n2814_lo;
  assign n2820_li = G118;
  assign n2823_li = n2820_lo;
  assign n2826_li = n2823_lo;
  assign n2829_li = n2826_lo;
  assign n2832_li = G119;
  assign n2835_li = n2832_lo;
  assign n2838_li = n2835_lo;
  assign n2841_li = n2838_lo;
  assign n2844_li = G120;
  assign n2847_li = n2844_lo;
  assign n2850_li = n2847_lo;
  assign n2853_li = n2850_lo;
  assign n2856_li = G121;
  assign n2859_li = n2856_lo;
  assign n2862_li = n2859_lo;
  assign n2865_li = n2862_lo;
  assign n2868_li = G122;
  assign n2871_li = n2868_lo;
  assign n2874_li = n2871_lo;
  assign n2877_li = n2874_lo;
  assign n2880_li = G123;
  assign n2883_li = n2880_lo;
  assign n2886_li = n2883_lo;
  assign n2889_li = n2886_lo;
  assign n2892_li = G124;
  assign n2895_li = n2892_lo;
  assign n2898_li = n2895_lo;
  assign n2901_li = n2898_lo;
  assign n2904_li = G125;
  assign n2907_li = n2904_lo;
  assign n2910_li = n2907_lo;
  assign n2913_li = n2910_lo;
  assign n2916_li = G126;
  assign n2919_li = n2916_lo;
  assign n2922_li = n2919_lo;
  assign n2925_li = n2922_lo;
  assign n2928_li = G127;
  assign n2931_li = n2928_lo;
  assign n2934_li = n2931_lo;
  assign n2937_li = n2934_lo;
  assign n2940_li = G128;
  assign n2943_li = n2940_lo;
  assign n2946_li = n2943_lo;
  assign n2949_li = n2946_lo;
  assign n2952_li = G129;
  assign n2955_li = n2952_lo;
  assign n2958_li = n2955_lo;
  assign n2961_li = n2958_lo;
  assign n2964_li = G130;
  assign n2967_li = n2964_lo;
  assign n2970_li = n2967_lo;
  assign n2973_li = n2970_lo;
  assign n2976_li = G131;
  assign n2979_li = n2976_lo;
  assign n2982_li = n2979_lo;
  assign n2985_li = n2982_lo;
  assign n2988_li = G132;
  assign n2991_li = n2988_lo;
  assign n2994_li = n2991_lo;
  assign n2997_li = n2994_lo;
  assign n3000_li = G133;
  assign n3003_li = n3000_lo;
  assign n3006_li = n3003_lo;
  assign n3009_li = n3006_lo;
  assign n3012_li = G134;
  assign n3015_li = n3012_lo;
  assign n3018_li = n3015_lo;
  assign n3021_li = n3018_lo;
  assign n3024_li = G135;
  assign n3027_li = n3024_lo;
  assign n3030_li = n3027_lo;
  assign n3033_li = n3030_lo;
  assign n3036_li = G136;
  assign n3039_li = n3036_lo;
  assign n3042_li = n3039_lo;
  assign n3045_li = n3042_lo;
  assign n3048_li = G137;
  assign n3051_li = n3048_lo;
  assign n3054_li = n3051_lo;
  assign n3057_li = n3054_lo;
  assign n3060_li = G138;
  assign n3063_li = n3060_lo;
  assign n3066_li = n3063_lo;
  assign n3069_li = n3066_lo;
  assign n3072_li = G139;
  assign n3075_li = n3072_lo;
  assign n3078_li = n3075_lo;
  assign n3081_li = n3078_lo;
  assign n3084_li = G140;
  assign n3087_li = n3084_lo;
  assign n3090_li = n3087_lo;
  assign n3093_li = n3090_lo;
  assign n3096_li = G141;
  assign n3099_li = n3096_lo;
  assign n3102_li = n3099_lo;
  assign n3105_li = n3102_lo;
  assign n3108_li = G142;
  assign n3111_li = n3108_lo;
  assign n3114_li = n3111_lo;
  assign n3117_li = n3114_lo;
  assign n3120_li = G143;
  assign n3123_li = n3120_lo;
  assign n3126_li = n3123_lo;
  assign n3129_li = n3126_lo;
  assign n3132_li = G144;
  assign n3135_li = n3132_lo;
  assign n3138_li = n3135_lo;
  assign n3141_li = n3138_lo;
  assign n3144_li = G145;
  assign n3147_li = n3144_lo;
  assign n3150_li = n3147_lo;
  assign n3153_li = n3150_lo;
  assign n3156_li = G146;
  assign n3159_li = n3156_lo;
  assign n3162_li = n3159_lo;
  assign n3165_li = n3162_lo;
  assign n3168_li = G147;
  assign n3171_li = n3168_lo;
  assign n3174_li = n3171_lo;
  assign n3177_li = n3174_lo;
  assign n3180_li = G148;
  assign n3183_li = n3180_lo;
  assign n3186_li = n3183_lo;
  assign n3189_li = n3186_lo;
  assign n3192_li = G149;
  assign n3195_li = n3192_lo;
  assign n3198_li = n3195_lo;
  assign n3201_li = n3198_lo;
  assign n3204_li = G150;
  assign n3207_li = n3204_lo;
  assign n3210_li = n3207_lo;
  assign n3213_li = n3210_lo;
  assign n3216_li = G151;
  assign n3219_li = n3216_lo;
  assign n3222_li = n3219_lo;
  assign n3225_li = n3222_lo;
  assign n3228_li = G152;
  assign n3231_li = n3228_lo;
  assign n3234_li = n3231_lo;
  assign n3237_li = n3234_lo;
  assign n3240_li = G153;
  assign n3243_li = n3240_lo;
  assign n3246_li = n3243_lo;
  assign n3249_li = n3246_lo;
  assign n3252_li = G154;
  assign n3255_li = n3252_lo;
  assign n3258_li = n3255_lo;
  assign n3261_li = n3258_lo;
  assign n3264_li = G155;
  assign n3267_li = n3264_lo;
  assign n3270_li = n3267_lo;
  assign n3273_li = n3270_lo;
  assign n3276_li = G156;
  assign n3279_li = n3276_lo;
  assign n3282_li = n3279_lo;
  assign n3285_li = n3282_lo;
  assign n3288_li = G157;
  assign n3291_li = n3288_lo;
  assign n3294_li = n3291_lo;
  assign n3297_li = n3294_lo;
  always @ (posedge clock) begin
    n1416_lo <= n1416_li;
    n1419_lo <= n1419_li;
    n1422_lo <= n1422_li;
    n1425_lo <= n1425_li;
    n1428_lo <= n1428_li;
    n1431_lo <= n1431_li;
    n1434_lo <= n1434_li;
    n1437_lo <= n1437_li;
    n1440_lo <= n1440_li;
    n1443_lo <= n1443_li;
    n1446_lo <= n1446_li;
    n1449_lo <= n1449_li;
    n1452_lo <= n1452_li;
    n1455_lo <= n1455_li;
    n1458_lo <= n1458_li;
    n1461_lo <= n1461_li;
    n1464_lo <= n1464_li;
    n1467_lo <= n1467_li;
    n1470_lo <= n1470_li;
    n1473_lo <= n1473_li;
    n1476_lo <= n1476_li;
    n1479_lo <= n1479_li;
    n1482_lo <= n1482_li;
    n1485_lo <= n1485_li;
    n1488_lo <= n1488_li;
    n1491_lo <= n1491_li;
    n1494_lo <= n1494_li;
    n1497_lo <= n1497_li;
    n1500_lo <= n1500_li;
    n1503_lo <= n1503_li;
    n1506_lo <= n1506_li;
    n1509_lo <= n1509_li;
    n1512_lo <= n1512_li;
    n1515_lo <= n1515_li;
    n1518_lo <= n1518_li;
    n1521_lo <= n1521_li;
    n1524_lo <= n1524_li;
    n1527_lo <= n1527_li;
    n1530_lo <= n1530_li;
    n1533_lo <= n1533_li;
    n1536_lo <= n1536_li;
    n1539_lo <= n1539_li;
    n1542_lo <= n1542_li;
    n1545_lo <= n1545_li;
    n1548_lo <= n1548_li;
    n1551_lo <= n1551_li;
    n1554_lo <= n1554_li;
    n1557_lo <= n1557_li;
    n1560_lo <= n1560_li;
    n1563_lo <= n1563_li;
    n1566_lo <= n1566_li;
    n1569_lo <= n1569_li;
    n1572_lo <= n1572_li;
    n1575_lo <= n1575_li;
    n1578_lo <= n1578_li;
    n1581_lo <= n1581_li;
    n1584_lo <= n1584_li;
    n1587_lo <= n1587_li;
    n1590_lo <= n1590_li;
    n1593_lo <= n1593_li;
    n1596_lo <= n1596_li;
    n1599_lo <= n1599_li;
    n1602_lo <= n1602_li;
    n1605_lo <= n1605_li;
    n1608_lo <= n1608_li;
    n1611_lo <= n1611_li;
    n1614_lo <= n1614_li;
    n1617_lo <= n1617_li;
    n1620_lo <= n1620_li;
    n1623_lo <= n1623_li;
    n1626_lo <= n1626_li;
    n1629_lo <= n1629_li;
    n1632_lo <= n1632_li;
    n1635_lo <= n1635_li;
    n1638_lo <= n1638_li;
    n1641_lo <= n1641_li;
    n1644_lo <= n1644_li;
    n1647_lo <= n1647_li;
    n1650_lo <= n1650_li;
    n1653_lo <= n1653_li;
    n1656_lo <= n1656_li;
    n1659_lo <= n1659_li;
    n1662_lo <= n1662_li;
    n1665_lo <= n1665_li;
    n1668_lo <= n1668_li;
    n1671_lo <= n1671_li;
    n1674_lo <= n1674_li;
    n1677_lo <= n1677_li;
    n1680_lo <= n1680_li;
    n1683_lo <= n1683_li;
    n1686_lo <= n1686_li;
    n1689_lo <= n1689_li;
    n1692_lo <= n1692_li;
    n1695_lo <= n1695_li;
    n1698_lo <= n1698_li;
    n1701_lo <= n1701_li;
    n1704_lo <= n1704_li;
    n1707_lo <= n1707_li;
    n1710_lo <= n1710_li;
    n1713_lo <= n1713_li;
    n1716_lo <= n1716_li;
    n1719_lo <= n1719_li;
    n1722_lo <= n1722_li;
    n1725_lo <= n1725_li;
    n1728_lo <= n1728_li;
    n1731_lo <= n1731_li;
    n1734_lo <= n1734_li;
    n1737_lo <= n1737_li;
    n1740_lo <= n1740_li;
    n1743_lo <= n1743_li;
    n1746_lo <= n1746_li;
    n1749_lo <= n1749_li;
    n1752_lo <= n1752_li;
    n1755_lo <= n1755_li;
    n1758_lo <= n1758_li;
    n1761_lo <= n1761_li;
    n1764_lo <= n1764_li;
    n1767_lo <= n1767_li;
    n1770_lo <= n1770_li;
    n1773_lo <= n1773_li;
    n1776_lo <= n1776_li;
    n1779_lo <= n1779_li;
    n1782_lo <= n1782_li;
    n1785_lo <= n1785_li;
    n1788_lo <= n1788_li;
    n1791_lo <= n1791_li;
    n1794_lo <= n1794_li;
    n1797_lo <= n1797_li;
    n1800_lo <= n1800_li;
    n1803_lo <= n1803_li;
    n1806_lo <= n1806_li;
    n1809_lo <= n1809_li;
    n1812_lo <= n1812_li;
    n1815_lo <= n1815_li;
    n1818_lo <= n1818_li;
    n1821_lo <= n1821_li;
    n1824_lo <= n1824_li;
    n1827_lo <= n1827_li;
    n1830_lo <= n1830_li;
    n1833_lo <= n1833_li;
    n1836_lo <= n1836_li;
    n1839_lo <= n1839_li;
    n1842_lo <= n1842_li;
    n1845_lo <= n1845_li;
    n1848_lo <= n1848_li;
    n1851_lo <= n1851_li;
    n1854_lo <= n1854_li;
    n1857_lo <= n1857_li;
    n1860_lo <= n1860_li;
    n1863_lo <= n1863_li;
    n1866_lo <= n1866_li;
    n1869_lo <= n1869_li;
    n1872_lo <= n1872_li;
    n1875_lo <= n1875_li;
    n1878_lo <= n1878_li;
    n1881_lo <= n1881_li;
    n1884_lo <= n1884_li;
    n1887_lo <= n1887_li;
    n1890_lo <= n1890_li;
    n1893_lo <= n1893_li;
    n1896_lo <= n1896_li;
    n1899_lo <= n1899_li;
    n1902_lo <= n1902_li;
    n1905_lo <= n1905_li;
    n1908_lo <= n1908_li;
    n1911_lo <= n1911_li;
    n1914_lo <= n1914_li;
    n1917_lo <= n1917_li;
    n1920_lo <= n1920_li;
    n1923_lo <= n1923_li;
    n1926_lo <= n1926_li;
    n1929_lo <= n1929_li;
    n1932_lo <= n1932_li;
    n1935_lo <= n1935_li;
    n1938_lo <= n1938_li;
    n1941_lo <= n1941_li;
    n1944_lo <= n1944_li;
    n1947_lo <= n1947_li;
    n1950_lo <= n1950_li;
    n1953_lo <= n1953_li;
    n1956_lo <= n1956_li;
    n1959_lo <= n1959_li;
    n1962_lo <= n1962_li;
    n1965_lo <= n1965_li;
    n1968_lo <= n1968_li;
    n1971_lo <= n1971_li;
    n1974_lo <= n1974_li;
    n1977_lo <= n1977_li;
    n1980_lo <= n1980_li;
    n1983_lo <= n1983_li;
    n1986_lo <= n1986_li;
    n1989_lo <= n1989_li;
    n1992_lo <= n1992_li;
    n1995_lo <= n1995_li;
    n1998_lo <= n1998_li;
    n2001_lo <= n2001_li;
    n2004_lo <= n2004_li;
    n2007_lo <= n2007_li;
    n2010_lo <= n2010_li;
    n2013_lo <= n2013_li;
    n2016_lo <= n2016_li;
    n2019_lo <= n2019_li;
    n2022_lo <= n2022_li;
    n2025_lo <= n2025_li;
    n2028_lo <= n2028_li;
    n2031_lo <= n2031_li;
    n2034_lo <= n2034_li;
    n2037_lo <= n2037_li;
    n2040_lo <= n2040_li;
    n2043_lo <= n2043_li;
    n2046_lo <= n2046_li;
    n2049_lo <= n2049_li;
    n2052_lo <= n2052_li;
    n2055_lo <= n2055_li;
    n2058_lo <= n2058_li;
    n2061_lo <= n2061_li;
    n2064_lo <= n2064_li;
    n2067_lo <= n2067_li;
    n2070_lo <= n2070_li;
    n2073_lo <= n2073_li;
    n2076_lo <= n2076_li;
    n2079_lo <= n2079_li;
    n2082_lo <= n2082_li;
    n2085_lo <= n2085_li;
    n2088_lo <= n2088_li;
    n2091_lo <= n2091_li;
    n2094_lo <= n2094_li;
    n2097_lo <= n2097_li;
    n2100_lo <= n2100_li;
    n2103_lo <= n2103_li;
    n2106_lo <= n2106_li;
    n2109_lo <= n2109_li;
    n2112_lo <= n2112_li;
    n2115_lo <= n2115_li;
    n2118_lo <= n2118_li;
    n2121_lo <= n2121_li;
    n2124_lo <= n2124_li;
    n2127_lo <= n2127_li;
    n2130_lo <= n2130_li;
    n2133_lo <= n2133_li;
    n2136_lo <= n2136_li;
    n2139_lo <= n2139_li;
    n2142_lo <= n2142_li;
    n2145_lo <= n2145_li;
    n2148_lo <= n2148_li;
    n2151_lo <= n2151_li;
    n2154_lo <= n2154_li;
    n2157_lo <= n2157_li;
    n2160_lo <= n2160_li;
    n2163_lo <= n2163_li;
    n2166_lo <= n2166_li;
    n2169_lo <= n2169_li;
    n2172_lo <= n2172_li;
    n2175_lo <= n2175_li;
    n2178_lo <= n2178_li;
    n2181_lo <= n2181_li;
    n2184_lo <= n2184_li;
    n2187_lo <= n2187_li;
    n2190_lo <= n2190_li;
    n2193_lo <= n2193_li;
    n2196_lo <= n2196_li;
    n2199_lo <= n2199_li;
    n2202_lo <= n2202_li;
    n2205_lo <= n2205_li;
    n2208_lo <= n2208_li;
    n2211_lo <= n2211_li;
    n2214_lo <= n2214_li;
    n2217_lo <= n2217_li;
    n2220_lo <= n2220_li;
    n2223_lo <= n2223_li;
    n2226_lo <= n2226_li;
    n2229_lo <= n2229_li;
    n2232_lo <= n2232_li;
    n2235_lo <= n2235_li;
    n2238_lo <= n2238_li;
    n2241_lo <= n2241_li;
    n2244_lo <= n2244_li;
    n2247_lo <= n2247_li;
    n2250_lo <= n2250_li;
    n2253_lo <= n2253_li;
    n2256_lo <= n2256_li;
    n2259_lo <= n2259_li;
    n2262_lo <= n2262_li;
    n2265_lo <= n2265_li;
    n2268_lo <= n2268_li;
    n2271_lo <= n2271_li;
    n2274_lo <= n2274_li;
    n2277_lo <= n2277_li;
    n2280_lo <= n2280_li;
    n2283_lo <= n2283_li;
    n2286_lo <= n2286_li;
    n2289_lo <= n2289_li;
    n2292_lo <= n2292_li;
    n2295_lo <= n2295_li;
    n2298_lo <= n2298_li;
    n2301_lo <= n2301_li;
    n2304_lo <= n2304_li;
    n2307_lo <= n2307_li;
    n2310_lo <= n2310_li;
    n2313_lo <= n2313_li;
    n2316_lo <= n2316_li;
    n2319_lo <= n2319_li;
    n2322_lo <= n2322_li;
    n2325_lo <= n2325_li;
    n2328_lo <= n2328_li;
    n2331_lo <= n2331_li;
    n2334_lo <= n2334_li;
    n2337_lo <= n2337_li;
    n2340_lo <= n2340_li;
    n2343_lo <= n2343_li;
    n2346_lo <= n2346_li;
    n2349_lo <= n2349_li;
    n2352_lo <= n2352_li;
    n2355_lo <= n2355_li;
    n2358_lo <= n2358_li;
    n2361_lo <= n2361_li;
    n2364_lo <= n2364_li;
    n2367_lo <= n2367_li;
    n2370_lo <= n2370_li;
    n2373_lo <= n2373_li;
    n2376_lo <= n2376_li;
    n2379_lo <= n2379_li;
    n2382_lo <= n2382_li;
    n2385_lo <= n2385_li;
    n2388_lo <= n2388_li;
    n2391_lo <= n2391_li;
    n2394_lo <= n2394_li;
    n2397_lo <= n2397_li;
    n2400_lo <= n2400_li;
    n2403_lo <= n2403_li;
    n2406_lo <= n2406_li;
    n2409_lo <= n2409_li;
    n2412_lo <= n2412_li;
    n2415_lo <= n2415_li;
    n2418_lo <= n2418_li;
    n2421_lo <= n2421_li;
    n2424_lo <= n2424_li;
    n2427_lo <= n2427_li;
    n2430_lo <= n2430_li;
    n2433_lo <= n2433_li;
    n2436_lo <= n2436_li;
    n2439_lo <= n2439_li;
    n2442_lo <= n2442_li;
    n2445_lo <= n2445_li;
    n2448_lo <= n2448_li;
    n2451_lo <= n2451_li;
    n2454_lo <= n2454_li;
    n2457_lo <= n2457_li;
    n2460_lo <= n2460_li;
    n2463_lo <= n2463_li;
    n2466_lo <= n2466_li;
    n2469_lo <= n2469_li;
    n2472_lo <= n2472_li;
    n2475_lo <= n2475_li;
    n2478_lo <= n2478_li;
    n2481_lo <= n2481_li;
    n2484_lo <= n2484_li;
    n2487_lo <= n2487_li;
    n2490_lo <= n2490_li;
    n2493_lo <= n2493_li;
    n2496_lo <= n2496_li;
    n2499_lo <= n2499_li;
    n2502_lo <= n2502_li;
    n2505_lo <= n2505_li;
    n2508_lo <= n2508_li;
    n2511_lo <= n2511_li;
    n2514_lo <= n2514_li;
    n2517_lo <= n2517_li;
    n2520_lo <= n2520_li;
    n2523_lo <= n2523_li;
    n2526_lo <= n2526_li;
    n2529_lo <= n2529_li;
    n2532_lo <= n2532_li;
    n2535_lo <= n2535_li;
    n2538_lo <= n2538_li;
    n2541_lo <= n2541_li;
    n2544_lo <= n2544_li;
    n2547_lo <= n2547_li;
    n2550_lo <= n2550_li;
    n2553_lo <= n2553_li;
    n2556_lo <= n2556_li;
    n2559_lo <= n2559_li;
    n2562_lo <= n2562_li;
    n2565_lo <= n2565_li;
    n2568_lo <= n2568_li;
    n2571_lo <= n2571_li;
    n2574_lo <= n2574_li;
    n2577_lo <= n2577_li;
    n2580_lo <= n2580_li;
    n2583_lo <= n2583_li;
    n2586_lo <= n2586_li;
    n2589_lo <= n2589_li;
    n2592_lo <= n2592_li;
    n2595_lo <= n2595_li;
    n2598_lo <= n2598_li;
    n2601_lo <= n2601_li;
    n2604_lo <= n2604_li;
    n2607_lo <= n2607_li;
    n2610_lo <= n2610_li;
    n2613_lo <= n2613_li;
    n2616_lo <= n2616_li;
    n2619_lo <= n2619_li;
    n2622_lo <= n2622_li;
    n2625_lo <= n2625_li;
    n2628_lo <= n2628_li;
    n2631_lo <= n2631_li;
    n2634_lo <= n2634_li;
    n2637_lo <= n2637_li;
    n2640_lo <= n2640_li;
    n2643_lo <= n2643_li;
    n2646_lo <= n2646_li;
    n2649_lo <= n2649_li;
    n2652_lo <= n2652_li;
    n2655_lo <= n2655_li;
    n2658_lo <= n2658_li;
    n2661_lo <= n2661_li;
    n2664_lo <= n2664_li;
    n2667_lo <= n2667_li;
    n2670_lo <= n2670_li;
    n2673_lo <= n2673_li;
    n2676_lo <= n2676_li;
    n2679_lo <= n2679_li;
    n2682_lo <= n2682_li;
    n2685_lo <= n2685_li;
    n2688_lo <= n2688_li;
    n2691_lo <= n2691_li;
    n2694_lo <= n2694_li;
    n2697_lo <= n2697_li;
    n2700_lo <= n2700_li;
    n2703_lo <= n2703_li;
    n2706_lo <= n2706_li;
    n2709_lo <= n2709_li;
    n2712_lo <= n2712_li;
    n2715_lo <= n2715_li;
    n2718_lo <= n2718_li;
    n2721_lo <= n2721_li;
    n2724_lo <= n2724_li;
    n2727_lo <= n2727_li;
    n2730_lo <= n2730_li;
    n2733_lo <= n2733_li;
    n2736_lo <= n2736_li;
    n2739_lo <= n2739_li;
    n2742_lo <= n2742_li;
    n2745_lo <= n2745_li;
    n2748_lo <= n2748_li;
    n2751_lo <= n2751_li;
    n2754_lo <= n2754_li;
    n2757_lo <= n2757_li;
    n2760_lo <= n2760_li;
    n2763_lo <= n2763_li;
    n2766_lo <= n2766_li;
    n2769_lo <= n2769_li;
    n2772_lo <= n2772_li;
    n2775_lo <= n2775_li;
    n2778_lo <= n2778_li;
    n2781_lo <= n2781_li;
    n2784_lo <= n2784_li;
    n2787_lo <= n2787_li;
    n2790_lo <= n2790_li;
    n2793_lo <= n2793_li;
    n2796_lo <= n2796_li;
    n2799_lo <= n2799_li;
    n2802_lo <= n2802_li;
    n2805_lo <= n2805_li;
    n2808_lo <= n2808_li;
    n2811_lo <= n2811_li;
    n2814_lo <= n2814_li;
    n2817_lo <= n2817_li;
    n2820_lo <= n2820_li;
    n2823_lo <= n2823_li;
    n2826_lo <= n2826_li;
    n2829_lo <= n2829_li;
    n2832_lo <= n2832_li;
    n2835_lo <= n2835_li;
    n2838_lo <= n2838_li;
    n2841_lo <= n2841_li;
    n2844_lo <= n2844_li;
    n2847_lo <= n2847_li;
    n2850_lo <= n2850_li;
    n2853_lo <= n2853_li;
    n2856_lo <= n2856_li;
    n2859_lo <= n2859_li;
    n2862_lo <= n2862_li;
    n2865_lo <= n2865_li;
    n2868_lo <= n2868_li;
    n2871_lo <= n2871_li;
    n2874_lo <= n2874_li;
    n2877_lo <= n2877_li;
    n2880_lo <= n2880_li;
    n2883_lo <= n2883_li;
    n2886_lo <= n2886_li;
    n2889_lo <= n2889_li;
    n2892_lo <= n2892_li;
    n2895_lo <= n2895_li;
    n2898_lo <= n2898_li;
    n2901_lo <= n2901_li;
    n2904_lo <= n2904_li;
    n2907_lo <= n2907_li;
    n2910_lo <= n2910_li;
    n2913_lo <= n2913_li;
    n2916_lo <= n2916_li;
    n2919_lo <= n2919_li;
    n2922_lo <= n2922_li;
    n2925_lo <= n2925_li;
    n2928_lo <= n2928_li;
    n2931_lo <= n2931_li;
    n2934_lo <= n2934_li;
    n2937_lo <= n2937_li;
    n2940_lo <= n2940_li;
    n2943_lo <= n2943_li;
    n2946_lo <= n2946_li;
    n2949_lo <= n2949_li;
    n2952_lo <= n2952_li;
    n2955_lo <= n2955_li;
    n2958_lo <= n2958_li;
    n2961_lo <= n2961_li;
    n2964_lo <= n2964_li;
    n2967_lo <= n2967_li;
    n2970_lo <= n2970_li;
    n2973_lo <= n2973_li;
    n2976_lo <= n2976_li;
    n2979_lo <= n2979_li;
    n2982_lo <= n2982_li;
    n2985_lo <= n2985_li;
    n2988_lo <= n2988_li;
    n2991_lo <= n2991_li;
    n2994_lo <= n2994_li;
    n2997_lo <= n2997_li;
    n3000_lo <= n3000_li;
    n3003_lo <= n3003_li;
    n3006_lo <= n3006_li;
    n3009_lo <= n3009_li;
    n3012_lo <= n3012_li;
    n3015_lo <= n3015_li;
    n3018_lo <= n3018_li;
    n3021_lo <= n3021_li;
    n3024_lo <= n3024_li;
    n3027_lo <= n3027_li;
    n3030_lo <= n3030_li;
    n3033_lo <= n3033_li;
    n3036_lo <= n3036_li;
    n3039_lo <= n3039_li;
    n3042_lo <= n3042_li;
    n3045_lo <= n3045_li;
    n3048_lo <= n3048_li;
    n3051_lo <= n3051_li;
    n3054_lo <= n3054_li;
    n3057_lo <= n3057_li;
    n3060_lo <= n3060_li;
    n3063_lo <= n3063_li;
    n3066_lo <= n3066_li;
    n3069_lo <= n3069_li;
    n3072_lo <= n3072_li;
    n3075_lo <= n3075_li;
    n3078_lo <= n3078_li;
    n3081_lo <= n3081_li;
    n3084_lo <= n3084_li;
    n3087_lo <= n3087_li;
    n3090_lo <= n3090_li;
    n3093_lo <= n3093_li;
    n3096_lo <= n3096_li;
    n3099_lo <= n3099_li;
    n3102_lo <= n3102_li;
    n3105_lo <= n3105_li;
    n3108_lo <= n3108_li;
    n3111_lo <= n3111_li;
    n3114_lo <= n3114_li;
    n3117_lo <= n3117_li;
    n3120_lo <= n3120_li;
    n3123_lo <= n3123_li;
    n3126_lo <= n3126_li;
    n3129_lo <= n3129_li;
    n3132_lo <= n3132_li;
    n3135_lo <= n3135_li;
    n3138_lo <= n3138_li;
    n3141_lo <= n3141_li;
    n3144_lo <= n3144_li;
    n3147_lo <= n3147_li;
    n3150_lo <= n3150_li;
    n3153_lo <= n3153_li;
    n3156_lo <= n3156_li;
    n3159_lo <= n3159_li;
    n3162_lo <= n3162_li;
    n3165_lo <= n3165_li;
    n3168_lo <= n3168_li;
    n3171_lo <= n3171_li;
    n3174_lo <= n3174_li;
    n3177_lo <= n3177_li;
    n3180_lo <= n3180_li;
    n3183_lo <= n3183_li;
    n3186_lo <= n3186_li;
    n3189_lo <= n3189_li;
    n3192_lo <= n3192_li;
    n3195_lo <= n3195_li;
    n3198_lo <= n3198_li;
    n3201_lo <= n3201_li;
    n3204_lo <= n3204_li;
    n3207_lo <= n3207_li;
    n3210_lo <= n3210_li;
    n3213_lo <= n3213_li;
    n3216_lo <= n3216_li;
    n3219_lo <= n3219_li;
    n3222_lo <= n3222_li;
    n3225_lo <= n3225_li;
    n3228_lo <= n3228_li;
    n3231_lo <= n3231_li;
    n3234_lo <= n3234_li;
    n3237_lo <= n3237_li;
    n3240_lo <= n3240_li;
    n3243_lo <= n3243_li;
    n3246_lo <= n3246_li;
    n3249_lo <= n3249_li;
    n3252_lo <= n3252_li;
    n3255_lo <= n3255_li;
    n3258_lo <= n3258_li;
    n3261_lo <= n3261_li;
    n3264_lo <= n3264_li;
    n3267_lo <= n3267_li;
    n3270_lo <= n3270_li;
    n3273_lo <= n3273_li;
    n3276_lo <= n3276_li;
    n3279_lo <= n3279_li;
    n3282_lo <= n3282_li;
    n3285_lo <= n3285_li;
    n3288_lo <= n3288_li;
    n3291_lo <= n3291_li;
    n3294_lo <= n3294_li;
    n3297_lo <= n3297_li;
  end
  initial begin
    n1416_lo <= 1'b0;
    n1419_lo <= 1'b0;
    n1422_lo <= 1'b0;
    n1425_lo <= 1'b0;
    n1428_lo <= 1'b0;
    n1431_lo <= 1'b0;
    n1434_lo <= 1'b0;
    n1437_lo <= 1'b0;
    n1440_lo <= 1'b0;
    n1443_lo <= 1'b0;
    n1446_lo <= 1'b0;
    n1449_lo <= 1'b0;
    n1452_lo <= 1'b0;
    n1455_lo <= 1'b0;
    n1458_lo <= 1'b0;
    n1461_lo <= 1'b0;
    n1464_lo <= 1'b0;
    n1467_lo <= 1'b0;
    n1470_lo <= 1'b0;
    n1473_lo <= 1'b0;
    n1476_lo <= 1'b0;
    n1479_lo <= 1'b0;
    n1482_lo <= 1'b0;
    n1485_lo <= 1'b0;
    n1488_lo <= 1'b0;
    n1491_lo <= 1'b0;
    n1494_lo <= 1'b0;
    n1497_lo <= 1'b0;
    n1500_lo <= 1'b0;
    n1503_lo <= 1'b0;
    n1506_lo <= 1'b0;
    n1509_lo <= 1'b0;
    n1512_lo <= 1'b0;
    n1515_lo <= 1'b0;
    n1518_lo <= 1'b0;
    n1521_lo <= 1'b0;
    n1524_lo <= 1'b0;
    n1527_lo <= 1'b0;
    n1530_lo <= 1'b0;
    n1533_lo <= 1'b0;
    n1536_lo <= 1'b0;
    n1539_lo <= 1'b0;
    n1542_lo <= 1'b0;
    n1545_lo <= 1'b0;
    n1548_lo <= 1'b0;
    n1551_lo <= 1'b0;
    n1554_lo <= 1'b0;
    n1557_lo <= 1'b0;
    n1560_lo <= 1'b0;
    n1563_lo <= 1'b0;
    n1566_lo <= 1'b0;
    n1569_lo <= 1'b0;
    n1572_lo <= 1'b0;
    n1575_lo <= 1'b0;
    n1578_lo <= 1'b0;
    n1581_lo <= 1'b0;
    n1584_lo <= 1'b0;
    n1587_lo <= 1'b0;
    n1590_lo <= 1'b0;
    n1593_lo <= 1'b0;
    n1596_lo <= 1'b0;
    n1599_lo <= 1'b0;
    n1602_lo <= 1'b0;
    n1605_lo <= 1'b0;
    n1608_lo <= 1'b0;
    n1611_lo <= 1'b0;
    n1614_lo <= 1'b0;
    n1617_lo <= 1'b0;
    n1620_lo <= 1'b0;
    n1623_lo <= 1'b0;
    n1626_lo <= 1'b0;
    n1629_lo <= 1'b0;
    n1632_lo <= 1'b0;
    n1635_lo <= 1'b0;
    n1638_lo <= 1'b0;
    n1641_lo <= 1'b0;
    n1644_lo <= 1'b0;
    n1647_lo <= 1'b0;
    n1650_lo <= 1'b0;
    n1653_lo <= 1'b0;
    n1656_lo <= 1'b0;
    n1659_lo <= 1'b0;
    n1662_lo <= 1'b0;
    n1665_lo <= 1'b0;
    n1668_lo <= 1'b0;
    n1671_lo <= 1'b0;
    n1674_lo <= 1'b0;
    n1677_lo <= 1'b0;
    n1680_lo <= 1'b0;
    n1683_lo <= 1'b0;
    n1686_lo <= 1'b0;
    n1689_lo <= 1'b0;
    n1692_lo <= 1'b0;
    n1695_lo <= 1'b0;
    n1698_lo <= 1'b0;
    n1701_lo <= 1'b0;
    n1704_lo <= 1'b0;
    n1707_lo <= 1'b0;
    n1710_lo <= 1'b0;
    n1713_lo <= 1'b0;
    n1716_lo <= 1'b0;
    n1719_lo <= 1'b0;
    n1722_lo <= 1'b0;
    n1725_lo <= 1'b0;
    n1728_lo <= 1'b0;
    n1731_lo <= 1'b0;
    n1734_lo <= 1'b0;
    n1737_lo <= 1'b0;
    n1740_lo <= 1'b0;
    n1743_lo <= 1'b0;
    n1746_lo <= 1'b0;
    n1749_lo <= 1'b0;
    n1752_lo <= 1'b0;
    n1755_lo <= 1'b0;
    n1758_lo <= 1'b0;
    n1761_lo <= 1'b0;
    n1764_lo <= 1'b0;
    n1767_lo <= 1'b0;
    n1770_lo <= 1'b0;
    n1773_lo <= 1'b0;
    n1776_lo <= 1'b0;
    n1779_lo <= 1'b0;
    n1782_lo <= 1'b0;
    n1785_lo <= 1'b0;
    n1788_lo <= 1'b0;
    n1791_lo <= 1'b0;
    n1794_lo <= 1'b0;
    n1797_lo <= 1'b0;
    n1800_lo <= 1'b0;
    n1803_lo <= 1'b0;
    n1806_lo <= 1'b0;
    n1809_lo <= 1'b0;
    n1812_lo <= 1'b0;
    n1815_lo <= 1'b0;
    n1818_lo <= 1'b0;
    n1821_lo <= 1'b0;
    n1824_lo <= 1'b0;
    n1827_lo <= 1'b0;
    n1830_lo <= 1'b0;
    n1833_lo <= 1'b0;
    n1836_lo <= 1'b0;
    n1839_lo <= 1'b0;
    n1842_lo <= 1'b0;
    n1845_lo <= 1'b0;
    n1848_lo <= 1'b0;
    n1851_lo <= 1'b0;
    n1854_lo <= 1'b0;
    n1857_lo <= 1'b0;
    n1860_lo <= 1'b0;
    n1863_lo <= 1'b0;
    n1866_lo <= 1'b0;
    n1869_lo <= 1'b0;
    n1872_lo <= 1'b0;
    n1875_lo <= 1'b0;
    n1878_lo <= 1'b0;
    n1881_lo <= 1'b0;
    n1884_lo <= 1'b0;
    n1887_lo <= 1'b0;
    n1890_lo <= 1'b0;
    n1893_lo <= 1'b0;
    n1896_lo <= 1'b0;
    n1899_lo <= 1'b0;
    n1902_lo <= 1'b0;
    n1905_lo <= 1'b0;
    n1908_lo <= 1'b0;
    n1911_lo <= 1'b0;
    n1914_lo <= 1'b0;
    n1917_lo <= 1'b0;
    n1920_lo <= 1'b0;
    n1923_lo <= 1'b0;
    n1926_lo <= 1'b0;
    n1929_lo <= 1'b0;
    n1932_lo <= 1'b0;
    n1935_lo <= 1'b0;
    n1938_lo <= 1'b0;
    n1941_lo <= 1'b0;
    n1944_lo <= 1'b0;
    n1947_lo <= 1'b0;
    n1950_lo <= 1'b0;
    n1953_lo <= 1'b0;
    n1956_lo <= 1'b0;
    n1959_lo <= 1'b0;
    n1962_lo <= 1'b0;
    n1965_lo <= 1'b0;
    n1968_lo <= 1'b0;
    n1971_lo <= 1'b0;
    n1974_lo <= 1'b0;
    n1977_lo <= 1'b0;
    n1980_lo <= 1'b0;
    n1983_lo <= 1'b0;
    n1986_lo <= 1'b0;
    n1989_lo <= 1'b0;
    n1992_lo <= 1'b0;
    n1995_lo <= 1'b0;
    n1998_lo <= 1'b0;
    n2001_lo <= 1'b0;
    n2004_lo <= 1'b0;
    n2007_lo <= 1'b0;
    n2010_lo <= 1'b0;
    n2013_lo <= 1'b0;
    n2016_lo <= 1'b0;
    n2019_lo <= 1'b0;
    n2022_lo <= 1'b0;
    n2025_lo <= 1'b0;
    n2028_lo <= 1'b0;
    n2031_lo <= 1'b0;
    n2034_lo <= 1'b0;
    n2037_lo <= 1'b0;
    n2040_lo <= 1'b0;
    n2043_lo <= 1'b0;
    n2046_lo <= 1'b0;
    n2049_lo <= 1'b0;
    n2052_lo <= 1'b0;
    n2055_lo <= 1'b0;
    n2058_lo <= 1'b0;
    n2061_lo <= 1'b0;
    n2064_lo <= 1'b0;
    n2067_lo <= 1'b0;
    n2070_lo <= 1'b0;
    n2073_lo <= 1'b0;
    n2076_lo <= 1'b0;
    n2079_lo <= 1'b0;
    n2082_lo <= 1'b0;
    n2085_lo <= 1'b0;
    n2088_lo <= 1'b0;
    n2091_lo <= 1'b0;
    n2094_lo <= 1'b0;
    n2097_lo <= 1'b0;
    n2100_lo <= 1'b0;
    n2103_lo <= 1'b0;
    n2106_lo <= 1'b0;
    n2109_lo <= 1'b0;
    n2112_lo <= 1'b0;
    n2115_lo <= 1'b0;
    n2118_lo <= 1'b0;
    n2121_lo <= 1'b0;
    n2124_lo <= 1'b0;
    n2127_lo <= 1'b0;
    n2130_lo <= 1'b0;
    n2133_lo <= 1'b0;
    n2136_lo <= 1'b0;
    n2139_lo <= 1'b0;
    n2142_lo <= 1'b0;
    n2145_lo <= 1'b0;
    n2148_lo <= 1'b0;
    n2151_lo <= 1'b0;
    n2154_lo <= 1'b0;
    n2157_lo <= 1'b0;
    n2160_lo <= 1'b0;
    n2163_lo <= 1'b0;
    n2166_lo <= 1'b0;
    n2169_lo <= 1'b0;
    n2172_lo <= 1'b0;
    n2175_lo <= 1'b0;
    n2178_lo <= 1'b0;
    n2181_lo <= 1'b0;
    n2184_lo <= 1'b0;
    n2187_lo <= 1'b0;
    n2190_lo <= 1'b0;
    n2193_lo <= 1'b0;
    n2196_lo <= 1'b0;
    n2199_lo <= 1'b0;
    n2202_lo <= 1'b0;
    n2205_lo <= 1'b0;
    n2208_lo <= 1'b0;
    n2211_lo <= 1'b0;
    n2214_lo <= 1'b0;
    n2217_lo <= 1'b0;
    n2220_lo <= 1'b0;
    n2223_lo <= 1'b0;
    n2226_lo <= 1'b0;
    n2229_lo <= 1'b0;
    n2232_lo <= 1'b0;
    n2235_lo <= 1'b0;
    n2238_lo <= 1'b0;
    n2241_lo <= 1'b0;
    n2244_lo <= 1'b0;
    n2247_lo <= 1'b0;
    n2250_lo <= 1'b0;
    n2253_lo <= 1'b0;
    n2256_lo <= 1'b0;
    n2259_lo <= 1'b0;
    n2262_lo <= 1'b0;
    n2265_lo <= 1'b0;
    n2268_lo <= 1'b0;
    n2271_lo <= 1'b0;
    n2274_lo <= 1'b0;
    n2277_lo <= 1'b0;
    n2280_lo <= 1'b0;
    n2283_lo <= 1'b0;
    n2286_lo <= 1'b0;
    n2289_lo <= 1'b0;
    n2292_lo <= 1'b0;
    n2295_lo <= 1'b0;
    n2298_lo <= 1'b0;
    n2301_lo <= 1'b0;
    n2304_lo <= 1'b0;
    n2307_lo <= 1'b0;
    n2310_lo <= 1'b0;
    n2313_lo <= 1'b0;
    n2316_lo <= 1'b0;
    n2319_lo <= 1'b0;
    n2322_lo <= 1'b0;
    n2325_lo <= 1'b0;
    n2328_lo <= 1'b0;
    n2331_lo <= 1'b0;
    n2334_lo <= 1'b0;
    n2337_lo <= 1'b0;
    n2340_lo <= 1'b0;
    n2343_lo <= 1'b0;
    n2346_lo <= 1'b0;
    n2349_lo <= 1'b0;
    n2352_lo <= 1'b0;
    n2355_lo <= 1'b0;
    n2358_lo <= 1'b0;
    n2361_lo <= 1'b0;
    n2364_lo <= 1'b0;
    n2367_lo <= 1'b0;
    n2370_lo <= 1'b0;
    n2373_lo <= 1'b0;
    n2376_lo <= 1'b0;
    n2379_lo <= 1'b0;
    n2382_lo <= 1'b0;
    n2385_lo <= 1'b0;
    n2388_lo <= 1'b0;
    n2391_lo <= 1'b0;
    n2394_lo <= 1'b0;
    n2397_lo <= 1'b0;
    n2400_lo <= 1'b0;
    n2403_lo <= 1'b0;
    n2406_lo <= 1'b0;
    n2409_lo <= 1'b0;
    n2412_lo <= 1'b0;
    n2415_lo <= 1'b0;
    n2418_lo <= 1'b0;
    n2421_lo <= 1'b0;
    n2424_lo <= 1'b0;
    n2427_lo <= 1'b0;
    n2430_lo <= 1'b0;
    n2433_lo <= 1'b0;
    n2436_lo <= 1'b0;
    n2439_lo <= 1'b0;
    n2442_lo <= 1'b0;
    n2445_lo <= 1'b0;
    n2448_lo <= 1'b0;
    n2451_lo <= 1'b0;
    n2454_lo <= 1'b0;
    n2457_lo <= 1'b0;
    n2460_lo <= 1'b0;
    n2463_lo <= 1'b0;
    n2466_lo <= 1'b0;
    n2469_lo <= 1'b0;
    n2472_lo <= 1'b0;
    n2475_lo <= 1'b0;
    n2478_lo <= 1'b0;
    n2481_lo <= 1'b0;
    n2484_lo <= 1'b0;
    n2487_lo <= 1'b0;
    n2490_lo <= 1'b0;
    n2493_lo <= 1'b0;
    n2496_lo <= 1'b0;
    n2499_lo <= 1'b0;
    n2502_lo <= 1'b0;
    n2505_lo <= 1'b0;
    n2508_lo <= 1'b0;
    n2511_lo <= 1'b0;
    n2514_lo <= 1'b0;
    n2517_lo <= 1'b0;
    n2520_lo <= 1'b0;
    n2523_lo <= 1'b0;
    n2526_lo <= 1'b0;
    n2529_lo <= 1'b0;
    n2532_lo <= 1'b0;
    n2535_lo <= 1'b0;
    n2538_lo <= 1'b0;
    n2541_lo <= 1'b0;
    n2544_lo <= 1'b0;
    n2547_lo <= 1'b0;
    n2550_lo <= 1'b0;
    n2553_lo <= 1'b0;
    n2556_lo <= 1'b0;
    n2559_lo <= 1'b0;
    n2562_lo <= 1'b0;
    n2565_lo <= 1'b0;
    n2568_lo <= 1'b0;
    n2571_lo <= 1'b0;
    n2574_lo <= 1'b0;
    n2577_lo <= 1'b0;
    n2580_lo <= 1'b0;
    n2583_lo <= 1'b0;
    n2586_lo <= 1'b0;
    n2589_lo <= 1'b0;
    n2592_lo <= 1'b0;
    n2595_lo <= 1'b0;
    n2598_lo <= 1'b0;
    n2601_lo <= 1'b0;
    n2604_lo <= 1'b0;
    n2607_lo <= 1'b0;
    n2610_lo <= 1'b0;
    n2613_lo <= 1'b0;
    n2616_lo <= 1'b0;
    n2619_lo <= 1'b0;
    n2622_lo <= 1'b0;
    n2625_lo <= 1'b0;
    n2628_lo <= 1'b0;
    n2631_lo <= 1'b0;
    n2634_lo <= 1'b0;
    n2637_lo <= 1'b0;
    n2640_lo <= 1'b0;
    n2643_lo <= 1'b0;
    n2646_lo <= 1'b0;
    n2649_lo <= 1'b0;
    n2652_lo <= 1'b0;
    n2655_lo <= 1'b0;
    n2658_lo <= 1'b0;
    n2661_lo <= 1'b0;
    n2664_lo <= 1'b0;
    n2667_lo <= 1'b0;
    n2670_lo <= 1'b0;
    n2673_lo <= 1'b0;
    n2676_lo <= 1'b0;
    n2679_lo <= 1'b0;
    n2682_lo <= 1'b0;
    n2685_lo <= 1'b0;
    n2688_lo <= 1'b0;
    n2691_lo <= 1'b0;
    n2694_lo <= 1'b0;
    n2697_lo <= 1'b0;
    n2700_lo <= 1'b0;
    n2703_lo <= 1'b0;
    n2706_lo <= 1'b0;
    n2709_lo <= 1'b0;
    n2712_lo <= 1'b0;
    n2715_lo <= 1'b0;
    n2718_lo <= 1'b0;
    n2721_lo <= 1'b0;
    n2724_lo <= 1'b0;
    n2727_lo <= 1'b0;
    n2730_lo <= 1'b0;
    n2733_lo <= 1'b0;
    n2736_lo <= 1'b0;
    n2739_lo <= 1'b0;
    n2742_lo <= 1'b0;
    n2745_lo <= 1'b0;
    n2748_lo <= 1'b0;
    n2751_lo <= 1'b0;
    n2754_lo <= 1'b0;
    n2757_lo <= 1'b0;
    n2760_lo <= 1'b0;
    n2763_lo <= 1'b0;
    n2766_lo <= 1'b0;
    n2769_lo <= 1'b0;
    n2772_lo <= 1'b0;
    n2775_lo <= 1'b0;
    n2778_lo <= 1'b0;
    n2781_lo <= 1'b0;
    n2784_lo <= 1'b0;
    n2787_lo <= 1'b0;
    n2790_lo <= 1'b0;
    n2793_lo <= 1'b0;
    n2796_lo <= 1'b0;
    n2799_lo <= 1'b0;
    n2802_lo <= 1'b0;
    n2805_lo <= 1'b0;
    n2808_lo <= 1'b0;
    n2811_lo <= 1'b0;
    n2814_lo <= 1'b0;
    n2817_lo <= 1'b0;
    n2820_lo <= 1'b0;
    n2823_lo <= 1'b0;
    n2826_lo <= 1'b0;
    n2829_lo <= 1'b0;
    n2832_lo <= 1'b0;
    n2835_lo <= 1'b0;
    n2838_lo <= 1'b0;
    n2841_lo <= 1'b0;
    n2844_lo <= 1'b0;
    n2847_lo <= 1'b0;
    n2850_lo <= 1'b0;
    n2853_lo <= 1'b0;
    n2856_lo <= 1'b0;
    n2859_lo <= 1'b0;
    n2862_lo <= 1'b0;
    n2865_lo <= 1'b0;
    n2868_lo <= 1'b0;
    n2871_lo <= 1'b0;
    n2874_lo <= 1'b0;
    n2877_lo <= 1'b0;
    n2880_lo <= 1'b0;
    n2883_lo <= 1'b0;
    n2886_lo <= 1'b0;
    n2889_lo <= 1'b0;
    n2892_lo <= 1'b0;
    n2895_lo <= 1'b0;
    n2898_lo <= 1'b0;
    n2901_lo <= 1'b0;
    n2904_lo <= 1'b0;
    n2907_lo <= 1'b0;
    n2910_lo <= 1'b0;
    n2913_lo <= 1'b0;
    n2916_lo <= 1'b0;
    n2919_lo <= 1'b0;
    n2922_lo <= 1'b0;
    n2925_lo <= 1'b0;
    n2928_lo <= 1'b0;
    n2931_lo <= 1'b0;
    n2934_lo <= 1'b0;
    n2937_lo <= 1'b0;
    n2940_lo <= 1'b0;
    n2943_lo <= 1'b0;
    n2946_lo <= 1'b0;
    n2949_lo <= 1'b0;
    n2952_lo <= 1'b0;
    n2955_lo <= 1'b0;
    n2958_lo <= 1'b0;
    n2961_lo <= 1'b0;
    n2964_lo <= 1'b0;
    n2967_lo <= 1'b0;
    n2970_lo <= 1'b0;
    n2973_lo <= 1'b0;
    n2976_lo <= 1'b0;
    n2979_lo <= 1'b0;
    n2982_lo <= 1'b0;
    n2985_lo <= 1'b0;
    n2988_lo <= 1'b0;
    n2991_lo <= 1'b0;
    n2994_lo <= 1'b0;
    n2997_lo <= 1'b0;
    n3000_lo <= 1'b0;
    n3003_lo <= 1'b0;
    n3006_lo <= 1'b0;
    n3009_lo <= 1'b0;
    n3012_lo <= 1'b0;
    n3015_lo <= 1'b0;
    n3018_lo <= 1'b0;
    n3021_lo <= 1'b0;
    n3024_lo <= 1'b0;
    n3027_lo <= 1'b0;
    n3030_lo <= 1'b0;
    n3033_lo <= 1'b0;
    n3036_lo <= 1'b0;
    n3039_lo <= 1'b0;
    n3042_lo <= 1'b0;
    n3045_lo <= 1'b0;
    n3048_lo <= 1'b0;
    n3051_lo <= 1'b0;
    n3054_lo <= 1'b0;
    n3057_lo <= 1'b0;
    n3060_lo <= 1'b0;
    n3063_lo <= 1'b0;
    n3066_lo <= 1'b0;
    n3069_lo <= 1'b0;
    n3072_lo <= 1'b0;
    n3075_lo <= 1'b0;
    n3078_lo <= 1'b0;
    n3081_lo <= 1'b0;
    n3084_lo <= 1'b0;
    n3087_lo <= 1'b0;
    n3090_lo <= 1'b0;
    n3093_lo <= 1'b0;
    n3096_lo <= 1'b0;
    n3099_lo <= 1'b0;
    n3102_lo <= 1'b0;
    n3105_lo <= 1'b0;
    n3108_lo <= 1'b0;
    n3111_lo <= 1'b0;
    n3114_lo <= 1'b0;
    n3117_lo <= 1'b0;
    n3120_lo <= 1'b0;
    n3123_lo <= 1'b0;
    n3126_lo <= 1'b0;
    n3129_lo <= 1'b0;
    n3132_lo <= 1'b0;
    n3135_lo <= 1'b0;
    n3138_lo <= 1'b0;
    n3141_lo <= 1'b0;
    n3144_lo <= 1'b0;
    n3147_lo <= 1'b0;
    n3150_lo <= 1'b0;
    n3153_lo <= 1'b0;
    n3156_lo <= 1'b0;
    n3159_lo <= 1'b0;
    n3162_lo <= 1'b0;
    n3165_lo <= 1'b0;
    n3168_lo <= 1'b0;
    n3171_lo <= 1'b0;
    n3174_lo <= 1'b0;
    n3177_lo <= 1'b0;
    n3180_lo <= 1'b0;
    n3183_lo <= 1'b0;
    n3186_lo <= 1'b0;
    n3189_lo <= 1'b0;
    n3192_lo <= 1'b0;
    n3195_lo <= 1'b0;
    n3198_lo <= 1'b0;
    n3201_lo <= 1'b0;
    n3204_lo <= 1'b0;
    n3207_lo <= 1'b0;
    n3210_lo <= 1'b0;
    n3213_lo <= 1'b0;
    n3216_lo <= 1'b0;
    n3219_lo <= 1'b0;
    n3222_lo <= 1'b0;
    n3225_lo <= 1'b0;
    n3228_lo <= 1'b0;
    n3231_lo <= 1'b0;
    n3234_lo <= 1'b0;
    n3237_lo <= 1'b0;
    n3240_lo <= 1'b0;
    n3243_lo <= 1'b0;
    n3246_lo <= 1'b0;
    n3249_lo <= 1'b0;
    n3252_lo <= 1'b0;
    n3255_lo <= 1'b0;
    n3258_lo <= 1'b0;
    n3261_lo <= 1'b0;
    n3264_lo <= 1'b0;
    n3267_lo <= 1'b0;
    n3270_lo <= 1'b0;
    n3273_lo <= 1'b0;
    n3276_lo <= 1'b0;
    n3279_lo <= 1'b0;
    n3282_lo <= 1'b0;
    n3285_lo <= 1'b0;
    n3288_lo <= 1'b0;
    n3291_lo <= 1'b0;
    n3294_lo <= 1'b0;
    n3297_lo <= 1'b0;
  end
endmodule


