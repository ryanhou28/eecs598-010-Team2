
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G6257,
  G6258,
  G6259,
  G6260,
  G6261,
  G6262,
  G6263,
  G6264,
  G6265,
  G6266,
  G6267,
  G6268,
  G6269,
  G6270,
  G6271,
  G6272,
  G6273,
  G6274,
  G6275,
  G6276,
  G6277,
  G6278,
  G6279,
  G6280,
  G6281,
  G6282,
  G6283,
  G6284,
  G6285,
  G6286,
  G6287,
  G6288
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;
  output G6257;output G6258;output G6259;output G6260;output G6261;output G6262;output G6263;output G6264;output G6265;output G6266;output G6267;output G6268;output G6269;output G6270;output G6271;output G6272;output G6273;output G6274;output G6275;output G6276;output G6277;output G6278;output G6279;output G6280;output G6281;output G6282;output G6283;output G6284;output G6285;output G6286;output G6287;output G6288;
  wire new_n66_;wire new_n67_;wire new_n68_;wire new_n69_;wire new_n71_;wire new_n72_;wire new_n73_;wire new_n74_;wire new_n75_;wire new_n76_;wire new_n77_;wire new_n78_;wire new_n79_;wire new_n80_;wire new_n81_;wire new_n83_;wire new_n84_;wire new_n85_;wire new_n86_;wire new_n87_;wire new_n88_;wire new_n89_;wire new_n90_;wire new_n91_;wire new_n92_;wire new_n93_;wire new_n94_;wire new_n95_;wire new_n96_;wire new_n97_;wire new_n98_;wire new_n99_;wire new_n100_;wire new_n101_;wire new_n103_;wire new_n104_;wire new_n105_;wire new_n106_;wire new_n107_;wire new_n108_;wire new_n109_;wire new_n110_;wire new_n111_;wire new_n112_;wire new_n113_;wire new_n114_;wire new_n115_;wire new_n116_;wire new_n117_;wire new_n118_;wire new_n119_;wire new_n120_;wire new_n121_;wire new_n122_;wire new_n123_;wire new_n124_;wire new_n125_;wire new_n126_;wire new_n127_;wire new_n128_;wire new_n129_;wire new_n131_;wire new_n132_;wire new_n133_;wire new_n134_;wire new_n135_;wire new_n136_;wire new_n137_;wire new_n138_;wire new_n139_;wire new_n140_;wire new_n141_;wire new_n142_;wire new_n143_;wire new_n144_;wire new_n145_;wire new_n146_;wire new_n147_;wire new_n148_;wire new_n149_;wire new_n150_;wire new_n151_;wire new_n152_;wire new_n153_;wire new_n154_;wire new_n155_;wire new_n156_;wire new_n157_;wire new_n158_;wire new_n159_;wire new_n160_;wire new_n161_;wire new_n162_;wire new_n163_;wire new_n164_;wire new_n165_;wire new_n167_;wire new_n168_;wire new_n169_;wire new_n170_;wire new_n171_;wire new_n172_;wire new_n173_;wire new_n174_;wire new_n175_;wire new_n176_;wire new_n177_;wire new_n178_;wire new_n179_;wire new_n180_;wire new_n181_;wire new_n182_;wire new_n183_;wire new_n184_;wire new_n185_;wire new_n186_;wire new_n187_;wire new_n188_;wire new_n189_;wire new_n190_;wire new_n191_;wire new_n192_;wire new_n193_;wire new_n194_;wire new_n195_;wire new_n196_;wire new_n197_;wire new_n198_;wire new_n199_;wire new_n200_;wire new_n201_;wire new_n202_;wire new_n203_;wire new_n204_;wire new_n205_;wire new_n206_;wire new_n207_;wire new_n208_;wire new_n209_;wire new_n211_;wire new_n212_;wire new_n213_;wire new_n214_;wire new_n215_;wire new_n216_;wire new_n217_;wire new_n218_;wire new_n219_;wire new_n220_;wire new_n221_;wire new_n222_;wire new_n223_;wire new_n224_;wire new_n225_;wire new_n226_;wire new_n227_;wire new_n228_;wire new_n229_;wire new_n230_;wire new_n231_;wire new_n232_;wire new_n233_;wire new_n234_;wire new_n235_;wire new_n236_;wire new_n237_;wire new_n238_;wire new_n239_;wire new_n240_;wire new_n241_;wire new_n242_;wire new_n243_;wire new_n244_;wire new_n245_;wire new_n246_;wire new_n247_;wire new_n248_;wire new_n249_;wire new_n250_;wire new_n251_;wire new_n252_;wire new_n253_;wire new_n254_;wire new_n255_;wire new_n256_;wire new_n257_;wire new_n258_;wire new_n259_;wire new_n260_;wire new_n261_;wire new_n263_;wire new_n264_;wire new_n265_;wire new_n266_;wire new_n267_;wire new_n268_;wire new_n269_;wire new_n270_;wire new_n271_;wire new_n272_;wire new_n273_;wire new_n274_;wire new_n275_;wire new_n276_;wire new_n277_;wire new_n278_;wire new_n279_;wire new_n280_;wire new_n281_;wire new_n282_;wire new_n283_;wire new_n284_;wire new_n285_;wire new_n286_;wire new_n287_;wire new_n288_;wire new_n289_;wire new_n290_;wire new_n291_;wire new_n292_;wire new_n293_;wire new_n294_;wire new_n295_;wire new_n296_;wire new_n297_;wire new_n298_;wire new_n299_;wire new_n300_;wire new_n301_;wire new_n302_;wire new_n303_;wire new_n304_;wire new_n305_;wire new_n306_;wire new_n307_;wire new_n308_;wire new_n309_;wire new_n310_;wire new_n311_;wire new_n312_;wire new_n313_;wire new_n314_;wire new_n315_;wire new_n316_;wire new_n317_;wire new_n318_;wire new_n319_;wire new_n320_;wire new_n321_;wire new_n323_;wire new_n324_;wire new_n325_;wire new_n326_;wire new_n327_;wire new_n328_;wire new_n329_;wire new_n330_;wire new_n331_;wire new_n332_;wire new_n333_;wire new_n334_;wire new_n335_;wire new_n336_;wire new_n337_;wire new_n338_;wire new_n339_;wire new_n340_;wire new_n341_;wire new_n342_;wire new_n343_;wire new_n344_;wire new_n345_;wire new_n346_;wire new_n347_;wire new_n348_;wire new_n349_;wire new_n350_;wire new_n351_;wire new_n352_;wire new_n353_;wire new_n354_;wire new_n355_;wire new_n356_;wire new_n357_;wire new_n358_;wire new_n359_;wire new_n360_;wire new_n361_;wire new_n362_;wire new_n363_;wire new_n364_;wire new_n365_;wire new_n366_;wire new_n367_;wire new_n368_;wire new_n369_;wire new_n370_;wire new_n371_;wire new_n372_;wire new_n373_;wire new_n374_;wire new_n375_;wire new_n376_;wire new_n377_;wire new_n378_;wire new_n379_;wire new_n380_;wire new_n381_;wire new_n382_;wire new_n383_;wire new_n384_;wire new_n385_;wire new_n386_;wire new_n387_;wire new_n388_;wire new_n389_;wire new_n391_;wire new_n392_;wire new_n393_;wire new_n394_;wire new_n395_;wire new_n396_;wire new_n397_;wire new_n398_;wire new_n399_;wire new_n400_;wire new_n401_;wire new_n402_;wire new_n403_;wire new_n404_;wire new_n405_;wire new_n406_;wire new_n407_;wire new_n408_;wire new_n409_;wire new_n410_;wire new_n411_;wire new_n412_;wire new_n413_;wire new_n414_;wire new_n415_;wire new_n416_;wire new_n417_;wire new_n418_;wire new_n419_;wire new_n420_;wire new_n421_;wire new_n422_;wire new_n423_;wire new_n424_;wire new_n425_;wire new_n426_;wire new_n427_;wire new_n428_;wire new_n429_;wire new_n430_;wire new_n431_;wire new_n432_;wire new_n433_;wire new_n434_;wire new_n435_;wire new_n436_;wire new_n437_;wire new_n438_;wire new_n439_;wire new_n440_;wire new_n441_;wire new_n442_;wire new_n443_;wire new_n444_;wire new_n445_;wire new_n446_;wire new_n447_;wire new_n448_;wire new_n449_;wire new_n450_;wire new_n451_;wire new_n452_;wire new_n453_;wire new_n454_;wire new_n455_;wire new_n456_;wire new_n457_;wire new_n458_;wire new_n459_;wire new_n460_;wire new_n461_;wire new_n462_;wire new_n463_;wire new_n464_;wire new_n465_;wire new_n467_;wire new_n468_;wire new_n469_;wire new_n470_;wire new_n471_;wire new_n472_;wire new_n473_;wire new_n474_;wire new_n475_;wire new_n476_;wire new_n477_;wire new_n478_;wire new_n479_;wire new_n480_;wire new_n481_;wire new_n482_;wire new_n483_;wire new_n484_;wire new_n485_;wire new_n486_;wire new_n487_;wire new_n488_;wire new_n489_;wire new_n490_;wire new_n491_;wire new_n492_;wire new_n493_;wire new_n494_;wire new_n495_;wire new_n496_;wire new_n497_;wire new_n498_;wire new_n499_;wire new_n500_;wire new_n501_;wire new_n502_;wire new_n503_;wire new_n504_;wire new_n505_;wire new_n506_;wire new_n507_;wire new_n508_;wire new_n509_;wire new_n510_;wire new_n511_;wire new_n512_;wire new_n513_;wire new_n514_;wire new_n515_;wire new_n516_;wire new_n517_;wire new_n518_;wire new_n519_;wire new_n520_;wire new_n521_;wire new_n522_;wire new_n523_;wire new_n524_;wire new_n525_;wire new_n526_;wire new_n527_;wire new_n528_;wire new_n529_;wire new_n530_;wire new_n531_;wire new_n532_;wire new_n533_;wire new_n534_;wire new_n535_;wire new_n536_;wire new_n537_;wire new_n538_;wire new_n539_;wire new_n540_;wire new_n541_;wire new_n542_;wire new_n543_;wire new_n544_;wire new_n545_;wire new_n546_;wire new_n547_;wire new_n548_;wire new_n549_;wire new_n551_;wire new_n552_;wire new_n553_;wire new_n554_;wire new_n555_;wire new_n556_;wire new_n557_;wire new_n558_;wire new_n559_;wire new_n560_;wire new_n561_;wire new_n562_;wire new_n563_;wire new_n564_;wire new_n565_;wire new_n566_;wire new_n567_;wire new_n568_;wire new_n569_;wire new_n570_;wire new_n571_;wire new_n572_;wire new_n573_;wire new_n574_;wire new_n575_;wire new_n576_;wire new_n577_;wire new_n578_;wire new_n579_;wire new_n580_;wire new_n581_;wire new_n582_;wire new_n583_;wire new_n584_;wire new_n585_;wire new_n586_;wire new_n587_;wire new_n588_;wire new_n589_;wire new_n590_;wire new_n591_;wire new_n592_;wire new_n593_;wire new_n594_;wire new_n595_;wire new_n596_;wire new_n597_;wire new_n598_;wire new_n599_;wire new_n600_;wire new_n601_;wire new_n602_;wire new_n603_;wire new_n604_;wire new_n605_;wire new_n606_;wire new_n607_;wire new_n608_;wire new_n609_;wire new_n610_;wire new_n611_;wire new_n612_;wire new_n613_;wire new_n614_;wire new_n615_;wire new_n616_;wire new_n617_;wire new_n618_;wire new_n619_;wire new_n620_;wire new_n621_;wire new_n622_;wire new_n623_;wire new_n624_;wire new_n625_;wire new_n626_;wire new_n627_;wire new_n628_;wire new_n629_;wire new_n630_;wire new_n631_;wire new_n632_;wire new_n633_;wire new_n634_;wire new_n635_;wire new_n636_;wire new_n637_;wire new_n638_;wire new_n639_;wire new_n640_;wire new_n641_;wire new_n643_;wire new_n644_;wire new_n645_;wire new_n646_;wire new_n647_;wire new_n648_;wire new_n649_;wire new_n650_;wire new_n651_;wire new_n652_;wire new_n653_;wire new_n654_;wire new_n655_;wire new_n656_;wire new_n657_;wire new_n658_;wire new_n659_;wire new_n660_;wire new_n661_;wire new_n662_;wire new_n663_;wire new_n664_;wire new_n665_;wire new_n666_;wire new_n667_;wire new_n668_;wire new_n669_;wire new_n670_;wire new_n671_;wire new_n672_;wire new_n673_;wire new_n674_;wire new_n675_;wire new_n676_;wire new_n677_;wire new_n678_;wire new_n679_;wire new_n680_;wire new_n681_;wire new_n682_;wire new_n683_;wire new_n684_;wire new_n685_;wire new_n686_;wire new_n687_;wire new_n688_;wire new_n689_;wire new_n690_;wire new_n691_;wire new_n692_;wire new_n693_;wire new_n694_;wire new_n695_;wire new_n696_;wire new_n697_;wire new_n698_;wire new_n699_;wire new_n700_;wire new_n701_;wire new_n702_;wire new_n703_;wire new_n704_;wire new_n705_;wire new_n706_;wire new_n707_;wire new_n708_;wire new_n709_;wire new_n710_;wire new_n711_;wire new_n712_;wire new_n713_;wire new_n714_;wire new_n715_;wire new_n716_;wire new_n717_;wire new_n718_;wire new_n719_;wire new_n720_;wire new_n721_;wire new_n722_;wire new_n723_;wire new_n724_;wire new_n725_;wire new_n726_;wire new_n727_;wire new_n728_;wire new_n729_;wire new_n730_;wire new_n731_;wire new_n732_;wire new_n733_;wire new_n734_;wire new_n735_;wire new_n736_;wire new_n737_;wire new_n738_;wire new_n739_;wire new_n740_;wire new_n741_;wire new_n743_;wire new_n744_;wire new_n745_;wire new_n746_;wire new_n747_;wire new_n748_;wire new_n749_;wire new_n750_;wire new_n751_;wire new_n752_;wire new_n753_;wire new_n754_;wire new_n755_;wire new_n756_;wire new_n757_;wire new_n758_;wire new_n759_;wire new_n760_;wire new_n761_;wire new_n762_;wire new_n763_;wire new_n764_;wire new_n765_;wire new_n766_;wire new_n767_;wire new_n768_;wire new_n769_;wire new_n770_;wire new_n771_;wire new_n772_;wire new_n773_;wire new_n774_;wire new_n775_;wire new_n776_;wire new_n777_;wire new_n778_;wire new_n779_;wire new_n780_;wire new_n781_;wire new_n782_;wire new_n783_;wire new_n784_;wire new_n785_;wire new_n786_;wire new_n787_;wire new_n788_;wire new_n789_;wire new_n790_;wire new_n791_;wire new_n792_;wire new_n793_;wire new_n794_;wire new_n795_;wire new_n796_;wire new_n797_;wire new_n798_;wire new_n799_;wire new_n800_;wire new_n801_;wire new_n802_;wire new_n803_;wire new_n804_;wire new_n805_;wire new_n806_;wire new_n807_;wire new_n808_;wire new_n809_;wire new_n810_;wire new_n811_;wire new_n812_;wire new_n813_;wire new_n814_;wire new_n815_;wire new_n816_;wire new_n817_;wire new_n818_;wire new_n819_;wire new_n820_;wire new_n821_;wire new_n822_;wire new_n823_;wire new_n824_;wire new_n825_;wire new_n826_;wire new_n827_;wire new_n828_;wire new_n829_;wire new_n830_;wire new_n831_;wire new_n832_;wire new_n833_;wire new_n834_;wire new_n835_;wire new_n836_;wire new_n837_;wire new_n838_;wire new_n839_;wire new_n840_;wire new_n841_;wire new_n842_;wire new_n843_;wire new_n844_;wire new_n845_;wire new_n846_;wire new_n847_;wire new_n848_;wire new_n849_;wire new_n851_;wire new_n852_;wire new_n853_;wire new_n854_;wire new_n855_;wire new_n856_;wire new_n857_;wire new_n858_;wire new_n859_;wire new_n860_;wire new_n861_;wire new_n862_;wire new_n863_;wire new_n864_;wire new_n865_;wire new_n866_;wire new_n867_;wire new_n868_;wire new_n869_;wire new_n870_;wire new_n871_;wire new_n872_;wire new_n873_;wire new_n874_;wire new_n875_;wire new_n876_;wire new_n877_;wire new_n878_;wire new_n879_;wire new_n880_;wire new_n881_;wire new_n882_;wire new_n883_;wire new_n884_;wire new_n885_;wire new_n886_;wire new_n887_;wire new_n888_;wire new_n889_;wire new_n890_;wire new_n891_;wire new_n892_;wire new_n893_;wire new_n894_;wire new_n895_;wire new_n896_;wire new_n897_;wire new_n898_;wire new_n899_;wire new_n900_;wire new_n901_;wire new_n902_;wire new_n903_;wire new_n904_;wire new_n905_;wire new_n906_;wire new_n907_;wire new_n908_;wire new_n909_;wire new_n910_;wire new_n911_;wire new_n912_;wire new_n913_;wire new_n914_;wire new_n915_;wire new_n916_;wire new_n917_;wire new_n918_;wire new_n919_;wire new_n920_;wire new_n921_;wire new_n922_;wire new_n923_;wire new_n924_;wire new_n925_;wire new_n926_;wire new_n927_;wire new_n928_;wire new_n929_;wire new_n930_;wire new_n931_;wire new_n932_;wire new_n933_;wire new_n934_;wire new_n935_;wire new_n936_;wire new_n937_;wire new_n938_;wire new_n939_;wire new_n940_;wire new_n941_;wire new_n942_;wire new_n943_;wire new_n944_;wire new_n945_;wire new_n946_;wire new_n947_;wire new_n948_;wire new_n949_;wire new_n950_;wire new_n951_;wire new_n952_;wire new_n953_;wire new_n954_;wire new_n955_;wire new_n956_;wire new_n957_;wire new_n958_;wire new_n959_;wire new_n960_;wire new_n961_;wire new_n962_;wire new_n963_;wire new_n964_;wire new_n965_;wire new_n967_;wire new_n968_;wire new_n969_;wire new_n970_;wire new_n971_;wire new_n972_;wire new_n973_;wire new_n974_;wire new_n975_;wire new_n976_;wire new_n977_;wire new_n978_;wire new_n979_;wire new_n980_;wire new_n981_;wire new_n982_;wire new_n983_;wire new_n984_;wire new_n985_;wire new_n986_;wire new_n987_;wire new_n988_;wire new_n989_;wire new_n990_;wire new_n991_;wire new_n992_;wire new_n993_;wire new_n994_;wire new_n995_;wire new_n996_;wire new_n997_;wire new_n998_;wire new_n999_;wire new_n1000_;wire new_n1001_;wire new_n1002_;wire new_n1003_;wire new_n1004_;wire new_n1005_;wire new_n1006_;wire new_n1007_;wire new_n1008_;wire new_n1009_;wire new_n1010_;wire new_n1011_;wire new_n1012_;wire new_n1013_;wire new_n1014_;wire new_n1015_;wire new_n1016_;wire new_n1017_;wire new_n1018_;wire new_n1019_;wire new_n1020_;wire new_n1021_;wire new_n1022_;wire new_n1023_;wire new_n1024_;wire new_n1025_;wire new_n1026_;wire new_n1027_;wire new_n1028_;wire new_n1029_;wire new_n1030_;wire new_n1031_;wire new_n1032_;wire new_n1033_;wire new_n1034_;wire new_n1035_;wire new_n1036_;wire new_n1037_;wire new_n1038_;wire new_n1039_;wire new_n1040_;wire new_n1041_;wire new_n1042_;wire new_n1043_;wire new_n1044_;wire new_n1045_;wire new_n1046_;wire new_n1047_;wire new_n1048_;wire new_n1049_;wire new_n1050_;wire new_n1051_;wire new_n1052_;wire new_n1053_;wire new_n1054_;wire new_n1055_;wire new_n1056_;wire new_n1057_;wire new_n1058_;wire new_n1059_;wire new_n1060_;wire new_n1061_;wire new_n1062_;wire new_n1063_;wire new_n1064_;wire new_n1065_;wire new_n1066_;wire new_n1067_;wire new_n1068_;wire new_n1069_;wire new_n1070_;wire new_n1071_;wire new_n1072_;wire new_n1073_;wire new_n1074_;wire new_n1075_;wire new_n1076_;wire new_n1077_;wire new_n1078_;wire new_n1079_;wire new_n1081_;wire new_n1082_;wire new_n1083_;wire new_n1084_;wire new_n1085_;wire new_n1086_;wire new_n1087_;wire new_n1088_;wire new_n1089_;wire new_n1090_;wire new_n1091_;wire new_n1092_;wire new_n1093_;wire new_n1094_;wire new_n1095_;wire new_n1096_;wire new_n1097_;wire new_n1098_;wire new_n1099_;wire new_n1100_;wire new_n1101_;wire new_n1102_;wire new_n1103_;wire new_n1104_;wire new_n1105_;wire new_n1106_;wire new_n1107_;wire new_n1108_;wire new_n1109_;wire new_n1110_;wire new_n1111_;wire new_n1112_;wire new_n1113_;wire new_n1114_;wire new_n1115_;wire new_n1116_;wire new_n1117_;wire new_n1118_;wire new_n1119_;wire new_n1120_;wire new_n1121_;wire new_n1122_;wire new_n1123_;wire new_n1124_;wire new_n1125_;wire new_n1126_;wire new_n1127_;wire new_n1128_;wire new_n1129_;wire new_n1130_;wire new_n1131_;wire new_n1132_;wire new_n1133_;wire new_n1134_;wire new_n1135_;wire new_n1136_;wire new_n1137_;wire new_n1138_;wire new_n1139_;wire new_n1140_;wire new_n1141_;wire new_n1142_;wire new_n1143_;wire new_n1144_;wire new_n1145_;wire new_n1146_;wire new_n1147_;wire new_n1148_;wire new_n1149_;wire new_n1150_;wire new_n1151_;wire new_n1152_;wire new_n1153_;wire new_n1154_;wire new_n1155_;wire new_n1156_;wire new_n1157_;wire new_n1158_;wire new_n1159_;wire new_n1160_;wire new_n1161_;wire new_n1162_;wire new_n1163_;wire new_n1164_;wire new_n1165_;wire new_n1166_;wire new_n1167_;wire new_n1168_;wire new_n1169_;wire new_n1170_;wire new_n1171_;wire new_n1172_;wire new_n1173_;wire new_n1174_;wire new_n1175_;wire new_n1176_;wire new_n1177_;wire new_n1178_;wire new_n1179_;wire new_n1180_;wire new_n1181_;wire new_n1182_;wire new_n1183_;wire new_n1184_;wire new_n1185_;wire new_n1186_;wire new_n1187_;wire new_n1188_;wire new_n1189_;wire new_n1190_;wire new_n1191_;wire new_n1193_;wire new_n1194_;wire new_n1195_;wire new_n1196_;wire new_n1197_;wire new_n1198_;wire new_n1199_;wire new_n1200_;wire new_n1201_;wire new_n1202_;wire new_n1203_;wire new_n1204_;wire new_n1205_;wire new_n1206_;wire new_n1207_;wire new_n1208_;wire new_n1209_;wire new_n1210_;wire new_n1211_;wire new_n1212_;wire new_n1213_;wire new_n1214_;wire new_n1215_;wire new_n1216_;wire new_n1217_;wire new_n1218_;wire new_n1219_;wire new_n1220_;wire new_n1221_;wire new_n1222_;wire new_n1223_;wire new_n1224_;wire new_n1225_;wire new_n1226_;wire new_n1227_;wire new_n1228_;wire new_n1229_;wire new_n1230_;wire new_n1231_;wire new_n1232_;wire new_n1233_;wire new_n1234_;wire new_n1235_;wire new_n1236_;wire new_n1237_;wire new_n1238_;wire new_n1239_;wire new_n1240_;wire new_n1241_;wire new_n1242_;wire new_n1243_;wire new_n1244_;wire new_n1245_;wire new_n1246_;wire new_n1247_;wire new_n1248_;wire new_n1249_;wire new_n1250_;wire new_n1251_;wire new_n1252_;wire new_n1253_;wire new_n1254_;wire new_n1255_;wire new_n1256_;wire new_n1257_;wire new_n1258_;wire new_n1259_;wire new_n1260_;wire new_n1261_;wire new_n1262_;wire new_n1263_;wire new_n1264_;wire new_n1265_;wire new_n1266_;wire new_n1267_;wire new_n1268_;wire new_n1269_;wire new_n1270_;wire new_n1271_;wire new_n1272_;wire new_n1273_;wire new_n1274_;wire new_n1275_;wire new_n1276_;wire new_n1277_;wire new_n1278_;wire new_n1279_;wire new_n1280_;wire new_n1281_;wire new_n1282_;wire new_n1283_;wire new_n1284_;wire new_n1285_;wire new_n1286_;wire new_n1287_;wire new_n1288_;wire new_n1289_;wire new_n1290_;wire new_n1291_;wire new_n1292_;wire new_n1293_;wire new_n1294_;wire new_n1295_;wire new_n1296_;wire new_n1298_;wire new_n1299_;wire new_n1300_;wire new_n1301_;wire new_n1302_;wire new_n1303_;wire new_n1304_;wire new_n1305_;wire new_n1306_;wire new_n1307_;wire new_n1308_;wire new_n1309_;wire new_n1310_;wire new_n1311_;wire new_n1312_;wire new_n1313_;wire new_n1314_;wire new_n1315_;wire new_n1316_;wire new_n1317_;wire new_n1318_;wire new_n1319_;wire new_n1320_;wire new_n1321_;wire new_n1322_;wire new_n1323_;wire new_n1324_;wire new_n1325_;wire new_n1326_;wire new_n1327_;wire new_n1328_;wire new_n1329_;wire new_n1330_;wire new_n1331_;wire new_n1332_;wire new_n1333_;wire new_n1334_;wire new_n1335_;wire new_n1336_;wire new_n1337_;wire new_n1338_;wire new_n1339_;wire new_n1340_;wire new_n1341_;wire new_n1342_;wire new_n1343_;wire new_n1344_;wire new_n1345_;wire new_n1346_;wire new_n1347_;wire new_n1348_;wire new_n1349_;wire new_n1350_;wire new_n1351_;wire new_n1352_;wire new_n1353_;wire new_n1354_;wire new_n1355_;wire new_n1356_;wire new_n1357_;wire new_n1358_;wire new_n1359_;wire new_n1360_;wire new_n1361_;wire new_n1362_;wire new_n1363_;wire new_n1364_;wire new_n1365_;wire new_n1366_;wire new_n1367_;wire new_n1368_;wire new_n1369_;wire new_n1370_;wire new_n1371_;wire new_n1372_;wire new_n1373_;wire new_n1374_;wire new_n1375_;wire new_n1376_;wire new_n1377_;wire new_n1378_;wire new_n1379_;wire new_n1380_;wire new_n1381_;wire new_n1382_;wire new_n1383_;wire new_n1384_;wire new_n1385_;wire new_n1386_;wire new_n1387_;wire new_n1388_;wire new_n1389_;wire new_n1390_;wire new_n1391_;wire new_n1392_;wire new_n1393_;wire new_n1395_;wire new_n1396_;wire new_n1397_;wire new_n1398_;wire new_n1399_;wire new_n1400_;wire new_n1401_;wire new_n1402_;wire new_n1403_;wire new_n1404_;wire new_n1405_;wire new_n1406_;wire new_n1407_;wire new_n1408_;wire new_n1409_;wire new_n1410_;wire new_n1411_;wire new_n1412_;wire new_n1413_;wire new_n1414_;wire new_n1415_;wire new_n1416_;wire new_n1417_;wire new_n1418_;wire new_n1419_;wire new_n1420_;wire new_n1421_;wire new_n1422_;wire new_n1423_;wire new_n1424_;wire new_n1425_;wire new_n1426_;wire new_n1427_;wire new_n1428_;wire new_n1429_;wire new_n1430_;wire new_n1431_;wire new_n1432_;wire new_n1433_;wire new_n1434_;wire new_n1435_;wire new_n1436_;wire new_n1437_;wire new_n1438_;wire new_n1439_;wire new_n1440_;wire new_n1441_;wire new_n1442_;wire new_n1443_;wire new_n1444_;wire new_n1445_;wire new_n1446_;wire new_n1447_;wire new_n1448_;wire new_n1449_;wire new_n1450_;wire new_n1451_;wire new_n1452_;wire new_n1453_;wire new_n1454_;wire new_n1455_;wire new_n1456_;wire new_n1457_;wire new_n1458_;wire new_n1459_;wire new_n1460_;wire new_n1461_;wire new_n1462_;wire new_n1463_;wire new_n1464_;wire new_n1465_;wire new_n1466_;wire new_n1467_;wire new_n1468_;wire new_n1469_;wire new_n1470_;wire new_n1471_;wire new_n1472_;wire new_n1473_;wire new_n1474_;wire new_n1475_;wire new_n1476_;wire new_n1477_;wire new_n1478_;wire new_n1479_;wire new_n1480_;wire new_n1481_;wire new_n1482_;wire new_n1484_;wire new_n1485_;wire new_n1486_;wire new_n1487_;wire new_n1488_;wire new_n1489_;wire new_n1490_;wire new_n1491_;wire new_n1492_;wire new_n1493_;wire new_n1494_;wire new_n1495_;wire new_n1496_;wire new_n1497_;wire new_n1498_;wire new_n1499_;wire new_n1500_;wire new_n1501_;wire new_n1502_;wire new_n1503_;wire new_n1504_;wire new_n1505_;wire new_n1506_;wire new_n1507_;wire new_n1508_;wire new_n1509_;wire new_n1510_;wire new_n1511_;wire new_n1512_;wire new_n1513_;wire new_n1514_;wire new_n1515_;wire new_n1516_;wire new_n1517_;wire new_n1518_;wire new_n1519_;wire new_n1520_;wire new_n1521_;wire new_n1522_;wire new_n1523_;wire new_n1524_;wire new_n1525_;wire new_n1526_;wire new_n1527_;wire new_n1528_;wire new_n1529_;wire new_n1530_;wire new_n1531_;wire new_n1532_;wire new_n1533_;wire new_n1534_;wire new_n1535_;wire new_n1536_;wire new_n1537_;wire new_n1538_;wire new_n1539_;wire new_n1540_;wire new_n1541_;wire new_n1542_;wire new_n1543_;wire new_n1544_;wire new_n1545_;wire new_n1546_;wire new_n1547_;wire new_n1548_;wire new_n1549_;wire new_n1550_;wire new_n1551_;wire new_n1552_;wire new_n1553_;wire new_n1554_;wire new_n1555_;wire new_n1556_;wire new_n1557_;wire new_n1558_;wire new_n1559_;wire new_n1560_;wire new_n1561_;wire new_n1562_;wire new_n1563_;wire new_n1565_;wire new_n1566_;wire new_n1567_;wire new_n1568_;wire new_n1569_;wire new_n1570_;wire new_n1571_;wire new_n1572_;wire new_n1573_;wire new_n1574_;wire new_n1575_;wire new_n1576_;wire new_n1577_;wire new_n1578_;wire new_n1579_;wire new_n1580_;wire new_n1581_;wire new_n1582_;wire new_n1583_;wire new_n1584_;wire new_n1585_;wire new_n1586_;wire new_n1587_;wire new_n1588_;wire new_n1589_;wire new_n1590_;wire new_n1591_;wire new_n1592_;wire new_n1593_;wire new_n1594_;wire new_n1595_;wire new_n1596_;wire new_n1597_;wire new_n1598_;wire new_n1599_;wire new_n1600_;wire new_n1601_;wire new_n1602_;wire new_n1603_;wire new_n1604_;wire new_n1605_;wire new_n1606_;wire new_n1607_;wire new_n1608_;wire new_n1609_;wire new_n1610_;wire new_n1611_;wire new_n1612_;wire new_n1613_;wire new_n1614_;wire new_n1615_;wire new_n1616_;wire new_n1617_;wire new_n1618_;wire new_n1619_;wire new_n1620_;wire new_n1621_;wire new_n1622_;wire new_n1623_;wire new_n1624_;wire new_n1625_;wire new_n1626_;wire new_n1627_;wire new_n1628_;wire new_n1629_;wire new_n1630_;wire new_n1631_;wire new_n1632_;wire new_n1633_;wire new_n1634_;wire new_n1635_;wire new_n1636_;wire new_n1638_;wire new_n1639_;wire new_n1640_;wire new_n1641_;wire new_n1642_;wire new_n1643_;wire new_n1644_;wire new_n1645_;wire new_n1646_;wire new_n1647_;wire new_n1648_;wire new_n1649_;wire new_n1650_;wire new_n1651_;wire new_n1652_;wire new_n1653_;wire new_n1654_;wire new_n1655_;wire new_n1656_;wire new_n1657_;wire new_n1658_;wire new_n1659_;wire new_n1660_;wire new_n1661_;wire new_n1662_;wire new_n1663_;wire new_n1664_;wire new_n1665_;wire new_n1666_;wire new_n1667_;wire new_n1668_;wire new_n1669_;wire new_n1670_;wire new_n1671_;wire new_n1672_;wire new_n1673_;wire new_n1674_;wire new_n1675_;wire new_n1676_;wire new_n1677_;wire new_n1678_;wire new_n1679_;wire new_n1680_;wire new_n1681_;wire new_n1682_;wire new_n1683_;wire new_n1684_;wire new_n1685_;wire new_n1686_;wire new_n1687_;wire new_n1688_;wire new_n1689_;wire new_n1690_;wire new_n1691_;wire new_n1692_;wire new_n1693_;wire new_n1694_;wire new_n1695_;wire new_n1696_;wire new_n1697_;wire new_n1698_;wire new_n1699_;wire new_n1700_;wire new_n1701_;wire new_n1703_;wire new_n1704_;wire new_n1705_;wire new_n1706_;wire new_n1707_;wire new_n1708_;wire new_n1709_;wire new_n1710_;wire new_n1711_;wire new_n1712_;wire new_n1713_;wire new_n1714_;wire new_n1715_;wire new_n1716_;wire new_n1717_;wire new_n1718_;wire new_n1719_;wire new_n1720_;wire new_n1721_;wire new_n1722_;wire new_n1723_;wire new_n1724_;wire new_n1725_;wire new_n1726_;wire new_n1727_;wire new_n1728_;wire new_n1729_;wire new_n1730_;wire new_n1731_;wire new_n1732_;wire new_n1733_;wire new_n1734_;wire new_n1735_;wire new_n1736_;wire new_n1737_;wire new_n1738_;wire new_n1739_;wire new_n1740_;wire new_n1741_;wire new_n1742_;wire new_n1743_;wire new_n1744_;wire new_n1745_;wire new_n1746_;wire new_n1747_;wire new_n1748_;wire new_n1749_;wire new_n1750_;wire new_n1751_;wire new_n1752_;wire new_n1753_;wire new_n1754_;wire new_n1755_;wire new_n1756_;wire new_n1757_;wire new_n1758_;wire new_n1760_;wire new_n1761_;wire new_n1762_;wire new_n1763_;wire new_n1764_;wire new_n1765_;wire new_n1766_;wire new_n1767_;wire new_n1768_;wire new_n1769_;wire new_n1770_;wire new_n1771_;wire new_n1772_;wire new_n1773_;wire new_n1774_;wire new_n1775_;wire new_n1776_;wire new_n1777_;wire new_n1778_;wire new_n1779_;wire new_n1780_;wire new_n1781_;wire new_n1782_;wire new_n1783_;wire new_n1784_;wire new_n1785_;wire new_n1786_;wire new_n1787_;wire new_n1788_;wire new_n1789_;wire new_n1790_;wire new_n1791_;wire new_n1792_;wire new_n1793_;wire new_n1794_;wire new_n1795_;wire new_n1796_;wire new_n1797_;wire new_n1798_;wire new_n1799_;wire new_n1800_;wire new_n1801_;wire new_n1802_;wire new_n1803_;wire new_n1804_;wire new_n1805_;wire new_n1806_;wire new_n1807_;wire new_n1809_;wire new_n1810_;wire new_n1811_;wire new_n1812_;wire new_n1813_;wire new_n1814_;wire new_n1815_;wire new_n1816_;wire new_n1817_;wire new_n1818_;wire new_n1819_;wire new_n1820_;wire new_n1821_;wire new_n1822_;wire new_n1823_;wire new_n1824_;wire new_n1825_;wire new_n1826_;wire new_n1827_;wire new_n1828_;wire new_n1829_;wire new_n1830_;wire new_n1831_;wire new_n1832_;wire new_n1833_;wire new_n1834_;wire new_n1835_;wire new_n1836_;wire new_n1837_;wire new_n1838_;wire new_n1839_;wire new_n1840_;wire new_n1841_;wire new_n1842_;wire new_n1843_;wire new_n1844_;wire new_n1845_;wire new_n1846_;wire new_n1847_;wire new_n1848_;wire new_n1850_;wire new_n1851_;wire new_n1852_;wire new_n1853_;wire new_n1854_;wire new_n1855_;wire new_n1856_;wire new_n1857_;wire new_n1858_;wire new_n1859_;wire new_n1860_;wire new_n1861_;wire new_n1862_;wire new_n1863_;wire new_n1864_;wire new_n1865_;wire new_n1866_;wire new_n1867_;wire new_n1868_;wire new_n1869_;wire new_n1870_;wire new_n1871_;wire new_n1872_;wire new_n1873_;wire new_n1874_;wire new_n1875_;wire new_n1876_;wire new_n1877_;wire new_n1878_;wire new_n1879_;wire new_n1880_;wire new_n1881_;wire new_n1883_;wire new_n1884_;wire new_n1885_;wire new_n1886_;wire new_n1887_;wire new_n1888_;wire new_n1889_;wire new_n1890_;wire new_n1891_;wire new_n1892_;wire new_n1893_;wire new_n1894_;wire new_n1895_;wire new_n1896_;wire new_n1897_;wire new_n1898_;wire new_n1899_;wire new_n1900_;wire new_n1901_;wire new_n1902_;wire new_n1903_;wire new_n1904_;wire new_n1905_;wire new_n1906_;wire new_n1908_;wire new_n1909_;wire new_n1910_;wire new_n1911_;wire new_n1912_;wire new_n1913_;wire new_n1914_;wire new_n1915_;wire new_n1916_;wire new_n1917_;wire new_n1918_;wire new_n1919_;wire new_n1920_;wire new_n1921_;wire new_n1922_;wire new_n1923_;wire new_n1925_;wire new_n1926_;wire new_n1927_;wire new_n1928_;wire new_n1929_;wire new_n1930_;wire new_n1931_;wire new_n1933_;
  wire G1_spl_;
  wire G1_spl_0;
  wire G1_spl_00;
  wire G1_spl_000;
  wire G1_spl_001;
  wire G1_spl_01;
  wire G1_spl_010;
  wire G1_spl_011;
  wire G1_spl_1;
  wire G1_spl_10;
  wire G1_spl_100;
  wire G1_spl_101;
  wire G1_spl_11;
  wire G1_spl_110;
  wire G1_spl_111;
  wire G17_spl_;
  wire G17_spl_0;
  wire G17_spl_00;
  wire G17_spl_000;
  wire G17_spl_001;
  wire G17_spl_01;
  wire G17_spl_010;
  wire G17_spl_011;
  wire G17_spl_1;
  wire G17_spl_10;
  wire G17_spl_100;
  wire G17_spl_101;
  wire G17_spl_11;
  wire G17_spl_110;
  wire G17_spl_111;
  wire G2_spl_;
  wire G2_spl_0;
  wire G2_spl_00;
  wire G2_spl_000;
  wire G2_spl_001;
  wire G2_spl_01;
  wire G2_spl_010;
  wire G2_spl_011;
  wire G2_spl_1;
  wire G2_spl_10;
  wire G2_spl_100;
  wire G2_spl_101;
  wire G2_spl_11;
  wire G2_spl_110;
  wire G2_spl_111;
  wire G18_spl_;
  wire G18_spl_0;
  wire G18_spl_00;
  wire G18_spl_000;
  wire G18_spl_001;
  wire G18_spl_01;
  wire G18_spl_010;
  wire G18_spl_011;
  wire G18_spl_1;
  wire G18_spl_10;
  wire G18_spl_100;
  wire G18_spl_101;
  wire G18_spl_11;
  wire G18_spl_110;
  wire G18_spl_111;
  wire new_n66__spl_;
  wire new_n67__spl_;
  wire new_n68__spl_;
  wire new_n68__spl_0;
  wire G19_spl_;
  wire G19_spl_0;
  wire G19_spl_00;
  wire G19_spl_000;
  wire G19_spl_001;
  wire G19_spl_01;
  wire G19_spl_010;
  wire G19_spl_011;
  wire G19_spl_1;
  wire G19_spl_10;
  wire G19_spl_100;
  wire G19_spl_101;
  wire G19_spl_11;
  wire G19_spl_110;
  wire G19_spl_111;
  wire G3_spl_;
  wire G3_spl_0;
  wire G3_spl_00;
  wire G3_spl_000;
  wire G3_spl_001;
  wire G3_spl_01;
  wire G3_spl_010;
  wire G3_spl_011;
  wire G3_spl_1;
  wire G3_spl_10;
  wire G3_spl_100;
  wire G3_spl_101;
  wire G3_spl_11;
  wire G3_spl_110;
  wire G3_spl_111;
  wire new_n72__spl_;
  wire new_n73__spl_;
  wire new_n74__spl_;
  wire new_n74__spl_0;
  wire new_n76__spl_;
  wire new_n77__spl_;
  wire new_n71__spl_;
  wire new_n79__spl_;
  wire new_n80__spl_;
  wire G20_spl_;
  wire G20_spl_0;
  wire G20_spl_00;
  wire G20_spl_000;
  wire G20_spl_001;
  wire G20_spl_01;
  wire G20_spl_010;
  wire G20_spl_011;
  wire G20_spl_1;
  wire G20_spl_10;
  wire G20_spl_100;
  wire G20_spl_101;
  wire G20_spl_11;
  wire G20_spl_110;
  wire G20_spl_111;
  wire G4_spl_;
  wire G4_spl_0;
  wire G4_spl_00;
  wire G4_spl_000;
  wire G4_spl_001;
  wire G4_spl_01;
  wire G4_spl_010;
  wire G4_spl_011;
  wire G4_spl_1;
  wire G4_spl_10;
  wire G4_spl_100;
  wire G4_spl_101;
  wire G4_spl_11;
  wire G4_spl_110;
  wire G4_spl_111;
  wire new_n86__spl_;
  wire new_n87__spl_;
  wire new_n88__spl_;
  wire new_n88__spl_0;
  wire new_n90__spl_;
  wire new_n91__spl_;
  wire new_n85__spl_;
  wire new_n93__spl_;
  wire new_n94__spl_;
  wire new_n84__spl_;
  wire new_n96__spl_;
  wire new_n97__spl_;
  wire new_n83__spl_;
  wire new_n99__spl_;
  wire new_n100__spl_;
  wire G21_spl_;
  wire G21_spl_0;
  wire G21_spl_00;
  wire G21_spl_000;
  wire G21_spl_001;
  wire G21_spl_01;
  wire G21_spl_010;
  wire G21_spl_011;
  wire G21_spl_1;
  wire G21_spl_10;
  wire G21_spl_100;
  wire G21_spl_101;
  wire G21_spl_11;
  wire G21_spl_110;
  wire G21_spl_111;
  wire G5_spl_;
  wire G5_spl_0;
  wire G5_spl_00;
  wire G5_spl_000;
  wire G5_spl_001;
  wire G5_spl_01;
  wire G5_spl_010;
  wire G5_spl_011;
  wire G5_spl_1;
  wire G5_spl_10;
  wire G5_spl_100;
  wire G5_spl_101;
  wire G5_spl_11;
  wire G5_spl_110;
  wire G5_spl_111;
  wire new_n108__spl_;
  wire new_n109__spl_;
  wire new_n110__spl_;
  wire new_n110__spl_0;
  wire new_n112__spl_;
  wire new_n113__spl_;
  wire new_n107__spl_;
  wire new_n115__spl_;
  wire new_n116__spl_;
  wire new_n106__spl_;
  wire new_n118__spl_;
  wire new_n119__spl_;
  wire new_n105__spl_;
  wire new_n121__spl_;
  wire new_n122__spl_;
  wire new_n104__spl_;
  wire new_n124__spl_;
  wire new_n125__spl_;
  wire new_n103__spl_;
  wire new_n127__spl_;
  wire new_n128__spl_;
  wire G22_spl_;
  wire G22_spl_0;
  wire G22_spl_00;
  wire G22_spl_000;
  wire G22_spl_001;
  wire G22_spl_01;
  wire G22_spl_010;
  wire G22_spl_011;
  wire G22_spl_1;
  wire G22_spl_10;
  wire G22_spl_100;
  wire G22_spl_101;
  wire G22_spl_11;
  wire G22_spl_110;
  wire G22_spl_111;
  wire G6_spl_;
  wire G6_spl_0;
  wire G6_spl_00;
  wire G6_spl_000;
  wire G6_spl_001;
  wire G6_spl_01;
  wire G6_spl_010;
  wire G6_spl_011;
  wire G6_spl_1;
  wire G6_spl_10;
  wire G6_spl_100;
  wire G6_spl_101;
  wire G6_spl_11;
  wire G6_spl_110;
  wire G6_spl_111;
  wire new_n138__spl_;
  wire new_n139__spl_;
  wire new_n140__spl_;
  wire new_n140__spl_0;
  wire new_n142__spl_;
  wire new_n143__spl_;
  wire new_n137__spl_;
  wire new_n145__spl_;
  wire new_n146__spl_;
  wire new_n136__spl_;
  wire new_n148__spl_;
  wire new_n149__spl_;
  wire new_n135__spl_;
  wire new_n151__spl_;
  wire new_n152__spl_;
  wire new_n134__spl_;
  wire new_n154__spl_;
  wire new_n155__spl_;
  wire new_n133__spl_;
  wire new_n157__spl_;
  wire new_n158__spl_;
  wire new_n132__spl_;
  wire new_n160__spl_;
  wire new_n161__spl_;
  wire new_n131__spl_;
  wire new_n163__spl_;
  wire new_n164__spl_;
  wire G23_spl_;
  wire G23_spl_0;
  wire G23_spl_00;
  wire G23_spl_000;
  wire G23_spl_001;
  wire G23_spl_01;
  wire G23_spl_010;
  wire G23_spl_011;
  wire G23_spl_1;
  wire G23_spl_10;
  wire G23_spl_100;
  wire G23_spl_101;
  wire G23_spl_11;
  wire G23_spl_110;
  wire G23_spl_111;
  wire G7_spl_;
  wire G7_spl_0;
  wire G7_spl_00;
  wire G7_spl_000;
  wire G7_spl_001;
  wire G7_spl_01;
  wire G7_spl_010;
  wire G7_spl_011;
  wire G7_spl_1;
  wire G7_spl_10;
  wire G7_spl_100;
  wire G7_spl_101;
  wire G7_spl_11;
  wire G7_spl_110;
  wire G7_spl_111;
  wire new_n176__spl_;
  wire new_n177__spl_;
  wire new_n178__spl_;
  wire new_n178__spl_0;
  wire new_n180__spl_;
  wire new_n181__spl_;
  wire new_n175__spl_;
  wire new_n183__spl_;
  wire new_n184__spl_;
  wire new_n174__spl_;
  wire new_n186__spl_;
  wire new_n187__spl_;
  wire new_n173__spl_;
  wire new_n189__spl_;
  wire new_n190__spl_;
  wire new_n172__spl_;
  wire new_n192__spl_;
  wire new_n193__spl_;
  wire new_n171__spl_;
  wire new_n195__spl_;
  wire new_n196__spl_;
  wire new_n170__spl_;
  wire new_n198__spl_;
  wire new_n199__spl_;
  wire new_n169__spl_;
  wire new_n201__spl_;
  wire new_n202__spl_;
  wire new_n168__spl_;
  wire new_n204__spl_;
  wire new_n205__spl_;
  wire new_n167__spl_;
  wire new_n207__spl_;
  wire new_n208__spl_;
  wire G24_spl_;
  wire G24_spl_0;
  wire G24_spl_00;
  wire G24_spl_000;
  wire G24_spl_001;
  wire G24_spl_01;
  wire G24_spl_010;
  wire G24_spl_011;
  wire G24_spl_1;
  wire G24_spl_10;
  wire G24_spl_100;
  wire G24_spl_101;
  wire G24_spl_11;
  wire G24_spl_110;
  wire G24_spl_111;
  wire G8_spl_;
  wire G8_spl_0;
  wire G8_spl_00;
  wire G8_spl_000;
  wire G8_spl_001;
  wire G8_spl_01;
  wire G8_spl_010;
  wire G8_spl_011;
  wire G8_spl_1;
  wire G8_spl_10;
  wire G8_spl_100;
  wire G8_spl_101;
  wire G8_spl_11;
  wire G8_spl_110;
  wire G8_spl_111;
  wire new_n222__spl_;
  wire new_n223__spl_;
  wire new_n224__spl_;
  wire new_n224__spl_0;
  wire new_n226__spl_;
  wire new_n227__spl_;
  wire new_n221__spl_;
  wire new_n229__spl_;
  wire new_n230__spl_;
  wire new_n220__spl_;
  wire new_n232__spl_;
  wire new_n233__spl_;
  wire new_n219__spl_;
  wire new_n235__spl_;
  wire new_n236__spl_;
  wire new_n218__spl_;
  wire new_n238__spl_;
  wire new_n239__spl_;
  wire new_n217__spl_;
  wire new_n241__spl_;
  wire new_n242__spl_;
  wire new_n216__spl_;
  wire new_n244__spl_;
  wire new_n245__spl_;
  wire new_n215__spl_;
  wire new_n247__spl_;
  wire new_n248__spl_;
  wire new_n214__spl_;
  wire new_n250__spl_;
  wire new_n251__spl_;
  wire new_n213__spl_;
  wire new_n253__spl_;
  wire new_n254__spl_;
  wire new_n212__spl_;
  wire new_n256__spl_;
  wire new_n257__spl_;
  wire new_n211__spl_;
  wire new_n259__spl_;
  wire new_n260__spl_;
  wire G25_spl_;
  wire G25_spl_0;
  wire G25_spl_00;
  wire G25_spl_000;
  wire G25_spl_001;
  wire G25_spl_01;
  wire G25_spl_010;
  wire G25_spl_011;
  wire G25_spl_1;
  wire G25_spl_10;
  wire G25_spl_100;
  wire G25_spl_101;
  wire G25_spl_11;
  wire G25_spl_110;
  wire G25_spl_111;
  wire G9_spl_;
  wire G9_spl_0;
  wire G9_spl_00;
  wire G9_spl_000;
  wire G9_spl_001;
  wire G9_spl_01;
  wire G9_spl_010;
  wire G9_spl_011;
  wire G9_spl_1;
  wire G9_spl_10;
  wire G9_spl_100;
  wire G9_spl_101;
  wire G9_spl_11;
  wire G9_spl_110;
  wire G9_spl_111;
  wire new_n276__spl_;
  wire new_n277__spl_;
  wire new_n278__spl_;
  wire new_n278__spl_0;
  wire new_n280__spl_;
  wire new_n281__spl_;
  wire new_n275__spl_;
  wire new_n283__spl_;
  wire new_n284__spl_;
  wire new_n274__spl_;
  wire new_n286__spl_;
  wire new_n287__spl_;
  wire new_n273__spl_;
  wire new_n289__spl_;
  wire new_n290__spl_;
  wire new_n272__spl_;
  wire new_n292__spl_;
  wire new_n293__spl_;
  wire new_n271__spl_;
  wire new_n295__spl_;
  wire new_n296__spl_;
  wire new_n270__spl_;
  wire new_n298__spl_;
  wire new_n299__spl_;
  wire new_n269__spl_;
  wire new_n301__spl_;
  wire new_n302__spl_;
  wire new_n268__spl_;
  wire new_n304__spl_;
  wire new_n305__spl_;
  wire new_n267__spl_;
  wire new_n307__spl_;
  wire new_n308__spl_;
  wire new_n266__spl_;
  wire new_n310__spl_;
  wire new_n311__spl_;
  wire new_n265__spl_;
  wire new_n313__spl_;
  wire new_n314__spl_;
  wire new_n264__spl_;
  wire new_n316__spl_;
  wire new_n317__spl_;
  wire new_n263__spl_;
  wire new_n319__spl_;
  wire new_n320__spl_;
  wire G26_spl_;
  wire G26_spl_0;
  wire G26_spl_00;
  wire G26_spl_000;
  wire G26_spl_001;
  wire G26_spl_01;
  wire G26_spl_010;
  wire G26_spl_011;
  wire G26_spl_1;
  wire G26_spl_10;
  wire G26_spl_100;
  wire G26_spl_101;
  wire G26_spl_11;
  wire G26_spl_110;
  wire G26_spl_111;
  wire G10_spl_;
  wire G10_spl_0;
  wire G10_spl_00;
  wire G10_spl_000;
  wire G10_spl_001;
  wire G10_spl_01;
  wire G10_spl_010;
  wire G10_spl_011;
  wire G10_spl_1;
  wire G10_spl_10;
  wire G10_spl_100;
  wire G10_spl_101;
  wire G10_spl_11;
  wire G10_spl_110;
  wire G10_spl_111;
  wire new_n338__spl_;
  wire new_n339__spl_;
  wire new_n340__spl_;
  wire new_n340__spl_0;
  wire new_n342__spl_;
  wire new_n343__spl_;
  wire new_n337__spl_;
  wire new_n345__spl_;
  wire new_n346__spl_;
  wire new_n336__spl_;
  wire new_n348__spl_;
  wire new_n349__spl_;
  wire new_n335__spl_;
  wire new_n351__spl_;
  wire new_n352__spl_;
  wire new_n334__spl_;
  wire new_n354__spl_;
  wire new_n355__spl_;
  wire new_n333__spl_;
  wire new_n357__spl_;
  wire new_n358__spl_;
  wire new_n332__spl_;
  wire new_n360__spl_;
  wire new_n361__spl_;
  wire new_n331__spl_;
  wire new_n363__spl_;
  wire new_n364__spl_;
  wire new_n330__spl_;
  wire new_n366__spl_;
  wire new_n367__spl_;
  wire new_n329__spl_;
  wire new_n369__spl_;
  wire new_n370__spl_;
  wire new_n328__spl_;
  wire new_n372__spl_;
  wire new_n373__spl_;
  wire new_n327__spl_;
  wire new_n375__spl_;
  wire new_n376__spl_;
  wire new_n326__spl_;
  wire new_n378__spl_;
  wire new_n379__spl_;
  wire new_n325__spl_;
  wire new_n381__spl_;
  wire new_n382__spl_;
  wire new_n324__spl_;
  wire new_n384__spl_;
  wire new_n385__spl_;
  wire new_n323__spl_;
  wire new_n387__spl_;
  wire new_n388__spl_;
  wire G27_spl_;
  wire G27_spl_0;
  wire G27_spl_00;
  wire G27_spl_000;
  wire G27_spl_001;
  wire G27_spl_01;
  wire G27_spl_010;
  wire G27_spl_011;
  wire G27_spl_1;
  wire G27_spl_10;
  wire G27_spl_100;
  wire G27_spl_101;
  wire G27_spl_11;
  wire G27_spl_110;
  wire G27_spl_111;
  wire G11_spl_;
  wire G11_spl_0;
  wire G11_spl_00;
  wire G11_spl_000;
  wire G11_spl_001;
  wire G11_spl_01;
  wire G11_spl_010;
  wire G11_spl_011;
  wire G11_spl_1;
  wire G11_spl_10;
  wire G11_spl_100;
  wire G11_spl_101;
  wire G11_spl_11;
  wire G11_spl_110;
  wire G11_spl_111;
  wire new_n408__spl_;
  wire new_n409__spl_;
  wire new_n410__spl_;
  wire new_n410__spl_0;
  wire new_n412__spl_;
  wire new_n413__spl_;
  wire new_n407__spl_;
  wire new_n415__spl_;
  wire new_n416__spl_;
  wire new_n406__spl_;
  wire new_n418__spl_;
  wire new_n419__spl_;
  wire new_n405__spl_;
  wire new_n421__spl_;
  wire new_n422__spl_;
  wire new_n404__spl_;
  wire new_n424__spl_;
  wire new_n425__spl_;
  wire new_n403__spl_;
  wire new_n427__spl_;
  wire new_n428__spl_;
  wire new_n402__spl_;
  wire new_n430__spl_;
  wire new_n431__spl_;
  wire new_n401__spl_;
  wire new_n433__spl_;
  wire new_n434__spl_;
  wire new_n400__spl_;
  wire new_n436__spl_;
  wire new_n437__spl_;
  wire new_n399__spl_;
  wire new_n439__spl_;
  wire new_n440__spl_;
  wire new_n398__spl_;
  wire new_n442__spl_;
  wire new_n443__spl_;
  wire new_n397__spl_;
  wire new_n445__spl_;
  wire new_n446__spl_;
  wire new_n396__spl_;
  wire new_n448__spl_;
  wire new_n449__spl_;
  wire new_n395__spl_;
  wire new_n451__spl_;
  wire new_n452__spl_;
  wire new_n394__spl_;
  wire new_n454__spl_;
  wire new_n455__spl_;
  wire new_n393__spl_;
  wire new_n457__spl_;
  wire new_n458__spl_;
  wire new_n392__spl_;
  wire new_n460__spl_;
  wire new_n461__spl_;
  wire new_n391__spl_;
  wire new_n463__spl_;
  wire new_n464__spl_;
  wire G28_spl_;
  wire G28_spl_0;
  wire G28_spl_00;
  wire G28_spl_000;
  wire G28_spl_001;
  wire G28_spl_01;
  wire G28_spl_010;
  wire G28_spl_011;
  wire G28_spl_1;
  wire G28_spl_10;
  wire G28_spl_100;
  wire G28_spl_101;
  wire G28_spl_11;
  wire G28_spl_110;
  wire G28_spl_111;
  wire G12_spl_;
  wire G12_spl_0;
  wire G12_spl_00;
  wire G12_spl_000;
  wire G12_spl_001;
  wire G12_spl_01;
  wire G12_spl_010;
  wire G12_spl_011;
  wire G12_spl_1;
  wire G12_spl_10;
  wire G12_spl_100;
  wire G12_spl_101;
  wire G12_spl_11;
  wire G12_spl_110;
  wire G12_spl_111;
  wire new_n486__spl_;
  wire new_n487__spl_;
  wire new_n488__spl_;
  wire new_n488__spl_0;
  wire new_n490__spl_;
  wire new_n491__spl_;
  wire new_n485__spl_;
  wire new_n493__spl_;
  wire new_n494__spl_;
  wire new_n484__spl_;
  wire new_n496__spl_;
  wire new_n497__spl_;
  wire new_n483__spl_;
  wire new_n499__spl_;
  wire new_n500__spl_;
  wire new_n482__spl_;
  wire new_n502__spl_;
  wire new_n503__spl_;
  wire new_n481__spl_;
  wire new_n505__spl_;
  wire new_n506__spl_;
  wire new_n480__spl_;
  wire new_n508__spl_;
  wire new_n509__spl_;
  wire new_n479__spl_;
  wire new_n511__spl_;
  wire new_n512__spl_;
  wire new_n478__spl_;
  wire new_n514__spl_;
  wire new_n515__spl_;
  wire new_n477__spl_;
  wire new_n517__spl_;
  wire new_n518__spl_;
  wire new_n476__spl_;
  wire new_n520__spl_;
  wire new_n521__spl_;
  wire new_n475__spl_;
  wire new_n523__spl_;
  wire new_n524__spl_;
  wire new_n474__spl_;
  wire new_n526__spl_;
  wire new_n527__spl_;
  wire new_n473__spl_;
  wire new_n529__spl_;
  wire new_n530__spl_;
  wire new_n472__spl_;
  wire new_n532__spl_;
  wire new_n533__spl_;
  wire new_n471__spl_;
  wire new_n535__spl_;
  wire new_n536__spl_;
  wire new_n470__spl_;
  wire new_n538__spl_;
  wire new_n539__spl_;
  wire new_n469__spl_;
  wire new_n541__spl_;
  wire new_n542__spl_;
  wire new_n468__spl_;
  wire new_n544__spl_;
  wire new_n545__spl_;
  wire new_n467__spl_;
  wire new_n547__spl_;
  wire new_n548__spl_;
  wire G29_spl_;
  wire G29_spl_0;
  wire G29_spl_00;
  wire G29_spl_000;
  wire G29_spl_001;
  wire G29_spl_01;
  wire G29_spl_010;
  wire G29_spl_011;
  wire G29_spl_1;
  wire G29_spl_10;
  wire G29_spl_100;
  wire G29_spl_101;
  wire G29_spl_11;
  wire G29_spl_110;
  wire G29_spl_111;
  wire G13_spl_;
  wire G13_spl_0;
  wire G13_spl_00;
  wire G13_spl_000;
  wire G13_spl_001;
  wire G13_spl_01;
  wire G13_spl_010;
  wire G13_spl_011;
  wire G13_spl_1;
  wire G13_spl_10;
  wire G13_spl_100;
  wire G13_spl_101;
  wire G13_spl_11;
  wire G13_spl_110;
  wire G13_spl_111;
  wire new_n572__spl_;
  wire new_n573__spl_;
  wire new_n574__spl_;
  wire new_n574__spl_0;
  wire new_n576__spl_;
  wire new_n577__spl_;
  wire new_n571__spl_;
  wire new_n579__spl_;
  wire new_n580__spl_;
  wire new_n570__spl_;
  wire new_n582__spl_;
  wire new_n583__spl_;
  wire new_n569__spl_;
  wire new_n585__spl_;
  wire new_n586__spl_;
  wire new_n568__spl_;
  wire new_n588__spl_;
  wire new_n589__spl_;
  wire new_n567__spl_;
  wire new_n591__spl_;
  wire new_n592__spl_;
  wire new_n566__spl_;
  wire new_n594__spl_;
  wire new_n595__spl_;
  wire new_n565__spl_;
  wire new_n597__spl_;
  wire new_n598__spl_;
  wire new_n564__spl_;
  wire new_n600__spl_;
  wire new_n601__spl_;
  wire new_n563__spl_;
  wire new_n603__spl_;
  wire new_n604__spl_;
  wire new_n562__spl_;
  wire new_n606__spl_;
  wire new_n607__spl_;
  wire new_n561__spl_;
  wire new_n609__spl_;
  wire new_n610__spl_;
  wire new_n560__spl_;
  wire new_n612__spl_;
  wire new_n613__spl_;
  wire new_n559__spl_;
  wire new_n615__spl_;
  wire new_n616__spl_;
  wire new_n558__spl_;
  wire new_n618__spl_;
  wire new_n619__spl_;
  wire new_n557__spl_;
  wire new_n621__spl_;
  wire new_n622__spl_;
  wire new_n556__spl_;
  wire new_n624__spl_;
  wire new_n625__spl_;
  wire new_n555__spl_;
  wire new_n627__spl_;
  wire new_n628__spl_;
  wire new_n554__spl_;
  wire new_n630__spl_;
  wire new_n631__spl_;
  wire new_n553__spl_;
  wire new_n633__spl_;
  wire new_n634__spl_;
  wire new_n552__spl_;
  wire new_n636__spl_;
  wire new_n637__spl_;
  wire new_n551__spl_;
  wire new_n639__spl_;
  wire new_n640__spl_;
  wire G30_spl_;
  wire G30_spl_0;
  wire G30_spl_00;
  wire G30_spl_000;
  wire G30_spl_001;
  wire G30_spl_01;
  wire G30_spl_010;
  wire G30_spl_011;
  wire G30_spl_1;
  wire G30_spl_10;
  wire G30_spl_100;
  wire G30_spl_101;
  wire G30_spl_11;
  wire G30_spl_110;
  wire G30_spl_111;
  wire G14_spl_;
  wire G14_spl_0;
  wire G14_spl_00;
  wire G14_spl_000;
  wire G14_spl_001;
  wire G14_spl_01;
  wire G14_spl_010;
  wire G14_spl_011;
  wire G14_spl_1;
  wire G14_spl_10;
  wire G14_spl_100;
  wire G14_spl_101;
  wire G14_spl_11;
  wire G14_spl_110;
  wire G14_spl_111;
  wire new_n666__spl_;
  wire new_n667__spl_;
  wire new_n668__spl_;
  wire new_n668__spl_0;
  wire new_n670__spl_;
  wire new_n671__spl_;
  wire new_n665__spl_;
  wire new_n673__spl_;
  wire new_n674__spl_;
  wire new_n664__spl_;
  wire new_n676__spl_;
  wire new_n677__spl_;
  wire new_n663__spl_;
  wire new_n679__spl_;
  wire new_n680__spl_;
  wire new_n662__spl_;
  wire new_n682__spl_;
  wire new_n683__spl_;
  wire new_n661__spl_;
  wire new_n685__spl_;
  wire new_n686__spl_;
  wire new_n660__spl_;
  wire new_n688__spl_;
  wire new_n689__spl_;
  wire new_n659__spl_;
  wire new_n691__spl_;
  wire new_n692__spl_;
  wire new_n658__spl_;
  wire new_n694__spl_;
  wire new_n695__spl_;
  wire new_n657__spl_;
  wire new_n697__spl_;
  wire new_n698__spl_;
  wire new_n656__spl_;
  wire new_n700__spl_;
  wire new_n701__spl_;
  wire new_n655__spl_;
  wire new_n703__spl_;
  wire new_n704__spl_;
  wire new_n654__spl_;
  wire new_n706__spl_;
  wire new_n707__spl_;
  wire new_n653__spl_;
  wire new_n709__spl_;
  wire new_n710__spl_;
  wire new_n652__spl_;
  wire new_n712__spl_;
  wire new_n713__spl_;
  wire new_n651__spl_;
  wire new_n715__spl_;
  wire new_n716__spl_;
  wire new_n650__spl_;
  wire new_n718__spl_;
  wire new_n719__spl_;
  wire new_n649__spl_;
  wire new_n721__spl_;
  wire new_n722__spl_;
  wire new_n648__spl_;
  wire new_n724__spl_;
  wire new_n725__spl_;
  wire new_n647__spl_;
  wire new_n727__spl_;
  wire new_n728__spl_;
  wire new_n646__spl_;
  wire new_n730__spl_;
  wire new_n731__spl_;
  wire new_n645__spl_;
  wire new_n733__spl_;
  wire new_n734__spl_;
  wire new_n644__spl_;
  wire new_n736__spl_;
  wire new_n737__spl_;
  wire new_n643__spl_;
  wire new_n739__spl_;
  wire new_n740__spl_;
  wire G31_spl_;
  wire G31_spl_0;
  wire G31_spl_00;
  wire G31_spl_000;
  wire G31_spl_001;
  wire G31_spl_01;
  wire G31_spl_010;
  wire G31_spl_011;
  wire G31_spl_1;
  wire G31_spl_10;
  wire G31_spl_100;
  wire G31_spl_101;
  wire G31_spl_11;
  wire G31_spl_110;
  wire G31_spl_111;
  wire G15_spl_;
  wire G15_spl_0;
  wire G15_spl_00;
  wire G15_spl_000;
  wire G15_spl_001;
  wire G15_spl_01;
  wire G15_spl_010;
  wire G15_spl_011;
  wire G15_spl_1;
  wire G15_spl_10;
  wire G15_spl_100;
  wire G15_spl_101;
  wire G15_spl_11;
  wire G15_spl_110;
  wire G15_spl_111;
  wire new_n768__spl_;
  wire new_n769__spl_;
  wire new_n770__spl_;
  wire new_n770__spl_0;
  wire new_n772__spl_;
  wire new_n773__spl_;
  wire new_n767__spl_;
  wire new_n775__spl_;
  wire new_n776__spl_;
  wire new_n766__spl_;
  wire new_n778__spl_;
  wire new_n779__spl_;
  wire new_n765__spl_;
  wire new_n781__spl_;
  wire new_n782__spl_;
  wire new_n764__spl_;
  wire new_n784__spl_;
  wire new_n785__spl_;
  wire new_n763__spl_;
  wire new_n787__spl_;
  wire new_n788__spl_;
  wire new_n762__spl_;
  wire new_n790__spl_;
  wire new_n791__spl_;
  wire new_n761__spl_;
  wire new_n793__spl_;
  wire new_n794__spl_;
  wire new_n760__spl_;
  wire new_n796__spl_;
  wire new_n797__spl_;
  wire new_n759__spl_;
  wire new_n799__spl_;
  wire new_n800__spl_;
  wire new_n758__spl_;
  wire new_n802__spl_;
  wire new_n803__spl_;
  wire new_n757__spl_;
  wire new_n805__spl_;
  wire new_n806__spl_;
  wire new_n756__spl_;
  wire new_n808__spl_;
  wire new_n809__spl_;
  wire new_n755__spl_;
  wire new_n811__spl_;
  wire new_n812__spl_;
  wire new_n754__spl_;
  wire new_n814__spl_;
  wire new_n815__spl_;
  wire new_n753__spl_;
  wire new_n817__spl_;
  wire new_n818__spl_;
  wire new_n752__spl_;
  wire new_n820__spl_;
  wire new_n821__spl_;
  wire new_n751__spl_;
  wire new_n823__spl_;
  wire new_n824__spl_;
  wire new_n750__spl_;
  wire new_n826__spl_;
  wire new_n827__spl_;
  wire new_n749__spl_;
  wire new_n829__spl_;
  wire new_n830__spl_;
  wire new_n748__spl_;
  wire new_n832__spl_;
  wire new_n833__spl_;
  wire new_n747__spl_;
  wire new_n835__spl_;
  wire new_n836__spl_;
  wire new_n746__spl_;
  wire new_n838__spl_;
  wire new_n839__spl_;
  wire new_n745__spl_;
  wire new_n841__spl_;
  wire new_n842__spl_;
  wire new_n744__spl_;
  wire new_n844__spl_;
  wire new_n845__spl_;
  wire new_n743__spl_;
  wire new_n847__spl_;
  wire new_n848__spl_;
  wire G32_spl_;
  wire G32_spl_0;
  wire G32_spl_00;
  wire G32_spl_000;
  wire G32_spl_001;
  wire G32_spl_01;
  wire G32_spl_010;
  wire G32_spl_011;
  wire G32_spl_1;
  wire G32_spl_10;
  wire G32_spl_100;
  wire G32_spl_101;
  wire G32_spl_11;
  wire G32_spl_110;
  wire G32_spl_111;
  wire G16_spl_;
  wire G16_spl_0;
  wire G16_spl_00;
  wire G16_spl_000;
  wire G16_spl_001;
  wire G16_spl_01;
  wire G16_spl_010;
  wire G16_spl_011;
  wire G16_spl_1;
  wire G16_spl_10;
  wire G16_spl_100;
  wire G16_spl_101;
  wire G16_spl_11;
  wire G16_spl_110;
  wire G16_spl_111;
  wire new_n878__spl_;
  wire new_n879__spl_;
  wire new_n880__spl_;
  wire new_n882__spl_;
  wire new_n883__spl_;
  wire new_n877__spl_;
  wire new_n885__spl_;
  wire new_n886__spl_;
  wire new_n876__spl_;
  wire new_n888__spl_;
  wire new_n889__spl_;
  wire new_n875__spl_;
  wire new_n891__spl_;
  wire new_n892__spl_;
  wire new_n874__spl_;
  wire new_n894__spl_;
  wire new_n895__spl_;
  wire new_n873__spl_;
  wire new_n897__spl_;
  wire new_n898__spl_;
  wire new_n872__spl_;
  wire new_n900__spl_;
  wire new_n901__spl_;
  wire new_n871__spl_;
  wire new_n903__spl_;
  wire new_n904__spl_;
  wire new_n870__spl_;
  wire new_n906__spl_;
  wire new_n907__spl_;
  wire new_n869__spl_;
  wire new_n909__spl_;
  wire new_n910__spl_;
  wire new_n868__spl_;
  wire new_n912__spl_;
  wire new_n913__spl_;
  wire new_n867__spl_;
  wire new_n915__spl_;
  wire new_n916__spl_;
  wire new_n866__spl_;
  wire new_n918__spl_;
  wire new_n919__spl_;
  wire new_n865__spl_;
  wire new_n921__spl_;
  wire new_n922__spl_;
  wire new_n864__spl_;
  wire new_n924__spl_;
  wire new_n925__spl_;
  wire new_n863__spl_;
  wire new_n927__spl_;
  wire new_n928__spl_;
  wire new_n862__spl_;
  wire new_n930__spl_;
  wire new_n931__spl_;
  wire new_n861__spl_;
  wire new_n933__spl_;
  wire new_n934__spl_;
  wire new_n860__spl_;
  wire new_n936__spl_;
  wire new_n937__spl_;
  wire new_n859__spl_;
  wire new_n939__spl_;
  wire new_n940__spl_;
  wire new_n858__spl_;
  wire new_n942__spl_;
  wire new_n943__spl_;
  wire new_n857__spl_;
  wire new_n945__spl_;
  wire new_n946__spl_;
  wire new_n856__spl_;
  wire new_n948__spl_;
  wire new_n949__spl_;
  wire new_n855__spl_;
  wire new_n951__spl_;
  wire new_n952__spl_;
  wire new_n854__spl_;
  wire new_n954__spl_;
  wire new_n955__spl_;
  wire new_n853__spl_;
  wire new_n957__spl_;
  wire new_n958__spl_;
  wire new_n852__spl_;
  wire new_n960__spl_;
  wire new_n961__spl_;
  wire new_n851__spl_;
  wire new_n963__spl_;
  wire new_n964__spl_;
  wire new_n994__spl_;
  wire new_n995__spl_;
  wire new_n996__spl_;
  wire new_n997__spl_;
  wire new_n993__spl_;
  wire new_n999__spl_;
  wire new_n1000__spl_;
  wire new_n992__spl_;
  wire new_n1002__spl_;
  wire new_n1003__spl_;
  wire new_n991__spl_;
  wire new_n1005__spl_;
  wire new_n1006__spl_;
  wire new_n990__spl_;
  wire new_n1008__spl_;
  wire new_n1009__spl_;
  wire new_n989__spl_;
  wire new_n1011__spl_;
  wire new_n1012__spl_;
  wire new_n988__spl_;
  wire new_n1014__spl_;
  wire new_n1015__spl_;
  wire new_n987__spl_;
  wire new_n1017__spl_;
  wire new_n1018__spl_;
  wire new_n986__spl_;
  wire new_n1020__spl_;
  wire new_n1021__spl_;
  wire new_n985__spl_;
  wire new_n1023__spl_;
  wire new_n1024__spl_;
  wire new_n984__spl_;
  wire new_n1026__spl_;
  wire new_n1027__spl_;
  wire new_n983__spl_;
  wire new_n1029__spl_;
  wire new_n1030__spl_;
  wire new_n982__spl_;
  wire new_n1032__spl_;
  wire new_n1033__spl_;
  wire new_n981__spl_;
  wire new_n1035__spl_;
  wire new_n1036__spl_;
  wire new_n980__spl_;
  wire new_n1038__spl_;
  wire new_n1039__spl_;
  wire new_n979__spl_;
  wire new_n1041__spl_;
  wire new_n1042__spl_;
  wire new_n978__spl_;
  wire new_n1044__spl_;
  wire new_n1045__spl_;
  wire new_n977__spl_;
  wire new_n1047__spl_;
  wire new_n1048__spl_;
  wire new_n976__spl_;
  wire new_n1050__spl_;
  wire new_n1051__spl_;
  wire new_n975__spl_;
  wire new_n1053__spl_;
  wire new_n1054__spl_;
  wire new_n974__spl_;
  wire new_n1056__spl_;
  wire new_n1057__spl_;
  wire new_n973__spl_;
  wire new_n1059__spl_;
  wire new_n1060__spl_;
  wire new_n972__spl_;
  wire new_n1062__spl_;
  wire new_n1063__spl_;
  wire new_n971__spl_;
  wire new_n1065__spl_;
  wire new_n1066__spl_;
  wire new_n970__spl_;
  wire new_n1068__spl_;
  wire new_n1069__spl_;
  wire new_n969__spl_;
  wire new_n1071__spl_;
  wire new_n1072__spl_;
  wire new_n968__spl_;
  wire new_n1074__spl_;
  wire new_n1075__spl_;
  wire new_n967__spl_;
  wire new_n1077__spl_;
  wire new_n1079__spl_;
  wire new_n1079__spl_0;
  wire new_n1107__spl_;
  wire new_n1108__spl_;
  wire new_n1109__spl_;
  wire new_n1106__spl_;
  wire new_n1111__spl_;
  wire new_n1112__spl_;
  wire new_n1105__spl_;
  wire new_n1114__spl_;
  wire new_n1115__spl_;
  wire new_n1104__spl_;
  wire new_n1117__spl_;
  wire new_n1118__spl_;
  wire new_n1103__spl_;
  wire new_n1120__spl_;
  wire new_n1121__spl_;
  wire new_n1102__spl_;
  wire new_n1123__spl_;
  wire new_n1124__spl_;
  wire new_n1101__spl_;
  wire new_n1126__spl_;
  wire new_n1127__spl_;
  wire new_n1100__spl_;
  wire new_n1129__spl_;
  wire new_n1130__spl_;
  wire new_n1099__spl_;
  wire new_n1132__spl_;
  wire new_n1133__spl_;
  wire new_n1098__spl_;
  wire new_n1135__spl_;
  wire new_n1136__spl_;
  wire new_n1097__spl_;
  wire new_n1138__spl_;
  wire new_n1139__spl_;
  wire new_n1096__spl_;
  wire new_n1141__spl_;
  wire new_n1142__spl_;
  wire new_n1095__spl_;
  wire new_n1144__spl_;
  wire new_n1145__spl_;
  wire new_n1094__spl_;
  wire new_n1147__spl_;
  wire new_n1148__spl_;
  wire new_n1093__spl_;
  wire new_n1150__spl_;
  wire new_n1151__spl_;
  wire new_n1092__spl_;
  wire new_n1153__spl_;
  wire new_n1154__spl_;
  wire new_n1091__spl_;
  wire new_n1156__spl_;
  wire new_n1157__spl_;
  wire new_n1090__spl_;
  wire new_n1159__spl_;
  wire new_n1160__spl_;
  wire new_n1089__spl_;
  wire new_n1162__spl_;
  wire new_n1163__spl_;
  wire new_n1088__spl_;
  wire new_n1165__spl_;
  wire new_n1166__spl_;
  wire new_n1087__spl_;
  wire new_n1168__spl_;
  wire new_n1169__spl_;
  wire new_n1086__spl_;
  wire new_n1171__spl_;
  wire new_n1172__spl_;
  wire new_n1085__spl_;
  wire new_n1174__spl_;
  wire new_n1175__spl_;
  wire new_n1084__spl_;
  wire new_n1177__spl_;
  wire new_n1178__spl_;
  wire new_n1083__spl_;
  wire new_n1180__spl_;
  wire new_n1181__spl_;
  wire new_n1082__spl_;
  wire new_n1183__spl_;
  wire new_n1184__spl_;
  wire new_n1081__spl_;
  wire new_n1186__spl_;
  wire new_n1187__spl_;
  wire new_n1189__spl_;
  wire new_n1190__spl_;
  wire new_n1218__spl_;
  wire new_n1219__spl_;
  wire new_n1220__spl_;
  wire new_n1217__spl_;
  wire new_n1222__spl_;
  wire new_n1223__spl_;
  wire new_n1216__spl_;
  wire new_n1225__spl_;
  wire new_n1226__spl_;
  wire new_n1215__spl_;
  wire new_n1228__spl_;
  wire new_n1229__spl_;
  wire new_n1214__spl_;
  wire new_n1231__spl_;
  wire new_n1232__spl_;
  wire new_n1213__spl_;
  wire new_n1234__spl_;
  wire new_n1235__spl_;
  wire new_n1212__spl_;
  wire new_n1237__spl_;
  wire new_n1238__spl_;
  wire new_n1211__spl_;
  wire new_n1240__spl_;
  wire new_n1241__spl_;
  wire new_n1210__spl_;
  wire new_n1243__spl_;
  wire new_n1244__spl_;
  wire new_n1209__spl_;
  wire new_n1246__spl_;
  wire new_n1247__spl_;
  wire new_n1208__spl_;
  wire new_n1249__spl_;
  wire new_n1250__spl_;
  wire new_n1207__spl_;
  wire new_n1252__spl_;
  wire new_n1253__spl_;
  wire new_n1206__spl_;
  wire new_n1255__spl_;
  wire new_n1256__spl_;
  wire new_n1205__spl_;
  wire new_n1258__spl_;
  wire new_n1259__spl_;
  wire new_n1204__spl_;
  wire new_n1261__spl_;
  wire new_n1262__spl_;
  wire new_n1203__spl_;
  wire new_n1264__spl_;
  wire new_n1265__spl_;
  wire new_n1202__spl_;
  wire new_n1267__spl_;
  wire new_n1268__spl_;
  wire new_n1201__spl_;
  wire new_n1270__spl_;
  wire new_n1271__spl_;
  wire new_n1200__spl_;
  wire new_n1273__spl_;
  wire new_n1274__spl_;
  wire new_n1199__spl_;
  wire new_n1276__spl_;
  wire new_n1277__spl_;
  wire new_n1198__spl_;
  wire new_n1279__spl_;
  wire new_n1280__spl_;
  wire new_n1197__spl_;
  wire new_n1282__spl_;
  wire new_n1283__spl_;
  wire new_n1196__spl_;
  wire new_n1285__spl_;
  wire new_n1286__spl_;
  wire new_n1195__spl_;
  wire new_n1288__spl_;
  wire new_n1289__spl_;
  wire new_n1194__spl_;
  wire new_n1291__spl_;
  wire new_n1292__spl_;
  wire new_n1193__spl_;
  wire new_n1294__spl_;
  wire new_n1295__spl_;
  wire new_n1321__spl_;
  wire new_n1322__spl_;
  wire new_n1323__spl_;
  wire new_n1320__spl_;
  wire new_n1325__spl_;
  wire new_n1326__spl_;
  wire new_n1319__spl_;
  wire new_n1328__spl_;
  wire new_n1329__spl_;
  wire new_n1318__spl_;
  wire new_n1331__spl_;
  wire new_n1332__spl_;
  wire new_n1317__spl_;
  wire new_n1334__spl_;
  wire new_n1335__spl_;
  wire new_n1316__spl_;
  wire new_n1337__spl_;
  wire new_n1338__spl_;
  wire new_n1315__spl_;
  wire new_n1340__spl_;
  wire new_n1341__spl_;
  wire new_n1314__spl_;
  wire new_n1343__spl_;
  wire new_n1344__spl_;
  wire new_n1313__spl_;
  wire new_n1346__spl_;
  wire new_n1347__spl_;
  wire new_n1312__spl_;
  wire new_n1349__spl_;
  wire new_n1350__spl_;
  wire new_n1311__spl_;
  wire new_n1352__spl_;
  wire new_n1353__spl_;
  wire new_n1310__spl_;
  wire new_n1355__spl_;
  wire new_n1356__spl_;
  wire new_n1309__spl_;
  wire new_n1358__spl_;
  wire new_n1359__spl_;
  wire new_n1308__spl_;
  wire new_n1361__spl_;
  wire new_n1362__spl_;
  wire new_n1307__spl_;
  wire new_n1364__spl_;
  wire new_n1365__spl_;
  wire new_n1306__spl_;
  wire new_n1367__spl_;
  wire new_n1368__spl_;
  wire new_n1305__spl_;
  wire new_n1370__spl_;
  wire new_n1371__spl_;
  wire new_n1304__spl_;
  wire new_n1373__spl_;
  wire new_n1374__spl_;
  wire new_n1303__spl_;
  wire new_n1376__spl_;
  wire new_n1377__spl_;
  wire new_n1302__spl_;
  wire new_n1379__spl_;
  wire new_n1380__spl_;
  wire new_n1301__spl_;
  wire new_n1382__spl_;
  wire new_n1383__spl_;
  wire new_n1300__spl_;
  wire new_n1385__spl_;
  wire new_n1386__spl_;
  wire new_n1299__spl_;
  wire new_n1388__spl_;
  wire new_n1389__spl_;
  wire new_n1298__spl_;
  wire new_n1391__spl_;
  wire new_n1392__spl_;
  wire new_n1416__spl_;
  wire new_n1417__spl_;
  wire new_n1418__spl_;
  wire new_n1415__spl_;
  wire new_n1420__spl_;
  wire new_n1421__spl_;
  wire new_n1414__spl_;
  wire new_n1423__spl_;
  wire new_n1424__spl_;
  wire new_n1413__spl_;
  wire new_n1426__spl_;
  wire new_n1427__spl_;
  wire new_n1412__spl_;
  wire new_n1429__spl_;
  wire new_n1430__spl_;
  wire new_n1411__spl_;
  wire new_n1432__spl_;
  wire new_n1433__spl_;
  wire new_n1410__spl_;
  wire new_n1435__spl_;
  wire new_n1436__spl_;
  wire new_n1409__spl_;
  wire new_n1438__spl_;
  wire new_n1439__spl_;
  wire new_n1408__spl_;
  wire new_n1441__spl_;
  wire new_n1442__spl_;
  wire new_n1407__spl_;
  wire new_n1444__spl_;
  wire new_n1445__spl_;
  wire new_n1406__spl_;
  wire new_n1447__spl_;
  wire new_n1448__spl_;
  wire new_n1405__spl_;
  wire new_n1450__spl_;
  wire new_n1451__spl_;
  wire new_n1404__spl_;
  wire new_n1453__spl_;
  wire new_n1454__spl_;
  wire new_n1403__spl_;
  wire new_n1456__spl_;
  wire new_n1457__spl_;
  wire new_n1402__spl_;
  wire new_n1459__spl_;
  wire new_n1460__spl_;
  wire new_n1401__spl_;
  wire new_n1462__spl_;
  wire new_n1463__spl_;
  wire new_n1400__spl_;
  wire new_n1465__spl_;
  wire new_n1466__spl_;
  wire new_n1399__spl_;
  wire new_n1468__spl_;
  wire new_n1469__spl_;
  wire new_n1398__spl_;
  wire new_n1471__spl_;
  wire new_n1472__spl_;
  wire new_n1397__spl_;
  wire new_n1474__spl_;
  wire new_n1475__spl_;
  wire new_n1396__spl_;
  wire new_n1477__spl_;
  wire new_n1478__spl_;
  wire new_n1395__spl_;
  wire new_n1480__spl_;
  wire new_n1481__spl_;
  wire new_n1503__spl_;
  wire new_n1504__spl_;
  wire new_n1505__spl_;
  wire new_n1502__spl_;
  wire new_n1507__spl_;
  wire new_n1508__spl_;
  wire new_n1501__spl_;
  wire new_n1510__spl_;
  wire new_n1511__spl_;
  wire new_n1500__spl_;
  wire new_n1513__spl_;
  wire new_n1514__spl_;
  wire new_n1499__spl_;
  wire new_n1516__spl_;
  wire new_n1517__spl_;
  wire new_n1498__spl_;
  wire new_n1519__spl_;
  wire new_n1520__spl_;
  wire new_n1497__spl_;
  wire new_n1522__spl_;
  wire new_n1523__spl_;
  wire new_n1496__spl_;
  wire new_n1525__spl_;
  wire new_n1526__spl_;
  wire new_n1495__spl_;
  wire new_n1528__spl_;
  wire new_n1529__spl_;
  wire new_n1494__spl_;
  wire new_n1531__spl_;
  wire new_n1532__spl_;
  wire new_n1493__spl_;
  wire new_n1534__spl_;
  wire new_n1535__spl_;
  wire new_n1492__spl_;
  wire new_n1537__spl_;
  wire new_n1538__spl_;
  wire new_n1491__spl_;
  wire new_n1540__spl_;
  wire new_n1541__spl_;
  wire new_n1490__spl_;
  wire new_n1543__spl_;
  wire new_n1544__spl_;
  wire new_n1489__spl_;
  wire new_n1546__spl_;
  wire new_n1547__spl_;
  wire new_n1488__spl_;
  wire new_n1549__spl_;
  wire new_n1550__spl_;
  wire new_n1487__spl_;
  wire new_n1552__spl_;
  wire new_n1553__spl_;
  wire new_n1486__spl_;
  wire new_n1555__spl_;
  wire new_n1556__spl_;
  wire new_n1485__spl_;
  wire new_n1558__spl_;
  wire new_n1559__spl_;
  wire new_n1484__spl_;
  wire new_n1561__spl_;
  wire new_n1562__spl_;
  wire new_n1582__spl_;
  wire new_n1583__spl_;
  wire new_n1584__spl_;
  wire new_n1581__spl_;
  wire new_n1586__spl_;
  wire new_n1587__spl_;
  wire new_n1580__spl_;
  wire new_n1589__spl_;
  wire new_n1590__spl_;
  wire new_n1579__spl_;
  wire new_n1592__spl_;
  wire new_n1593__spl_;
  wire new_n1578__spl_;
  wire new_n1595__spl_;
  wire new_n1596__spl_;
  wire new_n1577__spl_;
  wire new_n1598__spl_;
  wire new_n1599__spl_;
  wire new_n1576__spl_;
  wire new_n1601__spl_;
  wire new_n1602__spl_;
  wire new_n1575__spl_;
  wire new_n1604__spl_;
  wire new_n1605__spl_;
  wire new_n1574__spl_;
  wire new_n1607__spl_;
  wire new_n1608__spl_;
  wire new_n1573__spl_;
  wire new_n1610__spl_;
  wire new_n1611__spl_;
  wire new_n1572__spl_;
  wire new_n1613__spl_;
  wire new_n1614__spl_;
  wire new_n1571__spl_;
  wire new_n1616__spl_;
  wire new_n1617__spl_;
  wire new_n1570__spl_;
  wire new_n1619__spl_;
  wire new_n1620__spl_;
  wire new_n1569__spl_;
  wire new_n1622__spl_;
  wire new_n1623__spl_;
  wire new_n1568__spl_;
  wire new_n1625__spl_;
  wire new_n1626__spl_;
  wire new_n1567__spl_;
  wire new_n1628__spl_;
  wire new_n1629__spl_;
  wire new_n1566__spl_;
  wire new_n1631__spl_;
  wire new_n1632__spl_;
  wire new_n1565__spl_;
  wire new_n1634__spl_;
  wire new_n1635__spl_;
  wire new_n1653__spl_;
  wire new_n1654__spl_;
  wire new_n1655__spl_;
  wire new_n1652__spl_;
  wire new_n1657__spl_;
  wire new_n1658__spl_;
  wire new_n1651__spl_;
  wire new_n1660__spl_;
  wire new_n1661__spl_;
  wire new_n1650__spl_;
  wire new_n1663__spl_;
  wire new_n1664__spl_;
  wire new_n1649__spl_;
  wire new_n1666__spl_;
  wire new_n1667__spl_;
  wire new_n1648__spl_;
  wire new_n1669__spl_;
  wire new_n1670__spl_;
  wire new_n1647__spl_;
  wire new_n1672__spl_;
  wire new_n1673__spl_;
  wire new_n1646__spl_;
  wire new_n1675__spl_;
  wire new_n1676__spl_;
  wire new_n1645__spl_;
  wire new_n1678__spl_;
  wire new_n1679__spl_;
  wire new_n1644__spl_;
  wire new_n1681__spl_;
  wire new_n1682__spl_;
  wire new_n1643__spl_;
  wire new_n1684__spl_;
  wire new_n1685__spl_;
  wire new_n1642__spl_;
  wire new_n1687__spl_;
  wire new_n1688__spl_;
  wire new_n1641__spl_;
  wire new_n1690__spl_;
  wire new_n1691__spl_;
  wire new_n1640__spl_;
  wire new_n1693__spl_;
  wire new_n1694__spl_;
  wire new_n1639__spl_;
  wire new_n1696__spl_;
  wire new_n1697__spl_;
  wire new_n1638__spl_;
  wire new_n1699__spl_;
  wire new_n1700__spl_;
  wire new_n1716__spl_;
  wire new_n1717__spl_;
  wire new_n1718__spl_;
  wire new_n1715__spl_;
  wire new_n1720__spl_;
  wire new_n1721__spl_;
  wire new_n1714__spl_;
  wire new_n1723__spl_;
  wire new_n1724__spl_;
  wire new_n1713__spl_;
  wire new_n1726__spl_;
  wire new_n1727__spl_;
  wire new_n1712__spl_;
  wire new_n1729__spl_;
  wire new_n1730__spl_;
  wire new_n1711__spl_;
  wire new_n1732__spl_;
  wire new_n1733__spl_;
  wire new_n1710__spl_;
  wire new_n1735__spl_;
  wire new_n1736__spl_;
  wire new_n1709__spl_;
  wire new_n1738__spl_;
  wire new_n1739__spl_;
  wire new_n1708__spl_;
  wire new_n1741__spl_;
  wire new_n1742__spl_;
  wire new_n1707__spl_;
  wire new_n1744__spl_;
  wire new_n1745__spl_;
  wire new_n1706__spl_;
  wire new_n1747__spl_;
  wire new_n1748__spl_;
  wire new_n1705__spl_;
  wire new_n1750__spl_;
  wire new_n1751__spl_;
  wire new_n1704__spl_;
  wire new_n1753__spl_;
  wire new_n1754__spl_;
  wire new_n1703__spl_;
  wire new_n1756__spl_;
  wire new_n1757__spl_;
  wire new_n1771__spl_;
  wire new_n1772__spl_;
  wire new_n1773__spl_;
  wire new_n1770__spl_;
  wire new_n1775__spl_;
  wire new_n1776__spl_;
  wire new_n1769__spl_;
  wire new_n1778__spl_;
  wire new_n1779__spl_;
  wire new_n1768__spl_;
  wire new_n1781__spl_;
  wire new_n1782__spl_;
  wire new_n1767__spl_;
  wire new_n1784__spl_;
  wire new_n1785__spl_;
  wire new_n1766__spl_;
  wire new_n1787__spl_;
  wire new_n1788__spl_;
  wire new_n1765__spl_;
  wire new_n1790__spl_;
  wire new_n1791__spl_;
  wire new_n1764__spl_;
  wire new_n1793__spl_;
  wire new_n1794__spl_;
  wire new_n1763__spl_;
  wire new_n1796__spl_;
  wire new_n1797__spl_;
  wire new_n1762__spl_;
  wire new_n1799__spl_;
  wire new_n1800__spl_;
  wire new_n1761__spl_;
  wire new_n1802__spl_;
  wire new_n1803__spl_;
  wire new_n1760__spl_;
  wire new_n1805__spl_;
  wire new_n1806__spl_;
  wire new_n1818__spl_;
  wire new_n1819__spl_;
  wire new_n1820__spl_;
  wire new_n1817__spl_;
  wire new_n1822__spl_;
  wire new_n1823__spl_;
  wire new_n1816__spl_;
  wire new_n1825__spl_;
  wire new_n1826__spl_;
  wire new_n1815__spl_;
  wire new_n1828__spl_;
  wire new_n1829__spl_;
  wire new_n1814__spl_;
  wire new_n1831__spl_;
  wire new_n1832__spl_;
  wire new_n1813__spl_;
  wire new_n1834__spl_;
  wire new_n1835__spl_;
  wire new_n1812__spl_;
  wire new_n1837__spl_;
  wire new_n1838__spl_;
  wire new_n1811__spl_;
  wire new_n1840__spl_;
  wire new_n1841__spl_;
  wire new_n1810__spl_;
  wire new_n1843__spl_;
  wire new_n1844__spl_;
  wire new_n1809__spl_;
  wire new_n1846__spl_;
  wire new_n1847__spl_;
  wire new_n1857__spl_;
  wire new_n1858__spl_;
  wire new_n1859__spl_;
  wire new_n1856__spl_;
  wire new_n1861__spl_;
  wire new_n1862__spl_;
  wire new_n1855__spl_;
  wire new_n1864__spl_;
  wire new_n1865__spl_;
  wire new_n1854__spl_;
  wire new_n1867__spl_;
  wire new_n1868__spl_;
  wire new_n1853__spl_;
  wire new_n1870__spl_;
  wire new_n1871__spl_;
  wire new_n1852__spl_;
  wire new_n1873__spl_;
  wire new_n1874__spl_;
  wire new_n1851__spl_;
  wire new_n1876__spl_;
  wire new_n1877__spl_;
  wire new_n1850__spl_;
  wire new_n1879__spl_;
  wire new_n1880__spl_;
  wire new_n1888__spl_;
  wire new_n1889__spl_;
  wire new_n1890__spl_;
  wire new_n1887__spl_;
  wire new_n1892__spl_;
  wire new_n1893__spl_;
  wire new_n1886__spl_;
  wire new_n1895__spl_;
  wire new_n1896__spl_;
  wire new_n1885__spl_;
  wire new_n1898__spl_;
  wire new_n1899__spl_;
  wire new_n1884__spl_;
  wire new_n1901__spl_;
  wire new_n1902__spl_;
  wire new_n1883__spl_;
  wire new_n1904__spl_;
  wire new_n1905__spl_;
  wire new_n1911__spl_;
  wire new_n1912__spl_;
  wire new_n1913__spl_;
  wire new_n1910__spl_;
  wire new_n1915__spl_;
  wire new_n1916__spl_;
  wire new_n1909__spl_;
  wire new_n1918__spl_;
  wire new_n1919__spl_;
  wire new_n1908__spl_;
  wire new_n1921__spl_;
  wire new_n1922__spl_;
  wire new_n1925__spl_;
  wire new_n1926__spl_;
  wire new_n1927__spl_;
  wire new_n1928__spl_;
  wire new_n1930__spl_;
  wire new_n1931__spl_;

  and1
  g0000
  (
    .dina(G1_spl_000),
    .dinb(G17_spl_000),
    .dout(G6257)
  );


  nor2
  g0001
  (
    .dina(G2_spl_000),
    .dinb(G17_spl_000),
    .dout(new_n66_)
  );


  and1
  g0002
  (
    .dina(G1_spl_000),
    .dinb(G18_spl_000),
    .dout(new_n67_)
  );


  anb2
  g0003
  (
    .dina(new_n66__spl_),
    .dinb(new_n67__spl_),
    .dout(new_n68_)
  );


  anb1
  g0004
  (
    .dina(new_n66__spl_),
    .dinb(new_n67__spl_),
    .dout(new_n69_)
  );


  anb1
  g0005
  (
    .dina(new_n68__spl_0),
    .dinb(new_n69_),
    .dout(G6258)
  );


  nor2
  g0006
  (
    .dina(G1_spl_001),
    .dinb(G19_spl_000),
    .dout(new_n71_)
  );


  nor2
  g0007
  (
    .dina(G3_spl_000),
    .dinb(G17_spl_001),
    .dout(new_n72_)
  );


  and1
  g0008
  (
    .dina(G2_spl_000),
    .dinb(G18_spl_000),
    .dout(new_n73_)
  );


  anb2
  g0009
  (
    .dina(new_n72__spl_),
    .dinb(new_n73__spl_),
    .dout(new_n74_)
  );


  anb1
  g0010
  (
    .dina(new_n72__spl_),
    .dinb(new_n73__spl_),
    .dout(new_n75_)
  );


  anb1
  g0011
  (
    .dina(new_n74__spl_0),
    .dinb(new_n75_),
    .dout(new_n76_)
  );


  anb1
  g0012
  (
    .dina(new_n68__spl_0),
    .dinb(new_n76__spl_),
    .dout(new_n77_)
  );


  anb2
  g0013
  (
    .dina(new_n68__spl_),
    .dinb(new_n76__spl_),
    .dout(new_n78_)
  );


  anb2
  g0014
  (
    .dina(new_n77__spl_),
    .dinb(new_n78_),
    .dout(new_n79_)
  );


  anb1
  g0015
  (
    .dina(new_n71__spl_),
    .dinb(new_n79__spl_),
    .dout(new_n80_)
  );


  anb2
  g0016
  (
    .dina(new_n71__spl_),
    .dinb(new_n79__spl_),
    .dout(new_n81_)
  );


  anb2
  g0017
  (
    .dina(new_n80__spl_),
    .dinb(new_n81_),
    .dout(G6259)
  );


  nor2
  g0018
  (
    .dina(G1_spl_001),
    .dinb(G20_spl_000),
    .dout(new_n83_)
  );


  and2
  g0019
  (
    .dina(new_n77__spl_),
    .dinb(new_n80__spl_),
    .dout(new_n84_)
  );


  nor2
  g0020
  (
    .dina(G2_spl_001),
    .dinb(G19_spl_000),
    .dout(new_n85_)
  );


  nor2
  g0021
  (
    .dina(G4_spl_000),
    .dinb(G17_spl_001),
    .dout(new_n86_)
  );


  and1
  g0022
  (
    .dina(G3_spl_000),
    .dinb(G18_spl_001),
    .dout(new_n87_)
  );


  anb2
  g0023
  (
    .dina(new_n86__spl_),
    .dinb(new_n87__spl_),
    .dout(new_n88_)
  );


  anb1
  g0024
  (
    .dina(new_n86__spl_),
    .dinb(new_n87__spl_),
    .dout(new_n89_)
  );


  anb1
  g0025
  (
    .dina(new_n88__spl_0),
    .dinb(new_n89_),
    .dout(new_n90_)
  );


  anb1
  g0026
  (
    .dina(new_n74__spl_0),
    .dinb(new_n90__spl_),
    .dout(new_n91_)
  );


  anb2
  g0027
  (
    .dina(new_n74__spl_),
    .dinb(new_n90__spl_),
    .dout(new_n92_)
  );


  anb2
  g0028
  (
    .dina(new_n91__spl_),
    .dinb(new_n92_),
    .dout(new_n93_)
  );


  anb1
  g0029
  (
    .dina(new_n85__spl_),
    .dinb(new_n93__spl_),
    .dout(new_n94_)
  );


  anb2
  g0030
  (
    .dina(new_n85__spl_),
    .dinb(new_n93__spl_),
    .dout(new_n95_)
  );


  anb2
  g0031
  (
    .dina(new_n94__spl_),
    .dinb(new_n95_),
    .dout(new_n96_)
  );


  anb1
  g0032
  (
    .dina(new_n84__spl_),
    .dinb(new_n96__spl_),
    .dout(new_n97_)
  );


  anb2
  g0033
  (
    .dina(new_n84__spl_),
    .dinb(new_n96__spl_),
    .dout(new_n98_)
  );


  anb2
  g0034
  (
    .dina(new_n97__spl_),
    .dinb(new_n98_),
    .dout(new_n99_)
  );


  anb1
  g0035
  (
    .dina(new_n83__spl_),
    .dinb(new_n99__spl_),
    .dout(new_n100_)
  );


  anb2
  g0036
  (
    .dina(new_n83__spl_),
    .dinb(new_n99__spl_),
    .dout(new_n101_)
  );


  anb2
  g0037
  (
    .dina(new_n100__spl_),
    .dinb(new_n101_),
    .dout(G6260)
  );


  nor2
  g0038
  (
    .dina(G1_spl_010),
    .dinb(G21_spl_000),
    .dout(new_n103_)
  );


  and2
  g0039
  (
    .dina(new_n97__spl_),
    .dinb(new_n100__spl_),
    .dout(new_n104_)
  );


  nor2
  g0040
  (
    .dina(G2_spl_001),
    .dinb(G20_spl_000),
    .dout(new_n105_)
  );


  and2
  g0041
  (
    .dina(new_n91__spl_),
    .dinb(new_n94__spl_),
    .dout(new_n106_)
  );


  nor2
  g0042
  (
    .dina(G3_spl_001),
    .dinb(G19_spl_001),
    .dout(new_n107_)
  );


  and1
  g0043
  (
    .dina(G5_spl_000),
    .dinb(G17_spl_010),
    .dout(new_n108_)
  );


  nor2
  g0044
  (
    .dina(G4_spl_000),
    .dinb(G18_spl_001),
    .dout(new_n109_)
  );


  anb1
  g0045
  (
    .dina(new_n108__spl_),
    .dinb(new_n109__spl_),
    .dout(new_n110_)
  );


  anb2
  g0046
  (
    .dina(new_n108__spl_),
    .dinb(new_n109__spl_),
    .dout(new_n111_)
  );


  nab1
  g0047
  (
    .dina(new_n110__spl_0),
    .dinb(new_n111_),
    .dout(new_n112_)
  );


  anb1
  g0048
  (
    .dina(new_n88__spl_0),
    .dinb(new_n112__spl_),
    .dout(new_n113_)
  );


  anb2
  g0049
  (
    .dina(new_n88__spl_),
    .dinb(new_n112__spl_),
    .dout(new_n114_)
  );


  anb2
  g0050
  (
    .dina(new_n113__spl_),
    .dinb(new_n114_),
    .dout(new_n115_)
  );


  anb1
  g0051
  (
    .dina(new_n107__spl_),
    .dinb(new_n115__spl_),
    .dout(new_n116_)
  );


  anb2
  g0052
  (
    .dina(new_n107__spl_),
    .dinb(new_n115__spl_),
    .dout(new_n117_)
  );


  anb2
  g0053
  (
    .dina(new_n116__spl_),
    .dinb(new_n117_),
    .dout(new_n118_)
  );


  anb1
  g0054
  (
    .dina(new_n106__spl_),
    .dinb(new_n118__spl_),
    .dout(new_n119_)
  );


  anb2
  g0055
  (
    .dina(new_n106__spl_),
    .dinb(new_n118__spl_),
    .dout(new_n120_)
  );


  anb2
  g0056
  (
    .dina(new_n119__spl_),
    .dinb(new_n120_),
    .dout(new_n121_)
  );


  anb1
  g0057
  (
    .dina(new_n105__spl_),
    .dinb(new_n121__spl_),
    .dout(new_n122_)
  );


  anb2
  g0058
  (
    .dina(new_n105__spl_),
    .dinb(new_n121__spl_),
    .dout(new_n123_)
  );


  anb2
  g0059
  (
    .dina(new_n122__spl_),
    .dinb(new_n123_),
    .dout(new_n124_)
  );


  anb1
  g0060
  (
    .dina(new_n104__spl_),
    .dinb(new_n124__spl_),
    .dout(new_n125_)
  );


  anb2
  g0061
  (
    .dina(new_n104__spl_),
    .dinb(new_n124__spl_),
    .dout(new_n126_)
  );


  anb2
  g0062
  (
    .dina(new_n125__spl_),
    .dinb(new_n126_),
    .dout(new_n127_)
  );


  anb1
  g0063
  (
    .dina(new_n103__spl_),
    .dinb(new_n127__spl_),
    .dout(new_n128_)
  );


  anb2
  g0064
  (
    .dina(new_n103__spl_),
    .dinb(new_n127__spl_),
    .dout(new_n129_)
  );


  anb2
  g0065
  (
    .dina(new_n128__spl_),
    .dinb(new_n129_),
    .dout(G6261)
  );


  nor2
  g0066
  (
    .dina(G1_spl_010),
    .dinb(G22_spl_000),
    .dout(new_n131_)
  );


  and2
  g0067
  (
    .dina(new_n125__spl_),
    .dinb(new_n128__spl_),
    .dout(new_n132_)
  );


  nor2
  g0068
  (
    .dina(G2_spl_010),
    .dinb(G21_spl_000),
    .dout(new_n133_)
  );


  and2
  g0069
  (
    .dina(new_n119__spl_),
    .dinb(new_n122__spl_),
    .dout(new_n134_)
  );


  nor2
  g0070
  (
    .dina(G3_spl_001),
    .dinb(G20_spl_001),
    .dout(new_n135_)
  );


  and2
  g0071
  (
    .dina(new_n113__spl_),
    .dinb(new_n116__spl_),
    .dout(new_n136_)
  );


  nor2
  g0072
  (
    .dina(G4_spl_001),
    .dinb(G19_spl_001),
    .dout(new_n137_)
  );


  nor2
  g0073
  (
    .dina(G6_spl_000),
    .dinb(G17_spl_010),
    .dout(new_n138_)
  );


  and1
  g0074
  (
    .dina(G5_spl_000),
    .dinb(G18_spl_010),
    .dout(new_n139_)
  );


  anb2
  g0075
  (
    .dina(new_n138__spl_),
    .dinb(new_n139__spl_),
    .dout(new_n140_)
  );


  anb1
  g0076
  (
    .dina(new_n138__spl_),
    .dinb(new_n139__spl_),
    .dout(new_n141_)
  );


  nab2
  g0077
  (
    .dina(new_n140__spl_0),
    .dinb(new_n141_),
    .dout(new_n142_)
  );


  anb2
  g0078
  (
    .dina(new_n110__spl_0),
    .dinb(new_n142__spl_),
    .dout(new_n143_)
  );


  anb1
  g0079
  (
    .dina(new_n110__spl_),
    .dinb(new_n142__spl_),
    .dout(new_n144_)
  );


  nab2
  g0080
  (
    .dina(new_n143__spl_),
    .dinb(new_n144_),
    .dout(new_n145_)
  );


  anb1
  g0081
  (
    .dina(new_n137__spl_),
    .dinb(new_n145__spl_),
    .dout(new_n146_)
  );


  anb2
  g0082
  (
    .dina(new_n137__spl_),
    .dinb(new_n145__spl_),
    .dout(new_n147_)
  );


  anb2
  g0083
  (
    .dina(new_n146__spl_),
    .dinb(new_n147_),
    .dout(new_n148_)
  );


  anb1
  g0084
  (
    .dina(new_n136__spl_),
    .dinb(new_n148__spl_),
    .dout(new_n149_)
  );


  anb2
  g0085
  (
    .dina(new_n136__spl_),
    .dinb(new_n148__spl_),
    .dout(new_n150_)
  );


  anb2
  g0086
  (
    .dina(new_n149__spl_),
    .dinb(new_n150_),
    .dout(new_n151_)
  );


  anb1
  g0087
  (
    .dina(new_n135__spl_),
    .dinb(new_n151__spl_),
    .dout(new_n152_)
  );


  anb2
  g0088
  (
    .dina(new_n135__spl_),
    .dinb(new_n151__spl_),
    .dout(new_n153_)
  );


  anb2
  g0089
  (
    .dina(new_n152__spl_),
    .dinb(new_n153_),
    .dout(new_n154_)
  );


  anb1
  g0090
  (
    .dina(new_n134__spl_),
    .dinb(new_n154__spl_),
    .dout(new_n155_)
  );


  anb2
  g0091
  (
    .dina(new_n134__spl_),
    .dinb(new_n154__spl_),
    .dout(new_n156_)
  );


  anb2
  g0092
  (
    .dina(new_n155__spl_),
    .dinb(new_n156_),
    .dout(new_n157_)
  );


  anb1
  g0093
  (
    .dina(new_n133__spl_),
    .dinb(new_n157__spl_),
    .dout(new_n158_)
  );


  anb2
  g0094
  (
    .dina(new_n133__spl_),
    .dinb(new_n157__spl_),
    .dout(new_n159_)
  );


  anb2
  g0095
  (
    .dina(new_n158__spl_),
    .dinb(new_n159_),
    .dout(new_n160_)
  );


  anb1
  g0096
  (
    .dina(new_n132__spl_),
    .dinb(new_n160__spl_),
    .dout(new_n161_)
  );


  anb2
  g0097
  (
    .dina(new_n132__spl_),
    .dinb(new_n160__spl_),
    .dout(new_n162_)
  );


  anb2
  g0098
  (
    .dina(new_n161__spl_),
    .dinb(new_n162_),
    .dout(new_n163_)
  );


  anb1
  g0099
  (
    .dina(new_n131__spl_),
    .dinb(new_n163__spl_),
    .dout(new_n164_)
  );


  anb2
  g0100
  (
    .dina(new_n131__spl_),
    .dinb(new_n163__spl_),
    .dout(new_n165_)
  );


  anb2
  g0101
  (
    .dina(new_n164__spl_),
    .dinb(new_n165_),
    .dout(G6262)
  );


  nor2
  g0102
  (
    .dina(G1_spl_011),
    .dinb(G23_spl_000),
    .dout(new_n167_)
  );


  and2
  g0103
  (
    .dina(new_n161__spl_),
    .dinb(new_n164__spl_),
    .dout(new_n168_)
  );


  nor2
  g0104
  (
    .dina(G2_spl_010),
    .dinb(G22_spl_000),
    .dout(new_n169_)
  );


  and2
  g0105
  (
    .dina(new_n155__spl_),
    .dinb(new_n158__spl_),
    .dout(new_n170_)
  );


  nor2
  g0106
  (
    .dina(G3_spl_010),
    .dinb(G21_spl_001),
    .dout(new_n171_)
  );


  and2
  g0107
  (
    .dina(new_n149__spl_),
    .dinb(new_n152__spl_),
    .dout(new_n172_)
  );


  nor2
  g0108
  (
    .dina(G4_spl_001),
    .dinb(G20_spl_001),
    .dout(new_n173_)
  );


  anb1
  g0109
  (
    .dina(new_n143__spl_),
    .dinb(new_n146__spl_),
    .dout(new_n174_)
  );


  and1
  g0110
  (
    .dina(G5_spl_001),
    .dinb(G19_spl_010),
    .dout(new_n175_)
  );


  nor2
  g0111
  (
    .dina(G7_spl_000),
    .dinb(G17_spl_011),
    .dout(new_n176_)
  );


  and1
  g0112
  (
    .dina(G6_spl_000),
    .dinb(G18_spl_010),
    .dout(new_n177_)
  );


  anb2
  g0113
  (
    .dina(new_n176__spl_),
    .dinb(new_n177__spl_),
    .dout(new_n178_)
  );


  anb1
  g0114
  (
    .dina(new_n176__spl_),
    .dinb(new_n177__spl_),
    .dout(new_n179_)
  );


  anb1
  g0115
  (
    .dina(new_n178__spl_0),
    .dinb(new_n179_),
    .dout(new_n180_)
  );


  anb1
  g0116
  (
    .dina(new_n140__spl_0),
    .dinb(new_n180__spl_),
    .dout(new_n181_)
  );


  anb2
  g0117
  (
    .dina(new_n140__spl_),
    .dinb(new_n180__spl_),
    .dout(new_n182_)
  );


  nab1
  g0118
  (
    .dina(new_n181__spl_),
    .dinb(new_n182_),
    .dout(new_n183_)
  );


  anb2
  g0119
  (
    .dina(new_n175__spl_),
    .dinb(new_n183__spl_),
    .dout(new_n184_)
  );


  anb1
  g0120
  (
    .dina(new_n175__spl_),
    .dinb(new_n183__spl_),
    .dout(new_n185_)
  );


  anb1
  g0121
  (
    .dina(new_n184__spl_),
    .dinb(new_n185_),
    .dout(new_n186_)
  );


  anb2
  g0122
  (
    .dina(new_n174__spl_),
    .dinb(new_n186__spl_),
    .dout(new_n187_)
  );


  anb1
  g0123
  (
    .dina(new_n174__spl_),
    .dinb(new_n186__spl_),
    .dout(new_n188_)
  );


  nab2
  g0124
  (
    .dina(new_n187__spl_),
    .dinb(new_n188_),
    .dout(new_n189_)
  );


  anb1
  g0125
  (
    .dina(new_n173__spl_),
    .dinb(new_n189__spl_),
    .dout(new_n190_)
  );


  anb2
  g0126
  (
    .dina(new_n173__spl_),
    .dinb(new_n189__spl_),
    .dout(new_n191_)
  );


  anb2
  g0127
  (
    .dina(new_n190__spl_),
    .dinb(new_n191_),
    .dout(new_n192_)
  );


  anb1
  g0128
  (
    .dina(new_n172__spl_),
    .dinb(new_n192__spl_),
    .dout(new_n193_)
  );


  anb2
  g0129
  (
    .dina(new_n172__spl_),
    .dinb(new_n192__spl_),
    .dout(new_n194_)
  );


  anb2
  g0130
  (
    .dina(new_n193__spl_),
    .dinb(new_n194_),
    .dout(new_n195_)
  );


  anb1
  g0131
  (
    .dina(new_n171__spl_),
    .dinb(new_n195__spl_),
    .dout(new_n196_)
  );


  anb2
  g0132
  (
    .dina(new_n171__spl_),
    .dinb(new_n195__spl_),
    .dout(new_n197_)
  );


  anb2
  g0133
  (
    .dina(new_n196__spl_),
    .dinb(new_n197_),
    .dout(new_n198_)
  );


  anb1
  g0134
  (
    .dina(new_n170__spl_),
    .dinb(new_n198__spl_),
    .dout(new_n199_)
  );


  anb2
  g0135
  (
    .dina(new_n170__spl_),
    .dinb(new_n198__spl_),
    .dout(new_n200_)
  );


  anb2
  g0136
  (
    .dina(new_n199__spl_),
    .dinb(new_n200_),
    .dout(new_n201_)
  );


  anb1
  g0137
  (
    .dina(new_n169__spl_),
    .dinb(new_n201__spl_),
    .dout(new_n202_)
  );


  anb2
  g0138
  (
    .dina(new_n169__spl_),
    .dinb(new_n201__spl_),
    .dout(new_n203_)
  );


  anb2
  g0139
  (
    .dina(new_n202__spl_),
    .dinb(new_n203_),
    .dout(new_n204_)
  );


  anb1
  g0140
  (
    .dina(new_n168__spl_),
    .dinb(new_n204__spl_),
    .dout(new_n205_)
  );


  anb2
  g0141
  (
    .dina(new_n168__spl_),
    .dinb(new_n204__spl_),
    .dout(new_n206_)
  );


  anb2
  g0142
  (
    .dina(new_n205__spl_),
    .dinb(new_n206_),
    .dout(new_n207_)
  );


  anb1
  g0143
  (
    .dina(new_n167__spl_),
    .dinb(new_n207__spl_),
    .dout(new_n208_)
  );


  anb2
  g0144
  (
    .dina(new_n167__spl_),
    .dinb(new_n207__spl_),
    .dout(new_n209_)
  );


  anb2
  g0145
  (
    .dina(new_n208__spl_),
    .dinb(new_n209_),
    .dout(G6263)
  );


  nor2
  g0146
  (
    .dina(G1_spl_011),
    .dinb(G24_spl_000),
    .dout(new_n211_)
  );


  and2
  g0147
  (
    .dina(new_n205__spl_),
    .dinb(new_n208__spl_),
    .dout(new_n212_)
  );


  nor2
  g0148
  (
    .dina(G2_spl_011),
    .dinb(G23_spl_000),
    .dout(new_n213_)
  );


  and2
  g0149
  (
    .dina(new_n199__spl_),
    .dinb(new_n202__spl_),
    .dout(new_n214_)
  );


  nor2
  g0150
  (
    .dina(G3_spl_010),
    .dinb(G22_spl_001),
    .dout(new_n215_)
  );


  and2
  g0151
  (
    .dina(new_n193__spl_),
    .dinb(new_n196__spl_),
    .dout(new_n216_)
  );


  nor2
  g0152
  (
    .dina(G4_spl_010),
    .dinb(G21_spl_001),
    .dout(new_n217_)
  );


  anb1
  g0153
  (
    .dina(new_n187__spl_),
    .dinb(new_n190__spl_),
    .dout(new_n218_)
  );


  and1
  g0154
  (
    .dina(G5_spl_001),
    .dinb(G20_spl_010),
    .dout(new_n219_)
  );


  anb2
  g0155
  (
    .dina(new_n181__spl_),
    .dinb(new_n184__spl_),
    .dout(new_n220_)
  );


  and1
  g0156
  (
    .dina(G6_spl_001),
    .dinb(G19_spl_010),
    .dout(new_n221_)
  );


  nor2
  g0157
  (
    .dina(G8_spl_000),
    .dinb(G17_spl_011),
    .dout(new_n222_)
  );


  and1
  g0158
  (
    .dina(G7_spl_000),
    .dinb(G18_spl_011),
    .dout(new_n223_)
  );


  anb2
  g0159
  (
    .dina(new_n222__spl_),
    .dinb(new_n223__spl_),
    .dout(new_n224_)
  );


  anb1
  g0160
  (
    .dina(new_n222__spl_),
    .dinb(new_n223__spl_),
    .dout(new_n225_)
  );


  anb1
  g0161
  (
    .dina(new_n224__spl_0),
    .dinb(new_n225_),
    .dout(new_n226_)
  );


  anb1
  g0162
  (
    .dina(new_n178__spl_0),
    .dinb(new_n226__spl_),
    .dout(new_n227_)
  );


  anb2
  g0163
  (
    .dina(new_n178__spl_),
    .dinb(new_n226__spl_),
    .dout(new_n228_)
  );


  nab1
  g0164
  (
    .dina(new_n227__spl_),
    .dinb(new_n228_),
    .dout(new_n229_)
  );


  anb2
  g0165
  (
    .dina(new_n221__spl_),
    .dinb(new_n229__spl_),
    .dout(new_n230_)
  );


  anb1
  g0166
  (
    .dina(new_n221__spl_),
    .dinb(new_n229__spl_),
    .dout(new_n231_)
  );


  nab2
  g0167
  (
    .dina(new_n230__spl_),
    .dinb(new_n231_),
    .dout(new_n232_)
  );


  anb1
  g0168
  (
    .dina(new_n220__spl_),
    .dinb(new_n232__spl_),
    .dout(new_n233_)
  );


  anb2
  g0169
  (
    .dina(new_n220__spl_),
    .dinb(new_n232__spl_),
    .dout(new_n234_)
  );


  nab1
  g0170
  (
    .dina(new_n233__spl_),
    .dinb(new_n234_),
    .dout(new_n235_)
  );


  anb2
  g0171
  (
    .dina(new_n219__spl_),
    .dinb(new_n235__spl_),
    .dout(new_n236_)
  );


  anb1
  g0172
  (
    .dina(new_n219__spl_),
    .dinb(new_n235__spl_),
    .dout(new_n237_)
  );


  anb1
  g0173
  (
    .dina(new_n236__spl_),
    .dinb(new_n237_),
    .dout(new_n238_)
  );


  anb2
  g0174
  (
    .dina(new_n218__spl_),
    .dinb(new_n238__spl_),
    .dout(new_n239_)
  );


  anb1
  g0175
  (
    .dina(new_n218__spl_),
    .dinb(new_n238__spl_),
    .dout(new_n240_)
  );


  nab2
  g0176
  (
    .dina(new_n239__spl_),
    .dinb(new_n240_),
    .dout(new_n241_)
  );


  anb1
  g0177
  (
    .dina(new_n217__spl_),
    .dinb(new_n241__spl_),
    .dout(new_n242_)
  );


  anb2
  g0178
  (
    .dina(new_n217__spl_),
    .dinb(new_n241__spl_),
    .dout(new_n243_)
  );


  anb2
  g0179
  (
    .dina(new_n242__spl_),
    .dinb(new_n243_),
    .dout(new_n244_)
  );


  anb1
  g0180
  (
    .dina(new_n216__spl_),
    .dinb(new_n244__spl_),
    .dout(new_n245_)
  );


  anb2
  g0181
  (
    .dina(new_n216__spl_),
    .dinb(new_n244__spl_),
    .dout(new_n246_)
  );


  anb2
  g0182
  (
    .dina(new_n245__spl_),
    .dinb(new_n246_),
    .dout(new_n247_)
  );


  anb1
  g0183
  (
    .dina(new_n215__spl_),
    .dinb(new_n247__spl_),
    .dout(new_n248_)
  );


  anb2
  g0184
  (
    .dina(new_n215__spl_),
    .dinb(new_n247__spl_),
    .dout(new_n249_)
  );


  anb2
  g0185
  (
    .dina(new_n248__spl_),
    .dinb(new_n249_),
    .dout(new_n250_)
  );


  anb1
  g0186
  (
    .dina(new_n214__spl_),
    .dinb(new_n250__spl_),
    .dout(new_n251_)
  );


  anb2
  g0187
  (
    .dina(new_n214__spl_),
    .dinb(new_n250__spl_),
    .dout(new_n252_)
  );


  anb2
  g0188
  (
    .dina(new_n251__spl_),
    .dinb(new_n252_),
    .dout(new_n253_)
  );


  anb1
  g0189
  (
    .dina(new_n213__spl_),
    .dinb(new_n253__spl_),
    .dout(new_n254_)
  );


  anb2
  g0190
  (
    .dina(new_n213__spl_),
    .dinb(new_n253__spl_),
    .dout(new_n255_)
  );


  anb2
  g0191
  (
    .dina(new_n254__spl_),
    .dinb(new_n255_),
    .dout(new_n256_)
  );


  anb1
  g0192
  (
    .dina(new_n212__spl_),
    .dinb(new_n256__spl_),
    .dout(new_n257_)
  );


  anb2
  g0193
  (
    .dina(new_n212__spl_),
    .dinb(new_n256__spl_),
    .dout(new_n258_)
  );


  anb2
  g0194
  (
    .dina(new_n257__spl_),
    .dinb(new_n258_),
    .dout(new_n259_)
  );


  anb1
  g0195
  (
    .dina(new_n211__spl_),
    .dinb(new_n259__spl_),
    .dout(new_n260_)
  );


  anb2
  g0196
  (
    .dina(new_n211__spl_),
    .dinb(new_n259__spl_),
    .dout(new_n261_)
  );


  anb2
  g0197
  (
    .dina(new_n260__spl_),
    .dinb(new_n261_),
    .dout(G6264)
  );


  nor2
  g0198
  (
    .dina(G1_spl_100),
    .dinb(G25_spl_000),
    .dout(new_n263_)
  );


  and2
  g0199
  (
    .dina(new_n257__spl_),
    .dinb(new_n260__spl_),
    .dout(new_n264_)
  );


  nor2
  g0200
  (
    .dina(G2_spl_011),
    .dinb(G24_spl_000),
    .dout(new_n265_)
  );


  and2
  g0201
  (
    .dina(new_n251__spl_),
    .dinb(new_n254__spl_),
    .dout(new_n266_)
  );


  nor2
  g0202
  (
    .dina(G3_spl_011),
    .dinb(G23_spl_001),
    .dout(new_n267_)
  );


  and2
  g0203
  (
    .dina(new_n245__spl_),
    .dinb(new_n248__spl_),
    .dout(new_n268_)
  );


  nor2
  g0204
  (
    .dina(G4_spl_010),
    .dinb(G22_spl_001),
    .dout(new_n269_)
  );


  anb1
  g0205
  (
    .dina(new_n239__spl_),
    .dinb(new_n242__spl_),
    .dout(new_n270_)
  );


  and1
  g0206
  (
    .dina(G5_spl_010),
    .dinb(G21_spl_010),
    .dout(new_n271_)
  );


  anb2
  g0207
  (
    .dina(new_n233__spl_),
    .dinb(new_n236__spl_),
    .dout(new_n272_)
  );


  and1
  g0208
  (
    .dina(G6_spl_001),
    .dinb(G20_spl_010),
    .dout(new_n273_)
  );


  anb2
  g0209
  (
    .dina(new_n227__spl_),
    .dinb(new_n230__spl_),
    .dout(new_n274_)
  );


  and1
  g0210
  (
    .dina(G7_spl_001),
    .dinb(G19_spl_011),
    .dout(new_n275_)
  );


  nor2
  g0211
  (
    .dina(G9_spl_000),
    .dinb(G17_spl_100),
    .dout(new_n276_)
  );


  and1
  g0212
  (
    .dina(G8_spl_000),
    .dinb(G18_spl_011),
    .dout(new_n277_)
  );


  anb2
  g0213
  (
    .dina(new_n276__spl_),
    .dinb(new_n277__spl_),
    .dout(new_n278_)
  );


  anb1
  g0214
  (
    .dina(new_n276__spl_),
    .dinb(new_n277__spl_),
    .dout(new_n279_)
  );


  anb1
  g0215
  (
    .dina(new_n278__spl_0),
    .dinb(new_n279_),
    .dout(new_n280_)
  );


  anb1
  g0216
  (
    .dina(new_n224__spl_0),
    .dinb(new_n280__spl_),
    .dout(new_n281_)
  );


  anb2
  g0217
  (
    .dina(new_n224__spl_),
    .dinb(new_n280__spl_),
    .dout(new_n282_)
  );


  nab1
  g0218
  (
    .dina(new_n281__spl_),
    .dinb(new_n282_),
    .dout(new_n283_)
  );


  anb2
  g0219
  (
    .dina(new_n275__spl_),
    .dinb(new_n283__spl_),
    .dout(new_n284_)
  );


  anb1
  g0220
  (
    .dina(new_n275__spl_),
    .dinb(new_n283__spl_),
    .dout(new_n285_)
  );


  nab2
  g0221
  (
    .dina(new_n284__spl_),
    .dinb(new_n285_),
    .dout(new_n286_)
  );


  anb1
  g0222
  (
    .dina(new_n274__spl_),
    .dinb(new_n286__spl_),
    .dout(new_n287_)
  );


  anb2
  g0223
  (
    .dina(new_n274__spl_),
    .dinb(new_n286__spl_),
    .dout(new_n288_)
  );


  nab1
  g0224
  (
    .dina(new_n287__spl_),
    .dinb(new_n288_),
    .dout(new_n289_)
  );


  anb2
  g0225
  (
    .dina(new_n273__spl_),
    .dinb(new_n289__spl_),
    .dout(new_n290_)
  );


  anb1
  g0226
  (
    .dina(new_n273__spl_),
    .dinb(new_n289__spl_),
    .dout(new_n291_)
  );


  nab2
  g0227
  (
    .dina(new_n290__spl_),
    .dinb(new_n291_),
    .dout(new_n292_)
  );


  anb1
  g0228
  (
    .dina(new_n272__spl_),
    .dinb(new_n292__spl_),
    .dout(new_n293_)
  );


  anb2
  g0229
  (
    .dina(new_n272__spl_),
    .dinb(new_n292__spl_),
    .dout(new_n294_)
  );


  nab1
  g0230
  (
    .dina(new_n293__spl_),
    .dinb(new_n294_),
    .dout(new_n295_)
  );


  anb2
  g0231
  (
    .dina(new_n271__spl_),
    .dinb(new_n295__spl_),
    .dout(new_n296_)
  );


  anb1
  g0232
  (
    .dina(new_n271__spl_),
    .dinb(new_n295__spl_),
    .dout(new_n297_)
  );


  anb1
  g0233
  (
    .dina(new_n296__spl_),
    .dinb(new_n297_),
    .dout(new_n298_)
  );


  anb2
  g0234
  (
    .dina(new_n270__spl_),
    .dinb(new_n298__spl_),
    .dout(new_n299_)
  );


  anb1
  g0235
  (
    .dina(new_n270__spl_),
    .dinb(new_n298__spl_),
    .dout(new_n300_)
  );


  nab2
  g0236
  (
    .dina(new_n299__spl_),
    .dinb(new_n300_),
    .dout(new_n301_)
  );


  anb1
  g0237
  (
    .dina(new_n269__spl_),
    .dinb(new_n301__spl_),
    .dout(new_n302_)
  );


  anb2
  g0238
  (
    .dina(new_n269__spl_),
    .dinb(new_n301__spl_),
    .dout(new_n303_)
  );


  anb2
  g0239
  (
    .dina(new_n302__spl_),
    .dinb(new_n303_),
    .dout(new_n304_)
  );


  anb1
  g0240
  (
    .dina(new_n268__spl_),
    .dinb(new_n304__spl_),
    .dout(new_n305_)
  );


  anb2
  g0241
  (
    .dina(new_n268__spl_),
    .dinb(new_n304__spl_),
    .dout(new_n306_)
  );


  anb2
  g0242
  (
    .dina(new_n305__spl_),
    .dinb(new_n306_),
    .dout(new_n307_)
  );


  anb1
  g0243
  (
    .dina(new_n267__spl_),
    .dinb(new_n307__spl_),
    .dout(new_n308_)
  );


  anb2
  g0244
  (
    .dina(new_n267__spl_),
    .dinb(new_n307__spl_),
    .dout(new_n309_)
  );


  anb2
  g0245
  (
    .dina(new_n308__spl_),
    .dinb(new_n309_),
    .dout(new_n310_)
  );


  anb1
  g0246
  (
    .dina(new_n266__spl_),
    .dinb(new_n310__spl_),
    .dout(new_n311_)
  );


  anb2
  g0247
  (
    .dina(new_n266__spl_),
    .dinb(new_n310__spl_),
    .dout(new_n312_)
  );


  anb2
  g0248
  (
    .dina(new_n311__spl_),
    .dinb(new_n312_),
    .dout(new_n313_)
  );


  anb1
  g0249
  (
    .dina(new_n265__spl_),
    .dinb(new_n313__spl_),
    .dout(new_n314_)
  );


  anb2
  g0250
  (
    .dina(new_n265__spl_),
    .dinb(new_n313__spl_),
    .dout(new_n315_)
  );


  anb2
  g0251
  (
    .dina(new_n314__spl_),
    .dinb(new_n315_),
    .dout(new_n316_)
  );


  anb1
  g0252
  (
    .dina(new_n264__spl_),
    .dinb(new_n316__spl_),
    .dout(new_n317_)
  );


  anb2
  g0253
  (
    .dina(new_n264__spl_),
    .dinb(new_n316__spl_),
    .dout(new_n318_)
  );


  anb2
  g0254
  (
    .dina(new_n317__spl_),
    .dinb(new_n318_),
    .dout(new_n319_)
  );


  anb1
  g0255
  (
    .dina(new_n263__spl_),
    .dinb(new_n319__spl_),
    .dout(new_n320_)
  );


  anb2
  g0256
  (
    .dina(new_n263__spl_),
    .dinb(new_n319__spl_),
    .dout(new_n321_)
  );


  anb2
  g0257
  (
    .dina(new_n320__spl_),
    .dinb(new_n321_),
    .dout(G6265)
  );


  nor2
  g0258
  (
    .dina(G1_spl_100),
    .dinb(G26_spl_000),
    .dout(new_n323_)
  );


  and2
  g0259
  (
    .dina(new_n317__spl_),
    .dinb(new_n320__spl_),
    .dout(new_n324_)
  );


  nor2
  g0260
  (
    .dina(G2_spl_100),
    .dinb(G25_spl_000),
    .dout(new_n325_)
  );


  and2
  g0261
  (
    .dina(new_n311__spl_),
    .dinb(new_n314__spl_),
    .dout(new_n326_)
  );


  nor2
  g0262
  (
    .dina(G3_spl_011),
    .dinb(G24_spl_001),
    .dout(new_n327_)
  );


  and2
  g0263
  (
    .dina(new_n305__spl_),
    .dinb(new_n308__spl_),
    .dout(new_n328_)
  );


  nor2
  g0264
  (
    .dina(G4_spl_011),
    .dinb(G23_spl_001),
    .dout(new_n329_)
  );


  anb1
  g0265
  (
    .dina(new_n299__spl_),
    .dinb(new_n302__spl_),
    .dout(new_n330_)
  );


  and1
  g0266
  (
    .dina(G5_spl_010),
    .dinb(G22_spl_010),
    .dout(new_n331_)
  );


  anb2
  g0267
  (
    .dina(new_n293__spl_),
    .dinb(new_n296__spl_),
    .dout(new_n332_)
  );


  and1
  g0268
  (
    .dina(G6_spl_010),
    .dinb(G21_spl_010),
    .dout(new_n333_)
  );


  anb2
  g0269
  (
    .dina(new_n287__spl_),
    .dinb(new_n290__spl_),
    .dout(new_n334_)
  );


  and1
  g0270
  (
    .dina(G7_spl_001),
    .dinb(G20_spl_011),
    .dout(new_n335_)
  );


  anb2
  g0271
  (
    .dina(new_n281__spl_),
    .dinb(new_n284__spl_),
    .dout(new_n336_)
  );


  and1
  g0272
  (
    .dina(G8_spl_001),
    .dinb(G19_spl_011),
    .dout(new_n337_)
  );


  nor2
  g0273
  (
    .dina(G10_spl_000),
    .dinb(G17_spl_100),
    .dout(new_n338_)
  );


  and1
  g0274
  (
    .dina(G9_spl_000),
    .dinb(G18_spl_100),
    .dout(new_n339_)
  );


  anb2
  g0275
  (
    .dina(new_n338__spl_),
    .dinb(new_n339__spl_),
    .dout(new_n340_)
  );


  anb1
  g0276
  (
    .dina(new_n338__spl_),
    .dinb(new_n339__spl_),
    .dout(new_n341_)
  );


  anb1
  g0277
  (
    .dina(new_n340__spl_0),
    .dinb(new_n341_),
    .dout(new_n342_)
  );


  anb1
  g0278
  (
    .dina(new_n278__spl_0),
    .dinb(new_n342__spl_),
    .dout(new_n343_)
  );


  anb2
  g0279
  (
    .dina(new_n278__spl_),
    .dinb(new_n342__spl_),
    .dout(new_n344_)
  );


  nab1
  g0280
  (
    .dina(new_n343__spl_),
    .dinb(new_n344_),
    .dout(new_n345_)
  );


  anb2
  g0281
  (
    .dina(new_n337__spl_),
    .dinb(new_n345__spl_),
    .dout(new_n346_)
  );


  anb1
  g0282
  (
    .dina(new_n337__spl_),
    .dinb(new_n345__spl_),
    .dout(new_n347_)
  );


  nab2
  g0283
  (
    .dina(new_n346__spl_),
    .dinb(new_n347_),
    .dout(new_n348_)
  );


  anb1
  g0284
  (
    .dina(new_n336__spl_),
    .dinb(new_n348__spl_),
    .dout(new_n349_)
  );


  anb2
  g0285
  (
    .dina(new_n336__spl_),
    .dinb(new_n348__spl_),
    .dout(new_n350_)
  );


  nab1
  g0286
  (
    .dina(new_n349__spl_),
    .dinb(new_n350_),
    .dout(new_n351_)
  );


  anb2
  g0287
  (
    .dina(new_n335__spl_),
    .dinb(new_n351__spl_),
    .dout(new_n352_)
  );


  anb1
  g0288
  (
    .dina(new_n335__spl_),
    .dinb(new_n351__spl_),
    .dout(new_n353_)
  );


  nab2
  g0289
  (
    .dina(new_n352__spl_),
    .dinb(new_n353_),
    .dout(new_n354_)
  );


  anb1
  g0290
  (
    .dina(new_n334__spl_),
    .dinb(new_n354__spl_),
    .dout(new_n355_)
  );


  anb2
  g0291
  (
    .dina(new_n334__spl_),
    .dinb(new_n354__spl_),
    .dout(new_n356_)
  );


  nab1
  g0292
  (
    .dina(new_n355__spl_),
    .dinb(new_n356_),
    .dout(new_n357_)
  );


  anb2
  g0293
  (
    .dina(new_n333__spl_),
    .dinb(new_n357__spl_),
    .dout(new_n358_)
  );


  anb1
  g0294
  (
    .dina(new_n333__spl_),
    .dinb(new_n357__spl_),
    .dout(new_n359_)
  );


  nab2
  g0295
  (
    .dina(new_n358__spl_),
    .dinb(new_n359_),
    .dout(new_n360_)
  );


  anb1
  g0296
  (
    .dina(new_n332__spl_),
    .dinb(new_n360__spl_),
    .dout(new_n361_)
  );


  anb2
  g0297
  (
    .dina(new_n332__spl_),
    .dinb(new_n360__spl_),
    .dout(new_n362_)
  );


  nab1
  g0298
  (
    .dina(new_n361__spl_),
    .dinb(new_n362_),
    .dout(new_n363_)
  );


  anb2
  g0299
  (
    .dina(new_n331__spl_),
    .dinb(new_n363__spl_),
    .dout(new_n364_)
  );


  anb1
  g0300
  (
    .dina(new_n331__spl_),
    .dinb(new_n363__spl_),
    .dout(new_n365_)
  );


  anb1
  g0301
  (
    .dina(new_n364__spl_),
    .dinb(new_n365_),
    .dout(new_n366_)
  );


  anb2
  g0302
  (
    .dina(new_n330__spl_),
    .dinb(new_n366__spl_),
    .dout(new_n367_)
  );


  anb1
  g0303
  (
    .dina(new_n330__spl_),
    .dinb(new_n366__spl_),
    .dout(new_n368_)
  );


  nab2
  g0304
  (
    .dina(new_n367__spl_),
    .dinb(new_n368_),
    .dout(new_n369_)
  );


  anb1
  g0305
  (
    .dina(new_n329__spl_),
    .dinb(new_n369__spl_),
    .dout(new_n370_)
  );


  anb2
  g0306
  (
    .dina(new_n329__spl_),
    .dinb(new_n369__spl_),
    .dout(new_n371_)
  );


  anb2
  g0307
  (
    .dina(new_n370__spl_),
    .dinb(new_n371_),
    .dout(new_n372_)
  );


  anb1
  g0308
  (
    .dina(new_n328__spl_),
    .dinb(new_n372__spl_),
    .dout(new_n373_)
  );


  anb2
  g0309
  (
    .dina(new_n328__spl_),
    .dinb(new_n372__spl_),
    .dout(new_n374_)
  );


  anb2
  g0310
  (
    .dina(new_n373__spl_),
    .dinb(new_n374_),
    .dout(new_n375_)
  );


  anb1
  g0311
  (
    .dina(new_n327__spl_),
    .dinb(new_n375__spl_),
    .dout(new_n376_)
  );


  anb2
  g0312
  (
    .dina(new_n327__spl_),
    .dinb(new_n375__spl_),
    .dout(new_n377_)
  );


  anb2
  g0313
  (
    .dina(new_n376__spl_),
    .dinb(new_n377_),
    .dout(new_n378_)
  );


  anb1
  g0314
  (
    .dina(new_n326__spl_),
    .dinb(new_n378__spl_),
    .dout(new_n379_)
  );


  anb2
  g0315
  (
    .dina(new_n326__spl_),
    .dinb(new_n378__spl_),
    .dout(new_n380_)
  );


  anb2
  g0316
  (
    .dina(new_n379__spl_),
    .dinb(new_n380_),
    .dout(new_n381_)
  );


  anb1
  g0317
  (
    .dina(new_n325__spl_),
    .dinb(new_n381__spl_),
    .dout(new_n382_)
  );


  anb2
  g0318
  (
    .dina(new_n325__spl_),
    .dinb(new_n381__spl_),
    .dout(new_n383_)
  );


  anb2
  g0319
  (
    .dina(new_n382__spl_),
    .dinb(new_n383_),
    .dout(new_n384_)
  );


  anb1
  g0320
  (
    .dina(new_n324__spl_),
    .dinb(new_n384__spl_),
    .dout(new_n385_)
  );


  anb2
  g0321
  (
    .dina(new_n324__spl_),
    .dinb(new_n384__spl_),
    .dout(new_n386_)
  );


  anb2
  g0322
  (
    .dina(new_n385__spl_),
    .dinb(new_n386_),
    .dout(new_n387_)
  );


  anb1
  g0323
  (
    .dina(new_n323__spl_),
    .dinb(new_n387__spl_),
    .dout(new_n388_)
  );


  anb2
  g0324
  (
    .dina(new_n323__spl_),
    .dinb(new_n387__spl_),
    .dout(new_n389_)
  );


  anb2
  g0325
  (
    .dina(new_n388__spl_),
    .dinb(new_n389_),
    .dout(G6266)
  );


  nor2
  g0326
  (
    .dina(G1_spl_101),
    .dinb(G27_spl_000),
    .dout(new_n391_)
  );


  and2
  g0327
  (
    .dina(new_n385__spl_),
    .dinb(new_n388__spl_),
    .dout(new_n392_)
  );


  nor2
  g0328
  (
    .dina(G2_spl_100),
    .dinb(G26_spl_000),
    .dout(new_n393_)
  );


  and2
  g0329
  (
    .dina(new_n379__spl_),
    .dinb(new_n382__spl_),
    .dout(new_n394_)
  );


  nor2
  g0330
  (
    .dina(G3_spl_100),
    .dinb(G25_spl_001),
    .dout(new_n395_)
  );


  and2
  g0331
  (
    .dina(new_n373__spl_),
    .dinb(new_n376__spl_),
    .dout(new_n396_)
  );


  nor2
  g0332
  (
    .dina(G4_spl_011),
    .dinb(G24_spl_001),
    .dout(new_n397_)
  );


  anb1
  g0333
  (
    .dina(new_n367__spl_),
    .dinb(new_n370__spl_),
    .dout(new_n398_)
  );


  and1
  g0334
  (
    .dina(G5_spl_011),
    .dinb(G23_spl_010),
    .dout(new_n399_)
  );


  anb2
  g0335
  (
    .dina(new_n361__spl_),
    .dinb(new_n364__spl_),
    .dout(new_n400_)
  );


  and1
  g0336
  (
    .dina(G6_spl_010),
    .dinb(G22_spl_010),
    .dout(new_n401_)
  );


  anb2
  g0337
  (
    .dina(new_n355__spl_),
    .dinb(new_n358__spl_),
    .dout(new_n402_)
  );


  and1
  g0338
  (
    .dina(G7_spl_010),
    .dinb(G21_spl_011),
    .dout(new_n403_)
  );


  anb2
  g0339
  (
    .dina(new_n349__spl_),
    .dinb(new_n352__spl_),
    .dout(new_n404_)
  );


  and1
  g0340
  (
    .dina(G8_spl_001),
    .dinb(G20_spl_011),
    .dout(new_n405_)
  );


  anb2
  g0341
  (
    .dina(new_n343__spl_),
    .dinb(new_n346__spl_),
    .dout(new_n406_)
  );


  and1
  g0342
  (
    .dina(G9_spl_001),
    .dinb(G19_spl_100),
    .dout(new_n407_)
  );


  nor2
  g0343
  (
    .dina(G11_spl_000),
    .dinb(G17_spl_101),
    .dout(new_n408_)
  );


  and1
  g0344
  (
    .dina(G10_spl_000),
    .dinb(G18_spl_100),
    .dout(new_n409_)
  );


  anb2
  g0345
  (
    .dina(new_n408__spl_),
    .dinb(new_n409__spl_),
    .dout(new_n410_)
  );


  anb1
  g0346
  (
    .dina(new_n408__spl_),
    .dinb(new_n409__spl_),
    .dout(new_n411_)
  );


  anb1
  g0347
  (
    .dina(new_n410__spl_0),
    .dinb(new_n411_),
    .dout(new_n412_)
  );


  anb1
  g0348
  (
    .dina(new_n340__spl_0),
    .dinb(new_n412__spl_),
    .dout(new_n413_)
  );


  anb2
  g0349
  (
    .dina(new_n340__spl_),
    .dinb(new_n412__spl_),
    .dout(new_n414_)
  );


  nab1
  g0350
  (
    .dina(new_n413__spl_),
    .dinb(new_n414_),
    .dout(new_n415_)
  );


  anb2
  g0351
  (
    .dina(new_n407__spl_),
    .dinb(new_n415__spl_),
    .dout(new_n416_)
  );


  anb1
  g0352
  (
    .dina(new_n407__spl_),
    .dinb(new_n415__spl_),
    .dout(new_n417_)
  );


  nab2
  g0353
  (
    .dina(new_n416__spl_),
    .dinb(new_n417_),
    .dout(new_n418_)
  );


  anb1
  g0354
  (
    .dina(new_n406__spl_),
    .dinb(new_n418__spl_),
    .dout(new_n419_)
  );


  anb2
  g0355
  (
    .dina(new_n406__spl_),
    .dinb(new_n418__spl_),
    .dout(new_n420_)
  );


  nab1
  g0356
  (
    .dina(new_n419__spl_),
    .dinb(new_n420_),
    .dout(new_n421_)
  );


  anb2
  g0357
  (
    .dina(new_n405__spl_),
    .dinb(new_n421__spl_),
    .dout(new_n422_)
  );


  anb1
  g0358
  (
    .dina(new_n405__spl_),
    .dinb(new_n421__spl_),
    .dout(new_n423_)
  );


  nab2
  g0359
  (
    .dina(new_n422__spl_),
    .dinb(new_n423_),
    .dout(new_n424_)
  );


  anb1
  g0360
  (
    .dina(new_n404__spl_),
    .dinb(new_n424__spl_),
    .dout(new_n425_)
  );


  anb2
  g0361
  (
    .dina(new_n404__spl_),
    .dinb(new_n424__spl_),
    .dout(new_n426_)
  );


  nab1
  g0362
  (
    .dina(new_n425__spl_),
    .dinb(new_n426_),
    .dout(new_n427_)
  );


  anb2
  g0363
  (
    .dina(new_n403__spl_),
    .dinb(new_n427__spl_),
    .dout(new_n428_)
  );


  anb1
  g0364
  (
    .dina(new_n403__spl_),
    .dinb(new_n427__spl_),
    .dout(new_n429_)
  );


  nab2
  g0365
  (
    .dina(new_n428__spl_),
    .dinb(new_n429_),
    .dout(new_n430_)
  );


  anb1
  g0366
  (
    .dina(new_n402__spl_),
    .dinb(new_n430__spl_),
    .dout(new_n431_)
  );


  anb2
  g0367
  (
    .dina(new_n402__spl_),
    .dinb(new_n430__spl_),
    .dout(new_n432_)
  );


  nab1
  g0368
  (
    .dina(new_n431__spl_),
    .dinb(new_n432_),
    .dout(new_n433_)
  );


  anb2
  g0369
  (
    .dina(new_n401__spl_),
    .dinb(new_n433__spl_),
    .dout(new_n434_)
  );


  anb1
  g0370
  (
    .dina(new_n401__spl_),
    .dinb(new_n433__spl_),
    .dout(new_n435_)
  );


  nab2
  g0371
  (
    .dina(new_n434__spl_),
    .dinb(new_n435_),
    .dout(new_n436_)
  );


  anb1
  g0372
  (
    .dina(new_n400__spl_),
    .dinb(new_n436__spl_),
    .dout(new_n437_)
  );


  anb2
  g0373
  (
    .dina(new_n400__spl_),
    .dinb(new_n436__spl_),
    .dout(new_n438_)
  );


  nab1
  g0374
  (
    .dina(new_n437__spl_),
    .dinb(new_n438_),
    .dout(new_n439_)
  );


  anb2
  g0375
  (
    .dina(new_n399__spl_),
    .dinb(new_n439__spl_),
    .dout(new_n440_)
  );


  anb1
  g0376
  (
    .dina(new_n399__spl_),
    .dinb(new_n439__spl_),
    .dout(new_n441_)
  );


  anb1
  g0377
  (
    .dina(new_n440__spl_),
    .dinb(new_n441_),
    .dout(new_n442_)
  );


  anb2
  g0378
  (
    .dina(new_n398__spl_),
    .dinb(new_n442__spl_),
    .dout(new_n443_)
  );


  anb1
  g0379
  (
    .dina(new_n398__spl_),
    .dinb(new_n442__spl_),
    .dout(new_n444_)
  );


  nab2
  g0380
  (
    .dina(new_n443__spl_),
    .dinb(new_n444_),
    .dout(new_n445_)
  );


  anb1
  g0381
  (
    .dina(new_n397__spl_),
    .dinb(new_n445__spl_),
    .dout(new_n446_)
  );


  anb2
  g0382
  (
    .dina(new_n397__spl_),
    .dinb(new_n445__spl_),
    .dout(new_n447_)
  );


  anb2
  g0383
  (
    .dina(new_n446__spl_),
    .dinb(new_n447_),
    .dout(new_n448_)
  );


  anb1
  g0384
  (
    .dina(new_n396__spl_),
    .dinb(new_n448__spl_),
    .dout(new_n449_)
  );


  anb2
  g0385
  (
    .dina(new_n396__spl_),
    .dinb(new_n448__spl_),
    .dout(new_n450_)
  );


  anb2
  g0386
  (
    .dina(new_n449__spl_),
    .dinb(new_n450_),
    .dout(new_n451_)
  );


  anb1
  g0387
  (
    .dina(new_n395__spl_),
    .dinb(new_n451__spl_),
    .dout(new_n452_)
  );


  anb2
  g0388
  (
    .dina(new_n395__spl_),
    .dinb(new_n451__spl_),
    .dout(new_n453_)
  );


  anb2
  g0389
  (
    .dina(new_n452__spl_),
    .dinb(new_n453_),
    .dout(new_n454_)
  );


  anb1
  g0390
  (
    .dina(new_n394__spl_),
    .dinb(new_n454__spl_),
    .dout(new_n455_)
  );


  anb2
  g0391
  (
    .dina(new_n394__spl_),
    .dinb(new_n454__spl_),
    .dout(new_n456_)
  );


  anb2
  g0392
  (
    .dina(new_n455__spl_),
    .dinb(new_n456_),
    .dout(new_n457_)
  );


  anb1
  g0393
  (
    .dina(new_n393__spl_),
    .dinb(new_n457__spl_),
    .dout(new_n458_)
  );


  anb2
  g0394
  (
    .dina(new_n393__spl_),
    .dinb(new_n457__spl_),
    .dout(new_n459_)
  );


  anb2
  g0395
  (
    .dina(new_n458__spl_),
    .dinb(new_n459_),
    .dout(new_n460_)
  );


  anb1
  g0396
  (
    .dina(new_n392__spl_),
    .dinb(new_n460__spl_),
    .dout(new_n461_)
  );


  anb2
  g0397
  (
    .dina(new_n392__spl_),
    .dinb(new_n460__spl_),
    .dout(new_n462_)
  );


  anb2
  g0398
  (
    .dina(new_n461__spl_),
    .dinb(new_n462_),
    .dout(new_n463_)
  );


  anb1
  g0399
  (
    .dina(new_n391__spl_),
    .dinb(new_n463__spl_),
    .dout(new_n464_)
  );


  anb2
  g0400
  (
    .dina(new_n391__spl_),
    .dinb(new_n463__spl_),
    .dout(new_n465_)
  );


  anb2
  g0401
  (
    .dina(new_n464__spl_),
    .dinb(new_n465_),
    .dout(G6267)
  );


  nor2
  g0402
  (
    .dina(G1_spl_101),
    .dinb(G28_spl_000),
    .dout(new_n467_)
  );


  and2
  g0403
  (
    .dina(new_n461__spl_),
    .dinb(new_n464__spl_),
    .dout(new_n468_)
  );


  nor2
  g0404
  (
    .dina(G2_spl_101),
    .dinb(G27_spl_000),
    .dout(new_n469_)
  );


  and2
  g0405
  (
    .dina(new_n455__spl_),
    .dinb(new_n458__spl_),
    .dout(new_n470_)
  );


  nor2
  g0406
  (
    .dina(G3_spl_100),
    .dinb(G26_spl_001),
    .dout(new_n471_)
  );


  and2
  g0407
  (
    .dina(new_n449__spl_),
    .dinb(new_n452__spl_),
    .dout(new_n472_)
  );


  nor2
  g0408
  (
    .dina(G4_spl_100),
    .dinb(G25_spl_001),
    .dout(new_n473_)
  );


  anb1
  g0409
  (
    .dina(new_n443__spl_),
    .dinb(new_n446__spl_),
    .dout(new_n474_)
  );


  and1
  g0410
  (
    .dina(G5_spl_011),
    .dinb(G24_spl_010),
    .dout(new_n475_)
  );


  anb2
  g0411
  (
    .dina(new_n437__spl_),
    .dinb(new_n440__spl_),
    .dout(new_n476_)
  );


  and1
  g0412
  (
    .dina(G6_spl_011),
    .dinb(G23_spl_010),
    .dout(new_n477_)
  );


  anb2
  g0413
  (
    .dina(new_n431__spl_),
    .dinb(new_n434__spl_),
    .dout(new_n478_)
  );


  and1
  g0414
  (
    .dina(G7_spl_010),
    .dinb(G22_spl_011),
    .dout(new_n479_)
  );


  anb2
  g0415
  (
    .dina(new_n425__spl_),
    .dinb(new_n428__spl_),
    .dout(new_n480_)
  );


  and1
  g0416
  (
    .dina(G8_spl_010),
    .dinb(G21_spl_011),
    .dout(new_n481_)
  );


  anb2
  g0417
  (
    .dina(new_n419__spl_),
    .dinb(new_n422__spl_),
    .dout(new_n482_)
  );


  and1
  g0418
  (
    .dina(G9_spl_001),
    .dinb(G20_spl_100),
    .dout(new_n483_)
  );


  anb2
  g0419
  (
    .dina(new_n413__spl_),
    .dinb(new_n416__spl_),
    .dout(new_n484_)
  );


  and1
  g0420
  (
    .dina(G10_spl_001),
    .dinb(G19_spl_100),
    .dout(new_n485_)
  );


  nor2
  g0421
  (
    .dina(G12_spl_000),
    .dinb(G17_spl_101),
    .dout(new_n486_)
  );


  and1
  g0422
  (
    .dina(G11_spl_000),
    .dinb(G18_spl_101),
    .dout(new_n487_)
  );


  anb2
  g0423
  (
    .dina(new_n486__spl_),
    .dinb(new_n487__spl_),
    .dout(new_n488_)
  );


  anb1
  g0424
  (
    .dina(new_n486__spl_),
    .dinb(new_n487__spl_),
    .dout(new_n489_)
  );


  anb1
  g0425
  (
    .dina(new_n488__spl_0),
    .dinb(new_n489_),
    .dout(new_n490_)
  );


  anb1
  g0426
  (
    .dina(new_n410__spl_0),
    .dinb(new_n490__spl_),
    .dout(new_n491_)
  );


  anb2
  g0427
  (
    .dina(new_n410__spl_),
    .dinb(new_n490__spl_),
    .dout(new_n492_)
  );


  nab1
  g0428
  (
    .dina(new_n491__spl_),
    .dinb(new_n492_),
    .dout(new_n493_)
  );


  anb2
  g0429
  (
    .dina(new_n485__spl_),
    .dinb(new_n493__spl_),
    .dout(new_n494_)
  );


  anb1
  g0430
  (
    .dina(new_n485__spl_),
    .dinb(new_n493__spl_),
    .dout(new_n495_)
  );


  nab2
  g0431
  (
    .dina(new_n494__spl_),
    .dinb(new_n495_),
    .dout(new_n496_)
  );


  anb1
  g0432
  (
    .dina(new_n484__spl_),
    .dinb(new_n496__spl_),
    .dout(new_n497_)
  );


  anb2
  g0433
  (
    .dina(new_n484__spl_),
    .dinb(new_n496__spl_),
    .dout(new_n498_)
  );


  nab1
  g0434
  (
    .dina(new_n497__spl_),
    .dinb(new_n498_),
    .dout(new_n499_)
  );


  anb2
  g0435
  (
    .dina(new_n483__spl_),
    .dinb(new_n499__spl_),
    .dout(new_n500_)
  );


  anb1
  g0436
  (
    .dina(new_n483__spl_),
    .dinb(new_n499__spl_),
    .dout(new_n501_)
  );


  nab2
  g0437
  (
    .dina(new_n500__spl_),
    .dinb(new_n501_),
    .dout(new_n502_)
  );


  anb1
  g0438
  (
    .dina(new_n482__spl_),
    .dinb(new_n502__spl_),
    .dout(new_n503_)
  );


  anb2
  g0439
  (
    .dina(new_n482__spl_),
    .dinb(new_n502__spl_),
    .dout(new_n504_)
  );


  nab1
  g0440
  (
    .dina(new_n503__spl_),
    .dinb(new_n504_),
    .dout(new_n505_)
  );


  anb2
  g0441
  (
    .dina(new_n481__spl_),
    .dinb(new_n505__spl_),
    .dout(new_n506_)
  );


  anb1
  g0442
  (
    .dina(new_n481__spl_),
    .dinb(new_n505__spl_),
    .dout(new_n507_)
  );


  nab2
  g0443
  (
    .dina(new_n506__spl_),
    .dinb(new_n507_),
    .dout(new_n508_)
  );


  anb1
  g0444
  (
    .dina(new_n480__spl_),
    .dinb(new_n508__spl_),
    .dout(new_n509_)
  );


  anb2
  g0445
  (
    .dina(new_n480__spl_),
    .dinb(new_n508__spl_),
    .dout(new_n510_)
  );


  nab1
  g0446
  (
    .dina(new_n509__spl_),
    .dinb(new_n510_),
    .dout(new_n511_)
  );


  anb2
  g0447
  (
    .dina(new_n479__spl_),
    .dinb(new_n511__spl_),
    .dout(new_n512_)
  );


  anb1
  g0448
  (
    .dina(new_n479__spl_),
    .dinb(new_n511__spl_),
    .dout(new_n513_)
  );


  nab2
  g0449
  (
    .dina(new_n512__spl_),
    .dinb(new_n513_),
    .dout(new_n514_)
  );


  anb1
  g0450
  (
    .dina(new_n478__spl_),
    .dinb(new_n514__spl_),
    .dout(new_n515_)
  );


  anb2
  g0451
  (
    .dina(new_n478__spl_),
    .dinb(new_n514__spl_),
    .dout(new_n516_)
  );


  nab1
  g0452
  (
    .dina(new_n515__spl_),
    .dinb(new_n516_),
    .dout(new_n517_)
  );


  anb2
  g0453
  (
    .dina(new_n477__spl_),
    .dinb(new_n517__spl_),
    .dout(new_n518_)
  );


  anb1
  g0454
  (
    .dina(new_n477__spl_),
    .dinb(new_n517__spl_),
    .dout(new_n519_)
  );


  nab2
  g0455
  (
    .dina(new_n518__spl_),
    .dinb(new_n519_),
    .dout(new_n520_)
  );


  anb1
  g0456
  (
    .dina(new_n476__spl_),
    .dinb(new_n520__spl_),
    .dout(new_n521_)
  );


  anb2
  g0457
  (
    .dina(new_n476__spl_),
    .dinb(new_n520__spl_),
    .dout(new_n522_)
  );


  nab1
  g0458
  (
    .dina(new_n521__spl_),
    .dinb(new_n522_),
    .dout(new_n523_)
  );


  anb2
  g0459
  (
    .dina(new_n475__spl_),
    .dinb(new_n523__spl_),
    .dout(new_n524_)
  );


  anb1
  g0460
  (
    .dina(new_n475__spl_),
    .dinb(new_n523__spl_),
    .dout(new_n525_)
  );


  anb1
  g0461
  (
    .dina(new_n524__spl_),
    .dinb(new_n525_),
    .dout(new_n526_)
  );


  anb2
  g0462
  (
    .dina(new_n474__spl_),
    .dinb(new_n526__spl_),
    .dout(new_n527_)
  );


  anb1
  g0463
  (
    .dina(new_n474__spl_),
    .dinb(new_n526__spl_),
    .dout(new_n528_)
  );


  nab2
  g0464
  (
    .dina(new_n527__spl_),
    .dinb(new_n528_),
    .dout(new_n529_)
  );


  anb1
  g0465
  (
    .dina(new_n473__spl_),
    .dinb(new_n529__spl_),
    .dout(new_n530_)
  );


  anb2
  g0466
  (
    .dina(new_n473__spl_),
    .dinb(new_n529__spl_),
    .dout(new_n531_)
  );


  anb2
  g0467
  (
    .dina(new_n530__spl_),
    .dinb(new_n531_),
    .dout(new_n532_)
  );


  anb1
  g0468
  (
    .dina(new_n472__spl_),
    .dinb(new_n532__spl_),
    .dout(new_n533_)
  );


  anb2
  g0469
  (
    .dina(new_n472__spl_),
    .dinb(new_n532__spl_),
    .dout(new_n534_)
  );


  anb2
  g0470
  (
    .dina(new_n533__spl_),
    .dinb(new_n534_),
    .dout(new_n535_)
  );


  anb1
  g0471
  (
    .dina(new_n471__spl_),
    .dinb(new_n535__spl_),
    .dout(new_n536_)
  );


  anb2
  g0472
  (
    .dina(new_n471__spl_),
    .dinb(new_n535__spl_),
    .dout(new_n537_)
  );


  anb2
  g0473
  (
    .dina(new_n536__spl_),
    .dinb(new_n537_),
    .dout(new_n538_)
  );


  anb1
  g0474
  (
    .dina(new_n470__spl_),
    .dinb(new_n538__spl_),
    .dout(new_n539_)
  );


  anb2
  g0475
  (
    .dina(new_n470__spl_),
    .dinb(new_n538__spl_),
    .dout(new_n540_)
  );


  anb2
  g0476
  (
    .dina(new_n539__spl_),
    .dinb(new_n540_),
    .dout(new_n541_)
  );


  anb1
  g0477
  (
    .dina(new_n469__spl_),
    .dinb(new_n541__spl_),
    .dout(new_n542_)
  );


  anb2
  g0478
  (
    .dina(new_n469__spl_),
    .dinb(new_n541__spl_),
    .dout(new_n543_)
  );


  anb2
  g0479
  (
    .dina(new_n542__spl_),
    .dinb(new_n543_),
    .dout(new_n544_)
  );


  anb1
  g0480
  (
    .dina(new_n468__spl_),
    .dinb(new_n544__spl_),
    .dout(new_n545_)
  );


  anb2
  g0481
  (
    .dina(new_n468__spl_),
    .dinb(new_n544__spl_),
    .dout(new_n546_)
  );


  anb2
  g0482
  (
    .dina(new_n545__spl_),
    .dinb(new_n546_),
    .dout(new_n547_)
  );


  anb1
  g0483
  (
    .dina(new_n467__spl_),
    .dinb(new_n547__spl_),
    .dout(new_n548_)
  );


  anb2
  g0484
  (
    .dina(new_n467__spl_),
    .dinb(new_n547__spl_),
    .dout(new_n549_)
  );


  anb2
  g0485
  (
    .dina(new_n548__spl_),
    .dinb(new_n549_),
    .dout(G6268)
  );


  nor2
  g0486
  (
    .dina(G1_spl_110),
    .dinb(G29_spl_000),
    .dout(new_n551_)
  );


  and2
  g0487
  (
    .dina(new_n545__spl_),
    .dinb(new_n548__spl_),
    .dout(new_n552_)
  );


  nor2
  g0488
  (
    .dina(G2_spl_101),
    .dinb(G28_spl_000),
    .dout(new_n553_)
  );


  and2
  g0489
  (
    .dina(new_n539__spl_),
    .dinb(new_n542__spl_),
    .dout(new_n554_)
  );


  nor2
  g0490
  (
    .dina(G3_spl_101),
    .dinb(G27_spl_001),
    .dout(new_n555_)
  );


  and2
  g0491
  (
    .dina(new_n533__spl_),
    .dinb(new_n536__spl_),
    .dout(new_n556_)
  );


  nor2
  g0492
  (
    .dina(G4_spl_100),
    .dinb(G26_spl_001),
    .dout(new_n557_)
  );


  anb1
  g0493
  (
    .dina(new_n527__spl_),
    .dinb(new_n530__spl_),
    .dout(new_n558_)
  );


  and1
  g0494
  (
    .dina(G5_spl_100),
    .dinb(G25_spl_010),
    .dout(new_n559_)
  );


  anb2
  g0495
  (
    .dina(new_n521__spl_),
    .dinb(new_n524__spl_),
    .dout(new_n560_)
  );


  and1
  g0496
  (
    .dina(G6_spl_011),
    .dinb(G24_spl_010),
    .dout(new_n561_)
  );


  anb2
  g0497
  (
    .dina(new_n515__spl_),
    .dinb(new_n518__spl_),
    .dout(new_n562_)
  );


  and1
  g0498
  (
    .dina(G7_spl_011),
    .dinb(G23_spl_011),
    .dout(new_n563_)
  );


  anb2
  g0499
  (
    .dina(new_n509__spl_),
    .dinb(new_n512__spl_),
    .dout(new_n564_)
  );


  and1
  g0500
  (
    .dina(G8_spl_010),
    .dinb(G22_spl_011),
    .dout(new_n565_)
  );


  anb2
  g0501
  (
    .dina(new_n503__spl_),
    .dinb(new_n506__spl_),
    .dout(new_n566_)
  );


  and1
  g0502
  (
    .dina(G9_spl_010),
    .dinb(G21_spl_100),
    .dout(new_n567_)
  );


  anb2
  g0503
  (
    .dina(new_n497__spl_),
    .dinb(new_n500__spl_),
    .dout(new_n568_)
  );


  and1
  g0504
  (
    .dina(G10_spl_001),
    .dinb(G20_spl_100),
    .dout(new_n569_)
  );


  anb2
  g0505
  (
    .dina(new_n491__spl_),
    .dinb(new_n494__spl_),
    .dout(new_n570_)
  );


  and1
  g0506
  (
    .dina(G11_spl_001),
    .dinb(G19_spl_101),
    .dout(new_n571_)
  );


  nor2
  g0507
  (
    .dina(G13_spl_000),
    .dinb(G17_spl_110),
    .dout(new_n572_)
  );


  and1
  g0508
  (
    .dina(G12_spl_000),
    .dinb(G18_spl_101),
    .dout(new_n573_)
  );


  anb2
  g0509
  (
    .dina(new_n572__spl_),
    .dinb(new_n573__spl_),
    .dout(new_n574_)
  );


  anb1
  g0510
  (
    .dina(new_n572__spl_),
    .dinb(new_n573__spl_),
    .dout(new_n575_)
  );


  anb1
  g0511
  (
    .dina(new_n574__spl_0),
    .dinb(new_n575_),
    .dout(new_n576_)
  );


  anb1
  g0512
  (
    .dina(new_n488__spl_0),
    .dinb(new_n576__spl_),
    .dout(new_n577_)
  );


  anb2
  g0513
  (
    .dina(new_n488__spl_),
    .dinb(new_n576__spl_),
    .dout(new_n578_)
  );


  nab1
  g0514
  (
    .dina(new_n577__spl_),
    .dinb(new_n578_),
    .dout(new_n579_)
  );


  anb2
  g0515
  (
    .dina(new_n571__spl_),
    .dinb(new_n579__spl_),
    .dout(new_n580_)
  );


  anb1
  g0516
  (
    .dina(new_n571__spl_),
    .dinb(new_n579__spl_),
    .dout(new_n581_)
  );


  nab2
  g0517
  (
    .dina(new_n580__spl_),
    .dinb(new_n581_),
    .dout(new_n582_)
  );


  anb1
  g0518
  (
    .dina(new_n570__spl_),
    .dinb(new_n582__spl_),
    .dout(new_n583_)
  );


  anb2
  g0519
  (
    .dina(new_n570__spl_),
    .dinb(new_n582__spl_),
    .dout(new_n584_)
  );


  nab1
  g0520
  (
    .dina(new_n583__spl_),
    .dinb(new_n584_),
    .dout(new_n585_)
  );


  anb2
  g0521
  (
    .dina(new_n569__spl_),
    .dinb(new_n585__spl_),
    .dout(new_n586_)
  );


  anb1
  g0522
  (
    .dina(new_n569__spl_),
    .dinb(new_n585__spl_),
    .dout(new_n587_)
  );


  nab2
  g0523
  (
    .dina(new_n586__spl_),
    .dinb(new_n587_),
    .dout(new_n588_)
  );


  anb1
  g0524
  (
    .dina(new_n568__spl_),
    .dinb(new_n588__spl_),
    .dout(new_n589_)
  );


  anb2
  g0525
  (
    .dina(new_n568__spl_),
    .dinb(new_n588__spl_),
    .dout(new_n590_)
  );


  nab1
  g0526
  (
    .dina(new_n589__spl_),
    .dinb(new_n590_),
    .dout(new_n591_)
  );


  anb2
  g0527
  (
    .dina(new_n567__spl_),
    .dinb(new_n591__spl_),
    .dout(new_n592_)
  );


  anb1
  g0528
  (
    .dina(new_n567__spl_),
    .dinb(new_n591__spl_),
    .dout(new_n593_)
  );


  nab2
  g0529
  (
    .dina(new_n592__spl_),
    .dinb(new_n593_),
    .dout(new_n594_)
  );


  anb1
  g0530
  (
    .dina(new_n566__spl_),
    .dinb(new_n594__spl_),
    .dout(new_n595_)
  );


  anb2
  g0531
  (
    .dina(new_n566__spl_),
    .dinb(new_n594__spl_),
    .dout(new_n596_)
  );


  nab1
  g0532
  (
    .dina(new_n595__spl_),
    .dinb(new_n596_),
    .dout(new_n597_)
  );


  anb2
  g0533
  (
    .dina(new_n565__spl_),
    .dinb(new_n597__spl_),
    .dout(new_n598_)
  );


  anb1
  g0534
  (
    .dina(new_n565__spl_),
    .dinb(new_n597__spl_),
    .dout(new_n599_)
  );


  nab2
  g0535
  (
    .dina(new_n598__spl_),
    .dinb(new_n599_),
    .dout(new_n600_)
  );


  anb1
  g0536
  (
    .dina(new_n564__spl_),
    .dinb(new_n600__spl_),
    .dout(new_n601_)
  );


  anb2
  g0537
  (
    .dina(new_n564__spl_),
    .dinb(new_n600__spl_),
    .dout(new_n602_)
  );


  nab1
  g0538
  (
    .dina(new_n601__spl_),
    .dinb(new_n602_),
    .dout(new_n603_)
  );


  anb2
  g0539
  (
    .dina(new_n563__spl_),
    .dinb(new_n603__spl_),
    .dout(new_n604_)
  );


  anb1
  g0540
  (
    .dina(new_n563__spl_),
    .dinb(new_n603__spl_),
    .dout(new_n605_)
  );


  nab2
  g0541
  (
    .dina(new_n604__spl_),
    .dinb(new_n605_),
    .dout(new_n606_)
  );


  anb1
  g0542
  (
    .dina(new_n562__spl_),
    .dinb(new_n606__spl_),
    .dout(new_n607_)
  );


  anb2
  g0543
  (
    .dina(new_n562__spl_),
    .dinb(new_n606__spl_),
    .dout(new_n608_)
  );


  nab1
  g0544
  (
    .dina(new_n607__spl_),
    .dinb(new_n608_),
    .dout(new_n609_)
  );


  anb2
  g0545
  (
    .dina(new_n561__spl_),
    .dinb(new_n609__spl_),
    .dout(new_n610_)
  );


  anb1
  g0546
  (
    .dina(new_n561__spl_),
    .dinb(new_n609__spl_),
    .dout(new_n611_)
  );


  nab2
  g0547
  (
    .dina(new_n610__spl_),
    .dinb(new_n611_),
    .dout(new_n612_)
  );


  anb1
  g0548
  (
    .dina(new_n560__spl_),
    .dinb(new_n612__spl_),
    .dout(new_n613_)
  );


  anb2
  g0549
  (
    .dina(new_n560__spl_),
    .dinb(new_n612__spl_),
    .dout(new_n614_)
  );


  nab1
  g0550
  (
    .dina(new_n613__spl_),
    .dinb(new_n614_),
    .dout(new_n615_)
  );


  anb2
  g0551
  (
    .dina(new_n559__spl_),
    .dinb(new_n615__spl_),
    .dout(new_n616_)
  );


  anb1
  g0552
  (
    .dina(new_n559__spl_),
    .dinb(new_n615__spl_),
    .dout(new_n617_)
  );


  anb1
  g0553
  (
    .dina(new_n616__spl_),
    .dinb(new_n617_),
    .dout(new_n618_)
  );


  anb2
  g0554
  (
    .dina(new_n558__spl_),
    .dinb(new_n618__spl_),
    .dout(new_n619_)
  );


  anb1
  g0555
  (
    .dina(new_n558__spl_),
    .dinb(new_n618__spl_),
    .dout(new_n620_)
  );


  nab2
  g0556
  (
    .dina(new_n619__spl_),
    .dinb(new_n620_),
    .dout(new_n621_)
  );


  anb1
  g0557
  (
    .dina(new_n557__spl_),
    .dinb(new_n621__spl_),
    .dout(new_n622_)
  );


  anb2
  g0558
  (
    .dina(new_n557__spl_),
    .dinb(new_n621__spl_),
    .dout(new_n623_)
  );


  anb2
  g0559
  (
    .dina(new_n622__spl_),
    .dinb(new_n623_),
    .dout(new_n624_)
  );


  anb1
  g0560
  (
    .dina(new_n556__spl_),
    .dinb(new_n624__spl_),
    .dout(new_n625_)
  );


  anb2
  g0561
  (
    .dina(new_n556__spl_),
    .dinb(new_n624__spl_),
    .dout(new_n626_)
  );


  anb2
  g0562
  (
    .dina(new_n625__spl_),
    .dinb(new_n626_),
    .dout(new_n627_)
  );


  anb1
  g0563
  (
    .dina(new_n555__spl_),
    .dinb(new_n627__spl_),
    .dout(new_n628_)
  );


  anb2
  g0564
  (
    .dina(new_n555__spl_),
    .dinb(new_n627__spl_),
    .dout(new_n629_)
  );


  anb2
  g0565
  (
    .dina(new_n628__spl_),
    .dinb(new_n629_),
    .dout(new_n630_)
  );


  anb1
  g0566
  (
    .dina(new_n554__spl_),
    .dinb(new_n630__spl_),
    .dout(new_n631_)
  );


  anb2
  g0567
  (
    .dina(new_n554__spl_),
    .dinb(new_n630__spl_),
    .dout(new_n632_)
  );


  anb2
  g0568
  (
    .dina(new_n631__spl_),
    .dinb(new_n632_),
    .dout(new_n633_)
  );


  anb1
  g0569
  (
    .dina(new_n553__spl_),
    .dinb(new_n633__spl_),
    .dout(new_n634_)
  );


  anb2
  g0570
  (
    .dina(new_n553__spl_),
    .dinb(new_n633__spl_),
    .dout(new_n635_)
  );


  anb2
  g0571
  (
    .dina(new_n634__spl_),
    .dinb(new_n635_),
    .dout(new_n636_)
  );


  anb1
  g0572
  (
    .dina(new_n552__spl_),
    .dinb(new_n636__spl_),
    .dout(new_n637_)
  );


  anb2
  g0573
  (
    .dina(new_n552__spl_),
    .dinb(new_n636__spl_),
    .dout(new_n638_)
  );


  anb2
  g0574
  (
    .dina(new_n637__spl_),
    .dinb(new_n638_),
    .dout(new_n639_)
  );


  anb1
  g0575
  (
    .dina(new_n551__spl_),
    .dinb(new_n639__spl_),
    .dout(new_n640_)
  );


  anb2
  g0576
  (
    .dina(new_n551__spl_),
    .dinb(new_n639__spl_),
    .dout(new_n641_)
  );


  anb2
  g0577
  (
    .dina(new_n640__spl_),
    .dinb(new_n641_),
    .dout(G6269)
  );


  nor2
  g0578
  (
    .dina(G1_spl_110),
    .dinb(G30_spl_000),
    .dout(new_n643_)
  );


  and2
  g0579
  (
    .dina(new_n637__spl_),
    .dinb(new_n640__spl_),
    .dout(new_n644_)
  );


  nor2
  g0580
  (
    .dina(G2_spl_110),
    .dinb(G29_spl_000),
    .dout(new_n645_)
  );


  and2
  g0581
  (
    .dina(new_n631__spl_),
    .dinb(new_n634__spl_),
    .dout(new_n646_)
  );


  nor2
  g0582
  (
    .dina(G3_spl_101),
    .dinb(G28_spl_001),
    .dout(new_n647_)
  );


  and2
  g0583
  (
    .dina(new_n625__spl_),
    .dinb(new_n628__spl_),
    .dout(new_n648_)
  );


  nor2
  g0584
  (
    .dina(G4_spl_101),
    .dinb(G27_spl_001),
    .dout(new_n649_)
  );


  anb1
  g0585
  (
    .dina(new_n619__spl_),
    .dinb(new_n622__spl_),
    .dout(new_n650_)
  );


  and1
  g0586
  (
    .dina(G5_spl_100),
    .dinb(G26_spl_010),
    .dout(new_n651_)
  );


  anb2
  g0587
  (
    .dina(new_n613__spl_),
    .dinb(new_n616__spl_),
    .dout(new_n652_)
  );


  and1
  g0588
  (
    .dina(G6_spl_100),
    .dinb(G25_spl_010),
    .dout(new_n653_)
  );


  anb2
  g0589
  (
    .dina(new_n607__spl_),
    .dinb(new_n610__spl_),
    .dout(new_n654_)
  );


  and1
  g0590
  (
    .dina(G7_spl_011),
    .dinb(G24_spl_011),
    .dout(new_n655_)
  );


  anb2
  g0591
  (
    .dina(new_n601__spl_),
    .dinb(new_n604__spl_),
    .dout(new_n656_)
  );


  and1
  g0592
  (
    .dina(G8_spl_011),
    .dinb(G23_spl_011),
    .dout(new_n657_)
  );


  anb2
  g0593
  (
    .dina(new_n595__spl_),
    .dinb(new_n598__spl_),
    .dout(new_n658_)
  );


  and1
  g0594
  (
    .dina(G9_spl_010),
    .dinb(G22_spl_100),
    .dout(new_n659_)
  );


  anb2
  g0595
  (
    .dina(new_n589__spl_),
    .dinb(new_n592__spl_),
    .dout(new_n660_)
  );


  and1
  g0596
  (
    .dina(G10_spl_010),
    .dinb(G21_spl_100),
    .dout(new_n661_)
  );


  anb2
  g0597
  (
    .dina(new_n583__spl_),
    .dinb(new_n586__spl_),
    .dout(new_n662_)
  );


  and1
  g0598
  (
    .dina(G11_spl_001),
    .dinb(G20_spl_101),
    .dout(new_n663_)
  );


  anb2
  g0599
  (
    .dina(new_n577__spl_),
    .dinb(new_n580__spl_),
    .dout(new_n664_)
  );


  and1
  g0600
  (
    .dina(G12_spl_001),
    .dinb(G19_spl_101),
    .dout(new_n665_)
  );


  nor2
  g0601
  (
    .dina(G14_spl_000),
    .dinb(G17_spl_110),
    .dout(new_n666_)
  );


  and1
  g0602
  (
    .dina(G13_spl_000),
    .dinb(G18_spl_110),
    .dout(new_n667_)
  );


  anb2
  g0603
  (
    .dina(new_n666__spl_),
    .dinb(new_n667__spl_),
    .dout(new_n668_)
  );


  anb1
  g0604
  (
    .dina(new_n666__spl_),
    .dinb(new_n667__spl_),
    .dout(new_n669_)
  );


  anb1
  g0605
  (
    .dina(new_n668__spl_0),
    .dinb(new_n669_),
    .dout(new_n670_)
  );


  anb1
  g0606
  (
    .dina(new_n574__spl_0),
    .dinb(new_n670__spl_),
    .dout(new_n671_)
  );


  anb2
  g0607
  (
    .dina(new_n574__spl_),
    .dinb(new_n670__spl_),
    .dout(new_n672_)
  );


  nab1
  g0608
  (
    .dina(new_n671__spl_),
    .dinb(new_n672_),
    .dout(new_n673_)
  );


  anb2
  g0609
  (
    .dina(new_n665__spl_),
    .dinb(new_n673__spl_),
    .dout(new_n674_)
  );


  anb1
  g0610
  (
    .dina(new_n665__spl_),
    .dinb(new_n673__spl_),
    .dout(new_n675_)
  );


  nab2
  g0611
  (
    .dina(new_n674__spl_),
    .dinb(new_n675_),
    .dout(new_n676_)
  );


  anb1
  g0612
  (
    .dina(new_n664__spl_),
    .dinb(new_n676__spl_),
    .dout(new_n677_)
  );


  anb2
  g0613
  (
    .dina(new_n664__spl_),
    .dinb(new_n676__spl_),
    .dout(new_n678_)
  );


  nab1
  g0614
  (
    .dina(new_n677__spl_),
    .dinb(new_n678_),
    .dout(new_n679_)
  );


  anb2
  g0615
  (
    .dina(new_n663__spl_),
    .dinb(new_n679__spl_),
    .dout(new_n680_)
  );


  anb1
  g0616
  (
    .dina(new_n663__spl_),
    .dinb(new_n679__spl_),
    .dout(new_n681_)
  );


  nab2
  g0617
  (
    .dina(new_n680__spl_),
    .dinb(new_n681_),
    .dout(new_n682_)
  );


  anb1
  g0618
  (
    .dina(new_n662__spl_),
    .dinb(new_n682__spl_),
    .dout(new_n683_)
  );


  anb2
  g0619
  (
    .dina(new_n662__spl_),
    .dinb(new_n682__spl_),
    .dout(new_n684_)
  );


  nab1
  g0620
  (
    .dina(new_n683__spl_),
    .dinb(new_n684_),
    .dout(new_n685_)
  );


  anb2
  g0621
  (
    .dina(new_n661__spl_),
    .dinb(new_n685__spl_),
    .dout(new_n686_)
  );


  anb1
  g0622
  (
    .dina(new_n661__spl_),
    .dinb(new_n685__spl_),
    .dout(new_n687_)
  );


  nab2
  g0623
  (
    .dina(new_n686__spl_),
    .dinb(new_n687_),
    .dout(new_n688_)
  );


  anb1
  g0624
  (
    .dina(new_n660__spl_),
    .dinb(new_n688__spl_),
    .dout(new_n689_)
  );


  anb2
  g0625
  (
    .dina(new_n660__spl_),
    .dinb(new_n688__spl_),
    .dout(new_n690_)
  );


  nab1
  g0626
  (
    .dina(new_n689__spl_),
    .dinb(new_n690_),
    .dout(new_n691_)
  );


  anb2
  g0627
  (
    .dina(new_n659__spl_),
    .dinb(new_n691__spl_),
    .dout(new_n692_)
  );


  anb1
  g0628
  (
    .dina(new_n659__spl_),
    .dinb(new_n691__spl_),
    .dout(new_n693_)
  );


  nab2
  g0629
  (
    .dina(new_n692__spl_),
    .dinb(new_n693_),
    .dout(new_n694_)
  );


  anb1
  g0630
  (
    .dina(new_n658__spl_),
    .dinb(new_n694__spl_),
    .dout(new_n695_)
  );


  anb2
  g0631
  (
    .dina(new_n658__spl_),
    .dinb(new_n694__spl_),
    .dout(new_n696_)
  );


  nab1
  g0632
  (
    .dina(new_n695__spl_),
    .dinb(new_n696_),
    .dout(new_n697_)
  );


  anb2
  g0633
  (
    .dina(new_n657__spl_),
    .dinb(new_n697__spl_),
    .dout(new_n698_)
  );


  anb1
  g0634
  (
    .dina(new_n657__spl_),
    .dinb(new_n697__spl_),
    .dout(new_n699_)
  );


  nab2
  g0635
  (
    .dina(new_n698__spl_),
    .dinb(new_n699_),
    .dout(new_n700_)
  );


  anb1
  g0636
  (
    .dina(new_n656__spl_),
    .dinb(new_n700__spl_),
    .dout(new_n701_)
  );


  anb2
  g0637
  (
    .dina(new_n656__spl_),
    .dinb(new_n700__spl_),
    .dout(new_n702_)
  );


  nab1
  g0638
  (
    .dina(new_n701__spl_),
    .dinb(new_n702_),
    .dout(new_n703_)
  );


  anb2
  g0639
  (
    .dina(new_n655__spl_),
    .dinb(new_n703__spl_),
    .dout(new_n704_)
  );


  anb1
  g0640
  (
    .dina(new_n655__spl_),
    .dinb(new_n703__spl_),
    .dout(new_n705_)
  );


  nab2
  g0641
  (
    .dina(new_n704__spl_),
    .dinb(new_n705_),
    .dout(new_n706_)
  );


  anb1
  g0642
  (
    .dina(new_n654__spl_),
    .dinb(new_n706__spl_),
    .dout(new_n707_)
  );


  anb2
  g0643
  (
    .dina(new_n654__spl_),
    .dinb(new_n706__spl_),
    .dout(new_n708_)
  );


  nab1
  g0644
  (
    .dina(new_n707__spl_),
    .dinb(new_n708_),
    .dout(new_n709_)
  );


  anb2
  g0645
  (
    .dina(new_n653__spl_),
    .dinb(new_n709__spl_),
    .dout(new_n710_)
  );


  anb1
  g0646
  (
    .dina(new_n653__spl_),
    .dinb(new_n709__spl_),
    .dout(new_n711_)
  );


  nab2
  g0647
  (
    .dina(new_n710__spl_),
    .dinb(new_n711_),
    .dout(new_n712_)
  );


  anb1
  g0648
  (
    .dina(new_n652__spl_),
    .dinb(new_n712__spl_),
    .dout(new_n713_)
  );


  anb2
  g0649
  (
    .dina(new_n652__spl_),
    .dinb(new_n712__spl_),
    .dout(new_n714_)
  );


  nab1
  g0650
  (
    .dina(new_n713__spl_),
    .dinb(new_n714_),
    .dout(new_n715_)
  );


  anb2
  g0651
  (
    .dina(new_n651__spl_),
    .dinb(new_n715__spl_),
    .dout(new_n716_)
  );


  anb1
  g0652
  (
    .dina(new_n651__spl_),
    .dinb(new_n715__spl_),
    .dout(new_n717_)
  );


  anb1
  g0653
  (
    .dina(new_n716__spl_),
    .dinb(new_n717_),
    .dout(new_n718_)
  );


  anb2
  g0654
  (
    .dina(new_n650__spl_),
    .dinb(new_n718__spl_),
    .dout(new_n719_)
  );


  anb1
  g0655
  (
    .dina(new_n650__spl_),
    .dinb(new_n718__spl_),
    .dout(new_n720_)
  );


  nab2
  g0656
  (
    .dina(new_n719__spl_),
    .dinb(new_n720_),
    .dout(new_n721_)
  );


  anb1
  g0657
  (
    .dina(new_n649__spl_),
    .dinb(new_n721__spl_),
    .dout(new_n722_)
  );


  anb2
  g0658
  (
    .dina(new_n649__spl_),
    .dinb(new_n721__spl_),
    .dout(new_n723_)
  );


  anb2
  g0659
  (
    .dina(new_n722__spl_),
    .dinb(new_n723_),
    .dout(new_n724_)
  );


  anb1
  g0660
  (
    .dina(new_n648__spl_),
    .dinb(new_n724__spl_),
    .dout(new_n725_)
  );


  anb2
  g0661
  (
    .dina(new_n648__spl_),
    .dinb(new_n724__spl_),
    .dout(new_n726_)
  );


  anb2
  g0662
  (
    .dina(new_n725__spl_),
    .dinb(new_n726_),
    .dout(new_n727_)
  );


  anb1
  g0663
  (
    .dina(new_n647__spl_),
    .dinb(new_n727__spl_),
    .dout(new_n728_)
  );


  anb2
  g0664
  (
    .dina(new_n647__spl_),
    .dinb(new_n727__spl_),
    .dout(new_n729_)
  );


  anb2
  g0665
  (
    .dina(new_n728__spl_),
    .dinb(new_n729_),
    .dout(new_n730_)
  );


  anb1
  g0666
  (
    .dina(new_n646__spl_),
    .dinb(new_n730__spl_),
    .dout(new_n731_)
  );


  anb2
  g0667
  (
    .dina(new_n646__spl_),
    .dinb(new_n730__spl_),
    .dout(new_n732_)
  );


  anb2
  g0668
  (
    .dina(new_n731__spl_),
    .dinb(new_n732_),
    .dout(new_n733_)
  );


  anb1
  g0669
  (
    .dina(new_n645__spl_),
    .dinb(new_n733__spl_),
    .dout(new_n734_)
  );


  anb2
  g0670
  (
    .dina(new_n645__spl_),
    .dinb(new_n733__spl_),
    .dout(new_n735_)
  );


  anb2
  g0671
  (
    .dina(new_n734__spl_),
    .dinb(new_n735_),
    .dout(new_n736_)
  );


  anb1
  g0672
  (
    .dina(new_n644__spl_),
    .dinb(new_n736__spl_),
    .dout(new_n737_)
  );


  anb2
  g0673
  (
    .dina(new_n644__spl_),
    .dinb(new_n736__spl_),
    .dout(new_n738_)
  );


  anb2
  g0674
  (
    .dina(new_n737__spl_),
    .dinb(new_n738_),
    .dout(new_n739_)
  );


  anb1
  g0675
  (
    .dina(new_n643__spl_),
    .dinb(new_n739__spl_),
    .dout(new_n740_)
  );


  anb2
  g0676
  (
    .dina(new_n643__spl_),
    .dinb(new_n739__spl_),
    .dout(new_n741_)
  );


  anb2
  g0677
  (
    .dina(new_n740__spl_),
    .dinb(new_n741_),
    .dout(G6270)
  );


  nor2
  g0678
  (
    .dina(G1_spl_111),
    .dinb(G31_spl_000),
    .dout(new_n743_)
  );


  and2
  g0679
  (
    .dina(new_n737__spl_),
    .dinb(new_n740__spl_),
    .dout(new_n744_)
  );


  nor2
  g0680
  (
    .dina(G2_spl_110),
    .dinb(G30_spl_000),
    .dout(new_n745_)
  );


  and2
  g0681
  (
    .dina(new_n731__spl_),
    .dinb(new_n734__spl_),
    .dout(new_n746_)
  );


  nor2
  g0682
  (
    .dina(G3_spl_110),
    .dinb(G29_spl_001),
    .dout(new_n747_)
  );


  and2
  g0683
  (
    .dina(new_n725__spl_),
    .dinb(new_n728__spl_),
    .dout(new_n748_)
  );


  nor2
  g0684
  (
    .dina(G4_spl_101),
    .dinb(G28_spl_001),
    .dout(new_n749_)
  );


  anb1
  g0685
  (
    .dina(new_n719__spl_),
    .dinb(new_n722__spl_),
    .dout(new_n750_)
  );


  and1
  g0686
  (
    .dina(G5_spl_101),
    .dinb(G27_spl_010),
    .dout(new_n751_)
  );


  anb2
  g0687
  (
    .dina(new_n713__spl_),
    .dinb(new_n716__spl_),
    .dout(new_n752_)
  );


  and1
  g0688
  (
    .dina(G6_spl_100),
    .dinb(G26_spl_010),
    .dout(new_n753_)
  );


  anb2
  g0689
  (
    .dina(new_n707__spl_),
    .dinb(new_n710__spl_),
    .dout(new_n754_)
  );


  and1
  g0690
  (
    .dina(G7_spl_100),
    .dinb(G25_spl_011),
    .dout(new_n755_)
  );


  anb2
  g0691
  (
    .dina(new_n701__spl_),
    .dinb(new_n704__spl_),
    .dout(new_n756_)
  );


  and1
  g0692
  (
    .dina(G8_spl_011),
    .dinb(G24_spl_011),
    .dout(new_n757_)
  );


  anb2
  g0693
  (
    .dina(new_n695__spl_),
    .dinb(new_n698__spl_),
    .dout(new_n758_)
  );


  and1
  g0694
  (
    .dina(G9_spl_011),
    .dinb(G23_spl_100),
    .dout(new_n759_)
  );


  anb2
  g0695
  (
    .dina(new_n689__spl_),
    .dinb(new_n692__spl_),
    .dout(new_n760_)
  );


  and1
  g0696
  (
    .dina(G10_spl_010),
    .dinb(G22_spl_100),
    .dout(new_n761_)
  );


  anb2
  g0697
  (
    .dina(new_n683__spl_),
    .dinb(new_n686__spl_),
    .dout(new_n762_)
  );


  and1
  g0698
  (
    .dina(G11_spl_010),
    .dinb(G21_spl_101),
    .dout(new_n763_)
  );


  anb2
  g0699
  (
    .dina(new_n677__spl_),
    .dinb(new_n680__spl_),
    .dout(new_n764_)
  );


  and1
  g0700
  (
    .dina(G12_spl_001),
    .dinb(G20_spl_101),
    .dout(new_n765_)
  );


  anb2
  g0701
  (
    .dina(new_n671__spl_),
    .dinb(new_n674__spl_),
    .dout(new_n766_)
  );


  and1
  g0702
  (
    .dina(G13_spl_001),
    .dinb(G19_spl_110),
    .dout(new_n767_)
  );


  nor2
  g0703
  (
    .dina(G15_spl_000),
    .dinb(G17_spl_111),
    .dout(new_n768_)
  );


  and1
  g0704
  (
    .dina(G14_spl_000),
    .dinb(G18_spl_110),
    .dout(new_n769_)
  );


  anb2
  g0705
  (
    .dina(new_n768__spl_),
    .dinb(new_n769__spl_),
    .dout(new_n770_)
  );


  anb1
  g0706
  (
    .dina(new_n768__spl_),
    .dinb(new_n769__spl_),
    .dout(new_n771_)
  );


  anb1
  g0707
  (
    .dina(new_n770__spl_0),
    .dinb(new_n771_),
    .dout(new_n772_)
  );


  anb1
  g0708
  (
    .dina(new_n668__spl_0),
    .dinb(new_n772__spl_),
    .dout(new_n773_)
  );


  anb2
  g0709
  (
    .dina(new_n668__spl_),
    .dinb(new_n772__spl_),
    .dout(new_n774_)
  );


  nab1
  g0710
  (
    .dina(new_n773__spl_),
    .dinb(new_n774_),
    .dout(new_n775_)
  );


  anb2
  g0711
  (
    .dina(new_n767__spl_),
    .dinb(new_n775__spl_),
    .dout(new_n776_)
  );


  anb1
  g0712
  (
    .dina(new_n767__spl_),
    .dinb(new_n775__spl_),
    .dout(new_n777_)
  );


  nab2
  g0713
  (
    .dina(new_n776__spl_),
    .dinb(new_n777_),
    .dout(new_n778_)
  );


  anb1
  g0714
  (
    .dina(new_n766__spl_),
    .dinb(new_n778__spl_),
    .dout(new_n779_)
  );


  anb2
  g0715
  (
    .dina(new_n766__spl_),
    .dinb(new_n778__spl_),
    .dout(new_n780_)
  );


  nab1
  g0716
  (
    .dina(new_n779__spl_),
    .dinb(new_n780_),
    .dout(new_n781_)
  );


  anb2
  g0717
  (
    .dina(new_n765__spl_),
    .dinb(new_n781__spl_),
    .dout(new_n782_)
  );


  anb1
  g0718
  (
    .dina(new_n765__spl_),
    .dinb(new_n781__spl_),
    .dout(new_n783_)
  );


  nab2
  g0719
  (
    .dina(new_n782__spl_),
    .dinb(new_n783_),
    .dout(new_n784_)
  );


  anb1
  g0720
  (
    .dina(new_n764__spl_),
    .dinb(new_n784__spl_),
    .dout(new_n785_)
  );


  anb2
  g0721
  (
    .dina(new_n764__spl_),
    .dinb(new_n784__spl_),
    .dout(new_n786_)
  );


  nab1
  g0722
  (
    .dina(new_n785__spl_),
    .dinb(new_n786_),
    .dout(new_n787_)
  );


  anb2
  g0723
  (
    .dina(new_n763__spl_),
    .dinb(new_n787__spl_),
    .dout(new_n788_)
  );


  anb1
  g0724
  (
    .dina(new_n763__spl_),
    .dinb(new_n787__spl_),
    .dout(new_n789_)
  );


  nab2
  g0725
  (
    .dina(new_n788__spl_),
    .dinb(new_n789_),
    .dout(new_n790_)
  );


  anb1
  g0726
  (
    .dina(new_n762__spl_),
    .dinb(new_n790__spl_),
    .dout(new_n791_)
  );


  anb2
  g0727
  (
    .dina(new_n762__spl_),
    .dinb(new_n790__spl_),
    .dout(new_n792_)
  );


  nab1
  g0728
  (
    .dina(new_n791__spl_),
    .dinb(new_n792_),
    .dout(new_n793_)
  );


  anb2
  g0729
  (
    .dina(new_n761__spl_),
    .dinb(new_n793__spl_),
    .dout(new_n794_)
  );


  anb1
  g0730
  (
    .dina(new_n761__spl_),
    .dinb(new_n793__spl_),
    .dout(new_n795_)
  );


  nab2
  g0731
  (
    .dina(new_n794__spl_),
    .dinb(new_n795_),
    .dout(new_n796_)
  );


  anb1
  g0732
  (
    .dina(new_n760__spl_),
    .dinb(new_n796__spl_),
    .dout(new_n797_)
  );


  anb2
  g0733
  (
    .dina(new_n760__spl_),
    .dinb(new_n796__spl_),
    .dout(new_n798_)
  );


  nab1
  g0734
  (
    .dina(new_n797__spl_),
    .dinb(new_n798_),
    .dout(new_n799_)
  );


  anb2
  g0735
  (
    .dina(new_n759__spl_),
    .dinb(new_n799__spl_),
    .dout(new_n800_)
  );


  anb1
  g0736
  (
    .dina(new_n759__spl_),
    .dinb(new_n799__spl_),
    .dout(new_n801_)
  );


  nab2
  g0737
  (
    .dina(new_n800__spl_),
    .dinb(new_n801_),
    .dout(new_n802_)
  );


  anb1
  g0738
  (
    .dina(new_n758__spl_),
    .dinb(new_n802__spl_),
    .dout(new_n803_)
  );


  anb2
  g0739
  (
    .dina(new_n758__spl_),
    .dinb(new_n802__spl_),
    .dout(new_n804_)
  );


  nab1
  g0740
  (
    .dina(new_n803__spl_),
    .dinb(new_n804_),
    .dout(new_n805_)
  );


  anb2
  g0741
  (
    .dina(new_n757__spl_),
    .dinb(new_n805__spl_),
    .dout(new_n806_)
  );


  anb1
  g0742
  (
    .dina(new_n757__spl_),
    .dinb(new_n805__spl_),
    .dout(new_n807_)
  );


  nab2
  g0743
  (
    .dina(new_n806__spl_),
    .dinb(new_n807_),
    .dout(new_n808_)
  );


  anb1
  g0744
  (
    .dina(new_n756__spl_),
    .dinb(new_n808__spl_),
    .dout(new_n809_)
  );


  anb2
  g0745
  (
    .dina(new_n756__spl_),
    .dinb(new_n808__spl_),
    .dout(new_n810_)
  );


  nab1
  g0746
  (
    .dina(new_n809__spl_),
    .dinb(new_n810_),
    .dout(new_n811_)
  );


  anb2
  g0747
  (
    .dina(new_n755__spl_),
    .dinb(new_n811__spl_),
    .dout(new_n812_)
  );


  anb1
  g0748
  (
    .dina(new_n755__spl_),
    .dinb(new_n811__spl_),
    .dout(new_n813_)
  );


  nab2
  g0749
  (
    .dina(new_n812__spl_),
    .dinb(new_n813_),
    .dout(new_n814_)
  );


  anb1
  g0750
  (
    .dina(new_n754__spl_),
    .dinb(new_n814__spl_),
    .dout(new_n815_)
  );


  anb2
  g0751
  (
    .dina(new_n754__spl_),
    .dinb(new_n814__spl_),
    .dout(new_n816_)
  );


  nab1
  g0752
  (
    .dina(new_n815__spl_),
    .dinb(new_n816_),
    .dout(new_n817_)
  );


  anb2
  g0753
  (
    .dina(new_n753__spl_),
    .dinb(new_n817__spl_),
    .dout(new_n818_)
  );


  anb1
  g0754
  (
    .dina(new_n753__spl_),
    .dinb(new_n817__spl_),
    .dout(new_n819_)
  );


  nab2
  g0755
  (
    .dina(new_n818__spl_),
    .dinb(new_n819_),
    .dout(new_n820_)
  );


  anb1
  g0756
  (
    .dina(new_n752__spl_),
    .dinb(new_n820__spl_),
    .dout(new_n821_)
  );


  anb2
  g0757
  (
    .dina(new_n752__spl_),
    .dinb(new_n820__spl_),
    .dout(new_n822_)
  );


  nab1
  g0758
  (
    .dina(new_n821__spl_),
    .dinb(new_n822_),
    .dout(new_n823_)
  );


  anb2
  g0759
  (
    .dina(new_n751__spl_),
    .dinb(new_n823__spl_),
    .dout(new_n824_)
  );


  anb1
  g0760
  (
    .dina(new_n751__spl_),
    .dinb(new_n823__spl_),
    .dout(new_n825_)
  );


  anb1
  g0761
  (
    .dina(new_n824__spl_),
    .dinb(new_n825_),
    .dout(new_n826_)
  );


  anb2
  g0762
  (
    .dina(new_n750__spl_),
    .dinb(new_n826__spl_),
    .dout(new_n827_)
  );


  anb1
  g0763
  (
    .dina(new_n750__spl_),
    .dinb(new_n826__spl_),
    .dout(new_n828_)
  );


  nab2
  g0764
  (
    .dina(new_n827__spl_),
    .dinb(new_n828_),
    .dout(new_n829_)
  );


  anb1
  g0765
  (
    .dina(new_n749__spl_),
    .dinb(new_n829__spl_),
    .dout(new_n830_)
  );


  anb2
  g0766
  (
    .dina(new_n749__spl_),
    .dinb(new_n829__spl_),
    .dout(new_n831_)
  );


  anb2
  g0767
  (
    .dina(new_n830__spl_),
    .dinb(new_n831_),
    .dout(new_n832_)
  );


  anb1
  g0768
  (
    .dina(new_n748__spl_),
    .dinb(new_n832__spl_),
    .dout(new_n833_)
  );


  anb2
  g0769
  (
    .dina(new_n748__spl_),
    .dinb(new_n832__spl_),
    .dout(new_n834_)
  );


  anb2
  g0770
  (
    .dina(new_n833__spl_),
    .dinb(new_n834_),
    .dout(new_n835_)
  );


  anb1
  g0771
  (
    .dina(new_n747__spl_),
    .dinb(new_n835__spl_),
    .dout(new_n836_)
  );


  anb2
  g0772
  (
    .dina(new_n747__spl_),
    .dinb(new_n835__spl_),
    .dout(new_n837_)
  );


  anb2
  g0773
  (
    .dina(new_n836__spl_),
    .dinb(new_n837_),
    .dout(new_n838_)
  );


  anb1
  g0774
  (
    .dina(new_n746__spl_),
    .dinb(new_n838__spl_),
    .dout(new_n839_)
  );


  anb2
  g0775
  (
    .dina(new_n746__spl_),
    .dinb(new_n838__spl_),
    .dout(new_n840_)
  );


  anb2
  g0776
  (
    .dina(new_n839__spl_),
    .dinb(new_n840_),
    .dout(new_n841_)
  );


  anb1
  g0777
  (
    .dina(new_n745__spl_),
    .dinb(new_n841__spl_),
    .dout(new_n842_)
  );


  anb2
  g0778
  (
    .dina(new_n745__spl_),
    .dinb(new_n841__spl_),
    .dout(new_n843_)
  );


  anb2
  g0779
  (
    .dina(new_n842__spl_),
    .dinb(new_n843_),
    .dout(new_n844_)
  );


  anb1
  g0780
  (
    .dina(new_n744__spl_),
    .dinb(new_n844__spl_),
    .dout(new_n845_)
  );


  anb2
  g0781
  (
    .dina(new_n744__spl_),
    .dinb(new_n844__spl_),
    .dout(new_n846_)
  );


  anb2
  g0782
  (
    .dina(new_n845__spl_),
    .dinb(new_n846_),
    .dout(new_n847_)
  );


  anb1
  g0783
  (
    .dina(new_n743__spl_),
    .dinb(new_n847__spl_),
    .dout(new_n848_)
  );


  anb2
  g0784
  (
    .dina(new_n743__spl_),
    .dinb(new_n847__spl_),
    .dout(new_n849_)
  );


  anb2
  g0785
  (
    .dina(new_n848__spl_),
    .dinb(new_n849_),
    .dout(G6271)
  );


  nor2
  g0786
  (
    .dina(G1_spl_111),
    .dinb(G32_spl_000),
    .dout(new_n851_)
  );


  and2
  g0787
  (
    .dina(new_n845__spl_),
    .dinb(new_n848__spl_),
    .dout(new_n852_)
  );


  nor2
  g0788
  (
    .dina(G2_spl_111),
    .dinb(G31_spl_000),
    .dout(new_n853_)
  );


  and2
  g0789
  (
    .dina(new_n839__spl_),
    .dinb(new_n842__spl_),
    .dout(new_n854_)
  );


  nor2
  g0790
  (
    .dina(G3_spl_110),
    .dinb(G30_spl_001),
    .dout(new_n855_)
  );


  and2
  g0791
  (
    .dina(new_n833__spl_),
    .dinb(new_n836__spl_),
    .dout(new_n856_)
  );


  nor2
  g0792
  (
    .dina(G4_spl_110),
    .dinb(G29_spl_001),
    .dout(new_n857_)
  );


  anb1
  g0793
  (
    .dina(new_n827__spl_),
    .dinb(new_n830__spl_),
    .dout(new_n858_)
  );


  and1
  g0794
  (
    .dina(G5_spl_101),
    .dinb(G28_spl_010),
    .dout(new_n859_)
  );


  anb2
  g0795
  (
    .dina(new_n821__spl_),
    .dinb(new_n824__spl_),
    .dout(new_n860_)
  );


  and1
  g0796
  (
    .dina(G6_spl_101),
    .dinb(G27_spl_010),
    .dout(new_n861_)
  );


  anb2
  g0797
  (
    .dina(new_n815__spl_),
    .dinb(new_n818__spl_),
    .dout(new_n862_)
  );


  and1
  g0798
  (
    .dina(G7_spl_100),
    .dinb(G26_spl_011),
    .dout(new_n863_)
  );


  anb2
  g0799
  (
    .dina(new_n809__spl_),
    .dinb(new_n812__spl_),
    .dout(new_n864_)
  );


  and1
  g0800
  (
    .dina(G8_spl_100),
    .dinb(G25_spl_011),
    .dout(new_n865_)
  );


  anb2
  g0801
  (
    .dina(new_n803__spl_),
    .dinb(new_n806__spl_),
    .dout(new_n866_)
  );


  and1
  g0802
  (
    .dina(G9_spl_011),
    .dinb(G24_spl_100),
    .dout(new_n867_)
  );


  anb2
  g0803
  (
    .dina(new_n797__spl_),
    .dinb(new_n800__spl_),
    .dout(new_n868_)
  );


  and1
  g0804
  (
    .dina(G10_spl_011),
    .dinb(G23_spl_100),
    .dout(new_n869_)
  );


  anb2
  g0805
  (
    .dina(new_n791__spl_),
    .dinb(new_n794__spl_),
    .dout(new_n870_)
  );


  and1
  g0806
  (
    .dina(G11_spl_010),
    .dinb(G22_spl_101),
    .dout(new_n871_)
  );


  anb2
  g0807
  (
    .dina(new_n785__spl_),
    .dinb(new_n788__spl_),
    .dout(new_n872_)
  );


  and1
  g0808
  (
    .dina(G12_spl_010),
    .dinb(G21_spl_101),
    .dout(new_n873_)
  );


  anb2
  g0809
  (
    .dina(new_n779__spl_),
    .dinb(new_n782__spl_),
    .dout(new_n874_)
  );


  and1
  g0810
  (
    .dina(G13_spl_001),
    .dinb(G20_spl_110),
    .dout(new_n875_)
  );


  anb2
  g0811
  (
    .dina(new_n773__spl_),
    .dinb(new_n776__spl_),
    .dout(new_n876_)
  );


  and1
  g0812
  (
    .dina(G14_spl_001),
    .dinb(G19_spl_110),
    .dout(new_n877_)
  );


  and1
  g0813
  (
    .dina(G16_spl_000),
    .dinb(G17_spl_111),
    .dout(new_n878_)
  );


  nor2
  g0814
  (
    .dina(G15_spl_000),
    .dinb(G18_spl_111),
    .dout(new_n879_)
  );


  anb1
  g0815
  (
    .dina(new_n878__spl_),
    .dinb(new_n879__spl_),
    .dout(new_n880_)
  );


  anb2
  g0816
  (
    .dina(new_n878__spl_),
    .dinb(new_n879__spl_),
    .dout(new_n881_)
  );


  nab1
  g0817
  (
    .dina(new_n880__spl_),
    .dinb(new_n881_),
    .dout(new_n882_)
  );


  anb1
  g0818
  (
    .dina(new_n770__spl_0),
    .dinb(new_n882__spl_),
    .dout(new_n883_)
  );


  anb2
  g0819
  (
    .dina(new_n770__spl_),
    .dinb(new_n882__spl_),
    .dout(new_n884_)
  );


  nab1
  g0820
  (
    .dina(new_n883__spl_),
    .dinb(new_n884_),
    .dout(new_n885_)
  );


  anb2
  g0821
  (
    .dina(new_n877__spl_),
    .dinb(new_n885__spl_),
    .dout(new_n886_)
  );


  anb1
  g0822
  (
    .dina(new_n877__spl_),
    .dinb(new_n885__spl_),
    .dout(new_n887_)
  );


  nab2
  g0823
  (
    .dina(new_n886__spl_),
    .dinb(new_n887_),
    .dout(new_n888_)
  );


  anb1
  g0824
  (
    .dina(new_n876__spl_),
    .dinb(new_n888__spl_),
    .dout(new_n889_)
  );


  anb2
  g0825
  (
    .dina(new_n876__spl_),
    .dinb(new_n888__spl_),
    .dout(new_n890_)
  );


  nab1
  g0826
  (
    .dina(new_n889__spl_),
    .dinb(new_n890_),
    .dout(new_n891_)
  );


  anb2
  g0827
  (
    .dina(new_n875__spl_),
    .dinb(new_n891__spl_),
    .dout(new_n892_)
  );


  anb1
  g0828
  (
    .dina(new_n875__spl_),
    .dinb(new_n891__spl_),
    .dout(new_n893_)
  );


  nab2
  g0829
  (
    .dina(new_n892__spl_),
    .dinb(new_n893_),
    .dout(new_n894_)
  );


  anb1
  g0830
  (
    .dina(new_n874__spl_),
    .dinb(new_n894__spl_),
    .dout(new_n895_)
  );


  anb2
  g0831
  (
    .dina(new_n874__spl_),
    .dinb(new_n894__spl_),
    .dout(new_n896_)
  );


  nab1
  g0832
  (
    .dina(new_n895__spl_),
    .dinb(new_n896_),
    .dout(new_n897_)
  );


  anb2
  g0833
  (
    .dina(new_n873__spl_),
    .dinb(new_n897__spl_),
    .dout(new_n898_)
  );


  anb1
  g0834
  (
    .dina(new_n873__spl_),
    .dinb(new_n897__spl_),
    .dout(new_n899_)
  );


  nab2
  g0835
  (
    .dina(new_n898__spl_),
    .dinb(new_n899_),
    .dout(new_n900_)
  );


  anb1
  g0836
  (
    .dina(new_n872__spl_),
    .dinb(new_n900__spl_),
    .dout(new_n901_)
  );


  anb2
  g0837
  (
    .dina(new_n872__spl_),
    .dinb(new_n900__spl_),
    .dout(new_n902_)
  );


  nab1
  g0838
  (
    .dina(new_n901__spl_),
    .dinb(new_n902_),
    .dout(new_n903_)
  );


  anb2
  g0839
  (
    .dina(new_n871__spl_),
    .dinb(new_n903__spl_),
    .dout(new_n904_)
  );


  anb1
  g0840
  (
    .dina(new_n871__spl_),
    .dinb(new_n903__spl_),
    .dout(new_n905_)
  );


  nab2
  g0841
  (
    .dina(new_n904__spl_),
    .dinb(new_n905_),
    .dout(new_n906_)
  );


  anb1
  g0842
  (
    .dina(new_n870__spl_),
    .dinb(new_n906__spl_),
    .dout(new_n907_)
  );


  anb2
  g0843
  (
    .dina(new_n870__spl_),
    .dinb(new_n906__spl_),
    .dout(new_n908_)
  );


  nab1
  g0844
  (
    .dina(new_n907__spl_),
    .dinb(new_n908_),
    .dout(new_n909_)
  );


  anb2
  g0845
  (
    .dina(new_n869__spl_),
    .dinb(new_n909__spl_),
    .dout(new_n910_)
  );


  anb1
  g0846
  (
    .dina(new_n869__spl_),
    .dinb(new_n909__spl_),
    .dout(new_n911_)
  );


  nab2
  g0847
  (
    .dina(new_n910__spl_),
    .dinb(new_n911_),
    .dout(new_n912_)
  );


  anb1
  g0848
  (
    .dina(new_n868__spl_),
    .dinb(new_n912__spl_),
    .dout(new_n913_)
  );


  anb2
  g0849
  (
    .dina(new_n868__spl_),
    .dinb(new_n912__spl_),
    .dout(new_n914_)
  );


  nab1
  g0850
  (
    .dina(new_n913__spl_),
    .dinb(new_n914_),
    .dout(new_n915_)
  );


  anb2
  g0851
  (
    .dina(new_n867__spl_),
    .dinb(new_n915__spl_),
    .dout(new_n916_)
  );


  anb1
  g0852
  (
    .dina(new_n867__spl_),
    .dinb(new_n915__spl_),
    .dout(new_n917_)
  );


  nab2
  g0853
  (
    .dina(new_n916__spl_),
    .dinb(new_n917_),
    .dout(new_n918_)
  );


  anb1
  g0854
  (
    .dina(new_n866__spl_),
    .dinb(new_n918__spl_),
    .dout(new_n919_)
  );


  anb2
  g0855
  (
    .dina(new_n866__spl_),
    .dinb(new_n918__spl_),
    .dout(new_n920_)
  );


  nab1
  g0856
  (
    .dina(new_n919__spl_),
    .dinb(new_n920_),
    .dout(new_n921_)
  );


  anb2
  g0857
  (
    .dina(new_n865__spl_),
    .dinb(new_n921__spl_),
    .dout(new_n922_)
  );


  anb1
  g0858
  (
    .dina(new_n865__spl_),
    .dinb(new_n921__spl_),
    .dout(new_n923_)
  );


  nab2
  g0859
  (
    .dina(new_n922__spl_),
    .dinb(new_n923_),
    .dout(new_n924_)
  );


  anb1
  g0860
  (
    .dina(new_n864__spl_),
    .dinb(new_n924__spl_),
    .dout(new_n925_)
  );


  anb2
  g0861
  (
    .dina(new_n864__spl_),
    .dinb(new_n924__spl_),
    .dout(new_n926_)
  );


  nab1
  g0862
  (
    .dina(new_n925__spl_),
    .dinb(new_n926_),
    .dout(new_n927_)
  );


  anb2
  g0863
  (
    .dina(new_n863__spl_),
    .dinb(new_n927__spl_),
    .dout(new_n928_)
  );


  anb1
  g0864
  (
    .dina(new_n863__spl_),
    .dinb(new_n927__spl_),
    .dout(new_n929_)
  );


  nab2
  g0865
  (
    .dina(new_n928__spl_),
    .dinb(new_n929_),
    .dout(new_n930_)
  );


  anb1
  g0866
  (
    .dina(new_n862__spl_),
    .dinb(new_n930__spl_),
    .dout(new_n931_)
  );


  anb2
  g0867
  (
    .dina(new_n862__spl_),
    .dinb(new_n930__spl_),
    .dout(new_n932_)
  );


  nab1
  g0868
  (
    .dina(new_n931__spl_),
    .dinb(new_n932_),
    .dout(new_n933_)
  );


  anb2
  g0869
  (
    .dina(new_n861__spl_),
    .dinb(new_n933__spl_),
    .dout(new_n934_)
  );


  anb1
  g0870
  (
    .dina(new_n861__spl_),
    .dinb(new_n933__spl_),
    .dout(new_n935_)
  );


  nab2
  g0871
  (
    .dina(new_n934__spl_),
    .dinb(new_n935_),
    .dout(new_n936_)
  );


  anb1
  g0872
  (
    .dina(new_n860__spl_),
    .dinb(new_n936__spl_),
    .dout(new_n937_)
  );


  anb2
  g0873
  (
    .dina(new_n860__spl_),
    .dinb(new_n936__spl_),
    .dout(new_n938_)
  );


  nab1
  g0874
  (
    .dina(new_n937__spl_),
    .dinb(new_n938_),
    .dout(new_n939_)
  );


  anb2
  g0875
  (
    .dina(new_n859__spl_),
    .dinb(new_n939__spl_),
    .dout(new_n940_)
  );


  anb1
  g0876
  (
    .dina(new_n859__spl_),
    .dinb(new_n939__spl_),
    .dout(new_n941_)
  );


  anb1
  g0877
  (
    .dina(new_n940__spl_),
    .dinb(new_n941_),
    .dout(new_n942_)
  );


  anb2
  g0878
  (
    .dina(new_n858__spl_),
    .dinb(new_n942__spl_),
    .dout(new_n943_)
  );


  anb1
  g0879
  (
    .dina(new_n858__spl_),
    .dinb(new_n942__spl_),
    .dout(new_n944_)
  );


  nab2
  g0880
  (
    .dina(new_n943__spl_),
    .dinb(new_n944_),
    .dout(new_n945_)
  );


  anb1
  g0881
  (
    .dina(new_n857__spl_),
    .dinb(new_n945__spl_),
    .dout(new_n946_)
  );


  anb2
  g0882
  (
    .dina(new_n857__spl_),
    .dinb(new_n945__spl_),
    .dout(new_n947_)
  );


  anb2
  g0883
  (
    .dina(new_n946__spl_),
    .dinb(new_n947_),
    .dout(new_n948_)
  );


  anb1
  g0884
  (
    .dina(new_n856__spl_),
    .dinb(new_n948__spl_),
    .dout(new_n949_)
  );


  anb2
  g0885
  (
    .dina(new_n856__spl_),
    .dinb(new_n948__spl_),
    .dout(new_n950_)
  );


  anb2
  g0886
  (
    .dina(new_n949__spl_),
    .dinb(new_n950_),
    .dout(new_n951_)
  );


  anb1
  g0887
  (
    .dina(new_n855__spl_),
    .dinb(new_n951__spl_),
    .dout(new_n952_)
  );


  anb2
  g0888
  (
    .dina(new_n855__spl_),
    .dinb(new_n951__spl_),
    .dout(new_n953_)
  );


  anb2
  g0889
  (
    .dina(new_n952__spl_),
    .dinb(new_n953_),
    .dout(new_n954_)
  );


  anb1
  g0890
  (
    .dina(new_n854__spl_),
    .dinb(new_n954__spl_),
    .dout(new_n955_)
  );


  anb2
  g0891
  (
    .dina(new_n854__spl_),
    .dinb(new_n954__spl_),
    .dout(new_n956_)
  );


  anb2
  g0892
  (
    .dina(new_n955__spl_),
    .dinb(new_n956_),
    .dout(new_n957_)
  );


  anb1
  g0893
  (
    .dina(new_n853__spl_),
    .dinb(new_n957__spl_),
    .dout(new_n958_)
  );


  anb2
  g0894
  (
    .dina(new_n853__spl_),
    .dinb(new_n957__spl_),
    .dout(new_n959_)
  );


  anb2
  g0895
  (
    .dina(new_n958__spl_),
    .dinb(new_n959_),
    .dout(new_n960_)
  );


  anb1
  g0896
  (
    .dina(new_n852__spl_),
    .dinb(new_n960__spl_),
    .dout(new_n961_)
  );


  anb2
  g0897
  (
    .dina(new_n852__spl_),
    .dinb(new_n960__spl_),
    .dout(new_n962_)
  );


  anb2
  g0898
  (
    .dina(new_n961__spl_),
    .dinb(new_n962_),
    .dout(new_n963_)
  );


  anb1
  g0899
  (
    .dina(new_n851__spl_),
    .dinb(new_n963__spl_),
    .dout(new_n964_)
  );


  anb2
  g0900
  (
    .dina(new_n851__spl_),
    .dinb(new_n963__spl_),
    .dout(new_n965_)
  );


  anb2
  g0901
  (
    .dina(new_n964__spl_),
    .dinb(new_n965_),
    .dout(G6272)
  );


  nor1
  g0902
  (
    .dina(new_n961__spl_),
    .dinb(new_n964__spl_),
    .dout(new_n967_)
  );


  and1
  g0903
  (
    .dina(G2_spl_111),
    .dinb(G32_spl_000),
    .dout(new_n968_)
  );


  nor1
  g0904
  (
    .dina(new_n955__spl_),
    .dinb(new_n958__spl_),
    .dout(new_n969_)
  );


  and1
  g0905
  (
    .dina(G3_spl_111),
    .dinb(G31_spl_001),
    .dout(new_n970_)
  );


  nor1
  g0906
  (
    .dina(new_n949__spl_),
    .dinb(new_n952__spl_),
    .dout(new_n971_)
  );


  and1
  g0907
  (
    .dina(G4_spl_110),
    .dinb(G30_spl_001),
    .dout(new_n972_)
  );


  anb1
  g0908
  (
    .dina(new_n943__spl_),
    .dinb(new_n946__spl_),
    .dout(new_n973_)
  );


  and1
  g0909
  (
    .dina(G5_spl_110),
    .dinb(G29_spl_010),
    .dout(new_n974_)
  );


  anb2
  g0910
  (
    .dina(new_n937__spl_),
    .dinb(new_n940__spl_),
    .dout(new_n975_)
  );


  and1
  g0911
  (
    .dina(G6_spl_101),
    .dinb(G28_spl_010),
    .dout(new_n976_)
  );


  anb2
  g0912
  (
    .dina(new_n931__spl_),
    .dinb(new_n934__spl_),
    .dout(new_n977_)
  );


  and1
  g0913
  (
    .dina(G7_spl_101),
    .dinb(G27_spl_011),
    .dout(new_n978_)
  );


  anb2
  g0914
  (
    .dina(new_n925__spl_),
    .dinb(new_n928__spl_),
    .dout(new_n979_)
  );


  and1
  g0915
  (
    .dina(G8_spl_100),
    .dinb(G26_spl_011),
    .dout(new_n980_)
  );


  anb2
  g0916
  (
    .dina(new_n919__spl_),
    .dinb(new_n922__spl_),
    .dout(new_n981_)
  );


  and1
  g0917
  (
    .dina(G9_spl_100),
    .dinb(G25_spl_100),
    .dout(new_n982_)
  );


  anb2
  g0918
  (
    .dina(new_n913__spl_),
    .dinb(new_n916__spl_),
    .dout(new_n983_)
  );


  and1
  g0919
  (
    .dina(G10_spl_011),
    .dinb(G24_spl_100),
    .dout(new_n984_)
  );


  anb2
  g0920
  (
    .dina(new_n907__spl_),
    .dinb(new_n910__spl_),
    .dout(new_n985_)
  );


  and1
  g0921
  (
    .dina(G11_spl_011),
    .dinb(G23_spl_101),
    .dout(new_n986_)
  );


  anb2
  g0922
  (
    .dina(new_n901__spl_),
    .dinb(new_n904__spl_),
    .dout(new_n987_)
  );


  and1
  g0923
  (
    .dina(G12_spl_010),
    .dinb(G22_spl_101),
    .dout(new_n988_)
  );


  anb2
  g0924
  (
    .dina(new_n895__spl_),
    .dinb(new_n898__spl_),
    .dout(new_n989_)
  );


  and1
  g0925
  (
    .dina(G13_spl_010),
    .dinb(G21_spl_110),
    .dout(new_n990_)
  );


  anb2
  g0926
  (
    .dina(new_n889__spl_),
    .dinb(new_n892__spl_),
    .dout(new_n991_)
  );


  and1
  g0927
  (
    .dina(G14_spl_001),
    .dinb(G20_spl_110),
    .dout(new_n992_)
  );


  anb2
  g0928
  (
    .dina(new_n883__spl_),
    .dinb(new_n886__spl_),
    .dout(new_n993_)
  );


  and1
  g0929
  (
    .dina(G16_spl_000),
    .dinb(G18_spl_111),
    .dout(new_n994_)
  );


  anb1
  g0930
  (
    .dina(new_n994__spl_),
    .dinb(new_n880__spl_),
    .dout(new_n995_)
  );


  and1
  g0931
  (
    .dina(G15_spl_001),
    .dinb(G19_spl_111),
    .dout(new_n996_)
  );


  anb1
  g0932
  (
    .dina(new_n995__spl_),
    .dinb(new_n996__spl_),
    .dout(new_n997_)
  );


  anb2
  g0933
  (
    .dina(new_n995__spl_),
    .dinb(new_n996__spl_),
    .dout(new_n998_)
  );


  anb2
  g0934
  (
    .dina(new_n997__spl_),
    .dinb(new_n998_),
    .dout(new_n999_)
  );


  anb1
  g0935
  (
    .dina(new_n993__spl_),
    .dinb(new_n999__spl_),
    .dout(new_n1000_)
  );


  anb2
  g0936
  (
    .dina(new_n993__spl_),
    .dinb(new_n999__spl_),
    .dout(new_n1001_)
  );


  nab1
  g0937
  (
    .dina(new_n1000__spl_),
    .dinb(new_n1001_),
    .dout(new_n1002_)
  );


  anb2
  g0938
  (
    .dina(new_n992__spl_),
    .dinb(new_n1002__spl_),
    .dout(new_n1003_)
  );


  anb1
  g0939
  (
    .dina(new_n992__spl_),
    .dinb(new_n1002__spl_),
    .dout(new_n1004_)
  );


  nab2
  g0940
  (
    .dina(new_n1003__spl_),
    .dinb(new_n1004_),
    .dout(new_n1005_)
  );


  anb1
  g0941
  (
    .dina(new_n991__spl_),
    .dinb(new_n1005__spl_),
    .dout(new_n1006_)
  );


  anb2
  g0942
  (
    .dina(new_n991__spl_),
    .dinb(new_n1005__spl_),
    .dout(new_n1007_)
  );


  nab1
  g0943
  (
    .dina(new_n1006__spl_),
    .dinb(new_n1007_),
    .dout(new_n1008_)
  );


  anb2
  g0944
  (
    .dina(new_n990__spl_),
    .dinb(new_n1008__spl_),
    .dout(new_n1009_)
  );


  anb1
  g0945
  (
    .dina(new_n990__spl_),
    .dinb(new_n1008__spl_),
    .dout(new_n1010_)
  );


  nab2
  g0946
  (
    .dina(new_n1009__spl_),
    .dinb(new_n1010_),
    .dout(new_n1011_)
  );


  anb1
  g0947
  (
    .dina(new_n989__spl_),
    .dinb(new_n1011__spl_),
    .dout(new_n1012_)
  );


  anb2
  g0948
  (
    .dina(new_n989__spl_),
    .dinb(new_n1011__spl_),
    .dout(new_n1013_)
  );


  nab1
  g0949
  (
    .dina(new_n1012__spl_),
    .dinb(new_n1013_),
    .dout(new_n1014_)
  );


  anb2
  g0950
  (
    .dina(new_n988__spl_),
    .dinb(new_n1014__spl_),
    .dout(new_n1015_)
  );


  anb1
  g0951
  (
    .dina(new_n988__spl_),
    .dinb(new_n1014__spl_),
    .dout(new_n1016_)
  );


  nab2
  g0952
  (
    .dina(new_n1015__spl_),
    .dinb(new_n1016_),
    .dout(new_n1017_)
  );


  anb1
  g0953
  (
    .dina(new_n987__spl_),
    .dinb(new_n1017__spl_),
    .dout(new_n1018_)
  );


  anb2
  g0954
  (
    .dina(new_n987__spl_),
    .dinb(new_n1017__spl_),
    .dout(new_n1019_)
  );


  nab1
  g0955
  (
    .dina(new_n1018__spl_),
    .dinb(new_n1019_),
    .dout(new_n1020_)
  );


  anb2
  g0956
  (
    .dina(new_n986__spl_),
    .dinb(new_n1020__spl_),
    .dout(new_n1021_)
  );


  anb1
  g0957
  (
    .dina(new_n986__spl_),
    .dinb(new_n1020__spl_),
    .dout(new_n1022_)
  );


  nab2
  g0958
  (
    .dina(new_n1021__spl_),
    .dinb(new_n1022_),
    .dout(new_n1023_)
  );


  anb1
  g0959
  (
    .dina(new_n985__spl_),
    .dinb(new_n1023__spl_),
    .dout(new_n1024_)
  );


  anb2
  g0960
  (
    .dina(new_n985__spl_),
    .dinb(new_n1023__spl_),
    .dout(new_n1025_)
  );


  nab1
  g0961
  (
    .dina(new_n1024__spl_),
    .dinb(new_n1025_),
    .dout(new_n1026_)
  );


  anb2
  g0962
  (
    .dina(new_n984__spl_),
    .dinb(new_n1026__spl_),
    .dout(new_n1027_)
  );


  anb1
  g0963
  (
    .dina(new_n984__spl_),
    .dinb(new_n1026__spl_),
    .dout(new_n1028_)
  );


  nab2
  g0964
  (
    .dina(new_n1027__spl_),
    .dinb(new_n1028_),
    .dout(new_n1029_)
  );


  anb1
  g0965
  (
    .dina(new_n983__spl_),
    .dinb(new_n1029__spl_),
    .dout(new_n1030_)
  );


  anb2
  g0966
  (
    .dina(new_n983__spl_),
    .dinb(new_n1029__spl_),
    .dout(new_n1031_)
  );


  nab1
  g0967
  (
    .dina(new_n1030__spl_),
    .dinb(new_n1031_),
    .dout(new_n1032_)
  );


  anb2
  g0968
  (
    .dina(new_n982__spl_),
    .dinb(new_n1032__spl_),
    .dout(new_n1033_)
  );


  anb1
  g0969
  (
    .dina(new_n982__spl_),
    .dinb(new_n1032__spl_),
    .dout(new_n1034_)
  );


  nab2
  g0970
  (
    .dina(new_n1033__spl_),
    .dinb(new_n1034_),
    .dout(new_n1035_)
  );


  anb1
  g0971
  (
    .dina(new_n981__spl_),
    .dinb(new_n1035__spl_),
    .dout(new_n1036_)
  );


  anb2
  g0972
  (
    .dina(new_n981__spl_),
    .dinb(new_n1035__spl_),
    .dout(new_n1037_)
  );


  nab1
  g0973
  (
    .dina(new_n1036__spl_),
    .dinb(new_n1037_),
    .dout(new_n1038_)
  );


  anb2
  g0974
  (
    .dina(new_n980__spl_),
    .dinb(new_n1038__spl_),
    .dout(new_n1039_)
  );


  anb1
  g0975
  (
    .dina(new_n980__spl_),
    .dinb(new_n1038__spl_),
    .dout(new_n1040_)
  );


  nab2
  g0976
  (
    .dina(new_n1039__spl_),
    .dinb(new_n1040_),
    .dout(new_n1041_)
  );


  anb1
  g0977
  (
    .dina(new_n979__spl_),
    .dinb(new_n1041__spl_),
    .dout(new_n1042_)
  );


  anb2
  g0978
  (
    .dina(new_n979__spl_),
    .dinb(new_n1041__spl_),
    .dout(new_n1043_)
  );


  nab1
  g0979
  (
    .dina(new_n1042__spl_),
    .dinb(new_n1043_),
    .dout(new_n1044_)
  );


  anb2
  g0980
  (
    .dina(new_n978__spl_),
    .dinb(new_n1044__spl_),
    .dout(new_n1045_)
  );


  anb1
  g0981
  (
    .dina(new_n978__spl_),
    .dinb(new_n1044__spl_),
    .dout(new_n1046_)
  );


  nab2
  g0982
  (
    .dina(new_n1045__spl_),
    .dinb(new_n1046_),
    .dout(new_n1047_)
  );


  anb1
  g0983
  (
    .dina(new_n977__spl_),
    .dinb(new_n1047__spl_),
    .dout(new_n1048_)
  );


  anb2
  g0984
  (
    .dina(new_n977__spl_),
    .dinb(new_n1047__spl_),
    .dout(new_n1049_)
  );


  nab1
  g0985
  (
    .dina(new_n1048__spl_),
    .dinb(new_n1049_),
    .dout(new_n1050_)
  );


  anb2
  g0986
  (
    .dina(new_n976__spl_),
    .dinb(new_n1050__spl_),
    .dout(new_n1051_)
  );


  anb1
  g0987
  (
    .dina(new_n976__spl_),
    .dinb(new_n1050__spl_),
    .dout(new_n1052_)
  );


  nab2
  g0988
  (
    .dina(new_n1051__spl_),
    .dinb(new_n1052_),
    .dout(new_n1053_)
  );


  anb1
  g0989
  (
    .dina(new_n975__spl_),
    .dinb(new_n1053__spl_),
    .dout(new_n1054_)
  );


  anb2
  g0990
  (
    .dina(new_n975__spl_),
    .dinb(new_n1053__spl_),
    .dout(new_n1055_)
  );


  nab1
  g0991
  (
    .dina(new_n1054__spl_),
    .dinb(new_n1055_),
    .dout(new_n1056_)
  );


  anb2
  g0992
  (
    .dina(new_n974__spl_),
    .dinb(new_n1056__spl_),
    .dout(new_n1057_)
  );


  anb1
  g0993
  (
    .dina(new_n974__spl_),
    .dinb(new_n1056__spl_),
    .dout(new_n1058_)
  );


  anb1
  g0994
  (
    .dina(new_n1057__spl_),
    .dinb(new_n1058_),
    .dout(new_n1059_)
  );


  anb2
  g0995
  (
    .dina(new_n973__spl_),
    .dinb(new_n1059__spl_),
    .dout(new_n1060_)
  );


  anb1
  g0996
  (
    .dina(new_n973__spl_),
    .dinb(new_n1059__spl_),
    .dout(new_n1061_)
  );


  anb1
  g0997
  (
    .dina(new_n1060__spl_),
    .dinb(new_n1061_),
    .dout(new_n1062_)
  );


  anb2
  g0998
  (
    .dina(new_n972__spl_),
    .dinb(new_n1062__spl_),
    .dout(new_n1063_)
  );


  anb1
  g0999
  (
    .dina(new_n972__spl_),
    .dinb(new_n1062__spl_),
    .dout(new_n1064_)
  );


  anb1
  g1000
  (
    .dina(new_n1063__spl_),
    .dinb(new_n1064_),
    .dout(new_n1065_)
  );


  anb2
  g1001
  (
    .dina(new_n971__spl_),
    .dinb(new_n1065__spl_),
    .dout(new_n1066_)
  );


  anb1
  g1002
  (
    .dina(new_n971__spl_),
    .dinb(new_n1065__spl_),
    .dout(new_n1067_)
  );


  anb1
  g1003
  (
    .dina(new_n1066__spl_),
    .dinb(new_n1067_),
    .dout(new_n1068_)
  );


  anb2
  g1004
  (
    .dina(new_n970__spl_),
    .dinb(new_n1068__spl_),
    .dout(new_n1069_)
  );


  anb1
  g1005
  (
    .dina(new_n970__spl_),
    .dinb(new_n1068__spl_),
    .dout(new_n1070_)
  );


  anb1
  g1006
  (
    .dina(new_n1069__spl_),
    .dinb(new_n1070_),
    .dout(new_n1071_)
  );


  anb2
  g1007
  (
    .dina(new_n969__spl_),
    .dinb(new_n1071__spl_),
    .dout(new_n1072_)
  );


  anb1
  g1008
  (
    .dina(new_n969__spl_),
    .dinb(new_n1071__spl_),
    .dout(new_n1073_)
  );


  anb1
  g1009
  (
    .dina(new_n1072__spl_),
    .dinb(new_n1073_),
    .dout(new_n1074_)
  );


  anb2
  g1010
  (
    .dina(new_n968__spl_),
    .dinb(new_n1074__spl_),
    .dout(new_n1075_)
  );


  anb1
  g1011
  (
    .dina(new_n968__spl_),
    .dinb(new_n1074__spl_),
    .dout(new_n1076_)
  );


  anb1
  g1012
  (
    .dina(new_n1075__spl_),
    .dinb(new_n1076_),
    .dout(new_n1077_)
  );


  anb2
  g1013
  (
    .dina(new_n967__spl_),
    .dinb(new_n1077__spl_),
    .dout(new_n1078_)
  );


  anb2
  g1014
  (
    .dina(new_n1077__spl_),
    .dinb(new_n967__spl_),
    .dout(new_n1079_)
  );


  and1
  g1015
  (
    .dina(new_n1078_),
    .dinb(new_n1079__spl_0),
    .dout(G6273)
  );


  nor2
  g1016
  (
    .dina(new_n1072__spl_),
    .dinb(new_n1075__spl_),
    .dout(new_n1081_)
  );


  nor2
  g1017
  (
    .dina(G3_spl_111),
    .dinb(G32_spl_001),
    .dout(new_n1082_)
  );


  nor2
  g1018
  (
    .dina(new_n1066__spl_),
    .dinb(new_n1069__spl_),
    .dout(new_n1083_)
  );


  nor2
  g1019
  (
    .dina(G4_spl_111),
    .dinb(G31_spl_001),
    .dout(new_n1084_)
  );


  nor2
  g1020
  (
    .dina(new_n1060__spl_),
    .dinb(new_n1063__spl_),
    .dout(new_n1085_)
  );


  nor2
  g1021
  (
    .dina(G5_spl_110),
    .dinb(G30_spl_010),
    .dout(new_n1086_)
  );


  anb2
  g1022
  (
    .dina(new_n1054__spl_),
    .dinb(new_n1057__spl_),
    .dout(new_n1087_)
  );


  and1
  g1023
  (
    .dina(G6_spl_110),
    .dinb(G29_spl_010),
    .dout(new_n1088_)
  );


  anb2
  g1024
  (
    .dina(new_n1048__spl_),
    .dinb(new_n1051__spl_),
    .dout(new_n1089_)
  );


  and1
  g1025
  (
    .dina(G7_spl_101),
    .dinb(G28_spl_011),
    .dout(new_n1090_)
  );


  anb2
  g1026
  (
    .dina(new_n1042__spl_),
    .dinb(new_n1045__spl_),
    .dout(new_n1091_)
  );


  and1
  g1027
  (
    .dina(G8_spl_101),
    .dinb(G27_spl_011),
    .dout(new_n1092_)
  );


  anb2
  g1028
  (
    .dina(new_n1036__spl_),
    .dinb(new_n1039__spl_),
    .dout(new_n1093_)
  );


  and1
  g1029
  (
    .dina(G9_spl_100),
    .dinb(G26_spl_100),
    .dout(new_n1094_)
  );


  anb2
  g1030
  (
    .dina(new_n1030__spl_),
    .dinb(new_n1033__spl_),
    .dout(new_n1095_)
  );


  and1
  g1031
  (
    .dina(G10_spl_100),
    .dinb(G25_spl_100),
    .dout(new_n1096_)
  );


  anb2
  g1032
  (
    .dina(new_n1024__spl_),
    .dinb(new_n1027__spl_),
    .dout(new_n1097_)
  );


  and1
  g1033
  (
    .dina(G11_spl_011),
    .dinb(G24_spl_101),
    .dout(new_n1098_)
  );


  anb2
  g1034
  (
    .dina(new_n1018__spl_),
    .dinb(new_n1021__spl_),
    .dout(new_n1099_)
  );


  and1
  g1035
  (
    .dina(G12_spl_011),
    .dinb(G23_spl_101),
    .dout(new_n1100_)
  );


  anb2
  g1036
  (
    .dina(new_n1012__spl_),
    .dinb(new_n1015__spl_),
    .dout(new_n1101_)
  );


  and1
  g1037
  (
    .dina(G13_spl_010),
    .dinb(G22_spl_110),
    .dout(new_n1102_)
  );


  anb2
  g1038
  (
    .dina(new_n1006__spl_),
    .dinb(new_n1009__spl_),
    .dout(new_n1103_)
  );


  and1
  g1039
  (
    .dina(G14_spl_010),
    .dinb(G21_spl_110),
    .dout(new_n1104_)
  );


  anb2
  g1040
  (
    .dina(new_n1000__spl_),
    .dinb(new_n1003__spl_),
    .dout(new_n1105_)
  );


  and1
  g1041
  (
    .dina(G15_spl_001),
    .dinb(G20_spl_111),
    .dout(new_n1106_)
  );


  nor2
  g1042
  (
    .dina(G16_spl_001),
    .dinb(G19_spl_111),
    .dout(new_n1107_)
  );


  anb1
  g1043
  (
    .dina(new_n994__spl_),
    .dinb(new_n997__spl_),
    .dout(new_n1108_)
  );


  anb1
  g1044
  (
    .dina(new_n1107__spl_),
    .dinb(new_n1108__spl_),
    .dout(new_n1109_)
  );


  anb2
  g1045
  (
    .dina(new_n1107__spl_),
    .dinb(new_n1108__spl_),
    .dout(new_n1110_)
  );


  nab1
  g1046
  (
    .dina(new_n1109__spl_),
    .dinb(new_n1110_),
    .dout(new_n1111_)
  );


  anb2
  g1047
  (
    .dina(new_n1106__spl_),
    .dinb(new_n1111__spl_),
    .dout(new_n1112_)
  );


  anb1
  g1048
  (
    .dina(new_n1106__spl_),
    .dinb(new_n1111__spl_),
    .dout(new_n1113_)
  );


  nab2
  g1049
  (
    .dina(new_n1112__spl_),
    .dinb(new_n1113_),
    .dout(new_n1114_)
  );


  anb1
  g1050
  (
    .dina(new_n1105__spl_),
    .dinb(new_n1114__spl_),
    .dout(new_n1115_)
  );


  anb2
  g1051
  (
    .dina(new_n1105__spl_),
    .dinb(new_n1114__spl_),
    .dout(new_n1116_)
  );


  nab1
  g1052
  (
    .dina(new_n1115__spl_),
    .dinb(new_n1116_),
    .dout(new_n1117_)
  );


  anb2
  g1053
  (
    .dina(new_n1104__spl_),
    .dinb(new_n1117__spl_),
    .dout(new_n1118_)
  );


  anb1
  g1054
  (
    .dina(new_n1104__spl_),
    .dinb(new_n1117__spl_),
    .dout(new_n1119_)
  );


  nab2
  g1055
  (
    .dina(new_n1118__spl_),
    .dinb(new_n1119_),
    .dout(new_n1120_)
  );


  anb1
  g1056
  (
    .dina(new_n1103__spl_),
    .dinb(new_n1120__spl_),
    .dout(new_n1121_)
  );


  anb2
  g1057
  (
    .dina(new_n1103__spl_),
    .dinb(new_n1120__spl_),
    .dout(new_n1122_)
  );


  nab1
  g1058
  (
    .dina(new_n1121__spl_),
    .dinb(new_n1122_),
    .dout(new_n1123_)
  );


  anb2
  g1059
  (
    .dina(new_n1102__spl_),
    .dinb(new_n1123__spl_),
    .dout(new_n1124_)
  );


  anb1
  g1060
  (
    .dina(new_n1102__spl_),
    .dinb(new_n1123__spl_),
    .dout(new_n1125_)
  );


  nab2
  g1061
  (
    .dina(new_n1124__spl_),
    .dinb(new_n1125_),
    .dout(new_n1126_)
  );


  anb1
  g1062
  (
    .dina(new_n1101__spl_),
    .dinb(new_n1126__spl_),
    .dout(new_n1127_)
  );


  anb2
  g1063
  (
    .dina(new_n1101__spl_),
    .dinb(new_n1126__spl_),
    .dout(new_n1128_)
  );


  nab1
  g1064
  (
    .dina(new_n1127__spl_),
    .dinb(new_n1128_),
    .dout(new_n1129_)
  );


  anb2
  g1065
  (
    .dina(new_n1100__spl_),
    .dinb(new_n1129__spl_),
    .dout(new_n1130_)
  );


  anb1
  g1066
  (
    .dina(new_n1100__spl_),
    .dinb(new_n1129__spl_),
    .dout(new_n1131_)
  );


  nab2
  g1067
  (
    .dina(new_n1130__spl_),
    .dinb(new_n1131_),
    .dout(new_n1132_)
  );


  anb1
  g1068
  (
    .dina(new_n1099__spl_),
    .dinb(new_n1132__spl_),
    .dout(new_n1133_)
  );


  anb2
  g1069
  (
    .dina(new_n1099__spl_),
    .dinb(new_n1132__spl_),
    .dout(new_n1134_)
  );


  nab1
  g1070
  (
    .dina(new_n1133__spl_),
    .dinb(new_n1134_),
    .dout(new_n1135_)
  );


  anb2
  g1071
  (
    .dina(new_n1098__spl_),
    .dinb(new_n1135__spl_),
    .dout(new_n1136_)
  );


  anb1
  g1072
  (
    .dina(new_n1098__spl_),
    .dinb(new_n1135__spl_),
    .dout(new_n1137_)
  );


  nab2
  g1073
  (
    .dina(new_n1136__spl_),
    .dinb(new_n1137_),
    .dout(new_n1138_)
  );


  anb1
  g1074
  (
    .dina(new_n1097__spl_),
    .dinb(new_n1138__spl_),
    .dout(new_n1139_)
  );


  anb2
  g1075
  (
    .dina(new_n1097__spl_),
    .dinb(new_n1138__spl_),
    .dout(new_n1140_)
  );


  nab1
  g1076
  (
    .dina(new_n1139__spl_),
    .dinb(new_n1140_),
    .dout(new_n1141_)
  );


  anb2
  g1077
  (
    .dina(new_n1096__spl_),
    .dinb(new_n1141__spl_),
    .dout(new_n1142_)
  );


  anb1
  g1078
  (
    .dina(new_n1096__spl_),
    .dinb(new_n1141__spl_),
    .dout(new_n1143_)
  );


  nab2
  g1079
  (
    .dina(new_n1142__spl_),
    .dinb(new_n1143_),
    .dout(new_n1144_)
  );


  anb1
  g1080
  (
    .dina(new_n1095__spl_),
    .dinb(new_n1144__spl_),
    .dout(new_n1145_)
  );


  anb2
  g1081
  (
    .dina(new_n1095__spl_),
    .dinb(new_n1144__spl_),
    .dout(new_n1146_)
  );


  nab1
  g1082
  (
    .dina(new_n1145__spl_),
    .dinb(new_n1146_),
    .dout(new_n1147_)
  );


  anb2
  g1083
  (
    .dina(new_n1094__spl_),
    .dinb(new_n1147__spl_),
    .dout(new_n1148_)
  );


  anb1
  g1084
  (
    .dina(new_n1094__spl_),
    .dinb(new_n1147__spl_),
    .dout(new_n1149_)
  );


  nab2
  g1085
  (
    .dina(new_n1148__spl_),
    .dinb(new_n1149_),
    .dout(new_n1150_)
  );


  anb1
  g1086
  (
    .dina(new_n1093__spl_),
    .dinb(new_n1150__spl_),
    .dout(new_n1151_)
  );


  anb2
  g1087
  (
    .dina(new_n1093__spl_),
    .dinb(new_n1150__spl_),
    .dout(new_n1152_)
  );


  nab1
  g1088
  (
    .dina(new_n1151__spl_),
    .dinb(new_n1152_),
    .dout(new_n1153_)
  );


  anb2
  g1089
  (
    .dina(new_n1092__spl_),
    .dinb(new_n1153__spl_),
    .dout(new_n1154_)
  );


  anb1
  g1090
  (
    .dina(new_n1092__spl_),
    .dinb(new_n1153__spl_),
    .dout(new_n1155_)
  );


  nab2
  g1091
  (
    .dina(new_n1154__spl_),
    .dinb(new_n1155_),
    .dout(new_n1156_)
  );


  anb1
  g1092
  (
    .dina(new_n1091__spl_),
    .dinb(new_n1156__spl_),
    .dout(new_n1157_)
  );


  anb2
  g1093
  (
    .dina(new_n1091__spl_),
    .dinb(new_n1156__spl_),
    .dout(new_n1158_)
  );


  nab1
  g1094
  (
    .dina(new_n1157__spl_),
    .dinb(new_n1158_),
    .dout(new_n1159_)
  );


  anb2
  g1095
  (
    .dina(new_n1090__spl_),
    .dinb(new_n1159__spl_),
    .dout(new_n1160_)
  );


  anb1
  g1096
  (
    .dina(new_n1090__spl_),
    .dinb(new_n1159__spl_),
    .dout(new_n1161_)
  );


  nab2
  g1097
  (
    .dina(new_n1160__spl_),
    .dinb(new_n1161_),
    .dout(new_n1162_)
  );


  anb1
  g1098
  (
    .dina(new_n1089__spl_),
    .dinb(new_n1162__spl_),
    .dout(new_n1163_)
  );


  anb2
  g1099
  (
    .dina(new_n1089__spl_),
    .dinb(new_n1162__spl_),
    .dout(new_n1164_)
  );


  nab1
  g1100
  (
    .dina(new_n1163__spl_),
    .dinb(new_n1164_),
    .dout(new_n1165_)
  );


  anb2
  g1101
  (
    .dina(new_n1088__spl_),
    .dinb(new_n1165__spl_),
    .dout(new_n1166_)
  );


  anb1
  g1102
  (
    .dina(new_n1088__spl_),
    .dinb(new_n1165__spl_),
    .dout(new_n1167_)
  );


  nab2
  g1103
  (
    .dina(new_n1166__spl_),
    .dinb(new_n1167_),
    .dout(new_n1168_)
  );


  anb1
  g1104
  (
    .dina(new_n1087__spl_),
    .dinb(new_n1168__spl_),
    .dout(new_n1169_)
  );


  anb2
  g1105
  (
    .dina(new_n1087__spl_),
    .dinb(new_n1168__spl_),
    .dout(new_n1170_)
  );


  anb2
  g1106
  (
    .dina(new_n1169__spl_),
    .dinb(new_n1170_),
    .dout(new_n1171_)
  );


  anb1
  g1107
  (
    .dina(new_n1086__spl_),
    .dinb(new_n1171__spl_),
    .dout(new_n1172_)
  );


  anb2
  g1108
  (
    .dina(new_n1086__spl_),
    .dinb(new_n1171__spl_),
    .dout(new_n1173_)
  );


  anb2
  g1109
  (
    .dina(new_n1172__spl_),
    .dinb(new_n1173_),
    .dout(new_n1174_)
  );


  anb1
  g1110
  (
    .dina(new_n1085__spl_),
    .dinb(new_n1174__spl_),
    .dout(new_n1175_)
  );


  anb2
  g1111
  (
    .dina(new_n1085__spl_),
    .dinb(new_n1174__spl_),
    .dout(new_n1176_)
  );


  anb2
  g1112
  (
    .dina(new_n1175__spl_),
    .dinb(new_n1176_),
    .dout(new_n1177_)
  );


  anb1
  g1113
  (
    .dina(new_n1084__spl_),
    .dinb(new_n1177__spl_),
    .dout(new_n1178_)
  );


  anb2
  g1114
  (
    .dina(new_n1084__spl_),
    .dinb(new_n1177__spl_),
    .dout(new_n1179_)
  );


  anb2
  g1115
  (
    .dina(new_n1178__spl_),
    .dinb(new_n1179_),
    .dout(new_n1180_)
  );


  anb1
  g1116
  (
    .dina(new_n1083__spl_),
    .dinb(new_n1180__spl_),
    .dout(new_n1181_)
  );


  anb2
  g1117
  (
    .dina(new_n1083__spl_),
    .dinb(new_n1180__spl_),
    .dout(new_n1182_)
  );


  anb2
  g1118
  (
    .dina(new_n1181__spl_),
    .dinb(new_n1182_),
    .dout(new_n1183_)
  );


  anb1
  g1119
  (
    .dina(new_n1082__spl_),
    .dinb(new_n1183__spl_),
    .dout(new_n1184_)
  );


  anb2
  g1120
  (
    .dina(new_n1082__spl_),
    .dinb(new_n1183__spl_),
    .dout(new_n1185_)
  );


  anb2
  g1121
  (
    .dina(new_n1184__spl_),
    .dinb(new_n1185_),
    .dout(new_n1186_)
  );


  anb1
  g1122
  (
    .dina(new_n1081__spl_),
    .dinb(new_n1186__spl_),
    .dout(new_n1187_)
  );


  anb2
  g1123
  (
    .dina(new_n1081__spl_),
    .dinb(new_n1186__spl_),
    .dout(new_n1188_)
  );


  anb2
  g1124
  (
    .dina(new_n1187__spl_),
    .dinb(new_n1188_),
    .dout(new_n1189_)
  );


  anb1
  g1125
  (
    .dina(new_n1079__spl_0),
    .dinb(new_n1189__spl_),
    .dout(new_n1190_)
  );


  anb2
  g1126
  (
    .dina(new_n1079__spl_),
    .dinb(new_n1189__spl_),
    .dout(new_n1191_)
  );


  anb2
  g1127
  (
    .dina(new_n1190__spl_),
    .dinb(new_n1191_),
    .dout(G6274)
  );


  and2
  g1128
  (
    .dina(new_n1187__spl_),
    .dinb(new_n1190__spl_),
    .dout(new_n1193_)
  );


  and2
  g1129
  (
    .dina(new_n1181__spl_),
    .dinb(new_n1184__spl_),
    .dout(new_n1194_)
  );


  nor2
  g1130
  (
    .dina(G4_spl_111),
    .dinb(G32_spl_001),
    .dout(new_n1195_)
  );


  and2
  g1131
  (
    .dina(new_n1175__spl_),
    .dinb(new_n1178__spl_),
    .dout(new_n1196_)
  );


  nor2
  g1132
  (
    .dina(G5_spl_111),
    .dinb(G31_spl_010),
    .dout(new_n1197_)
  );


  and2
  g1133
  (
    .dina(new_n1169__spl_),
    .dinb(new_n1172__spl_),
    .dout(new_n1198_)
  );


  nor2
  g1134
  (
    .dina(G6_spl_110),
    .dinb(G30_spl_010),
    .dout(new_n1199_)
  );


  anb2
  g1135
  (
    .dina(new_n1163__spl_),
    .dinb(new_n1166__spl_),
    .dout(new_n1200_)
  );


  and1
  g1136
  (
    .dina(G7_spl_110),
    .dinb(G29_spl_011),
    .dout(new_n1201_)
  );


  anb2
  g1137
  (
    .dina(new_n1157__spl_),
    .dinb(new_n1160__spl_),
    .dout(new_n1202_)
  );


  and1
  g1138
  (
    .dina(G8_spl_101),
    .dinb(G28_spl_011),
    .dout(new_n1203_)
  );


  anb2
  g1139
  (
    .dina(new_n1151__spl_),
    .dinb(new_n1154__spl_),
    .dout(new_n1204_)
  );


  and1
  g1140
  (
    .dina(G9_spl_101),
    .dinb(G27_spl_100),
    .dout(new_n1205_)
  );


  anb2
  g1141
  (
    .dina(new_n1145__spl_),
    .dinb(new_n1148__spl_),
    .dout(new_n1206_)
  );


  and1
  g1142
  (
    .dina(G10_spl_100),
    .dinb(G26_spl_100),
    .dout(new_n1207_)
  );


  anb2
  g1143
  (
    .dina(new_n1139__spl_),
    .dinb(new_n1142__spl_),
    .dout(new_n1208_)
  );


  and1
  g1144
  (
    .dina(G11_spl_100),
    .dinb(G25_spl_101),
    .dout(new_n1209_)
  );


  anb2
  g1145
  (
    .dina(new_n1133__spl_),
    .dinb(new_n1136__spl_),
    .dout(new_n1210_)
  );


  and1
  g1146
  (
    .dina(G12_spl_011),
    .dinb(G24_spl_101),
    .dout(new_n1211_)
  );


  anb2
  g1147
  (
    .dina(new_n1127__spl_),
    .dinb(new_n1130__spl_),
    .dout(new_n1212_)
  );


  and1
  g1148
  (
    .dina(G13_spl_011),
    .dinb(G23_spl_110),
    .dout(new_n1213_)
  );


  anb2
  g1149
  (
    .dina(new_n1121__spl_),
    .dinb(new_n1124__spl_),
    .dout(new_n1214_)
  );


  and1
  g1150
  (
    .dina(G14_spl_010),
    .dinb(G22_spl_110),
    .dout(new_n1215_)
  );


  anb2
  g1151
  (
    .dina(new_n1115__spl_),
    .dinb(new_n1118__spl_),
    .dout(new_n1216_)
  );


  nor2
  g1152
  (
    .dina(G15_spl_010),
    .dinb(G21_spl_111),
    .dout(new_n1217_)
  );


  and1
  g1153
  (
    .dina(G16_spl_001),
    .dinb(G20_spl_111),
    .dout(new_n1218_)
  );


  anb2
  g1154
  (
    .dina(new_n1109__spl_),
    .dinb(new_n1112__spl_),
    .dout(new_n1219_)
  );


  anb2
  g1155
  (
    .dina(new_n1218__spl_),
    .dinb(new_n1219__spl_),
    .dout(new_n1220_)
  );


  anb1
  g1156
  (
    .dina(new_n1218__spl_),
    .dinb(new_n1219__spl_),
    .dout(new_n1221_)
  );


  nab2
  g1157
  (
    .dina(new_n1220__spl_),
    .dinb(new_n1221_),
    .dout(new_n1222_)
  );


  anb1
  g1158
  (
    .dina(new_n1217__spl_),
    .dinb(new_n1222__spl_),
    .dout(new_n1223_)
  );


  anb2
  g1159
  (
    .dina(new_n1217__spl_),
    .dinb(new_n1222__spl_),
    .dout(new_n1224_)
  );


  anb2
  g1160
  (
    .dina(new_n1223__spl_),
    .dinb(new_n1224_),
    .dout(new_n1225_)
  );


  anb1
  g1161
  (
    .dina(new_n1216__spl_),
    .dinb(new_n1225__spl_),
    .dout(new_n1226_)
  );


  anb2
  g1162
  (
    .dina(new_n1216__spl_),
    .dinb(new_n1225__spl_),
    .dout(new_n1227_)
  );


  nab1
  g1163
  (
    .dina(new_n1226__spl_),
    .dinb(new_n1227_),
    .dout(new_n1228_)
  );


  anb2
  g1164
  (
    .dina(new_n1215__spl_),
    .dinb(new_n1228__spl_),
    .dout(new_n1229_)
  );


  anb1
  g1165
  (
    .dina(new_n1215__spl_),
    .dinb(new_n1228__spl_),
    .dout(new_n1230_)
  );


  nab2
  g1166
  (
    .dina(new_n1229__spl_),
    .dinb(new_n1230_),
    .dout(new_n1231_)
  );


  anb1
  g1167
  (
    .dina(new_n1214__spl_),
    .dinb(new_n1231__spl_),
    .dout(new_n1232_)
  );


  anb2
  g1168
  (
    .dina(new_n1214__spl_),
    .dinb(new_n1231__spl_),
    .dout(new_n1233_)
  );


  nab1
  g1169
  (
    .dina(new_n1232__spl_),
    .dinb(new_n1233_),
    .dout(new_n1234_)
  );


  anb2
  g1170
  (
    .dina(new_n1213__spl_),
    .dinb(new_n1234__spl_),
    .dout(new_n1235_)
  );


  anb1
  g1171
  (
    .dina(new_n1213__spl_),
    .dinb(new_n1234__spl_),
    .dout(new_n1236_)
  );


  nab2
  g1172
  (
    .dina(new_n1235__spl_),
    .dinb(new_n1236_),
    .dout(new_n1237_)
  );


  anb1
  g1173
  (
    .dina(new_n1212__spl_),
    .dinb(new_n1237__spl_),
    .dout(new_n1238_)
  );


  anb2
  g1174
  (
    .dina(new_n1212__spl_),
    .dinb(new_n1237__spl_),
    .dout(new_n1239_)
  );


  nab1
  g1175
  (
    .dina(new_n1238__spl_),
    .dinb(new_n1239_),
    .dout(new_n1240_)
  );


  anb2
  g1176
  (
    .dina(new_n1211__spl_),
    .dinb(new_n1240__spl_),
    .dout(new_n1241_)
  );


  anb1
  g1177
  (
    .dina(new_n1211__spl_),
    .dinb(new_n1240__spl_),
    .dout(new_n1242_)
  );


  nab2
  g1178
  (
    .dina(new_n1241__spl_),
    .dinb(new_n1242_),
    .dout(new_n1243_)
  );


  anb1
  g1179
  (
    .dina(new_n1210__spl_),
    .dinb(new_n1243__spl_),
    .dout(new_n1244_)
  );


  anb2
  g1180
  (
    .dina(new_n1210__spl_),
    .dinb(new_n1243__spl_),
    .dout(new_n1245_)
  );


  nab1
  g1181
  (
    .dina(new_n1244__spl_),
    .dinb(new_n1245_),
    .dout(new_n1246_)
  );


  anb2
  g1182
  (
    .dina(new_n1209__spl_),
    .dinb(new_n1246__spl_),
    .dout(new_n1247_)
  );


  anb1
  g1183
  (
    .dina(new_n1209__spl_),
    .dinb(new_n1246__spl_),
    .dout(new_n1248_)
  );


  nab2
  g1184
  (
    .dina(new_n1247__spl_),
    .dinb(new_n1248_),
    .dout(new_n1249_)
  );


  anb1
  g1185
  (
    .dina(new_n1208__spl_),
    .dinb(new_n1249__spl_),
    .dout(new_n1250_)
  );


  anb2
  g1186
  (
    .dina(new_n1208__spl_),
    .dinb(new_n1249__spl_),
    .dout(new_n1251_)
  );


  nab1
  g1187
  (
    .dina(new_n1250__spl_),
    .dinb(new_n1251_),
    .dout(new_n1252_)
  );


  anb2
  g1188
  (
    .dina(new_n1207__spl_),
    .dinb(new_n1252__spl_),
    .dout(new_n1253_)
  );


  anb1
  g1189
  (
    .dina(new_n1207__spl_),
    .dinb(new_n1252__spl_),
    .dout(new_n1254_)
  );


  nab2
  g1190
  (
    .dina(new_n1253__spl_),
    .dinb(new_n1254_),
    .dout(new_n1255_)
  );


  anb1
  g1191
  (
    .dina(new_n1206__spl_),
    .dinb(new_n1255__spl_),
    .dout(new_n1256_)
  );


  anb2
  g1192
  (
    .dina(new_n1206__spl_),
    .dinb(new_n1255__spl_),
    .dout(new_n1257_)
  );


  nab1
  g1193
  (
    .dina(new_n1256__spl_),
    .dinb(new_n1257_),
    .dout(new_n1258_)
  );


  anb2
  g1194
  (
    .dina(new_n1205__spl_),
    .dinb(new_n1258__spl_),
    .dout(new_n1259_)
  );


  anb1
  g1195
  (
    .dina(new_n1205__spl_),
    .dinb(new_n1258__spl_),
    .dout(new_n1260_)
  );


  nab2
  g1196
  (
    .dina(new_n1259__spl_),
    .dinb(new_n1260_),
    .dout(new_n1261_)
  );


  anb1
  g1197
  (
    .dina(new_n1204__spl_),
    .dinb(new_n1261__spl_),
    .dout(new_n1262_)
  );


  anb2
  g1198
  (
    .dina(new_n1204__spl_),
    .dinb(new_n1261__spl_),
    .dout(new_n1263_)
  );


  nab1
  g1199
  (
    .dina(new_n1262__spl_),
    .dinb(new_n1263_),
    .dout(new_n1264_)
  );


  anb2
  g1200
  (
    .dina(new_n1203__spl_),
    .dinb(new_n1264__spl_),
    .dout(new_n1265_)
  );


  anb1
  g1201
  (
    .dina(new_n1203__spl_),
    .dinb(new_n1264__spl_),
    .dout(new_n1266_)
  );


  nab2
  g1202
  (
    .dina(new_n1265__spl_),
    .dinb(new_n1266_),
    .dout(new_n1267_)
  );


  anb1
  g1203
  (
    .dina(new_n1202__spl_),
    .dinb(new_n1267__spl_),
    .dout(new_n1268_)
  );


  anb2
  g1204
  (
    .dina(new_n1202__spl_),
    .dinb(new_n1267__spl_),
    .dout(new_n1269_)
  );


  nab1
  g1205
  (
    .dina(new_n1268__spl_),
    .dinb(new_n1269_),
    .dout(new_n1270_)
  );


  anb2
  g1206
  (
    .dina(new_n1201__spl_),
    .dinb(new_n1270__spl_),
    .dout(new_n1271_)
  );


  anb1
  g1207
  (
    .dina(new_n1201__spl_),
    .dinb(new_n1270__spl_),
    .dout(new_n1272_)
  );


  nab2
  g1208
  (
    .dina(new_n1271__spl_),
    .dinb(new_n1272_),
    .dout(new_n1273_)
  );


  anb1
  g1209
  (
    .dina(new_n1200__spl_),
    .dinb(new_n1273__spl_),
    .dout(new_n1274_)
  );


  anb2
  g1210
  (
    .dina(new_n1200__spl_),
    .dinb(new_n1273__spl_),
    .dout(new_n1275_)
  );


  anb2
  g1211
  (
    .dina(new_n1274__spl_),
    .dinb(new_n1275_),
    .dout(new_n1276_)
  );


  anb1
  g1212
  (
    .dina(new_n1199__spl_),
    .dinb(new_n1276__spl_),
    .dout(new_n1277_)
  );


  anb2
  g1213
  (
    .dina(new_n1199__spl_),
    .dinb(new_n1276__spl_),
    .dout(new_n1278_)
  );


  anb2
  g1214
  (
    .dina(new_n1277__spl_),
    .dinb(new_n1278_),
    .dout(new_n1279_)
  );


  anb1
  g1215
  (
    .dina(new_n1198__spl_),
    .dinb(new_n1279__spl_),
    .dout(new_n1280_)
  );


  anb2
  g1216
  (
    .dina(new_n1198__spl_),
    .dinb(new_n1279__spl_),
    .dout(new_n1281_)
  );


  anb2
  g1217
  (
    .dina(new_n1280__spl_),
    .dinb(new_n1281_),
    .dout(new_n1282_)
  );


  anb1
  g1218
  (
    .dina(new_n1197__spl_),
    .dinb(new_n1282__spl_),
    .dout(new_n1283_)
  );


  anb2
  g1219
  (
    .dina(new_n1197__spl_),
    .dinb(new_n1282__spl_),
    .dout(new_n1284_)
  );


  anb2
  g1220
  (
    .dina(new_n1283__spl_),
    .dinb(new_n1284_),
    .dout(new_n1285_)
  );


  anb1
  g1221
  (
    .dina(new_n1196__spl_),
    .dinb(new_n1285__spl_),
    .dout(new_n1286_)
  );


  anb2
  g1222
  (
    .dina(new_n1196__spl_),
    .dinb(new_n1285__spl_),
    .dout(new_n1287_)
  );


  anb2
  g1223
  (
    .dina(new_n1286__spl_),
    .dinb(new_n1287_),
    .dout(new_n1288_)
  );


  anb1
  g1224
  (
    .dina(new_n1195__spl_),
    .dinb(new_n1288__spl_),
    .dout(new_n1289_)
  );


  anb2
  g1225
  (
    .dina(new_n1195__spl_),
    .dinb(new_n1288__spl_),
    .dout(new_n1290_)
  );


  anb2
  g1226
  (
    .dina(new_n1289__spl_),
    .dinb(new_n1290_),
    .dout(new_n1291_)
  );


  anb1
  g1227
  (
    .dina(new_n1194__spl_),
    .dinb(new_n1291__spl_),
    .dout(new_n1292_)
  );


  anb2
  g1228
  (
    .dina(new_n1194__spl_),
    .dinb(new_n1291__spl_),
    .dout(new_n1293_)
  );


  anb2
  g1229
  (
    .dina(new_n1292__spl_),
    .dinb(new_n1293_),
    .dout(new_n1294_)
  );


  anb1
  g1230
  (
    .dina(new_n1193__spl_),
    .dinb(new_n1294__spl_),
    .dout(new_n1295_)
  );


  anb2
  g1231
  (
    .dina(new_n1193__spl_),
    .dinb(new_n1294__spl_),
    .dout(new_n1296_)
  );


  anb2
  g1232
  (
    .dina(new_n1295__spl_),
    .dinb(new_n1296_),
    .dout(G6275)
  );


  and2
  g1233
  (
    .dina(new_n1292__spl_),
    .dinb(new_n1295__spl_),
    .dout(new_n1298_)
  );


  and2
  g1234
  (
    .dina(new_n1286__spl_),
    .dinb(new_n1289__spl_),
    .dout(new_n1299_)
  );


  nor2
  g1235
  (
    .dina(G5_spl_111),
    .dinb(G32_spl_010),
    .dout(new_n1300_)
  );


  and2
  g1236
  (
    .dina(new_n1280__spl_),
    .dinb(new_n1283__spl_),
    .dout(new_n1301_)
  );


  nor2
  g1237
  (
    .dina(G6_spl_111),
    .dinb(G31_spl_010),
    .dout(new_n1302_)
  );


  and2
  g1238
  (
    .dina(new_n1274__spl_),
    .dinb(new_n1277__spl_),
    .dout(new_n1303_)
  );


  nor2
  g1239
  (
    .dina(G7_spl_110),
    .dinb(G30_spl_011),
    .dout(new_n1304_)
  );


  anb2
  g1240
  (
    .dina(new_n1268__spl_),
    .dinb(new_n1271__spl_),
    .dout(new_n1305_)
  );


  and1
  g1241
  (
    .dina(G8_spl_110),
    .dinb(G29_spl_011),
    .dout(new_n1306_)
  );


  anb2
  g1242
  (
    .dina(new_n1262__spl_),
    .dinb(new_n1265__spl_),
    .dout(new_n1307_)
  );


  and1
  g1243
  (
    .dina(G9_spl_101),
    .dinb(G28_spl_100),
    .dout(new_n1308_)
  );


  anb2
  g1244
  (
    .dina(new_n1256__spl_),
    .dinb(new_n1259__spl_),
    .dout(new_n1309_)
  );


  and1
  g1245
  (
    .dina(G10_spl_101),
    .dinb(G27_spl_100),
    .dout(new_n1310_)
  );


  anb2
  g1246
  (
    .dina(new_n1250__spl_),
    .dinb(new_n1253__spl_),
    .dout(new_n1311_)
  );


  and1
  g1247
  (
    .dina(G11_spl_100),
    .dinb(G26_spl_101),
    .dout(new_n1312_)
  );


  anb2
  g1248
  (
    .dina(new_n1244__spl_),
    .dinb(new_n1247__spl_),
    .dout(new_n1313_)
  );


  and1
  g1249
  (
    .dina(G12_spl_100),
    .dinb(G25_spl_101),
    .dout(new_n1314_)
  );


  anb2
  g1250
  (
    .dina(new_n1238__spl_),
    .dinb(new_n1241__spl_),
    .dout(new_n1315_)
  );


  and1
  g1251
  (
    .dina(G13_spl_011),
    .dinb(G24_spl_110),
    .dout(new_n1316_)
  );


  anb2
  g1252
  (
    .dina(new_n1232__spl_),
    .dinb(new_n1235__spl_),
    .dout(new_n1317_)
  );


  and1
  g1253
  (
    .dina(G14_spl_011),
    .dinb(G23_spl_110),
    .dout(new_n1318_)
  );


  anb2
  g1254
  (
    .dina(new_n1226__spl_),
    .dinb(new_n1229__spl_),
    .dout(new_n1319_)
  );


  and1
  g1255
  (
    .dina(G15_spl_010),
    .dinb(G22_spl_111),
    .dout(new_n1320_)
  );


  nor2
  g1256
  (
    .dina(G16_spl_010),
    .dinb(G21_spl_111),
    .dout(new_n1321_)
  );


  anb1
  g1257
  (
    .dina(new_n1220__spl_),
    .dinb(new_n1223__spl_),
    .dout(new_n1322_)
  );


  anb1
  g1258
  (
    .dina(new_n1321__spl_),
    .dinb(new_n1322__spl_),
    .dout(new_n1323_)
  );


  anb2
  g1259
  (
    .dina(new_n1321__spl_),
    .dinb(new_n1322__spl_),
    .dout(new_n1324_)
  );


  nab1
  g1260
  (
    .dina(new_n1323__spl_),
    .dinb(new_n1324_),
    .dout(new_n1325_)
  );


  anb2
  g1261
  (
    .dina(new_n1320__spl_),
    .dinb(new_n1325__spl_),
    .dout(new_n1326_)
  );


  anb1
  g1262
  (
    .dina(new_n1320__spl_),
    .dinb(new_n1325__spl_),
    .dout(new_n1327_)
  );


  nab2
  g1263
  (
    .dina(new_n1326__spl_),
    .dinb(new_n1327_),
    .dout(new_n1328_)
  );


  anb1
  g1264
  (
    .dina(new_n1319__spl_),
    .dinb(new_n1328__spl_),
    .dout(new_n1329_)
  );


  anb2
  g1265
  (
    .dina(new_n1319__spl_),
    .dinb(new_n1328__spl_),
    .dout(new_n1330_)
  );


  nab1
  g1266
  (
    .dina(new_n1329__spl_),
    .dinb(new_n1330_),
    .dout(new_n1331_)
  );


  anb2
  g1267
  (
    .dina(new_n1318__spl_),
    .dinb(new_n1331__spl_),
    .dout(new_n1332_)
  );


  anb1
  g1268
  (
    .dina(new_n1318__spl_),
    .dinb(new_n1331__spl_),
    .dout(new_n1333_)
  );


  nab2
  g1269
  (
    .dina(new_n1332__spl_),
    .dinb(new_n1333_),
    .dout(new_n1334_)
  );


  anb1
  g1270
  (
    .dina(new_n1317__spl_),
    .dinb(new_n1334__spl_),
    .dout(new_n1335_)
  );


  anb2
  g1271
  (
    .dina(new_n1317__spl_),
    .dinb(new_n1334__spl_),
    .dout(new_n1336_)
  );


  nab1
  g1272
  (
    .dina(new_n1335__spl_),
    .dinb(new_n1336_),
    .dout(new_n1337_)
  );


  anb2
  g1273
  (
    .dina(new_n1316__spl_),
    .dinb(new_n1337__spl_),
    .dout(new_n1338_)
  );


  anb1
  g1274
  (
    .dina(new_n1316__spl_),
    .dinb(new_n1337__spl_),
    .dout(new_n1339_)
  );


  nab2
  g1275
  (
    .dina(new_n1338__spl_),
    .dinb(new_n1339_),
    .dout(new_n1340_)
  );


  anb1
  g1276
  (
    .dina(new_n1315__spl_),
    .dinb(new_n1340__spl_),
    .dout(new_n1341_)
  );


  anb2
  g1277
  (
    .dina(new_n1315__spl_),
    .dinb(new_n1340__spl_),
    .dout(new_n1342_)
  );


  nab1
  g1278
  (
    .dina(new_n1341__spl_),
    .dinb(new_n1342_),
    .dout(new_n1343_)
  );


  anb2
  g1279
  (
    .dina(new_n1314__spl_),
    .dinb(new_n1343__spl_),
    .dout(new_n1344_)
  );


  anb1
  g1280
  (
    .dina(new_n1314__spl_),
    .dinb(new_n1343__spl_),
    .dout(new_n1345_)
  );


  nab2
  g1281
  (
    .dina(new_n1344__spl_),
    .dinb(new_n1345_),
    .dout(new_n1346_)
  );


  anb1
  g1282
  (
    .dina(new_n1313__spl_),
    .dinb(new_n1346__spl_),
    .dout(new_n1347_)
  );


  anb2
  g1283
  (
    .dina(new_n1313__spl_),
    .dinb(new_n1346__spl_),
    .dout(new_n1348_)
  );


  nab1
  g1284
  (
    .dina(new_n1347__spl_),
    .dinb(new_n1348_),
    .dout(new_n1349_)
  );


  anb2
  g1285
  (
    .dina(new_n1312__spl_),
    .dinb(new_n1349__spl_),
    .dout(new_n1350_)
  );


  anb1
  g1286
  (
    .dina(new_n1312__spl_),
    .dinb(new_n1349__spl_),
    .dout(new_n1351_)
  );


  nab2
  g1287
  (
    .dina(new_n1350__spl_),
    .dinb(new_n1351_),
    .dout(new_n1352_)
  );


  anb1
  g1288
  (
    .dina(new_n1311__spl_),
    .dinb(new_n1352__spl_),
    .dout(new_n1353_)
  );


  anb2
  g1289
  (
    .dina(new_n1311__spl_),
    .dinb(new_n1352__spl_),
    .dout(new_n1354_)
  );


  nab1
  g1290
  (
    .dina(new_n1353__spl_),
    .dinb(new_n1354_),
    .dout(new_n1355_)
  );


  anb2
  g1291
  (
    .dina(new_n1310__spl_),
    .dinb(new_n1355__spl_),
    .dout(new_n1356_)
  );


  anb1
  g1292
  (
    .dina(new_n1310__spl_),
    .dinb(new_n1355__spl_),
    .dout(new_n1357_)
  );


  nab2
  g1293
  (
    .dina(new_n1356__spl_),
    .dinb(new_n1357_),
    .dout(new_n1358_)
  );


  anb1
  g1294
  (
    .dina(new_n1309__spl_),
    .dinb(new_n1358__spl_),
    .dout(new_n1359_)
  );


  anb2
  g1295
  (
    .dina(new_n1309__spl_),
    .dinb(new_n1358__spl_),
    .dout(new_n1360_)
  );


  nab1
  g1296
  (
    .dina(new_n1359__spl_),
    .dinb(new_n1360_),
    .dout(new_n1361_)
  );


  anb2
  g1297
  (
    .dina(new_n1308__spl_),
    .dinb(new_n1361__spl_),
    .dout(new_n1362_)
  );


  anb1
  g1298
  (
    .dina(new_n1308__spl_),
    .dinb(new_n1361__spl_),
    .dout(new_n1363_)
  );


  nab2
  g1299
  (
    .dina(new_n1362__spl_),
    .dinb(new_n1363_),
    .dout(new_n1364_)
  );


  anb1
  g1300
  (
    .dina(new_n1307__spl_),
    .dinb(new_n1364__spl_),
    .dout(new_n1365_)
  );


  anb2
  g1301
  (
    .dina(new_n1307__spl_),
    .dinb(new_n1364__spl_),
    .dout(new_n1366_)
  );


  nab1
  g1302
  (
    .dina(new_n1365__spl_),
    .dinb(new_n1366_),
    .dout(new_n1367_)
  );


  anb2
  g1303
  (
    .dina(new_n1306__spl_),
    .dinb(new_n1367__spl_),
    .dout(new_n1368_)
  );


  anb1
  g1304
  (
    .dina(new_n1306__spl_),
    .dinb(new_n1367__spl_),
    .dout(new_n1369_)
  );


  nab2
  g1305
  (
    .dina(new_n1368__spl_),
    .dinb(new_n1369_),
    .dout(new_n1370_)
  );


  anb1
  g1306
  (
    .dina(new_n1305__spl_),
    .dinb(new_n1370__spl_),
    .dout(new_n1371_)
  );


  anb2
  g1307
  (
    .dina(new_n1305__spl_),
    .dinb(new_n1370__spl_),
    .dout(new_n1372_)
  );


  anb2
  g1308
  (
    .dina(new_n1371__spl_),
    .dinb(new_n1372_),
    .dout(new_n1373_)
  );


  anb1
  g1309
  (
    .dina(new_n1304__spl_),
    .dinb(new_n1373__spl_),
    .dout(new_n1374_)
  );


  anb2
  g1310
  (
    .dina(new_n1304__spl_),
    .dinb(new_n1373__spl_),
    .dout(new_n1375_)
  );


  anb2
  g1311
  (
    .dina(new_n1374__spl_),
    .dinb(new_n1375_),
    .dout(new_n1376_)
  );


  anb1
  g1312
  (
    .dina(new_n1303__spl_),
    .dinb(new_n1376__spl_),
    .dout(new_n1377_)
  );


  anb2
  g1313
  (
    .dina(new_n1303__spl_),
    .dinb(new_n1376__spl_),
    .dout(new_n1378_)
  );


  anb2
  g1314
  (
    .dina(new_n1377__spl_),
    .dinb(new_n1378_),
    .dout(new_n1379_)
  );


  anb1
  g1315
  (
    .dina(new_n1302__spl_),
    .dinb(new_n1379__spl_),
    .dout(new_n1380_)
  );


  anb2
  g1316
  (
    .dina(new_n1302__spl_),
    .dinb(new_n1379__spl_),
    .dout(new_n1381_)
  );


  anb2
  g1317
  (
    .dina(new_n1380__spl_),
    .dinb(new_n1381_),
    .dout(new_n1382_)
  );


  anb1
  g1318
  (
    .dina(new_n1301__spl_),
    .dinb(new_n1382__spl_),
    .dout(new_n1383_)
  );


  anb2
  g1319
  (
    .dina(new_n1301__spl_),
    .dinb(new_n1382__spl_),
    .dout(new_n1384_)
  );


  anb2
  g1320
  (
    .dina(new_n1383__spl_),
    .dinb(new_n1384_),
    .dout(new_n1385_)
  );


  anb1
  g1321
  (
    .dina(new_n1300__spl_),
    .dinb(new_n1385__spl_),
    .dout(new_n1386_)
  );


  anb2
  g1322
  (
    .dina(new_n1300__spl_),
    .dinb(new_n1385__spl_),
    .dout(new_n1387_)
  );


  anb2
  g1323
  (
    .dina(new_n1386__spl_),
    .dinb(new_n1387_),
    .dout(new_n1388_)
  );


  anb1
  g1324
  (
    .dina(new_n1299__spl_),
    .dinb(new_n1388__spl_),
    .dout(new_n1389_)
  );


  anb2
  g1325
  (
    .dina(new_n1299__spl_),
    .dinb(new_n1388__spl_),
    .dout(new_n1390_)
  );


  anb2
  g1326
  (
    .dina(new_n1389__spl_),
    .dinb(new_n1390_),
    .dout(new_n1391_)
  );


  anb1
  g1327
  (
    .dina(new_n1298__spl_),
    .dinb(new_n1391__spl_),
    .dout(new_n1392_)
  );


  anb2
  g1328
  (
    .dina(new_n1298__spl_),
    .dinb(new_n1391__spl_),
    .dout(new_n1393_)
  );


  anb2
  g1329
  (
    .dina(new_n1392__spl_),
    .dinb(new_n1393_),
    .dout(G6276)
  );


  and2
  g1330
  (
    .dina(new_n1389__spl_),
    .dinb(new_n1392__spl_),
    .dout(new_n1395_)
  );


  and2
  g1331
  (
    .dina(new_n1383__spl_),
    .dinb(new_n1386__spl_),
    .dout(new_n1396_)
  );


  nor2
  g1332
  (
    .dina(G6_spl_111),
    .dinb(G32_spl_010),
    .dout(new_n1397_)
  );


  and2
  g1333
  (
    .dina(new_n1377__spl_),
    .dinb(new_n1380__spl_),
    .dout(new_n1398_)
  );


  nor2
  g1334
  (
    .dina(G7_spl_111),
    .dinb(G31_spl_011),
    .dout(new_n1399_)
  );


  and2
  g1335
  (
    .dina(new_n1371__spl_),
    .dinb(new_n1374__spl_),
    .dout(new_n1400_)
  );


  nor2
  g1336
  (
    .dina(G8_spl_110),
    .dinb(G30_spl_011),
    .dout(new_n1401_)
  );


  anb2
  g1337
  (
    .dina(new_n1365__spl_),
    .dinb(new_n1368__spl_),
    .dout(new_n1402_)
  );


  and1
  g1338
  (
    .dina(G9_spl_110),
    .dinb(G29_spl_100),
    .dout(new_n1403_)
  );


  anb2
  g1339
  (
    .dina(new_n1359__spl_),
    .dinb(new_n1362__spl_),
    .dout(new_n1404_)
  );


  and1
  g1340
  (
    .dina(G10_spl_101),
    .dinb(G28_spl_100),
    .dout(new_n1405_)
  );


  anb2
  g1341
  (
    .dina(new_n1353__spl_),
    .dinb(new_n1356__spl_),
    .dout(new_n1406_)
  );


  and1
  g1342
  (
    .dina(G11_spl_101),
    .dinb(G27_spl_101),
    .dout(new_n1407_)
  );


  anb2
  g1343
  (
    .dina(new_n1347__spl_),
    .dinb(new_n1350__spl_),
    .dout(new_n1408_)
  );


  and1
  g1344
  (
    .dina(G12_spl_100),
    .dinb(G26_spl_101),
    .dout(new_n1409_)
  );


  anb2
  g1345
  (
    .dina(new_n1341__spl_),
    .dinb(new_n1344__spl_),
    .dout(new_n1410_)
  );


  and1
  g1346
  (
    .dina(G13_spl_100),
    .dinb(G25_spl_110),
    .dout(new_n1411_)
  );


  anb2
  g1347
  (
    .dina(new_n1335__spl_),
    .dinb(new_n1338__spl_),
    .dout(new_n1412_)
  );


  and1
  g1348
  (
    .dina(G14_spl_011),
    .dinb(G24_spl_110),
    .dout(new_n1413_)
  );


  anb2
  g1349
  (
    .dina(new_n1329__spl_),
    .dinb(new_n1332__spl_),
    .dout(new_n1414_)
  );


  nor2
  g1350
  (
    .dina(G15_spl_011),
    .dinb(G23_spl_111),
    .dout(new_n1415_)
  );


  and1
  g1351
  (
    .dina(G16_spl_010),
    .dinb(G22_spl_111),
    .dout(new_n1416_)
  );


  anb2
  g1352
  (
    .dina(new_n1323__spl_),
    .dinb(new_n1326__spl_),
    .dout(new_n1417_)
  );


  anb2
  g1353
  (
    .dina(new_n1416__spl_),
    .dinb(new_n1417__spl_),
    .dout(new_n1418_)
  );


  anb1
  g1354
  (
    .dina(new_n1416__spl_),
    .dinb(new_n1417__spl_),
    .dout(new_n1419_)
  );


  nab2
  g1355
  (
    .dina(new_n1418__spl_),
    .dinb(new_n1419_),
    .dout(new_n1420_)
  );


  anb1
  g1356
  (
    .dina(new_n1415__spl_),
    .dinb(new_n1420__spl_),
    .dout(new_n1421_)
  );


  anb2
  g1357
  (
    .dina(new_n1415__spl_),
    .dinb(new_n1420__spl_),
    .dout(new_n1422_)
  );


  anb2
  g1358
  (
    .dina(new_n1421__spl_),
    .dinb(new_n1422_),
    .dout(new_n1423_)
  );


  anb1
  g1359
  (
    .dina(new_n1414__spl_),
    .dinb(new_n1423__spl_),
    .dout(new_n1424_)
  );


  anb2
  g1360
  (
    .dina(new_n1414__spl_),
    .dinb(new_n1423__spl_),
    .dout(new_n1425_)
  );


  nab1
  g1361
  (
    .dina(new_n1424__spl_),
    .dinb(new_n1425_),
    .dout(new_n1426_)
  );


  anb2
  g1362
  (
    .dina(new_n1413__spl_),
    .dinb(new_n1426__spl_),
    .dout(new_n1427_)
  );


  anb1
  g1363
  (
    .dina(new_n1413__spl_),
    .dinb(new_n1426__spl_),
    .dout(new_n1428_)
  );


  nab2
  g1364
  (
    .dina(new_n1427__spl_),
    .dinb(new_n1428_),
    .dout(new_n1429_)
  );


  anb1
  g1365
  (
    .dina(new_n1412__spl_),
    .dinb(new_n1429__spl_),
    .dout(new_n1430_)
  );


  anb2
  g1366
  (
    .dina(new_n1412__spl_),
    .dinb(new_n1429__spl_),
    .dout(new_n1431_)
  );


  nab1
  g1367
  (
    .dina(new_n1430__spl_),
    .dinb(new_n1431_),
    .dout(new_n1432_)
  );


  anb2
  g1368
  (
    .dina(new_n1411__spl_),
    .dinb(new_n1432__spl_),
    .dout(new_n1433_)
  );


  anb1
  g1369
  (
    .dina(new_n1411__spl_),
    .dinb(new_n1432__spl_),
    .dout(new_n1434_)
  );


  nab2
  g1370
  (
    .dina(new_n1433__spl_),
    .dinb(new_n1434_),
    .dout(new_n1435_)
  );


  anb1
  g1371
  (
    .dina(new_n1410__spl_),
    .dinb(new_n1435__spl_),
    .dout(new_n1436_)
  );


  anb2
  g1372
  (
    .dina(new_n1410__spl_),
    .dinb(new_n1435__spl_),
    .dout(new_n1437_)
  );


  nab1
  g1373
  (
    .dina(new_n1436__spl_),
    .dinb(new_n1437_),
    .dout(new_n1438_)
  );


  anb2
  g1374
  (
    .dina(new_n1409__spl_),
    .dinb(new_n1438__spl_),
    .dout(new_n1439_)
  );


  anb1
  g1375
  (
    .dina(new_n1409__spl_),
    .dinb(new_n1438__spl_),
    .dout(new_n1440_)
  );


  nab2
  g1376
  (
    .dina(new_n1439__spl_),
    .dinb(new_n1440_),
    .dout(new_n1441_)
  );


  anb1
  g1377
  (
    .dina(new_n1408__spl_),
    .dinb(new_n1441__spl_),
    .dout(new_n1442_)
  );


  anb2
  g1378
  (
    .dina(new_n1408__spl_),
    .dinb(new_n1441__spl_),
    .dout(new_n1443_)
  );


  nab1
  g1379
  (
    .dina(new_n1442__spl_),
    .dinb(new_n1443_),
    .dout(new_n1444_)
  );


  anb2
  g1380
  (
    .dina(new_n1407__spl_),
    .dinb(new_n1444__spl_),
    .dout(new_n1445_)
  );


  anb1
  g1381
  (
    .dina(new_n1407__spl_),
    .dinb(new_n1444__spl_),
    .dout(new_n1446_)
  );


  nab2
  g1382
  (
    .dina(new_n1445__spl_),
    .dinb(new_n1446_),
    .dout(new_n1447_)
  );


  anb1
  g1383
  (
    .dina(new_n1406__spl_),
    .dinb(new_n1447__spl_),
    .dout(new_n1448_)
  );


  anb2
  g1384
  (
    .dina(new_n1406__spl_),
    .dinb(new_n1447__spl_),
    .dout(new_n1449_)
  );


  nab1
  g1385
  (
    .dina(new_n1448__spl_),
    .dinb(new_n1449_),
    .dout(new_n1450_)
  );


  anb2
  g1386
  (
    .dina(new_n1405__spl_),
    .dinb(new_n1450__spl_),
    .dout(new_n1451_)
  );


  anb1
  g1387
  (
    .dina(new_n1405__spl_),
    .dinb(new_n1450__spl_),
    .dout(new_n1452_)
  );


  nab2
  g1388
  (
    .dina(new_n1451__spl_),
    .dinb(new_n1452_),
    .dout(new_n1453_)
  );


  anb1
  g1389
  (
    .dina(new_n1404__spl_),
    .dinb(new_n1453__spl_),
    .dout(new_n1454_)
  );


  anb2
  g1390
  (
    .dina(new_n1404__spl_),
    .dinb(new_n1453__spl_),
    .dout(new_n1455_)
  );


  nab1
  g1391
  (
    .dina(new_n1454__spl_),
    .dinb(new_n1455_),
    .dout(new_n1456_)
  );


  anb2
  g1392
  (
    .dina(new_n1403__spl_),
    .dinb(new_n1456__spl_),
    .dout(new_n1457_)
  );


  anb1
  g1393
  (
    .dina(new_n1403__spl_),
    .dinb(new_n1456__spl_),
    .dout(new_n1458_)
  );


  nab2
  g1394
  (
    .dina(new_n1457__spl_),
    .dinb(new_n1458_),
    .dout(new_n1459_)
  );


  anb1
  g1395
  (
    .dina(new_n1402__spl_),
    .dinb(new_n1459__spl_),
    .dout(new_n1460_)
  );


  anb2
  g1396
  (
    .dina(new_n1402__spl_),
    .dinb(new_n1459__spl_),
    .dout(new_n1461_)
  );


  anb2
  g1397
  (
    .dina(new_n1460__spl_),
    .dinb(new_n1461_),
    .dout(new_n1462_)
  );


  anb1
  g1398
  (
    .dina(new_n1401__spl_),
    .dinb(new_n1462__spl_),
    .dout(new_n1463_)
  );


  anb2
  g1399
  (
    .dina(new_n1401__spl_),
    .dinb(new_n1462__spl_),
    .dout(new_n1464_)
  );


  anb2
  g1400
  (
    .dina(new_n1463__spl_),
    .dinb(new_n1464_),
    .dout(new_n1465_)
  );


  anb1
  g1401
  (
    .dina(new_n1400__spl_),
    .dinb(new_n1465__spl_),
    .dout(new_n1466_)
  );


  anb2
  g1402
  (
    .dina(new_n1400__spl_),
    .dinb(new_n1465__spl_),
    .dout(new_n1467_)
  );


  anb2
  g1403
  (
    .dina(new_n1466__spl_),
    .dinb(new_n1467_),
    .dout(new_n1468_)
  );


  anb1
  g1404
  (
    .dina(new_n1399__spl_),
    .dinb(new_n1468__spl_),
    .dout(new_n1469_)
  );


  anb2
  g1405
  (
    .dina(new_n1399__spl_),
    .dinb(new_n1468__spl_),
    .dout(new_n1470_)
  );


  anb2
  g1406
  (
    .dina(new_n1469__spl_),
    .dinb(new_n1470_),
    .dout(new_n1471_)
  );


  anb1
  g1407
  (
    .dina(new_n1398__spl_),
    .dinb(new_n1471__spl_),
    .dout(new_n1472_)
  );


  anb2
  g1408
  (
    .dina(new_n1398__spl_),
    .dinb(new_n1471__spl_),
    .dout(new_n1473_)
  );


  anb2
  g1409
  (
    .dina(new_n1472__spl_),
    .dinb(new_n1473_),
    .dout(new_n1474_)
  );


  anb1
  g1410
  (
    .dina(new_n1397__spl_),
    .dinb(new_n1474__spl_),
    .dout(new_n1475_)
  );


  anb2
  g1411
  (
    .dina(new_n1397__spl_),
    .dinb(new_n1474__spl_),
    .dout(new_n1476_)
  );


  anb2
  g1412
  (
    .dina(new_n1475__spl_),
    .dinb(new_n1476_),
    .dout(new_n1477_)
  );


  anb1
  g1413
  (
    .dina(new_n1396__spl_),
    .dinb(new_n1477__spl_),
    .dout(new_n1478_)
  );


  anb2
  g1414
  (
    .dina(new_n1396__spl_),
    .dinb(new_n1477__spl_),
    .dout(new_n1479_)
  );


  anb2
  g1415
  (
    .dina(new_n1478__spl_),
    .dinb(new_n1479_),
    .dout(new_n1480_)
  );


  anb1
  g1416
  (
    .dina(new_n1395__spl_),
    .dinb(new_n1480__spl_),
    .dout(new_n1481_)
  );


  anb2
  g1417
  (
    .dina(new_n1395__spl_),
    .dinb(new_n1480__spl_),
    .dout(new_n1482_)
  );


  anb2
  g1418
  (
    .dina(new_n1481__spl_),
    .dinb(new_n1482_),
    .dout(G6277)
  );


  and2
  g1419
  (
    .dina(new_n1478__spl_),
    .dinb(new_n1481__spl_),
    .dout(new_n1484_)
  );


  and2
  g1420
  (
    .dina(new_n1472__spl_),
    .dinb(new_n1475__spl_),
    .dout(new_n1485_)
  );


  nor2
  g1421
  (
    .dina(G7_spl_111),
    .dinb(G32_spl_011),
    .dout(new_n1486_)
  );


  and2
  g1422
  (
    .dina(new_n1466__spl_),
    .dinb(new_n1469__spl_),
    .dout(new_n1487_)
  );


  nor2
  g1423
  (
    .dina(G8_spl_111),
    .dinb(G31_spl_011),
    .dout(new_n1488_)
  );


  and2
  g1424
  (
    .dina(new_n1460__spl_),
    .dinb(new_n1463__spl_),
    .dout(new_n1489_)
  );


  nor2
  g1425
  (
    .dina(G9_spl_110),
    .dinb(G30_spl_100),
    .dout(new_n1490_)
  );


  anb2
  g1426
  (
    .dina(new_n1454__spl_),
    .dinb(new_n1457__spl_),
    .dout(new_n1491_)
  );


  and1
  g1427
  (
    .dina(G10_spl_110),
    .dinb(G29_spl_100),
    .dout(new_n1492_)
  );


  anb2
  g1428
  (
    .dina(new_n1448__spl_),
    .dinb(new_n1451__spl_),
    .dout(new_n1493_)
  );


  and1
  g1429
  (
    .dina(G11_spl_101),
    .dinb(G28_spl_101),
    .dout(new_n1494_)
  );


  anb2
  g1430
  (
    .dina(new_n1442__spl_),
    .dinb(new_n1445__spl_),
    .dout(new_n1495_)
  );


  and1
  g1431
  (
    .dina(G12_spl_101),
    .dinb(G27_spl_101),
    .dout(new_n1496_)
  );


  anb2
  g1432
  (
    .dina(new_n1436__spl_),
    .dinb(new_n1439__spl_),
    .dout(new_n1497_)
  );


  and1
  g1433
  (
    .dina(G13_spl_100),
    .dinb(G26_spl_110),
    .dout(new_n1498_)
  );


  anb2
  g1434
  (
    .dina(new_n1430__spl_),
    .dinb(new_n1433__spl_),
    .dout(new_n1499_)
  );


  and1
  g1435
  (
    .dina(G14_spl_100),
    .dinb(G25_spl_110),
    .dout(new_n1500_)
  );


  anb2
  g1436
  (
    .dina(new_n1424__spl_),
    .dinb(new_n1427__spl_),
    .dout(new_n1501_)
  );


  and1
  g1437
  (
    .dina(G15_spl_011),
    .dinb(G24_spl_111),
    .dout(new_n1502_)
  );


  nor2
  g1438
  (
    .dina(G16_spl_011),
    .dinb(G23_spl_111),
    .dout(new_n1503_)
  );


  anb1
  g1439
  (
    .dina(new_n1418__spl_),
    .dinb(new_n1421__spl_),
    .dout(new_n1504_)
  );


  anb1
  g1440
  (
    .dina(new_n1503__spl_),
    .dinb(new_n1504__spl_),
    .dout(new_n1505_)
  );


  anb2
  g1441
  (
    .dina(new_n1503__spl_),
    .dinb(new_n1504__spl_),
    .dout(new_n1506_)
  );


  nab1
  g1442
  (
    .dina(new_n1505__spl_),
    .dinb(new_n1506_),
    .dout(new_n1507_)
  );


  anb2
  g1443
  (
    .dina(new_n1502__spl_),
    .dinb(new_n1507__spl_),
    .dout(new_n1508_)
  );


  anb1
  g1444
  (
    .dina(new_n1502__spl_),
    .dinb(new_n1507__spl_),
    .dout(new_n1509_)
  );


  nab2
  g1445
  (
    .dina(new_n1508__spl_),
    .dinb(new_n1509_),
    .dout(new_n1510_)
  );


  anb1
  g1446
  (
    .dina(new_n1501__spl_),
    .dinb(new_n1510__spl_),
    .dout(new_n1511_)
  );


  anb2
  g1447
  (
    .dina(new_n1501__spl_),
    .dinb(new_n1510__spl_),
    .dout(new_n1512_)
  );


  nab1
  g1448
  (
    .dina(new_n1511__spl_),
    .dinb(new_n1512_),
    .dout(new_n1513_)
  );


  anb2
  g1449
  (
    .dina(new_n1500__spl_),
    .dinb(new_n1513__spl_),
    .dout(new_n1514_)
  );


  anb1
  g1450
  (
    .dina(new_n1500__spl_),
    .dinb(new_n1513__spl_),
    .dout(new_n1515_)
  );


  nab2
  g1451
  (
    .dina(new_n1514__spl_),
    .dinb(new_n1515_),
    .dout(new_n1516_)
  );


  anb1
  g1452
  (
    .dina(new_n1499__spl_),
    .dinb(new_n1516__spl_),
    .dout(new_n1517_)
  );


  anb2
  g1453
  (
    .dina(new_n1499__spl_),
    .dinb(new_n1516__spl_),
    .dout(new_n1518_)
  );


  nab1
  g1454
  (
    .dina(new_n1517__spl_),
    .dinb(new_n1518_),
    .dout(new_n1519_)
  );


  anb2
  g1455
  (
    .dina(new_n1498__spl_),
    .dinb(new_n1519__spl_),
    .dout(new_n1520_)
  );


  anb1
  g1456
  (
    .dina(new_n1498__spl_),
    .dinb(new_n1519__spl_),
    .dout(new_n1521_)
  );


  nab2
  g1457
  (
    .dina(new_n1520__spl_),
    .dinb(new_n1521_),
    .dout(new_n1522_)
  );


  anb1
  g1458
  (
    .dina(new_n1497__spl_),
    .dinb(new_n1522__spl_),
    .dout(new_n1523_)
  );


  anb2
  g1459
  (
    .dina(new_n1497__spl_),
    .dinb(new_n1522__spl_),
    .dout(new_n1524_)
  );


  nab1
  g1460
  (
    .dina(new_n1523__spl_),
    .dinb(new_n1524_),
    .dout(new_n1525_)
  );


  anb2
  g1461
  (
    .dina(new_n1496__spl_),
    .dinb(new_n1525__spl_),
    .dout(new_n1526_)
  );


  anb1
  g1462
  (
    .dina(new_n1496__spl_),
    .dinb(new_n1525__spl_),
    .dout(new_n1527_)
  );


  nab2
  g1463
  (
    .dina(new_n1526__spl_),
    .dinb(new_n1527_),
    .dout(new_n1528_)
  );


  anb1
  g1464
  (
    .dina(new_n1495__spl_),
    .dinb(new_n1528__spl_),
    .dout(new_n1529_)
  );


  anb2
  g1465
  (
    .dina(new_n1495__spl_),
    .dinb(new_n1528__spl_),
    .dout(new_n1530_)
  );


  nab1
  g1466
  (
    .dina(new_n1529__spl_),
    .dinb(new_n1530_),
    .dout(new_n1531_)
  );


  anb2
  g1467
  (
    .dina(new_n1494__spl_),
    .dinb(new_n1531__spl_),
    .dout(new_n1532_)
  );


  anb1
  g1468
  (
    .dina(new_n1494__spl_),
    .dinb(new_n1531__spl_),
    .dout(new_n1533_)
  );


  nab2
  g1469
  (
    .dina(new_n1532__spl_),
    .dinb(new_n1533_),
    .dout(new_n1534_)
  );


  anb1
  g1470
  (
    .dina(new_n1493__spl_),
    .dinb(new_n1534__spl_),
    .dout(new_n1535_)
  );


  anb2
  g1471
  (
    .dina(new_n1493__spl_),
    .dinb(new_n1534__spl_),
    .dout(new_n1536_)
  );


  nab1
  g1472
  (
    .dina(new_n1535__spl_),
    .dinb(new_n1536_),
    .dout(new_n1537_)
  );


  anb2
  g1473
  (
    .dina(new_n1492__spl_),
    .dinb(new_n1537__spl_),
    .dout(new_n1538_)
  );


  anb1
  g1474
  (
    .dina(new_n1492__spl_),
    .dinb(new_n1537__spl_),
    .dout(new_n1539_)
  );


  nab2
  g1475
  (
    .dina(new_n1538__spl_),
    .dinb(new_n1539_),
    .dout(new_n1540_)
  );


  anb1
  g1476
  (
    .dina(new_n1491__spl_),
    .dinb(new_n1540__spl_),
    .dout(new_n1541_)
  );


  anb2
  g1477
  (
    .dina(new_n1491__spl_),
    .dinb(new_n1540__spl_),
    .dout(new_n1542_)
  );


  anb2
  g1478
  (
    .dina(new_n1541__spl_),
    .dinb(new_n1542_),
    .dout(new_n1543_)
  );


  anb1
  g1479
  (
    .dina(new_n1490__spl_),
    .dinb(new_n1543__spl_),
    .dout(new_n1544_)
  );


  anb2
  g1480
  (
    .dina(new_n1490__spl_),
    .dinb(new_n1543__spl_),
    .dout(new_n1545_)
  );


  anb2
  g1481
  (
    .dina(new_n1544__spl_),
    .dinb(new_n1545_),
    .dout(new_n1546_)
  );


  anb1
  g1482
  (
    .dina(new_n1489__spl_),
    .dinb(new_n1546__spl_),
    .dout(new_n1547_)
  );


  anb2
  g1483
  (
    .dina(new_n1489__spl_),
    .dinb(new_n1546__spl_),
    .dout(new_n1548_)
  );


  anb2
  g1484
  (
    .dina(new_n1547__spl_),
    .dinb(new_n1548_),
    .dout(new_n1549_)
  );


  anb1
  g1485
  (
    .dina(new_n1488__spl_),
    .dinb(new_n1549__spl_),
    .dout(new_n1550_)
  );


  anb2
  g1486
  (
    .dina(new_n1488__spl_),
    .dinb(new_n1549__spl_),
    .dout(new_n1551_)
  );


  anb2
  g1487
  (
    .dina(new_n1550__spl_),
    .dinb(new_n1551_),
    .dout(new_n1552_)
  );


  anb1
  g1488
  (
    .dina(new_n1487__spl_),
    .dinb(new_n1552__spl_),
    .dout(new_n1553_)
  );


  anb2
  g1489
  (
    .dina(new_n1487__spl_),
    .dinb(new_n1552__spl_),
    .dout(new_n1554_)
  );


  anb2
  g1490
  (
    .dina(new_n1553__spl_),
    .dinb(new_n1554_),
    .dout(new_n1555_)
  );


  anb1
  g1491
  (
    .dina(new_n1486__spl_),
    .dinb(new_n1555__spl_),
    .dout(new_n1556_)
  );


  anb2
  g1492
  (
    .dina(new_n1486__spl_),
    .dinb(new_n1555__spl_),
    .dout(new_n1557_)
  );


  anb2
  g1493
  (
    .dina(new_n1556__spl_),
    .dinb(new_n1557_),
    .dout(new_n1558_)
  );


  anb1
  g1494
  (
    .dina(new_n1485__spl_),
    .dinb(new_n1558__spl_),
    .dout(new_n1559_)
  );


  anb2
  g1495
  (
    .dina(new_n1485__spl_),
    .dinb(new_n1558__spl_),
    .dout(new_n1560_)
  );


  anb2
  g1496
  (
    .dina(new_n1559__spl_),
    .dinb(new_n1560_),
    .dout(new_n1561_)
  );


  anb1
  g1497
  (
    .dina(new_n1484__spl_),
    .dinb(new_n1561__spl_),
    .dout(new_n1562_)
  );


  anb2
  g1498
  (
    .dina(new_n1484__spl_),
    .dinb(new_n1561__spl_),
    .dout(new_n1563_)
  );


  anb2
  g1499
  (
    .dina(new_n1562__spl_),
    .dinb(new_n1563_),
    .dout(G6278)
  );


  and2
  g1500
  (
    .dina(new_n1559__spl_),
    .dinb(new_n1562__spl_),
    .dout(new_n1565_)
  );


  and2
  g1501
  (
    .dina(new_n1553__spl_),
    .dinb(new_n1556__spl_),
    .dout(new_n1566_)
  );


  nor2
  g1502
  (
    .dina(G8_spl_111),
    .dinb(G32_spl_011),
    .dout(new_n1567_)
  );


  and2
  g1503
  (
    .dina(new_n1547__spl_),
    .dinb(new_n1550__spl_),
    .dout(new_n1568_)
  );


  nor2
  g1504
  (
    .dina(G9_spl_111),
    .dinb(G31_spl_100),
    .dout(new_n1569_)
  );


  and2
  g1505
  (
    .dina(new_n1541__spl_),
    .dinb(new_n1544__spl_),
    .dout(new_n1570_)
  );


  nor2
  g1506
  (
    .dina(G10_spl_110),
    .dinb(G30_spl_100),
    .dout(new_n1571_)
  );


  anb2
  g1507
  (
    .dina(new_n1535__spl_),
    .dinb(new_n1538__spl_),
    .dout(new_n1572_)
  );


  and1
  g1508
  (
    .dina(G11_spl_110),
    .dinb(G29_spl_101),
    .dout(new_n1573_)
  );


  anb2
  g1509
  (
    .dina(new_n1529__spl_),
    .dinb(new_n1532__spl_),
    .dout(new_n1574_)
  );


  and1
  g1510
  (
    .dina(G12_spl_101),
    .dinb(G28_spl_101),
    .dout(new_n1575_)
  );


  anb2
  g1511
  (
    .dina(new_n1523__spl_),
    .dinb(new_n1526__spl_),
    .dout(new_n1576_)
  );


  and1
  g1512
  (
    .dina(G13_spl_101),
    .dinb(G27_spl_110),
    .dout(new_n1577_)
  );


  anb2
  g1513
  (
    .dina(new_n1517__spl_),
    .dinb(new_n1520__spl_),
    .dout(new_n1578_)
  );


  and1
  g1514
  (
    .dina(G14_spl_100),
    .dinb(G26_spl_110),
    .dout(new_n1579_)
  );


  anb2
  g1515
  (
    .dina(new_n1511__spl_),
    .dinb(new_n1514__spl_),
    .dout(new_n1580_)
  );


  nor2
  g1516
  (
    .dina(G15_spl_100),
    .dinb(G25_spl_111),
    .dout(new_n1581_)
  );


  and1
  g1517
  (
    .dina(G16_spl_011),
    .dinb(G24_spl_111),
    .dout(new_n1582_)
  );


  anb2
  g1518
  (
    .dina(new_n1505__spl_),
    .dinb(new_n1508__spl_),
    .dout(new_n1583_)
  );


  anb2
  g1519
  (
    .dina(new_n1582__spl_),
    .dinb(new_n1583__spl_),
    .dout(new_n1584_)
  );


  anb1
  g1520
  (
    .dina(new_n1582__spl_),
    .dinb(new_n1583__spl_),
    .dout(new_n1585_)
  );


  nab2
  g1521
  (
    .dina(new_n1584__spl_),
    .dinb(new_n1585_),
    .dout(new_n1586_)
  );


  anb1
  g1522
  (
    .dina(new_n1581__spl_),
    .dinb(new_n1586__spl_),
    .dout(new_n1587_)
  );


  anb2
  g1523
  (
    .dina(new_n1581__spl_),
    .dinb(new_n1586__spl_),
    .dout(new_n1588_)
  );


  anb2
  g1524
  (
    .dina(new_n1587__spl_),
    .dinb(new_n1588_),
    .dout(new_n1589_)
  );


  anb1
  g1525
  (
    .dina(new_n1580__spl_),
    .dinb(new_n1589__spl_),
    .dout(new_n1590_)
  );


  anb2
  g1526
  (
    .dina(new_n1580__spl_),
    .dinb(new_n1589__spl_),
    .dout(new_n1591_)
  );


  nab1
  g1527
  (
    .dina(new_n1590__spl_),
    .dinb(new_n1591_),
    .dout(new_n1592_)
  );


  anb2
  g1528
  (
    .dina(new_n1579__spl_),
    .dinb(new_n1592__spl_),
    .dout(new_n1593_)
  );


  anb1
  g1529
  (
    .dina(new_n1579__spl_),
    .dinb(new_n1592__spl_),
    .dout(new_n1594_)
  );


  nab2
  g1530
  (
    .dina(new_n1593__spl_),
    .dinb(new_n1594_),
    .dout(new_n1595_)
  );


  anb1
  g1531
  (
    .dina(new_n1578__spl_),
    .dinb(new_n1595__spl_),
    .dout(new_n1596_)
  );


  anb2
  g1532
  (
    .dina(new_n1578__spl_),
    .dinb(new_n1595__spl_),
    .dout(new_n1597_)
  );


  nab1
  g1533
  (
    .dina(new_n1596__spl_),
    .dinb(new_n1597_),
    .dout(new_n1598_)
  );


  anb2
  g1534
  (
    .dina(new_n1577__spl_),
    .dinb(new_n1598__spl_),
    .dout(new_n1599_)
  );


  anb1
  g1535
  (
    .dina(new_n1577__spl_),
    .dinb(new_n1598__spl_),
    .dout(new_n1600_)
  );


  nab2
  g1536
  (
    .dina(new_n1599__spl_),
    .dinb(new_n1600_),
    .dout(new_n1601_)
  );


  anb1
  g1537
  (
    .dina(new_n1576__spl_),
    .dinb(new_n1601__spl_),
    .dout(new_n1602_)
  );


  anb2
  g1538
  (
    .dina(new_n1576__spl_),
    .dinb(new_n1601__spl_),
    .dout(new_n1603_)
  );


  nab1
  g1539
  (
    .dina(new_n1602__spl_),
    .dinb(new_n1603_),
    .dout(new_n1604_)
  );


  anb2
  g1540
  (
    .dina(new_n1575__spl_),
    .dinb(new_n1604__spl_),
    .dout(new_n1605_)
  );


  anb1
  g1541
  (
    .dina(new_n1575__spl_),
    .dinb(new_n1604__spl_),
    .dout(new_n1606_)
  );


  nab2
  g1542
  (
    .dina(new_n1605__spl_),
    .dinb(new_n1606_),
    .dout(new_n1607_)
  );


  anb1
  g1543
  (
    .dina(new_n1574__spl_),
    .dinb(new_n1607__spl_),
    .dout(new_n1608_)
  );


  anb2
  g1544
  (
    .dina(new_n1574__spl_),
    .dinb(new_n1607__spl_),
    .dout(new_n1609_)
  );


  nab1
  g1545
  (
    .dina(new_n1608__spl_),
    .dinb(new_n1609_),
    .dout(new_n1610_)
  );


  anb2
  g1546
  (
    .dina(new_n1573__spl_),
    .dinb(new_n1610__spl_),
    .dout(new_n1611_)
  );


  anb1
  g1547
  (
    .dina(new_n1573__spl_),
    .dinb(new_n1610__spl_),
    .dout(new_n1612_)
  );


  nab2
  g1548
  (
    .dina(new_n1611__spl_),
    .dinb(new_n1612_),
    .dout(new_n1613_)
  );


  anb1
  g1549
  (
    .dina(new_n1572__spl_),
    .dinb(new_n1613__spl_),
    .dout(new_n1614_)
  );


  anb2
  g1550
  (
    .dina(new_n1572__spl_),
    .dinb(new_n1613__spl_),
    .dout(new_n1615_)
  );


  anb2
  g1551
  (
    .dina(new_n1614__spl_),
    .dinb(new_n1615_),
    .dout(new_n1616_)
  );


  anb1
  g1552
  (
    .dina(new_n1571__spl_),
    .dinb(new_n1616__spl_),
    .dout(new_n1617_)
  );


  anb2
  g1553
  (
    .dina(new_n1571__spl_),
    .dinb(new_n1616__spl_),
    .dout(new_n1618_)
  );


  anb2
  g1554
  (
    .dina(new_n1617__spl_),
    .dinb(new_n1618_),
    .dout(new_n1619_)
  );


  anb1
  g1555
  (
    .dina(new_n1570__spl_),
    .dinb(new_n1619__spl_),
    .dout(new_n1620_)
  );


  anb2
  g1556
  (
    .dina(new_n1570__spl_),
    .dinb(new_n1619__spl_),
    .dout(new_n1621_)
  );


  anb2
  g1557
  (
    .dina(new_n1620__spl_),
    .dinb(new_n1621_),
    .dout(new_n1622_)
  );


  anb1
  g1558
  (
    .dina(new_n1569__spl_),
    .dinb(new_n1622__spl_),
    .dout(new_n1623_)
  );


  anb2
  g1559
  (
    .dina(new_n1569__spl_),
    .dinb(new_n1622__spl_),
    .dout(new_n1624_)
  );


  anb2
  g1560
  (
    .dina(new_n1623__spl_),
    .dinb(new_n1624_),
    .dout(new_n1625_)
  );


  anb1
  g1561
  (
    .dina(new_n1568__spl_),
    .dinb(new_n1625__spl_),
    .dout(new_n1626_)
  );


  anb2
  g1562
  (
    .dina(new_n1568__spl_),
    .dinb(new_n1625__spl_),
    .dout(new_n1627_)
  );


  anb2
  g1563
  (
    .dina(new_n1626__spl_),
    .dinb(new_n1627_),
    .dout(new_n1628_)
  );


  anb1
  g1564
  (
    .dina(new_n1567__spl_),
    .dinb(new_n1628__spl_),
    .dout(new_n1629_)
  );


  anb2
  g1565
  (
    .dina(new_n1567__spl_),
    .dinb(new_n1628__spl_),
    .dout(new_n1630_)
  );


  anb2
  g1566
  (
    .dina(new_n1629__spl_),
    .dinb(new_n1630_),
    .dout(new_n1631_)
  );


  anb1
  g1567
  (
    .dina(new_n1566__spl_),
    .dinb(new_n1631__spl_),
    .dout(new_n1632_)
  );


  anb2
  g1568
  (
    .dina(new_n1566__spl_),
    .dinb(new_n1631__spl_),
    .dout(new_n1633_)
  );


  anb2
  g1569
  (
    .dina(new_n1632__spl_),
    .dinb(new_n1633_),
    .dout(new_n1634_)
  );


  anb1
  g1570
  (
    .dina(new_n1565__spl_),
    .dinb(new_n1634__spl_),
    .dout(new_n1635_)
  );


  anb2
  g1571
  (
    .dina(new_n1565__spl_),
    .dinb(new_n1634__spl_),
    .dout(new_n1636_)
  );


  anb2
  g1572
  (
    .dina(new_n1635__spl_),
    .dinb(new_n1636_),
    .dout(G6279)
  );


  and2
  g1573
  (
    .dina(new_n1632__spl_),
    .dinb(new_n1635__spl_),
    .dout(new_n1638_)
  );


  and2
  g1574
  (
    .dina(new_n1626__spl_),
    .dinb(new_n1629__spl_),
    .dout(new_n1639_)
  );


  nor2
  g1575
  (
    .dina(G9_spl_111),
    .dinb(G32_spl_100),
    .dout(new_n1640_)
  );


  and2
  g1576
  (
    .dina(new_n1620__spl_),
    .dinb(new_n1623__spl_),
    .dout(new_n1641_)
  );


  nor2
  g1577
  (
    .dina(G10_spl_111),
    .dinb(G31_spl_100),
    .dout(new_n1642_)
  );


  and2
  g1578
  (
    .dina(new_n1614__spl_),
    .dinb(new_n1617__spl_),
    .dout(new_n1643_)
  );


  nor2
  g1579
  (
    .dina(G11_spl_110),
    .dinb(G30_spl_101),
    .dout(new_n1644_)
  );


  anb2
  g1580
  (
    .dina(new_n1608__spl_),
    .dinb(new_n1611__spl_),
    .dout(new_n1645_)
  );


  and1
  g1581
  (
    .dina(G12_spl_110),
    .dinb(G29_spl_101),
    .dout(new_n1646_)
  );


  anb2
  g1582
  (
    .dina(new_n1602__spl_),
    .dinb(new_n1605__spl_),
    .dout(new_n1647_)
  );


  and1
  g1583
  (
    .dina(G13_spl_101),
    .dinb(G28_spl_110),
    .dout(new_n1648_)
  );


  anb2
  g1584
  (
    .dina(new_n1596__spl_),
    .dinb(new_n1599__spl_),
    .dout(new_n1649_)
  );


  and1
  g1585
  (
    .dina(G14_spl_101),
    .dinb(G27_spl_110),
    .dout(new_n1650_)
  );


  anb2
  g1586
  (
    .dina(new_n1590__spl_),
    .dinb(new_n1593__spl_),
    .dout(new_n1651_)
  );


  and1
  g1587
  (
    .dina(G15_spl_100),
    .dinb(G26_spl_111),
    .dout(new_n1652_)
  );


  nor2
  g1588
  (
    .dina(G16_spl_100),
    .dinb(G25_spl_111),
    .dout(new_n1653_)
  );


  anb1
  g1589
  (
    .dina(new_n1584__spl_),
    .dinb(new_n1587__spl_),
    .dout(new_n1654_)
  );


  anb1
  g1590
  (
    .dina(new_n1653__spl_),
    .dinb(new_n1654__spl_),
    .dout(new_n1655_)
  );


  anb2
  g1591
  (
    .dina(new_n1653__spl_),
    .dinb(new_n1654__spl_),
    .dout(new_n1656_)
  );


  nab1
  g1592
  (
    .dina(new_n1655__spl_),
    .dinb(new_n1656_),
    .dout(new_n1657_)
  );


  anb2
  g1593
  (
    .dina(new_n1652__spl_),
    .dinb(new_n1657__spl_),
    .dout(new_n1658_)
  );


  anb1
  g1594
  (
    .dina(new_n1652__spl_),
    .dinb(new_n1657__spl_),
    .dout(new_n1659_)
  );


  nab2
  g1595
  (
    .dina(new_n1658__spl_),
    .dinb(new_n1659_),
    .dout(new_n1660_)
  );


  anb1
  g1596
  (
    .dina(new_n1651__spl_),
    .dinb(new_n1660__spl_),
    .dout(new_n1661_)
  );


  anb2
  g1597
  (
    .dina(new_n1651__spl_),
    .dinb(new_n1660__spl_),
    .dout(new_n1662_)
  );


  nab1
  g1598
  (
    .dina(new_n1661__spl_),
    .dinb(new_n1662_),
    .dout(new_n1663_)
  );


  anb2
  g1599
  (
    .dina(new_n1650__spl_),
    .dinb(new_n1663__spl_),
    .dout(new_n1664_)
  );


  anb1
  g1600
  (
    .dina(new_n1650__spl_),
    .dinb(new_n1663__spl_),
    .dout(new_n1665_)
  );


  nab2
  g1601
  (
    .dina(new_n1664__spl_),
    .dinb(new_n1665_),
    .dout(new_n1666_)
  );


  anb1
  g1602
  (
    .dina(new_n1649__spl_),
    .dinb(new_n1666__spl_),
    .dout(new_n1667_)
  );


  anb2
  g1603
  (
    .dina(new_n1649__spl_),
    .dinb(new_n1666__spl_),
    .dout(new_n1668_)
  );


  nab1
  g1604
  (
    .dina(new_n1667__spl_),
    .dinb(new_n1668_),
    .dout(new_n1669_)
  );


  anb2
  g1605
  (
    .dina(new_n1648__spl_),
    .dinb(new_n1669__spl_),
    .dout(new_n1670_)
  );


  anb1
  g1606
  (
    .dina(new_n1648__spl_),
    .dinb(new_n1669__spl_),
    .dout(new_n1671_)
  );


  nab2
  g1607
  (
    .dina(new_n1670__spl_),
    .dinb(new_n1671_),
    .dout(new_n1672_)
  );


  anb1
  g1608
  (
    .dina(new_n1647__spl_),
    .dinb(new_n1672__spl_),
    .dout(new_n1673_)
  );


  anb2
  g1609
  (
    .dina(new_n1647__spl_),
    .dinb(new_n1672__spl_),
    .dout(new_n1674_)
  );


  nab1
  g1610
  (
    .dina(new_n1673__spl_),
    .dinb(new_n1674_),
    .dout(new_n1675_)
  );


  anb2
  g1611
  (
    .dina(new_n1646__spl_),
    .dinb(new_n1675__spl_),
    .dout(new_n1676_)
  );


  anb1
  g1612
  (
    .dina(new_n1646__spl_),
    .dinb(new_n1675__spl_),
    .dout(new_n1677_)
  );


  nab2
  g1613
  (
    .dina(new_n1676__spl_),
    .dinb(new_n1677_),
    .dout(new_n1678_)
  );


  anb1
  g1614
  (
    .dina(new_n1645__spl_),
    .dinb(new_n1678__spl_),
    .dout(new_n1679_)
  );


  anb2
  g1615
  (
    .dina(new_n1645__spl_),
    .dinb(new_n1678__spl_),
    .dout(new_n1680_)
  );


  anb2
  g1616
  (
    .dina(new_n1679__spl_),
    .dinb(new_n1680_),
    .dout(new_n1681_)
  );


  anb1
  g1617
  (
    .dina(new_n1644__spl_),
    .dinb(new_n1681__spl_),
    .dout(new_n1682_)
  );


  anb2
  g1618
  (
    .dina(new_n1644__spl_),
    .dinb(new_n1681__spl_),
    .dout(new_n1683_)
  );


  anb2
  g1619
  (
    .dina(new_n1682__spl_),
    .dinb(new_n1683_),
    .dout(new_n1684_)
  );


  anb1
  g1620
  (
    .dina(new_n1643__spl_),
    .dinb(new_n1684__spl_),
    .dout(new_n1685_)
  );


  anb2
  g1621
  (
    .dina(new_n1643__spl_),
    .dinb(new_n1684__spl_),
    .dout(new_n1686_)
  );


  anb2
  g1622
  (
    .dina(new_n1685__spl_),
    .dinb(new_n1686_),
    .dout(new_n1687_)
  );


  anb1
  g1623
  (
    .dina(new_n1642__spl_),
    .dinb(new_n1687__spl_),
    .dout(new_n1688_)
  );


  anb2
  g1624
  (
    .dina(new_n1642__spl_),
    .dinb(new_n1687__spl_),
    .dout(new_n1689_)
  );


  anb2
  g1625
  (
    .dina(new_n1688__spl_),
    .dinb(new_n1689_),
    .dout(new_n1690_)
  );


  anb1
  g1626
  (
    .dina(new_n1641__spl_),
    .dinb(new_n1690__spl_),
    .dout(new_n1691_)
  );


  anb2
  g1627
  (
    .dina(new_n1641__spl_),
    .dinb(new_n1690__spl_),
    .dout(new_n1692_)
  );


  anb2
  g1628
  (
    .dina(new_n1691__spl_),
    .dinb(new_n1692_),
    .dout(new_n1693_)
  );


  anb1
  g1629
  (
    .dina(new_n1640__spl_),
    .dinb(new_n1693__spl_),
    .dout(new_n1694_)
  );


  anb2
  g1630
  (
    .dina(new_n1640__spl_),
    .dinb(new_n1693__spl_),
    .dout(new_n1695_)
  );


  anb2
  g1631
  (
    .dina(new_n1694__spl_),
    .dinb(new_n1695_),
    .dout(new_n1696_)
  );


  anb1
  g1632
  (
    .dina(new_n1639__spl_),
    .dinb(new_n1696__spl_),
    .dout(new_n1697_)
  );


  anb2
  g1633
  (
    .dina(new_n1639__spl_),
    .dinb(new_n1696__spl_),
    .dout(new_n1698_)
  );


  anb2
  g1634
  (
    .dina(new_n1697__spl_),
    .dinb(new_n1698_),
    .dout(new_n1699_)
  );


  anb1
  g1635
  (
    .dina(new_n1638__spl_),
    .dinb(new_n1699__spl_),
    .dout(new_n1700_)
  );


  anb2
  g1636
  (
    .dina(new_n1638__spl_),
    .dinb(new_n1699__spl_),
    .dout(new_n1701_)
  );


  anb2
  g1637
  (
    .dina(new_n1700__spl_),
    .dinb(new_n1701_),
    .dout(G6280)
  );


  and2
  g1638
  (
    .dina(new_n1697__spl_),
    .dinb(new_n1700__spl_),
    .dout(new_n1703_)
  );


  and2
  g1639
  (
    .dina(new_n1691__spl_),
    .dinb(new_n1694__spl_),
    .dout(new_n1704_)
  );


  nor2
  g1640
  (
    .dina(G10_spl_111),
    .dinb(G32_spl_100),
    .dout(new_n1705_)
  );


  and2
  g1641
  (
    .dina(new_n1685__spl_),
    .dinb(new_n1688__spl_),
    .dout(new_n1706_)
  );


  nor2
  g1642
  (
    .dina(G11_spl_111),
    .dinb(G31_spl_101),
    .dout(new_n1707_)
  );


  and2
  g1643
  (
    .dina(new_n1679__spl_),
    .dinb(new_n1682__spl_),
    .dout(new_n1708_)
  );


  nor2
  g1644
  (
    .dina(G12_spl_110),
    .dinb(G30_spl_101),
    .dout(new_n1709_)
  );


  anb2
  g1645
  (
    .dina(new_n1673__spl_),
    .dinb(new_n1676__spl_),
    .dout(new_n1710_)
  );


  and1
  g1646
  (
    .dina(G13_spl_110),
    .dinb(G29_spl_110),
    .dout(new_n1711_)
  );


  anb2
  g1647
  (
    .dina(new_n1667__spl_),
    .dinb(new_n1670__spl_),
    .dout(new_n1712_)
  );


  and1
  g1648
  (
    .dina(G14_spl_101),
    .dinb(G28_spl_110),
    .dout(new_n1713_)
  );


  anb2
  g1649
  (
    .dina(new_n1661__spl_),
    .dinb(new_n1664__spl_),
    .dout(new_n1714_)
  );


  nor2
  g1650
  (
    .dina(G15_spl_101),
    .dinb(G27_spl_111),
    .dout(new_n1715_)
  );


  and1
  g1651
  (
    .dina(G16_spl_100),
    .dinb(G26_spl_111),
    .dout(new_n1716_)
  );


  anb2
  g1652
  (
    .dina(new_n1655__spl_),
    .dinb(new_n1658__spl_),
    .dout(new_n1717_)
  );


  anb2
  g1653
  (
    .dina(new_n1716__spl_),
    .dinb(new_n1717__spl_),
    .dout(new_n1718_)
  );


  anb1
  g1654
  (
    .dina(new_n1716__spl_),
    .dinb(new_n1717__spl_),
    .dout(new_n1719_)
  );


  nab2
  g1655
  (
    .dina(new_n1718__spl_),
    .dinb(new_n1719_),
    .dout(new_n1720_)
  );


  anb1
  g1656
  (
    .dina(new_n1715__spl_),
    .dinb(new_n1720__spl_),
    .dout(new_n1721_)
  );


  anb2
  g1657
  (
    .dina(new_n1715__spl_),
    .dinb(new_n1720__spl_),
    .dout(new_n1722_)
  );


  anb2
  g1658
  (
    .dina(new_n1721__spl_),
    .dinb(new_n1722_),
    .dout(new_n1723_)
  );


  anb1
  g1659
  (
    .dina(new_n1714__spl_),
    .dinb(new_n1723__spl_),
    .dout(new_n1724_)
  );


  anb2
  g1660
  (
    .dina(new_n1714__spl_),
    .dinb(new_n1723__spl_),
    .dout(new_n1725_)
  );


  nab1
  g1661
  (
    .dina(new_n1724__spl_),
    .dinb(new_n1725_),
    .dout(new_n1726_)
  );


  anb2
  g1662
  (
    .dina(new_n1713__spl_),
    .dinb(new_n1726__spl_),
    .dout(new_n1727_)
  );


  anb1
  g1663
  (
    .dina(new_n1713__spl_),
    .dinb(new_n1726__spl_),
    .dout(new_n1728_)
  );


  nab2
  g1664
  (
    .dina(new_n1727__spl_),
    .dinb(new_n1728_),
    .dout(new_n1729_)
  );


  anb1
  g1665
  (
    .dina(new_n1712__spl_),
    .dinb(new_n1729__spl_),
    .dout(new_n1730_)
  );


  anb2
  g1666
  (
    .dina(new_n1712__spl_),
    .dinb(new_n1729__spl_),
    .dout(new_n1731_)
  );


  nab1
  g1667
  (
    .dina(new_n1730__spl_),
    .dinb(new_n1731_),
    .dout(new_n1732_)
  );


  anb2
  g1668
  (
    .dina(new_n1711__spl_),
    .dinb(new_n1732__spl_),
    .dout(new_n1733_)
  );


  anb1
  g1669
  (
    .dina(new_n1711__spl_),
    .dinb(new_n1732__spl_),
    .dout(new_n1734_)
  );


  nab2
  g1670
  (
    .dina(new_n1733__spl_),
    .dinb(new_n1734_),
    .dout(new_n1735_)
  );


  anb1
  g1671
  (
    .dina(new_n1710__spl_),
    .dinb(new_n1735__spl_),
    .dout(new_n1736_)
  );


  anb2
  g1672
  (
    .dina(new_n1710__spl_),
    .dinb(new_n1735__spl_),
    .dout(new_n1737_)
  );


  anb2
  g1673
  (
    .dina(new_n1736__spl_),
    .dinb(new_n1737_),
    .dout(new_n1738_)
  );


  anb1
  g1674
  (
    .dina(new_n1709__spl_),
    .dinb(new_n1738__spl_),
    .dout(new_n1739_)
  );


  anb2
  g1675
  (
    .dina(new_n1709__spl_),
    .dinb(new_n1738__spl_),
    .dout(new_n1740_)
  );


  anb2
  g1676
  (
    .dina(new_n1739__spl_),
    .dinb(new_n1740_),
    .dout(new_n1741_)
  );


  anb1
  g1677
  (
    .dina(new_n1708__spl_),
    .dinb(new_n1741__spl_),
    .dout(new_n1742_)
  );


  anb2
  g1678
  (
    .dina(new_n1708__spl_),
    .dinb(new_n1741__spl_),
    .dout(new_n1743_)
  );


  anb2
  g1679
  (
    .dina(new_n1742__spl_),
    .dinb(new_n1743_),
    .dout(new_n1744_)
  );


  anb1
  g1680
  (
    .dina(new_n1707__spl_),
    .dinb(new_n1744__spl_),
    .dout(new_n1745_)
  );


  anb2
  g1681
  (
    .dina(new_n1707__spl_),
    .dinb(new_n1744__spl_),
    .dout(new_n1746_)
  );


  anb2
  g1682
  (
    .dina(new_n1745__spl_),
    .dinb(new_n1746_),
    .dout(new_n1747_)
  );


  anb1
  g1683
  (
    .dina(new_n1706__spl_),
    .dinb(new_n1747__spl_),
    .dout(new_n1748_)
  );


  anb2
  g1684
  (
    .dina(new_n1706__spl_),
    .dinb(new_n1747__spl_),
    .dout(new_n1749_)
  );


  anb2
  g1685
  (
    .dina(new_n1748__spl_),
    .dinb(new_n1749_),
    .dout(new_n1750_)
  );


  anb1
  g1686
  (
    .dina(new_n1705__spl_),
    .dinb(new_n1750__spl_),
    .dout(new_n1751_)
  );


  anb2
  g1687
  (
    .dina(new_n1705__spl_),
    .dinb(new_n1750__spl_),
    .dout(new_n1752_)
  );


  anb2
  g1688
  (
    .dina(new_n1751__spl_),
    .dinb(new_n1752_),
    .dout(new_n1753_)
  );


  anb1
  g1689
  (
    .dina(new_n1704__spl_),
    .dinb(new_n1753__spl_),
    .dout(new_n1754_)
  );


  anb2
  g1690
  (
    .dina(new_n1704__spl_),
    .dinb(new_n1753__spl_),
    .dout(new_n1755_)
  );


  anb2
  g1691
  (
    .dina(new_n1754__spl_),
    .dinb(new_n1755_),
    .dout(new_n1756_)
  );


  anb1
  g1692
  (
    .dina(new_n1703__spl_),
    .dinb(new_n1756__spl_),
    .dout(new_n1757_)
  );


  anb2
  g1693
  (
    .dina(new_n1703__spl_),
    .dinb(new_n1756__spl_),
    .dout(new_n1758_)
  );


  anb2
  g1694
  (
    .dina(new_n1757__spl_),
    .dinb(new_n1758_),
    .dout(G6281)
  );


  and2
  g1695
  (
    .dina(new_n1754__spl_),
    .dinb(new_n1757__spl_),
    .dout(new_n1760_)
  );


  and2
  g1696
  (
    .dina(new_n1748__spl_),
    .dinb(new_n1751__spl_),
    .dout(new_n1761_)
  );


  nor2
  g1697
  (
    .dina(G11_spl_111),
    .dinb(G32_spl_101),
    .dout(new_n1762_)
  );


  and2
  g1698
  (
    .dina(new_n1742__spl_),
    .dinb(new_n1745__spl_),
    .dout(new_n1763_)
  );


  nor2
  g1699
  (
    .dina(G12_spl_111),
    .dinb(G31_spl_101),
    .dout(new_n1764_)
  );


  and2
  g1700
  (
    .dina(new_n1736__spl_),
    .dinb(new_n1739__spl_),
    .dout(new_n1765_)
  );


  nor2
  g1701
  (
    .dina(G13_spl_110),
    .dinb(G30_spl_110),
    .dout(new_n1766_)
  );


  anb2
  g1702
  (
    .dina(new_n1730__spl_),
    .dinb(new_n1733__spl_),
    .dout(new_n1767_)
  );


  and1
  g1703
  (
    .dina(G14_spl_110),
    .dinb(G29_spl_110),
    .dout(new_n1768_)
  );


  anb2
  g1704
  (
    .dina(new_n1724__spl_),
    .dinb(new_n1727__spl_),
    .dout(new_n1769_)
  );


  and1
  g1705
  (
    .dina(G15_spl_101),
    .dinb(G28_spl_111),
    .dout(new_n1770_)
  );


  nor2
  g1706
  (
    .dina(G16_spl_101),
    .dinb(G27_spl_111),
    .dout(new_n1771_)
  );


  anb1
  g1707
  (
    .dina(new_n1718__spl_),
    .dinb(new_n1721__spl_),
    .dout(new_n1772_)
  );


  anb1
  g1708
  (
    .dina(new_n1771__spl_),
    .dinb(new_n1772__spl_),
    .dout(new_n1773_)
  );


  anb2
  g1709
  (
    .dina(new_n1771__spl_),
    .dinb(new_n1772__spl_),
    .dout(new_n1774_)
  );


  nab1
  g1710
  (
    .dina(new_n1773__spl_),
    .dinb(new_n1774_),
    .dout(new_n1775_)
  );


  anb2
  g1711
  (
    .dina(new_n1770__spl_),
    .dinb(new_n1775__spl_),
    .dout(new_n1776_)
  );


  anb1
  g1712
  (
    .dina(new_n1770__spl_),
    .dinb(new_n1775__spl_),
    .dout(new_n1777_)
  );


  nab2
  g1713
  (
    .dina(new_n1776__spl_),
    .dinb(new_n1777_),
    .dout(new_n1778_)
  );


  anb1
  g1714
  (
    .dina(new_n1769__spl_),
    .dinb(new_n1778__spl_),
    .dout(new_n1779_)
  );


  anb2
  g1715
  (
    .dina(new_n1769__spl_),
    .dinb(new_n1778__spl_),
    .dout(new_n1780_)
  );


  nab1
  g1716
  (
    .dina(new_n1779__spl_),
    .dinb(new_n1780_),
    .dout(new_n1781_)
  );


  anb2
  g1717
  (
    .dina(new_n1768__spl_),
    .dinb(new_n1781__spl_),
    .dout(new_n1782_)
  );


  anb1
  g1718
  (
    .dina(new_n1768__spl_),
    .dinb(new_n1781__spl_),
    .dout(new_n1783_)
  );


  nab2
  g1719
  (
    .dina(new_n1782__spl_),
    .dinb(new_n1783_),
    .dout(new_n1784_)
  );


  anb1
  g1720
  (
    .dina(new_n1767__spl_),
    .dinb(new_n1784__spl_),
    .dout(new_n1785_)
  );


  anb2
  g1721
  (
    .dina(new_n1767__spl_),
    .dinb(new_n1784__spl_),
    .dout(new_n1786_)
  );


  anb2
  g1722
  (
    .dina(new_n1785__spl_),
    .dinb(new_n1786_),
    .dout(new_n1787_)
  );


  anb1
  g1723
  (
    .dina(new_n1766__spl_),
    .dinb(new_n1787__spl_),
    .dout(new_n1788_)
  );


  anb2
  g1724
  (
    .dina(new_n1766__spl_),
    .dinb(new_n1787__spl_),
    .dout(new_n1789_)
  );


  anb2
  g1725
  (
    .dina(new_n1788__spl_),
    .dinb(new_n1789_),
    .dout(new_n1790_)
  );


  anb1
  g1726
  (
    .dina(new_n1765__spl_),
    .dinb(new_n1790__spl_),
    .dout(new_n1791_)
  );


  anb2
  g1727
  (
    .dina(new_n1765__spl_),
    .dinb(new_n1790__spl_),
    .dout(new_n1792_)
  );


  anb2
  g1728
  (
    .dina(new_n1791__spl_),
    .dinb(new_n1792_),
    .dout(new_n1793_)
  );


  anb1
  g1729
  (
    .dina(new_n1764__spl_),
    .dinb(new_n1793__spl_),
    .dout(new_n1794_)
  );


  anb2
  g1730
  (
    .dina(new_n1764__spl_),
    .dinb(new_n1793__spl_),
    .dout(new_n1795_)
  );


  anb2
  g1731
  (
    .dina(new_n1794__spl_),
    .dinb(new_n1795_),
    .dout(new_n1796_)
  );


  anb1
  g1732
  (
    .dina(new_n1763__spl_),
    .dinb(new_n1796__spl_),
    .dout(new_n1797_)
  );


  anb2
  g1733
  (
    .dina(new_n1763__spl_),
    .dinb(new_n1796__spl_),
    .dout(new_n1798_)
  );


  anb2
  g1734
  (
    .dina(new_n1797__spl_),
    .dinb(new_n1798_),
    .dout(new_n1799_)
  );


  anb1
  g1735
  (
    .dina(new_n1762__spl_),
    .dinb(new_n1799__spl_),
    .dout(new_n1800_)
  );


  anb2
  g1736
  (
    .dina(new_n1762__spl_),
    .dinb(new_n1799__spl_),
    .dout(new_n1801_)
  );


  anb2
  g1737
  (
    .dina(new_n1800__spl_),
    .dinb(new_n1801_),
    .dout(new_n1802_)
  );


  anb1
  g1738
  (
    .dina(new_n1761__spl_),
    .dinb(new_n1802__spl_),
    .dout(new_n1803_)
  );


  anb2
  g1739
  (
    .dina(new_n1761__spl_),
    .dinb(new_n1802__spl_),
    .dout(new_n1804_)
  );


  anb2
  g1740
  (
    .dina(new_n1803__spl_),
    .dinb(new_n1804_),
    .dout(new_n1805_)
  );


  anb1
  g1741
  (
    .dina(new_n1760__spl_),
    .dinb(new_n1805__spl_),
    .dout(new_n1806_)
  );


  anb2
  g1742
  (
    .dina(new_n1760__spl_),
    .dinb(new_n1805__spl_),
    .dout(new_n1807_)
  );


  anb2
  g1743
  (
    .dina(new_n1806__spl_),
    .dinb(new_n1807_),
    .dout(G6282)
  );


  and2
  g1744
  (
    .dina(new_n1803__spl_),
    .dinb(new_n1806__spl_),
    .dout(new_n1809_)
  );


  and2
  g1745
  (
    .dina(new_n1797__spl_),
    .dinb(new_n1800__spl_),
    .dout(new_n1810_)
  );


  nor2
  g1746
  (
    .dina(G12_spl_111),
    .dinb(G32_spl_101),
    .dout(new_n1811_)
  );


  and2
  g1747
  (
    .dina(new_n1791__spl_),
    .dinb(new_n1794__spl_),
    .dout(new_n1812_)
  );


  nor2
  g1748
  (
    .dina(G13_spl_111),
    .dinb(G31_spl_110),
    .dout(new_n1813_)
  );


  and2
  g1749
  (
    .dina(new_n1785__spl_),
    .dinb(new_n1788__spl_),
    .dout(new_n1814_)
  );


  nor2
  g1750
  (
    .dina(G14_spl_110),
    .dinb(G30_spl_110),
    .dout(new_n1815_)
  );


  anb2
  g1751
  (
    .dina(new_n1779__spl_),
    .dinb(new_n1782__spl_),
    .dout(new_n1816_)
  );


  nor2
  g1752
  (
    .dina(G15_spl_110),
    .dinb(G29_spl_111),
    .dout(new_n1817_)
  );


  and1
  g1753
  (
    .dina(G16_spl_101),
    .dinb(G28_spl_111),
    .dout(new_n1818_)
  );


  anb2
  g1754
  (
    .dina(new_n1773__spl_),
    .dinb(new_n1776__spl_),
    .dout(new_n1819_)
  );


  anb2
  g1755
  (
    .dina(new_n1818__spl_),
    .dinb(new_n1819__spl_),
    .dout(new_n1820_)
  );


  anb1
  g1756
  (
    .dina(new_n1818__spl_),
    .dinb(new_n1819__spl_),
    .dout(new_n1821_)
  );


  nab2
  g1757
  (
    .dina(new_n1820__spl_),
    .dinb(new_n1821_),
    .dout(new_n1822_)
  );


  anb1
  g1758
  (
    .dina(new_n1817__spl_),
    .dinb(new_n1822__spl_),
    .dout(new_n1823_)
  );


  anb2
  g1759
  (
    .dina(new_n1817__spl_),
    .dinb(new_n1822__spl_),
    .dout(new_n1824_)
  );


  anb2
  g1760
  (
    .dina(new_n1823__spl_),
    .dinb(new_n1824_),
    .dout(new_n1825_)
  );


  anb1
  g1761
  (
    .dina(new_n1816__spl_),
    .dinb(new_n1825__spl_),
    .dout(new_n1826_)
  );


  anb2
  g1762
  (
    .dina(new_n1816__spl_),
    .dinb(new_n1825__spl_),
    .dout(new_n1827_)
  );


  anb2
  g1763
  (
    .dina(new_n1826__spl_),
    .dinb(new_n1827_),
    .dout(new_n1828_)
  );


  anb1
  g1764
  (
    .dina(new_n1815__spl_),
    .dinb(new_n1828__spl_),
    .dout(new_n1829_)
  );


  anb2
  g1765
  (
    .dina(new_n1815__spl_),
    .dinb(new_n1828__spl_),
    .dout(new_n1830_)
  );


  anb2
  g1766
  (
    .dina(new_n1829__spl_),
    .dinb(new_n1830_),
    .dout(new_n1831_)
  );


  anb1
  g1767
  (
    .dina(new_n1814__spl_),
    .dinb(new_n1831__spl_),
    .dout(new_n1832_)
  );


  anb2
  g1768
  (
    .dina(new_n1814__spl_),
    .dinb(new_n1831__spl_),
    .dout(new_n1833_)
  );


  anb2
  g1769
  (
    .dina(new_n1832__spl_),
    .dinb(new_n1833_),
    .dout(new_n1834_)
  );


  anb1
  g1770
  (
    .dina(new_n1813__spl_),
    .dinb(new_n1834__spl_),
    .dout(new_n1835_)
  );


  anb2
  g1771
  (
    .dina(new_n1813__spl_),
    .dinb(new_n1834__spl_),
    .dout(new_n1836_)
  );


  anb2
  g1772
  (
    .dina(new_n1835__spl_),
    .dinb(new_n1836_),
    .dout(new_n1837_)
  );


  anb1
  g1773
  (
    .dina(new_n1812__spl_),
    .dinb(new_n1837__spl_),
    .dout(new_n1838_)
  );


  anb2
  g1774
  (
    .dina(new_n1812__spl_),
    .dinb(new_n1837__spl_),
    .dout(new_n1839_)
  );


  anb2
  g1775
  (
    .dina(new_n1838__spl_),
    .dinb(new_n1839_),
    .dout(new_n1840_)
  );


  anb1
  g1776
  (
    .dina(new_n1811__spl_),
    .dinb(new_n1840__spl_),
    .dout(new_n1841_)
  );


  anb2
  g1777
  (
    .dina(new_n1811__spl_),
    .dinb(new_n1840__spl_),
    .dout(new_n1842_)
  );


  anb2
  g1778
  (
    .dina(new_n1841__spl_),
    .dinb(new_n1842_),
    .dout(new_n1843_)
  );


  anb1
  g1779
  (
    .dina(new_n1810__spl_),
    .dinb(new_n1843__spl_),
    .dout(new_n1844_)
  );


  anb2
  g1780
  (
    .dina(new_n1810__spl_),
    .dinb(new_n1843__spl_),
    .dout(new_n1845_)
  );


  anb2
  g1781
  (
    .dina(new_n1844__spl_),
    .dinb(new_n1845_),
    .dout(new_n1846_)
  );


  anb1
  g1782
  (
    .dina(new_n1809__spl_),
    .dinb(new_n1846__spl_),
    .dout(new_n1847_)
  );


  anb2
  g1783
  (
    .dina(new_n1809__spl_),
    .dinb(new_n1846__spl_),
    .dout(new_n1848_)
  );


  anb2
  g1784
  (
    .dina(new_n1847__spl_),
    .dinb(new_n1848_),
    .dout(G6283)
  );


  and2
  g1785
  (
    .dina(new_n1844__spl_),
    .dinb(new_n1847__spl_),
    .dout(new_n1850_)
  );


  and2
  g1786
  (
    .dina(new_n1838__spl_),
    .dinb(new_n1841__spl_),
    .dout(new_n1851_)
  );


  nor2
  g1787
  (
    .dina(G13_spl_111),
    .dinb(G32_spl_110),
    .dout(new_n1852_)
  );


  and2
  g1788
  (
    .dina(new_n1832__spl_),
    .dinb(new_n1835__spl_),
    .dout(new_n1853_)
  );


  nor2
  g1789
  (
    .dina(G14_spl_111),
    .dinb(G31_spl_110),
    .dout(new_n1854_)
  );


  and2
  g1790
  (
    .dina(new_n1826__spl_),
    .dinb(new_n1829__spl_),
    .dout(new_n1855_)
  );


  nor2
  g1791
  (
    .dina(G15_spl_110),
    .dinb(G30_spl_111),
    .dout(new_n1856_)
  );


  nor2
  g1792
  (
    .dina(G16_spl_110),
    .dinb(G29_spl_111),
    .dout(new_n1857_)
  );


  anb1
  g1793
  (
    .dina(new_n1820__spl_),
    .dinb(new_n1823__spl_),
    .dout(new_n1858_)
  );


  anb1
  g1794
  (
    .dina(new_n1857__spl_),
    .dinb(new_n1858__spl_),
    .dout(new_n1859_)
  );


  anb2
  g1795
  (
    .dina(new_n1857__spl_),
    .dinb(new_n1858__spl_),
    .dout(new_n1860_)
  );


  anb2
  g1796
  (
    .dina(new_n1859__spl_),
    .dinb(new_n1860_),
    .dout(new_n1861_)
  );


  anb1
  g1797
  (
    .dina(new_n1856__spl_),
    .dinb(new_n1861__spl_),
    .dout(new_n1862_)
  );


  anb2
  g1798
  (
    .dina(new_n1856__spl_),
    .dinb(new_n1861__spl_),
    .dout(new_n1863_)
  );


  anb2
  g1799
  (
    .dina(new_n1862__spl_),
    .dinb(new_n1863_),
    .dout(new_n1864_)
  );


  anb1
  g1800
  (
    .dina(new_n1855__spl_),
    .dinb(new_n1864__spl_),
    .dout(new_n1865_)
  );


  anb2
  g1801
  (
    .dina(new_n1855__spl_),
    .dinb(new_n1864__spl_),
    .dout(new_n1866_)
  );


  anb2
  g1802
  (
    .dina(new_n1865__spl_),
    .dinb(new_n1866_),
    .dout(new_n1867_)
  );


  anb1
  g1803
  (
    .dina(new_n1854__spl_),
    .dinb(new_n1867__spl_),
    .dout(new_n1868_)
  );


  anb2
  g1804
  (
    .dina(new_n1854__spl_),
    .dinb(new_n1867__spl_),
    .dout(new_n1869_)
  );


  anb2
  g1805
  (
    .dina(new_n1868__spl_),
    .dinb(new_n1869_),
    .dout(new_n1870_)
  );


  anb1
  g1806
  (
    .dina(new_n1853__spl_),
    .dinb(new_n1870__spl_),
    .dout(new_n1871_)
  );


  anb2
  g1807
  (
    .dina(new_n1853__spl_),
    .dinb(new_n1870__spl_),
    .dout(new_n1872_)
  );


  anb2
  g1808
  (
    .dina(new_n1871__spl_),
    .dinb(new_n1872_),
    .dout(new_n1873_)
  );


  anb1
  g1809
  (
    .dina(new_n1852__spl_),
    .dinb(new_n1873__spl_),
    .dout(new_n1874_)
  );


  anb2
  g1810
  (
    .dina(new_n1852__spl_),
    .dinb(new_n1873__spl_),
    .dout(new_n1875_)
  );


  anb2
  g1811
  (
    .dina(new_n1874__spl_),
    .dinb(new_n1875_),
    .dout(new_n1876_)
  );


  anb1
  g1812
  (
    .dina(new_n1851__spl_),
    .dinb(new_n1876__spl_),
    .dout(new_n1877_)
  );


  anb2
  g1813
  (
    .dina(new_n1851__spl_),
    .dinb(new_n1876__spl_),
    .dout(new_n1878_)
  );


  anb2
  g1814
  (
    .dina(new_n1877__spl_),
    .dinb(new_n1878_),
    .dout(new_n1879_)
  );


  anb1
  g1815
  (
    .dina(new_n1850__spl_),
    .dinb(new_n1879__spl_),
    .dout(new_n1880_)
  );


  anb2
  g1816
  (
    .dina(new_n1850__spl_),
    .dinb(new_n1879__spl_),
    .dout(new_n1881_)
  );


  anb2
  g1817
  (
    .dina(new_n1880__spl_),
    .dinb(new_n1881_),
    .dout(G6284)
  );


  and2
  g1818
  (
    .dina(new_n1877__spl_),
    .dinb(new_n1880__spl_),
    .dout(new_n1883_)
  );


  and2
  g1819
  (
    .dina(new_n1871__spl_),
    .dinb(new_n1874__spl_),
    .dout(new_n1884_)
  );


  nor2
  g1820
  (
    .dina(G14_spl_111),
    .dinb(G32_spl_110),
    .dout(new_n1885_)
  );


  and2
  g1821
  (
    .dina(new_n1865__spl_),
    .dinb(new_n1868__spl_),
    .dout(new_n1886_)
  );


  nor2
  g1822
  (
    .dina(G15_spl_111),
    .dinb(G31_spl_111),
    .dout(new_n1887_)
  );


  nor2
  g1823
  (
    .dina(G16_spl_110),
    .dinb(G30_spl_111),
    .dout(new_n1888_)
  );


  nor1
  g1824
  (
    .dina(new_n1859__spl_),
    .dinb(new_n1862__spl_),
    .dout(new_n1889_)
  );


  anb1
  g1825
  (
    .dina(new_n1888__spl_),
    .dinb(new_n1889__spl_),
    .dout(new_n1890_)
  );


  anb2
  g1826
  (
    .dina(new_n1888__spl_),
    .dinb(new_n1889__spl_),
    .dout(new_n1891_)
  );


  anb2
  g1827
  (
    .dina(new_n1890__spl_),
    .dinb(new_n1891_),
    .dout(new_n1892_)
  );


  anb1
  g1828
  (
    .dina(new_n1887__spl_),
    .dinb(new_n1892__spl_),
    .dout(new_n1893_)
  );


  anb2
  g1829
  (
    .dina(new_n1887__spl_),
    .dinb(new_n1892__spl_),
    .dout(new_n1894_)
  );


  anb2
  g1830
  (
    .dina(new_n1893__spl_),
    .dinb(new_n1894_),
    .dout(new_n1895_)
  );


  anb1
  g1831
  (
    .dina(new_n1886__spl_),
    .dinb(new_n1895__spl_),
    .dout(new_n1896_)
  );


  anb2
  g1832
  (
    .dina(new_n1886__spl_),
    .dinb(new_n1895__spl_),
    .dout(new_n1897_)
  );


  anb2
  g1833
  (
    .dina(new_n1896__spl_),
    .dinb(new_n1897_),
    .dout(new_n1898_)
  );


  anb1
  g1834
  (
    .dina(new_n1885__spl_),
    .dinb(new_n1898__spl_),
    .dout(new_n1899_)
  );


  anb2
  g1835
  (
    .dina(new_n1885__spl_),
    .dinb(new_n1898__spl_),
    .dout(new_n1900_)
  );


  anb2
  g1836
  (
    .dina(new_n1899__spl_),
    .dinb(new_n1900_),
    .dout(new_n1901_)
  );


  anb1
  g1837
  (
    .dina(new_n1884__spl_),
    .dinb(new_n1901__spl_),
    .dout(new_n1902_)
  );


  anb2
  g1838
  (
    .dina(new_n1884__spl_),
    .dinb(new_n1901__spl_),
    .dout(new_n1903_)
  );


  anb2
  g1839
  (
    .dina(new_n1902__spl_),
    .dinb(new_n1903_),
    .dout(new_n1904_)
  );


  anb1
  g1840
  (
    .dina(new_n1883__spl_),
    .dinb(new_n1904__spl_),
    .dout(new_n1905_)
  );


  anb2
  g1841
  (
    .dina(new_n1883__spl_),
    .dinb(new_n1904__spl_),
    .dout(new_n1906_)
  );


  anb2
  g1842
  (
    .dina(new_n1905__spl_),
    .dinb(new_n1906_),
    .dout(G6285)
  );


  and2
  g1843
  (
    .dina(new_n1902__spl_),
    .dinb(new_n1905__spl_),
    .dout(new_n1908_)
  );


  and2
  g1844
  (
    .dina(new_n1896__spl_),
    .dinb(new_n1899__spl_),
    .dout(new_n1909_)
  );


  nor2
  g1845
  (
    .dina(G15_spl_111),
    .dinb(G32_spl_111),
    .dout(new_n1910_)
  );


  nor2
  g1846
  (
    .dina(G16_spl_111),
    .dinb(G31_spl_111),
    .dout(new_n1911_)
  );


  nor1
  g1847
  (
    .dina(new_n1890__spl_),
    .dinb(new_n1893__spl_),
    .dout(new_n1912_)
  );


  anb1
  g1848
  (
    .dina(new_n1911__spl_),
    .dinb(new_n1912__spl_),
    .dout(new_n1913_)
  );


  anb2
  g1849
  (
    .dina(new_n1911__spl_),
    .dinb(new_n1912__spl_),
    .dout(new_n1914_)
  );


  anb2
  g1850
  (
    .dina(new_n1913__spl_),
    .dinb(new_n1914_),
    .dout(new_n1915_)
  );


  anb1
  g1851
  (
    .dina(new_n1910__spl_),
    .dinb(new_n1915__spl_),
    .dout(new_n1916_)
  );


  anb2
  g1852
  (
    .dina(new_n1910__spl_),
    .dinb(new_n1915__spl_),
    .dout(new_n1917_)
  );


  anb2
  g1853
  (
    .dina(new_n1916__spl_),
    .dinb(new_n1917_),
    .dout(new_n1918_)
  );


  anb1
  g1854
  (
    .dina(new_n1909__spl_),
    .dinb(new_n1918__spl_),
    .dout(new_n1919_)
  );


  anb2
  g1855
  (
    .dina(new_n1909__spl_),
    .dinb(new_n1918__spl_),
    .dout(new_n1920_)
  );


  anb2
  g1856
  (
    .dina(new_n1919__spl_),
    .dinb(new_n1920_),
    .dout(new_n1921_)
  );


  anb1
  g1857
  (
    .dina(new_n1908__spl_),
    .dinb(new_n1921__spl_),
    .dout(new_n1922_)
  );


  anb2
  g1858
  (
    .dina(new_n1908__spl_),
    .dinb(new_n1921__spl_),
    .dout(new_n1923_)
  );


  anb2
  g1859
  (
    .dina(new_n1922__spl_),
    .dinb(new_n1923_),
    .dout(G6286)
  );


  nor2
  g1860
  (
    .dina(G16_spl_111),
    .dinb(G32_spl_111),
    .dout(new_n1925_)
  );


  nor1
  g1861
  (
    .dina(new_n1913__spl_),
    .dinb(new_n1916__spl_),
    .dout(new_n1926_)
  );


  anb1
  g1862
  (
    .dina(new_n1925__spl_),
    .dinb(new_n1926__spl_),
    .dout(new_n1927_)
  );


  and2
  g1863
  (
    .dina(new_n1919__spl_),
    .dinb(new_n1922__spl_),
    .dout(new_n1928_)
  );


  anb2
  g1864
  (
    .dina(new_n1925__spl_),
    .dinb(new_n1926__spl_),
    .dout(new_n1929_)
  );


  anb2
  g1865
  (
    .dina(new_n1927__spl_),
    .dinb(new_n1929_),
    .dout(new_n1930_)
  );


  anb1
  g1866
  (
    .dina(new_n1928__spl_),
    .dinb(new_n1930__spl_),
    .dout(new_n1931_)
  );


  nor1
  g1867
  (
    .dina(new_n1927__spl_),
    .dinb(new_n1931__spl_),
    .dout(G6287)
  );


  anb2
  g1868
  (
    .dina(new_n1928__spl_),
    .dinb(new_n1930__spl_),
    .dout(new_n1933_)
  );


  anb2
  g1869
  (
    .dina(new_n1931__spl_),
    .dinb(new_n1933_),
    .dout(G6288)
  );


  splt
  gG1
  (
    .dout(G1_spl_),
    .din(G1)
  );


  splt
  gG1_spl_
  (
    .dout(G1_spl_0),
    .din(G1_spl_)
  );


  splt
  gG1_spl_0
  (
    .dout(G1_spl_00),
    .din(G1_spl_0)
  );


  splt
  gG1_spl_00
  (
    .dout(G1_spl_000),
    .din(G1_spl_00)
  );


  splt
  gG1_spl_00
  (
    .dout(G1_spl_001),
    .din(G1_spl_00)
  );


  splt
  gG1_spl_0
  (
    .dout(G1_spl_01),
    .din(G1_spl_0)
  );


  splt
  gG1_spl_01
  (
    .dout(G1_spl_010),
    .din(G1_spl_01)
  );


  splt
  gG1_spl_01
  (
    .dout(G1_spl_011),
    .din(G1_spl_01)
  );


  splt
  gG1_spl_
  (
    .dout(G1_spl_1),
    .din(G1_spl_)
  );


  splt
  gG1_spl_1
  (
    .dout(G1_spl_10),
    .din(G1_spl_1)
  );


  splt
  gG1_spl_10
  (
    .dout(G1_spl_100),
    .din(G1_spl_10)
  );


  splt
  gG1_spl_10
  (
    .dout(G1_spl_101),
    .din(G1_spl_10)
  );


  splt
  gG1_spl_1
  (
    .dout(G1_spl_11),
    .din(G1_spl_1)
  );


  splt
  gG1_spl_11
  (
    .dout(G1_spl_110),
    .din(G1_spl_11)
  );


  splt
  gG1_spl_11
  (
    .dout(G1_spl_111),
    .din(G1_spl_11)
  );


  splt
  gG17
  (
    .dout(G17_spl_),
    .din(G17)
  );


  splt
  gG17_spl_
  (
    .dout(G17_spl_0),
    .din(G17_spl_)
  );


  splt
  gG17_spl_0
  (
    .dout(G17_spl_00),
    .din(G17_spl_0)
  );


  splt
  gG17_spl_00
  (
    .dout(G17_spl_000),
    .din(G17_spl_00)
  );


  splt
  gG17_spl_00
  (
    .dout(G17_spl_001),
    .din(G17_spl_00)
  );


  splt
  gG17_spl_0
  (
    .dout(G17_spl_01),
    .din(G17_spl_0)
  );


  splt
  gG17_spl_01
  (
    .dout(G17_spl_010),
    .din(G17_spl_01)
  );


  splt
  gG17_spl_01
  (
    .dout(G17_spl_011),
    .din(G17_spl_01)
  );


  splt
  gG17_spl_
  (
    .dout(G17_spl_1),
    .din(G17_spl_)
  );


  splt
  gG17_spl_1
  (
    .dout(G17_spl_10),
    .din(G17_spl_1)
  );


  splt
  gG17_spl_10
  (
    .dout(G17_spl_100),
    .din(G17_spl_10)
  );


  splt
  gG17_spl_10
  (
    .dout(G17_spl_101),
    .din(G17_spl_10)
  );


  splt
  gG17_spl_1
  (
    .dout(G17_spl_11),
    .din(G17_spl_1)
  );


  splt
  gG17_spl_11
  (
    .dout(G17_spl_110),
    .din(G17_spl_11)
  );


  splt
  gG17_spl_11
  (
    .dout(G17_spl_111),
    .din(G17_spl_11)
  );


  splt
  gG2
  (
    .dout(G2_spl_),
    .din(G2)
  );


  splt
  gG2_spl_
  (
    .dout(G2_spl_0),
    .din(G2_spl_)
  );


  splt
  gG2_spl_0
  (
    .dout(G2_spl_00),
    .din(G2_spl_0)
  );


  splt
  gG2_spl_00
  (
    .dout(G2_spl_000),
    .din(G2_spl_00)
  );


  splt
  gG2_spl_00
  (
    .dout(G2_spl_001),
    .din(G2_spl_00)
  );


  splt
  gG2_spl_0
  (
    .dout(G2_spl_01),
    .din(G2_spl_0)
  );


  splt
  gG2_spl_01
  (
    .dout(G2_spl_010),
    .din(G2_spl_01)
  );


  splt
  gG2_spl_01
  (
    .dout(G2_spl_011),
    .din(G2_spl_01)
  );


  splt
  gG2_spl_
  (
    .dout(G2_spl_1),
    .din(G2_spl_)
  );


  splt
  gG2_spl_1
  (
    .dout(G2_spl_10),
    .din(G2_spl_1)
  );


  splt
  gG2_spl_10
  (
    .dout(G2_spl_100),
    .din(G2_spl_10)
  );


  splt
  gG2_spl_10
  (
    .dout(G2_spl_101),
    .din(G2_spl_10)
  );


  splt
  gG2_spl_1
  (
    .dout(G2_spl_11),
    .din(G2_spl_1)
  );


  splt
  gG2_spl_11
  (
    .dout(G2_spl_110),
    .din(G2_spl_11)
  );


  splt
  gG2_spl_11
  (
    .dout(G2_spl_111),
    .din(G2_spl_11)
  );


  splt
  gG18
  (
    .dout(G18_spl_),
    .din(G18)
  );


  splt
  gG18_spl_
  (
    .dout(G18_spl_0),
    .din(G18_spl_)
  );


  splt
  gG18_spl_0
  (
    .dout(G18_spl_00),
    .din(G18_spl_0)
  );


  splt
  gG18_spl_00
  (
    .dout(G18_spl_000),
    .din(G18_spl_00)
  );


  splt
  gG18_spl_00
  (
    .dout(G18_spl_001),
    .din(G18_spl_00)
  );


  splt
  gG18_spl_0
  (
    .dout(G18_spl_01),
    .din(G18_spl_0)
  );


  splt
  gG18_spl_01
  (
    .dout(G18_spl_010),
    .din(G18_spl_01)
  );


  splt
  gG18_spl_01
  (
    .dout(G18_spl_011),
    .din(G18_spl_01)
  );


  splt
  gG18_spl_
  (
    .dout(G18_spl_1),
    .din(G18_spl_)
  );


  splt
  gG18_spl_1
  (
    .dout(G18_spl_10),
    .din(G18_spl_1)
  );


  splt
  gG18_spl_10
  (
    .dout(G18_spl_100),
    .din(G18_spl_10)
  );


  splt
  gG18_spl_10
  (
    .dout(G18_spl_101),
    .din(G18_spl_10)
  );


  splt
  gG18_spl_1
  (
    .dout(G18_spl_11),
    .din(G18_spl_1)
  );


  splt
  gG18_spl_11
  (
    .dout(G18_spl_110),
    .din(G18_spl_11)
  );


  splt
  gG18_spl_11
  (
    .dout(G18_spl_111),
    .din(G18_spl_11)
  );


  splt
  gnew_n66_
  (
    .dout(new_n66__spl_),
    .din(new_n66_)
  );


  splt
  gnew_n67_
  (
    .dout(new_n67__spl_),
    .din(new_n67_)
  );


  splt
  gnew_n68_
  (
    .dout(new_n68__spl_),
    .din(new_n68_)
  );


  splt
  gnew_n68__spl_
  (
    .dout(new_n68__spl_0),
    .din(new_n68__spl_)
  );


  splt
  gG19
  (
    .dout(G19_spl_),
    .din(G19)
  );


  splt
  gG19_spl_
  (
    .dout(G19_spl_0),
    .din(G19_spl_)
  );


  splt
  gG19_spl_0
  (
    .dout(G19_spl_00),
    .din(G19_spl_0)
  );


  splt
  gG19_spl_00
  (
    .dout(G19_spl_000),
    .din(G19_spl_00)
  );


  splt
  gG19_spl_00
  (
    .dout(G19_spl_001),
    .din(G19_spl_00)
  );


  splt
  gG19_spl_0
  (
    .dout(G19_spl_01),
    .din(G19_spl_0)
  );


  splt
  gG19_spl_01
  (
    .dout(G19_spl_010),
    .din(G19_spl_01)
  );


  splt
  gG19_spl_01
  (
    .dout(G19_spl_011),
    .din(G19_spl_01)
  );


  splt
  gG19_spl_
  (
    .dout(G19_spl_1),
    .din(G19_spl_)
  );


  splt
  gG19_spl_1
  (
    .dout(G19_spl_10),
    .din(G19_spl_1)
  );


  splt
  gG19_spl_10
  (
    .dout(G19_spl_100),
    .din(G19_spl_10)
  );


  splt
  gG19_spl_10
  (
    .dout(G19_spl_101),
    .din(G19_spl_10)
  );


  splt
  gG19_spl_1
  (
    .dout(G19_spl_11),
    .din(G19_spl_1)
  );


  splt
  gG19_spl_11
  (
    .dout(G19_spl_110),
    .din(G19_spl_11)
  );


  splt
  gG19_spl_11
  (
    .dout(G19_spl_111),
    .din(G19_spl_11)
  );


  splt
  gG3
  (
    .dout(G3_spl_),
    .din(G3)
  );


  splt
  gG3_spl_
  (
    .dout(G3_spl_0),
    .din(G3_spl_)
  );


  splt
  gG3_spl_0
  (
    .dout(G3_spl_00),
    .din(G3_spl_0)
  );


  splt
  gG3_spl_00
  (
    .dout(G3_spl_000),
    .din(G3_spl_00)
  );


  splt
  gG3_spl_00
  (
    .dout(G3_spl_001),
    .din(G3_spl_00)
  );


  splt
  gG3_spl_0
  (
    .dout(G3_spl_01),
    .din(G3_spl_0)
  );


  splt
  gG3_spl_01
  (
    .dout(G3_spl_010),
    .din(G3_spl_01)
  );


  splt
  gG3_spl_01
  (
    .dout(G3_spl_011),
    .din(G3_spl_01)
  );


  splt
  gG3_spl_
  (
    .dout(G3_spl_1),
    .din(G3_spl_)
  );


  splt
  gG3_spl_1
  (
    .dout(G3_spl_10),
    .din(G3_spl_1)
  );


  splt
  gG3_spl_10
  (
    .dout(G3_spl_100),
    .din(G3_spl_10)
  );


  splt
  gG3_spl_10
  (
    .dout(G3_spl_101),
    .din(G3_spl_10)
  );


  splt
  gG3_spl_1
  (
    .dout(G3_spl_11),
    .din(G3_spl_1)
  );


  splt
  gG3_spl_11
  (
    .dout(G3_spl_110),
    .din(G3_spl_11)
  );


  splt
  gG3_spl_11
  (
    .dout(G3_spl_111),
    .din(G3_spl_11)
  );


  splt
  gnew_n72_
  (
    .dout(new_n72__spl_),
    .din(new_n72_)
  );


  splt
  gnew_n73_
  (
    .dout(new_n73__spl_),
    .din(new_n73_)
  );


  splt
  gnew_n74_
  (
    .dout(new_n74__spl_),
    .din(new_n74_)
  );


  splt
  gnew_n74__spl_
  (
    .dout(new_n74__spl_0),
    .din(new_n74__spl_)
  );


  splt
  gnew_n76_
  (
    .dout(new_n76__spl_),
    .din(new_n76_)
  );


  splt
  gnew_n77_
  (
    .dout(new_n77__spl_),
    .din(new_n77_)
  );


  splt
  gnew_n71_
  (
    .dout(new_n71__spl_),
    .din(new_n71_)
  );


  splt
  gnew_n79_
  (
    .dout(new_n79__spl_),
    .din(new_n79_)
  );


  splt
  gnew_n80_
  (
    .dout(new_n80__spl_),
    .din(new_n80_)
  );


  splt
  gG20
  (
    .dout(G20_spl_),
    .din(G20)
  );


  splt
  gG20_spl_
  (
    .dout(G20_spl_0),
    .din(G20_spl_)
  );


  splt
  gG20_spl_0
  (
    .dout(G20_spl_00),
    .din(G20_spl_0)
  );


  splt
  gG20_spl_00
  (
    .dout(G20_spl_000),
    .din(G20_spl_00)
  );


  splt
  gG20_spl_00
  (
    .dout(G20_spl_001),
    .din(G20_spl_00)
  );


  splt
  gG20_spl_0
  (
    .dout(G20_spl_01),
    .din(G20_spl_0)
  );


  splt
  gG20_spl_01
  (
    .dout(G20_spl_010),
    .din(G20_spl_01)
  );


  splt
  gG20_spl_01
  (
    .dout(G20_spl_011),
    .din(G20_spl_01)
  );


  splt
  gG20_spl_
  (
    .dout(G20_spl_1),
    .din(G20_spl_)
  );


  splt
  gG20_spl_1
  (
    .dout(G20_spl_10),
    .din(G20_spl_1)
  );


  splt
  gG20_spl_10
  (
    .dout(G20_spl_100),
    .din(G20_spl_10)
  );


  splt
  gG20_spl_10
  (
    .dout(G20_spl_101),
    .din(G20_spl_10)
  );


  splt
  gG20_spl_1
  (
    .dout(G20_spl_11),
    .din(G20_spl_1)
  );


  splt
  gG20_spl_11
  (
    .dout(G20_spl_110),
    .din(G20_spl_11)
  );


  splt
  gG20_spl_11
  (
    .dout(G20_spl_111),
    .din(G20_spl_11)
  );


  splt
  gG4
  (
    .dout(G4_spl_),
    .din(G4)
  );


  splt
  gG4_spl_
  (
    .dout(G4_spl_0),
    .din(G4_spl_)
  );


  splt
  gG4_spl_0
  (
    .dout(G4_spl_00),
    .din(G4_spl_0)
  );


  splt
  gG4_spl_00
  (
    .dout(G4_spl_000),
    .din(G4_spl_00)
  );


  splt
  gG4_spl_00
  (
    .dout(G4_spl_001),
    .din(G4_spl_00)
  );


  splt
  gG4_spl_0
  (
    .dout(G4_spl_01),
    .din(G4_spl_0)
  );


  splt
  gG4_spl_01
  (
    .dout(G4_spl_010),
    .din(G4_spl_01)
  );


  splt
  gG4_spl_01
  (
    .dout(G4_spl_011),
    .din(G4_spl_01)
  );


  splt
  gG4_spl_
  (
    .dout(G4_spl_1),
    .din(G4_spl_)
  );


  splt
  gG4_spl_1
  (
    .dout(G4_spl_10),
    .din(G4_spl_1)
  );


  splt
  gG4_spl_10
  (
    .dout(G4_spl_100),
    .din(G4_spl_10)
  );


  splt
  gG4_spl_10
  (
    .dout(G4_spl_101),
    .din(G4_spl_10)
  );


  splt
  gG4_spl_1
  (
    .dout(G4_spl_11),
    .din(G4_spl_1)
  );


  splt
  gG4_spl_11
  (
    .dout(G4_spl_110),
    .din(G4_spl_11)
  );


  splt
  gG4_spl_11
  (
    .dout(G4_spl_111),
    .din(G4_spl_11)
  );


  splt
  gnew_n86_
  (
    .dout(new_n86__spl_),
    .din(new_n86_)
  );


  splt
  gnew_n87_
  (
    .dout(new_n87__spl_),
    .din(new_n87_)
  );


  splt
  gnew_n88_
  (
    .dout(new_n88__spl_),
    .din(new_n88_)
  );


  splt
  gnew_n88__spl_
  (
    .dout(new_n88__spl_0),
    .din(new_n88__spl_)
  );


  splt
  gnew_n90_
  (
    .dout(new_n90__spl_),
    .din(new_n90_)
  );


  splt
  gnew_n91_
  (
    .dout(new_n91__spl_),
    .din(new_n91_)
  );


  splt
  gnew_n85_
  (
    .dout(new_n85__spl_),
    .din(new_n85_)
  );


  splt
  gnew_n93_
  (
    .dout(new_n93__spl_),
    .din(new_n93_)
  );


  splt
  gnew_n94_
  (
    .dout(new_n94__spl_),
    .din(new_n94_)
  );


  splt
  gnew_n84_
  (
    .dout(new_n84__spl_),
    .din(new_n84_)
  );


  splt
  gnew_n96_
  (
    .dout(new_n96__spl_),
    .din(new_n96_)
  );


  splt
  gnew_n97_
  (
    .dout(new_n97__spl_),
    .din(new_n97_)
  );


  splt
  gnew_n83_
  (
    .dout(new_n83__spl_),
    .din(new_n83_)
  );


  splt
  gnew_n99_
  (
    .dout(new_n99__spl_),
    .din(new_n99_)
  );


  splt
  gnew_n100_
  (
    .dout(new_n100__spl_),
    .din(new_n100_)
  );


  splt
  gG21
  (
    .dout(G21_spl_),
    .din(G21)
  );


  splt
  gG21_spl_
  (
    .dout(G21_spl_0),
    .din(G21_spl_)
  );


  splt
  gG21_spl_0
  (
    .dout(G21_spl_00),
    .din(G21_spl_0)
  );


  splt
  gG21_spl_00
  (
    .dout(G21_spl_000),
    .din(G21_spl_00)
  );


  splt
  gG21_spl_00
  (
    .dout(G21_spl_001),
    .din(G21_spl_00)
  );


  splt
  gG21_spl_0
  (
    .dout(G21_spl_01),
    .din(G21_spl_0)
  );


  splt
  gG21_spl_01
  (
    .dout(G21_spl_010),
    .din(G21_spl_01)
  );


  splt
  gG21_spl_01
  (
    .dout(G21_spl_011),
    .din(G21_spl_01)
  );


  splt
  gG21_spl_
  (
    .dout(G21_spl_1),
    .din(G21_spl_)
  );


  splt
  gG21_spl_1
  (
    .dout(G21_spl_10),
    .din(G21_spl_1)
  );


  splt
  gG21_spl_10
  (
    .dout(G21_spl_100),
    .din(G21_spl_10)
  );


  splt
  gG21_spl_10
  (
    .dout(G21_spl_101),
    .din(G21_spl_10)
  );


  splt
  gG21_spl_1
  (
    .dout(G21_spl_11),
    .din(G21_spl_1)
  );


  splt
  gG21_spl_11
  (
    .dout(G21_spl_110),
    .din(G21_spl_11)
  );


  splt
  gG21_spl_11
  (
    .dout(G21_spl_111),
    .din(G21_spl_11)
  );


  splt
  gG5
  (
    .dout(G5_spl_),
    .din(G5)
  );


  splt
  gG5_spl_
  (
    .dout(G5_spl_0),
    .din(G5_spl_)
  );


  splt
  gG5_spl_0
  (
    .dout(G5_spl_00),
    .din(G5_spl_0)
  );


  splt
  gG5_spl_00
  (
    .dout(G5_spl_000),
    .din(G5_spl_00)
  );


  splt
  gG5_spl_00
  (
    .dout(G5_spl_001),
    .din(G5_spl_00)
  );


  splt
  gG5_spl_0
  (
    .dout(G5_spl_01),
    .din(G5_spl_0)
  );


  splt
  gG5_spl_01
  (
    .dout(G5_spl_010),
    .din(G5_spl_01)
  );


  splt
  gG5_spl_01
  (
    .dout(G5_spl_011),
    .din(G5_spl_01)
  );


  splt
  gG5_spl_
  (
    .dout(G5_spl_1),
    .din(G5_spl_)
  );


  splt
  gG5_spl_1
  (
    .dout(G5_spl_10),
    .din(G5_spl_1)
  );


  splt
  gG5_spl_10
  (
    .dout(G5_spl_100),
    .din(G5_spl_10)
  );


  splt
  gG5_spl_10
  (
    .dout(G5_spl_101),
    .din(G5_spl_10)
  );


  splt
  gG5_spl_1
  (
    .dout(G5_spl_11),
    .din(G5_spl_1)
  );


  splt
  gG5_spl_11
  (
    .dout(G5_spl_110),
    .din(G5_spl_11)
  );


  splt
  gG5_spl_11
  (
    .dout(G5_spl_111),
    .din(G5_spl_11)
  );


  splt
  gnew_n108_
  (
    .dout(new_n108__spl_),
    .din(new_n108_)
  );


  splt
  gnew_n109_
  (
    .dout(new_n109__spl_),
    .din(new_n109_)
  );


  splt
  gnew_n110_
  (
    .dout(new_n110__spl_),
    .din(new_n110_)
  );


  splt
  gnew_n110__spl_
  (
    .dout(new_n110__spl_0),
    .din(new_n110__spl_)
  );


  splt
  gnew_n112_
  (
    .dout(new_n112__spl_),
    .din(new_n112_)
  );


  splt
  gnew_n113_
  (
    .dout(new_n113__spl_),
    .din(new_n113_)
  );


  splt
  gnew_n107_
  (
    .dout(new_n107__spl_),
    .din(new_n107_)
  );


  splt
  gnew_n115_
  (
    .dout(new_n115__spl_),
    .din(new_n115_)
  );


  splt
  gnew_n116_
  (
    .dout(new_n116__spl_),
    .din(new_n116_)
  );


  splt
  gnew_n106_
  (
    .dout(new_n106__spl_),
    .din(new_n106_)
  );


  splt
  gnew_n118_
  (
    .dout(new_n118__spl_),
    .din(new_n118_)
  );


  splt
  gnew_n119_
  (
    .dout(new_n119__spl_),
    .din(new_n119_)
  );


  splt
  gnew_n105_
  (
    .dout(new_n105__spl_),
    .din(new_n105_)
  );


  splt
  gnew_n121_
  (
    .dout(new_n121__spl_),
    .din(new_n121_)
  );


  splt
  gnew_n122_
  (
    .dout(new_n122__spl_),
    .din(new_n122_)
  );


  splt
  gnew_n104_
  (
    .dout(new_n104__spl_),
    .din(new_n104_)
  );


  splt
  gnew_n124_
  (
    .dout(new_n124__spl_),
    .din(new_n124_)
  );


  splt
  gnew_n125_
  (
    .dout(new_n125__spl_),
    .din(new_n125_)
  );


  splt
  gnew_n103_
  (
    .dout(new_n103__spl_),
    .din(new_n103_)
  );


  splt
  gnew_n127_
  (
    .dout(new_n127__spl_),
    .din(new_n127_)
  );


  splt
  gnew_n128_
  (
    .dout(new_n128__spl_),
    .din(new_n128_)
  );


  splt
  gG22
  (
    .dout(G22_spl_),
    .din(G22)
  );


  splt
  gG22_spl_
  (
    .dout(G22_spl_0),
    .din(G22_spl_)
  );


  splt
  gG22_spl_0
  (
    .dout(G22_spl_00),
    .din(G22_spl_0)
  );


  splt
  gG22_spl_00
  (
    .dout(G22_spl_000),
    .din(G22_spl_00)
  );


  splt
  gG22_spl_00
  (
    .dout(G22_spl_001),
    .din(G22_spl_00)
  );


  splt
  gG22_spl_0
  (
    .dout(G22_spl_01),
    .din(G22_spl_0)
  );


  splt
  gG22_spl_01
  (
    .dout(G22_spl_010),
    .din(G22_spl_01)
  );


  splt
  gG22_spl_01
  (
    .dout(G22_spl_011),
    .din(G22_spl_01)
  );


  splt
  gG22_spl_
  (
    .dout(G22_spl_1),
    .din(G22_spl_)
  );


  splt
  gG22_spl_1
  (
    .dout(G22_spl_10),
    .din(G22_spl_1)
  );


  splt
  gG22_spl_10
  (
    .dout(G22_spl_100),
    .din(G22_spl_10)
  );


  splt
  gG22_spl_10
  (
    .dout(G22_spl_101),
    .din(G22_spl_10)
  );


  splt
  gG22_spl_1
  (
    .dout(G22_spl_11),
    .din(G22_spl_1)
  );


  splt
  gG22_spl_11
  (
    .dout(G22_spl_110),
    .din(G22_spl_11)
  );


  splt
  gG22_spl_11
  (
    .dout(G22_spl_111),
    .din(G22_spl_11)
  );


  splt
  gG6
  (
    .dout(G6_spl_),
    .din(G6)
  );


  splt
  gG6_spl_
  (
    .dout(G6_spl_0),
    .din(G6_spl_)
  );


  splt
  gG6_spl_0
  (
    .dout(G6_spl_00),
    .din(G6_spl_0)
  );


  splt
  gG6_spl_00
  (
    .dout(G6_spl_000),
    .din(G6_spl_00)
  );


  splt
  gG6_spl_00
  (
    .dout(G6_spl_001),
    .din(G6_spl_00)
  );


  splt
  gG6_spl_0
  (
    .dout(G6_spl_01),
    .din(G6_spl_0)
  );


  splt
  gG6_spl_01
  (
    .dout(G6_spl_010),
    .din(G6_spl_01)
  );


  splt
  gG6_spl_01
  (
    .dout(G6_spl_011),
    .din(G6_spl_01)
  );


  splt
  gG6_spl_
  (
    .dout(G6_spl_1),
    .din(G6_spl_)
  );


  splt
  gG6_spl_1
  (
    .dout(G6_spl_10),
    .din(G6_spl_1)
  );


  splt
  gG6_spl_10
  (
    .dout(G6_spl_100),
    .din(G6_spl_10)
  );


  splt
  gG6_spl_10
  (
    .dout(G6_spl_101),
    .din(G6_spl_10)
  );


  splt
  gG6_spl_1
  (
    .dout(G6_spl_11),
    .din(G6_spl_1)
  );


  splt
  gG6_spl_11
  (
    .dout(G6_spl_110),
    .din(G6_spl_11)
  );


  splt
  gG6_spl_11
  (
    .dout(G6_spl_111),
    .din(G6_spl_11)
  );


  splt
  gnew_n138_
  (
    .dout(new_n138__spl_),
    .din(new_n138_)
  );


  splt
  gnew_n139_
  (
    .dout(new_n139__spl_),
    .din(new_n139_)
  );


  splt
  gnew_n140_
  (
    .dout(new_n140__spl_),
    .din(new_n140_)
  );


  splt
  gnew_n140__spl_
  (
    .dout(new_n140__spl_0),
    .din(new_n140__spl_)
  );


  splt
  gnew_n142_
  (
    .dout(new_n142__spl_),
    .din(new_n142_)
  );


  splt
  gnew_n143_
  (
    .dout(new_n143__spl_),
    .din(new_n143_)
  );


  splt
  gnew_n137_
  (
    .dout(new_n137__spl_),
    .din(new_n137_)
  );


  splt
  gnew_n145_
  (
    .dout(new_n145__spl_),
    .din(new_n145_)
  );


  splt
  gnew_n146_
  (
    .dout(new_n146__spl_),
    .din(new_n146_)
  );


  splt
  gnew_n136_
  (
    .dout(new_n136__spl_),
    .din(new_n136_)
  );


  splt
  gnew_n148_
  (
    .dout(new_n148__spl_),
    .din(new_n148_)
  );


  splt
  gnew_n149_
  (
    .dout(new_n149__spl_),
    .din(new_n149_)
  );


  splt
  gnew_n135_
  (
    .dout(new_n135__spl_),
    .din(new_n135_)
  );


  splt
  gnew_n151_
  (
    .dout(new_n151__spl_),
    .din(new_n151_)
  );


  splt
  gnew_n152_
  (
    .dout(new_n152__spl_),
    .din(new_n152_)
  );


  splt
  gnew_n134_
  (
    .dout(new_n134__spl_),
    .din(new_n134_)
  );


  splt
  gnew_n154_
  (
    .dout(new_n154__spl_),
    .din(new_n154_)
  );


  splt
  gnew_n155_
  (
    .dout(new_n155__spl_),
    .din(new_n155_)
  );


  splt
  gnew_n133_
  (
    .dout(new_n133__spl_),
    .din(new_n133_)
  );


  splt
  gnew_n157_
  (
    .dout(new_n157__spl_),
    .din(new_n157_)
  );


  splt
  gnew_n158_
  (
    .dout(new_n158__spl_),
    .din(new_n158_)
  );


  splt
  gnew_n132_
  (
    .dout(new_n132__spl_),
    .din(new_n132_)
  );


  splt
  gnew_n160_
  (
    .dout(new_n160__spl_),
    .din(new_n160_)
  );


  splt
  gnew_n161_
  (
    .dout(new_n161__spl_),
    .din(new_n161_)
  );


  splt
  gnew_n131_
  (
    .dout(new_n131__spl_),
    .din(new_n131_)
  );


  splt
  gnew_n163_
  (
    .dout(new_n163__spl_),
    .din(new_n163_)
  );


  splt
  gnew_n164_
  (
    .dout(new_n164__spl_),
    .din(new_n164_)
  );


  splt
  gG23
  (
    .dout(G23_spl_),
    .din(G23)
  );


  splt
  gG23_spl_
  (
    .dout(G23_spl_0),
    .din(G23_spl_)
  );


  splt
  gG23_spl_0
  (
    .dout(G23_spl_00),
    .din(G23_spl_0)
  );


  splt
  gG23_spl_00
  (
    .dout(G23_spl_000),
    .din(G23_spl_00)
  );


  splt
  gG23_spl_00
  (
    .dout(G23_spl_001),
    .din(G23_spl_00)
  );


  splt
  gG23_spl_0
  (
    .dout(G23_spl_01),
    .din(G23_spl_0)
  );


  splt
  gG23_spl_01
  (
    .dout(G23_spl_010),
    .din(G23_spl_01)
  );


  splt
  gG23_spl_01
  (
    .dout(G23_spl_011),
    .din(G23_spl_01)
  );


  splt
  gG23_spl_
  (
    .dout(G23_spl_1),
    .din(G23_spl_)
  );


  splt
  gG23_spl_1
  (
    .dout(G23_spl_10),
    .din(G23_spl_1)
  );


  splt
  gG23_spl_10
  (
    .dout(G23_spl_100),
    .din(G23_spl_10)
  );


  splt
  gG23_spl_10
  (
    .dout(G23_spl_101),
    .din(G23_spl_10)
  );


  splt
  gG23_spl_1
  (
    .dout(G23_spl_11),
    .din(G23_spl_1)
  );


  splt
  gG23_spl_11
  (
    .dout(G23_spl_110),
    .din(G23_spl_11)
  );


  splt
  gG23_spl_11
  (
    .dout(G23_spl_111),
    .din(G23_spl_11)
  );


  splt
  gG7
  (
    .dout(G7_spl_),
    .din(G7)
  );


  splt
  gG7_spl_
  (
    .dout(G7_spl_0),
    .din(G7_spl_)
  );


  splt
  gG7_spl_0
  (
    .dout(G7_spl_00),
    .din(G7_spl_0)
  );


  splt
  gG7_spl_00
  (
    .dout(G7_spl_000),
    .din(G7_spl_00)
  );


  splt
  gG7_spl_00
  (
    .dout(G7_spl_001),
    .din(G7_spl_00)
  );


  splt
  gG7_spl_0
  (
    .dout(G7_spl_01),
    .din(G7_spl_0)
  );


  splt
  gG7_spl_01
  (
    .dout(G7_spl_010),
    .din(G7_spl_01)
  );


  splt
  gG7_spl_01
  (
    .dout(G7_spl_011),
    .din(G7_spl_01)
  );


  splt
  gG7_spl_
  (
    .dout(G7_spl_1),
    .din(G7_spl_)
  );


  splt
  gG7_spl_1
  (
    .dout(G7_spl_10),
    .din(G7_spl_1)
  );


  splt
  gG7_spl_10
  (
    .dout(G7_spl_100),
    .din(G7_spl_10)
  );


  splt
  gG7_spl_10
  (
    .dout(G7_spl_101),
    .din(G7_spl_10)
  );


  splt
  gG7_spl_1
  (
    .dout(G7_spl_11),
    .din(G7_spl_1)
  );


  splt
  gG7_spl_11
  (
    .dout(G7_spl_110),
    .din(G7_spl_11)
  );


  splt
  gG7_spl_11
  (
    .dout(G7_spl_111),
    .din(G7_spl_11)
  );


  splt
  gnew_n176_
  (
    .dout(new_n176__spl_),
    .din(new_n176_)
  );


  splt
  gnew_n177_
  (
    .dout(new_n177__spl_),
    .din(new_n177_)
  );


  splt
  gnew_n178_
  (
    .dout(new_n178__spl_),
    .din(new_n178_)
  );


  splt
  gnew_n178__spl_
  (
    .dout(new_n178__spl_0),
    .din(new_n178__spl_)
  );


  splt
  gnew_n180_
  (
    .dout(new_n180__spl_),
    .din(new_n180_)
  );


  splt
  gnew_n181_
  (
    .dout(new_n181__spl_),
    .din(new_n181_)
  );


  splt
  gnew_n175_
  (
    .dout(new_n175__spl_),
    .din(new_n175_)
  );


  splt
  gnew_n183_
  (
    .dout(new_n183__spl_),
    .din(new_n183_)
  );


  splt
  gnew_n184_
  (
    .dout(new_n184__spl_),
    .din(new_n184_)
  );


  splt
  gnew_n174_
  (
    .dout(new_n174__spl_),
    .din(new_n174_)
  );


  splt
  gnew_n186_
  (
    .dout(new_n186__spl_),
    .din(new_n186_)
  );


  splt
  gnew_n187_
  (
    .dout(new_n187__spl_),
    .din(new_n187_)
  );


  splt
  gnew_n173_
  (
    .dout(new_n173__spl_),
    .din(new_n173_)
  );


  splt
  gnew_n189_
  (
    .dout(new_n189__spl_),
    .din(new_n189_)
  );


  splt
  gnew_n190_
  (
    .dout(new_n190__spl_),
    .din(new_n190_)
  );


  splt
  gnew_n172_
  (
    .dout(new_n172__spl_),
    .din(new_n172_)
  );


  splt
  gnew_n192_
  (
    .dout(new_n192__spl_),
    .din(new_n192_)
  );


  splt
  gnew_n193_
  (
    .dout(new_n193__spl_),
    .din(new_n193_)
  );


  splt
  gnew_n171_
  (
    .dout(new_n171__spl_),
    .din(new_n171_)
  );


  splt
  gnew_n195_
  (
    .dout(new_n195__spl_),
    .din(new_n195_)
  );


  splt
  gnew_n196_
  (
    .dout(new_n196__spl_),
    .din(new_n196_)
  );


  splt
  gnew_n170_
  (
    .dout(new_n170__spl_),
    .din(new_n170_)
  );


  splt
  gnew_n198_
  (
    .dout(new_n198__spl_),
    .din(new_n198_)
  );


  splt
  gnew_n199_
  (
    .dout(new_n199__spl_),
    .din(new_n199_)
  );


  splt
  gnew_n169_
  (
    .dout(new_n169__spl_),
    .din(new_n169_)
  );


  splt
  gnew_n201_
  (
    .dout(new_n201__spl_),
    .din(new_n201_)
  );


  splt
  gnew_n202_
  (
    .dout(new_n202__spl_),
    .din(new_n202_)
  );


  splt
  gnew_n168_
  (
    .dout(new_n168__spl_),
    .din(new_n168_)
  );


  splt
  gnew_n204_
  (
    .dout(new_n204__spl_),
    .din(new_n204_)
  );


  splt
  gnew_n205_
  (
    .dout(new_n205__spl_),
    .din(new_n205_)
  );


  splt
  gnew_n167_
  (
    .dout(new_n167__spl_),
    .din(new_n167_)
  );


  splt
  gnew_n207_
  (
    .dout(new_n207__spl_),
    .din(new_n207_)
  );


  splt
  gnew_n208_
  (
    .dout(new_n208__spl_),
    .din(new_n208_)
  );


  splt
  gG24
  (
    .dout(G24_spl_),
    .din(G24)
  );


  splt
  gG24_spl_
  (
    .dout(G24_spl_0),
    .din(G24_spl_)
  );


  splt
  gG24_spl_0
  (
    .dout(G24_spl_00),
    .din(G24_spl_0)
  );


  splt
  gG24_spl_00
  (
    .dout(G24_spl_000),
    .din(G24_spl_00)
  );


  splt
  gG24_spl_00
  (
    .dout(G24_spl_001),
    .din(G24_spl_00)
  );


  splt
  gG24_spl_0
  (
    .dout(G24_spl_01),
    .din(G24_spl_0)
  );


  splt
  gG24_spl_01
  (
    .dout(G24_spl_010),
    .din(G24_spl_01)
  );


  splt
  gG24_spl_01
  (
    .dout(G24_spl_011),
    .din(G24_spl_01)
  );


  splt
  gG24_spl_
  (
    .dout(G24_spl_1),
    .din(G24_spl_)
  );


  splt
  gG24_spl_1
  (
    .dout(G24_spl_10),
    .din(G24_spl_1)
  );


  splt
  gG24_spl_10
  (
    .dout(G24_spl_100),
    .din(G24_spl_10)
  );


  splt
  gG24_spl_10
  (
    .dout(G24_spl_101),
    .din(G24_spl_10)
  );


  splt
  gG24_spl_1
  (
    .dout(G24_spl_11),
    .din(G24_spl_1)
  );


  splt
  gG24_spl_11
  (
    .dout(G24_spl_110),
    .din(G24_spl_11)
  );


  splt
  gG24_spl_11
  (
    .dout(G24_spl_111),
    .din(G24_spl_11)
  );


  splt
  gG8
  (
    .dout(G8_spl_),
    .din(G8)
  );


  splt
  gG8_spl_
  (
    .dout(G8_spl_0),
    .din(G8_spl_)
  );


  splt
  gG8_spl_0
  (
    .dout(G8_spl_00),
    .din(G8_spl_0)
  );


  splt
  gG8_spl_00
  (
    .dout(G8_spl_000),
    .din(G8_spl_00)
  );


  splt
  gG8_spl_00
  (
    .dout(G8_spl_001),
    .din(G8_spl_00)
  );


  splt
  gG8_spl_0
  (
    .dout(G8_spl_01),
    .din(G8_spl_0)
  );


  splt
  gG8_spl_01
  (
    .dout(G8_spl_010),
    .din(G8_spl_01)
  );


  splt
  gG8_spl_01
  (
    .dout(G8_spl_011),
    .din(G8_spl_01)
  );


  splt
  gG8_spl_
  (
    .dout(G8_spl_1),
    .din(G8_spl_)
  );


  splt
  gG8_spl_1
  (
    .dout(G8_spl_10),
    .din(G8_spl_1)
  );


  splt
  gG8_spl_10
  (
    .dout(G8_spl_100),
    .din(G8_spl_10)
  );


  splt
  gG8_spl_10
  (
    .dout(G8_spl_101),
    .din(G8_spl_10)
  );


  splt
  gG8_spl_1
  (
    .dout(G8_spl_11),
    .din(G8_spl_1)
  );


  splt
  gG8_spl_11
  (
    .dout(G8_spl_110),
    .din(G8_spl_11)
  );


  splt
  gG8_spl_11
  (
    .dout(G8_spl_111),
    .din(G8_spl_11)
  );


  splt
  gnew_n222_
  (
    .dout(new_n222__spl_),
    .din(new_n222_)
  );


  splt
  gnew_n223_
  (
    .dout(new_n223__spl_),
    .din(new_n223_)
  );


  splt
  gnew_n224_
  (
    .dout(new_n224__spl_),
    .din(new_n224_)
  );


  splt
  gnew_n224__spl_
  (
    .dout(new_n224__spl_0),
    .din(new_n224__spl_)
  );


  splt
  gnew_n226_
  (
    .dout(new_n226__spl_),
    .din(new_n226_)
  );


  splt
  gnew_n227_
  (
    .dout(new_n227__spl_),
    .din(new_n227_)
  );


  splt
  gnew_n221_
  (
    .dout(new_n221__spl_),
    .din(new_n221_)
  );


  splt
  gnew_n229_
  (
    .dout(new_n229__spl_),
    .din(new_n229_)
  );


  splt
  gnew_n230_
  (
    .dout(new_n230__spl_),
    .din(new_n230_)
  );


  splt
  gnew_n220_
  (
    .dout(new_n220__spl_),
    .din(new_n220_)
  );


  splt
  gnew_n232_
  (
    .dout(new_n232__spl_),
    .din(new_n232_)
  );


  splt
  gnew_n233_
  (
    .dout(new_n233__spl_),
    .din(new_n233_)
  );


  splt
  gnew_n219_
  (
    .dout(new_n219__spl_),
    .din(new_n219_)
  );


  splt
  gnew_n235_
  (
    .dout(new_n235__spl_),
    .din(new_n235_)
  );


  splt
  gnew_n236_
  (
    .dout(new_n236__spl_),
    .din(new_n236_)
  );


  splt
  gnew_n218_
  (
    .dout(new_n218__spl_),
    .din(new_n218_)
  );


  splt
  gnew_n238_
  (
    .dout(new_n238__spl_),
    .din(new_n238_)
  );


  splt
  gnew_n239_
  (
    .dout(new_n239__spl_),
    .din(new_n239_)
  );


  splt
  gnew_n217_
  (
    .dout(new_n217__spl_),
    .din(new_n217_)
  );


  splt
  gnew_n241_
  (
    .dout(new_n241__spl_),
    .din(new_n241_)
  );


  splt
  gnew_n242_
  (
    .dout(new_n242__spl_),
    .din(new_n242_)
  );


  splt
  gnew_n216_
  (
    .dout(new_n216__spl_),
    .din(new_n216_)
  );


  splt
  gnew_n244_
  (
    .dout(new_n244__spl_),
    .din(new_n244_)
  );


  splt
  gnew_n245_
  (
    .dout(new_n245__spl_),
    .din(new_n245_)
  );


  splt
  gnew_n215_
  (
    .dout(new_n215__spl_),
    .din(new_n215_)
  );


  splt
  gnew_n247_
  (
    .dout(new_n247__spl_),
    .din(new_n247_)
  );


  splt
  gnew_n248_
  (
    .dout(new_n248__spl_),
    .din(new_n248_)
  );


  splt
  gnew_n214_
  (
    .dout(new_n214__spl_),
    .din(new_n214_)
  );


  splt
  gnew_n250_
  (
    .dout(new_n250__spl_),
    .din(new_n250_)
  );


  splt
  gnew_n251_
  (
    .dout(new_n251__spl_),
    .din(new_n251_)
  );


  splt
  gnew_n213_
  (
    .dout(new_n213__spl_),
    .din(new_n213_)
  );


  splt
  gnew_n253_
  (
    .dout(new_n253__spl_),
    .din(new_n253_)
  );


  splt
  gnew_n254_
  (
    .dout(new_n254__spl_),
    .din(new_n254_)
  );


  splt
  gnew_n212_
  (
    .dout(new_n212__spl_),
    .din(new_n212_)
  );


  splt
  gnew_n256_
  (
    .dout(new_n256__spl_),
    .din(new_n256_)
  );


  splt
  gnew_n257_
  (
    .dout(new_n257__spl_),
    .din(new_n257_)
  );


  splt
  gnew_n211_
  (
    .dout(new_n211__spl_),
    .din(new_n211_)
  );


  splt
  gnew_n259_
  (
    .dout(new_n259__spl_),
    .din(new_n259_)
  );


  splt
  gnew_n260_
  (
    .dout(new_n260__spl_),
    .din(new_n260_)
  );


  splt
  gG25
  (
    .dout(G25_spl_),
    .din(G25)
  );


  splt
  gG25_spl_
  (
    .dout(G25_spl_0),
    .din(G25_spl_)
  );


  splt
  gG25_spl_0
  (
    .dout(G25_spl_00),
    .din(G25_spl_0)
  );


  splt
  gG25_spl_00
  (
    .dout(G25_spl_000),
    .din(G25_spl_00)
  );


  splt
  gG25_spl_00
  (
    .dout(G25_spl_001),
    .din(G25_spl_00)
  );


  splt
  gG25_spl_0
  (
    .dout(G25_spl_01),
    .din(G25_spl_0)
  );


  splt
  gG25_spl_01
  (
    .dout(G25_spl_010),
    .din(G25_spl_01)
  );


  splt
  gG25_spl_01
  (
    .dout(G25_spl_011),
    .din(G25_spl_01)
  );


  splt
  gG25_spl_
  (
    .dout(G25_spl_1),
    .din(G25_spl_)
  );


  splt
  gG25_spl_1
  (
    .dout(G25_spl_10),
    .din(G25_spl_1)
  );


  splt
  gG25_spl_10
  (
    .dout(G25_spl_100),
    .din(G25_spl_10)
  );


  splt
  gG25_spl_10
  (
    .dout(G25_spl_101),
    .din(G25_spl_10)
  );


  splt
  gG25_spl_1
  (
    .dout(G25_spl_11),
    .din(G25_spl_1)
  );


  splt
  gG25_spl_11
  (
    .dout(G25_spl_110),
    .din(G25_spl_11)
  );


  splt
  gG25_spl_11
  (
    .dout(G25_spl_111),
    .din(G25_spl_11)
  );


  splt
  gG9
  (
    .dout(G9_spl_),
    .din(G9)
  );


  splt
  gG9_spl_
  (
    .dout(G9_spl_0),
    .din(G9_spl_)
  );


  splt
  gG9_spl_0
  (
    .dout(G9_spl_00),
    .din(G9_spl_0)
  );


  splt
  gG9_spl_00
  (
    .dout(G9_spl_000),
    .din(G9_spl_00)
  );


  splt
  gG9_spl_00
  (
    .dout(G9_spl_001),
    .din(G9_spl_00)
  );


  splt
  gG9_spl_0
  (
    .dout(G9_spl_01),
    .din(G9_spl_0)
  );


  splt
  gG9_spl_01
  (
    .dout(G9_spl_010),
    .din(G9_spl_01)
  );


  splt
  gG9_spl_01
  (
    .dout(G9_spl_011),
    .din(G9_spl_01)
  );


  splt
  gG9_spl_
  (
    .dout(G9_spl_1),
    .din(G9_spl_)
  );


  splt
  gG9_spl_1
  (
    .dout(G9_spl_10),
    .din(G9_spl_1)
  );


  splt
  gG9_spl_10
  (
    .dout(G9_spl_100),
    .din(G9_spl_10)
  );


  splt
  gG9_spl_10
  (
    .dout(G9_spl_101),
    .din(G9_spl_10)
  );


  splt
  gG9_spl_1
  (
    .dout(G9_spl_11),
    .din(G9_spl_1)
  );


  splt
  gG9_spl_11
  (
    .dout(G9_spl_110),
    .din(G9_spl_11)
  );


  splt
  gG9_spl_11
  (
    .dout(G9_spl_111),
    .din(G9_spl_11)
  );


  splt
  gnew_n276_
  (
    .dout(new_n276__spl_),
    .din(new_n276_)
  );


  splt
  gnew_n277_
  (
    .dout(new_n277__spl_),
    .din(new_n277_)
  );


  splt
  gnew_n278_
  (
    .dout(new_n278__spl_),
    .din(new_n278_)
  );


  splt
  gnew_n278__spl_
  (
    .dout(new_n278__spl_0),
    .din(new_n278__spl_)
  );


  splt
  gnew_n280_
  (
    .dout(new_n280__spl_),
    .din(new_n280_)
  );


  splt
  gnew_n281_
  (
    .dout(new_n281__spl_),
    .din(new_n281_)
  );


  splt
  gnew_n275_
  (
    .dout(new_n275__spl_),
    .din(new_n275_)
  );


  splt
  gnew_n283_
  (
    .dout(new_n283__spl_),
    .din(new_n283_)
  );


  splt
  gnew_n284_
  (
    .dout(new_n284__spl_),
    .din(new_n284_)
  );


  splt
  gnew_n274_
  (
    .dout(new_n274__spl_),
    .din(new_n274_)
  );


  splt
  gnew_n286_
  (
    .dout(new_n286__spl_),
    .din(new_n286_)
  );


  splt
  gnew_n287_
  (
    .dout(new_n287__spl_),
    .din(new_n287_)
  );


  splt
  gnew_n273_
  (
    .dout(new_n273__spl_),
    .din(new_n273_)
  );


  splt
  gnew_n289_
  (
    .dout(new_n289__spl_),
    .din(new_n289_)
  );


  splt
  gnew_n290_
  (
    .dout(new_n290__spl_),
    .din(new_n290_)
  );


  splt
  gnew_n272_
  (
    .dout(new_n272__spl_),
    .din(new_n272_)
  );


  splt
  gnew_n292_
  (
    .dout(new_n292__spl_),
    .din(new_n292_)
  );


  splt
  gnew_n293_
  (
    .dout(new_n293__spl_),
    .din(new_n293_)
  );


  splt
  gnew_n271_
  (
    .dout(new_n271__spl_),
    .din(new_n271_)
  );


  splt
  gnew_n295_
  (
    .dout(new_n295__spl_),
    .din(new_n295_)
  );


  splt
  gnew_n296_
  (
    .dout(new_n296__spl_),
    .din(new_n296_)
  );


  splt
  gnew_n270_
  (
    .dout(new_n270__spl_),
    .din(new_n270_)
  );


  splt
  gnew_n298_
  (
    .dout(new_n298__spl_),
    .din(new_n298_)
  );


  splt
  gnew_n299_
  (
    .dout(new_n299__spl_),
    .din(new_n299_)
  );


  splt
  gnew_n269_
  (
    .dout(new_n269__spl_),
    .din(new_n269_)
  );


  splt
  gnew_n301_
  (
    .dout(new_n301__spl_),
    .din(new_n301_)
  );


  splt
  gnew_n302_
  (
    .dout(new_n302__spl_),
    .din(new_n302_)
  );


  splt
  gnew_n268_
  (
    .dout(new_n268__spl_),
    .din(new_n268_)
  );


  splt
  gnew_n304_
  (
    .dout(new_n304__spl_),
    .din(new_n304_)
  );


  splt
  gnew_n305_
  (
    .dout(new_n305__spl_),
    .din(new_n305_)
  );


  splt
  gnew_n267_
  (
    .dout(new_n267__spl_),
    .din(new_n267_)
  );


  splt
  gnew_n307_
  (
    .dout(new_n307__spl_),
    .din(new_n307_)
  );


  splt
  gnew_n308_
  (
    .dout(new_n308__spl_),
    .din(new_n308_)
  );


  splt
  gnew_n266_
  (
    .dout(new_n266__spl_),
    .din(new_n266_)
  );


  splt
  gnew_n310_
  (
    .dout(new_n310__spl_),
    .din(new_n310_)
  );


  splt
  gnew_n311_
  (
    .dout(new_n311__spl_),
    .din(new_n311_)
  );


  splt
  gnew_n265_
  (
    .dout(new_n265__spl_),
    .din(new_n265_)
  );


  splt
  gnew_n313_
  (
    .dout(new_n313__spl_),
    .din(new_n313_)
  );


  splt
  gnew_n314_
  (
    .dout(new_n314__spl_),
    .din(new_n314_)
  );


  splt
  gnew_n264_
  (
    .dout(new_n264__spl_),
    .din(new_n264_)
  );


  splt
  gnew_n316_
  (
    .dout(new_n316__spl_),
    .din(new_n316_)
  );


  splt
  gnew_n317_
  (
    .dout(new_n317__spl_),
    .din(new_n317_)
  );


  splt
  gnew_n263_
  (
    .dout(new_n263__spl_),
    .din(new_n263_)
  );


  splt
  gnew_n319_
  (
    .dout(new_n319__spl_),
    .din(new_n319_)
  );


  splt
  gnew_n320_
  (
    .dout(new_n320__spl_),
    .din(new_n320_)
  );


  splt
  gG26
  (
    .dout(G26_spl_),
    .din(G26)
  );


  splt
  gG26_spl_
  (
    .dout(G26_spl_0),
    .din(G26_spl_)
  );


  splt
  gG26_spl_0
  (
    .dout(G26_spl_00),
    .din(G26_spl_0)
  );


  splt
  gG26_spl_00
  (
    .dout(G26_spl_000),
    .din(G26_spl_00)
  );


  splt
  gG26_spl_00
  (
    .dout(G26_spl_001),
    .din(G26_spl_00)
  );


  splt
  gG26_spl_0
  (
    .dout(G26_spl_01),
    .din(G26_spl_0)
  );


  splt
  gG26_spl_01
  (
    .dout(G26_spl_010),
    .din(G26_spl_01)
  );


  splt
  gG26_spl_01
  (
    .dout(G26_spl_011),
    .din(G26_spl_01)
  );


  splt
  gG26_spl_
  (
    .dout(G26_spl_1),
    .din(G26_spl_)
  );


  splt
  gG26_spl_1
  (
    .dout(G26_spl_10),
    .din(G26_spl_1)
  );


  splt
  gG26_spl_10
  (
    .dout(G26_spl_100),
    .din(G26_spl_10)
  );


  splt
  gG26_spl_10
  (
    .dout(G26_spl_101),
    .din(G26_spl_10)
  );


  splt
  gG26_spl_1
  (
    .dout(G26_spl_11),
    .din(G26_spl_1)
  );


  splt
  gG26_spl_11
  (
    .dout(G26_spl_110),
    .din(G26_spl_11)
  );


  splt
  gG26_spl_11
  (
    .dout(G26_spl_111),
    .din(G26_spl_11)
  );


  splt
  gG10
  (
    .dout(G10_spl_),
    .din(G10)
  );


  splt
  gG10_spl_
  (
    .dout(G10_spl_0),
    .din(G10_spl_)
  );


  splt
  gG10_spl_0
  (
    .dout(G10_spl_00),
    .din(G10_spl_0)
  );


  splt
  gG10_spl_00
  (
    .dout(G10_spl_000),
    .din(G10_spl_00)
  );


  splt
  gG10_spl_00
  (
    .dout(G10_spl_001),
    .din(G10_spl_00)
  );


  splt
  gG10_spl_0
  (
    .dout(G10_spl_01),
    .din(G10_spl_0)
  );


  splt
  gG10_spl_01
  (
    .dout(G10_spl_010),
    .din(G10_spl_01)
  );


  splt
  gG10_spl_01
  (
    .dout(G10_spl_011),
    .din(G10_spl_01)
  );


  splt
  gG10_spl_
  (
    .dout(G10_spl_1),
    .din(G10_spl_)
  );


  splt
  gG10_spl_1
  (
    .dout(G10_spl_10),
    .din(G10_spl_1)
  );


  splt
  gG10_spl_10
  (
    .dout(G10_spl_100),
    .din(G10_spl_10)
  );


  splt
  gG10_spl_10
  (
    .dout(G10_spl_101),
    .din(G10_spl_10)
  );


  splt
  gG10_spl_1
  (
    .dout(G10_spl_11),
    .din(G10_spl_1)
  );


  splt
  gG10_spl_11
  (
    .dout(G10_spl_110),
    .din(G10_spl_11)
  );


  splt
  gG10_spl_11
  (
    .dout(G10_spl_111),
    .din(G10_spl_11)
  );


  splt
  gnew_n338_
  (
    .dout(new_n338__spl_),
    .din(new_n338_)
  );


  splt
  gnew_n339_
  (
    .dout(new_n339__spl_),
    .din(new_n339_)
  );


  splt
  gnew_n340_
  (
    .dout(new_n340__spl_),
    .din(new_n340_)
  );


  splt
  gnew_n340__spl_
  (
    .dout(new_n340__spl_0),
    .din(new_n340__spl_)
  );


  splt
  gnew_n342_
  (
    .dout(new_n342__spl_),
    .din(new_n342_)
  );


  splt
  gnew_n343_
  (
    .dout(new_n343__spl_),
    .din(new_n343_)
  );


  splt
  gnew_n337_
  (
    .dout(new_n337__spl_),
    .din(new_n337_)
  );


  splt
  gnew_n345_
  (
    .dout(new_n345__spl_),
    .din(new_n345_)
  );


  splt
  gnew_n346_
  (
    .dout(new_n346__spl_),
    .din(new_n346_)
  );


  splt
  gnew_n336_
  (
    .dout(new_n336__spl_),
    .din(new_n336_)
  );


  splt
  gnew_n348_
  (
    .dout(new_n348__spl_),
    .din(new_n348_)
  );


  splt
  gnew_n349_
  (
    .dout(new_n349__spl_),
    .din(new_n349_)
  );


  splt
  gnew_n335_
  (
    .dout(new_n335__spl_),
    .din(new_n335_)
  );


  splt
  gnew_n351_
  (
    .dout(new_n351__spl_),
    .din(new_n351_)
  );


  splt
  gnew_n352_
  (
    .dout(new_n352__spl_),
    .din(new_n352_)
  );


  splt
  gnew_n334_
  (
    .dout(new_n334__spl_),
    .din(new_n334_)
  );


  splt
  gnew_n354_
  (
    .dout(new_n354__spl_),
    .din(new_n354_)
  );


  splt
  gnew_n355_
  (
    .dout(new_n355__spl_),
    .din(new_n355_)
  );


  splt
  gnew_n333_
  (
    .dout(new_n333__spl_),
    .din(new_n333_)
  );


  splt
  gnew_n357_
  (
    .dout(new_n357__spl_),
    .din(new_n357_)
  );


  splt
  gnew_n358_
  (
    .dout(new_n358__spl_),
    .din(new_n358_)
  );


  splt
  gnew_n332_
  (
    .dout(new_n332__spl_),
    .din(new_n332_)
  );


  splt
  gnew_n360_
  (
    .dout(new_n360__spl_),
    .din(new_n360_)
  );


  splt
  gnew_n361_
  (
    .dout(new_n361__spl_),
    .din(new_n361_)
  );


  splt
  gnew_n331_
  (
    .dout(new_n331__spl_),
    .din(new_n331_)
  );


  splt
  gnew_n363_
  (
    .dout(new_n363__spl_),
    .din(new_n363_)
  );


  splt
  gnew_n364_
  (
    .dout(new_n364__spl_),
    .din(new_n364_)
  );


  splt
  gnew_n330_
  (
    .dout(new_n330__spl_),
    .din(new_n330_)
  );


  splt
  gnew_n366_
  (
    .dout(new_n366__spl_),
    .din(new_n366_)
  );


  splt
  gnew_n367_
  (
    .dout(new_n367__spl_),
    .din(new_n367_)
  );


  splt
  gnew_n329_
  (
    .dout(new_n329__spl_),
    .din(new_n329_)
  );


  splt
  gnew_n369_
  (
    .dout(new_n369__spl_),
    .din(new_n369_)
  );


  splt
  gnew_n370_
  (
    .dout(new_n370__spl_),
    .din(new_n370_)
  );


  splt
  gnew_n328_
  (
    .dout(new_n328__spl_),
    .din(new_n328_)
  );


  splt
  gnew_n372_
  (
    .dout(new_n372__spl_),
    .din(new_n372_)
  );


  splt
  gnew_n373_
  (
    .dout(new_n373__spl_),
    .din(new_n373_)
  );


  splt
  gnew_n327_
  (
    .dout(new_n327__spl_),
    .din(new_n327_)
  );


  splt
  gnew_n375_
  (
    .dout(new_n375__spl_),
    .din(new_n375_)
  );


  splt
  gnew_n376_
  (
    .dout(new_n376__spl_),
    .din(new_n376_)
  );


  splt
  gnew_n326_
  (
    .dout(new_n326__spl_),
    .din(new_n326_)
  );


  splt
  gnew_n378_
  (
    .dout(new_n378__spl_),
    .din(new_n378_)
  );


  splt
  gnew_n379_
  (
    .dout(new_n379__spl_),
    .din(new_n379_)
  );


  splt
  gnew_n325_
  (
    .dout(new_n325__spl_),
    .din(new_n325_)
  );


  splt
  gnew_n381_
  (
    .dout(new_n381__spl_),
    .din(new_n381_)
  );


  splt
  gnew_n382_
  (
    .dout(new_n382__spl_),
    .din(new_n382_)
  );


  splt
  gnew_n324_
  (
    .dout(new_n324__spl_),
    .din(new_n324_)
  );


  splt
  gnew_n384_
  (
    .dout(new_n384__spl_),
    .din(new_n384_)
  );


  splt
  gnew_n385_
  (
    .dout(new_n385__spl_),
    .din(new_n385_)
  );


  splt
  gnew_n323_
  (
    .dout(new_n323__spl_),
    .din(new_n323_)
  );


  splt
  gnew_n387_
  (
    .dout(new_n387__spl_),
    .din(new_n387_)
  );


  splt
  gnew_n388_
  (
    .dout(new_n388__spl_),
    .din(new_n388_)
  );


  splt
  gG27
  (
    .dout(G27_spl_),
    .din(G27)
  );


  splt
  gG27_spl_
  (
    .dout(G27_spl_0),
    .din(G27_spl_)
  );


  splt
  gG27_spl_0
  (
    .dout(G27_spl_00),
    .din(G27_spl_0)
  );


  splt
  gG27_spl_00
  (
    .dout(G27_spl_000),
    .din(G27_spl_00)
  );


  splt
  gG27_spl_00
  (
    .dout(G27_spl_001),
    .din(G27_spl_00)
  );


  splt
  gG27_spl_0
  (
    .dout(G27_spl_01),
    .din(G27_spl_0)
  );


  splt
  gG27_spl_01
  (
    .dout(G27_spl_010),
    .din(G27_spl_01)
  );


  splt
  gG27_spl_01
  (
    .dout(G27_spl_011),
    .din(G27_spl_01)
  );


  splt
  gG27_spl_
  (
    .dout(G27_spl_1),
    .din(G27_spl_)
  );


  splt
  gG27_spl_1
  (
    .dout(G27_spl_10),
    .din(G27_spl_1)
  );


  splt
  gG27_spl_10
  (
    .dout(G27_spl_100),
    .din(G27_spl_10)
  );


  splt
  gG27_spl_10
  (
    .dout(G27_spl_101),
    .din(G27_spl_10)
  );


  splt
  gG27_spl_1
  (
    .dout(G27_spl_11),
    .din(G27_spl_1)
  );


  splt
  gG27_spl_11
  (
    .dout(G27_spl_110),
    .din(G27_spl_11)
  );


  splt
  gG27_spl_11
  (
    .dout(G27_spl_111),
    .din(G27_spl_11)
  );


  splt
  gG11
  (
    .dout(G11_spl_),
    .din(G11)
  );


  splt
  gG11_spl_
  (
    .dout(G11_spl_0),
    .din(G11_spl_)
  );


  splt
  gG11_spl_0
  (
    .dout(G11_spl_00),
    .din(G11_spl_0)
  );


  splt
  gG11_spl_00
  (
    .dout(G11_spl_000),
    .din(G11_spl_00)
  );


  splt
  gG11_spl_00
  (
    .dout(G11_spl_001),
    .din(G11_spl_00)
  );


  splt
  gG11_spl_0
  (
    .dout(G11_spl_01),
    .din(G11_spl_0)
  );


  splt
  gG11_spl_01
  (
    .dout(G11_spl_010),
    .din(G11_spl_01)
  );


  splt
  gG11_spl_01
  (
    .dout(G11_spl_011),
    .din(G11_spl_01)
  );


  splt
  gG11_spl_
  (
    .dout(G11_spl_1),
    .din(G11_spl_)
  );


  splt
  gG11_spl_1
  (
    .dout(G11_spl_10),
    .din(G11_spl_1)
  );


  splt
  gG11_spl_10
  (
    .dout(G11_spl_100),
    .din(G11_spl_10)
  );


  splt
  gG11_spl_10
  (
    .dout(G11_spl_101),
    .din(G11_spl_10)
  );


  splt
  gG11_spl_1
  (
    .dout(G11_spl_11),
    .din(G11_spl_1)
  );


  splt
  gG11_spl_11
  (
    .dout(G11_spl_110),
    .din(G11_spl_11)
  );


  splt
  gG11_spl_11
  (
    .dout(G11_spl_111),
    .din(G11_spl_11)
  );


  splt
  gnew_n408_
  (
    .dout(new_n408__spl_),
    .din(new_n408_)
  );


  splt
  gnew_n409_
  (
    .dout(new_n409__spl_),
    .din(new_n409_)
  );


  splt
  gnew_n410_
  (
    .dout(new_n410__spl_),
    .din(new_n410_)
  );


  splt
  gnew_n410__spl_
  (
    .dout(new_n410__spl_0),
    .din(new_n410__spl_)
  );


  splt
  gnew_n412_
  (
    .dout(new_n412__spl_),
    .din(new_n412_)
  );


  splt
  gnew_n413_
  (
    .dout(new_n413__spl_),
    .din(new_n413_)
  );


  splt
  gnew_n407_
  (
    .dout(new_n407__spl_),
    .din(new_n407_)
  );


  splt
  gnew_n415_
  (
    .dout(new_n415__spl_),
    .din(new_n415_)
  );


  splt
  gnew_n416_
  (
    .dout(new_n416__spl_),
    .din(new_n416_)
  );


  splt
  gnew_n406_
  (
    .dout(new_n406__spl_),
    .din(new_n406_)
  );


  splt
  gnew_n418_
  (
    .dout(new_n418__spl_),
    .din(new_n418_)
  );


  splt
  gnew_n419_
  (
    .dout(new_n419__spl_),
    .din(new_n419_)
  );


  splt
  gnew_n405_
  (
    .dout(new_n405__spl_),
    .din(new_n405_)
  );


  splt
  gnew_n421_
  (
    .dout(new_n421__spl_),
    .din(new_n421_)
  );


  splt
  gnew_n422_
  (
    .dout(new_n422__spl_),
    .din(new_n422_)
  );


  splt
  gnew_n404_
  (
    .dout(new_n404__spl_),
    .din(new_n404_)
  );


  splt
  gnew_n424_
  (
    .dout(new_n424__spl_),
    .din(new_n424_)
  );


  splt
  gnew_n425_
  (
    .dout(new_n425__spl_),
    .din(new_n425_)
  );


  splt
  gnew_n403_
  (
    .dout(new_n403__spl_),
    .din(new_n403_)
  );


  splt
  gnew_n427_
  (
    .dout(new_n427__spl_),
    .din(new_n427_)
  );


  splt
  gnew_n428_
  (
    .dout(new_n428__spl_),
    .din(new_n428_)
  );


  splt
  gnew_n402_
  (
    .dout(new_n402__spl_),
    .din(new_n402_)
  );


  splt
  gnew_n430_
  (
    .dout(new_n430__spl_),
    .din(new_n430_)
  );


  splt
  gnew_n431_
  (
    .dout(new_n431__spl_),
    .din(new_n431_)
  );


  splt
  gnew_n401_
  (
    .dout(new_n401__spl_),
    .din(new_n401_)
  );


  splt
  gnew_n433_
  (
    .dout(new_n433__spl_),
    .din(new_n433_)
  );


  splt
  gnew_n434_
  (
    .dout(new_n434__spl_),
    .din(new_n434_)
  );


  splt
  gnew_n400_
  (
    .dout(new_n400__spl_),
    .din(new_n400_)
  );


  splt
  gnew_n436_
  (
    .dout(new_n436__spl_),
    .din(new_n436_)
  );


  splt
  gnew_n437_
  (
    .dout(new_n437__spl_),
    .din(new_n437_)
  );


  splt
  gnew_n399_
  (
    .dout(new_n399__spl_),
    .din(new_n399_)
  );


  splt
  gnew_n439_
  (
    .dout(new_n439__spl_),
    .din(new_n439_)
  );


  splt
  gnew_n440_
  (
    .dout(new_n440__spl_),
    .din(new_n440_)
  );


  splt
  gnew_n398_
  (
    .dout(new_n398__spl_),
    .din(new_n398_)
  );


  splt
  gnew_n442_
  (
    .dout(new_n442__spl_),
    .din(new_n442_)
  );


  splt
  gnew_n443_
  (
    .dout(new_n443__spl_),
    .din(new_n443_)
  );


  splt
  gnew_n397_
  (
    .dout(new_n397__spl_),
    .din(new_n397_)
  );


  splt
  gnew_n445_
  (
    .dout(new_n445__spl_),
    .din(new_n445_)
  );


  splt
  gnew_n446_
  (
    .dout(new_n446__spl_),
    .din(new_n446_)
  );


  splt
  gnew_n396_
  (
    .dout(new_n396__spl_),
    .din(new_n396_)
  );


  splt
  gnew_n448_
  (
    .dout(new_n448__spl_),
    .din(new_n448_)
  );


  splt
  gnew_n449_
  (
    .dout(new_n449__spl_),
    .din(new_n449_)
  );


  splt
  gnew_n395_
  (
    .dout(new_n395__spl_),
    .din(new_n395_)
  );


  splt
  gnew_n451_
  (
    .dout(new_n451__spl_),
    .din(new_n451_)
  );


  splt
  gnew_n452_
  (
    .dout(new_n452__spl_),
    .din(new_n452_)
  );


  splt
  gnew_n394_
  (
    .dout(new_n394__spl_),
    .din(new_n394_)
  );


  splt
  gnew_n454_
  (
    .dout(new_n454__spl_),
    .din(new_n454_)
  );


  splt
  gnew_n455_
  (
    .dout(new_n455__spl_),
    .din(new_n455_)
  );


  splt
  gnew_n393_
  (
    .dout(new_n393__spl_),
    .din(new_n393_)
  );


  splt
  gnew_n457_
  (
    .dout(new_n457__spl_),
    .din(new_n457_)
  );


  splt
  gnew_n458_
  (
    .dout(new_n458__spl_),
    .din(new_n458_)
  );


  splt
  gnew_n392_
  (
    .dout(new_n392__spl_),
    .din(new_n392_)
  );


  splt
  gnew_n460_
  (
    .dout(new_n460__spl_),
    .din(new_n460_)
  );


  splt
  gnew_n461_
  (
    .dout(new_n461__spl_),
    .din(new_n461_)
  );


  splt
  gnew_n391_
  (
    .dout(new_n391__spl_),
    .din(new_n391_)
  );


  splt
  gnew_n463_
  (
    .dout(new_n463__spl_),
    .din(new_n463_)
  );


  splt
  gnew_n464_
  (
    .dout(new_n464__spl_),
    .din(new_n464_)
  );


  splt
  gG28
  (
    .dout(G28_spl_),
    .din(G28)
  );


  splt
  gG28_spl_
  (
    .dout(G28_spl_0),
    .din(G28_spl_)
  );


  splt
  gG28_spl_0
  (
    .dout(G28_spl_00),
    .din(G28_spl_0)
  );


  splt
  gG28_spl_00
  (
    .dout(G28_spl_000),
    .din(G28_spl_00)
  );


  splt
  gG28_spl_00
  (
    .dout(G28_spl_001),
    .din(G28_spl_00)
  );


  splt
  gG28_spl_0
  (
    .dout(G28_spl_01),
    .din(G28_spl_0)
  );


  splt
  gG28_spl_01
  (
    .dout(G28_spl_010),
    .din(G28_spl_01)
  );


  splt
  gG28_spl_01
  (
    .dout(G28_spl_011),
    .din(G28_spl_01)
  );


  splt
  gG28_spl_
  (
    .dout(G28_spl_1),
    .din(G28_spl_)
  );


  splt
  gG28_spl_1
  (
    .dout(G28_spl_10),
    .din(G28_spl_1)
  );


  splt
  gG28_spl_10
  (
    .dout(G28_spl_100),
    .din(G28_spl_10)
  );


  splt
  gG28_spl_10
  (
    .dout(G28_spl_101),
    .din(G28_spl_10)
  );


  splt
  gG28_spl_1
  (
    .dout(G28_spl_11),
    .din(G28_spl_1)
  );


  splt
  gG28_spl_11
  (
    .dout(G28_spl_110),
    .din(G28_spl_11)
  );


  splt
  gG28_spl_11
  (
    .dout(G28_spl_111),
    .din(G28_spl_11)
  );


  splt
  gG12
  (
    .dout(G12_spl_),
    .din(G12)
  );


  splt
  gG12_spl_
  (
    .dout(G12_spl_0),
    .din(G12_spl_)
  );


  splt
  gG12_spl_0
  (
    .dout(G12_spl_00),
    .din(G12_spl_0)
  );


  splt
  gG12_spl_00
  (
    .dout(G12_spl_000),
    .din(G12_spl_00)
  );


  splt
  gG12_spl_00
  (
    .dout(G12_spl_001),
    .din(G12_spl_00)
  );


  splt
  gG12_spl_0
  (
    .dout(G12_spl_01),
    .din(G12_spl_0)
  );


  splt
  gG12_spl_01
  (
    .dout(G12_spl_010),
    .din(G12_spl_01)
  );


  splt
  gG12_spl_01
  (
    .dout(G12_spl_011),
    .din(G12_spl_01)
  );


  splt
  gG12_spl_
  (
    .dout(G12_spl_1),
    .din(G12_spl_)
  );


  splt
  gG12_spl_1
  (
    .dout(G12_spl_10),
    .din(G12_spl_1)
  );


  splt
  gG12_spl_10
  (
    .dout(G12_spl_100),
    .din(G12_spl_10)
  );


  splt
  gG12_spl_10
  (
    .dout(G12_spl_101),
    .din(G12_spl_10)
  );


  splt
  gG12_spl_1
  (
    .dout(G12_spl_11),
    .din(G12_spl_1)
  );


  splt
  gG12_spl_11
  (
    .dout(G12_spl_110),
    .din(G12_spl_11)
  );


  splt
  gG12_spl_11
  (
    .dout(G12_spl_111),
    .din(G12_spl_11)
  );


  splt
  gnew_n486_
  (
    .dout(new_n486__spl_),
    .din(new_n486_)
  );


  splt
  gnew_n487_
  (
    .dout(new_n487__spl_),
    .din(new_n487_)
  );


  splt
  gnew_n488_
  (
    .dout(new_n488__spl_),
    .din(new_n488_)
  );


  splt
  gnew_n488__spl_
  (
    .dout(new_n488__spl_0),
    .din(new_n488__spl_)
  );


  splt
  gnew_n490_
  (
    .dout(new_n490__spl_),
    .din(new_n490_)
  );


  splt
  gnew_n491_
  (
    .dout(new_n491__spl_),
    .din(new_n491_)
  );


  splt
  gnew_n485_
  (
    .dout(new_n485__spl_),
    .din(new_n485_)
  );


  splt
  gnew_n493_
  (
    .dout(new_n493__spl_),
    .din(new_n493_)
  );


  splt
  gnew_n494_
  (
    .dout(new_n494__spl_),
    .din(new_n494_)
  );


  splt
  gnew_n484_
  (
    .dout(new_n484__spl_),
    .din(new_n484_)
  );


  splt
  gnew_n496_
  (
    .dout(new_n496__spl_),
    .din(new_n496_)
  );


  splt
  gnew_n497_
  (
    .dout(new_n497__spl_),
    .din(new_n497_)
  );


  splt
  gnew_n483_
  (
    .dout(new_n483__spl_),
    .din(new_n483_)
  );


  splt
  gnew_n499_
  (
    .dout(new_n499__spl_),
    .din(new_n499_)
  );


  splt
  gnew_n500_
  (
    .dout(new_n500__spl_),
    .din(new_n500_)
  );


  splt
  gnew_n482_
  (
    .dout(new_n482__spl_),
    .din(new_n482_)
  );


  splt
  gnew_n502_
  (
    .dout(new_n502__spl_),
    .din(new_n502_)
  );


  splt
  gnew_n503_
  (
    .dout(new_n503__spl_),
    .din(new_n503_)
  );


  splt
  gnew_n481_
  (
    .dout(new_n481__spl_),
    .din(new_n481_)
  );


  splt
  gnew_n505_
  (
    .dout(new_n505__spl_),
    .din(new_n505_)
  );


  splt
  gnew_n506_
  (
    .dout(new_n506__spl_),
    .din(new_n506_)
  );


  splt
  gnew_n480_
  (
    .dout(new_n480__spl_),
    .din(new_n480_)
  );


  splt
  gnew_n508_
  (
    .dout(new_n508__spl_),
    .din(new_n508_)
  );


  splt
  gnew_n509_
  (
    .dout(new_n509__spl_),
    .din(new_n509_)
  );


  splt
  gnew_n479_
  (
    .dout(new_n479__spl_),
    .din(new_n479_)
  );


  splt
  gnew_n511_
  (
    .dout(new_n511__spl_),
    .din(new_n511_)
  );


  splt
  gnew_n512_
  (
    .dout(new_n512__spl_),
    .din(new_n512_)
  );


  splt
  gnew_n478_
  (
    .dout(new_n478__spl_),
    .din(new_n478_)
  );


  splt
  gnew_n514_
  (
    .dout(new_n514__spl_),
    .din(new_n514_)
  );


  splt
  gnew_n515_
  (
    .dout(new_n515__spl_),
    .din(new_n515_)
  );


  splt
  gnew_n477_
  (
    .dout(new_n477__spl_),
    .din(new_n477_)
  );


  splt
  gnew_n517_
  (
    .dout(new_n517__spl_),
    .din(new_n517_)
  );


  splt
  gnew_n518_
  (
    .dout(new_n518__spl_),
    .din(new_n518_)
  );


  splt
  gnew_n476_
  (
    .dout(new_n476__spl_),
    .din(new_n476_)
  );


  splt
  gnew_n520_
  (
    .dout(new_n520__spl_),
    .din(new_n520_)
  );


  splt
  gnew_n521_
  (
    .dout(new_n521__spl_),
    .din(new_n521_)
  );


  splt
  gnew_n475_
  (
    .dout(new_n475__spl_),
    .din(new_n475_)
  );


  splt
  gnew_n523_
  (
    .dout(new_n523__spl_),
    .din(new_n523_)
  );


  splt
  gnew_n524_
  (
    .dout(new_n524__spl_),
    .din(new_n524_)
  );


  splt
  gnew_n474_
  (
    .dout(new_n474__spl_),
    .din(new_n474_)
  );


  splt
  gnew_n526_
  (
    .dout(new_n526__spl_),
    .din(new_n526_)
  );


  splt
  gnew_n527_
  (
    .dout(new_n527__spl_),
    .din(new_n527_)
  );


  splt
  gnew_n473_
  (
    .dout(new_n473__spl_),
    .din(new_n473_)
  );


  splt
  gnew_n529_
  (
    .dout(new_n529__spl_),
    .din(new_n529_)
  );


  splt
  gnew_n530_
  (
    .dout(new_n530__spl_),
    .din(new_n530_)
  );


  splt
  gnew_n472_
  (
    .dout(new_n472__spl_),
    .din(new_n472_)
  );


  splt
  gnew_n532_
  (
    .dout(new_n532__spl_),
    .din(new_n532_)
  );


  splt
  gnew_n533_
  (
    .dout(new_n533__spl_),
    .din(new_n533_)
  );


  splt
  gnew_n471_
  (
    .dout(new_n471__spl_),
    .din(new_n471_)
  );


  splt
  gnew_n535_
  (
    .dout(new_n535__spl_),
    .din(new_n535_)
  );


  splt
  gnew_n536_
  (
    .dout(new_n536__spl_),
    .din(new_n536_)
  );


  splt
  gnew_n470_
  (
    .dout(new_n470__spl_),
    .din(new_n470_)
  );


  splt
  gnew_n538_
  (
    .dout(new_n538__spl_),
    .din(new_n538_)
  );


  splt
  gnew_n539_
  (
    .dout(new_n539__spl_),
    .din(new_n539_)
  );


  splt
  gnew_n469_
  (
    .dout(new_n469__spl_),
    .din(new_n469_)
  );


  splt
  gnew_n541_
  (
    .dout(new_n541__spl_),
    .din(new_n541_)
  );


  splt
  gnew_n542_
  (
    .dout(new_n542__spl_),
    .din(new_n542_)
  );


  splt
  gnew_n468_
  (
    .dout(new_n468__spl_),
    .din(new_n468_)
  );


  splt
  gnew_n544_
  (
    .dout(new_n544__spl_),
    .din(new_n544_)
  );


  splt
  gnew_n545_
  (
    .dout(new_n545__spl_),
    .din(new_n545_)
  );


  splt
  gnew_n467_
  (
    .dout(new_n467__spl_),
    .din(new_n467_)
  );


  splt
  gnew_n547_
  (
    .dout(new_n547__spl_),
    .din(new_n547_)
  );


  splt
  gnew_n548_
  (
    .dout(new_n548__spl_),
    .din(new_n548_)
  );


  splt
  gG29
  (
    .dout(G29_spl_),
    .din(G29)
  );


  splt
  gG29_spl_
  (
    .dout(G29_spl_0),
    .din(G29_spl_)
  );


  splt
  gG29_spl_0
  (
    .dout(G29_spl_00),
    .din(G29_spl_0)
  );


  splt
  gG29_spl_00
  (
    .dout(G29_spl_000),
    .din(G29_spl_00)
  );


  splt
  gG29_spl_00
  (
    .dout(G29_spl_001),
    .din(G29_spl_00)
  );


  splt
  gG29_spl_0
  (
    .dout(G29_spl_01),
    .din(G29_spl_0)
  );


  splt
  gG29_spl_01
  (
    .dout(G29_spl_010),
    .din(G29_spl_01)
  );


  splt
  gG29_spl_01
  (
    .dout(G29_spl_011),
    .din(G29_spl_01)
  );


  splt
  gG29_spl_
  (
    .dout(G29_spl_1),
    .din(G29_spl_)
  );


  splt
  gG29_spl_1
  (
    .dout(G29_spl_10),
    .din(G29_spl_1)
  );


  splt
  gG29_spl_10
  (
    .dout(G29_spl_100),
    .din(G29_spl_10)
  );


  splt
  gG29_spl_10
  (
    .dout(G29_spl_101),
    .din(G29_spl_10)
  );


  splt
  gG29_spl_1
  (
    .dout(G29_spl_11),
    .din(G29_spl_1)
  );


  splt
  gG29_spl_11
  (
    .dout(G29_spl_110),
    .din(G29_spl_11)
  );


  splt
  gG29_spl_11
  (
    .dout(G29_spl_111),
    .din(G29_spl_11)
  );


  splt
  gG13
  (
    .dout(G13_spl_),
    .din(G13)
  );


  splt
  gG13_spl_
  (
    .dout(G13_spl_0),
    .din(G13_spl_)
  );


  splt
  gG13_spl_0
  (
    .dout(G13_spl_00),
    .din(G13_spl_0)
  );


  splt
  gG13_spl_00
  (
    .dout(G13_spl_000),
    .din(G13_spl_00)
  );


  splt
  gG13_spl_00
  (
    .dout(G13_spl_001),
    .din(G13_spl_00)
  );


  splt
  gG13_spl_0
  (
    .dout(G13_spl_01),
    .din(G13_spl_0)
  );


  splt
  gG13_spl_01
  (
    .dout(G13_spl_010),
    .din(G13_spl_01)
  );


  splt
  gG13_spl_01
  (
    .dout(G13_spl_011),
    .din(G13_spl_01)
  );


  splt
  gG13_spl_
  (
    .dout(G13_spl_1),
    .din(G13_spl_)
  );


  splt
  gG13_spl_1
  (
    .dout(G13_spl_10),
    .din(G13_spl_1)
  );


  splt
  gG13_spl_10
  (
    .dout(G13_spl_100),
    .din(G13_spl_10)
  );


  splt
  gG13_spl_10
  (
    .dout(G13_spl_101),
    .din(G13_spl_10)
  );


  splt
  gG13_spl_1
  (
    .dout(G13_spl_11),
    .din(G13_spl_1)
  );


  splt
  gG13_spl_11
  (
    .dout(G13_spl_110),
    .din(G13_spl_11)
  );


  splt
  gG13_spl_11
  (
    .dout(G13_spl_111),
    .din(G13_spl_11)
  );


  splt
  gnew_n572_
  (
    .dout(new_n572__spl_),
    .din(new_n572_)
  );


  splt
  gnew_n573_
  (
    .dout(new_n573__spl_),
    .din(new_n573_)
  );


  splt
  gnew_n574_
  (
    .dout(new_n574__spl_),
    .din(new_n574_)
  );


  splt
  gnew_n574__spl_
  (
    .dout(new_n574__spl_0),
    .din(new_n574__spl_)
  );


  splt
  gnew_n576_
  (
    .dout(new_n576__spl_),
    .din(new_n576_)
  );


  splt
  gnew_n577_
  (
    .dout(new_n577__spl_),
    .din(new_n577_)
  );


  splt
  gnew_n571_
  (
    .dout(new_n571__spl_),
    .din(new_n571_)
  );


  splt
  gnew_n579_
  (
    .dout(new_n579__spl_),
    .din(new_n579_)
  );


  splt
  gnew_n580_
  (
    .dout(new_n580__spl_),
    .din(new_n580_)
  );


  splt
  gnew_n570_
  (
    .dout(new_n570__spl_),
    .din(new_n570_)
  );


  splt
  gnew_n582_
  (
    .dout(new_n582__spl_),
    .din(new_n582_)
  );


  splt
  gnew_n583_
  (
    .dout(new_n583__spl_),
    .din(new_n583_)
  );


  splt
  gnew_n569_
  (
    .dout(new_n569__spl_),
    .din(new_n569_)
  );


  splt
  gnew_n585_
  (
    .dout(new_n585__spl_),
    .din(new_n585_)
  );


  splt
  gnew_n586_
  (
    .dout(new_n586__spl_),
    .din(new_n586_)
  );


  splt
  gnew_n568_
  (
    .dout(new_n568__spl_),
    .din(new_n568_)
  );


  splt
  gnew_n588_
  (
    .dout(new_n588__spl_),
    .din(new_n588_)
  );


  splt
  gnew_n589_
  (
    .dout(new_n589__spl_),
    .din(new_n589_)
  );


  splt
  gnew_n567_
  (
    .dout(new_n567__spl_),
    .din(new_n567_)
  );


  splt
  gnew_n591_
  (
    .dout(new_n591__spl_),
    .din(new_n591_)
  );


  splt
  gnew_n592_
  (
    .dout(new_n592__spl_),
    .din(new_n592_)
  );


  splt
  gnew_n566_
  (
    .dout(new_n566__spl_),
    .din(new_n566_)
  );


  splt
  gnew_n594_
  (
    .dout(new_n594__spl_),
    .din(new_n594_)
  );


  splt
  gnew_n595_
  (
    .dout(new_n595__spl_),
    .din(new_n595_)
  );


  splt
  gnew_n565_
  (
    .dout(new_n565__spl_),
    .din(new_n565_)
  );


  splt
  gnew_n597_
  (
    .dout(new_n597__spl_),
    .din(new_n597_)
  );


  splt
  gnew_n598_
  (
    .dout(new_n598__spl_),
    .din(new_n598_)
  );


  splt
  gnew_n564_
  (
    .dout(new_n564__spl_),
    .din(new_n564_)
  );


  splt
  gnew_n600_
  (
    .dout(new_n600__spl_),
    .din(new_n600_)
  );


  splt
  gnew_n601_
  (
    .dout(new_n601__spl_),
    .din(new_n601_)
  );


  splt
  gnew_n563_
  (
    .dout(new_n563__spl_),
    .din(new_n563_)
  );


  splt
  gnew_n603_
  (
    .dout(new_n603__spl_),
    .din(new_n603_)
  );


  splt
  gnew_n604_
  (
    .dout(new_n604__spl_),
    .din(new_n604_)
  );


  splt
  gnew_n562_
  (
    .dout(new_n562__spl_),
    .din(new_n562_)
  );


  splt
  gnew_n606_
  (
    .dout(new_n606__spl_),
    .din(new_n606_)
  );


  splt
  gnew_n607_
  (
    .dout(new_n607__spl_),
    .din(new_n607_)
  );


  splt
  gnew_n561_
  (
    .dout(new_n561__spl_),
    .din(new_n561_)
  );


  splt
  gnew_n609_
  (
    .dout(new_n609__spl_),
    .din(new_n609_)
  );


  splt
  gnew_n610_
  (
    .dout(new_n610__spl_),
    .din(new_n610_)
  );


  splt
  gnew_n560_
  (
    .dout(new_n560__spl_),
    .din(new_n560_)
  );


  splt
  gnew_n612_
  (
    .dout(new_n612__spl_),
    .din(new_n612_)
  );


  splt
  gnew_n613_
  (
    .dout(new_n613__spl_),
    .din(new_n613_)
  );


  splt
  gnew_n559_
  (
    .dout(new_n559__spl_),
    .din(new_n559_)
  );


  splt
  gnew_n615_
  (
    .dout(new_n615__spl_),
    .din(new_n615_)
  );


  splt
  gnew_n616_
  (
    .dout(new_n616__spl_),
    .din(new_n616_)
  );


  splt
  gnew_n558_
  (
    .dout(new_n558__spl_),
    .din(new_n558_)
  );


  splt
  gnew_n618_
  (
    .dout(new_n618__spl_),
    .din(new_n618_)
  );


  splt
  gnew_n619_
  (
    .dout(new_n619__spl_),
    .din(new_n619_)
  );


  splt
  gnew_n557_
  (
    .dout(new_n557__spl_),
    .din(new_n557_)
  );


  splt
  gnew_n621_
  (
    .dout(new_n621__spl_),
    .din(new_n621_)
  );


  splt
  gnew_n622_
  (
    .dout(new_n622__spl_),
    .din(new_n622_)
  );


  splt
  gnew_n556_
  (
    .dout(new_n556__spl_),
    .din(new_n556_)
  );


  splt
  gnew_n624_
  (
    .dout(new_n624__spl_),
    .din(new_n624_)
  );


  splt
  gnew_n625_
  (
    .dout(new_n625__spl_),
    .din(new_n625_)
  );


  splt
  gnew_n555_
  (
    .dout(new_n555__spl_),
    .din(new_n555_)
  );


  splt
  gnew_n627_
  (
    .dout(new_n627__spl_),
    .din(new_n627_)
  );


  splt
  gnew_n628_
  (
    .dout(new_n628__spl_),
    .din(new_n628_)
  );


  splt
  gnew_n554_
  (
    .dout(new_n554__spl_),
    .din(new_n554_)
  );


  splt
  gnew_n630_
  (
    .dout(new_n630__spl_),
    .din(new_n630_)
  );


  splt
  gnew_n631_
  (
    .dout(new_n631__spl_),
    .din(new_n631_)
  );


  splt
  gnew_n553_
  (
    .dout(new_n553__spl_),
    .din(new_n553_)
  );


  splt
  gnew_n633_
  (
    .dout(new_n633__spl_),
    .din(new_n633_)
  );


  splt
  gnew_n634_
  (
    .dout(new_n634__spl_),
    .din(new_n634_)
  );


  splt
  gnew_n552_
  (
    .dout(new_n552__spl_),
    .din(new_n552_)
  );


  splt
  gnew_n636_
  (
    .dout(new_n636__spl_),
    .din(new_n636_)
  );


  splt
  gnew_n637_
  (
    .dout(new_n637__spl_),
    .din(new_n637_)
  );


  splt
  gnew_n551_
  (
    .dout(new_n551__spl_),
    .din(new_n551_)
  );


  splt
  gnew_n639_
  (
    .dout(new_n639__spl_),
    .din(new_n639_)
  );


  splt
  gnew_n640_
  (
    .dout(new_n640__spl_),
    .din(new_n640_)
  );


  splt
  gG30
  (
    .dout(G30_spl_),
    .din(G30)
  );


  splt
  gG30_spl_
  (
    .dout(G30_spl_0),
    .din(G30_spl_)
  );


  splt
  gG30_spl_0
  (
    .dout(G30_spl_00),
    .din(G30_spl_0)
  );


  splt
  gG30_spl_00
  (
    .dout(G30_spl_000),
    .din(G30_spl_00)
  );


  splt
  gG30_spl_00
  (
    .dout(G30_spl_001),
    .din(G30_spl_00)
  );


  splt
  gG30_spl_0
  (
    .dout(G30_spl_01),
    .din(G30_spl_0)
  );


  splt
  gG30_spl_01
  (
    .dout(G30_spl_010),
    .din(G30_spl_01)
  );


  splt
  gG30_spl_01
  (
    .dout(G30_spl_011),
    .din(G30_spl_01)
  );


  splt
  gG30_spl_
  (
    .dout(G30_spl_1),
    .din(G30_spl_)
  );


  splt
  gG30_spl_1
  (
    .dout(G30_spl_10),
    .din(G30_spl_1)
  );


  splt
  gG30_spl_10
  (
    .dout(G30_spl_100),
    .din(G30_spl_10)
  );


  splt
  gG30_spl_10
  (
    .dout(G30_spl_101),
    .din(G30_spl_10)
  );


  splt
  gG30_spl_1
  (
    .dout(G30_spl_11),
    .din(G30_spl_1)
  );


  splt
  gG30_spl_11
  (
    .dout(G30_spl_110),
    .din(G30_spl_11)
  );


  splt
  gG30_spl_11
  (
    .dout(G30_spl_111),
    .din(G30_spl_11)
  );


  splt
  gG14
  (
    .dout(G14_spl_),
    .din(G14)
  );


  splt
  gG14_spl_
  (
    .dout(G14_spl_0),
    .din(G14_spl_)
  );


  splt
  gG14_spl_0
  (
    .dout(G14_spl_00),
    .din(G14_spl_0)
  );


  splt
  gG14_spl_00
  (
    .dout(G14_spl_000),
    .din(G14_spl_00)
  );


  splt
  gG14_spl_00
  (
    .dout(G14_spl_001),
    .din(G14_spl_00)
  );


  splt
  gG14_spl_0
  (
    .dout(G14_spl_01),
    .din(G14_spl_0)
  );


  splt
  gG14_spl_01
  (
    .dout(G14_spl_010),
    .din(G14_spl_01)
  );


  splt
  gG14_spl_01
  (
    .dout(G14_spl_011),
    .din(G14_spl_01)
  );


  splt
  gG14_spl_
  (
    .dout(G14_spl_1),
    .din(G14_spl_)
  );


  splt
  gG14_spl_1
  (
    .dout(G14_spl_10),
    .din(G14_spl_1)
  );


  splt
  gG14_spl_10
  (
    .dout(G14_spl_100),
    .din(G14_spl_10)
  );


  splt
  gG14_spl_10
  (
    .dout(G14_spl_101),
    .din(G14_spl_10)
  );


  splt
  gG14_spl_1
  (
    .dout(G14_spl_11),
    .din(G14_spl_1)
  );


  splt
  gG14_spl_11
  (
    .dout(G14_spl_110),
    .din(G14_spl_11)
  );


  splt
  gG14_spl_11
  (
    .dout(G14_spl_111),
    .din(G14_spl_11)
  );


  splt
  gnew_n666_
  (
    .dout(new_n666__spl_),
    .din(new_n666_)
  );


  splt
  gnew_n667_
  (
    .dout(new_n667__spl_),
    .din(new_n667_)
  );


  splt
  gnew_n668_
  (
    .dout(new_n668__spl_),
    .din(new_n668_)
  );


  splt
  gnew_n668__spl_
  (
    .dout(new_n668__spl_0),
    .din(new_n668__spl_)
  );


  splt
  gnew_n670_
  (
    .dout(new_n670__spl_),
    .din(new_n670_)
  );


  splt
  gnew_n671_
  (
    .dout(new_n671__spl_),
    .din(new_n671_)
  );


  splt
  gnew_n665_
  (
    .dout(new_n665__spl_),
    .din(new_n665_)
  );


  splt
  gnew_n673_
  (
    .dout(new_n673__spl_),
    .din(new_n673_)
  );


  splt
  gnew_n674_
  (
    .dout(new_n674__spl_),
    .din(new_n674_)
  );


  splt
  gnew_n664_
  (
    .dout(new_n664__spl_),
    .din(new_n664_)
  );


  splt
  gnew_n676_
  (
    .dout(new_n676__spl_),
    .din(new_n676_)
  );


  splt
  gnew_n677_
  (
    .dout(new_n677__spl_),
    .din(new_n677_)
  );


  splt
  gnew_n663_
  (
    .dout(new_n663__spl_),
    .din(new_n663_)
  );


  splt
  gnew_n679_
  (
    .dout(new_n679__spl_),
    .din(new_n679_)
  );


  splt
  gnew_n680_
  (
    .dout(new_n680__spl_),
    .din(new_n680_)
  );


  splt
  gnew_n662_
  (
    .dout(new_n662__spl_),
    .din(new_n662_)
  );


  splt
  gnew_n682_
  (
    .dout(new_n682__spl_),
    .din(new_n682_)
  );


  splt
  gnew_n683_
  (
    .dout(new_n683__spl_),
    .din(new_n683_)
  );


  splt
  gnew_n661_
  (
    .dout(new_n661__spl_),
    .din(new_n661_)
  );


  splt
  gnew_n685_
  (
    .dout(new_n685__spl_),
    .din(new_n685_)
  );


  splt
  gnew_n686_
  (
    .dout(new_n686__spl_),
    .din(new_n686_)
  );


  splt
  gnew_n660_
  (
    .dout(new_n660__spl_),
    .din(new_n660_)
  );


  splt
  gnew_n688_
  (
    .dout(new_n688__spl_),
    .din(new_n688_)
  );


  splt
  gnew_n689_
  (
    .dout(new_n689__spl_),
    .din(new_n689_)
  );


  splt
  gnew_n659_
  (
    .dout(new_n659__spl_),
    .din(new_n659_)
  );


  splt
  gnew_n691_
  (
    .dout(new_n691__spl_),
    .din(new_n691_)
  );


  splt
  gnew_n692_
  (
    .dout(new_n692__spl_),
    .din(new_n692_)
  );


  splt
  gnew_n658_
  (
    .dout(new_n658__spl_),
    .din(new_n658_)
  );


  splt
  gnew_n694_
  (
    .dout(new_n694__spl_),
    .din(new_n694_)
  );


  splt
  gnew_n695_
  (
    .dout(new_n695__spl_),
    .din(new_n695_)
  );


  splt
  gnew_n657_
  (
    .dout(new_n657__spl_),
    .din(new_n657_)
  );


  splt
  gnew_n697_
  (
    .dout(new_n697__spl_),
    .din(new_n697_)
  );


  splt
  gnew_n698_
  (
    .dout(new_n698__spl_),
    .din(new_n698_)
  );


  splt
  gnew_n656_
  (
    .dout(new_n656__spl_),
    .din(new_n656_)
  );


  splt
  gnew_n700_
  (
    .dout(new_n700__spl_),
    .din(new_n700_)
  );


  splt
  gnew_n701_
  (
    .dout(new_n701__spl_),
    .din(new_n701_)
  );


  splt
  gnew_n655_
  (
    .dout(new_n655__spl_),
    .din(new_n655_)
  );


  splt
  gnew_n703_
  (
    .dout(new_n703__spl_),
    .din(new_n703_)
  );


  splt
  gnew_n704_
  (
    .dout(new_n704__spl_),
    .din(new_n704_)
  );


  splt
  gnew_n654_
  (
    .dout(new_n654__spl_),
    .din(new_n654_)
  );


  splt
  gnew_n706_
  (
    .dout(new_n706__spl_),
    .din(new_n706_)
  );


  splt
  gnew_n707_
  (
    .dout(new_n707__spl_),
    .din(new_n707_)
  );


  splt
  gnew_n653_
  (
    .dout(new_n653__spl_),
    .din(new_n653_)
  );


  splt
  gnew_n709_
  (
    .dout(new_n709__spl_),
    .din(new_n709_)
  );


  splt
  gnew_n710_
  (
    .dout(new_n710__spl_),
    .din(new_n710_)
  );


  splt
  gnew_n652_
  (
    .dout(new_n652__spl_),
    .din(new_n652_)
  );


  splt
  gnew_n712_
  (
    .dout(new_n712__spl_),
    .din(new_n712_)
  );


  splt
  gnew_n713_
  (
    .dout(new_n713__spl_),
    .din(new_n713_)
  );


  splt
  gnew_n651_
  (
    .dout(new_n651__spl_),
    .din(new_n651_)
  );


  splt
  gnew_n715_
  (
    .dout(new_n715__spl_),
    .din(new_n715_)
  );


  splt
  gnew_n716_
  (
    .dout(new_n716__spl_),
    .din(new_n716_)
  );


  splt
  gnew_n650_
  (
    .dout(new_n650__spl_),
    .din(new_n650_)
  );


  splt
  gnew_n718_
  (
    .dout(new_n718__spl_),
    .din(new_n718_)
  );


  splt
  gnew_n719_
  (
    .dout(new_n719__spl_),
    .din(new_n719_)
  );


  splt
  gnew_n649_
  (
    .dout(new_n649__spl_),
    .din(new_n649_)
  );


  splt
  gnew_n721_
  (
    .dout(new_n721__spl_),
    .din(new_n721_)
  );


  splt
  gnew_n722_
  (
    .dout(new_n722__spl_),
    .din(new_n722_)
  );


  splt
  gnew_n648_
  (
    .dout(new_n648__spl_),
    .din(new_n648_)
  );


  splt
  gnew_n724_
  (
    .dout(new_n724__spl_),
    .din(new_n724_)
  );


  splt
  gnew_n725_
  (
    .dout(new_n725__spl_),
    .din(new_n725_)
  );


  splt
  gnew_n647_
  (
    .dout(new_n647__spl_),
    .din(new_n647_)
  );


  splt
  gnew_n727_
  (
    .dout(new_n727__spl_),
    .din(new_n727_)
  );


  splt
  gnew_n728_
  (
    .dout(new_n728__spl_),
    .din(new_n728_)
  );


  splt
  gnew_n646_
  (
    .dout(new_n646__spl_),
    .din(new_n646_)
  );


  splt
  gnew_n730_
  (
    .dout(new_n730__spl_),
    .din(new_n730_)
  );


  splt
  gnew_n731_
  (
    .dout(new_n731__spl_),
    .din(new_n731_)
  );


  splt
  gnew_n645_
  (
    .dout(new_n645__spl_),
    .din(new_n645_)
  );


  splt
  gnew_n733_
  (
    .dout(new_n733__spl_),
    .din(new_n733_)
  );


  splt
  gnew_n734_
  (
    .dout(new_n734__spl_),
    .din(new_n734_)
  );


  splt
  gnew_n644_
  (
    .dout(new_n644__spl_),
    .din(new_n644_)
  );


  splt
  gnew_n736_
  (
    .dout(new_n736__spl_),
    .din(new_n736_)
  );


  splt
  gnew_n737_
  (
    .dout(new_n737__spl_),
    .din(new_n737_)
  );


  splt
  gnew_n643_
  (
    .dout(new_n643__spl_),
    .din(new_n643_)
  );


  splt
  gnew_n739_
  (
    .dout(new_n739__spl_),
    .din(new_n739_)
  );


  splt
  gnew_n740_
  (
    .dout(new_n740__spl_),
    .din(new_n740_)
  );


  splt
  gG31
  (
    .dout(G31_spl_),
    .din(G31)
  );


  splt
  gG31_spl_
  (
    .dout(G31_spl_0),
    .din(G31_spl_)
  );


  splt
  gG31_spl_0
  (
    .dout(G31_spl_00),
    .din(G31_spl_0)
  );


  splt
  gG31_spl_00
  (
    .dout(G31_spl_000),
    .din(G31_spl_00)
  );


  splt
  gG31_spl_00
  (
    .dout(G31_spl_001),
    .din(G31_spl_00)
  );


  splt
  gG31_spl_0
  (
    .dout(G31_spl_01),
    .din(G31_spl_0)
  );


  splt
  gG31_spl_01
  (
    .dout(G31_spl_010),
    .din(G31_spl_01)
  );


  splt
  gG31_spl_01
  (
    .dout(G31_spl_011),
    .din(G31_spl_01)
  );


  splt
  gG31_spl_
  (
    .dout(G31_spl_1),
    .din(G31_spl_)
  );


  splt
  gG31_spl_1
  (
    .dout(G31_spl_10),
    .din(G31_spl_1)
  );


  splt
  gG31_spl_10
  (
    .dout(G31_spl_100),
    .din(G31_spl_10)
  );


  splt
  gG31_spl_10
  (
    .dout(G31_spl_101),
    .din(G31_spl_10)
  );


  splt
  gG31_spl_1
  (
    .dout(G31_spl_11),
    .din(G31_spl_1)
  );


  splt
  gG31_spl_11
  (
    .dout(G31_spl_110),
    .din(G31_spl_11)
  );


  splt
  gG31_spl_11
  (
    .dout(G31_spl_111),
    .din(G31_spl_11)
  );


  splt
  gG15
  (
    .dout(G15_spl_),
    .din(G15)
  );


  splt
  gG15_spl_
  (
    .dout(G15_spl_0),
    .din(G15_spl_)
  );


  splt
  gG15_spl_0
  (
    .dout(G15_spl_00),
    .din(G15_spl_0)
  );


  splt
  gG15_spl_00
  (
    .dout(G15_spl_000),
    .din(G15_spl_00)
  );


  splt
  gG15_spl_00
  (
    .dout(G15_spl_001),
    .din(G15_spl_00)
  );


  splt
  gG15_spl_0
  (
    .dout(G15_spl_01),
    .din(G15_spl_0)
  );


  splt
  gG15_spl_01
  (
    .dout(G15_spl_010),
    .din(G15_spl_01)
  );


  splt
  gG15_spl_01
  (
    .dout(G15_spl_011),
    .din(G15_spl_01)
  );


  splt
  gG15_spl_
  (
    .dout(G15_spl_1),
    .din(G15_spl_)
  );


  splt
  gG15_spl_1
  (
    .dout(G15_spl_10),
    .din(G15_spl_1)
  );


  splt
  gG15_spl_10
  (
    .dout(G15_spl_100),
    .din(G15_spl_10)
  );


  splt
  gG15_spl_10
  (
    .dout(G15_spl_101),
    .din(G15_spl_10)
  );


  splt
  gG15_spl_1
  (
    .dout(G15_spl_11),
    .din(G15_spl_1)
  );


  splt
  gG15_spl_11
  (
    .dout(G15_spl_110),
    .din(G15_spl_11)
  );


  splt
  gG15_spl_11
  (
    .dout(G15_spl_111),
    .din(G15_spl_11)
  );


  splt
  gnew_n768_
  (
    .dout(new_n768__spl_),
    .din(new_n768_)
  );


  splt
  gnew_n769_
  (
    .dout(new_n769__spl_),
    .din(new_n769_)
  );


  splt
  gnew_n770_
  (
    .dout(new_n770__spl_),
    .din(new_n770_)
  );


  splt
  gnew_n770__spl_
  (
    .dout(new_n770__spl_0),
    .din(new_n770__spl_)
  );


  splt
  gnew_n772_
  (
    .dout(new_n772__spl_),
    .din(new_n772_)
  );


  splt
  gnew_n773_
  (
    .dout(new_n773__spl_),
    .din(new_n773_)
  );


  splt
  gnew_n767_
  (
    .dout(new_n767__spl_),
    .din(new_n767_)
  );


  splt
  gnew_n775_
  (
    .dout(new_n775__spl_),
    .din(new_n775_)
  );


  splt
  gnew_n776_
  (
    .dout(new_n776__spl_),
    .din(new_n776_)
  );


  splt
  gnew_n766_
  (
    .dout(new_n766__spl_),
    .din(new_n766_)
  );


  splt
  gnew_n778_
  (
    .dout(new_n778__spl_),
    .din(new_n778_)
  );


  splt
  gnew_n779_
  (
    .dout(new_n779__spl_),
    .din(new_n779_)
  );


  splt
  gnew_n765_
  (
    .dout(new_n765__spl_),
    .din(new_n765_)
  );


  splt
  gnew_n781_
  (
    .dout(new_n781__spl_),
    .din(new_n781_)
  );


  splt
  gnew_n782_
  (
    .dout(new_n782__spl_),
    .din(new_n782_)
  );


  splt
  gnew_n764_
  (
    .dout(new_n764__spl_),
    .din(new_n764_)
  );


  splt
  gnew_n784_
  (
    .dout(new_n784__spl_),
    .din(new_n784_)
  );


  splt
  gnew_n785_
  (
    .dout(new_n785__spl_),
    .din(new_n785_)
  );


  splt
  gnew_n763_
  (
    .dout(new_n763__spl_),
    .din(new_n763_)
  );


  splt
  gnew_n787_
  (
    .dout(new_n787__spl_),
    .din(new_n787_)
  );


  splt
  gnew_n788_
  (
    .dout(new_n788__spl_),
    .din(new_n788_)
  );


  splt
  gnew_n762_
  (
    .dout(new_n762__spl_),
    .din(new_n762_)
  );


  splt
  gnew_n790_
  (
    .dout(new_n790__spl_),
    .din(new_n790_)
  );


  splt
  gnew_n791_
  (
    .dout(new_n791__spl_),
    .din(new_n791_)
  );


  splt
  gnew_n761_
  (
    .dout(new_n761__spl_),
    .din(new_n761_)
  );


  splt
  gnew_n793_
  (
    .dout(new_n793__spl_),
    .din(new_n793_)
  );


  splt
  gnew_n794_
  (
    .dout(new_n794__spl_),
    .din(new_n794_)
  );


  splt
  gnew_n760_
  (
    .dout(new_n760__spl_),
    .din(new_n760_)
  );


  splt
  gnew_n796_
  (
    .dout(new_n796__spl_),
    .din(new_n796_)
  );


  splt
  gnew_n797_
  (
    .dout(new_n797__spl_),
    .din(new_n797_)
  );


  splt
  gnew_n759_
  (
    .dout(new_n759__spl_),
    .din(new_n759_)
  );


  splt
  gnew_n799_
  (
    .dout(new_n799__spl_),
    .din(new_n799_)
  );


  splt
  gnew_n800_
  (
    .dout(new_n800__spl_),
    .din(new_n800_)
  );


  splt
  gnew_n758_
  (
    .dout(new_n758__spl_),
    .din(new_n758_)
  );


  splt
  gnew_n802_
  (
    .dout(new_n802__spl_),
    .din(new_n802_)
  );


  splt
  gnew_n803_
  (
    .dout(new_n803__spl_),
    .din(new_n803_)
  );


  splt
  gnew_n757_
  (
    .dout(new_n757__spl_),
    .din(new_n757_)
  );


  splt
  gnew_n805_
  (
    .dout(new_n805__spl_),
    .din(new_n805_)
  );


  splt
  gnew_n806_
  (
    .dout(new_n806__spl_),
    .din(new_n806_)
  );


  splt
  gnew_n756_
  (
    .dout(new_n756__spl_),
    .din(new_n756_)
  );


  splt
  gnew_n808_
  (
    .dout(new_n808__spl_),
    .din(new_n808_)
  );


  splt
  gnew_n809_
  (
    .dout(new_n809__spl_),
    .din(new_n809_)
  );


  splt
  gnew_n755_
  (
    .dout(new_n755__spl_),
    .din(new_n755_)
  );


  splt
  gnew_n811_
  (
    .dout(new_n811__spl_),
    .din(new_n811_)
  );


  splt
  gnew_n812_
  (
    .dout(new_n812__spl_),
    .din(new_n812_)
  );


  splt
  gnew_n754_
  (
    .dout(new_n754__spl_),
    .din(new_n754_)
  );


  splt
  gnew_n814_
  (
    .dout(new_n814__spl_),
    .din(new_n814_)
  );


  splt
  gnew_n815_
  (
    .dout(new_n815__spl_),
    .din(new_n815_)
  );


  splt
  gnew_n753_
  (
    .dout(new_n753__spl_),
    .din(new_n753_)
  );


  splt
  gnew_n817_
  (
    .dout(new_n817__spl_),
    .din(new_n817_)
  );


  splt
  gnew_n818_
  (
    .dout(new_n818__spl_),
    .din(new_n818_)
  );


  splt
  gnew_n752_
  (
    .dout(new_n752__spl_),
    .din(new_n752_)
  );


  splt
  gnew_n820_
  (
    .dout(new_n820__spl_),
    .din(new_n820_)
  );


  splt
  gnew_n821_
  (
    .dout(new_n821__spl_),
    .din(new_n821_)
  );


  splt
  gnew_n751_
  (
    .dout(new_n751__spl_),
    .din(new_n751_)
  );


  splt
  gnew_n823_
  (
    .dout(new_n823__spl_),
    .din(new_n823_)
  );


  splt
  gnew_n824_
  (
    .dout(new_n824__spl_),
    .din(new_n824_)
  );


  splt
  gnew_n750_
  (
    .dout(new_n750__spl_),
    .din(new_n750_)
  );


  splt
  gnew_n826_
  (
    .dout(new_n826__spl_),
    .din(new_n826_)
  );


  splt
  gnew_n827_
  (
    .dout(new_n827__spl_),
    .din(new_n827_)
  );


  splt
  gnew_n749_
  (
    .dout(new_n749__spl_),
    .din(new_n749_)
  );


  splt
  gnew_n829_
  (
    .dout(new_n829__spl_),
    .din(new_n829_)
  );


  splt
  gnew_n830_
  (
    .dout(new_n830__spl_),
    .din(new_n830_)
  );


  splt
  gnew_n748_
  (
    .dout(new_n748__spl_),
    .din(new_n748_)
  );


  splt
  gnew_n832_
  (
    .dout(new_n832__spl_),
    .din(new_n832_)
  );


  splt
  gnew_n833_
  (
    .dout(new_n833__spl_),
    .din(new_n833_)
  );


  splt
  gnew_n747_
  (
    .dout(new_n747__spl_),
    .din(new_n747_)
  );


  splt
  gnew_n835_
  (
    .dout(new_n835__spl_),
    .din(new_n835_)
  );


  splt
  gnew_n836_
  (
    .dout(new_n836__spl_),
    .din(new_n836_)
  );


  splt
  gnew_n746_
  (
    .dout(new_n746__spl_),
    .din(new_n746_)
  );


  splt
  gnew_n838_
  (
    .dout(new_n838__spl_),
    .din(new_n838_)
  );


  splt
  gnew_n839_
  (
    .dout(new_n839__spl_),
    .din(new_n839_)
  );


  splt
  gnew_n745_
  (
    .dout(new_n745__spl_),
    .din(new_n745_)
  );


  splt
  gnew_n841_
  (
    .dout(new_n841__spl_),
    .din(new_n841_)
  );


  splt
  gnew_n842_
  (
    .dout(new_n842__spl_),
    .din(new_n842_)
  );


  splt
  gnew_n744_
  (
    .dout(new_n744__spl_),
    .din(new_n744_)
  );


  splt
  gnew_n844_
  (
    .dout(new_n844__spl_),
    .din(new_n844_)
  );


  splt
  gnew_n845_
  (
    .dout(new_n845__spl_),
    .din(new_n845_)
  );


  splt
  gnew_n743_
  (
    .dout(new_n743__spl_),
    .din(new_n743_)
  );


  splt
  gnew_n847_
  (
    .dout(new_n847__spl_),
    .din(new_n847_)
  );


  splt
  gnew_n848_
  (
    .dout(new_n848__spl_),
    .din(new_n848_)
  );


  splt
  gG32
  (
    .dout(G32_spl_),
    .din(G32)
  );


  splt
  gG32_spl_
  (
    .dout(G32_spl_0),
    .din(G32_spl_)
  );


  splt
  gG32_spl_0
  (
    .dout(G32_spl_00),
    .din(G32_spl_0)
  );


  splt
  gG32_spl_00
  (
    .dout(G32_spl_000),
    .din(G32_spl_00)
  );


  splt
  gG32_spl_00
  (
    .dout(G32_spl_001),
    .din(G32_spl_00)
  );


  splt
  gG32_spl_0
  (
    .dout(G32_spl_01),
    .din(G32_spl_0)
  );


  splt
  gG32_spl_01
  (
    .dout(G32_spl_010),
    .din(G32_spl_01)
  );


  splt
  gG32_spl_01
  (
    .dout(G32_spl_011),
    .din(G32_spl_01)
  );


  splt
  gG32_spl_
  (
    .dout(G32_spl_1),
    .din(G32_spl_)
  );


  splt
  gG32_spl_1
  (
    .dout(G32_spl_10),
    .din(G32_spl_1)
  );


  splt
  gG32_spl_10
  (
    .dout(G32_spl_100),
    .din(G32_spl_10)
  );


  splt
  gG32_spl_10
  (
    .dout(G32_spl_101),
    .din(G32_spl_10)
  );


  splt
  gG32_spl_1
  (
    .dout(G32_spl_11),
    .din(G32_spl_1)
  );


  splt
  gG32_spl_11
  (
    .dout(G32_spl_110),
    .din(G32_spl_11)
  );


  splt
  gG32_spl_11
  (
    .dout(G32_spl_111),
    .din(G32_spl_11)
  );


  splt
  gG16
  (
    .dout(G16_spl_),
    .din(G16)
  );


  splt
  gG16_spl_
  (
    .dout(G16_spl_0),
    .din(G16_spl_)
  );


  splt
  gG16_spl_0
  (
    .dout(G16_spl_00),
    .din(G16_spl_0)
  );


  splt
  gG16_spl_00
  (
    .dout(G16_spl_000),
    .din(G16_spl_00)
  );


  splt
  gG16_spl_00
  (
    .dout(G16_spl_001),
    .din(G16_spl_00)
  );


  splt
  gG16_spl_0
  (
    .dout(G16_spl_01),
    .din(G16_spl_0)
  );


  splt
  gG16_spl_01
  (
    .dout(G16_spl_010),
    .din(G16_spl_01)
  );


  splt
  gG16_spl_01
  (
    .dout(G16_spl_011),
    .din(G16_spl_01)
  );


  splt
  gG16_spl_
  (
    .dout(G16_spl_1),
    .din(G16_spl_)
  );


  splt
  gG16_spl_1
  (
    .dout(G16_spl_10),
    .din(G16_spl_1)
  );


  splt
  gG16_spl_10
  (
    .dout(G16_spl_100),
    .din(G16_spl_10)
  );


  splt
  gG16_spl_10
  (
    .dout(G16_spl_101),
    .din(G16_spl_10)
  );


  splt
  gG16_spl_1
  (
    .dout(G16_spl_11),
    .din(G16_spl_1)
  );


  splt
  gG16_spl_11
  (
    .dout(G16_spl_110),
    .din(G16_spl_11)
  );


  splt
  gG16_spl_11
  (
    .dout(G16_spl_111),
    .din(G16_spl_11)
  );


  splt
  gnew_n878_
  (
    .dout(new_n878__spl_),
    .din(new_n878_)
  );


  splt
  gnew_n879_
  (
    .dout(new_n879__spl_),
    .din(new_n879_)
  );


  splt
  gnew_n880_
  (
    .dout(new_n880__spl_),
    .din(new_n880_)
  );


  splt
  gnew_n882_
  (
    .dout(new_n882__spl_),
    .din(new_n882_)
  );


  splt
  gnew_n883_
  (
    .dout(new_n883__spl_),
    .din(new_n883_)
  );


  splt
  gnew_n877_
  (
    .dout(new_n877__spl_),
    .din(new_n877_)
  );


  splt
  gnew_n885_
  (
    .dout(new_n885__spl_),
    .din(new_n885_)
  );


  splt
  gnew_n886_
  (
    .dout(new_n886__spl_),
    .din(new_n886_)
  );


  splt
  gnew_n876_
  (
    .dout(new_n876__spl_),
    .din(new_n876_)
  );


  splt
  gnew_n888_
  (
    .dout(new_n888__spl_),
    .din(new_n888_)
  );


  splt
  gnew_n889_
  (
    .dout(new_n889__spl_),
    .din(new_n889_)
  );


  splt
  gnew_n875_
  (
    .dout(new_n875__spl_),
    .din(new_n875_)
  );


  splt
  gnew_n891_
  (
    .dout(new_n891__spl_),
    .din(new_n891_)
  );


  splt
  gnew_n892_
  (
    .dout(new_n892__spl_),
    .din(new_n892_)
  );


  splt
  gnew_n874_
  (
    .dout(new_n874__spl_),
    .din(new_n874_)
  );


  splt
  gnew_n894_
  (
    .dout(new_n894__spl_),
    .din(new_n894_)
  );


  splt
  gnew_n895_
  (
    .dout(new_n895__spl_),
    .din(new_n895_)
  );


  splt
  gnew_n873_
  (
    .dout(new_n873__spl_),
    .din(new_n873_)
  );


  splt
  gnew_n897_
  (
    .dout(new_n897__spl_),
    .din(new_n897_)
  );


  splt
  gnew_n898_
  (
    .dout(new_n898__spl_),
    .din(new_n898_)
  );


  splt
  gnew_n872_
  (
    .dout(new_n872__spl_),
    .din(new_n872_)
  );


  splt
  gnew_n900_
  (
    .dout(new_n900__spl_),
    .din(new_n900_)
  );


  splt
  gnew_n901_
  (
    .dout(new_n901__spl_),
    .din(new_n901_)
  );


  splt
  gnew_n871_
  (
    .dout(new_n871__spl_),
    .din(new_n871_)
  );


  splt
  gnew_n903_
  (
    .dout(new_n903__spl_),
    .din(new_n903_)
  );


  splt
  gnew_n904_
  (
    .dout(new_n904__spl_),
    .din(new_n904_)
  );


  splt
  gnew_n870_
  (
    .dout(new_n870__spl_),
    .din(new_n870_)
  );


  splt
  gnew_n906_
  (
    .dout(new_n906__spl_),
    .din(new_n906_)
  );


  splt
  gnew_n907_
  (
    .dout(new_n907__spl_),
    .din(new_n907_)
  );


  splt
  gnew_n869_
  (
    .dout(new_n869__spl_),
    .din(new_n869_)
  );


  splt
  gnew_n909_
  (
    .dout(new_n909__spl_),
    .din(new_n909_)
  );


  splt
  gnew_n910_
  (
    .dout(new_n910__spl_),
    .din(new_n910_)
  );


  splt
  gnew_n868_
  (
    .dout(new_n868__spl_),
    .din(new_n868_)
  );


  splt
  gnew_n912_
  (
    .dout(new_n912__spl_),
    .din(new_n912_)
  );


  splt
  gnew_n913_
  (
    .dout(new_n913__spl_),
    .din(new_n913_)
  );


  splt
  gnew_n867_
  (
    .dout(new_n867__spl_),
    .din(new_n867_)
  );


  splt
  gnew_n915_
  (
    .dout(new_n915__spl_),
    .din(new_n915_)
  );


  splt
  gnew_n916_
  (
    .dout(new_n916__spl_),
    .din(new_n916_)
  );


  splt
  gnew_n866_
  (
    .dout(new_n866__spl_),
    .din(new_n866_)
  );


  splt
  gnew_n918_
  (
    .dout(new_n918__spl_),
    .din(new_n918_)
  );


  splt
  gnew_n919_
  (
    .dout(new_n919__spl_),
    .din(new_n919_)
  );


  splt
  gnew_n865_
  (
    .dout(new_n865__spl_),
    .din(new_n865_)
  );


  splt
  gnew_n921_
  (
    .dout(new_n921__spl_),
    .din(new_n921_)
  );


  splt
  gnew_n922_
  (
    .dout(new_n922__spl_),
    .din(new_n922_)
  );


  splt
  gnew_n864_
  (
    .dout(new_n864__spl_),
    .din(new_n864_)
  );


  splt
  gnew_n924_
  (
    .dout(new_n924__spl_),
    .din(new_n924_)
  );


  splt
  gnew_n925_
  (
    .dout(new_n925__spl_),
    .din(new_n925_)
  );


  splt
  gnew_n863_
  (
    .dout(new_n863__spl_),
    .din(new_n863_)
  );


  splt
  gnew_n927_
  (
    .dout(new_n927__spl_),
    .din(new_n927_)
  );


  splt
  gnew_n928_
  (
    .dout(new_n928__spl_),
    .din(new_n928_)
  );


  splt
  gnew_n862_
  (
    .dout(new_n862__spl_),
    .din(new_n862_)
  );


  splt
  gnew_n930_
  (
    .dout(new_n930__spl_),
    .din(new_n930_)
  );


  splt
  gnew_n931_
  (
    .dout(new_n931__spl_),
    .din(new_n931_)
  );


  splt
  gnew_n861_
  (
    .dout(new_n861__spl_),
    .din(new_n861_)
  );


  splt
  gnew_n933_
  (
    .dout(new_n933__spl_),
    .din(new_n933_)
  );


  splt
  gnew_n934_
  (
    .dout(new_n934__spl_),
    .din(new_n934_)
  );


  splt
  gnew_n860_
  (
    .dout(new_n860__spl_),
    .din(new_n860_)
  );


  splt
  gnew_n936_
  (
    .dout(new_n936__spl_),
    .din(new_n936_)
  );


  splt
  gnew_n937_
  (
    .dout(new_n937__spl_),
    .din(new_n937_)
  );


  splt
  gnew_n859_
  (
    .dout(new_n859__spl_),
    .din(new_n859_)
  );


  splt
  gnew_n939_
  (
    .dout(new_n939__spl_),
    .din(new_n939_)
  );


  splt
  gnew_n940_
  (
    .dout(new_n940__spl_),
    .din(new_n940_)
  );


  splt
  gnew_n858_
  (
    .dout(new_n858__spl_),
    .din(new_n858_)
  );


  splt
  gnew_n942_
  (
    .dout(new_n942__spl_),
    .din(new_n942_)
  );


  splt
  gnew_n943_
  (
    .dout(new_n943__spl_),
    .din(new_n943_)
  );


  splt
  gnew_n857_
  (
    .dout(new_n857__spl_),
    .din(new_n857_)
  );


  splt
  gnew_n945_
  (
    .dout(new_n945__spl_),
    .din(new_n945_)
  );


  splt
  gnew_n946_
  (
    .dout(new_n946__spl_),
    .din(new_n946_)
  );


  splt
  gnew_n856_
  (
    .dout(new_n856__spl_),
    .din(new_n856_)
  );


  splt
  gnew_n948_
  (
    .dout(new_n948__spl_),
    .din(new_n948_)
  );


  splt
  gnew_n949_
  (
    .dout(new_n949__spl_),
    .din(new_n949_)
  );


  splt
  gnew_n855_
  (
    .dout(new_n855__spl_),
    .din(new_n855_)
  );


  splt
  gnew_n951_
  (
    .dout(new_n951__spl_),
    .din(new_n951_)
  );


  splt
  gnew_n952_
  (
    .dout(new_n952__spl_),
    .din(new_n952_)
  );


  splt
  gnew_n854_
  (
    .dout(new_n854__spl_),
    .din(new_n854_)
  );


  splt
  gnew_n954_
  (
    .dout(new_n954__spl_),
    .din(new_n954_)
  );


  splt
  gnew_n955_
  (
    .dout(new_n955__spl_),
    .din(new_n955_)
  );


  splt
  gnew_n853_
  (
    .dout(new_n853__spl_),
    .din(new_n853_)
  );


  splt
  gnew_n957_
  (
    .dout(new_n957__spl_),
    .din(new_n957_)
  );


  splt
  gnew_n958_
  (
    .dout(new_n958__spl_),
    .din(new_n958_)
  );


  splt
  gnew_n852_
  (
    .dout(new_n852__spl_),
    .din(new_n852_)
  );


  splt
  gnew_n960_
  (
    .dout(new_n960__spl_),
    .din(new_n960_)
  );


  splt
  gnew_n961_
  (
    .dout(new_n961__spl_),
    .din(new_n961_)
  );


  splt
  gnew_n851_
  (
    .dout(new_n851__spl_),
    .din(new_n851_)
  );


  splt
  gnew_n963_
  (
    .dout(new_n963__spl_),
    .din(new_n963_)
  );


  splt
  gnew_n964_
  (
    .dout(new_n964__spl_),
    .din(new_n964_)
  );


  splt
  gnew_n994_
  (
    .dout(new_n994__spl_),
    .din(new_n994_)
  );


  splt
  gnew_n995_
  (
    .dout(new_n995__spl_),
    .din(new_n995_)
  );


  splt
  gnew_n996_
  (
    .dout(new_n996__spl_),
    .din(new_n996_)
  );


  splt
  gnew_n997_
  (
    .dout(new_n997__spl_),
    .din(new_n997_)
  );


  splt
  gnew_n993_
  (
    .dout(new_n993__spl_),
    .din(new_n993_)
  );


  splt
  gnew_n999_
  (
    .dout(new_n999__spl_),
    .din(new_n999_)
  );


  splt
  gnew_n1000_
  (
    .dout(new_n1000__spl_),
    .din(new_n1000_)
  );


  splt
  gnew_n992_
  (
    .dout(new_n992__spl_),
    .din(new_n992_)
  );


  splt
  gnew_n1002_
  (
    .dout(new_n1002__spl_),
    .din(new_n1002_)
  );


  splt
  gnew_n1003_
  (
    .dout(new_n1003__spl_),
    .din(new_n1003_)
  );


  splt
  gnew_n991_
  (
    .dout(new_n991__spl_),
    .din(new_n991_)
  );


  splt
  gnew_n1005_
  (
    .dout(new_n1005__spl_),
    .din(new_n1005_)
  );


  splt
  gnew_n1006_
  (
    .dout(new_n1006__spl_),
    .din(new_n1006_)
  );


  splt
  gnew_n990_
  (
    .dout(new_n990__spl_),
    .din(new_n990_)
  );


  splt
  gnew_n1008_
  (
    .dout(new_n1008__spl_),
    .din(new_n1008_)
  );


  splt
  gnew_n1009_
  (
    .dout(new_n1009__spl_),
    .din(new_n1009_)
  );


  splt
  gnew_n989_
  (
    .dout(new_n989__spl_),
    .din(new_n989_)
  );


  splt
  gnew_n1011_
  (
    .dout(new_n1011__spl_),
    .din(new_n1011_)
  );


  splt
  gnew_n1012_
  (
    .dout(new_n1012__spl_),
    .din(new_n1012_)
  );


  splt
  gnew_n988_
  (
    .dout(new_n988__spl_),
    .din(new_n988_)
  );


  splt
  gnew_n1014_
  (
    .dout(new_n1014__spl_),
    .din(new_n1014_)
  );


  splt
  gnew_n1015_
  (
    .dout(new_n1015__spl_),
    .din(new_n1015_)
  );


  splt
  gnew_n987_
  (
    .dout(new_n987__spl_),
    .din(new_n987_)
  );


  splt
  gnew_n1017_
  (
    .dout(new_n1017__spl_),
    .din(new_n1017_)
  );


  splt
  gnew_n1018_
  (
    .dout(new_n1018__spl_),
    .din(new_n1018_)
  );


  splt
  gnew_n986_
  (
    .dout(new_n986__spl_),
    .din(new_n986_)
  );


  splt
  gnew_n1020_
  (
    .dout(new_n1020__spl_),
    .din(new_n1020_)
  );


  splt
  gnew_n1021_
  (
    .dout(new_n1021__spl_),
    .din(new_n1021_)
  );


  splt
  gnew_n985_
  (
    .dout(new_n985__spl_),
    .din(new_n985_)
  );


  splt
  gnew_n1023_
  (
    .dout(new_n1023__spl_),
    .din(new_n1023_)
  );


  splt
  gnew_n1024_
  (
    .dout(new_n1024__spl_),
    .din(new_n1024_)
  );


  splt
  gnew_n984_
  (
    .dout(new_n984__spl_),
    .din(new_n984_)
  );


  splt
  gnew_n1026_
  (
    .dout(new_n1026__spl_),
    .din(new_n1026_)
  );


  splt
  gnew_n1027_
  (
    .dout(new_n1027__spl_),
    .din(new_n1027_)
  );


  splt
  gnew_n983_
  (
    .dout(new_n983__spl_),
    .din(new_n983_)
  );


  splt
  gnew_n1029_
  (
    .dout(new_n1029__spl_),
    .din(new_n1029_)
  );


  splt
  gnew_n1030_
  (
    .dout(new_n1030__spl_),
    .din(new_n1030_)
  );


  splt
  gnew_n982_
  (
    .dout(new_n982__spl_),
    .din(new_n982_)
  );


  splt
  gnew_n1032_
  (
    .dout(new_n1032__spl_),
    .din(new_n1032_)
  );


  splt
  gnew_n1033_
  (
    .dout(new_n1033__spl_),
    .din(new_n1033_)
  );


  splt
  gnew_n981_
  (
    .dout(new_n981__spl_),
    .din(new_n981_)
  );


  splt
  gnew_n1035_
  (
    .dout(new_n1035__spl_),
    .din(new_n1035_)
  );


  splt
  gnew_n1036_
  (
    .dout(new_n1036__spl_),
    .din(new_n1036_)
  );


  splt
  gnew_n980_
  (
    .dout(new_n980__spl_),
    .din(new_n980_)
  );


  splt
  gnew_n1038_
  (
    .dout(new_n1038__spl_),
    .din(new_n1038_)
  );


  splt
  gnew_n1039_
  (
    .dout(new_n1039__spl_),
    .din(new_n1039_)
  );


  splt
  gnew_n979_
  (
    .dout(new_n979__spl_),
    .din(new_n979_)
  );


  splt
  gnew_n1041_
  (
    .dout(new_n1041__spl_),
    .din(new_n1041_)
  );


  splt
  gnew_n1042_
  (
    .dout(new_n1042__spl_),
    .din(new_n1042_)
  );


  splt
  gnew_n978_
  (
    .dout(new_n978__spl_),
    .din(new_n978_)
  );


  splt
  gnew_n1044_
  (
    .dout(new_n1044__spl_),
    .din(new_n1044_)
  );


  splt
  gnew_n1045_
  (
    .dout(new_n1045__spl_),
    .din(new_n1045_)
  );


  splt
  gnew_n977_
  (
    .dout(new_n977__spl_),
    .din(new_n977_)
  );


  splt
  gnew_n1047_
  (
    .dout(new_n1047__spl_),
    .din(new_n1047_)
  );


  splt
  gnew_n1048_
  (
    .dout(new_n1048__spl_),
    .din(new_n1048_)
  );


  splt
  gnew_n976_
  (
    .dout(new_n976__spl_),
    .din(new_n976_)
  );


  splt
  gnew_n1050_
  (
    .dout(new_n1050__spl_),
    .din(new_n1050_)
  );


  splt
  gnew_n1051_
  (
    .dout(new_n1051__spl_),
    .din(new_n1051_)
  );


  splt
  gnew_n975_
  (
    .dout(new_n975__spl_),
    .din(new_n975_)
  );


  splt
  gnew_n1053_
  (
    .dout(new_n1053__spl_),
    .din(new_n1053_)
  );


  splt
  gnew_n1054_
  (
    .dout(new_n1054__spl_),
    .din(new_n1054_)
  );


  splt
  gnew_n974_
  (
    .dout(new_n974__spl_),
    .din(new_n974_)
  );


  splt
  gnew_n1056_
  (
    .dout(new_n1056__spl_),
    .din(new_n1056_)
  );


  splt
  gnew_n1057_
  (
    .dout(new_n1057__spl_),
    .din(new_n1057_)
  );


  splt
  gnew_n973_
  (
    .dout(new_n973__spl_),
    .din(new_n973_)
  );


  splt
  gnew_n1059_
  (
    .dout(new_n1059__spl_),
    .din(new_n1059_)
  );


  splt
  gnew_n1060_
  (
    .dout(new_n1060__spl_),
    .din(new_n1060_)
  );


  splt
  gnew_n972_
  (
    .dout(new_n972__spl_),
    .din(new_n972_)
  );


  splt
  gnew_n1062_
  (
    .dout(new_n1062__spl_),
    .din(new_n1062_)
  );


  splt
  gnew_n1063_
  (
    .dout(new_n1063__spl_),
    .din(new_n1063_)
  );


  splt
  gnew_n971_
  (
    .dout(new_n971__spl_),
    .din(new_n971_)
  );


  splt
  gnew_n1065_
  (
    .dout(new_n1065__spl_),
    .din(new_n1065_)
  );


  splt
  gnew_n1066_
  (
    .dout(new_n1066__spl_),
    .din(new_n1066_)
  );


  splt
  gnew_n970_
  (
    .dout(new_n970__spl_),
    .din(new_n970_)
  );


  splt
  gnew_n1068_
  (
    .dout(new_n1068__spl_),
    .din(new_n1068_)
  );


  splt
  gnew_n1069_
  (
    .dout(new_n1069__spl_),
    .din(new_n1069_)
  );


  splt
  gnew_n969_
  (
    .dout(new_n969__spl_),
    .din(new_n969_)
  );


  splt
  gnew_n1071_
  (
    .dout(new_n1071__spl_),
    .din(new_n1071_)
  );


  splt
  gnew_n1072_
  (
    .dout(new_n1072__spl_),
    .din(new_n1072_)
  );


  splt
  gnew_n968_
  (
    .dout(new_n968__spl_),
    .din(new_n968_)
  );


  splt
  gnew_n1074_
  (
    .dout(new_n1074__spl_),
    .din(new_n1074_)
  );


  splt
  gnew_n1075_
  (
    .dout(new_n1075__spl_),
    .din(new_n1075_)
  );


  splt
  gnew_n967_
  (
    .dout(new_n967__spl_),
    .din(new_n967_)
  );


  splt
  gnew_n1077_
  (
    .dout(new_n1077__spl_),
    .din(new_n1077_)
  );


  splt
  gnew_n1079_
  (
    .dout(new_n1079__spl_),
    .din(new_n1079_)
  );


  splt
  gnew_n1079__spl_
  (
    .dout(new_n1079__spl_0),
    .din(new_n1079__spl_)
  );


  splt
  gnew_n1107_
  (
    .dout(new_n1107__spl_),
    .din(new_n1107_)
  );


  splt
  gnew_n1108_
  (
    .dout(new_n1108__spl_),
    .din(new_n1108_)
  );


  splt
  gnew_n1109_
  (
    .dout(new_n1109__spl_),
    .din(new_n1109_)
  );


  splt
  gnew_n1106_
  (
    .dout(new_n1106__spl_),
    .din(new_n1106_)
  );


  splt
  gnew_n1111_
  (
    .dout(new_n1111__spl_),
    .din(new_n1111_)
  );


  splt
  gnew_n1112_
  (
    .dout(new_n1112__spl_),
    .din(new_n1112_)
  );


  splt
  gnew_n1105_
  (
    .dout(new_n1105__spl_),
    .din(new_n1105_)
  );


  splt
  gnew_n1114_
  (
    .dout(new_n1114__spl_),
    .din(new_n1114_)
  );


  splt
  gnew_n1115_
  (
    .dout(new_n1115__spl_),
    .din(new_n1115_)
  );


  splt
  gnew_n1104_
  (
    .dout(new_n1104__spl_),
    .din(new_n1104_)
  );


  splt
  gnew_n1117_
  (
    .dout(new_n1117__spl_),
    .din(new_n1117_)
  );


  splt
  gnew_n1118_
  (
    .dout(new_n1118__spl_),
    .din(new_n1118_)
  );


  splt
  gnew_n1103_
  (
    .dout(new_n1103__spl_),
    .din(new_n1103_)
  );


  splt
  gnew_n1120_
  (
    .dout(new_n1120__spl_),
    .din(new_n1120_)
  );


  splt
  gnew_n1121_
  (
    .dout(new_n1121__spl_),
    .din(new_n1121_)
  );


  splt
  gnew_n1102_
  (
    .dout(new_n1102__spl_),
    .din(new_n1102_)
  );


  splt
  gnew_n1123_
  (
    .dout(new_n1123__spl_),
    .din(new_n1123_)
  );


  splt
  gnew_n1124_
  (
    .dout(new_n1124__spl_),
    .din(new_n1124_)
  );


  splt
  gnew_n1101_
  (
    .dout(new_n1101__spl_),
    .din(new_n1101_)
  );


  splt
  gnew_n1126_
  (
    .dout(new_n1126__spl_),
    .din(new_n1126_)
  );


  splt
  gnew_n1127_
  (
    .dout(new_n1127__spl_),
    .din(new_n1127_)
  );


  splt
  gnew_n1100_
  (
    .dout(new_n1100__spl_),
    .din(new_n1100_)
  );


  splt
  gnew_n1129_
  (
    .dout(new_n1129__spl_),
    .din(new_n1129_)
  );


  splt
  gnew_n1130_
  (
    .dout(new_n1130__spl_),
    .din(new_n1130_)
  );


  splt
  gnew_n1099_
  (
    .dout(new_n1099__spl_),
    .din(new_n1099_)
  );


  splt
  gnew_n1132_
  (
    .dout(new_n1132__spl_),
    .din(new_n1132_)
  );


  splt
  gnew_n1133_
  (
    .dout(new_n1133__spl_),
    .din(new_n1133_)
  );


  splt
  gnew_n1098_
  (
    .dout(new_n1098__spl_),
    .din(new_n1098_)
  );


  splt
  gnew_n1135_
  (
    .dout(new_n1135__spl_),
    .din(new_n1135_)
  );


  splt
  gnew_n1136_
  (
    .dout(new_n1136__spl_),
    .din(new_n1136_)
  );


  splt
  gnew_n1097_
  (
    .dout(new_n1097__spl_),
    .din(new_n1097_)
  );


  splt
  gnew_n1138_
  (
    .dout(new_n1138__spl_),
    .din(new_n1138_)
  );


  splt
  gnew_n1139_
  (
    .dout(new_n1139__spl_),
    .din(new_n1139_)
  );


  splt
  gnew_n1096_
  (
    .dout(new_n1096__spl_),
    .din(new_n1096_)
  );


  splt
  gnew_n1141_
  (
    .dout(new_n1141__spl_),
    .din(new_n1141_)
  );


  splt
  gnew_n1142_
  (
    .dout(new_n1142__spl_),
    .din(new_n1142_)
  );


  splt
  gnew_n1095_
  (
    .dout(new_n1095__spl_),
    .din(new_n1095_)
  );


  splt
  gnew_n1144_
  (
    .dout(new_n1144__spl_),
    .din(new_n1144_)
  );


  splt
  gnew_n1145_
  (
    .dout(new_n1145__spl_),
    .din(new_n1145_)
  );


  splt
  gnew_n1094_
  (
    .dout(new_n1094__spl_),
    .din(new_n1094_)
  );


  splt
  gnew_n1147_
  (
    .dout(new_n1147__spl_),
    .din(new_n1147_)
  );


  splt
  gnew_n1148_
  (
    .dout(new_n1148__spl_),
    .din(new_n1148_)
  );


  splt
  gnew_n1093_
  (
    .dout(new_n1093__spl_),
    .din(new_n1093_)
  );


  splt
  gnew_n1150_
  (
    .dout(new_n1150__spl_),
    .din(new_n1150_)
  );


  splt
  gnew_n1151_
  (
    .dout(new_n1151__spl_),
    .din(new_n1151_)
  );


  splt
  gnew_n1092_
  (
    .dout(new_n1092__spl_),
    .din(new_n1092_)
  );


  splt
  gnew_n1153_
  (
    .dout(new_n1153__spl_),
    .din(new_n1153_)
  );


  splt
  gnew_n1154_
  (
    .dout(new_n1154__spl_),
    .din(new_n1154_)
  );


  splt
  gnew_n1091_
  (
    .dout(new_n1091__spl_),
    .din(new_n1091_)
  );


  splt
  gnew_n1156_
  (
    .dout(new_n1156__spl_),
    .din(new_n1156_)
  );


  splt
  gnew_n1157_
  (
    .dout(new_n1157__spl_),
    .din(new_n1157_)
  );


  splt
  gnew_n1090_
  (
    .dout(new_n1090__spl_),
    .din(new_n1090_)
  );


  splt
  gnew_n1159_
  (
    .dout(new_n1159__spl_),
    .din(new_n1159_)
  );


  splt
  gnew_n1160_
  (
    .dout(new_n1160__spl_),
    .din(new_n1160_)
  );


  splt
  gnew_n1089_
  (
    .dout(new_n1089__spl_),
    .din(new_n1089_)
  );


  splt
  gnew_n1162_
  (
    .dout(new_n1162__spl_),
    .din(new_n1162_)
  );


  splt
  gnew_n1163_
  (
    .dout(new_n1163__spl_),
    .din(new_n1163_)
  );


  splt
  gnew_n1088_
  (
    .dout(new_n1088__spl_),
    .din(new_n1088_)
  );


  splt
  gnew_n1165_
  (
    .dout(new_n1165__spl_),
    .din(new_n1165_)
  );


  splt
  gnew_n1166_
  (
    .dout(new_n1166__spl_),
    .din(new_n1166_)
  );


  splt
  gnew_n1087_
  (
    .dout(new_n1087__spl_),
    .din(new_n1087_)
  );


  splt
  gnew_n1168_
  (
    .dout(new_n1168__spl_),
    .din(new_n1168_)
  );


  splt
  gnew_n1169_
  (
    .dout(new_n1169__spl_),
    .din(new_n1169_)
  );


  splt
  gnew_n1086_
  (
    .dout(new_n1086__spl_),
    .din(new_n1086_)
  );


  splt
  gnew_n1171_
  (
    .dout(new_n1171__spl_),
    .din(new_n1171_)
  );


  splt
  gnew_n1172_
  (
    .dout(new_n1172__spl_),
    .din(new_n1172_)
  );


  splt
  gnew_n1085_
  (
    .dout(new_n1085__spl_),
    .din(new_n1085_)
  );


  splt
  gnew_n1174_
  (
    .dout(new_n1174__spl_),
    .din(new_n1174_)
  );


  splt
  gnew_n1175_
  (
    .dout(new_n1175__spl_),
    .din(new_n1175_)
  );


  splt
  gnew_n1084_
  (
    .dout(new_n1084__spl_),
    .din(new_n1084_)
  );


  splt
  gnew_n1177_
  (
    .dout(new_n1177__spl_),
    .din(new_n1177_)
  );


  splt
  gnew_n1178_
  (
    .dout(new_n1178__spl_),
    .din(new_n1178_)
  );


  splt
  gnew_n1083_
  (
    .dout(new_n1083__spl_),
    .din(new_n1083_)
  );


  splt
  gnew_n1180_
  (
    .dout(new_n1180__spl_),
    .din(new_n1180_)
  );


  splt
  gnew_n1181_
  (
    .dout(new_n1181__spl_),
    .din(new_n1181_)
  );


  splt
  gnew_n1082_
  (
    .dout(new_n1082__spl_),
    .din(new_n1082_)
  );


  splt
  gnew_n1183_
  (
    .dout(new_n1183__spl_),
    .din(new_n1183_)
  );


  splt
  gnew_n1184_
  (
    .dout(new_n1184__spl_),
    .din(new_n1184_)
  );


  splt
  gnew_n1081_
  (
    .dout(new_n1081__spl_),
    .din(new_n1081_)
  );


  splt
  gnew_n1186_
  (
    .dout(new_n1186__spl_),
    .din(new_n1186_)
  );


  splt
  gnew_n1187_
  (
    .dout(new_n1187__spl_),
    .din(new_n1187_)
  );


  splt
  gnew_n1189_
  (
    .dout(new_n1189__spl_),
    .din(new_n1189_)
  );


  splt
  gnew_n1190_
  (
    .dout(new_n1190__spl_),
    .din(new_n1190_)
  );


  splt
  gnew_n1218_
  (
    .dout(new_n1218__spl_),
    .din(new_n1218_)
  );


  splt
  gnew_n1219_
  (
    .dout(new_n1219__spl_),
    .din(new_n1219_)
  );


  splt
  gnew_n1220_
  (
    .dout(new_n1220__spl_),
    .din(new_n1220_)
  );


  splt
  gnew_n1217_
  (
    .dout(new_n1217__spl_),
    .din(new_n1217_)
  );


  splt
  gnew_n1222_
  (
    .dout(new_n1222__spl_),
    .din(new_n1222_)
  );


  splt
  gnew_n1223_
  (
    .dout(new_n1223__spl_),
    .din(new_n1223_)
  );


  splt
  gnew_n1216_
  (
    .dout(new_n1216__spl_),
    .din(new_n1216_)
  );


  splt
  gnew_n1225_
  (
    .dout(new_n1225__spl_),
    .din(new_n1225_)
  );


  splt
  gnew_n1226_
  (
    .dout(new_n1226__spl_),
    .din(new_n1226_)
  );


  splt
  gnew_n1215_
  (
    .dout(new_n1215__spl_),
    .din(new_n1215_)
  );


  splt
  gnew_n1228_
  (
    .dout(new_n1228__spl_),
    .din(new_n1228_)
  );


  splt
  gnew_n1229_
  (
    .dout(new_n1229__spl_),
    .din(new_n1229_)
  );


  splt
  gnew_n1214_
  (
    .dout(new_n1214__spl_),
    .din(new_n1214_)
  );


  splt
  gnew_n1231_
  (
    .dout(new_n1231__spl_),
    .din(new_n1231_)
  );


  splt
  gnew_n1232_
  (
    .dout(new_n1232__spl_),
    .din(new_n1232_)
  );


  splt
  gnew_n1213_
  (
    .dout(new_n1213__spl_),
    .din(new_n1213_)
  );


  splt
  gnew_n1234_
  (
    .dout(new_n1234__spl_),
    .din(new_n1234_)
  );


  splt
  gnew_n1235_
  (
    .dout(new_n1235__spl_),
    .din(new_n1235_)
  );


  splt
  gnew_n1212_
  (
    .dout(new_n1212__spl_),
    .din(new_n1212_)
  );


  splt
  gnew_n1237_
  (
    .dout(new_n1237__spl_),
    .din(new_n1237_)
  );


  splt
  gnew_n1238_
  (
    .dout(new_n1238__spl_),
    .din(new_n1238_)
  );


  splt
  gnew_n1211_
  (
    .dout(new_n1211__spl_),
    .din(new_n1211_)
  );


  splt
  gnew_n1240_
  (
    .dout(new_n1240__spl_),
    .din(new_n1240_)
  );


  splt
  gnew_n1241_
  (
    .dout(new_n1241__spl_),
    .din(new_n1241_)
  );


  splt
  gnew_n1210_
  (
    .dout(new_n1210__spl_),
    .din(new_n1210_)
  );


  splt
  gnew_n1243_
  (
    .dout(new_n1243__spl_),
    .din(new_n1243_)
  );


  splt
  gnew_n1244_
  (
    .dout(new_n1244__spl_),
    .din(new_n1244_)
  );


  splt
  gnew_n1209_
  (
    .dout(new_n1209__spl_),
    .din(new_n1209_)
  );


  splt
  gnew_n1246_
  (
    .dout(new_n1246__spl_),
    .din(new_n1246_)
  );


  splt
  gnew_n1247_
  (
    .dout(new_n1247__spl_),
    .din(new_n1247_)
  );


  splt
  gnew_n1208_
  (
    .dout(new_n1208__spl_),
    .din(new_n1208_)
  );


  splt
  gnew_n1249_
  (
    .dout(new_n1249__spl_),
    .din(new_n1249_)
  );


  splt
  gnew_n1250_
  (
    .dout(new_n1250__spl_),
    .din(new_n1250_)
  );


  splt
  gnew_n1207_
  (
    .dout(new_n1207__spl_),
    .din(new_n1207_)
  );


  splt
  gnew_n1252_
  (
    .dout(new_n1252__spl_),
    .din(new_n1252_)
  );


  splt
  gnew_n1253_
  (
    .dout(new_n1253__spl_),
    .din(new_n1253_)
  );


  splt
  gnew_n1206_
  (
    .dout(new_n1206__spl_),
    .din(new_n1206_)
  );


  splt
  gnew_n1255_
  (
    .dout(new_n1255__spl_),
    .din(new_n1255_)
  );


  splt
  gnew_n1256_
  (
    .dout(new_n1256__spl_),
    .din(new_n1256_)
  );


  splt
  gnew_n1205_
  (
    .dout(new_n1205__spl_),
    .din(new_n1205_)
  );


  splt
  gnew_n1258_
  (
    .dout(new_n1258__spl_),
    .din(new_n1258_)
  );


  splt
  gnew_n1259_
  (
    .dout(new_n1259__spl_),
    .din(new_n1259_)
  );


  splt
  gnew_n1204_
  (
    .dout(new_n1204__spl_),
    .din(new_n1204_)
  );


  splt
  gnew_n1261_
  (
    .dout(new_n1261__spl_),
    .din(new_n1261_)
  );


  splt
  gnew_n1262_
  (
    .dout(new_n1262__spl_),
    .din(new_n1262_)
  );


  splt
  gnew_n1203_
  (
    .dout(new_n1203__spl_),
    .din(new_n1203_)
  );


  splt
  gnew_n1264_
  (
    .dout(new_n1264__spl_),
    .din(new_n1264_)
  );


  splt
  gnew_n1265_
  (
    .dout(new_n1265__spl_),
    .din(new_n1265_)
  );


  splt
  gnew_n1202_
  (
    .dout(new_n1202__spl_),
    .din(new_n1202_)
  );


  splt
  gnew_n1267_
  (
    .dout(new_n1267__spl_),
    .din(new_n1267_)
  );


  splt
  gnew_n1268_
  (
    .dout(new_n1268__spl_),
    .din(new_n1268_)
  );


  splt
  gnew_n1201_
  (
    .dout(new_n1201__spl_),
    .din(new_n1201_)
  );


  splt
  gnew_n1270_
  (
    .dout(new_n1270__spl_),
    .din(new_n1270_)
  );


  splt
  gnew_n1271_
  (
    .dout(new_n1271__spl_),
    .din(new_n1271_)
  );


  splt
  gnew_n1200_
  (
    .dout(new_n1200__spl_),
    .din(new_n1200_)
  );


  splt
  gnew_n1273_
  (
    .dout(new_n1273__spl_),
    .din(new_n1273_)
  );


  splt
  gnew_n1274_
  (
    .dout(new_n1274__spl_),
    .din(new_n1274_)
  );


  splt
  gnew_n1199_
  (
    .dout(new_n1199__spl_),
    .din(new_n1199_)
  );


  splt
  gnew_n1276_
  (
    .dout(new_n1276__spl_),
    .din(new_n1276_)
  );


  splt
  gnew_n1277_
  (
    .dout(new_n1277__spl_),
    .din(new_n1277_)
  );


  splt
  gnew_n1198_
  (
    .dout(new_n1198__spl_),
    .din(new_n1198_)
  );


  splt
  gnew_n1279_
  (
    .dout(new_n1279__spl_),
    .din(new_n1279_)
  );


  splt
  gnew_n1280_
  (
    .dout(new_n1280__spl_),
    .din(new_n1280_)
  );


  splt
  gnew_n1197_
  (
    .dout(new_n1197__spl_),
    .din(new_n1197_)
  );


  splt
  gnew_n1282_
  (
    .dout(new_n1282__spl_),
    .din(new_n1282_)
  );


  splt
  gnew_n1283_
  (
    .dout(new_n1283__spl_),
    .din(new_n1283_)
  );


  splt
  gnew_n1196_
  (
    .dout(new_n1196__spl_),
    .din(new_n1196_)
  );


  splt
  gnew_n1285_
  (
    .dout(new_n1285__spl_),
    .din(new_n1285_)
  );


  splt
  gnew_n1286_
  (
    .dout(new_n1286__spl_),
    .din(new_n1286_)
  );


  splt
  gnew_n1195_
  (
    .dout(new_n1195__spl_),
    .din(new_n1195_)
  );


  splt
  gnew_n1288_
  (
    .dout(new_n1288__spl_),
    .din(new_n1288_)
  );


  splt
  gnew_n1289_
  (
    .dout(new_n1289__spl_),
    .din(new_n1289_)
  );


  splt
  gnew_n1194_
  (
    .dout(new_n1194__spl_),
    .din(new_n1194_)
  );


  splt
  gnew_n1291_
  (
    .dout(new_n1291__spl_),
    .din(new_n1291_)
  );


  splt
  gnew_n1292_
  (
    .dout(new_n1292__spl_),
    .din(new_n1292_)
  );


  splt
  gnew_n1193_
  (
    .dout(new_n1193__spl_),
    .din(new_n1193_)
  );


  splt
  gnew_n1294_
  (
    .dout(new_n1294__spl_),
    .din(new_n1294_)
  );


  splt
  gnew_n1295_
  (
    .dout(new_n1295__spl_),
    .din(new_n1295_)
  );


  splt
  gnew_n1321_
  (
    .dout(new_n1321__spl_),
    .din(new_n1321_)
  );


  splt
  gnew_n1322_
  (
    .dout(new_n1322__spl_),
    .din(new_n1322_)
  );


  splt
  gnew_n1323_
  (
    .dout(new_n1323__spl_),
    .din(new_n1323_)
  );


  splt
  gnew_n1320_
  (
    .dout(new_n1320__spl_),
    .din(new_n1320_)
  );


  splt
  gnew_n1325_
  (
    .dout(new_n1325__spl_),
    .din(new_n1325_)
  );


  splt
  gnew_n1326_
  (
    .dout(new_n1326__spl_),
    .din(new_n1326_)
  );


  splt
  gnew_n1319_
  (
    .dout(new_n1319__spl_),
    .din(new_n1319_)
  );


  splt
  gnew_n1328_
  (
    .dout(new_n1328__spl_),
    .din(new_n1328_)
  );


  splt
  gnew_n1329_
  (
    .dout(new_n1329__spl_),
    .din(new_n1329_)
  );


  splt
  gnew_n1318_
  (
    .dout(new_n1318__spl_),
    .din(new_n1318_)
  );


  splt
  gnew_n1331_
  (
    .dout(new_n1331__spl_),
    .din(new_n1331_)
  );


  splt
  gnew_n1332_
  (
    .dout(new_n1332__spl_),
    .din(new_n1332_)
  );


  splt
  gnew_n1317_
  (
    .dout(new_n1317__spl_),
    .din(new_n1317_)
  );


  splt
  gnew_n1334_
  (
    .dout(new_n1334__spl_),
    .din(new_n1334_)
  );


  splt
  gnew_n1335_
  (
    .dout(new_n1335__spl_),
    .din(new_n1335_)
  );


  splt
  gnew_n1316_
  (
    .dout(new_n1316__spl_),
    .din(new_n1316_)
  );


  splt
  gnew_n1337_
  (
    .dout(new_n1337__spl_),
    .din(new_n1337_)
  );


  splt
  gnew_n1338_
  (
    .dout(new_n1338__spl_),
    .din(new_n1338_)
  );


  splt
  gnew_n1315_
  (
    .dout(new_n1315__spl_),
    .din(new_n1315_)
  );


  splt
  gnew_n1340_
  (
    .dout(new_n1340__spl_),
    .din(new_n1340_)
  );


  splt
  gnew_n1341_
  (
    .dout(new_n1341__spl_),
    .din(new_n1341_)
  );


  splt
  gnew_n1314_
  (
    .dout(new_n1314__spl_),
    .din(new_n1314_)
  );


  splt
  gnew_n1343_
  (
    .dout(new_n1343__spl_),
    .din(new_n1343_)
  );


  splt
  gnew_n1344_
  (
    .dout(new_n1344__spl_),
    .din(new_n1344_)
  );


  splt
  gnew_n1313_
  (
    .dout(new_n1313__spl_),
    .din(new_n1313_)
  );


  splt
  gnew_n1346_
  (
    .dout(new_n1346__spl_),
    .din(new_n1346_)
  );


  splt
  gnew_n1347_
  (
    .dout(new_n1347__spl_),
    .din(new_n1347_)
  );


  splt
  gnew_n1312_
  (
    .dout(new_n1312__spl_),
    .din(new_n1312_)
  );


  splt
  gnew_n1349_
  (
    .dout(new_n1349__spl_),
    .din(new_n1349_)
  );


  splt
  gnew_n1350_
  (
    .dout(new_n1350__spl_),
    .din(new_n1350_)
  );


  splt
  gnew_n1311_
  (
    .dout(new_n1311__spl_),
    .din(new_n1311_)
  );


  splt
  gnew_n1352_
  (
    .dout(new_n1352__spl_),
    .din(new_n1352_)
  );


  splt
  gnew_n1353_
  (
    .dout(new_n1353__spl_),
    .din(new_n1353_)
  );


  splt
  gnew_n1310_
  (
    .dout(new_n1310__spl_),
    .din(new_n1310_)
  );


  splt
  gnew_n1355_
  (
    .dout(new_n1355__spl_),
    .din(new_n1355_)
  );


  splt
  gnew_n1356_
  (
    .dout(new_n1356__spl_),
    .din(new_n1356_)
  );


  splt
  gnew_n1309_
  (
    .dout(new_n1309__spl_),
    .din(new_n1309_)
  );


  splt
  gnew_n1358_
  (
    .dout(new_n1358__spl_),
    .din(new_n1358_)
  );


  splt
  gnew_n1359_
  (
    .dout(new_n1359__spl_),
    .din(new_n1359_)
  );


  splt
  gnew_n1308_
  (
    .dout(new_n1308__spl_),
    .din(new_n1308_)
  );


  splt
  gnew_n1361_
  (
    .dout(new_n1361__spl_),
    .din(new_n1361_)
  );


  splt
  gnew_n1362_
  (
    .dout(new_n1362__spl_),
    .din(new_n1362_)
  );


  splt
  gnew_n1307_
  (
    .dout(new_n1307__spl_),
    .din(new_n1307_)
  );


  splt
  gnew_n1364_
  (
    .dout(new_n1364__spl_),
    .din(new_n1364_)
  );


  splt
  gnew_n1365_
  (
    .dout(new_n1365__spl_),
    .din(new_n1365_)
  );


  splt
  gnew_n1306_
  (
    .dout(new_n1306__spl_),
    .din(new_n1306_)
  );


  splt
  gnew_n1367_
  (
    .dout(new_n1367__spl_),
    .din(new_n1367_)
  );


  splt
  gnew_n1368_
  (
    .dout(new_n1368__spl_),
    .din(new_n1368_)
  );


  splt
  gnew_n1305_
  (
    .dout(new_n1305__spl_),
    .din(new_n1305_)
  );


  splt
  gnew_n1370_
  (
    .dout(new_n1370__spl_),
    .din(new_n1370_)
  );


  splt
  gnew_n1371_
  (
    .dout(new_n1371__spl_),
    .din(new_n1371_)
  );


  splt
  gnew_n1304_
  (
    .dout(new_n1304__spl_),
    .din(new_n1304_)
  );


  splt
  gnew_n1373_
  (
    .dout(new_n1373__spl_),
    .din(new_n1373_)
  );


  splt
  gnew_n1374_
  (
    .dout(new_n1374__spl_),
    .din(new_n1374_)
  );


  splt
  gnew_n1303_
  (
    .dout(new_n1303__spl_),
    .din(new_n1303_)
  );


  splt
  gnew_n1376_
  (
    .dout(new_n1376__spl_),
    .din(new_n1376_)
  );


  splt
  gnew_n1377_
  (
    .dout(new_n1377__spl_),
    .din(new_n1377_)
  );


  splt
  gnew_n1302_
  (
    .dout(new_n1302__spl_),
    .din(new_n1302_)
  );


  splt
  gnew_n1379_
  (
    .dout(new_n1379__spl_),
    .din(new_n1379_)
  );


  splt
  gnew_n1380_
  (
    .dout(new_n1380__spl_),
    .din(new_n1380_)
  );


  splt
  gnew_n1301_
  (
    .dout(new_n1301__spl_),
    .din(new_n1301_)
  );


  splt
  gnew_n1382_
  (
    .dout(new_n1382__spl_),
    .din(new_n1382_)
  );


  splt
  gnew_n1383_
  (
    .dout(new_n1383__spl_),
    .din(new_n1383_)
  );


  splt
  gnew_n1300_
  (
    .dout(new_n1300__spl_),
    .din(new_n1300_)
  );


  splt
  gnew_n1385_
  (
    .dout(new_n1385__spl_),
    .din(new_n1385_)
  );


  splt
  gnew_n1386_
  (
    .dout(new_n1386__spl_),
    .din(new_n1386_)
  );


  splt
  gnew_n1299_
  (
    .dout(new_n1299__spl_),
    .din(new_n1299_)
  );


  splt
  gnew_n1388_
  (
    .dout(new_n1388__spl_),
    .din(new_n1388_)
  );


  splt
  gnew_n1389_
  (
    .dout(new_n1389__spl_),
    .din(new_n1389_)
  );


  splt
  gnew_n1298_
  (
    .dout(new_n1298__spl_),
    .din(new_n1298_)
  );


  splt
  gnew_n1391_
  (
    .dout(new_n1391__spl_),
    .din(new_n1391_)
  );


  splt
  gnew_n1392_
  (
    .dout(new_n1392__spl_),
    .din(new_n1392_)
  );


  splt
  gnew_n1416_
  (
    .dout(new_n1416__spl_),
    .din(new_n1416_)
  );


  splt
  gnew_n1417_
  (
    .dout(new_n1417__spl_),
    .din(new_n1417_)
  );


  splt
  gnew_n1418_
  (
    .dout(new_n1418__spl_),
    .din(new_n1418_)
  );


  splt
  gnew_n1415_
  (
    .dout(new_n1415__spl_),
    .din(new_n1415_)
  );


  splt
  gnew_n1420_
  (
    .dout(new_n1420__spl_),
    .din(new_n1420_)
  );


  splt
  gnew_n1421_
  (
    .dout(new_n1421__spl_),
    .din(new_n1421_)
  );


  splt
  gnew_n1414_
  (
    .dout(new_n1414__spl_),
    .din(new_n1414_)
  );


  splt
  gnew_n1423_
  (
    .dout(new_n1423__spl_),
    .din(new_n1423_)
  );


  splt
  gnew_n1424_
  (
    .dout(new_n1424__spl_),
    .din(new_n1424_)
  );


  splt
  gnew_n1413_
  (
    .dout(new_n1413__spl_),
    .din(new_n1413_)
  );


  splt
  gnew_n1426_
  (
    .dout(new_n1426__spl_),
    .din(new_n1426_)
  );


  splt
  gnew_n1427_
  (
    .dout(new_n1427__spl_),
    .din(new_n1427_)
  );


  splt
  gnew_n1412_
  (
    .dout(new_n1412__spl_),
    .din(new_n1412_)
  );


  splt
  gnew_n1429_
  (
    .dout(new_n1429__spl_),
    .din(new_n1429_)
  );


  splt
  gnew_n1430_
  (
    .dout(new_n1430__spl_),
    .din(new_n1430_)
  );


  splt
  gnew_n1411_
  (
    .dout(new_n1411__spl_),
    .din(new_n1411_)
  );


  splt
  gnew_n1432_
  (
    .dout(new_n1432__spl_),
    .din(new_n1432_)
  );


  splt
  gnew_n1433_
  (
    .dout(new_n1433__spl_),
    .din(new_n1433_)
  );


  splt
  gnew_n1410_
  (
    .dout(new_n1410__spl_),
    .din(new_n1410_)
  );


  splt
  gnew_n1435_
  (
    .dout(new_n1435__spl_),
    .din(new_n1435_)
  );


  splt
  gnew_n1436_
  (
    .dout(new_n1436__spl_),
    .din(new_n1436_)
  );


  splt
  gnew_n1409_
  (
    .dout(new_n1409__spl_),
    .din(new_n1409_)
  );


  splt
  gnew_n1438_
  (
    .dout(new_n1438__spl_),
    .din(new_n1438_)
  );


  splt
  gnew_n1439_
  (
    .dout(new_n1439__spl_),
    .din(new_n1439_)
  );


  splt
  gnew_n1408_
  (
    .dout(new_n1408__spl_),
    .din(new_n1408_)
  );


  splt
  gnew_n1441_
  (
    .dout(new_n1441__spl_),
    .din(new_n1441_)
  );


  splt
  gnew_n1442_
  (
    .dout(new_n1442__spl_),
    .din(new_n1442_)
  );


  splt
  gnew_n1407_
  (
    .dout(new_n1407__spl_),
    .din(new_n1407_)
  );


  splt
  gnew_n1444_
  (
    .dout(new_n1444__spl_),
    .din(new_n1444_)
  );


  splt
  gnew_n1445_
  (
    .dout(new_n1445__spl_),
    .din(new_n1445_)
  );


  splt
  gnew_n1406_
  (
    .dout(new_n1406__spl_),
    .din(new_n1406_)
  );


  splt
  gnew_n1447_
  (
    .dout(new_n1447__spl_),
    .din(new_n1447_)
  );


  splt
  gnew_n1448_
  (
    .dout(new_n1448__spl_),
    .din(new_n1448_)
  );


  splt
  gnew_n1405_
  (
    .dout(new_n1405__spl_),
    .din(new_n1405_)
  );


  splt
  gnew_n1450_
  (
    .dout(new_n1450__spl_),
    .din(new_n1450_)
  );


  splt
  gnew_n1451_
  (
    .dout(new_n1451__spl_),
    .din(new_n1451_)
  );


  splt
  gnew_n1404_
  (
    .dout(new_n1404__spl_),
    .din(new_n1404_)
  );


  splt
  gnew_n1453_
  (
    .dout(new_n1453__spl_),
    .din(new_n1453_)
  );


  splt
  gnew_n1454_
  (
    .dout(new_n1454__spl_),
    .din(new_n1454_)
  );


  splt
  gnew_n1403_
  (
    .dout(new_n1403__spl_),
    .din(new_n1403_)
  );


  splt
  gnew_n1456_
  (
    .dout(new_n1456__spl_),
    .din(new_n1456_)
  );


  splt
  gnew_n1457_
  (
    .dout(new_n1457__spl_),
    .din(new_n1457_)
  );


  splt
  gnew_n1402_
  (
    .dout(new_n1402__spl_),
    .din(new_n1402_)
  );


  splt
  gnew_n1459_
  (
    .dout(new_n1459__spl_),
    .din(new_n1459_)
  );


  splt
  gnew_n1460_
  (
    .dout(new_n1460__spl_),
    .din(new_n1460_)
  );


  splt
  gnew_n1401_
  (
    .dout(new_n1401__spl_),
    .din(new_n1401_)
  );


  splt
  gnew_n1462_
  (
    .dout(new_n1462__spl_),
    .din(new_n1462_)
  );


  splt
  gnew_n1463_
  (
    .dout(new_n1463__spl_),
    .din(new_n1463_)
  );


  splt
  gnew_n1400_
  (
    .dout(new_n1400__spl_),
    .din(new_n1400_)
  );


  splt
  gnew_n1465_
  (
    .dout(new_n1465__spl_),
    .din(new_n1465_)
  );


  splt
  gnew_n1466_
  (
    .dout(new_n1466__spl_),
    .din(new_n1466_)
  );


  splt
  gnew_n1399_
  (
    .dout(new_n1399__spl_),
    .din(new_n1399_)
  );


  splt
  gnew_n1468_
  (
    .dout(new_n1468__spl_),
    .din(new_n1468_)
  );


  splt
  gnew_n1469_
  (
    .dout(new_n1469__spl_),
    .din(new_n1469_)
  );


  splt
  gnew_n1398_
  (
    .dout(new_n1398__spl_),
    .din(new_n1398_)
  );


  splt
  gnew_n1471_
  (
    .dout(new_n1471__spl_),
    .din(new_n1471_)
  );


  splt
  gnew_n1472_
  (
    .dout(new_n1472__spl_),
    .din(new_n1472_)
  );


  splt
  gnew_n1397_
  (
    .dout(new_n1397__spl_),
    .din(new_n1397_)
  );


  splt
  gnew_n1474_
  (
    .dout(new_n1474__spl_),
    .din(new_n1474_)
  );


  splt
  gnew_n1475_
  (
    .dout(new_n1475__spl_),
    .din(new_n1475_)
  );


  splt
  gnew_n1396_
  (
    .dout(new_n1396__spl_),
    .din(new_n1396_)
  );


  splt
  gnew_n1477_
  (
    .dout(new_n1477__spl_),
    .din(new_n1477_)
  );


  splt
  gnew_n1478_
  (
    .dout(new_n1478__spl_),
    .din(new_n1478_)
  );


  splt
  gnew_n1395_
  (
    .dout(new_n1395__spl_),
    .din(new_n1395_)
  );


  splt
  gnew_n1480_
  (
    .dout(new_n1480__spl_),
    .din(new_n1480_)
  );


  splt
  gnew_n1481_
  (
    .dout(new_n1481__spl_),
    .din(new_n1481_)
  );


  splt
  gnew_n1503_
  (
    .dout(new_n1503__spl_),
    .din(new_n1503_)
  );


  splt
  gnew_n1504_
  (
    .dout(new_n1504__spl_),
    .din(new_n1504_)
  );


  splt
  gnew_n1505_
  (
    .dout(new_n1505__spl_),
    .din(new_n1505_)
  );


  splt
  gnew_n1502_
  (
    .dout(new_n1502__spl_),
    .din(new_n1502_)
  );


  splt
  gnew_n1507_
  (
    .dout(new_n1507__spl_),
    .din(new_n1507_)
  );


  splt
  gnew_n1508_
  (
    .dout(new_n1508__spl_),
    .din(new_n1508_)
  );


  splt
  gnew_n1501_
  (
    .dout(new_n1501__spl_),
    .din(new_n1501_)
  );


  splt
  gnew_n1510_
  (
    .dout(new_n1510__spl_),
    .din(new_n1510_)
  );


  splt
  gnew_n1511_
  (
    .dout(new_n1511__spl_),
    .din(new_n1511_)
  );


  splt
  gnew_n1500_
  (
    .dout(new_n1500__spl_),
    .din(new_n1500_)
  );


  splt
  gnew_n1513_
  (
    .dout(new_n1513__spl_),
    .din(new_n1513_)
  );


  splt
  gnew_n1514_
  (
    .dout(new_n1514__spl_),
    .din(new_n1514_)
  );


  splt
  gnew_n1499_
  (
    .dout(new_n1499__spl_),
    .din(new_n1499_)
  );


  splt
  gnew_n1516_
  (
    .dout(new_n1516__spl_),
    .din(new_n1516_)
  );


  splt
  gnew_n1517_
  (
    .dout(new_n1517__spl_),
    .din(new_n1517_)
  );


  splt
  gnew_n1498_
  (
    .dout(new_n1498__spl_),
    .din(new_n1498_)
  );


  splt
  gnew_n1519_
  (
    .dout(new_n1519__spl_),
    .din(new_n1519_)
  );


  splt
  gnew_n1520_
  (
    .dout(new_n1520__spl_),
    .din(new_n1520_)
  );


  splt
  gnew_n1497_
  (
    .dout(new_n1497__spl_),
    .din(new_n1497_)
  );


  splt
  gnew_n1522_
  (
    .dout(new_n1522__spl_),
    .din(new_n1522_)
  );


  splt
  gnew_n1523_
  (
    .dout(new_n1523__spl_),
    .din(new_n1523_)
  );


  splt
  gnew_n1496_
  (
    .dout(new_n1496__spl_),
    .din(new_n1496_)
  );


  splt
  gnew_n1525_
  (
    .dout(new_n1525__spl_),
    .din(new_n1525_)
  );


  splt
  gnew_n1526_
  (
    .dout(new_n1526__spl_),
    .din(new_n1526_)
  );


  splt
  gnew_n1495_
  (
    .dout(new_n1495__spl_),
    .din(new_n1495_)
  );


  splt
  gnew_n1528_
  (
    .dout(new_n1528__spl_),
    .din(new_n1528_)
  );


  splt
  gnew_n1529_
  (
    .dout(new_n1529__spl_),
    .din(new_n1529_)
  );


  splt
  gnew_n1494_
  (
    .dout(new_n1494__spl_),
    .din(new_n1494_)
  );


  splt
  gnew_n1531_
  (
    .dout(new_n1531__spl_),
    .din(new_n1531_)
  );


  splt
  gnew_n1532_
  (
    .dout(new_n1532__spl_),
    .din(new_n1532_)
  );


  splt
  gnew_n1493_
  (
    .dout(new_n1493__spl_),
    .din(new_n1493_)
  );


  splt
  gnew_n1534_
  (
    .dout(new_n1534__spl_),
    .din(new_n1534_)
  );


  splt
  gnew_n1535_
  (
    .dout(new_n1535__spl_),
    .din(new_n1535_)
  );


  splt
  gnew_n1492_
  (
    .dout(new_n1492__spl_),
    .din(new_n1492_)
  );


  splt
  gnew_n1537_
  (
    .dout(new_n1537__spl_),
    .din(new_n1537_)
  );


  splt
  gnew_n1538_
  (
    .dout(new_n1538__spl_),
    .din(new_n1538_)
  );


  splt
  gnew_n1491_
  (
    .dout(new_n1491__spl_),
    .din(new_n1491_)
  );


  splt
  gnew_n1540_
  (
    .dout(new_n1540__spl_),
    .din(new_n1540_)
  );


  splt
  gnew_n1541_
  (
    .dout(new_n1541__spl_),
    .din(new_n1541_)
  );


  splt
  gnew_n1490_
  (
    .dout(new_n1490__spl_),
    .din(new_n1490_)
  );


  splt
  gnew_n1543_
  (
    .dout(new_n1543__spl_),
    .din(new_n1543_)
  );


  splt
  gnew_n1544_
  (
    .dout(new_n1544__spl_),
    .din(new_n1544_)
  );


  splt
  gnew_n1489_
  (
    .dout(new_n1489__spl_),
    .din(new_n1489_)
  );


  splt
  gnew_n1546_
  (
    .dout(new_n1546__spl_),
    .din(new_n1546_)
  );


  splt
  gnew_n1547_
  (
    .dout(new_n1547__spl_),
    .din(new_n1547_)
  );


  splt
  gnew_n1488_
  (
    .dout(new_n1488__spl_),
    .din(new_n1488_)
  );


  splt
  gnew_n1549_
  (
    .dout(new_n1549__spl_),
    .din(new_n1549_)
  );


  splt
  gnew_n1550_
  (
    .dout(new_n1550__spl_),
    .din(new_n1550_)
  );


  splt
  gnew_n1487_
  (
    .dout(new_n1487__spl_),
    .din(new_n1487_)
  );


  splt
  gnew_n1552_
  (
    .dout(new_n1552__spl_),
    .din(new_n1552_)
  );


  splt
  gnew_n1553_
  (
    .dout(new_n1553__spl_),
    .din(new_n1553_)
  );


  splt
  gnew_n1486_
  (
    .dout(new_n1486__spl_),
    .din(new_n1486_)
  );


  splt
  gnew_n1555_
  (
    .dout(new_n1555__spl_),
    .din(new_n1555_)
  );


  splt
  gnew_n1556_
  (
    .dout(new_n1556__spl_),
    .din(new_n1556_)
  );


  splt
  gnew_n1485_
  (
    .dout(new_n1485__spl_),
    .din(new_n1485_)
  );


  splt
  gnew_n1558_
  (
    .dout(new_n1558__spl_),
    .din(new_n1558_)
  );


  splt
  gnew_n1559_
  (
    .dout(new_n1559__spl_),
    .din(new_n1559_)
  );


  splt
  gnew_n1484_
  (
    .dout(new_n1484__spl_),
    .din(new_n1484_)
  );


  splt
  gnew_n1561_
  (
    .dout(new_n1561__spl_),
    .din(new_n1561_)
  );


  splt
  gnew_n1562_
  (
    .dout(new_n1562__spl_),
    .din(new_n1562_)
  );


  splt
  gnew_n1582_
  (
    .dout(new_n1582__spl_),
    .din(new_n1582_)
  );


  splt
  gnew_n1583_
  (
    .dout(new_n1583__spl_),
    .din(new_n1583_)
  );


  splt
  gnew_n1584_
  (
    .dout(new_n1584__spl_),
    .din(new_n1584_)
  );


  splt
  gnew_n1581_
  (
    .dout(new_n1581__spl_),
    .din(new_n1581_)
  );


  splt
  gnew_n1586_
  (
    .dout(new_n1586__spl_),
    .din(new_n1586_)
  );


  splt
  gnew_n1587_
  (
    .dout(new_n1587__spl_),
    .din(new_n1587_)
  );


  splt
  gnew_n1580_
  (
    .dout(new_n1580__spl_),
    .din(new_n1580_)
  );


  splt
  gnew_n1589_
  (
    .dout(new_n1589__spl_),
    .din(new_n1589_)
  );


  splt
  gnew_n1590_
  (
    .dout(new_n1590__spl_),
    .din(new_n1590_)
  );


  splt
  gnew_n1579_
  (
    .dout(new_n1579__spl_),
    .din(new_n1579_)
  );


  splt
  gnew_n1592_
  (
    .dout(new_n1592__spl_),
    .din(new_n1592_)
  );


  splt
  gnew_n1593_
  (
    .dout(new_n1593__spl_),
    .din(new_n1593_)
  );


  splt
  gnew_n1578_
  (
    .dout(new_n1578__spl_),
    .din(new_n1578_)
  );


  splt
  gnew_n1595_
  (
    .dout(new_n1595__spl_),
    .din(new_n1595_)
  );


  splt
  gnew_n1596_
  (
    .dout(new_n1596__spl_),
    .din(new_n1596_)
  );


  splt
  gnew_n1577_
  (
    .dout(new_n1577__spl_),
    .din(new_n1577_)
  );


  splt
  gnew_n1598_
  (
    .dout(new_n1598__spl_),
    .din(new_n1598_)
  );


  splt
  gnew_n1599_
  (
    .dout(new_n1599__spl_),
    .din(new_n1599_)
  );


  splt
  gnew_n1576_
  (
    .dout(new_n1576__spl_),
    .din(new_n1576_)
  );


  splt
  gnew_n1601_
  (
    .dout(new_n1601__spl_),
    .din(new_n1601_)
  );


  splt
  gnew_n1602_
  (
    .dout(new_n1602__spl_),
    .din(new_n1602_)
  );


  splt
  gnew_n1575_
  (
    .dout(new_n1575__spl_),
    .din(new_n1575_)
  );


  splt
  gnew_n1604_
  (
    .dout(new_n1604__spl_),
    .din(new_n1604_)
  );


  splt
  gnew_n1605_
  (
    .dout(new_n1605__spl_),
    .din(new_n1605_)
  );


  splt
  gnew_n1574_
  (
    .dout(new_n1574__spl_),
    .din(new_n1574_)
  );


  splt
  gnew_n1607_
  (
    .dout(new_n1607__spl_),
    .din(new_n1607_)
  );


  splt
  gnew_n1608_
  (
    .dout(new_n1608__spl_),
    .din(new_n1608_)
  );


  splt
  gnew_n1573_
  (
    .dout(new_n1573__spl_),
    .din(new_n1573_)
  );


  splt
  gnew_n1610_
  (
    .dout(new_n1610__spl_),
    .din(new_n1610_)
  );


  splt
  gnew_n1611_
  (
    .dout(new_n1611__spl_),
    .din(new_n1611_)
  );


  splt
  gnew_n1572_
  (
    .dout(new_n1572__spl_),
    .din(new_n1572_)
  );


  splt
  gnew_n1613_
  (
    .dout(new_n1613__spl_),
    .din(new_n1613_)
  );


  splt
  gnew_n1614_
  (
    .dout(new_n1614__spl_),
    .din(new_n1614_)
  );


  splt
  gnew_n1571_
  (
    .dout(new_n1571__spl_),
    .din(new_n1571_)
  );


  splt
  gnew_n1616_
  (
    .dout(new_n1616__spl_),
    .din(new_n1616_)
  );


  splt
  gnew_n1617_
  (
    .dout(new_n1617__spl_),
    .din(new_n1617_)
  );


  splt
  gnew_n1570_
  (
    .dout(new_n1570__spl_),
    .din(new_n1570_)
  );


  splt
  gnew_n1619_
  (
    .dout(new_n1619__spl_),
    .din(new_n1619_)
  );


  splt
  gnew_n1620_
  (
    .dout(new_n1620__spl_),
    .din(new_n1620_)
  );


  splt
  gnew_n1569_
  (
    .dout(new_n1569__spl_),
    .din(new_n1569_)
  );


  splt
  gnew_n1622_
  (
    .dout(new_n1622__spl_),
    .din(new_n1622_)
  );


  splt
  gnew_n1623_
  (
    .dout(new_n1623__spl_),
    .din(new_n1623_)
  );


  splt
  gnew_n1568_
  (
    .dout(new_n1568__spl_),
    .din(new_n1568_)
  );


  splt
  gnew_n1625_
  (
    .dout(new_n1625__spl_),
    .din(new_n1625_)
  );


  splt
  gnew_n1626_
  (
    .dout(new_n1626__spl_),
    .din(new_n1626_)
  );


  splt
  gnew_n1567_
  (
    .dout(new_n1567__spl_),
    .din(new_n1567_)
  );


  splt
  gnew_n1628_
  (
    .dout(new_n1628__spl_),
    .din(new_n1628_)
  );


  splt
  gnew_n1629_
  (
    .dout(new_n1629__spl_),
    .din(new_n1629_)
  );


  splt
  gnew_n1566_
  (
    .dout(new_n1566__spl_),
    .din(new_n1566_)
  );


  splt
  gnew_n1631_
  (
    .dout(new_n1631__spl_),
    .din(new_n1631_)
  );


  splt
  gnew_n1632_
  (
    .dout(new_n1632__spl_),
    .din(new_n1632_)
  );


  splt
  gnew_n1565_
  (
    .dout(new_n1565__spl_),
    .din(new_n1565_)
  );


  splt
  gnew_n1634_
  (
    .dout(new_n1634__spl_),
    .din(new_n1634_)
  );


  splt
  gnew_n1635_
  (
    .dout(new_n1635__spl_),
    .din(new_n1635_)
  );


  splt
  gnew_n1653_
  (
    .dout(new_n1653__spl_),
    .din(new_n1653_)
  );


  splt
  gnew_n1654_
  (
    .dout(new_n1654__spl_),
    .din(new_n1654_)
  );


  splt
  gnew_n1655_
  (
    .dout(new_n1655__spl_),
    .din(new_n1655_)
  );


  splt
  gnew_n1652_
  (
    .dout(new_n1652__spl_),
    .din(new_n1652_)
  );


  splt
  gnew_n1657_
  (
    .dout(new_n1657__spl_),
    .din(new_n1657_)
  );


  splt
  gnew_n1658_
  (
    .dout(new_n1658__spl_),
    .din(new_n1658_)
  );


  splt
  gnew_n1651_
  (
    .dout(new_n1651__spl_),
    .din(new_n1651_)
  );


  splt
  gnew_n1660_
  (
    .dout(new_n1660__spl_),
    .din(new_n1660_)
  );


  splt
  gnew_n1661_
  (
    .dout(new_n1661__spl_),
    .din(new_n1661_)
  );


  splt
  gnew_n1650_
  (
    .dout(new_n1650__spl_),
    .din(new_n1650_)
  );


  splt
  gnew_n1663_
  (
    .dout(new_n1663__spl_),
    .din(new_n1663_)
  );


  splt
  gnew_n1664_
  (
    .dout(new_n1664__spl_),
    .din(new_n1664_)
  );


  splt
  gnew_n1649_
  (
    .dout(new_n1649__spl_),
    .din(new_n1649_)
  );


  splt
  gnew_n1666_
  (
    .dout(new_n1666__spl_),
    .din(new_n1666_)
  );


  splt
  gnew_n1667_
  (
    .dout(new_n1667__spl_),
    .din(new_n1667_)
  );


  splt
  gnew_n1648_
  (
    .dout(new_n1648__spl_),
    .din(new_n1648_)
  );


  splt
  gnew_n1669_
  (
    .dout(new_n1669__spl_),
    .din(new_n1669_)
  );


  splt
  gnew_n1670_
  (
    .dout(new_n1670__spl_),
    .din(new_n1670_)
  );


  splt
  gnew_n1647_
  (
    .dout(new_n1647__spl_),
    .din(new_n1647_)
  );


  splt
  gnew_n1672_
  (
    .dout(new_n1672__spl_),
    .din(new_n1672_)
  );


  splt
  gnew_n1673_
  (
    .dout(new_n1673__spl_),
    .din(new_n1673_)
  );


  splt
  gnew_n1646_
  (
    .dout(new_n1646__spl_),
    .din(new_n1646_)
  );


  splt
  gnew_n1675_
  (
    .dout(new_n1675__spl_),
    .din(new_n1675_)
  );


  splt
  gnew_n1676_
  (
    .dout(new_n1676__spl_),
    .din(new_n1676_)
  );


  splt
  gnew_n1645_
  (
    .dout(new_n1645__spl_),
    .din(new_n1645_)
  );


  splt
  gnew_n1678_
  (
    .dout(new_n1678__spl_),
    .din(new_n1678_)
  );


  splt
  gnew_n1679_
  (
    .dout(new_n1679__spl_),
    .din(new_n1679_)
  );


  splt
  gnew_n1644_
  (
    .dout(new_n1644__spl_),
    .din(new_n1644_)
  );


  splt
  gnew_n1681_
  (
    .dout(new_n1681__spl_),
    .din(new_n1681_)
  );


  splt
  gnew_n1682_
  (
    .dout(new_n1682__spl_),
    .din(new_n1682_)
  );


  splt
  gnew_n1643_
  (
    .dout(new_n1643__spl_),
    .din(new_n1643_)
  );


  splt
  gnew_n1684_
  (
    .dout(new_n1684__spl_),
    .din(new_n1684_)
  );


  splt
  gnew_n1685_
  (
    .dout(new_n1685__spl_),
    .din(new_n1685_)
  );


  splt
  gnew_n1642_
  (
    .dout(new_n1642__spl_),
    .din(new_n1642_)
  );


  splt
  gnew_n1687_
  (
    .dout(new_n1687__spl_),
    .din(new_n1687_)
  );


  splt
  gnew_n1688_
  (
    .dout(new_n1688__spl_),
    .din(new_n1688_)
  );


  splt
  gnew_n1641_
  (
    .dout(new_n1641__spl_),
    .din(new_n1641_)
  );


  splt
  gnew_n1690_
  (
    .dout(new_n1690__spl_),
    .din(new_n1690_)
  );


  splt
  gnew_n1691_
  (
    .dout(new_n1691__spl_),
    .din(new_n1691_)
  );


  splt
  gnew_n1640_
  (
    .dout(new_n1640__spl_),
    .din(new_n1640_)
  );


  splt
  gnew_n1693_
  (
    .dout(new_n1693__spl_),
    .din(new_n1693_)
  );


  splt
  gnew_n1694_
  (
    .dout(new_n1694__spl_),
    .din(new_n1694_)
  );


  splt
  gnew_n1639_
  (
    .dout(new_n1639__spl_),
    .din(new_n1639_)
  );


  splt
  gnew_n1696_
  (
    .dout(new_n1696__spl_),
    .din(new_n1696_)
  );


  splt
  gnew_n1697_
  (
    .dout(new_n1697__spl_),
    .din(new_n1697_)
  );


  splt
  gnew_n1638_
  (
    .dout(new_n1638__spl_),
    .din(new_n1638_)
  );


  splt
  gnew_n1699_
  (
    .dout(new_n1699__spl_),
    .din(new_n1699_)
  );


  splt
  gnew_n1700_
  (
    .dout(new_n1700__spl_),
    .din(new_n1700_)
  );


  splt
  gnew_n1716_
  (
    .dout(new_n1716__spl_),
    .din(new_n1716_)
  );


  splt
  gnew_n1717_
  (
    .dout(new_n1717__spl_),
    .din(new_n1717_)
  );


  splt
  gnew_n1718_
  (
    .dout(new_n1718__spl_),
    .din(new_n1718_)
  );


  splt
  gnew_n1715_
  (
    .dout(new_n1715__spl_),
    .din(new_n1715_)
  );


  splt
  gnew_n1720_
  (
    .dout(new_n1720__spl_),
    .din(new_n1720_)
  );


  splt
  gnew_n1721_
  (
    .dout(new_n1721__spl_),
    .din(new_n1721_)
  );


  splt
  gnew_n1714_
  (
    .dout(new_n1714__spl_),
    .din(new_n1714_)
  );


  splt
  gnew_n1723_
  (
    .dout(new_n1723__spl_),
    .din(new_n1723_)
  );


  splt
  gnew_n1724_
  (
    .dout(new_n1724__spl_),
    .din(new_n1724_)
  );


  splt
  gnew_n1713_
  (
    .dout(new_n1713__spl_),
    .din(new_n1713_)
  );


  splt
  gnew_n1726_
  (
    .dout(new_n1726__spl_),
    .din(new_n1726_)
  );


  splt
  gnew_n1727_
  (
    .dout(new_n1727__spl_),
    .din(new_n1727_)
  );


  splt
  gnew_n1712_
  (
    .dout(new_n1712__spl_),
    .din(new_n1712_)
  );


  splt
  gnew_n1729_
  (
    .dout(new_n1729__spl_),
    .din(new_n1729_)
  );


  splt
  gnew_n1730_
  (
    .dout(new_n1730__spl_),
    .din(new_n1730_)
  );


  splt
  gnew_n1711_
  (
    .dout(new_n1711__spl_),
    .din(new_n1711_)
  );


  splt
  gnew_n1732_
  (
    .dout(new_n1732__spl_),
    .din(new_n1732_)
  );


  splt
  gnew_n1733_
  (
    .dout(new_n1733__spl_),
    .din(new_n1733_)
  );


  splt
  gnew_n1710_
  (
    .dout(new_n1710__spl_),
    .din(new_n1710_)
  );


  splt
  gnew_n1735_
  (
    .dout(new_n1735__spl_),
    .din(new_n1735_)
  );


  splt
  gnew_n1736_
  (
    .dout(new_n1736__spl_),
    .din(new_n1736_)
  );


  splt
  gnew_n1709_
  (
    .dout(new_n1709__spl_),
    .din(new_n1709_)
  );


  splt
  gnew_n1738_
  (
    .dout(new_n1738__spl_),
    .din(new_n1738_)
  );


  splt
  gnew_n1739_
  (
    .dout(new_n1739__spl_),
    .din(new_n1739_)
  );


  splt
  gnew_n1708_
  (
    .dout(new_n1708__spl_),
    .din(new_n1708_)
  );


  splt
  gnew_n1741_
  (
    .dout(new_n1741__spl_),
    .din(new_n1741_)
  );


  splt
  gnew_n1742_
  (
    .dout(new_n1742__spl_),
    .din(new_n1742_)
  );


  splt
  gnew_n1707_
  (
    .dout(new_n1707__spl_),
    .din(new_n1707_)
  );


  splt
  gnew_n1744_
  (
    .dout(new_n1744__spl_),
    .din(new_n1744_)
  );


  splt
  gnew_n1745_
  (
    .dout(new_n1745__spl_),
    .din(new_n1745_)
  );


  splt
  gnew_n1706_
  (
    .dout(new_n1706__spl_),
    .din(new_n1706_)
  );


  splt
  gnew_n1747_
  (
    .dout(new_n1747__spl_),
    .din(new_n1747_)
  );


  splt
  gnew_n1748_
  (
    .dout(new_n1748__spl_),
    .din(new_n1748_)
  );


  splt
  gnew_n1705_
  (
    .dout(new_n1705__spl_),
    .din(new_n1705_)
  );


  splt
  gnew_n1750_
  (
    .dout(new_n1750__spl_),
    .din(new_n1750_)
  );


  splt
  gnew_n1751_
  (
    .dout(new_n1751__spl_),
    .din(new_n1751_)
  );


  splt
  gnew_n1704_
  (
    .dout(new_n1704__spl_),
    .din(new_n1704_)
  );


  splt
  gnew_n1753_
  (
    .dout(new_n1753__spl_),
    .din(new_n1753_)
  );


  splt
  gnew_n1754_
  (
    .dout(new_n1754__spl_),
    .din(new_n1754_)
  );


  splt
  gnew_n1703_
  (
    .dout(new_n1703__spl_),
    .din(new_n1703_)
  );


  splt
  gnew_n1756_
  (
    .dout(new_n1756__spl_),
    .din(new_n1756_)
  );


  splt
  gnew_n1757_
  (
    .dout(new_n1757__spl_),
    .din(new_n1757_)
  );


  splt
  gnew_n1771_
  (
    .dout(new_n1771__spl_),
    .din(new_n1771_)
  );


  splt
  gnew_n1772_
  (
    .dout(new_n1772__spl_),
    .din(new_n1772_)
  );


  splt
  gnew_n1773_
  (
    .dout(new_n1773__spl_),
    .din(new_n1773_)
  );


  splt
  gnew_n1770_
  (
    .dout(new_n1770__spl_),
    .din(new_n1770_)
  );


  splt
  gnew_n1775_
  (
    .dout(new_n1775__spl_),
    .din(new_n1775_)
  );


  splt
  gnew_n1776_
  (
    .dout(new_n1776__spl_),
    .din(new_n1776_)
  );


  splt
  gnew_n1769_
  (
    .dout(new_n1769__spl_),
    .din(new_n1769_)
  );


  splt
  gnew_n1778_
  (
    .dout(new_n1778__spl_),
    .din(new_n1778_)
  );


  splt
  gnew_n1779_
  (
    .dout(new_n1779__spl_),
    .din(new_n1779_)
  );


  splt
  gnew_n1768_
  (
    .dout(new_n1768__spl_),
    .din(new_n1768_)
  );


  splt
  gnew_n1781_
  (
    .dout(new_n1781__spl_),
    .din(new_n1781_)
  );


  splt
  gnew_n1782_
  (
    .dout(new_n1782__spl_),
    .din(new_n1782_)
  );


  splt
  gnew_n1767_
  (
    .dout(new_n1767__spl_),
    .din(new_n1767_)
  );


  splt
  gnew_n1784_
  (
    .dout(new_n1784__spl_),
    .din(new_n1784_)
  );


  splt
  gnew_n1785_
  (
    .dout(new_n1785__spl_),
    .din(new_n1785_)
  );


  splt
  gnew_n1766_
  (
    .dout(new_n1766__spl_),
    .din(new_n1766_)
  );


  splt
  gnew_n1787_
  (
    .dout(new_n1787__spl_),
    .din(new_n1787_)
  );


  splt
  gnew_n1788_
  (
    .dout(new_n1788__spl_),
    .din(new_n1788_)
  );


  splt
  gnew_n1765_
  (
    .dout(new_n1765__spl_),
    .din(new_n1765_)
  );


  splt
  gnew_n1790_
  (
    .dout(new_n1790__spl_),
    .din(new_n1790_)
  );


  splt
  gnew_n1791_
  (
    .dout(new_n1791__spl_),
    .din(new_n1791_)
  );


  splt
  gnew_n1764_
  (
    .dout(new_n1764__spl_),
    .din(new_n1764_)
  );


  splt
  gnew_n1793_
  (
    .dout(new_n1793__spl_),
    .din(new_n1793_)
  );


  splt
  gnew_n1794_
  (
    .dout(new_n1794__spl_),
    .din(new_n1794_)
  );


  splt
  gnew_n1763_
  (
    .dout(new_n1763__spl_),
    .din(new_n1763_)
  );


  splt
  gnew_n1796_
  (
    .dout(new_n1796__spl_),
    .din(new_n1796_)
  );


  splt
  gnew_n1797_
  (
    .dout(new_n1797__spl_),
    .din(new_n1797_)
  );


  splt
  gnew_n1762_
  (
    .dout(new_n1762__spl_),
    .din(new_n1762_)
  );


  splt
  gnew_n1799_
  (
    .dout(new_n1799__spl_),
    .din(new_n1799_)
  );


  splt
  gnew_n1800_
  (
    .dout(new_n1800__spl_),
    .din(new_n1800_)
  );


  splt
  gnew_n1761_
  (
    .dout(new_n1761__spl_),
    .din(new_n1761_)
  );


  splt
  gnew_n1802_
  (
    .dout(new_n1802__spl_),
    .din(new_n1802_)
  );


  splt
  gnew_n1803_
  (
    .dout(new_n1803__spl_),
    .din(new_n1803_)
  );


  splt
  gnew_n1760_
  (
    .dout(new_n1760__spl_),
    .din(new_n1760_)
  );


  splt
  gnew_n1805_
  (
    .dout(new_n1805__spl_),
    .din(new_n1805_)
  );


  splt
  gnew_n1806_
  (
    .dout(new_n1806__spl_),
    .din(new_n1806_)
  );


  splt
  gnew_n1818_
  (
    .dout(new_n1818__spl_),
    .din(new_n1818_)
  );


  splt
  gnew_n1819_
  (
    .dout(new_n1819__spl_),
    .din(new_n1819_)
  );


  splt
  gnew_n1820_
  (
    .dout(new_n1820__spl_),
    .din(new_n1820_)
  );


  splt
  gnew_n1817_
  (
    .dout(new_n1817__spl_),
    .din(new_n1817_)
  );


  splt
  gnew_n1822_
  (
    .dout(new_n1822__spl_),
    .din(new_n1822_)
  );


  splt
  gnew_n1823_
  (
    .dout(new_n1823__spl_),
    .din(new_n1823_)
  );


  splt
  gnew_n1816_
  (
    .dout(new_n1816__spl_),
    .din(new_n1816_)
  );


  splt
  gnew_n1825_
  (
    .dout(new_n1825__spl_),
    .din(new_n1825_)
  );


  splt
  gnew_n1826_
  (
    .dout(new_n1826__spl_),
    .din(new_n1826_)
  );


  splt
  gnew_n1815_
  (
    .dout(new_n1815__spl_),
    .din(new_n1815_)
  );


  splt
  gnew_n1828_
  (
    .dout(new_n1828__spl_),
    .din(new_n1828_)
  );


  splt
  gnew_n1829_
  (
    .dout(new_n1829__spl_),
    .din(new_n1829_)
  );


  splt
  gnew_n1814_
  (
    .dout(new_n1814__spl_),
    .din(new_n1814_)
  );


  splt
  gnew_n1831_
  (
    .dout(new_n1831__spl_),
    .din(new_n1831_)
  );


  splt
  gnew_n1832_
  (
    .dout(new_n1832__spl_),
    .din(new_n1832_)
  );


  splt
  gnew_n1813_
  (
    .dout(new_n1813__spl_),
    .din(new_n1813_)
  );


  splt
  gnew_n1834_
  (
    .dout(new_n1834__spl_),
    .din(new_n1834_)
  );


  splt
  gnew_n1835_
  (
    .dout(new_n1835__spl_),
    .din(new_n1835_)
  );


  splt
  gnew_n1812_
  (
    .dout(new_n1812__spl_),
    .din(new_n1812_)
  );


  splt
  gnew_n1837_
  (
    .dout(new_n1837__spl_),
    .din(new_n1837_)
  );


  splt
  gnew_n1838_
  (
    .dout(new_n1838__spl_),
    .din(new_n1838_)
  );


  splt
  gnew_n1811_
  (
    .dout(new_n1811__spl_),
    .din(new_n1811_)
  );


  splt
  gnew_n1840_
  (
    .dout(new_n1840__spl_),
    .din(new_n1840_)
  );


  splt
  gnew_n1841_
  (
    .dout(new_n1841__spl_),
    .din(new_n1841_)
  );


  splt
  gnew_n1810_
  (
    .dout(new_n1810__spl_),
    .din(new_n1810_)
  );


  splt
  gnew_n1843_
  (
    .dout(new_n1843__spl_),
    .din(new_n1843_)
  );


  splt
  gnew_n1844_
  (
    .dout(new_n1844__spl_),
    .din(new_n1844_)
  );


  splt
  gnew_n1809_
  (
    .dout(new_n1809__spl_),
    .din(new_n1809_)
  );


  splt
  gnew_n1846_
  (
    .dout(new_n1846__spl_),
    .din(new_n1846_)
  );


  splt
  gnew_n1847_
  (
    .dout(new_n1847__spl_),
    .din(new_n1847_)
  );


  splt
  gnew_n1857_
  (
    .dout(new_n1857__spl_),
    .din(new_n1857_)
  );


  splt
  gnew_n1858_
  (
    .dout(new_n1858__spl_),
    .din(new_n1858_)
  );


  splt
  gnew_n1859_
  (
    .dout(new_n1859__spl_),
    .din(new_n1859_)
  );


  splt
  gnew_n1856_
  (
    .dout(new_n1856__spl_),
    .din(new_n1856_)
  );


  splt
  gnew_n1861_
  (
    .dout(new_n1861__spl_),
    .din(new_n1861_)
  );


  splt
  gnew_n1862_
  (
    .dout(new_n1862__spl_),
    .din(new_n1862_)
  );


  splt
  gnew_n1855_
  (
    .dout(new_n1855__spl_),
    .din(new_n1855_)
  );


  splt
  gnew_n1864_
  (
    .dout(new_n1864__spl_),
    .din(new_n1864_)
  );


  splt
  gnew_n1865_
  (
    .dout(new_n1865__spl_),
    .din(new_n1865_)
  );


  splt
  gnew_n1854_
  (
    .dout(new_n1854__spl_),
    .din(new_n1854_)
  );


  splt
  gnew_n1867_
  (
    .dout(new_n1867__spl_),
    .din(new_n1867_)
  );


  splt
  gnew_n1868_
  (
    .dout(new_n1868__spl_),
    .din(new_n1868_)
  );


  splt
  gnew_n1853_
  (
    .dout(new_n1853__spl_),
    .din(new_n1853_)
  );


  splt
  gnew_n1870_
  (
    .dout(new_n1870__spl_),
    .din(new_n1870_)
  );


  splt
  gnew_n1871_
  (
    .dout(new_n1871__spl_),
    .din(new_n1871_)
  );


  splt
  gnew_n1852_
  (
    .dout(new_n1852__spl_),
    .din(new_n1852_)
  );


  splt
  gnew_n1873_
  (
    .dout(new_n1873__spl_),
    .din(new_n1873_)
  );


  splt
  gnew_n1874_
  (
    .dout(new_n1874__spl_),
    .din(new_n1874_)
  );


  splt
  gnew_n1851_
  (
    .dout(new_n1851__spl_),
    .din(new_n1851_)
  );


  splt
  gnew_n1876_
  (
    .dout(new_n1876__spl_),
    .din(new_n1876_)
  );


  splt
  gnew_n1877_
  (
    .dout(new_n1877__spl_),
    .din(new_n1877_)
  );


  splt
  gnew_n1850_
  (
    .dout(new_n1850__spl_),
    .din(new_n1850_)
  );


  splt
  gnew_n1879_
  (
    .dout(new_n1879__spl_),
    .din(new_n1879_)
  );


  splt
  gnew_n1880_
  (
    .dout(new_n1880__spl_),
    .din(new_n1880_)
  );


  splt
  gnew_n1888_
  (
    .dout(new_n1888__spl_),
    .din(new_n1888_)
  );


  splt
  gnew_n1889_
  (
    .dout(new_n1889__spl_),
    .din(new_n1889_)
  );


  splt
  gnew_n1890_
  (
    .dout(new_n1890__spl_),
    .din(new_n1890_)
  );


  splt
  gnew_n1887_
  (
    .dout(new_n1887__spl_),
    .din(new_n1887_)
  );


  splt
  gnew_n1892_
  (
    .dout(new_n1892__spl_),
    .din(new_n1892_)
  );


  splt
  gnew_n1893_
  (
    .dout(new_n1893__spl_),
    .din(new_n1893_)
  );


  splt
  gnew_n1886_
  (
    .dout(new_n1886__spl_),
    .din(new_n1886_)
  );


  splt
  gnew_n1895_
  (
    .dout(new_n1895__spl_),
    .din(new_n1895_)
  );


  splt
  gnew_n1896_
  (
    .dout(new_n1896__spl_),
    .din(new_n1896_)
  );


  splt
  gnew_n1885_
  (
    .dout(new_n1885__spl_),
    .din(new_n1885_)
  );


  splt
  gnew_n1898_
  (
    .dout(new_n1898__spl_),
    .din(new_n1898_)
  );


  splt
  gnew_n1899_
  (
    .dout(new_n1899__spl_),
    .din(new_n1899_)
  );


  splt
  gnew_n1884_
  (
    .dout(new_n1884__spl_),
    .din(new_n1884_)
  );


  splt
  gnew_n1901_
  (
    .dout(new_n1901__spl_),
    .din(new_n1901_)
  );


  splt
  gnew_n1902_
  (
    .dout(new_n1902__spl_),
    .din(new_n1902_)
  );


  splt
  gnew_n1883_
  (
    .dout(new_n1883__spl_),
    .din(new_n1883_)
  );


  splt
  gnew_n1904_
  (
    .dout(new_n1904__spl_),
    .din(new_n1904_)
  );


  splt
  gnew_n1905_
  (
    .dout(new_n1905__spl_),
    .din(new_n1905_)
  );


  splt
  gnew_n1911_
  (
    .dout(new_n1911__spl_),
    .din(new_n1911_)
  );


  splt
  gnew_n1912_
  (
    .dout(new_n1912__spl_),
    .din(new_n1912_)
  );


  splt
  gnew_n1913_
  (
    .dout(new_n1913__spl_),
    .din(new_n1913_)
  );


  splt
  gnew_n1910_
  (
    .dout(new_n1910__spl_),
    .din(new_n1910_)
  );


  splt
  gnew_n1915_
  (
    .dout(new_n1915__spl_),
    .din(new_n1915_)
  );


  splt
  gnew_n1916_
  (
    .dout(new_n1916__spl_),
    .din(new_n1916_)
  );


  splt
  gnew_n1909_
  (
    .dout(new_n1909__spl_),
    .din(new_n1909_)
  );


  splt
  gnew_n1918_
  (
    .dout(new_n1918__spl_),
    .din(new_n1918_)
  );


  splt
  gnew_n1919_
  (
    .dout(new_n1919__spl_),
    .din(new_n1919_)
  );


  splt
  gnew_n1908_
  (
    .dout(new_n1908__spl_),
    .din(new_n1908_)
  );


  splt
  gnew_n1921_
  (
    .dout(new_n1921__spl_),
    .din(new_n1921_)
  );


  splt
  gnew_n1922_
  (
    .dout(new_n1922__spl_),
    .din(new_n1922_)
  );


  splt
  gnew_n1925_
  (
    .dout(new_n1925__spl_),
    .din(new_n1925_)
  );


  splt
  gnew_n1926_
  (
    .dout(new_n1926__spl_),
    .din(new_n1926_)
  );


  splt
  gnew_n1927_
  (
    .dout(new_n1927__spl_),
    .din(new_n1927_)
  );


  splt
  gnew_n1928_
  (
    .dout(new_n1928__spl_),
    .din(new_n1928_)
  );


  splt
  gnew_n1930_
  (
    .dout(new_n1930__spl_),
    .din(new_n1930_)
  );


  splt
  gnew_n1931_
  (
    .dout(new_n1931__spl_),
    .din(new_n1931_)
  );


endmodule
