
module mymod
(
  G1_p,
  G1_n,
  G2_p,
  G2_n,
  G3_p,
  G3_n,
  G4_p,
  G4_n,
  G5_p,
  G5_n,
  G6_p,
  G6_n,
  G7_p,
  G7_n,
  G8_p,
  G8_n,
  G9_p,
  G9_n,
  G10_p,
  G10_n,
  G11_p,
  G11_n,
  G12_p,
  G12_n,
  G13_p,
  G13_n,
  G14_p,
  G14_n,
  G15_p,
  G15_n,
  G16_p,
  G16_n,
  G17_p,
  G17_n,
  G18_p,
  G18_n,
  G19_p,
  G19_n,
  G20_p,
  G20_n,
  G21_p,
  G21_n,
  G22_p,
  G22_n,
  G23_p,
  G23_n,
  G24_p,
  G24_n,
  G25_p,
  G25_n,
  G26_p,
  G26_n,
  G27_p,
  G27_n,
  G28_p,
  G28_n,
  G29_p,
  G29_n,
  G30_p,
  G30_n,
  G31_p,
  G31_n,
  G32_p,
  G32_n,
  G33_p,
  G33_n,
  G34_p,
  G34_n,
  G35_p,
  G35_n,
  G36_p,
  G36_n,
  G426_p,
  G427_p,
  G428_p,
  G429_n,
  G430_n,
  G431_n,
  G432_n
);

  input G1_p;input G1_n;input G2_p;input G2_n;input G3_p;input G3_n;input G4_p;input G4_n;input G5_p;input G5_n;input G6_p;input G6_n;input G7_p;input G7_n;input G8_p;input G8_n;input G9_p;input G9_n;input G10_p;input G10_n;input G11_p;input G11_n;input G12_p;input G12_n;input G13_p;input G13_n;input G14_p;input G14_n;input G15_p;input G15_n;input G16_p;input G16_n;input G17_p;input G17_n;input G18_p;input G18_n;input G19_p;input G19_n;input G20_p;input G20_n;input G21_p;input G21_n;input G22_p;input G22_n;input G23_p;input G23_n;input G24_p;input G24_n;input G25_p;input G25_n;input G26_p;input G26_n;input G27_p;input G27_n;input G28_p;input G28_n;input G29_p;input G29_n;input G30_p;input G30_n;input G31_p;input G31_n;input G32_p;input G32_n;input G33_p;input G33_n;input G34_p;input G34_n;input G35_p;input G35_n;input G36_p;input G36_n;
  output G426_p;output G427_p;output G428_p;output G429_n;output G430_n;output G431_n;output G432_n;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire g37_p;
  wire g37_n;
  wire g38_p;
  wire g38_n;
  wire g39_p;
  wire g39_n;
  wire g40_p;
  wire g40_n;
  wire g41_p;
  wire g41_n;
  wire g42_p;
  wire g42_n;
  wire g43_p;
  wire g43_n;
  wire g44_p;
  wire g44_n;
  wire g45_p;
  wire g45_n;
  wire g46_p;
  wire g46_n;
  wire g47_p;
  wire g47_n;
  wire g48_p;
  wire g48_n;
  wire g49_p;
  wire g49_n;
  wire g50_p;
  wire g50_n;
  wire g51_p;
  wire g51_n;
  wire g52_p;
  wire g52_n;
  wire g53_p;
  wire g53_n;
  wire g54_p;
  wire g54_n;
  wire g55_p;
  wire g55_n;
  wire g56_p;
  wire g56_n;
  wire g57_p;
  wire g57_n;
  wire g58_p;
  wire g58_n;
  wire g59_p;
  wire g59_n;
  wire g60_p;
  wire g60_n;
  wire g61_p;
  wire g61_n;
  wire g62_p;
  wire g62_n;
  wire g63_p;
  wire g63_n;
  wire g64_p;
  wire g64_n;
  wire g65_p;
  wire g65_n;
  wire g66_p;
  wire g66_n;
  wire g67_p;
  wire g67_n;
  wire g68_p;
  wire g68_n;
  wire g69_p;
  wire g69_n;
  wire g70_p;
  wire g70_n;
  wire g71_p;
  wire g71_n;
  wire g72_p;
  wire g72_n;
  wire g73_p;
  wire g73_n;
  wire g74_p;
  wire g74_n;
  wire g75_p;
  wire g75_n;
  wire g76_p;
  wire g76_n;
  wire g77_p;
  wire g77_n;
  wire g78_p;
  wire g78_n;
  wire g79_p;
  wire g79_n;
  wire g80_p;
  wire g80_n;
  wire g81_p;
  wire g81_n;
  wire g82_p;
  wire g82_n;
  wire g83_p;
  wire g83_n;
  wire g84_p;
  wire g84_n;
  wire g85_p;
  wire g85_n;
  wire g86_p;
  wire g86_n;
  wire g87_p;
  wire g87_n;
  wire g88_p;
  wire g88_n;
  wire g89_p;
  wire g89_n;
  wire g90_p;
  wire g90_n;
  wire g91_p;
  wire g91_n;
  wire g92_p;
  wire g92_n;
  wire g93_p;
  wire g93_n;
  wire g94_p;
  wire g94_n;
  wire g95_p;
  wire g95_n;
  wire g96_p;
  wire g96_n;
  wire g97_p;
  wire g97_n;
  wire g98_p;
  wire g98_n;
  wire g99_p;
  wire g99_n;
  wire g100_p;
  wire g100_n;
  wire g101_p;
  wire g101_n;
  wire g102_p;
  wire g102_n;
  wire g103_p;
  wire g103_n;
  wire g104_p;
  wire g104_n;
  wire g105_p;
  wire g105_n;
  wire g106_p;
  wire g106_n;
  wire g107_p;
  wire g107_n;
  wire g108_p;
  wire g108_n;
  wire g109_p;
  wire g109_n;
  wire g110_p;
  wire g110_n;
  wire g111_p;
  wire g111_n;
  wire g112_p;
  wire g112_n;
  wire g113_p;
  wire g113_n;
  wire g114_p;
  wire g114_n;
  wire g115_p;
  wire g115_n;
  wire g116_p;
  wire g116_n;
  wire g117_p;
  wire g117_n;
  wire g118_p;
  wire g118_n;
  wire g119_p;
  wire g119_n;
  wire g120_p;
  wire g120_n;
  wire g121_p;
  wire g121_n;
  wire g122_p;
  wire g122_n;
  wire g123_p;
  wire g123_n;
  wire g124_p;
  wire g124_n;
  wire g125_p;
  wire g125_n;
  wire g126_p;
  wire g126_n;
  wire g127_p;
  wire g127_n;
  wire g128_p;
  wire g128_n;
  wire g129_p;
  wire g129_n;
  wire g130_p;
  wire g130_n;
  wire g131_p;
  wire g131_n;
  wire g132_p;
  wire g132_n;
  wire g133_p;
  wire g133_n;
  wire g134_p;
  wire g134_n;
  wire g135_p;
  wire g135_n;
  wire g136_p;
  wire g136_n;
  wire g137_p;
  wire g137_n;
  wire g138_p;
  wire g138_n;
  wire g139_p;
  wire g139_n;
  wire g140_p;
  wire g140_n;
  wire g141_p;
  wire g141_n;
  wire g142_p;
  wire g142_n;
  wire g143_p;
  wire g143_n;
  wire g144_p;
  wire g144_n;
  wire g145_p;
  wire g145_n;
  wire g146_p;
  wire g146_n;
  wire g147_p;
  wire g147_n;
  wire g148_p;
  wire g148_n;
  wire g149_p;
  wire g149_n;
  wire g150_p;
  wire g150_n;
  wire g151_p;
  wire g151_n;
  wire g152_p;
  wire g152_n;
  wire g153_p;
  wire g153_n;
  wire g154_p;
  wire g154_n;
  wire g155_p;
  wire g155_n;
  wire g156_p;
  wire g156_n;
  wire g157_p;
  wire g157_n;
  wire g158_p;
  wire g158_n;
  wire g159_p;
  wire g159_n;
  wire g160_p;
  wire g160_n;
  wire G16_n_spl_;
  wire G18_p_spl_;
  wire G16_p_spl_;
  wire G18_n_spl_;
  wire G12_n_spl_;
  wire G14_p_spl_;
  wire G12_p_spl_;
  wire G14_n_spl_;
  wire G1_n_spl_;
  wire G2_p_spl_;
  wire G1_p_spl_;
  wire G2_n_spl_;
  wire G28_n_spl_;
  wire G30_p_spl_;
  wire G28_p_spl_;
  wire G30_n_spl_;
  wire G32_n_spl_;
  wire G34_p_spl_;
  wire G32_p_spl_;
  wire G34_n_spl_;
  wire G20_n_spl_;
  wire G22_p_spl_;
  wire G20_p_spl_;
  wire G22_n_spl_;
  wire G24_n_spl_;
  wire G26_p_spl_;
  wire G24_p_spl_;
  wire G26_n_spl_;
  wire G4_n_spl_;
  wire G6_p_spl_;
  wire G4_p_spl_;
  wire G6_n_spl_;
  wire G8_n_spl_;
  wire G10_p_spl_;
  wire G8_p_spl_;
  wire G10_n_spl_;
  wire g53_n_spl_;
  wire g53_n_spl_0;
  wire g53_n_spl_00;
  wire g53_n_spl_000;
  wire g53_n_spl_001;
  wire g53_n_spl_01;
  wire g53_n_spl_1;
  wire g53_n_spl_10;
  wire g53_n_spl_11;
  wire g53_p_spl_;
  wire g53_p_spl_0;
  wire g53_p_spl_00;
  wire g53_p_spl_000;
  wire g53_p_spl_01;
  wire g53_p_spl_1;
  wire g53_p_spl_10;
  wire g53_p_spl_11;
  wire G11_n_spl_;
  wire g55_p_spl_;
  wire G11_p_spl_;
  wire g55_n_spl_;
  wire G35_n_spl_;
  wire g58_p_spl_;
  wire G35_p_spl_;
  wire g58_n_spl_;
  wire G7_n_spl_;
  wire g62_p_spl_;
  wire G7_p_spl_;
  wire g62_n_spl_;
  wire G23_n_spl_;
  wire g65_p_spl_;
  wire G23_p_spl_;
  wire g65_n_spl_;
  wire G15_n_spl_;
  wire g70_p_spl_;
  wire G15_p_spl_;
  wire g70_n_spl_;
  wire G3_n_spl_;
  wire g73_p_spl_;
  wire G3_p_spl_;
  wire g73_n_spl_;
  wire G19_n_spl_;
  wire g77_p_spl_;
  wire G19_p_spl_;
  wire g77_n_spl_;
  wire G31_n_spl_;
  wire g80_p_spl_;
  wire G31_p_spl_;
  wire g80_n_spl_;
  wire G27_n_spl_;
  wire g83_p_spl_;
  wire G27_p_spl_;
  wire g83_n_spl_;
  wire g88_n_spl_;
  wire g88_n_spl_0;
  wire g88_n_spl_00;
  wire g88_n_spl_000;
  wire g88_n_spl_001;
  wire g88_n_spl_01;
  wire g88_n_spl_1;
  wire g88_n_spl_10;
  wire g88_n_spl_11;
  wire g88_p_spl_;
  wire g88_p_spl_0;
  wire g88_p_spl_00;
  wire g88_p_spl_000;
  wire g88_p_spl_01;
  wire g88_p_spl_1;
  wire g88_p_spl_10;
  wire g88_p_spl_11;
  wire G13_n_spl_;
  wire g90_p_spl_;
  wire G13_p_spl_;
  wire g90_n_spl_;
  wire G36_p_spl_;
  wire g93_n_spl_;
  wire G9_p_spl_;
  wire g97_n_spl_;
  wire G25_p_spl_;
  wire g100_n_spl_;
  wire G17_n_spl_;
  wire g105_p_spl_;
  wire G17_p_spl_;
  wire g105_n_spl_;
  wire G5_n_spl_;
  wire g108_p_spl_;
  wire G21_n_spl_;
  wire g112_p_spl_;
  wire G21_p_spl_;
  wire g112_n_spl_;
  wire G33_p_spl_;
  wire g115_n_spl_;
  wire G29_n_spl_;
  wire g118_p_spl_;
  wire G29_p_spl_;
  wire g118_n_spl_;
  wire g123_p_spl_;
  wire g123_p_spl_0;
  wire g123_p_spl_00;
  wire g123_p_spl_1;
  wire g123_n_spl_;
  wire g123_n_spl_0;
  wire g123_n_spl_00;
  wire g123_n_spl_000;
  wire g123_n_spl_01;
  wire g123_n_spl_1;
  wire g123_n_spl_10;
  wire g123_n_spl_11;
  wire g131_n_spl_;
  wire g138_n_spl_;
  wire g136_p_spl_;
  wire g138_p_spl_;
  wire g134_p_spl_;
  wire g144_n_spl_;
  wire g140_p_spl_;
  wire g129_n_spl_;
  wire g127_n_spl_;
  wire g133_p_spl_;
  wire g153_n_spl_;

  LA
  g_g37_p
  (
    .dout(g37_p),
    .din1(G16_n_spl_),
    .din2(G18_p_spl_)
  );


  FA
  g_g37_n
  (
    .dout(g37_n),
    .din1(G16_p_spl_),
    .din2(G18_n_spl_)
  );


  LA
  g_g38_p
  (
    .dout(g38_p),
    .din1(G12_n_spl_),
    .din2(G14_p_spl_)
  );


  FA
  g_g38_n
  (
    .dout(g38_n),
    .din1(G12_p_spl_),
    .din2(G14_n_spl_)
  );


  LA
  g_g39_p
  (
    .dout(g39_p),
    .din1(g37_n),
    .din2(g38_n)
  );


  FA
  g_g39_n
  (
    .dout(g39_n),
    .din1(g37_p),
    .din2(g38_p)
  );


  LA
  g_g40_p
  (
    .dout(g40_p),
    .din1(G1_n_spl_),
    .din2(G2_p_spl_)
  );


  FA
  g_g40_n
  (
    .dout(g40_n),
    .din1(G1_p_spl_),
    .din2(G2_n_spl_)
  );


  LA
  g_g41_p
  (
    .dout(g41_p),
    .din1(G28_n_spl_),
    .din2(G30_p_spl_)
  );


  FA
  g_g41_n
  (
    .dout(g41_n),
    .din1(G28_p_spl_),
    .din2(G30_n_spl_)
  );


  LA
  g_g42_p
  (
    .dout(g42_p),
    .din1(g40_n),
    .din2(g41_n)
  );


  FA
  g_g42_n
  (
    .dout(g42_n),
    .din1(g40_p),
    .din2(g41_p)
  );


  LA
  g_g43_p
  (
    .dout(g43_p),
    .din1(g39_p),
    .din2(g42_p)
  );


  FA
  g_g43_n
  (
    .dout(g43_n),
    .din1(g39_n),
    .din2(g42_n)
  );


  LA
  g_g44_p
  (
    .dout(g44_p),
    .din1(G32_n_spl_),
    .din2(G34_p_spl_)
  );


  FA
  g_g44_n
  (
    .dout(g44_n),
    .din1(G32_p_spl_),
    .din2(G34_n_spl_)
  );


  LA
  g_g45_p
  (
    .dout(g45_p),
    .din1(G20_n_spl_),
    .din2(G22_p_spl_)
  );


  FA
  g_g45_n
  (
    .dout(g45_n),
    .din1(G20_p_spl_),
    .din2(G22_n_spl_)
  );


  LA
  g_g46_p
  (
    .dout(g46_p),
    .din1(g44_n),
    .din2(g45_n)
  );


  FA
  g_g46_n
  (
    .dout(g46_n),
    .din1(g44_p),
    .din2(g45_p)
  );


  LA
  g_g47_p
  (
    .dout(g47_p),
    .din1(G24_n_spl_),
    .din2(G26_p_spl_)
  );


  FA
  g_g47_n
  (
    .dout(g47_n),
    .din1(G24_p_spl_),
    .din2(G26_n_spl_)
  );


  LA
  g_g48_p
  (
    .dout(g48_p),
    .din1(G4_n_spl_),
    .din2(G6_p_spl_)
  );


  FA
  g_g48_n
  (
    .dout(g48_n),
    .din1(G4_p_spl_),
    .din2(G6_n_spl_)
  );


  LA
  g_g49_p
  (
    .dout(g49_p),
    .din1(G8_n_spl_),
    .din2(G10_p_spl_)
  );


  FA
  g_g49_n
  (
    .dout(g49_n),
    .din1(G8_p_spl_),
    .din2(G10_n_spl_)
  );


  LA
  g_g50_p
  (
    .dout(g50_p),
    .din1(g48_n),
    .din2(g49_n)
  );


  FA
  g_g50_n
  (
    .dout(g50_n),
    .din1(g48_p),
    .din2(g49_p)
  );


  LA
  g_g51_p
  (
    .dout(g51_p),
    .din1(g47_n),
    .din2(g50_p)
  );


  FA
  g_g51_n
  (
    .dout(g51_n),
    .din1(g47_p),
    .din2(g50_n)
  );


  LA
  g_g52_p
  (
    .dout(g52_p),
    .din1(g46_p),
    .din2(g51_p)
  );


  FA
  g_g52_n
  (
    .dout(g52_n),
    .din1(g46_n),
    .din2(g51_n)
  );


  LA
  g_g53_p
  (
    .dout(g53_p),
    .din1(g43_p),
    .din2(g52_p)
  );


  FA
  g_g53_n
  (
    .dout(g53_n),
    .din1(g43_n),
    .din2(g52_n)
  );


  LA
  g_g54_p
  (
    .dout(g54_p),
    .din1(G8_p_spl_),
    .din2(g53_n_spl_000)
  );


  FA
  g_g54_n
  (
    .dout(g54_n),
    .din1(G8_n_spl_),
    .din2(g53_p_spl_000)
  );


  LA
  g_g55_p
  (
    .dout(g55_p),
    .din1(G10_p_spl_),
    .din2(g54_n)
  );


  FA
  g_g55_n
  (
    .dout(g55_n),
    .din1(G10_n_spl_),
    .din2(g54_p)
  );


  LA
  g_g56_p
  (
    .dout(g56_p),
    .din1(G11_n_spl_),
    .din2(g55_p_spl_)
  );


  FA
  g_g56_n
  (
    .dout(g56_n),
    .din1(G11_p_spl_),
    .din2(g55_n_spl_)
  );


  LA
  g_g57_p
  (
    .dout(g57_p),
    .din1(G32_p_spl_),
    .din2(g53_n_spl_000)
  );


  FA
  g_g57_n
  (
    .dout(g57_n),
    .din1(G32_n_spl_),
    .din2(g53_p_spl_000)
  );


  LA
  g_g58_p
  (
    .dout(g58_p),
    .din1(G34_p_spl_),
    .din2(g57_n)
  );


  FA
  g_g58_n
  (
    .dout(g58_n),
    .din1(G34_n_spl_),
    .din2(g57_p)
  );


  LA
  g_g59_p
  (
    .dout(g59_p),
    .din1(G35_n_spl_),
    .din2(g58_p_spl_)
  );


  FA
  g_g59_n
  (
    .dout(g59_n),
    .din1(G35_p_spl_),
    .din2(g58_n_spl_)
  );


  LA
  g_g60_p
  (
    .dout(g60_p),
    .din1(g56_n),
    .din2(g59_n)
  );


  FA
  g_g60_n
  (
    .dout(g60_n),
    .din1(g56_p),
    .din2(g59_p)
  );


  LA
  g_g61_p
  (
    .dout(g61_p),
    .din1(G4_p_spl_),
    .din2(g53_n_spl_001)
  );


  FA
  g_g61_n
  (
    .dout(g61_n),
    .din1(G4_n_spl_),
    .din2(g53_p_spl_00)
  );


  LA
  g_g62_p
  (
    .dout(g62_p),
    .din1(G6_p_spl_),
    .din2(g61_n)
  );


  FA
  g_g62_n
  (
    .dout(g62_n),
    .din1(G6_n_spl_),
    .din2(g61_p)
  );


  LA
  g_g63_p
  (
    .dout(g63_p),
    .din1(G7_n_spl_),
    .din2(g62_p_spl_)
  );


  FA
  g_g63_n
  (
    .dout(g63_n),
    .din1(G7_p_spl_),
    .din2(g62_n_spl_)
  );


  LA
  g_g64_p
  (
    .dout(g64_p),
    .din1(G20_p_spl_),
    .din2(g53_n_spl_001)
  );


  FA
  g_g64_n
  (
    .dout(g64_n),
    .din1(G20_n_spl_),
    .din2(g53_p_spl_01)
  );


  LA
  g_g65_p
  (
    .dout(g65_p),
    .din1(G22_p_spl_),
    .din2(g64_n)
  );


  FA
  g_g65_n
  (
    .dout(g65_n),
    .din1(G22_n_spl_),
    .din2(g64_p)
  );


  LA
  g_g66_p
  (
    .dout(g66_p),
    .din1(G23_n_spl_),
    .din2(g65_p_spl_)
  );


  FA
  g_g66_n
  (
    .dout(g66_n),
    .din1(G23_p_spl_),
    .din2(g65_n_spl_)
  );


  LA
  g_g67_p
  (
    .dout(g67_p),
    .din1(g63_n),
    .din2(g66_n)
  );


  FA
  g_g67_n
  (
    .dout(g67_n),
    .din1(g63_p),
    .din2(g66_p)
  );


  LA
  g_g68_p
  (
    .dout(g68_p),
    .din1(g60_p),
    .din2(g67_p)
  );


  FA
  g_g68_n
  (
    .dout(g68_n),
    .din1(g60_n),
    .din2(g67_n)
  );


  LA
  g_g69_p
  (
    .dout(g69_p),
    .din1(G12_p_spl_),
    .din2(g53_n_spl_01)
  );


  FA
  g_g69_n
  (
    .dout(g69_n),
    .din1(G12_n_spl_),
    .din2(g53_p_spl_01)
  );


  LA
  g_g70_p
  (
    .dout(g70_p),
    .din1(G14_p_spl_),
    .din2(g69_n)
  );


  FA
  g_g70_n
  (
    .dout(g70_n),
    .din1(G14_n_spl_),
    .din2(g69_p)
  );


  LA
  g_g71_p
  (
    .dout(g71_p),
    .din1(G15_n_spl_),
    .din2(g70_p_spl_)
  );


  FA
  g_g71_n
  (
    .dout(g71_n),
    .din1(G15_p_spl_),
    .din2(g70_n_spl_)
  );


  LA
  g_g72_p
  (
    .dout(g72_p),
    .din1(G1_p_spl_),
    .din2(g53_n_spl_01)
  );


  FA
  g_g72_n
  (
    .dout(g72_n),
    .din1(G1_n_spl_),
    .din2(g53_p_spl_10)
  );


  LA
  g_g73_p
  (
    .dout(g73_p),
    .din1(G2_p_spl_),
    .din2(g72_n)
  );


  FA
  g_g73_n
  (
    .dout(g73_n),
    .din1(G2_n_spl_),
    .din2(g72_p)
  );


  LA
  g_g74_p
  (
    .dout(g74_p),
    .din1(G3_n_spl_),
    .din2(g73_p_spl_)
  );


  FA
  g_g74_n
  (
    .dout(g74_n),
    .din1(G3_p_spl_),
    .din2(g73_n_spl_)
  );


  LA
  g_g75_p
  (
    .dout(g75_p),
    .din1(g71_n),
    .din2(g74_n)
  );


  FA
  g_g75_n
  (
    .dout(g75_n),
    .din1(g71_p),
    .din2(g74_p)
  );


  LA
  g_g76_p
  (
    .dout(g76_p),
    .din1(G16_p_spl_),
    .din2(g53_n_spl_10)
  );


  FA
  g_g76_n
  (
    .dout(g76_n),
    .din1(G16_n_spl_),
    .din2(g53_p_spl_10)
  );


  LA
  g_g77_p
  (
    .dout(g77_p),
    .din1(G18_p_spl_),
    .din2(g76_n)
  );


  FA
  g_g77_n
  (
    .dout(g77_n),
    .din1(G18_n_spl_),
    .din2(g76_p)
  );


  LA
  g_g78_p
  (
    .dout(g78_p),
    .din1(G19_n_spl_),
    .din2(g77_p_spl_)
  );


  FA
  g_g78_n
  (
    .dout(g78_n),
    .din1(G19_p_spl_),
    .din2(g77_n_spl_)
  );


  LA
  g_g79_p
  (
    .dout(g79_p),
    .din1(G28_p_spl_),
    .din2(g53_n_spl_10)
  );


  FA
  g_g79_n
  (
    .dout(g79_n),
    .din1(G28_n_spl_),
    .din2(g53_p_spl_11)
  );


  LA
  g_g80_p
  (
    .dout(g80_p),
    .din1(G30_p_spl_),
    .din2(g79_n)
  );


  FA
  g_g80_n
  (
    .dout(g80_n),
    .din1(G30_n_spl_),
    .din2(g79_p)
  );


  LA
  g_g81_p
  (
    .dout(g81_p),
    .din1(G31_n_spl_),
    .din2(g80_p_spl_)
  );


  FA
  g_g81_n
  (
    .dout(g81_n),
    .din1(G31_p_spl_),
    .din2(g80_n_spl_)
  );


  LA
  g_g82_p
  (
    .dout(g82_p),
    .din1(G24_p_spl_),
    .din2(g53_n_spl_11)
  );


  FA
  g_g82_n
  (
    .dout(g82_n),
    .din1(G24_n_spl_),
    .din2(g53_p_spl_11)
  );


  LA
  g_g83_p
  (
    .dout(g83_p),
    .din1(G26_p_spl_),
    .din2(g82_n)
  );


  FA
  g_g83_n
  (
    .dout(g83_n),
    .din1(G26_n_spl_),
    .din2(g82_p)
  );


  LA
  g_g84_p
  (
    .dout(g84_p),
    .din1(G27_n_spl_),
    .din2(g83_p_spl_)
  );


  FA
  g_g84_n
  (
    .dout(g84_n),
    .din1(G27_p_spl_),
    .din2(g83_n_spl_)
  );


  LA
  g_g85_p
  (
    .dout(g85_p),
    .din1(g81_n),
    .din2(g84_n)
  );


  FA
  g_g85_n
  (
    .dout(g85_n),
    .din1(g81_p),
    .din2(g84_p)
  );


  LA
  g_g86_p
  (
    .dout(g86_p),
    .din1(g78_n),
    .din2(g85_p)
  );


  FA
  g_g86_n
  (
    .dout(g86_n),
    .din1(g78_p),
    .din2(g85_n)
  );


  LA
  g_g87_p
  (
    .dout(g87_p),
    .din1(g75_p),
    .din2(g86_p)
  );


  FA
  g_g87_n
  (
    .dout(g87_n),
    .din1(g75_n),
    .din2(g86_n)
  );


  LA
  g_g88_p
  (
    .dout(g88_p),
    .din1(g68_p),
    .din2(g87_p)
  );


  FA
  g_g88_n
  (
    .dout(g88_n),
    .din1(g68_n),
    .din2(g87_n)
  );


  LA
  g_g89_p
  (
    .dout(g89_p),
    .din1(G11_p_spl_),
    .din2(g88_n_spl_000)
  );


  FA
  g_g89_n
  (
    .dout(g89_n),
    .din1(G11_n_spl_),
    .din2(g88_p_spl_000)
  );


  LA
  g_g90_p
  (
    .dout(g90_p),
    .din1(g55_p_spl_),
    .din2(g89_n)
  );


  FA
  g_g90_n
  (
    .dout(g90_n),
    .din1(g55_n_spl_),
    .din2(g89_p)
  );


  LA
  g_g91_p
  (
    .dout(g91_p),
    .din1(G13_n_spl_),
    .din2(g90_p_spl_)
  );


  FA
  g_g91_n
  (
    .dout(g91_n),
    .din1(G13_p_spl_),
    .din2(g90_n_spl_)
  );


  LA
  g_g92_p
  (
    .dout(g92_p),
    .din1(G35_p_spl_),
    .din2(g88_n_spl_000)
  );


  FA
  g_g92_n
  (
    .dout(g92_n),
    .din1(G35_n_spl_),
    .din2(g88_p_spl_000)
  );


  LA
  g_g93_p
  (
    .dout(g93_p),
    .din1(g58_p_spl_),
    .din2(g92_n)
  );


  FA
  g_g93_n
  (
    .dout(g93_n),
    .din1(g58_n_spl_),
    .din2(g92_p)
  );


  LA
  g_g94_p
  (
    .dout(g94_p),
    .din1(G36_n),
    .din2(g93_p)
  );


  FA
  g_g94_n
  (
    .dout(g94_n),
    .din1(G36_p_spl_),
    .din2(g93_n_spl_)
  );


  LA
  g_g95_p
  (
    .dout(g95_p),
    .din1(g91_n),
    .din2(g94_n)
  );


  FA
  g_g95_n
  (
    .dout(g95_n),
    .din1(g91_p),
    .din2(g94_p)
  );


  LA
  g_g96_p
  (
    .dout(g96_p),
    .din1(G7_p_spl_),
    .din2(g88_n_spl_001)
  );


  FA
  g_g96_n
  (
    .dout(g96_n),
    .din1(G7_n_spl_),
    .din2(g88_p_spl_00)
  );


  LA
  g_g97_p
  (
    .dout(g97_p),
    .din1(g62_p_spl_),
    .din2(g96_n)
  );


  FA
  g_g97_n
  (
    .dout(g97_n),
    .din1(g62_n_spl_),
    .din2(g96_p)
  );


  LA
  g_g98_p
  (
    .dout(g98_p),
    .din1(G9_n),
    .din2(g97_p)
  );


  FA
  g_g98_n
  (
    .dout(g98_n),
    .din1(G9_p_spl_),
    .din2(g97_n_spl_)
  );


  LA
  g_g99_p
  (
    .dout(g99_p),
    .din1(G23_p_spl_),
    .din2(g88_n_spl_001)
  );


  FA
  g_g99_n
  (
    .dout(g99_n),
    .din1(G23_n_spl_),
    .din2(g88_p_spl_01)
  );


  LA
  g_g100_p
  (
    .dout(g100_p),
    .din1(g65_p_spl_),
    .din2(g99_n)
  );


  FA
  g_g100_n
  (
    .dout(g100_n),
    .din1(g65_n_spl_),
    .din2(g99_p)
  );


  LA
  g_g101_p
  (
    .dout(g101_p),
    .din1(G25_n),
    .din2(g100_p)
  );


  FA
  g_g101_n
  (
    .dout(g101_n),
    .din1(G25_p_spl_),
    .din2(g100_n_spl_)
  );


  LA
  g_g102_p
  (
    .dout(g102_p),
    .din1(g98_n),
    .din2(g101_n)
  );


  FA
  g_g102_n
  (
    .dout(g102_n),
    .din1(g98_p),
    .din2(g101_p)
  );


  LA
  g_g103_p
  (
    .dout(g103_p),
    .din1(g95_p),
    .din2(g102_p)
  );


  FA
  g_g103_n
  (
    .dout(g103_n),
    .din1(g95_n),
    .din2(g102_n)
  );


  LA
  g_g104_p
  (
    .dout(g104_p),
    .din1(G15_p_spl_),
    .din2(g88_n_spl_01)
  );


  FA
  g_g104_n
  (
    .dout(g104_n),
    .din1(G15_n_spl_),
    .din2(g88_p_spl_01)
  );


  LA
  g_g105_p
  (
    .dout(g105_p),
    .din1(g70_p_spl_),
    .din2(g104_n)
  );


  FA
  g_g105_n
  (
    .dout(g105_n),
    .din1(g70_n_spl_),
    .din2(g104_p)
  );


  LA
  g_g106_p
  (
    .dout(g106_p),
    .din1(G17_n_spl_),
    .din2(g105_p_spl_)
  );


  FA
  g_g106_n
  (
    .dout(g106_n),
    .din1(G17_p_spl_),
    .din2(g105_n_spl_)
  );


  LA
  g_g107_p
  (
    .dout(g107_p),
    .din1(G3_p_spl_),
    .din2(g88_n_spl_01)
  );


  FA
  g_g107_n
  (
    .dout(g107_n),
    .din1(G3_n_spl_),
    .din2(g88_p_spl_10)
  );


  LA
  g_g108_p
  (
    .dout(g108_p),
    .din1(g73_p_spl_),
    .din2(g107_n)
  );


  FA
  g_g108_n
  (
    .dout(g108_n),
    .din1(g73_n_spl_),
    .din2(g107_p)
  );


  LA
  g_g109_p
  (
    .dout(g109_p),
    .din1(G5_n_spl_),
    .din2(g108_p_spl_)
  );


  FA
  g_g109_n
  (
    .dout(g109_n),
    .din1(G5_p),
    .din2(g108_n)
  );


  LA
  g_g110_p
  (
    .dout(g110_p),
    .din1(g106_n),
    .din2(g109_n)
  );


  FA
  g_g110_n
  (
    .dout(g110_n),
    .din1(g106_p),
    .din2(g109_p)
  );


  LA
  g_g111_p
  (
    .dout(g111_p),
    .din1(G19_p_spl_),
    .din2(g88_n_spl_10)
  );


  FA
  g_g111_n
  (
    .dout(g111_n),
    .din1(G19_n_spl_),
    .din2(g88_p_spl_10)
  );


  LA
  g_g112_p
  (
    .dout(g112_p),
    .din1(g77_p_spl_),
    .din2(g111_n)
  );


  FA
  g_g112_n
  (
    .dout(g112_n),
    .din1(g77_n_spl_),
    .din2(g111_p)
  );


  LA
  g_g113_p
  (
    .dout(g113_p),
    .din1(G21_n_spl_),
    .din2(g112_p_spl_)
  );


  FA
  g_g113_n
  (
    .dout(g113_n),
    .din1(G21_p_spl_),
    .din2(g112_n_spl_)
  );


  LA
  g_g114_p
  (
    .dout(g114_p),
    .din1(G31_p_spl_),
    .din2(g88_n_spl_10)
  );


  FA
  g_g114_n
  (
    .dout(g114_n),
    .din1(G31_n_spl_),
    .din2(g88_p_spl_11)
  );


  LA
  g_g115_p
  (
    .dout(g115_p),
    .din1(g80_p_spl_),
    .din2(g114_n)
  );


  FA
  g_g115_n
  (
    .dout(g115_n),
    .din1(g80_n_spl_),
    .din2(g114_p)
  );


  LA
  g_g116_p
  (
    .dout(g116_p),
    .din1(G33_n),
    .din2(g115_p)
  );


  FA
  g_g116_n
  (
    .dout(g116_n),
    .din1(G33_p_spl_),
    .din2(g115_n_spl_)
  );


  LA
  g_g117_p
  (
    .dout(g117_p),
    .din1(G27_p_spl_),
    .din2(g88_n_spl_11)
  );


  FA
  g_g117_n
  (
    .dout(g117_n),
    .din1(G27_n_spl_),
    .din2(g88_p_spl_11)
  );


  LA
  g_g118_p
  (
    .dout(g118_p),
    .din1(g83_p_spl_),
    .din2(g117_n)
  );


  FA
  g_g118_n
  (
    .dout(g118_n),
    .din1(g83_n_spl_),
    .din2(g117_p)
  );


  LA
  g_g119_p
  (
    .dout(g119_p),
    .din1(G29_n_spl_),
    .din2(g118_p_spl_)
  );


  FA
  g_g119_n
  (
    .dout(g119_n),
    .din1(G29_p_spl_),
    .din2(g118_n_spl_)
  );


  LA
  g_g120_p
  (
    .dout(g120_p),
    .din1(g116_n),
    .din2(g119_n)
  );


  FA
  g_g120_n
  (
    .dout(g120_n),
    .din1(g116_p),
    .din2(g119_p)
  );


  LA
  g_g121_p
  (
    .dout(g121_p),
    .din1(g113_n),
    .din2(g120_p)
  );


  FA
  g_g121_n
  (
    .dout(g121_n),
    .din1(g113_p),
    .din2(g120_n)
  );


  LA
  g_g122_p
  (
    .dout(g122_p),
    .din1(g110_p),
    .din2(g121_p)
  );


  FA
  g_g122_n
  (
    .dout(g122_n),
    .din1(g110_n),
    .din2(g121_n)
  );


  LA
  g_g123_p
  (
    .dout(g123_p),
    .din1(g103_p),
    .din2(g122_p)
  );


  FA
  g_g123_n
  (
    .dout(g123_n),
    .din1(g103_n),
    .din2(g122_n)
  );


  FA
  g_g124_n
  (
    .dout(g124_n),
    .din1(G5_n_spl_),
    .din2(g123_p_spl_00)
  );


  LA
  g_g125_p
  (
    .dout(g125_p),
    .din1(g108_p_spl_),
    .din2(g124_n)
  );


  LA
  g_g126_p
  (
    .dout(g126_p),
    .din1(G29_p_spl_),
    .din2(g123_n_spl_000)
  );


  FA
  g_g126_n
  (
    .dout(g126_n),
    .din1(G29_n_spl_),
    .din2(g123_p_spl_00)
  );


  LA
  g_g127_p
  (
    .dout(g127_p),
    .din1(g118_p_spl_),
    .din2(g126_n)
  );


  FA
  g_g127_n
  (
    .dout(g127_n),
    .din1(g118_n_spl_),
    .din2(g126_p)
  );


  LA
  g_g128_p
  (
    .dout(g128_p),
    .din1(G25_p_spl_),
    .din2(g123_n_spl_000)
  );


  FA
  g_g129_n
  (
    .dout(g129_n),
    .din1(g100_n_spl_),
    .din2(g128_p)
  );


  LA
  g_g130_p
  (
    .dout(g130_p),
    .din1(G9_p_spl_),
    .din2(g123_n_spl_00)
  );


  FA
  g_g131_n
  (
    .dout(g131_n),
    .din1(g97_n_spl_),
    .din2(g130_p)
  );


  LA
  g_g132_p
  (
    .dout(g132_p),
    .din1(G13_p_spl_),
    .din2(g123_n_spl_01)
  );


  FA
  g_g132_n
  (
    .dout(g132_n),
    .din1(G13_n_spl_),
    .din2(g123_p_spl_0)
  );


  LA
  g_g133_p
  (
    .dout(g133_p),
    .din1(g90_p_spl_),
    .din2(g132_n)
  );


  FA
  g_g133_n
  (
    .dout(g133_n),
    .din1(g90_n_spl_),
    .din2(g132_p)
  );


  LA
  g_g134_p
  (
    .dout(g134_p),
    .din1(g131_n_spl_),
    .din2(g133_n)
  );


  LA
  g_g135_p
  (
    .dout(g135_p),
    .din1(G21_p_spl_),
    .din2(g123_n_spl_01)
  );


  FA
  g_g135_n
  (
    .dout(g135_n),
    .din1(G21_n_spl_),
    .din2(g123_p_spl_1)
  );


  LA
  g_g136_p
  (
    .dout(g136_p),
    .din1(g112_p_spl_),
    .din2(g135_n)
  );


  FA
  g_g136_n
  (
    .dout(g136_n),
    .din1(g112_n_spl_),
    .din2(g135_p)
  );


  LA
  g_g137_p
  (
    .dout(g137_p),
    .din1(G17_p_spl_),
    .din2(g123_n_spl_10)
  );


  FA
  g_g137_n
  (
    .dout(g137_n),
    .din1(G17_n_spl_),
    .din2(g123_p_spl_1)
  );


  LA
  g_g138_p
  (
    .dout(g138_p),
    .din1(g105_p_spl_),
    .din2(g137_n)
  );


  FA
  g_g138_n
  (
    .dout(g138_n),
    .din1(g105_n_spl_),
    .din2(g137_p)
  );


  LA
  g_g139_p
  (
    .dout(g139_p),
    .din1(g136_n),
    .din2(g138_n_spl_)
  );


  FA
  g_g139_n
  (
    .dout(g139_n),
    .din1(g136_p_spl_),
    .din2(g138_p_spl_)
  );


  LA
  g_g140_p
  (
    .dout(g140_p),
    .din1(g134_p_spl_),
    .din2(g139_p)
  );


  LA
  g_g141_p
  (
    .dout(g141_p),
    .din1(G36_p_spl_),
    .din2(g123_n_spl_10)
  );


  FA
  g_g142_n
  (
    .dout(g142_n),
    .din1(g93_n_spl_),
    .din2(g141_p)
  );


  LA
  g_g143_p
  (
    .dout(g143_p),
    .din1(G33_p_spl_),
    .din2(g123_n_spl_11)
  );


  FA
  g_g144_n
  (
    .dout(g144_n),
    .din1(g115_n_spl_),
    .din2(g143_p)
  );


  LA
  g_g145_p
  (
    .dout(g145_p),
    .din1(g142_n),
    .din2(g144_n_spl_)
  );


  LA
  g_g146_p
  (
    .dout(g146_p),
    .din1(g140_p_spl_),
    .din2(g145_p)
  );


  LA
  g_g147_p
  (
    .dout(g147_p),
    .din1(g129_n_spl_),
    .din2(g146_p)
  );


  LA
  g_g148_p
  (
    .dout(g148_p),
    .din1(g127_n_spl_),
    .din2(g147_p)
  );


  FA
  g_g149_n
  (
    .dout(g149_n),
    .din1(g125_p),
    .din2(g148_p)
  );


  FA
  g_g150_n
  (
    .dout(g150_n),
    .din1(g127_n_spl_),
    .din2(g139_n)
  );


  FA
  g_g151_n
  (
    .dout(g151_n),
    .din1(g133_p_spl_),
    .din2(g138_p_spl_)
  );


  FA
  g_g152_n
  (
    .dout(g152_n),
    .din1(g136_p_spl_),
    .din2(g151_n)
  );


  FA
  g_g153_n
  (
    .dout(g153_n),
    .din1(g129_n_spl_),
    .din2(g152_n)
  );


  LA
  g_g154_p
  (
    .dout(g154_p),
    .din1(g134_p_spl_),
    .din2(g153_n_spl_)
  );


  LA
  g_g155_p
  (
    .dout(g155_p),
    .din1(g150_n),
    .din2(g154_p)
  );


  FA
  g_g156_n
  (
    .dout(g156_n),
    .din1(g127_p),
    .din2(g144_n_spl_)
  );


  LA
  g_g157_p
  (
    .dout(g157_p),
    .din1(g138_n_spl_),
    .din2(g156_n)
  );


  FA
  g_g158_n
  (
    .dout(g158_n),
    .din1(g133_p_spl_),
    .din2(g157_p)
  );


  LA
  g_g159_p
  (
    .dout(g159_p),
    .din1(g153_n_spl_),
    .din2(g158_n)
  );


  LA
  g_g160_p
  (
    .dout(g160_p),
    .din1(g131_n_spl_),
    .din2(g159_p)
  );


  buf

  (
    G426_p,
    g53_n_spl_11
  );


  buf

  (
    G427_p,
    g88_n_spl_11
  );


  buf

  (
    G428_p,
    g123_n_spl_11
  );


  buf

  (
    G429_n,
    g149_n
  );


  buf

  (
    G430_n,
    g140_p_spl_
  );


  buf

  (
    G431_n,
    g155_p
  );


  buf

  (
    G432_n,
    g160_p
  );


  buf

  (
    G16_n_spl_,
    G16_n
  );


  buf

  (
    G18_p_spl_,
    G18_p
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    G18_n_spl_,
    G18_n
  );


  buf

  (
    G12_n_spl_,
    G12_n
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G14_n_spl_,
    G14_n
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G28_n_spl_,
    G28_n
  );


  buf

  (
    G30_p_spl_,
    G30_p
  );


  buf

  (
    G28_p_spl_,
    G28_p
  );


  buf

  (
    G30_n_spl_,
    G30_n
  );


  buf

  (
    G32_n_spl_,
    G32_n
  );


  buf

  (
    G34_p_spl_,
    G34_p
  );


  buf

  (
    G32_p_spl_,
    G32_p
  );


  buf

  (
    G34_n_spl_,
    G34_n
  );


  buf

  (
    G20_n_spl_,
    G20_n
  );


  buf

  (
    G22_p_spl_,
    G22_p
  );


  buf

  (
    G20_p_spl_,
    G20_p
  );


  buf

  (
    G22_n_spl_,
    G22_n
  );


  buf

  (
    G24_n_spl_,
    G24_n
  );


  buf

  (
    G26_p_spl_,
    G26_p
  );


  buf

  (
    G24_p_spl_,
    G24_p
  );


  buf

  (
    G26_n_spl_,
    G26_n
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G6_n_spl_,
    G6_n
  );


  buf

  (
    G8_n_spl_,
    G8_n
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G10_n_spl_,
    G10_n
  );


  buf

  (
    g53_n_spl_,
    g53_n
  );


  buf

  (
    g53_n_spl_0,
    g53_n_spl_
  );


  buf

  (
    g53_n_spl_00,
    g53_n_spl_0
  );


  buf

  (
    g53_n_spl_000,
    g53_n_spl_00
  );


  buf

  (
    g53_n_spl_001,
    g53_n_spl_00
  );


  buf

  (
    g53_n_spl_01,
    g53_n_spl_0
  );


  buf

  (
    g53_n_spl_1,
    g53_n_spl_
  );


  buf

  (
    g53_n_spl_10,
    g53_n_spl_1
  );


  buf

  (
    g53_n_spl_11,
    g53_n_spl_1
  );


  buf

  (
    g53_p_spl_,
    g53_p
  );


  buf

  (
    g53_p_spl_0,
    g53_p_spl_
  );


  buf

  (
    g53_p_spl_00,
    g53_p_spl_0
  );


  buf

  (
    g53_p_spl_000,
    g53_p_spl_00
  );


  buf

  (
    g53_p_spl_01,
    g53_p_spl_0
  );


  buf

  (
    g53_p_spl_1,
    g53_p_spl_
  );


  buf

  (
    g53_p_spl_10,
    g53_p_spl_1
  );


  buf

  (
    g53_p_spl_11,
    g53_p_spl_1
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    g55_p_spl_,
    g55_p
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    g55_n_spl_,
    g55_n
  );


  buf

  (
    G35_n_spl_,
    G35_n
  );


  buf

  (
    g58_p_spl_,
    g58_p
  );


  buf

  (
    G35_p_spl_,
    G35_p
  );


  buf

  (
    g58_n_spl_,
    g58_n
  );


  buf

  (
    G7_n_spl_,
    G7_n
  );


  buf

  (
    g62_p_spl_,
    g62_p
  );


  buf

  (
    G7_p_spl_,
    G7_p
  );


  buf

  (
    g62_n_spl_,
    g62_n
  );


  buf

  (
    G23_n_spl_,
    G23_n
  );


  buf

  (
    g65_p_spl_,
    g65_p
  );


  buf

  (
    G23_p_spl_,
    G23_p
  );


  buf

  (
    g65_n_spl_,
    g65_n
  );


  buf

  (
    G15_n_spl_,
    G15_n
  );


  buf

  (
    g70_p_spl_,
    g70_p
  );


  buf

  (
    G15_p_spl_,
    G15_p
  );


  buf

  (
    g70_n_spl_,
    g70_n
  );


  buf

  (
    G3_n_spl_,
    G3_n
  );


  buf

  (
    g73_p_spl_,
    g73_p
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    g73_n_spl_,
    g73_n
  );


  buf

  (
    G19_n_spl_,
    G19_n
  );


  buf

  (
    g77_p_spl_,
    g77_p
  );


  buf

  (
    G19_p_spl_,
    G19_p
  );


  buf

  (
    g77_n_spl_,
    g77_n
  );


  buf

  (
    G31_n_spl_,
    G31_n
  );


  buf

  (
    g80_p_spl_,
    g80_p
  );


  buf

  (
    G31_p_spl_,
    G31_p
  );


  buf

  (
    g80_n_spl_,
    g80_n
  );


  buf

  (
    G27_n_spl_,
    G27_n
  );


  buf

  (
    g83_p_spl_,
    g83_p
  );


  buf

  (
    G27_p_spl_,
    G27_p
  );


  buf

  (
    g83_n_spl_,
    g83_n
  );


  buf

  (
    g88_n_spl_,
    g88_n
  );


  buf

  (
    g88_n_spl_0,
    g88_n_spl_
  );


  buf

  (
    g88_n_spl_00,
    g88_n_spl_0
  );


  buf

  (
    g88_n_spl_000,
    g88_n_spl_00
  );


  buf

  (
    g88_n_spl_001,
    g88_n_spl_00
  );


  buf

  (
    g88_n_spl_01,
    g88_n_spl_0
  );


  buf

  (
    g88_n_spl_1,
    g88_n_spl_
  );


  buf

  (
    g88_n_spl_10,
    g88_n_spl_1
  );


  buf

  (
    g88_n_spl_11,
    g88_n_spl_1
  );


  buf

  (
    g88_p_spl_,
    g88_p
  );


  buf

  (
    g88_p_spl_0,
    g88_p_spl_
  );


  buf

  (
    g88_p_spl_00,
    g88_p_spl_0
  );


  buf

  (
    g88_p_spl_000,
    g88_p_spl_00
  );


  buf

  (
    g88_p_spl_01,
    g88_p_spl_0
  );


  buf

  (
    g88_p_spl_1,
    g88_p_spl_
  );


  buf

  (
    g88_p_spl_10,
    g88_p_spl_1
  );


  buf

  (
    g88_p_spl_11,
    g88_p_spl_1
  );


  buf

  (
    G13_n_spl_,
    G13_n
  );


  buf

  (
    g90_p_spl_,
    g90_p
  );


  buf

  (
    G13_p_spl_,
    G13_p
  );


  buf

  (
    g90_n_spl_,
    g90_n
  );


  buf

  (
    G36_p_spl_,
    G36_p
  );


  buf

  (
    g93_n_spl_,
    g93_n
  );


  buf

  (
    G9_p_spl_,
    G9_p
  );


  buf

  (
    g97_n_spl_,
    g97_n
  );


  buf

  (
    G25_p_spl_,
    G25_p
  );


  buf

  (
    g100_n_spl_,
    g100_n
  );


  buf

  (
    G17_n_spl_,
    G17_n
  );


  buf

  (
    g105_p_spl_,
    g105_p
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    g105_n_spl_,
    g105_n
  );


  buf

  (
    G5_n_spl_,
    G5_n
  );


  buf

  (
    g108_p_spl_,
    g108_p
  );


  buf

  (
    G21_n_spl_,
    G21_n
  );


  buf

  (
    g112_p_spl_,
    g112_p
  );


  buf

  (
    G21_p_spl_,
    G21_p
  );


  buf

  (
    g112_n_spl_,
    g112_n
  );


  buf

  (
    G33_p_spl_,
    G33_p
  );


  buf

  (
    g115_n_spl_,
    g115_n
  );


  buf

  (
    G29_n_spl_,
    G29_n
  );


  buf

  (
    g118_p_spl_,
    g118_p
  );


  buf

  (
    G29_p_spl_,
    G29_p
  );


  buf

  (
    g118_n_spl_,
    g118_n
  );


  buf

  (
    g123_p_spl_,
    g123_p
  );


  buf

  (
    g123_p_spl_0,
    g123_p_spl_
  );


  buf

  (
    g123_p_spl_00,
    g123_p_spl_0
  );


  buf

  (
    g123_p_spl_1,
    g123_p_spl_
  );


  buf

  (
    g123_n_spl_,
    g123_n
  );


  buf

  (
    g123_n_spl_0,
    g123_n_spl_
  );


  buf

  (
    g123_n_spl_00,
    g123_n_spl_0
  );


  buf

  (
    g123_n_spl_000,
    g123_n_spl_00
  );


  buf

  (
    g123_n_spl_01,
    g123_n_spl_0
  );


  buf

  (
    g123_n_spl_1,
    g123_n_spl_
  );


  buf

  (
    g123_n_spl_10,
    g123_n_spl_1
  );


  buf

  (
    g123_n_spl_11,
    g123_n_spl_1
  );


  buf

  (
    g131_n_spl_,
    g131_n
  );


  buf

  (
    g138_n_spl_,
    g138_n
  );


  buf

  (
    g136_p_spl_,
    g136_p
  );


  buf

  (
    g138_p_spl_,
    g138_p
  );


  buf

  (
    g134_p_spl_,
    g134_p
  );


  buf

  (
    g144_n_spl_,
    g144_n
  );


  buf

  (
    g140_p_spl_,
    g140_p
  );


  buf

  (
    g129_n_spl_,
    g129_n
  );


  buf

  (
    g127_n_spl_,
    g127_n
  );


  buf

  (
    g133_p_spl_,
    g133_p
  );


  buf

  (
    g153_n_spl_,
    g153_n
  );


endmodule
