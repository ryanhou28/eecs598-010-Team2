// Benchmark "mymod" written by ABC on Sun Oct 29 19:31:48 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41,
    G468, G469, G470, G471, G472, G473, G474, G475, G476, G477, G478, G479,
    G480, G481, G482, G483, G484, G485, G486, G487, G488, G489, G490, G491,
    G492, G493, G494, G495, G496, G497, G498, G499  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41;
  output G468, G469, G470, G471, G472, G473, G474, G475, G476, G477, G478,
    G479, G480, G481, G482, G483, G484, G485, G486, G487, G488, G489, G490,
    G491, G492, G493, G494, G495, G496, G497, G498, G499;
  reg n286_lo, n298_lo, n310_lo, n322_lo, n334_lo, n346_lo, n358_lo,
    n370_lo, n382_lo, n394_lo, n406_lo, n418_lo, n430_lo, n442_lo, n454_lo,
    n466_lo, n478_lo, n490_lo, n502_lo, n514_lo, n526_lo, n538_lo, n550_lo,
    n562_lo, n574_lo, n586_lo, n598_lo, n610_lo, n622_lo, n634_lo, n646_lo,
    n658_lo, n661_lo, n673_lo, n685_lo, n697_lo, n709_lo, n721_lo, n733_lo,
    n745_lo, n757_lo, n1248_o2, n1249_o2, n1250_o2, n1251_o2, n1252_o2,
    n1253_o2, n1254_o2, n1255_o2, n1207_o2, n1208_o2, n1209_o2, n1210_o2,
    n1211_o2, n1212_o2, n1213_o2, n1214_o2, n1215_o2, n1216_o2, n1217_o2,
    n1218_o2, n1219_o2, n1220_o2, n1221_o2, n1222_o2, n1223_o2, n1224_o2,
    n1225_o2, n1226_o2, n1227_o2, n1228_o2, n1229_o2, n1230_o2, n1231_o2,
    n1232_o2, n1233_o2, n1234_o2, n1235_o2, n1236_o2, n1237_o2, n1238_o2,
    G374_o2, G376_o2, G370_o2, G372_o2, G373_o2, G377_o2, G371_o2, G375_o2,
    G354_o2, G356_o2, G350_o2, G352_o2, G353_o2, G357_o2, G351_o2, G355_o2,
    G386_o2, G391_o2, n283_lo_buf_o2, n295_lo_buf_o2, n307_lo_buf_o2,
    n319_lo_buf_o2, n331_lo_buf_o2, n343_lo_buf_o2, n355_lo_buf_o2,
    n367_lo_buf_o2, n379_lo_buf_o2, n391_lo_buf_o2, n403_lo_buf_o2,
    n415_lo_buf_o2, n427_lo_buf_o2, n439_lo_buf_o2, n451_lo_buf_o2,
    n463_lo_buf_o2, n475_lo_buf_o2, n487_lo_buf_o2, n499_lo_buf_o2,
    n511_lo_buf_o2, n523_lo_buf_o2, n535_lo_buf_o2, n547_lo_buf_o2,
    n559_lo_buf_o2, n571_lo_buf_o2, n583_lo_buf_o2, n595_lo_buf_o2,
    n607_lo_buf_o2, n619_lo_buf_o2, n631_lo_buf_o2, n643_lo_buf_o2,
    n655_lo_buf_o2, G234_o2, G247_o2, G260_o2, G273_o2, G286_o2, G299_o2,
    G312_o2, G325_o2, n667_lo_buf_o2, n679_lo_buf_o2, n691_lo_buf_o2,
    n703_lo_buf_o2, n715_lo_buf_o2, n727_lo_buf_o2, n739_lo_buf_o2,
    n751_lo_buf_o2, n763_lo_buf_o2, G186_o2, G189_o2, G192_o2, G195_o2,
    G198_o2, G201_o2, G204_o2, G207_o2, n280_lo_buf_o2, n292_lo_buf_o2,
    n304_lo_buf_o2, n316_lo_buf_o2, n328_lo_buf_o2, n340_lo_buf_o2,
    n352_lo_buf_o2, n364_lo_buf_o2, n376_lo_buf_o2, n388_lo_buf_o2,
    n400_lo_buf_o2, n412_lo_buf_o2, n424_lo_buf_o2, n436_lo_buf_o2,
    n448_lo_buf_o2, n460_lo_buf_o2, n472_lo_buf_o2, n484_lo_buf_o2,
    n496_lo_buf_o2, n508_lo_buf_o2, n520_lo_buf_o2, n532_lo_buf_o2,
    n544_lo_buf_o2, n556_lo_buf_o2, n568_lo_buf_o2, n580_lo_buf_o2,
    n592_lo_buf_o2, n604_lo_buf_o2, n616_lo_buf_o2, n628_lo_buf_o2,
    n640_lo_buf_o2, n652_lo_buf_o2;
  wire new_n451_, new_n453_, new_n455_, new_n457_, new_n459_, new_n461_,
    new_n463_, new_n465_, new_n467_, new_n469_, new_n471_, new_n473_,
    new_n475_, new_n477_, new_n479_, new_n481_, new_n483_, new_n485_,
    new_n487_, new_n489_, new_n491_, new_n493_, new_n495_, new_n497_,
    new_n499_, new_n501_, new_n503_, new_n505_, new_n507_, new_n509_,
    new_n511_, new_n513_, new_n515_, new_n517_, new_n519_, new_n521_,
    new_n523_, new_n525_, new_n527_, new_n529_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n597_, new_n599_, new_n601_,
    new_n603_, new_n605_, new_n607_, new_n609_, new_n611_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n631_, new_n633_,
    new_n635_, new_n637_, new_n639_, new_n641_, new_n643_, new_n645_,
    new_n647_, new_n649_, new_n651_, new_n653_, new_n655_, new_n657_,
    new_n659_, new_n661_, new_n663_, new_n665_, new_n667_, new_n669_,
    new_n671_, new_n673_, new_n675_, new_n677_, new_n679_, new_n681_,
    new_n683_, new_n685_, new_n687_, new_n689_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_,
    new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_,
    new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_,
    new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_,
    new_n1558_, new_n1559_, new_n1780_, new_n1781_, new_n1782_, new_n1783_,
    new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_,
    new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_,
    new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_,
    new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_,
    new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_,
    new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_,
    new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_,
    new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_,
    new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_,
    new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_,
    new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_,
    new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_,
    new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_,
    new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_,
    new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_,
    new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_,
    new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_,
    new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_,
    new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_,
    new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_,
    new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_,
    new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_,
    new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_,
    new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_,
    new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_,
    new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_,
    new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_,
    new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_,
    new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_,
    new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_,
    new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_,
    new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_,
    new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_,
    new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_,
    new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_,
    new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_,
    new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_,
    new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_,
    new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_,
    new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_,
    new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_,
    new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_,
    new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_,
    new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_,
    new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_,
    new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_,
    new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_,
    new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_,
    new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_,
    new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_,
    new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_,
    new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_,
    new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_,
    new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_,
    new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_,
    new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_,
    new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_,
    new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_,
    new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_,
    new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_,
    new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_,
    new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_,
    new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_,
    new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_,
    new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_,
    new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_,
    new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_,
    new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_,
    new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_,
    new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_,
    new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_,
    new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_,
    new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_,
    new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_,
    new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_,
    new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_,
    n286_li, n298_li, n310_li, n322_li, n334_li, n346_li, n358_li, n370_li,
    n382_li, n394_li, n406_li, n418_li, n430_li, n442_li, n454_li, n466_li,
    n478_li, n490_li, n502_li, n514_li, n526_li, n538_li, n550_li, n562_li,
    n574_li, n586_li, n598_li, n610_li, n622_li, n634_li, n646_li, n658_li,
    n661_li, n673_li, n685_li, n697_li, n709_li, n721_li, n733_li, n745_li,
    n757_li, n1248_i2, n1249_i2, n1250_i2, n1251_i2, n1252_i2, n1253_i2,
    n1254_i2, n1255_i2, n1207_i2, n1208_i2, n1209_i2, n1210_i2, n1211_i2,
    n1212_i2, n1213_i2, n1214_i2, n1215_i2, n1216_i2, n1217_i2, n1218_i2,
    n1219_i2, n1220_i2, n1221_i2, n1222_i2, n1223_i2, n1224_i2, n1225_i2,
    n1226_i2, n1227_i2, n1228_i2, n1229_i2, n1230_i2, n1231_i2, n1232_i2,
    n1233_i2, n1234_i2, n1235_i2, n1236_i2, n1237_i2, n1238_i2, G374_i2,
    G376_i2, G370_i2, G372_i2, G373_i2, G377_i2, G371_i2, G375_i2, G354_i2,
    G356_i2, G350_i2, G352_i2, G353_i2, G357_i2, G351_i2, G355_i2, G386_i2,
    G391_i2, n283_lo_buf_i2, n295_lo_buf_i2, n307_lo_buf_i2,
    n319_lo_buf_i2, n331_lo_buf_i2, n343_lo_buf_i2, n355_lo_buf_i2,
    n367_lo_buf_i2, n379_lo_buf_i2, n391_lo_buf_i2, n403_lo_buf_i2,
    n415_lo_buf_i2, n427_lo_buf_i2, n439_lo_buf_i2, n451_lo_buf_i2,
    n463_lo_buf_i2, n475_lo_buf_i2, n487_lo_buf_i2, n499_lo_buf_i2,
    n511_lo_buf_i2, n523_lo_buf_i2, n535_lo_buf_i2, n547_lo_buf_i2,
    n559_lo_buf_i2, n571_lo_buf_i2, n583_lo_buf_i2, n595_lo_buf_i2,
    n607_lo_buf_i2, n619_lo_buf_i2, n631_lo_buf_i2, n643_lo_buf_i2,
    n655_lo_buf_i2, G234_i2, G247_i2, G260_i2, G273_i2, G286_i2, G299_i2,
    G312_i2, G325_i2, n667_lo_buf_i2, n679_lo_buf_i2, n691_lo_buf_i2,
    n703_lo_buf_i2, n715_lo_buf_i2, n727_lo_buf_i2, n739_lo_buf_i2,
    n751_lo_buf_i2, n763_lo_buf_i2, G186_i2, G189_i2, G192_i2, G195_i2,
    G198_i2, G201_i2, G204_i2, G207_i2, n280_lo_buf_i2, n292_lo_buf_i2,
    n304_lo_buf_i2, n316_lo_buf_i2, n328_lo_buf_i2, n340_lo_buf_i2,
    n352_lo_buf_i2, n364_lo_buf_i2, n376_lo_buf_i2, n388_lo_buf_i2,
    n400_lo_buf_i2, n412_lo_buf_i2, n424_lo_buf_i2, n436_lo_buf_i2,
    n448_lo_buf_i2, n460_lo_buf_i2, n472_lo_buf_i2, n484_lo_buf_i2,
    n496_lo_buf_i2, n508_lo_buf_i2, n520_lo_buf_i2, n532_lo_buf_i2,
    n544_lo_buf_i2, n556_lo_buf_i2, n568_lo_buf_i2, n580_lo_buf_i2,
    n592_lo_buf_i2, n604_lo_buf_i2, n616_lo_buf_i2, n628_lo_buf_i2,
    n640_lo_buf_i2, n652_lo_buf_i2;
  assign new_n451_ = ~G1;
  assign new_n453_ = ~G2;
  assign new_n455_ = ~G3;
  assign new_n457_ = ~G4;
  assign new_n459_ = ~G5;
  assign new_n461_ = ~G6;
  assign new_n463_ = ~G7;
  assign new_n465_ = ~G8;
  assign new_n467_ = ~G9;
  assign new_n469_ = ~G10;
  assign new_n471_ = ~G11;
  assign new_n473_ = ~G12;
  assign new_n475_ = ~G13;
  assign new_n477_ = ~G14;
  assign new_n479_ = ~G15;
  assign new_n481_ = ~G16;
  assign new_n483_ = ~G17;
  assign new_n485_ = ~G18;
  assign new_n487_ = ~G19;
  assign new_n489_ = ~G20;
  assign new_n491_ = ~G21;
  assign new_n493_ = ~G22;
  assign new_n495_ = ~G23;
  assign new_n497_ = ~G24;
  assign new_n499_ = ~G25;
  assign new_n501_ = ~G26;
  assign new_n503_ = ~G27;
  assign new_n505_ = ~G28;
  assign new_n507_ = ~G29;
  assign new_n509_ = ~G30;
  assign new_n511_ = ~G31;
  assign new_n513_ = ~G32;
  assign new_n515_ = ~G33;
  assign new_n517_ = ~G34;
  assign new_n519_ = ~G35;
  assign new_n521_ = ~G36;
  assign new_n523_ = ~G37;
  assign new_n525_ = ~G38;
  assign new_n527_ = ~G39;
  assign new_n529_ = ~G40;
  assign new_n531_ = ~G41;
  assign new_n532_ = n286_lo;
  assign new_n533_ = ~n286_lo;
  assign new_n534_ = n298_lo;
  assign new_n535_ = ~n298_lo;
  assign new_n536_ = n310_lo;
  assign new_n537_ = ~n310_lo;
  assign new_n538_ = n322_lo;
  assign new_n539_ = ~n322_lo;
  assign new_n540_ = n334_lo;
  assign new_n541_ = ~n334_lo;
  assign new_n542_ = n346_lo;
  assign new_n543_ = ~n346_lo;
  assign new_n544_ = n358_lo;
  assign new_n545_ = ~n358_lo;
  assign new_n546_ = n370_lo;
  assign new_n547_ = ~n370_lo;
  assign new_n548_ = n382_lo;
  assign new_n549_ = ~n382_lo;
  assign new_n550_ = n394_lo;
  assign new_n551_ = ~n394_lo;
  assign new_n552_ = n406_lo;
  assign new_n553_ = ~n406_lo;
  assign new_n554_ = n418_lo;
  assign new_n555_ = ~n418_lo;
  assign new_n556_ = n430_lo;
  assign new_n557_ = ~n430_lo;
  assign new_n558_ = n442_lo;
  assign new_n559_ = ~n442_lo;
  assign new_n560_ = n454_lo;
  assign new_n561_ = ~n454_lo;
  assign new_n562_ = n466_lo;
  assign new_n563_ = ~n466_lo;
  assign new_n564_ = n478_lo;
  assign new_n565_ = ~n478_lo;
  assign new_n566_ = n490_lo;
  assign new_n567_ = ~n490_lo;
  assign new_n568_ = n502_lo;
  assign new_n569_ = ~n502_lo;
  assign new_n570_ = n514_lo;
  assign new_n571_ = ~n514_lo;
  assign new_n572_ = n526_lo;
  assign new_n573_ = ~n526_lo;
  assign new_n574_ = n538_lo;
  assign new_n575_ = ~n538_lo;
  assign new_n576_ = n550_lo;
  assign new_n577_ = ~n550_lo;
  assign new_n578_ = n562_lo;
  assign new_n579_ = ~n562_lo;
  assign new_n580_ = n574_lo;
  assign new_n581_ = ~n574_lo;
  assign new_n582_ = n586_lo;
  assign new_n583_ = ~n586_lo;
  assign new_n584_ = n598_lo;
  assign new_n585_ = ~n598_lo;
  assign new_n586_ = n610_lo;
  assign new_n587_ = ~n610_lo;
  assign new_n588_ = n622_lo;
  assign new_n589_ = ~n622_lo;
  assign new_n590_ = n634_lo;
  assign new_n591_ = ~n634_lo;
  assign new_n592_ = n646_lo;
  assign new_n593_ = ~n646_lo;
  assign new_n594_ = n658_lo;
  assign new_n595_ = ~n658_lo;
  assign new_n597_ = ~n661_lo;
  assign new_n599_ = ~n673_lo;
  assign new_n601_ = ~n685_lo;
  assign new_n603_ = ~n697_lo;
  assign new_n605_ = ~n709_lo;
  assign new_n607_ = ~n721_lo;
  assign new_n609_ = ~n733_lo;
  assign new_n611_ = ~n745_lo;
  assign new_n613_ = ~n757_lo;
  assign new_n614_ = n1248_o2;
  assign new_n615_ = ~n1248_o2;
  assign new_n616_ = n1249_o2;
  assign new_n617_ = ~n1249_o2;
  assign new_n618_ = n1250_o2;
  assign new_n619_ = ~n1250_o2;
  assign new_n620_ = n1251_o2;
  assign new_n621_ = ~n1251_o2;
  assign new_n622_ = n1252_o2;
  assign new_n623_ = ~n1252_o2;
  assign new_n624_ = n1253_o2;
  assign new_n625_ = ~n1253_o2;
  assign new_n626_ = n1254_o2;
  assign new_n627_ = ~n1254_o2;
  assign new_n628_ = n1255_o2;
  assign new_n629_ = ~n1255_o2;
  assign new_n631_ = ~n1207_o2;
  assign new_n633_ = ~n1208_o2;
  assign new_n635_ = ~n1209_o2;
  assign new_n637_ = ~n1210_o2;
  assign new_n639_ = ~n1211_o2;
  assign new_n641_ = ~n1212_o2;
  assign new_n643_ = ~n1213_o2;
  assign new_n645_ = ~n1214_o2;
  assign new_n647_ = ~n1215_o2;
  assign new_n649_ = ~n1216_o2;
  assign new_n651_ = ~n1217_o2;
  assign new_n653_ = ~n1218_o2;
  assign new_n655_ = ~n1219_o2;
  assign new_n657_ = ~n1220_o2;
  assign new_n659_ = ~n1221_o2;
  assign new_n661_ = ~n1222_o2;
  assign new_n663_ = ~n1223_o2;
  assign new_n665_ = ~n1224_o2;
  assign new_n667_ = ~n1225_o2;
  assign new_n669_ = ~n1226_o2;
  assign new_n671_ = ~n1227_o2;
  assign new_n673_ = ~n1228_o2;
  assign new_n675_ = ~n1229_o2;
  assign new_n677_ = ~n1230_o2;
  assign new_n679_ = ~n1231_o2;
  assign new_n681_ = ~n1232_o2;
  assign new_n683_ = ~n1233_o2;
  assign new_n685_ = ~n1234_o2;
  assign new_n687_ = ~n1235_o2;
  assign new_n689_ = ~n1236_o2;
  assign new_n691_ = ~n1237_o2;
  assign new_n693_ = ~n1238_o2;
  assign new_n694_ = G374_o2;
  assign new_n695_ = ~G374_o2;
  assign new_n696_ = G376_o2;
  assign new_n697_ = ~G376_o2;
  assign new_n698_ = G370_o2;
  assign new_n699_ = ~G370_o2;
  assign new_n700_ = G372_o2;
  assign new_n701_ = ~G372_o2;
  assign new_n702_ = G373_o2;
  assign new_n703_ = ~G373_o2;
  assign new_n704_ = G377_o2;
  assign new_n705_ = ~G377_o2;
  assign new_n706_ = G371_o2;
  assign new_n707_ = ~G371_o2;
  assign new_n708_ = G375_o2;
  assign new_n709_ = ~G375_o2;
  assign new_n710_ = G354_o2;
  assign new_n711_ = ~G354_o2;
  assign new_n712_ = G356_o2;
  assign new_n713_ = ~G356_o2;
  assign new_n714_ = G350_o2;
  assign new_n715_ = ~G350_o2;
  assign new_n716_ = G352_o2;
  assign new_n717_ = ~G352_o2;
  assign new_n718_ = G353_o2;
  assign new_n719_ = ~G353_o2;
  assign new_n720_ = G357_o2;
  assign new_n721_ = ~G357_o2;
  assign new_n722_ = G351_o2;
  assign new_n723_ = ~G351_o2;
  assign new_n724_ = G355_o2;
  assign new_n725_ = ~G355_o2;
  assign new_n726_ = G386_o2;
  assign new_n727_ = ~G386_o2;
  assign new_n728_ = G391_o2;
  assign new_n729_ = ~G391_o2;
  assign new_n730_ = n283_lo_buf_o2;
  assign new_n731_ = ~n283_lo_buf_o2;
  assign new_n732_ = n295_lo_buf_o2;
  assign new_n733_ = ~n295_lo_buf_o2;
  assign new_n734_ = n307_lo_buf_o2;
  assign new_n735_ = ~n307_lo_buf_o2;
  assign new_n736_ = n319_lo_buf_o2;
  assign new_n737_ = ~n319_lo_buf_o2;
  assign new_n738_ = n331_lo_buf_o2;
  assign new_n739_ = ~n331_lo_buf_o2;
  assign new_n740_ = n343_lo_buf_o2;
  assign new_n741_ = ~n343_lo_buf_o2;
  assign new_n742_ = n355_lo_buf_o2;
  assign new_n743_ = ~n355_lo_buf_o2;
  assign new_n744_ = n367_lo_buf_o2;
  assign new_n745_ = ~n367_lo_buf_o2;
  assign new_n746_ = n379_lo_buf_o2;
  assign new_n747_ = ~n379_lo_buf_o2;
  assign new_n748_ = n391_lo_buf_o2;
  assign new_n749_ = ~n391_lo_buf_o2;
  assign new_n750_ = n403_lo_buf_o2;
  assign new_n751_ = ~n403_lo_buf_o2;
  assign new_n752_ = n415_lo_buf_o2;
  assign new_n753_ = ~n415_lo_buf_o2;
  assign new_n754_ = n427_lo_buf_o2;
  assign new_n755_ = ~n427_lo_buf_o2;
  assign new_n756_ = n439_lo_buf_o2;
  assign new_n757_ = ~n439_lo_buf_o2;
  assign new_n758_ = n451_lo_buf_o2;
  assign new_n759_ = ~n451_lo_buf_o2;
  assign new_n760_ = n463_lo_buf_o2;
  assign new_n761_ = ~n463_lo_buf_o2;
  assign new_n762_ = n475_lo_buf_o2;
  assign new_n763_ = ~n475_lo_buf_o2;
  assign new_n764_ = n487_lo_buf_o2;
  assign new_n765_ = ~n487_lo_buf_o2;
  assign new_n766_ = n499_lo_buf_o2;
  assign new_n767_ = ~n499_lo_buf_o2;
  assign new_n768_ = n511_lo_buf_o2;
  assign new_n769_ = ~n511_lo_buf_o2;
  assign new_n770_ = n523_lo_buf_o2;
  assign new_n771_ = ~n523_lo_buf_o2;
  assign new_n772_ = n535_lo_buf_o2;
  assign new_n773_ = ~n535_lo_buf_o2;
  assign new_n774_ = n547_lo_buf_o2;
  assign new_n775_ = ~n547_lo_buf_o2;
  assign new_n776_ = n559_lo_buf_o2;
  assign new_n777_ = ~n559_lo_buf_o2;
  assign new_n778_ = n571_lo_buf_o2;
  assign new_n779_ = ~n571_lo_buf_o2;
  assign new_n780_ = n583_lo_buf_o2;
  assign new_n781_ = ~n583_lo_buf_o2;
  assign new_n782_ = n595_lo_buf_o2;
  assign new_n783_ = ~n595_lo_buf_o2;
  assign new_n784_ = n607_lo_buf_o2;
  assign new_n785_ = ~n607_lo_buf_o2;
  assign new_n786_ = n619_lo_buf_o2;
  assign new_n787_ = ~n619_lo_buf_o2;
  assign new_n788_ = n631_lo_buf_o2;
  assign new_n789_ = ~n631_lo_buf_o2;
  assign new_n790_ = n643_lo_buf_o2;
  assign new_n791_ = ~n643_lo_buf_o2;
  assign new_n792_ = n655_lo_buf_o2;
  assign new_n793_ = ~n655_lo_buf_o2;
  assign new_n794_ = G234_o2;
  assign new_n795_ = ~G234_o2;
  assign new_n796_ = G247_o2;
  assign new_n797_ = ~G247_o2;
  assign new_n798_ = G260_o2;
  assign new_n799_ = ~G260_o2;
  assign new_n800_ = G273_o2;
  assign new_n801_ = ~G273_o2;
  assign new_n802_ = G286_o2;
  assign new_n803_ = ~G286_o2;
  assign new_n804_ = G299_o2;
  assign new_n805_ = ~G299_o2;
  assign new_n806_ = G312_o2;
  assign new_n807_ = ~G312_o2;
  assign new_n808_ = G325_o2;
  assign new_n809_ = ~G325_o2;
  assign new_n810_ = n667_lo_buf_o2;
  assign new_n811_ = ~n667_lo_buf_o2;
  assign new_n812_ = n679_lo_buf_o2;
  assign new_n813_ = ~n679_lo_buf_o2;
  assign new_n814_ = n691_lo_buf_o2;
  assign new_n815_ = ~n691_lo_buf_o2;
  assign new_n816_ = n703_lo_buf_o2;
  assign new_n817_ = ~n703_lo_buf_o2;
  assign new_n818_ = n715_lo_buf_o2;
  assign new_n819_ = ~n715_lo_buf_o2;
  assign new_n820_ = n727_lo_buf_o2;
  assign new_n821_ = ~n727_lo_buf_o2;
  assign new_n822_ = n739_lo_buf_o2;
  assign new_n823_ = ~n739_lo_buf_o2;
  assign new_n824_ = n751_lo_buf_o2;
  assign new_n825_ = ~n751_lo_buf_o2;
  assign new_n826_ = n763_lo_buf_o2;
  assign new_n827_ = ~n763_lo_buf_o2;
  assign new_n828_ = G186_o2;
  assign new_n829_ = ~G186_o2;
  assign new_n830_ = G189_o2;
  assign new_n831_ = ~G189_o2;
  assign new_n832_ = G192_o2;
  assign new_n833_ = ~G192_o2;
  assign new_n834_ = G195_o2;
  assign new_n835_ = ~G195_o2;
  assign new_n836_ = G198_o2;
  assign new_n837_ = ~G198_o2;
  assign new_n838_ = G201_o2;
  assign new_n839_ = ~G201_o2;
  assign new_n840_ = G204_o2;
  assign new_n841_ = ~G204_o2;
  assign new_n842_ = G207_o2;
  assign new_n843_ = ~G207_o2;
  assign new_n844_ = n280_lo_buf_o2;
  assign new_n845_ = ~n280_lo_buf_o2;
  assign new_n846_ = n292_lo_buf_o2;
  assign new_n847_ = ~n292_lo_buf_o2;
  assign new_n848_ = n304_lo_buf_o2;
  assign new_n849_ = ~n304_lo_buf_o2;
  assign new_n850_ = n316_lo_buf_o2;
  assign new_n851_ = ~n316_lo_buf_o2;
  assign new_n852_ = n328_lo_buf_o2;
  assign new_n853_ = ~n328_lo_buf_o2;
  assign new_n854_ = n340_lo_buf_o2;
  assign new_n855_ = ~n340_lo_buf_o2;
  assign new_n856_ = n352_lo_buf_o2;
  assign new_n857_ = ~n352_lo_buf_o2;
  assign new_n858_ = n364_lo_buf_o2;
  assign new_n859_ = ~n364_lo_buf_o2;
  assign new_n860_ = n376_lo_buf_o2;
  assign new_n861_ = ~n376_lo_buf_o2;
  assign new_n862_ = n388_lo_buf_o2;
  assign new_n863_ = ~n388_lo_buf_o2;
  assign new_n864_ = n400_lo_buf_o2;
  assign new_n865_ = ~n400_lo_buf_o2;
  assign new_n866_ = n412_lo_buf_o2;
  assign new_n867_ = ~n412_lo_buf_o2;
  assign new_n868_ = n424_lo_buf_o2;
  assign new_n869_ = ~n424_lo_buf_o2;
  assign new_n870_ = n436_lo_buf_o2;
  assign new_n871_ = ~n436_lo_buf_o2;
  assign new_n872_ = n448_lo_buf_o2;
  assign new_n873_ = ~n448_lo_buf_o2;
  assign new_n874_ = n460_lo_buf_o2;
  assign new_n875_ = ~n460_lo_buf_o2;
  assign new_n876_ = n472_lo_buf_o2;
  assign new_n877_ = ~n472_lo_buf_o2;
  assign new_n878_ = n484_lo_buf_o2;
  assign new_n879_ = ~n484_lo_buf_o2;
  assign new_n880_ = n496_lo_buf_o2;
  assign new_n881_ = ~n496_lo_buf_o2;
  assign new_n882_ = n508_lo_buf_o2;
  assign new_n883_ = ~n508_lo_buf_o2;
  assign new_n884_ = n520_lo_buf_o2;
  assign new_n885_ = ~n520_lo_buf_o2;
  assign new_n886_ = n532_lo_buf_o2;
  assign new_n887_ = ~n532_lo_buf_o2;
  assign new_n888_ = n544_lo_buf_o2;
  assign new_n889_ = ~n544_lo_buf_o2;
  assign new_n890_ = n556_lo_buf_o2;
  assign new_n891_ = ~n556_lo_buf_o2;
  assign new_n892_ = n568_lo_buf_o2;
  assign new_n893_ = ~n568_lo_buf_o2;
  assign new_n894_ = n580_lo_buf_o2;
  assign new_n895_ = ~n580_lo_buf_o2;
  assign new_n896_ = n592_lo_buf_o2;
  assign new_n897_ = ~n592_lo_buf_o2;
  assign new_n898_ = n604_lo_buf_o2;
  assign new_n899_ = ~n604_lo_buf_o2;
  assign new_n900_ = n616_lo_buf_o2;
  assign new_n901_ = ~n616_lo_buf_o2;
  assign new_n902_ = n628_lo_buf_o2;
  assign new_n903_ = ~n628_lo_buf_o2;
  assign new_n904_ = n640_lo_buf_o2;
  assign new_n905_ = ~n640_lo_buf_o2;
  assign new_n906_ = n652_lo_buf_o2;
  assign new_n907_ = ~n652_lo_buf_o2;
  assign new_n908_ = new_n715_ & new_n1782_;
  assign new_n909_ = new_n714_ | new_n1787_;
  assign new_n910_ = new_n908_ & new_n1792_;
  assign new_n911_ = new_n909_ | new_n1797_;
  assign new_n912_ = new_n910_ & new_n723_;
  assign new_n913_ = new_n911_ | new_n722_;
  assign new_n914_ = new_n912_ & new_n1801_;
  assign new_n915_ = new_n913_ | new_n1804_;
  assign new_n916_ = new_n1807_ & new_n1811_;
  assign new_n917_ = new_n1815_ | new_n1819_;
  assign new_n918_ = new_n917_ | new_n532_;
  assign new_n919_ = new_n916_ | new_n533_;
  assign new_n920_ = new_n919_ & new_n918_;
  assign new_n921_ = new_n1807_ & new_n1824_;
  assign new_n922_ = new_n1815_ | new_n1829_;
  assign new_n923_ = new_n922_ | new_n534_;
  assign new_n924_ = new_n921_ | new_n535_;
  assign new_n925_ = new_n924_ & new_n923_;
  assign new_n926_ = new_n1808_ & new_n1834_;
  assign new_n927_ = new_n1816_ | new_n1839_;
  assign new_n928_ = new_n927_ | new_n536_;
  assign new_n929_ = new_n926_ | new_n537_;
  assign new_n930_ = new_n929_ & new_n928_;
  assign new_n931_ = new_n1808_ & new_n1844_;
  assign new_n932_ = new_n1816_ | new_n1849_;
  assign new_n933_ = new_n932_ | new_n538_;
  assign new_n934_ = new_n931_ | new_n539_;
  assign new_n935_ = new_n934_ & new_n933_;
  assign new_n936_ = new_n717_ & new_n1782_;
  assign new_n937_ = new_n716_ | new_n1787_;
  assign new_n938_ = new_n936_ & new_n719_;
  assign new_n939_ = new_n937_ | new_n718_;
  assign new_n940_ = new_n938_ & new_n1854_;
  assign new_n941_ = new_n939_ | new_n1859_;
  assign new_n942_ = new_n940_ & new_n1801_;
  assign new_n943_ = new_n941_ | new_n1804_;
  assign new_n944_ = new_n1863_ & new_n1811_;
  assign new_n945_ = new_n1866_ | new_n1819_;
  assign new_n946_ = new_n945_ | new_n540_;
  assign new_n947_ = new_n944_ | new_n541_;
  assign new_n948_ = new_n947_ & new_n946_;
  assign new_n949_ = new_n1863_ & new_n1824_;
  assign new_n950_ = new_n1866_ | new_n1829_;
  assign new_n951_ = new_n950_ | new_n542_;
  assign new_n952_ = new_n949_ | new_n543_;
  assign new_n953_ = new_n952_ & new_n951_;
  assign new_n954_ = new_n1864_ & new_n1834_;
  assign new_n955_ = new_n1867_ | new_n1839_;
  assign new_n956_ = new_n955_ | new_n544_;
  assign new_n957_ = new_n954_ | new_n545_;
  assign new_n958_ = new_n957_ & new_n956_;
  assign new_n959_ = new_n1864_ & new_n1844_;
  assign new_n960_ = new_n1867_ | new_n1849_;
  assign new_n961_ = new_n960_ | new_n546_;
  assign new_n962_ = new_n959_ | new_n547_;
  assign new_n963_ = new_n962_ & new_n961_;
  assign new_n964_ = new_n711_ & new_n1870_;
  assign new_n965_ = new_n710_ | new_n1875_;
  assign new_n966_ = new_n964_ & new_n1792_;
  assign new_n967_ = new_n965_ | new_n1797_;
  assign new_n968_ = new_n966_ & new_n725_;
  assign new_n969_ = new_n967_ | new_n724_;
  assign new_n970_ = new_n968_ & new_n1802_;
  assign new_n971_ = new_n969_ | new_n1805_;
  assign new_n972_ = new_n1879_ & new_n1812_;
  assign new_n973_ = new_n1882_ | new_n1820_;
  assign new_n974_ = new_n973_ | new_n548_;
  assign new_n975_ = new_n972_ | new_n549_;
  assign new_n976_ = new_n975_ & new_n974_;
  assign new_n977_ = new_n1879_ & new_n1825_;
  assign new_n978_ = new_n1882_ | new_n1830_;
  assign new_n979_ = new_n978_ | new_n550_;
  assign new_n980_ = new_n977_ | new_n551_;
  assign new_n981_ = new_n980_ & new_n979_;
  assign new_n982_ = new_n1880_ & new_n1835_;
  assign new_n983_ = new_n1883_ | new_n1840_;
  assign new_n984_ = new_n983_ | new_n552_;
  assign new_n985_ = new_n982_ | new_n553_;
  assign new_n986_ = new_n985_ & new_n984_;
  assign new_n987_ = new_n1880_ & new_n1845_;
  assign new_n988_ = new_n1883_ | new_n1850_;
  assign new_n989_ = new_n988_ | new_n554_;
  assign new_n990_ = new_n987_ | new_n555_;
  assign new_n991_ = new_n990_ & new_n989_;
  assign new_n992_ = new_n713_ & new_n1870_;
  assign new_n993_ = new_n712_ | new_n1875_;
  assign new_n994_ = new_n992_ & new_n721_;
  assign new_n995_ = new_n993_ | new_n720_;
  assign new_n996_ = new_n994_ & new_n1854_;
  assign new_n997_ = new_n995_ | new_n1859_;
  assign new_n998_ = new_n996_ & new_n1802_;
  assign new_n999_ = new_n997_ | new_n1805_;
  assign new_n1000_ = new_n1885_ & new_n1812_;
  assign new_n1001_ = new_n1888_ | new_n1820_;
  assign new_n1002_ = new_n1001_ | new_n556_;
  assign new_n1003_ = new_n1000_ | new_n557_;
  assign new_n1004_ = new_n1003_ & new_n1002_;
  assign new_n1005_ = new_n1885_ & new_n1825_;
  assign new_n1006_ = new_n1888_ | new_n1830_;
  assign new_n1007_ = new_n1006_ | new_n558_;
  assign new_n1008_ = new_n1005_ | new_n559_;
  assign new_n1009_ = new_n1008_ & new_n1007_;
  assign new_n1010_ = new_n1886_ & new_n1835_;
  assign new_n1011_ = new_n1889_ | new_n1840_;
  assign new_n1012_ = new_n1011_ | new_n560_;
  assign new_n1013_ = new_n1010_ | new_n561_;
  assign new_n1014_ = new_n1013_ & new_n1012_;
  assign new_n1015_ = new_n1886_ & new_n1845_;
  assign new_n1016_ = new_n1889_ | new_n1850_;
  assign new_n1017_ = new_n1016_ | new_n562_;
  assign new_n1018_ = new_n1015_ | new_n563_;
  assign new_n1019_ = new_n1018_ & new_n1017_;
  assign new_n1020_ = new_n699_ & new_n1813_;
  assign new_n1021_ = new_n698_ | new_n1821_;
  assign new_n1022_ = new_n1020_ & new_n1836_;
  assign new_n1023_ = new_n1021_ | new_n1841_;
  assign new_n1024_ = new_n1022_ & new_n707_;
  assign new_n1025_ = new_n1023_ | new_n706_;
  assign new_n1026_ = new_n1024_ & new_n1891_;
  assign new_n1027_ = new_n1025_ | new_n1894_;
  assign new_n1028_ = new_n1897_ & new_n1783_;
  assign new_n1029_ = new_n1900_ | new_n1788_;
  assign new_n1030_ = new_n1029_ | new_n564_;
  assign new_n1031_ = new_n1028_ | new_n565_;
  assign new_n1032_ = new_n1031_ & new_n1030_;
  assign new_n1033_ = new_n1897_ & new_n1871_;
  assign new_n1034_ = new_n1900_ | new_n1876_;
  assign new_n1035_ = new_n1034_ | new_n566_;
  assign new_n1036_ = new_n1033_ | new_n567_;
  assign new_n1037_ = new_n1036_ & new_n1035_;
  assign new_n1038_ = new_n1898_ & new_n1793_;
  assign new_n1039_ = new_n1901_ | new_n1798_;
  assign new_n1040_ = new_n1039_ | new_n568_;
  assign new_n1041_ = new_n1038_ | new_n569_;
  assign new_n1042_ = new_n1041_ & new_n1040_;
  assign new_n1043_ = new_n1898_ & new_n1855_;
  assign new_n1044_ = new_n1901_ | new_n1860_;
  assign new_n1045_ = new_n1044_ | new_n570_;
  assign new_n1046_ = new_n1043_ | new_n571_;
  assign new_n1047_ = new_n1046_ & new_n1045_;
  assign new_n1048_ = new_n701_ & new_n1813_;
  assign new_n1049_ = new_n700_ | new_n1821_;
  assign new_n1050_ = new_n1048_ & new_n703_;
  assign new_n1051_ = new_n1049_ | new_n702_;
  assign new_n1052_ = new_n1050_ & new_n1846_;
  assign new_n1053_ = new_n1051_ | new_n1851_;
  assign new_n1054_ = new_n1052_ & new_n1891_;
  assign new_n1055_ = new_n1053_ | new_n1894_;
  assign new_n1056_ = new_n1903_ & new_n1783_;
  assign new_n1057_ = new_n1906_ | new_n1788_;
  assign new_n1058_ = new_n1057_ | new_n572_;
  assign new_n1059_ = new_n1056_ | new_n573_;
  assign new_n1060_ = new_n1059_ & new_n1058_;
  assign new_n1061_ = new_n1903_ & new_n1871_;
  assign new_n1062_ = new_n1906_ | new_n1876_;
  assign new_n1063_ = new_n1062_ | new_n574_;
  assign new_n1064_ = new_n1061_ | new_n575_;
  assign new_n1065_ = new_n1064_ & new_n1063_;
  assign new_n1066_ = new_n1904_ & new_n1793_;
  assign new_n1067_ = new_n1907_ | new_n1798_;
  assign new_n1068_ = new_n1067_ | new_n576_;
  assign new_n1069_ = new_n1066_ | new_n577_;
  assign new_n1070_ = new_n1069_ & new_n1068_;
  assign new_n1071_ = new_n1904_ & new_n1855_;
  assign new_n1072_ = new_n1907_ | new_n1860_;
  assign new_n1073_ = new_n1072_ | new_n578_;
  assign new_n1074_ = new_n1071_ | new_n579_;
  assign new_n1075_ = new_n1074_ & new_n1073_;
  assign new_n1076_ = new_n695_ & new_n1826_;
  assign new_n1077_ = new_n694_ | new_n1831_;
  assign new_n1078_ = new_n1076_ & new_n1836_;
  assign new_n1079_ = new_n1077_ | new_n1841_;
  assign new_n1080_ = new_n1078_ & new_n709_;
  assign new_n1081_ = new_n1079_ | new_n708_;
  assign new_n1082_ = new_n1080_ & new_n1892_;
  assign new_n1083_ = new_n1081_ | new_n1895_;
  assign new_n1084_ = new_n1909_ & new_n1784_;
  assign new_n1085_ = new_n1912_ | new_n1789_;
  assign new_n1086_ = new_n1085_ | new_n580_;
  assign new_n1087_ = new_n1084_ | new_n581_;
  assign new_n1088_ = new_n1087_ & new_n1086_;
  assign new_n1089_ = new_n1909_ & new_n1872_;
  assign new_n1090_ = new_n1912_ | new_n1877_;
  assign new_n1091_ = new_n1090_ | new_n582_;
  assign new_n1092_ = new_n1089_ | new_n583_;
  assign new_n1093_ = new_n1092_ & new_n1091_;
  assign new_n1094_ = new_n1910_ & new_n1794_;
  assign new_n1095_ = new_n1913_ | new_n1799_;
  assign new_n1096_ = new_n1095_ | new_n584_;
  assign new_n1097_ = new_n1094_ | new_n585_;
  assign new_n1098_ = new_n1097_ & new_n1096_;
  assign new_n1099_ = new_n1910_ & new_n1856_;
  assign new_n1100_ = new_n1913_ | new_n1861_;
  assign new_n1101_ = new_n1100_ | new_n586_;
  assign new_n1102_ = new_n1099_ | new_n587_;
  assign new_n1103_ = new_n1102_ & new_n1101_;
  assign new_n1104_ = new_n697_ & new_n1826_;
  assign new_n1105_ = new_n696_ | new_n1831_;
  assign new_n1106_ = new_n1104_ & new_n705_;
  assign new_n1107_ = new_n1105_ | new_n704_;
  assign new_n1108_ = new_n1106_ & new_n1846_;
  assign new_n1109_ = new_n1107_ | new_n1851_;
  assign new_n1110_ = new_n1108_ & new_n1892_;
  assign new_n1111_ = new_n1109_ | new_n1895_;
  assign new_n1112_ = new_n1915_ & new_n1784_;
  assign new_n1113_ = new_n1918_ | new_n1789_;
  assign new_n1114_ = new_n1113_ | new_n588_;
  assign new_n1115_ = new_n1112_ | new_n589_;
  assign new_n1116_ = new_n1115_ & new_n1114_;
  assign new_n1117_ = new_n1915_ & new_n1872_;
  assign new_n1118_ = new_n1918_ | new_n1877_;
  assign new_n1119_ = new_n1118_ | new_n590_;
  assign new_n1120_ = new_n1117_ | new_n591_;
  assign new_n1121_ = new_n1120_ & new_n1119_;
  assign new_n1122_ = new_n1916_ & new_n1794_;
  assign new_n1123_ = new_n1919_ | new_n1799_;
  assign new_n1124_ = new_n1123_ | new_n592_;
  assign new_n1125_ = new_n1122_ | new_n593_;
  assign new_n1126_ = new_n1125_ & new_n1124_;
  assign new_n1127_ = new_n1916_ & new_n1856_;
  assign new_n1128_ = new_n1919_ | new_n1861_;
  assign new_n1129_ = new_n1128_ | new_n594_;
  assign new_n1130_ = new_n1127_ | new_n595_;
  assign new_n1131_ = new_n1130_ & new_n1129_;
  assign new_n1132_ = new_n1920_ | new_n1921_;
  assign new_n1133_ = new_n1922_ | new_n1924_;
  assign new_n1134_ = new_n1133_ | new_n1926_;
  assign new_n1135_ = new_n1922_ | new_n1929_;
  assign new_n1136_ = new_n1135_ | new_n1932_;
  assign new_n1137_ = new_n1934_ | new_n1921_;
  assign new_n1138_ = new_n1137_ | new_n1924_;
  assign new_n1139_ = new_n1138_ | new_n1932_;
  assign new_n1140_ = new_n1920_ | new_n1937_;
  assign new_n1141_ = new_n1140_ | new_n1923_;
  assign new_n1142_ = new_n1141_ | new_n1931_;
  assign new_n1143_ = new_n1136_ & new_n1134_;
  assign new_n1144_ = new_n1143_ & new_n1139_;
  assign new_n1145_ = new_n1144_ & new_n1142_;
  assign new_n1146_ = new_n1939_ | new_n1940_;
  assign new_n1147_ = new_n1941_ | new_n1943_;
  assign new_n1148_ = new_n1147_ | new_n1945_;
  assign new_n1149_ = new_n1941_ | new_n1948_;
  assign new_n1150_ = new_n1149_ | new_n1951_;
  assign new_n1151_ = new_n1953_ | new_n1940_;
  assign new_n1152_ = new_n1151_ | new_n1943_;
  assign new_n1153_ = new_n1152_ | new_n1951_;
  assign new_n1154_ = new_n1939_ | new_n1956_;
  assign new_n1155_ = new_n1154_ | new_n1942_;
  assign new_n1156_ = new_n1155_ | new_n1950_;
  assign new_n1157_ = new_n1150_ & new_n1148_;
  assign new_n1158_ = new_n1157_ & new_n1153_;
  assign new_n1159_ = new_n1158_ & new_n1156_;
  assign new_n1160_ = new_n1958_ & new_n1960_;
  assign new_n1161_ = new_n1962_ | new_n1963_;
  assign new_n1162_ = new_n1962_ & new_n1963_;
  assign new_n1163_ = new_n1958_ | new_n1960_;
  assign new_n1164_ = new_n1163_ & new_n1161_;
  assign new_n1165_ = new_n1162_ | new_n1160_;
  assign new_n1166_ = new_n1964_ & new_n1966_;
  assign new_n1167_ = new_n1968_ | new_n1969_;
  assign new_n1168_ = new_n1968_ & new_n1969_;
  assign new_n1169_ = new_n1964_ | new_n1966_;
  assign new_n1170_ = new_n1169_ & new_n1167_;
  assign new_n1171_ = new_n1168_ | new_n1166_;
  assign new_n1172_ = new_n1970_ & new_n1971_;
  assign new_n1173_ = new_n1972_ | new_n1973_;
  assign new_n1174_ = new_n1972_ & new_n1973_;
  assign new_n1175_ = new_n1970_ | new_n1971_;
  assign new_n1176_ = new_n1175_ & new_n1173_;
  assign new_n1177_ = new_n1174_ | new_n1172_;
  assign new_n1178_ = new_n1976_ & new_n810_;
  assign new_n1179_ = new_n1983_ | new_n811_;
  assign new_n1180_ = new_n1989_ & new_n1992_;
  assign new_n1181_ = new_n1995_ | new_n1998_;
  assign new_n1182_ = new_n1995_ & new_n1998_;
  assign new_n1183_ = new_n1989_ | new_n1992_;
  assign new_n1184_ = new_n1183_ & new_n1181_;
  assign new_n1185_ = new_n1182_ | new_n1180_;
  assign new_n1186_ = new_n2000_ & new_n2001_;
  assign new_n1187_ = new_n2002_ | new_n2003_;
  assign new_n1188_ = new_n2002_ & new_n2003_;
  assign new_n1189_ = new_n2000_ | new_n2001_;
  assign new_n1190_ = new_n1189_ & new_n1187_;
  assign new_n1191_ = new_n1188_ | new_n1186_;
  assign new_n1192_ = new_n1190_ | new_n1177_;
  assign new_n1193_ = new_n1191_ | new_n1176_;
  assign new_n1194_ = new_n1193_ & new_n1192_;
  assign new_n1195_ = new_n2004_ & new_n2006_;
  assign new_n1196_ = new_n2008_ | new_n2009_;
  assign new_n1197_ = new_n2008_ & new_n2009_;
  assign new_n1198_ = new_n2004_ | new_n2006_;
  assign new_n1199_ = new_n1198_ & new_n1196_;
  assign new_n1200_ = new_n1197_ | new_n1195_;
  assign new_n1201_ = new_n2010_ & new_n2012_;
  assign new_n1202_ = new_n2014_ | new_n2015_;
  assign new_n1203_ = new_n2014_ & new_n2015_;
  assign new_n1204_ = new_n2010_ | new_n2012_;
  assign new_n1205_ = new_n1204_ & new_n1202_;
  assign new_n1206_ = new_n1203_ | new_n1201_;
  assign new_n1207_ = new_n2016_ & new_n2017_;
  assign new_n1208_ = new_n2018_ | new_n2019_;
  assign new_n1209_ = new_n2018_ & new_n2019_;
  assign new_n1210_ = new_n2016_ | new_n2017_;
  assign new_n1211_ = new_n1210_ & new_n1208_;
  assign new_n1212_ = new_n1209_ | new_n1207_;
  assign new_n1213_ = new_n1976_ & new_n812_;
  assign new_n1214_ = new_n1983_ | new_n813_;
  assign new_n1215_ = new_n2021_ & new_n2024_;
  assign new_n1216_ = new_n2027_ | new_n2030_;
  assign new_n1217_ = new_n2027_ & new_n2030_;
  assign new_n1218_ = new_n2021_ | new_n2024_;
  assign new_n1219_ = new_n1218_ & new_n1216_;
  assign new_n1220_ = new_n1217_ | new_n1215_;
  assign new_n1221_ = new_n2032_ & new_n2033_;
  assign new_n1222_ = new_n2034_ | new_n2035_;
  assign new_n1223_ = new_n2034_ & new_n2035_;
  assign new_n1224_ = new_n2032_ | new_n2033_;
  assign new_n1225_ = new_n1224_ & new_n1222_;
  assign new_n1226_ = new_n1223_ | new_n1221_;
  assign new_n1227_ = new_n1225_ | new_n1212_;
  assign new_n1228_ = new_n1226_ | new_n1211_;
  assign new_n1229_ = new_n1228_ & new_n1227_;
  assign new_n1230_ = new_n2036_ & new_n2038_;
  assign new_n1231_ = new_n2040_ | new_n2041_;
  assign new_n1232_ = new_n2040_ & new_n2041_;
  assign new_n1233_ = new_n2036_ | new_n2038_;
  assign new_n1234_ = new_n1233_ & new_n1231_;
  assign new_n1235_ = new_n1232_ | new_n1230_;
  assign new_n1236_ = new_n2042_ & new_n2044_;
  assign new_n1237_ = new_n2046_ | new_n2047_;
  assign new_n1238_ = new_n2046_ & new_n2047_;
  assign new_n1239_ = new_n2042_ | new_n2044_;
  assign new_n1240_ = new_n1239_ & new_n1237_;
  assign new_n1241_ = new_n1238_ | new_n1236_;
  assign new_n1242_ = new_n2048_ & new_n2049_;
  assign new_n1243_ = new_n2050_ | new_n2051_;
  assign new_n1244_ = new_n2050_ & new_n2051_;
  assign new_n1245_ = new_n2048_ | new_n2049_;
  assign new_n1246_ = new_n1245_ & new_n1243_;
  assign new_n1247_ = new_n1244_ | new_n1242_;
  assign new_n1248_ = new_n1977_ & new_n814_;
  assign new_n1249_ = new_n1984_ | new_n815_;
  assign new_n1250_ = new_n2031_ & new_n1993_;
  assign new_n1251_ = new_n2025_ | new_n1999_;
  assign new_n1252_ = new_n2025_ & new_n1999_;
  assign new_n1253_ = new_n2031_ | new_n1993_;
  assign new_n1254_ = new_n1253_ & new_n1251_;
  assign new_n1255_ = new_n1252_ | new_n1250_;
  assign new_n1256_ = new_n2052_ & new_n2053_;
  assign new_n1257_ = new_n2054_ | new_n2055_;
  assign new_n1258_ = new_n2054_ & new_n2055_;
  assign new_n1259_ = new_n2052_ | new_n2053_;
  assign new_n1260_ = new_n1259_ & new_n1257_;
  assign new_n1261_ = new_n1258_ | new_n1256_;
  assign new_n1262_ = new_n1260_ | new_n1247_;
  assign new_n1263_ = new_n1261_ | new_n1246_;
  assign new_n1264_ = new_n1263_ & new_n1262_;
  assign new_n1265_ = new_n2056_ & new_n2058_;
  assign new_n1266_ = new_n2060_ | new_n2061_;
  assign new_n1267_ = new_n2060_ & new_n2061_;
  assign new_n1268_ = new_n2056_ | new_n2058_;
  assign new_n1269_ = new_n1268_ & new_n1266_;
  assign new_n1270_ = new_n1267_ | new_n1265_;
  assign new_n1271_ = new_n2062_ & new_n2064_;
  assign new_n1272_ = new_n2066_ | new_n2067_;
  assign new_n1273_ = new_n2066_ & new_n2067_;
  assign new_n1274_ = new_n2062_ | new_n2064_;
  assign new_n1275_ = new_n1274_ & new_n1272_;
  assign new_n1276_ = new_n1273_ | new_n1271_;
  assign new_n1277_ = new_n2068_ & new_n2069_;
  assign new_n1278_ = new_n2070_ | new_n2071_;
  assign new_n1279_ = new_n2070_ & new_n2071_;
  assign new_n1280_ = new_n2068_ | new_n2069_;
  assign new_n1281_ = new_n1280_ & new_n1278_;
  assign new_n1282_ = new_n1279_ | new_n1277_;
  assign new_n1283_ = new_n1977_ & new_n816_;
  assign new_n1284_ = new_n1984_ | new_n817_;
  assign new_n1285_ = new_n2022_ & new_n1996_;
  assign new_n1286_ = new_n2028_ | new_n1990_;
  assign new_n1287_ = new_n2028_ & new_n1990_;
  assign new_n1288_ = new_n2022_ | new_n1996_;
  assign new_n1289_ = new_n1288_ & new_n1286_;
  assign new_n1290_ = new_n1287_ | new_n1285_;
  assign new_n1291_ = new_n2072_ & new_n2073_;
  assign new_n1292_ = new_n2074_ | new_n2075_;
  assign new_n1293_ = new_n2074_ & new_n2075_;
  assign new_n1294_ = new_n2072_ | new_n2073_;
  assign new_n1295_ = new_n1294_ & new_n1292_;
  assign new_n1296_ = new_n1293_ | new_n1291_;
  assign new_n1297_ = new_n1295_ | new_n1282_;
  assign new_n1298_ = new_n1296_ | new_n1281_;
  assign new_n1299_ = new_n1298_ & new_n1297_;
  assign new_n1300_ = new_n2076_ & new_n2078_;
  assign new_n1301_ = new_n2080_ | new_n2081_;
  assign new_n1302_ = new_n2080_ & new_n2081_;
  assign new_n1303_ = new_n2076_ | new_n2078_;
  assign new_n1304_ = new_n1303_ & new_n1301_;
  assign new_n1305_ = new_n1302_ | new_n1300_;
  assign new_n1306_ = new_n2082_ & new_n2084_;
  assign new_n1307_ = new_n2086_ | new_n2087_;
  assign new_n1308_ = new_n2086_ & new_n2087_;
  assign new_n1309_ = new_n2082_ | new_n2084_;
  assign new_n1310_ = new_n1309_ & new_n1307_;
  assign new_n1311_ = new_n1308_ | new_n1306_;
  assign new_n1312_ = new_n2088_ & new_n2089_;
  assign new_n1313_ = new_n2090_ | new_n2091_;
  assign new_n1314_ = new_n2090_ & new_n2091_;
  assign new_n1315_ = new_n2088_ | new_n2089_;
  assign new_n1316_ = new_n1315_ & new_n1313_;
  assign new_n1317_ = new_n1314_ | new_n1312_;
  assign new_n1318_ = new_n1979_ & new_n818_;
  assign new_n1319_ = new_n1986_ | new_n819_;
  assign new_n1320_ = new_n2093_ & new_n2096_;
  assign new_n1321_ = new_n2099_ | new_n2102_;
  assign new_n1322_ = new_n2099_ & new_n2102_;
  assign new_n1323_ = new_n2093_ | new_n2096_;
  assign new_n1324_ = new_n1323_ & new_n1321_;
  assign new_n1325_ = new_n1322_ | new_n1320_;
  assign new_n1326_ = new_n2104_ & new_n2105_;
  assign new_n1327_ = new_n2106_ | new_n2107_;
  assign new_n1328_ = new_n2106_ & new_n2107_;
  assign new_n1329_ = new_n2104_ | new_n2105_;
  assign new_n1330_ = new_n1329_ & new_n1327_;
  assign new_n1331_ = new_n1328_ | new_n1326_;
  assign new_n1332_ = new_n1330_ | new_n1317_;
  assign new_n1333_ = new_n1331_ | new_n1316_;
  assign new_n1334_ = new_n1333_ & new_n1332_;
  assign new_n1335_ = new_n2108_ & new_n2110_;
  assign new_n1336_ = new_n2112_ | new_n2113_;
  assign new_n1337_ = new_n2112_ & new_n2113_;
  assign new_n1338_ = new_n2108_ | new_n2110_;
  assign new_n1339_ = new_n1338_ & new_n1336_;
  assign new_n1340_ = new_n1337_ | new_n1335_;
  assign new_n1341_ = new_n2114_ & new_n2116_;
  assign new_n1342_ = new_n2118_ | new_n2119_;
  assign new_n1343_ = new_n2118_ & new_n2119_;
  assign new_n1344_ = new_n2114_ | new_n2116_;
  assign new_n1345_ = new_n1344_ & new_n1342_;
  assign new_n1346_ = new_n1343_ | new_n1341_;
  assign new_n1347_ = new_n2120_ & new_n2121_;
  assign new_n1348_ = new_n2122_ | new_n2123_;
  assign new_n1349_ = new_n2122_ & new_n2123_;
  assign new_n1350_ = new_n2120_ | new_n2121_;
  assign new_n1351_ = new_n1350_ & new_n1348_;
  assign new_n1352_ = new_n1349_ | new_n1347_;
  assign new_n1353_ = new_n1979_ & new_n820_;
  assign new_n1354_ = new_n1986_ | new_n821_;
  assign new_n1355_ = new_n2125_ & new_n2128_;
  assign new_n1356_ = new_n2131_ | new_n2134_;
  assign new_n1357_ = new_n2131_ & new_n2134_;
  assign new_n1358_ = new_n2125_ | new_n2128_;
  assign new_n1359_ = new_n1358_ & new_n1356_;
  assign new_n1360_ = new_n1357_ | new_n1355_;
  assign new_n1361_ = new_n2136_ & new_n2137_;
  assign new_n1362_ = new_n2138_ | new_n2139_;
  assign new_n1363_ = new_n2138_ & new_n2139_;
  assign new_n1364_ = new_n2136_ | new_n2137_;
  assign new_n1365_ = new_n1364_ & new_n1362_;
  assign new_n1366_ = new_n1363_ | new_n1361_;
  assign new_n1367_ = new_n1365_ | new_n1352_;
  assign new_n1368_ = new_n1366_ | new_n1351_;
  assign new_n1369_ = new_n1368_ & new_n1367_;
  assign new_n1370_ = new_n2140_ & new_n2142_;
  assign new_n1371_ = new_n2144_ | new_n2145_;
  assign new_n1372_ = new_n2144_ & new_n2145_;
  assign new_n1373_ = new_n2140_ | new_n2142_;
  assign new_n1374_ = new_n1373_ & new_n1371_;
  assign new_n1375_ = new_n1372_ | new_n1370_;
  assign new_n1376_ = new_n2146_ & new_n2148_;
  assign new_n1377_ = new_n2150_ | new_n2151_;
  assign new_n1378_ = new_n2150_ & new_n2151_;
  assign new_n1379_ = new_n2146_ | new_n2148_;
  assign new_n1380_ = new_n1379_ & new_n1377_;
  assign new_n1381_ = new_n1378_ | new_n1376_;
  assign new_n1382_ = new_n2152_ & new_n2153_;
  assign new_n1383_ = new_n2154_ | new_n2155_;
  assign new_n1384_ = new_n2154_ & new_n2155_;
  assign new_n1385_ = new_n2152_ | new_n2153_;
  assign new_n1386_ = new_n1385_ & new_n1383_;
  assign new_n1387_ = new_n1384_ | new_n1382_;
  assign new_n1388_ = new_n1980_ & new_n822_;
  assign new_n1389_ = new_n1987_ | new_n823_;
  assign new_n1390_ = new_n2135_ & new_n2097_;
  assign new_n1391_ = new_n2129_ | new_n2103_;
  assign new_n1392_ = new_n2129_ & new_n2103_;
  assign new_n1393_ = new_n2135_ | new_n2097_;
  assign new_n1394_ = new_n1393_ & new_n1391_;
  assign new_n1395_ = new_n1392_ | new_n1390_;
  assign new_n1396_ = new_n2156_ & new_n2157_;
  assign new_n1397_ = new_n2158_ | new_n2159_;
  assign new_n1398_ = new_n2158_ & new_n2159_;
  assign new_n1399_ = new_n2156_ | new_n2157_;
  assign new_n1400_ = new_n1399_ & new_n1397_;
  assign new_n1401_ = new_n1398_ | new_n1396_;
  assign new_n1402_ = new_n1400_ | new_n1387_;
  assign new_n1403_ = new_n1401_ | new_n1386_;
  assign new_n1404_ = new_n1403_ & new_n1402_;
  assign new_n1405_ = new_n2160_ & new_n2162_;
  assign new_n1406_ = new_n2164_ | new_n2165_;
  assign new_n1407_ = new_n2164_ & new_n2165_;
  assign new_n1408_ = new_n2160_ | new_n2162_;
  assign new_n1409_ = new_n1408_ & new_n1406_;
  assign new_n1410_ = new_n1407_ | new_n1405_;
  assign new_n1411_ = new_n2166_ & new_n2168_;
  assign new_n1412_ = new_n2170_ | new_n2171_;
  assign new_n1413_ = new_n2170_ & new_n2171_;
  assign new_n1414_ = new_n2166_ | new_n2168_;
  assign new_n1415_ = new_n1414_ & new_n1412_;
  assign new_n1416_ = new_n1413_ | new_n1411_;
  assign new_n1417_ = new_n2172_ & new_n2173_;
  assign new_n1418_ = new_n2174_ | new_n2175_;
  assign new_n1419_ = new_n2174_ & new_n2175_;
  assign new_n1420_ = new_n2172_ | new_n2173_;
  assign new_n1421_ = new_n1420_ & new_n1418_;
  assign new_n1422_ = new_n1419_ | new_n1417_;
  assign new_n1423_ = new_n1980_ & new_n824_;
  assign new_n1424_ = new_n1987_ | new_n825_;
  assign new_n1425_ = new_n2126_ & new_n2100_;
  assign new_n1426_ = new_n2132_ | new_n2094_;
  assign new_n1427_ = new_n2132_ & new_n2094_;
  assign new_n1428_ = new_n2126_ | new_n2100_;
  assign new_n1429_ = new_n1428_ & new_n1426_;
  assign new_n1430_ = new_n1427_ | new_n1425_;
  assign new_n1431_ = new_n2176_ & new_n2177_;
  assign new_n1432_ = new_n2178_ | new_n2179_;
  assign new_n1433_ = new_n2178_ & new_n2179_;
  assign new_n1434_ = new_n2176_ | new_n2177_;
  assign new_n1435_ = new_n1434_ & new_n1432_;
  assign new_n1436_ = new_n1433_ | new_n1431_;
  assign new_n1437_ = new_n1435_ | new_n1422_;
  assign new_n1438_ = new_n1436_ | new_n1421_;
  assign new_n1439_ = new_n1438_ & new_n1437_;
  assign new_n1440_ = new_n2180_ & new_n2182_;
  assign new_n1441_ = new_n2184_ | new_n2185_;
  assign new_n1442_ = new_n2184_ & new_n2185_;
  assign new_n1443_ = new_n2180_ | new_n2182_;
  assign new_n1444_ = new_n1443_ & new_n1441_;
  assign new_n1445_ = new_n1442_ | new_n1440_;
  assign new_n1446_ = new_n2186_ & new_n2188_;
  assign new_n1447_ = new_n2190_ | new_n2191_;
  assign new_n1448_ = new_n2190_ & new_n2191_;
  assign new_n1449_ = new_n2186_ | new_n2188_;
  assign new_n1450_ = new_n1449_ & new_n1447_;
  assign new_n1451_ = new_n1448_ | new_n1446_;
  assign new_n1452_ = new_n1450_ | new_n1445_;
  assign new_n1453_ = new_n1451_ | new_n1444_;
  assign new_n1454_ = new_n1453_ & new_n1452_;
  assign new_n1455_ = new_n2192_ & new_n2194_;
  assign new_n1456_ = new_n2196_ | new_n2197_;
  assign new_n1457_ = new_n2196_ & new_n2197_;
  assign new_n1458_ = new_n2192_ | new_n2194_;
  assign new_n1459_ = new_n1458_ & new_n1456_;
  assign new_n1460_ = new_n1457_ | new_n1455_;
  assign new_n1461_ = new_n2198_ & new_n2200_;
  assign new_n1462_ = new_n2202_ | new_n2203_;
  assign new_n1463_ = new_n2202_ & new_n2203_;
  assign new_n1464_ = new_n2198_ | new_n2200_;
  assign new_n1465_ = new_n1464_ & new_n1462_;
  assign new_n1466_ = new_n1463_ | new_n1461_;
  assign new_n1467_ = new_n1465_ | new_n1460_;
  assign new_n1468_ = new_n1466_ | new_n1459_;
  assign new_n1469_ = new_n1468_ & new_n1467_;
  assign new_n1470_ = new_n2204_ & new_n2206_;
  assign new_n1471_ = new_n2208_ | new_n2209_;
  assign new_n1472_ = new_n2208_ & new_n2209_;
  assign new_n1473_ = new_n2204_ | new_n2206_;
  assign new_n1474_ = new_n1473_ & new_n1471_;
  assign new_n1475_ = new_n1472_ | new_n1470_;
  assign new_n1476_ = new_n2210_ & new_n2212_;
  assign new_n1477_ = new_n2214_ | new_n2215_;
  assign new_n1478_ = new_n2214_ & new_n2215_;
  assign new_n1479_ = new_n2210_ | new_n2212_;
  assign new_n1480_ = new_n1479_ & new_n1477_;
  assign new_n1481_ = new_n1478_ | new_n1476_;
  assign new_n1482_ = new_n1480_ | new_n1475_;
  assign new_n1483_ = new_n1481_ | new_n1474_;
  assign new_n1484_ = new_n1483_ & new_n1482_;
  assign new_n1485_ = new_n2216_ & new_n2218_;
  assign new_n1486_ = new_n2220_ | new_n2221_;
  assign new_n1487_ = new_n2220_ & new_n2221_;
  assign new_n1488_ = new_n2216_ | new_n2218_;
  assign new_n1489_ = new_n1488_ & new_n1486_;
  assign new_n1490_ = new_n1487_ | new_n1485_;
  assign new_n1491_ = new_n2222_ & new_n2224_;
  assign new_n1492_ = new_n2226_ | new_n2227_;
  assign new_n1493_ = new_n2226_ & new_n2227_;
  assign new_n1494_ = new_n2222_ | new_n2224_;
  assign new_n1495_ = new_n1494_ & new_n1492_;
  assign new_n1496_ = new_n1493_ | new_n1491_;
  assign new_n1497_ = new_n1495_ | new_n1490_;
  assign new_n1498_ = new_n1496_ | new_n1489_;
  assign new_n1499_ = new_n1498_ & new_n1497_;
  assign new_n1500_ = new_n2228_ & new_n2230_;
  assign new_n1501_ = new_n2232_ | new_n2233_;
  assign new_n1502_ = new_n2232_ & new_n2233_;
  assign new_n1503_ = new_n2228_ | new_n2230_;
  assign new_n1504_ = new_n1503_ & new_n1501_;
  assign new_n1505_ = new_n1502_ | new_n1500_;
  assign new_n1506_ = new_n2234_ & new_n2236_;
  assign new_n1507_ = new_n2238_ | new_n2239_;
  assign new_n1508_ = new_n2238_ & new_n2239_;
  assign new_n1509_ = new_n2234_ | new_n2236_;
  assign new_n1510_ = new_n1509_ & new_n1507_;
  assign new_n1511_ = new_n1508_ | new_n1506_;
  assign new_n1512_ = new_n1510_ | new_n1505_;
  assign new_n1513_ = new_n1511_ | new_n1504_;
  assign new_n1514_ = new_n1513_ & new_n1512_;
  assign new_n1515_ = new_n2240_ & new_n2242_;
  assign new_n1516_ = new_n2244_ | new_n2245_;
  assign new_n1517_ = new_n2244_ & new_n2245_;
  assign new_n1518_ = new_n2240_ | new_n2242_;
  assign new_n1519_ = new_n1518_ & new_n1516_;
  assign new_n1520_ = new_n1517_ | new_n1515_;
  assign new_n1521_ = new_n2246_ & new_n2248_;
  assign new_n1522_ = new_n2250_ | new_n2251_;
  assign new_n1523_ = new_n2250_ & new_n2251_;
  assign new_n1524_ = new_n2246_ | new_n2248_;
  assign new_n1525_ = new_n1524_ & new_n1522_;
  assign new_n1526_ = new_n1523_ | new_n1521_;
  assign new_n1527_ = new_n1525_ | new_n1520_;
  assign new_n1528_ = new_n1526_ | new_n1519_;
  assign new_n1529_ = new_n1528_ & new_n1527_;
  assign new_n1530_ = new_n2252_ & new_n2254_;
  assign new_n1531_ = new_n2256_ | new_n2257_;
  assign new_n1532_ = new_n2256_ & new_n2257_;
  assign new_n1533_ = new_n2252_ | new_n2254_;
  assign new_n1534_ = new_n1533_ & new_n1531_;
  assign new_n1535_ = new_n1532_ | new_n1530_;
  assign new_n1536_ = new_n2258_ & new_n2260_;
  assign new_n1537_ = new_n2262_ | new_n2263_;
  assign new_n1538_ = new_n2262_ & new_n2263_;
  assign new_n1539_ = new_n2258_ | new_n2260_;
  assign new_n1540_ = new_n1539_ & new_n1537_;
  assign new_n1541_ = new_n1538_ | new_n1536_;
  assign new_n1542_ = new_n1540_ | new_n1535_;
  assign new_n1543_ = new_n1541_ | new_n1534_;
  assign new_n1544_ = new_n1543_ & new_n1542_;
  assign new_n1545_ = new_n2264_ & new_n2266_;
  assign new_n1546_ = new_n2268_ | new_n2269_;
  assign new_n1547_ = new_n2268_ & new_n2269_;
  assign new_n1548_ = new_n2264_ | new_n2266_;
  assign new_n1549_ = new_n1548_ & new_n1546_;
  assign new_n1550_ = new_n1547_ | new_n1545_;
  assign new_n1551_ = new_n2270_ & new_n2272_;
  assign new_n1552_ = new_n2274_ | new_n2275_;
  assign new_n1553_ = new_n2274_ & new_n2275_;
  assign new_n1554_ = new_n2270_ | new_n2272_;
  assign new_n1555_ = new_n1554_ & new_n1552_;
  assign new_n1556_ = new_n1553_ | new_n1551_;
  assign new_n1557_ = new_n1555_ | new_n1550_;
  assign new_n1558_ = new_n1556_ | new_n1549_;
  assign new_n1559_ = new_n1558_ & new_n1557_;
  assign G468 = ~new_n920_;
  assign G469 = ~new_n925_;
  assign G470 = ~new_n930_;
  assign G471 = ~new_n935_;
  assign G472 = ~new_n948_;
  assign G473 = ~new_n953_;
  assign G474 = ~new_n958_;
  assign G475 = ~new_n963_;
  assign G476 = ~new_n976_;
  assign G477 = ~new_n981_;
  assign G478 = ~new_n986_;
  assign G479 = ~new_n991_;
  assign G480 = ~new_n1004_;
  assign G481 = ~new_n1009_;
  assign G482 = ~new_n1014_;
  assign G483 = ~new_n1019_;
  assign G484 = ~new_n1032_;
  assign G485 = ~new_n1037_;
  assign G486 = ~new_n1042_;
  assign G487 = ~new_n1047_;
  assign G488 = ~new_n1060_;
  assign G489 = ~new_n1065_;
  assign G490 = ~new_n1070_;
  assign G491 = ~new_n1075_;
  assign G492 = ~new_n1088_;
  assign G493 = ~new_n1093_;
  assign G494 = ~new_n1098_;
  assign G495 = ~new_n1103_;
  assign G496 = ~new_n1116_;
  assign G497 = ~new_n1121_;
  assign G498 = ~new_n1126_;
  assign G499 = ~new_n1131_;
  assign n286_li = ~new_n631_;
  assign n298_li = ~new_n633_;
  assign n310_li = ~new_n635_;
  assign n322_li = ~new_n637_;
  assign n334_li = ~new_n639_;
  assign n346_li = ~new_n641_;
  assign n358_li = ~new_n643_;
  assign n370_li = ~new_n645_;
  assign n382_li = ~new_n647_;
  assign n394_li = ~new_n649_;
  assign n406_li = ~new_n651_;
  assign n418_li = ~new_n653_;
  assign n430_li = ~new_n655_;
  assign n442_li = ~new_n657_;
  assign n454_li = ~new_n659_;
  assign n466_li = ~new_n661_;
  assign n478_li = ~new_n663_;
  assign n490_li = ~new_n665_;
  assign n502_li = ~new_n667_;
  assign n514_li = ~new_n669_;
  assign n526_li = ~new_n671_;
  assign n538_li = ~new_n673_;
  assign n550_li = ~new_n675_;
  assign n562_li = ~new_n677_;
  assign n574_li = ~new_n679_;
  assign n586_li = ~new_n681_;
  assign n598_li = ~new_n683_;
  assign n610_li = ~new_n685_;
  assign n622_li = ~new_n687_;
  assign n634_li = ~new_n689_;
  assign n646_li = ~new_n691_;
  assign n658_li = ~new_n693_;
  assign n661_li = ~new_n515_;
  assign n673_li = ~new_n517_;
  assign n685_li = ~new_n519_;
  assign n697_li = ~new_n521_;
  assign n709_li = ~new_n523_;
  assign n721_li = ~new_n525_;
  assign n733_li = ~new_n527_;
  assign n745_li = ~new_n529_;
  assign n757_li = ~new_n531_;
  assign n1248_i2 = ~new_n1937_;
  assign n1249_i2 = ~new_n1934_;
  assign n1250_i2 = ~new_n1929_;
  assign n1251_i2 = ~new_n1926_;
  assign n1252_i2 = ~new_n1956_;
  assign n1253_i2 = ~new_n1953_;
  assign n1254_i2 = ~new_n1948_;
  assign n1255_i2 = ~new_n1945_;
  assign n1207_i2 = ~new_n1959_;
  assign n1208_i2 = ~new_n2005_;
  assign n1209_i2 = ~new_n2037_;
  assign n1210_i2 = ~new_n2057_;
  assign n1211_i2 = ~new_n1961_;
  assign n1212_i2 = ~new_n2007_;
  assign n1213_i2 = ~new_n2039_;
  assign n1214_i2 = ~new_n2059_;
  assign n1215_i2 = ~new_n1965_;
  assign n1216_i2 = ~new_n2011_;
  assign n1217_i2 = ~new_n2043_;
  assign n1218_i2 = ~new_n2063_;
  assign n1219_i2 = ~new_n1967_;
  assign n1220_i2 = ~new_n2013_;
  assign n1221_i2 = ~new_n2045_;
  assign n1222_i2 = ~new_n2065_;
  assign n1223_i2 = ~new_n2077_;
  assign n1224_i2 = ~new_n2109_;
  assign n1225_i2 = ~new_n2141_;
  assign n1226_i2 = ~new_n2161_;
  assign n1227_i2 = ~new_n2079_;
  assign n1228_i2 = ~new_n2111_;
  assign n1229_i2 = ~new_n2143_;
  assign n1230_i2 = ~new_n2163_;
  assign n1231_i2 = ~new_n2083_;
  assign n1232_i2 = ~new_n2115_;
  assign n1233_i2 = ~new_n2147_;
  assign n1234_i2 = ~new_n2167_;
  assign n1235_i2 = ~new_n2085_;
  assign n1236_i2 = ~new_n2117_;
  assign n1237_i2 = ~new_n2149_;
  assign n1238_i2 = ~new_n2169_;
  assign G374_i2 = ~new_n1938_;
  assign G376_i2 = G374_i2;
  assign G370_i2 = ~new_n1935_;
  assign G372_i2 = G370_i2;
  assign G373_i2 = ~new_n1930_;
  assign G377_i2 = G373_i2;
  assign G371_i2 = ~new_n1927_;
  assign G375_i2 = G371_i2;
  assign G354_i2 = ~new_n1957_;
  assign G356_i2 = G354_i2;
  assign G350_i2 = ~new_n1954_;
  assign G352_i2 = G350_i2;
  assign G353_i2 = ~new_n1949_;
  assign G357_i2 = G353_i2;
  assign G351_i2 = ~new_n1946_;
  assign G355_i2 = G351_i2;
  assign G386_i2 = ~new_n1145_;
  assign G391_i2 = ~new_n1159_;
  assign n283_lo_buf_i2 = ~new_n2181_;
  assign n295_lo_buf_i2 = ~new_n2183_;
  assign n307_lo_buf_i2 = ~new_n2187_;
  assign n319_lo_buf_i2 = ~new_n2189_;
  assign n331_lo_buf_i2 = ~new_n2193_;
  assign n343_lo_buf_i2 = ~new_n2195_;
  assign n355_lo_buf_i2 = ~new_n2199_;
  assign n367_lo_buf_i2 = ~new_n2201_;
  assign n379_lo_buf_i2 = ~new_n2205_;
  assign n391_lo_buf_i2 = ~new_n2207_;
  assign n403_lo_buf_i2 = ~new_n2211_;
  assign n415_lo_buf_i2 = ~new_n2213_;
  assign n427_lo_buf_i2 = ~new_n2217_;
  assign n439_lo_buf_i2 = ~new_n2219_;
  assign n451_lo_buf_i2 = ~new_n2223_;
  assign n463_lo_buf_i2 = ~new_n2225_;
  assign n475_lo_buf_i2 = ~new_n2229_;
  assign n487_lo_buf_i2 = ~new_n2231_;
  assign n499_lo_buf_i2 = ~new_n2235_;
  assign n511_lo_buf_i2 = ~new_n2237_;
  assign n523_lo_buf_i2 = ~new_n2241_;
  assign n535_lo_buf_i2 = ~new_n2243_;
  assign n547_lo_buf_i2 = ~new_n2247_;
  assign n559_lo_buf_i2 = ~new_n2249_;
  assign n571_lo_buf_i2 = ~new_n2253_;
  assign n583_lo_buf_i2 = ~new_n2255_;
  assign n595_lo_buf_i2 = ~new_n2259_;
  assign n607_lo_buf_i2 = ~new_n2261_;
  assign n619_lo_buf_i2 = ~new_n2265_;
  assign n631_lo_buf_i2 = ~new_n2267_;
  assign n643_lo_buf_i2 = ~new_n2271_;
  assign n655_lo_buf_i2 = ~new_n2273_;
  assign G234_i2 = ~new_n1194_;
  assign G247_i2 = ~new_n1229_;
  assign G260_i2 = ~new_n1264_;
  assign G273_i2 = ~new_n1299_;
  assign G286_i2 = ~new_n1334_;
  assign G299_i2 = ~new_n1369_;
  assign G312_i2 = ~new_n1404_;
  assign G325_i2 = ~new_n1439_;
  assign n667_lo_buf_i2 = ~new_n597_;
  assign n679_lo_buf_i2 = ~new_n599_;
  assign n691_lo_buf_i2 = ~new_n601_;
  assign n703_lo_buf_i2 = ~new_n603_;
  assign n715_lo_buf_i2 = ~new_n605_;
  assign n727_lo_buf_i2 = ~new_n607_;
  assign n739_lo_buf_i2 = ~new_n609_;
  assign n751_lo_buf_i2 = ~new_n611_;
  assign n763_lo_buf_i2 = ~new_n613_;
  assign G186_i2 = ~new_n1454_;
  assign G189_i2 = ~new_n1469_;
  assign G192_i2 = ~new_n1484_;
  assign G195_i2 = ~new_n1499_;
  assign G198_i2 = ~new_n1514_;
  assign G201_i2 = ~new_n1529_;
  assign G204_i2 = ~new_n1544_;
  assign G207_i2 = ~new_n1559_;
  assign n280_lo_buf_i2 = ~new_n451_;
  assign n292_lo_buf_i2 = ~new_n453_;
  assign n304_lo_buf_i2 = ~new_n455_;
  assign n316_lo_buf_i2 = ~new_n457_;
  assign n328_lo_buf_i2 = ~new_n459_;
  assign n340_lo_buf_i2 = ~new_n461_;
  assign n352_lo_buf_i2 = ~new_n463_;
  assign n364_lo_buf_i2 = ~new_n465_;
  assign n376_lo_buf_i2 = ~new_n467_;
  assign n388_lo_buf_i2 = ~new_n469_;
  assign n400_lo_buf_i2 = ~new_n471_;
  assign n412_lo_buf_i2 = ~new_n473_;
  assign n424_lo_buf_i2 = ~new_n475_;
  assign n436_lo_buf_i2 = ~new_n477_;
  assign n448_lo_buf_i2 = ~new_n479_;
  assign n460_lo_buf_i2 = ~new_n481_;
  assign n472_lo_buf_i2 = ~new_n483_;
  assign n484_lo_buf_i2 = ~new_n485_;
  assign n496_lo_buf_i2 = ~new_n487_;
  assign n508_lo_buf_i2 = ~new_n489_;
  assign n520_lo_buf_i2 = ~new_n491_;
  assign n532_lo_buf_i2 = ~new_n493_;
  assign n544_lo_buf_i2 = ~new_n495_;
  assign n556_lo_buf_i2 = ~new_n497_;
  assign n568_lo_buf_i2 = ~new_n499_;
  assign n580_lo_buf_i2 = ~new_n501_;
  assign n592_lo_buf_i2 = ~new_n503_;
  assign n604_lo_buf_i2 = ~new_n505_;
  assign n616_lo_buf_i2 = ~new_n507_;
  assign n628_lo_buf_i2 = ~new_n509_;
  assign n640_lo_buf_i2 = ~new_n511_;
  assign n652_lo_buf_i2 = ~new_n513_;
  assign new_n1780_ = new_n622_;
  assign new_n1781_ = new_n1780_;
  assign new_n1782_ = new_n1781_;
  assign new_n1783_ = new_n1781_;
  assign new_n1784_ = new_n1780_;
  assign new_n1785_ = new_n623_;
  assign new_n1786_ = new_n1785_;
  assign new_n1787_ = new_n1786_;
  assign new_n1788_ = new_n1786_;
  assign new_n1789_ = new_n1785_;
  assign new_n1790_ = new_n626_;
  assign new_n1791_ = new_n1790_;
  assign new_n1792_ = new_n1791_;
  assign new_n1793_ = new_n1791_;
  assign new_n1794_ = new_n1790_;
  assign new_n1795_ = new_n627_;
  assign new_n1796_ = new_n1795_;
  assign new_n1797_ = new_n1796_;
  assign new_n1798_ = new_n1796_;
  assign new_n1799_ = new_n1795_;
  assign new_n1800_ = new_n726_;
  assign new_n1801_ = new_n1800_;
  assign new_n1802_ = new_n1800_;
  assign new_n1803_ = new_n727_;
  assign new_n1804_ = new_n1803_;
  assign new_n1805_ = new_n1803_;
  assign new_n1806_ = new_n914_;
  assign new_n1807_ = new_n1806_;
  assign new_n1808_ = new_n1806_;
  assign new_n1809_ = new_n614_;
  assign new_n1810_ = new_n1809_;
  assign new_n1811_ = new_n1810_;
  assign new_n1812_ = new_n1810_;
  assign new_n1813_ = new_n1809_;
  assign new_n1814_ = new_n915_;
  assign new_n1815_ = new_n1814_;
  assign new_n1816_ = new_n1814_;
  assign new_n1817_ = new_n615_;
  assign new_n1818_ = new_n1817_;
  assign new_n1819_ = new_n1818_;
  assign new_n1820_ = new_n1818_;
  assign new_n1821_ = new_n1817_;
  assign new_n1822_ = new_n616_;
  assign new_n1823_ = new_n1822_;
  assign new_n1824_ = new_n1823_;
  assign new_n1825_ = new_n1823_;
  assign new_n1826_ = new_n1822_;
  assign new_n1827_ = new_n617_;
  assign new_n1828_ = new_n1827_;
  assign new_n1829_ = new_n1828_;
  assign new_n1830_ = new_n1828_;
  assign new_n1831_ = new_n1827_;
  assign new_n1832_ = new_n618_;
  assign new_n1833_ = new_n1832_;
  assign new_n1834_ = new_n1833_;
  assign new_n1835_ = new_n1833_;
  assign new_n1836_ = new_n1832_;
  assign new_n1837_ = new_n619_;
  assign new_n1838_ = new_n1837_;
  assign new_n1839_ = new_n1838_;
  assign new_n1840_ = new_n1838_;
  assign new_n1841_ = new_n1837_;
  assign new_n1842_ = new_n620_;
  assign new_n1843_ = new_n1842_;
  assign new_n1844_ = new_n1843_;
  assign new_n1845_ = new_n1843_;
  assign new_n1846_ = new_n1842_;
  assign new_n1847_ = new_n621_;
  assign new_n1848_ = new_n1847_;
  assign new_n1849_ = new_n1848_;
  assign new_n1850_ = new_n1848_;
  assign new_n1851_ = new_n1847_;
  assign new_n1852_ = new_n628_;
  assign new_n1853_ = new_n1852_;
  assign new_n1854_ = new_n1853_;
  assign new_n1855_ = new_n1853_;
  assign new_n1856_ = new_n1852_;
  assign new_n1857_ = new_n629_;
  assign new_n1858_ = new_n1857_;
  assign new_n1859_ = new_n1858_;
  assign new_n1860_ = new_n1858_;
  assign new_n1861_ = new_n1857_;
  assign new_n1862_ = new_n942_;
  assign new_n1863_ = new_n1862_;
  assign new_n1864_ = new_n1862_;
  assign new_n1865_ = new_n943_;
  assign new_n1866_ = new_n1865_;
  assign new_n1867_ = new_n1865_;
  assign new_n1868_ = new_n624_;
  assign new_n1869_ = new_n1868_;
  assign new_n1870_ = new_n1869_;
  assign new_n1871_ = new_n1869_;
  assign new_n1872_ = new_n1868_;
  assign new_n1873_ = new_n625_;
  assign new_n1874_ = new_n1873_;
  assign new_n1875_ = new_n1874_;
  assign new_n1876_ = new_n1874_;
  assign new_n1877_ = new_n1873_;
  assign new_n1878_ = new_n970_;
  assign new_n1879_ = new_n1878_;
  assign new_n1880_ = new_n1878_;
  assign new_n1881_ = new_n971_;
  assign new_n1882_ = new_n1881_;
  assign new_n1883_ = new_n1881_;
  assign new_n1884_ = new_n998_;
  assign new_n1885_ = new_n1884_;
  assign new_n1886_ = new_n1884_;
  assign new_n1887_ = new_n999_;
  assign new_n1888_ = new_n1887_;
  assign new_n1889_ = new_n1887_;
  assign new_n1890_ = new_n728_;
  assign new_n1891_ = new_n1890_;
  assign new_n1892_ = new_n1890_;
  assign new_n1893_ = new_n729_;
  assign new_n1894_ = new_n1893_;
  assign new_n1895_ = new_n1893_;
  assign new_n1896_ = new_n1026_;
  assign new_n1897_ = new_n1896_;
  assign new_n1898_ = new_n1896_;
  assign new_n1899_ = new_n1027_;
  assign new_n1900_ = new_n1899_;
  assign new_n1901_ = new_n1899_;
  assign new_n1902_ = new_n1054_;
  assign new_n1903_ = new_n1902_;
  assign new_n1904_ = new_n1902_;
  assign new_n1905_ = new_n1055_;
  assign new_n1906_ = new_n1905_;
  assign new_n1907_ = new_n1905_;
  assign new_n1908_ = new_n1082_;
  assign new_n1909_ = new_n1908_;
  assign new_n1910_ = new_n1908_;
  assign new_n1911_ = new_n1083_;
  assign new_n1912_ = new_n1911_;
  assign new_n1913_ = new_n1911_;
  assign new_n1914_ = new_n1110_;
  assign new_n1915_ = new_n1914_;
  assign new_n1916_ = new_n1914_;
  assign new_n1917_ = new_n1111_;
  assign new_n1918_ = new_n1917_;
  assign new_n1919_ = new_n1917_;
  assign new_n1920_ = new_n796_;
  assign new_n1921_ = new_n794_;
  assign new_n1922_ = new_n1132_;
  assign new_n1923_ = new_n798_;
  assign new_n1924_ = new_n1923_;
  assign new_n1925_ = new_n801_;
  assign new_n1926_ = new_n1925_;
  assign new_n1927_ = new_n1925_;
  assign new_n1928_ = new_n799_;
  assign new_n1929_ = new_n1928_;
  assign new_n1930_ = new_n1928_;
  assign new_n1931_ = new_n800_;
  assign new_n1932_ = new_n1931_;
  assign new_n1933_ = new_n797_;
  assign new_n1934_ = new_n1933_;
  assign new_n1935_ = new_n1933_;
  assign new_n1936_ = new_n795_;
  assign new_n1937_ = new_n1936_;
  assign new_n1938_ = new_n1936_;
  assign new_n1939_ = new_n804_;
  assign new_n1940_ = new_n802_;
  assign new_n1941_ = new_n1146_;
  assign new_n1942_ = new_n806_;
  assign new_n1943_ = new_n1942_;
  assign new_n1944_ = new_n809_;
  assign new_n1945_ = new_n1944_;
  assign new_n1946_ = new_n1944_;
  assign new_n1947_ = new_n807_;
  assign new_n1948_ = new_n1947_;
  assign new_n1949_ = new_n1947_;
  assign new_n1950_ = new_n808_;
  assign new_n1951_ = new_n1950_;
  assign new_n1952_ = new_n805_;
  assign new_n1953_ = new_n1952_;
  assign new_n1954_ = new_n1952_;
  assign new_n1955_ = new_n803_;
  assign new_n1956_ = new_n1955_;
  assign new_n1957_ = new_n1955_;
  assign new_n1958_ = new_n738_;
  assign new_n1959_ = new_n731_;
  assign new_n1960_ = new_n1959_;
  assign new_n1961_ = new_n739_;
  assign new_n1962_ = new_n1961_;
  assign new_n1963_ = new_n730_;
  assign new_n1964_ = new_n754_;
  assign new_n1965_ = new_n747_;
  assign new_n1966_ = new_n1965_;
  assign new_n1967_ = new_n755_;
  assign new_n1968_ = new_n1967_;
  assign new_n1969_ = new_n746_;
  assign new_n1970_ = new_n1171_;
  assign new_n1971_ = new_n1164_;
  assign new_n1972_ = new_n1170_;
  assign new_n1973_ = new_n1165_;
  assign new_n1974_ = new_n826_;
  assign new_n1975_ = new_n1974_;
  assign new_n1976_ = new_n1975_;
  assign new_n1977_ = new_n1975_;
  assign new_n1978_ = new_n1974_;
  assign new_n1979_ = new_n1978_;
  assign new_n1980_ = new_n1978_;
  assign new_n1981_ = new_n827_;
  assign new_n1982_ = new_n1981_;
  assign new_n1983_ = new_n1982_;
  assign new_n1984_ = new_n1982_;
  assign new_n1985_ = new_n1981_;
  assign new_n1986_ = new_n1985_;
  assign new_n1987_ = new_n1985_;
  assign new_n1988_ = new_n838_;
  assign new_n1989_ = new_n1988_;
  assign new_n1990_ = new_n1988_;
  assign new_n1991_ = new_n837_;
  assign new_n1992_ = new_n1991_;
  assign new_n1993_ = new_n1991_;
  assign new_n1994_ = new_n839_;
  assign new_n1995_ = new_n1994_;
  assign new_n1996_ = new_n1994_;
  assign new_n1997_ = new_n836_;
  assign new_n1998_ = new_n1997_;
  assign new_n1999_ = new_n1997_;
  assign new_n2000_ = new_n1185_;
  assign new_n2001_ = new_n1179_;
  assign new_n2002_ = new_n1184_;
  assign new_n2003_ = new_n1178_;
  assign new_n2004_ = new_n740_;
  assign new_n2005_ = new_n733_;
  assign new_n2006_ = new_n2005_;
  assign new_n2007_ = new_n741_;
  assign new_n2008_ = new_n2007_;
  assign new_n2009_ = new_n732_;
  assign new_n2010_ = new_n756_;
  assign new_n2011_ = new_n749_;
  assign new_n2012_ = new_n2011_;
  assign new_n2013_ = new_n757_;
  assign new_n2014_ = new_n2013_;
  assign new_n2015_ = new_n748_;
  assign new_n2016_ = new_n1206_;
  assign new_n2017_ = new_n1199_;
  assign new_n2018_ = new_n1205_;
  assign new_n2019_ = new_n1200_;
  assign new_n2020_ = new_n842_;
  assign new_n2021_ = new_n2020_;
  assign new_n2022_ = new_n2020_;
  assign new_n2023_ = new_n841_;
  assign new_n2024_ = new_n2023_;
  assign new_n2025_ = new_n2023_;
  assign new_n2026_ = new_n843_;
  assign new_n2027_ = new_n2026_;
  assign new_n2028_ = new_n2026_;
  assign new_n2029_ = new_n840_;
  assign new_n2030_ = new_n2029_;
  assign new_n2031_ = new_n2029_;
  assign new_n2032_ = new_n1220_;
  assign new_n2033_ = new_n1214_;
  assign new_n2034_ = new_n1219_;
  assign new_n2035_ = new_n1213_;
  assign new_n2036_ = new_n742_;
  assign new_n2037_ = new_n735_;
  assign new_n2038_ = new_n2037_;
  assign new_n2039_ = new_n743_;
  assign new_n2040_ = new_n2039_;
  assign new_n2041_ = new_n734_;
  assign new_n2042_ = new_n758_;
  assign new_n2043_ = new_n751_;
  assign new_n2044_ = new_n2043_;
  assign new_n2045_ = new_n759_;
  assign new_n2046_ = new_n2045_;
  assign new_n2047_ = new_n750_;
  assign new_n2048_ = new_n1241_;
  assign new_n2049_ = new_n1234_;
  assign new_n2050_ = new_n1240_;
  assign new_n2051_ = new_n1235_;
  assign new_n2052_ = new_n1255_;
  assign new_n2053_ = new_n1249_;
  assign new_n2054_ = new_n1254_;
  assign new_n2055_ = new_n1248_;
  assign new_n2056_ = new_n744_;
  assign new_n2057_ = new_n737_;
  assign new_n2058_ = new_n2057_;
  assign new_n2059_ = new_n745_;
  assign new_n2060_ = new_n2059_;
  assign new_n2061_ = new_n736_;
  assign new_n2062_ = new_n760_;
  assign new_n2063_ = new_n753_;
  assign new_n2064_ = new_n2063_;
  assign new_n2065_ = new_n761_;
  assign new_n2066_ = new_n2065_;
  assign new_n2067_ = new_n752_;
  assign new_n2068_ = new_n1276_;
  assign new_n2069_ = new_n1269_;
  assign new_n2070_ = new_n1275_;
  assign new_n2071_ = new_n1270_;
  assign new_n2072_ = new_n1290_;
  assign new_n2073_ = new_n1284_;
  assign new_n2074_ = new_n1289_;
  assign new_n2075_ = new_n1283_;
  assign new_n2076_ = new_n770_;
  assign new_n2077_ = new_n763_;
  assign new_n2078_ = new_n2077_;
  assign new_n2079_ = new_n771_;
  assign new_n2080_ = new_n2079_;
  assign new_n2081_ = new_n762_;
  assign new_n2082_ = new_n786_;
  assign new_n2083_ = new_n779_;
  assign new_n2084_ = new_n2083_;
  assign new_n2085_ = new_n787_;
  assign new_n2086_ = new_n2085_;
  assign new_n2087_ = new_n778_;
  assign new_n2088_ = new_n1311_;
  assign new_n2089_ = new_n1304_;
  assign new_n2090_ = new_n1310_;
  assign new_n2091_ = new_n1305_;
  assign new_n2092_ = new_n830_;
  assign new_n2093_ = new_n2092_;
  assign new_n2094_ = new_n2092_;
  assign new_n2095_ = new_n829_;
  assign new_n2096_ = new_n2095_;
  assign new_n2097_ = new_n2095_;
  assign new_n2098_ = new_n831_;
  assign new_n2099_ = new_n2098_;
  assign new_n2100_ = new_n2098_;
  assign new_n2101_ = new_n828_;
  assign new_n2102_ = new_n2101_;
  assign new_n2103_ = new_n2101_;
  assign new_n2104_ = new_n1325_;
  assign new_n2105_ = new_n1319_;
  assign new_n2106_ = new_n1324_;
  assign new_n2107_ = new_n1318_;
  assign new_n2108_ = new_n772_;
  assign new_n2109_ = new_n765_;
  assign new_n2110_ = new_n2109_;
  assign new_n2111_ = new_n773_;
  assign new_n2112_ = new_n2111_;
  assign new_n2113_ = new_n764_;
  assign new_n2114_ = new_n788_;
  assign new_n2115_ = new_n781_;
  assign new_n2116_ = new_n2115_;
  assign new_n2117_ = new_n789_;
  assign new_n2118_ = new_n2117_;
  assign new_n2119_ = new_n780_;
  assign new_n2120_ = new_n1346_;
  assign new_n2121_ = new_n1339_;
  assign new_n2122_ = new_n1345_;
  assign new_n2123_ = new_n1340_;
  assign new_n2124_ = new_n834_;
  assign new_n2125_ = new_n2124_;
  assign new_n2126_ = new_n2124_;
  assign new_n2127_ = new_n833_;
  assign new_n2128_ = new_n2127_;
  assign new_n2129_ = new_n2127_;
  assign new_n2130_ = new_n835_;
  assign new_n2131_ = new_n2130_;
  assign new_n2132_ = new_n2130_;
  assign new_n2133_ = new_n832_;
  assign new_n2134_ = new_n2133_;
  assign new_n2135_ = new_n2133_;
  assign new_n2136_ = new_n1360_;
  assign new_n2137_ = new_n1354_;
  assign new_n2138_ = new_n1359_;
  assign new_n2139_ = new_n1353_;
  assign new_n2140_ = new_n774_;
  assign new_n2141_ = new_n767_;
  assign new_n2142_ = new_n2141_;
  assign new_n2143_ = new_n775_;
  assign new_n2144_ = new_n2143_;
  assign new_n2145_ = new_n766_;
  assign new_n2146_ = new_n790_;
  assign new_n2147_ = new_n783_;
  assign new_n2148_ = new_n2147_;
  assign new_n2149_ = new_n791_;
  assign new_n2150_ = new_n2149_;
  assign new_n2151_ = new_n782_;
  assign new_n2152_ = new_n1381_;
  assign new_n2153_ = new_n1374_;
  assign new_n2154_ = new_n1380_;
  assign new_n2155_ = new_n1375_;
  assign new_n2156_ = new_n1395_;
  assign new_n2157_ = new_n1389_;
  assign new_n2158_ = new_n1394_;
  assign new_n2159_ = new_n1388_;
  assign new_n2160_ = new_n776_;
  assign new_n2161_ = new_n769_;
  assign new_n2162_ = new_n2161_;
  assign new_n2163_ = new_n777_;
  assign new_n2164_ = new_n2163_;
  assign new_n2165_ = new_n768_;
  assign new_n2166_ = new_n792_;
  assign new_n2167_ = new_n785_;
  assign new_n2168_ = new_n2167_;
  assign new_n2169_ = new_n793_;
  assign new_n2170_ = new_n2169_;
  assign new_n2171_ = new_n784_;
  assign new_n2172_ = new_n1416_;
  assign new_n2173_ = new_n1409_;
  assign new_n2174_ = new_n1415_;
  assign new_n2175_ = new_n1410_;
  assign new_n2176_ = new_n1430_;
  assign new_n2177_ = new_n1424_;
  assign new_n2178_ = new_n1429_;
  assign new_n2179_ = new_n1423_;
  assign new_n2180_ = new_n846_;
  assign new_n2181_ = new_n845_;
  assign new_n2182_ = new_n2181_;
  assign new_n2183_ = new_n847_;
  assign new_n2184_ = new_n2183_;
  assign new_n2185_ = new_n844_;
  assign new_n2186_ = new_n850_;
  assign new_n2187_ = new_n849_;
  assign new_n2188_ = new_n2187_;
  assign new_n2189_ = new_n851_;
  assign new_n2190_ = new_n2189_;
  assign new_n2191_ = new_n848_;
  assign new_n2192_ = new_n854_;
  assign new_n2193_ = new_n853_;
  assign new_n2194_ = new_n2193_;
  assign new_n2195_ = new_n855_;
  assign new_n2196_ = new_n2195_;
  assign new_n2197_ = new_n852_;
  assign new_n2198_ = new_n858_;
  assign new_n2199_ = new_n857_;
  assign new_n2200_ = new_n2199_;
  assign new_n2201_ = new_n859_;
  assign new_n2202_ = new_n2201_;
  assign new_n2203_ = new_n856_;
  assign new_n2204_ = new_n862_;
  assign new_n2205_ = new_n861_;
  assign new_n2206_ = new_n2205_;
  assign new_n2207_ = new_n863_;
  assign new_n2208_ = new_n2207_;
  assign new_n2209_ = new_n860_;
  assign new_n2210_ = new_n866_;
  assign new_n2211_ = new_n865_;
  assign new_n2212_ = new_n2211_;
  assign new_n2213_ = new_n867_;
  assign new_n2214_ = new_n2213_;
  assign new_n2215_ = new_n864_;
  assign new_n2216_ = new_n870_;
  assign new_n2217_ = new_n869_;
  assign new_n2218_ = new_n2217_;
  assign new_n2219_ = new_n871_;
  assign new_n2220_ = new_n2219_;
  assign new_n2221_ = new_n868_;
  assign new_n2222_ = new_n874_;
  assign new_n2223_ = new_n873_;
  assign new_n2224_ = new_n2223_;
  assign new_n2225_ = new_n875_;
  assign new_n2226_ = new_n2225_;
  assign new_n2227_ = new_n872_;
  assign new_n2228_ = new_n878_;
  assign new_n2229_ = new_n877_;
  assign new_n2230_ = new_n2229_;
  assign new_n2231_ = new_n879_;
  assign new_n2232_ = new_n2231_;
  assign new_n2233_ = new_n876_;
  assign new_n2234_ = new_n882_;
  assign new_n2235_ = new_n881_;
  assign new_n2236_ = new_n2235_;
  assign new_n2237_ = new_n883_;
  assign new_n2238_ = new_n2237_;
  assign new_n2239_ = new_n880_;
  assign new_n2240_ = new_n886_;
  assign new_n2241_ = new_n885_;
  assign new_n2242_ = new_n2241_;
  assign new_n2243_ = new_n887_;
  assign new_n2244_ = new_n2243_;
  assign new_n2245_ = new_n884_;
  assign new_n2246_ = new_n890_;
  assign new_n2247_ = new_n889_;
  assign new_n2248_ = new_n2247_;
  assign new_n2249_ = new_n891_;
  assign new_n2250_ = new_n2249_;
  assign new_n2251_ = new_n888_;
  assign new_n2252_ = new_n894_;
  assign new_n2253_ = new_n893_;
  assign new_n2254_ = new_n2253_;
  assign new_n2255_ = new_n895_;
  assign new_n2256_ = new_n2255_;
  assign new_n2257_ = new_n892_;
  assign new_n2258_ = new_n898_;
  assign new_n2259_ = new_n897_;
  assign new_n2260_ = new_n2259_;
  assign new_n2261_ = new_n899_;
  assign new_n2262_ = new_n2261_;
  assign new_n2263_ = new_n896_;
  assign new_n2264_ = new_n902_;
  assign new_n2265_ = new_n901_;
  assign new_n2266_ = new_n2265_;
  assign new_n2267_ = new_n903_;
  assign new_n2268_ = new_n2267_;
  assign new_n2269_ = new_n900_;
  assign new_n2270_ = new_n906_;
  assign new_n2271_ = new_n905_;
  assign new_n2272_ = new_n2271_;
  assign new_n2273_ = new_n907_;
  assign new_n2274_ = new_n2273_;
  assign new_n2275_ = new_n904_;
  always @ (posedge clock) begin
    n286_lo <= n286_li;
    n298_lo <= n298_li;
    n310_lo <= n310_li;
    n322_lo <= n322_li;
    n334_lo <= n334_li;
    n346_lo <= n346_li;
    n358_lo <= n358_li;
    n370_lo <= n370_li;
    n382_lo <= n382_li;
    n394_lo <= n394_li;
    n406_lo <= n406_li;
    n418_lo <= n418_li;
    n430_lo <= n430_li;
    n442_lo <= n442_li;
    n454_lo <= n454_li;
    n466_lo <= n466_li;
    n478_lo <= n478_li;
    n490_lo <= n490_li;
    n502_lo <= n502_li;
    n514_lo <= n514_li;
    n526_lo <= n526_li;
    n538_lo <= n538_li;
    n550_lo <= n550_li;
    n562_lo <= n562_li;
    n574_lo <= n574_li;
    n586_lo <= n586_li;
    n598_lo <= n598_li;
    n610_lo <= n610_li;
    n622_lo <= n622_li;
    n634_lo <= n634_li;
    n646_lo <= n646_li;
    n658_lo <= n658_li;
    n661_lo <= n661_li;
    n673_lo <= n673_li;
    n685_lo <= n685_li;
    n697_lo <= n697_li;
    n709_lo <= n709_li;
    n721_lo <= n721_li;
    n733_lo <= n733_li;
    n745_lo <= n745_li;
    n757_lo <= n757_li;
    n1248_o2 <= n1248_i2;
    n1249_o2 <= n1249_i2;
    n1250_o2 <= n1250_i2;
    n1251_o2 <= n1251_i2;
    n1252_o2 <= n1252_i2;
    n1253_o2 <= n1253_i2;
    n1254_o2 <= n1254_i2;
    n1255_o2 <= n1255_i2;
    n1207_o2 <= n1207_i2;
    n1208_o2 <= n1208_i2;
    n1209_o2 <= n1209_i2;
    n1210_o2 <= n1210_i2;
    n1211_o2 <= n1211_i2;
    n1212_o2 <= n1212_i2;
    n1213_o2 <= n1213_i2;
    n1214_o2 <= n1214_i2;
    n1215_o2 <= n1215_i2;
    n1216_o2 <= n1216_i2;
    n1217_o2 <= n1217_i2;
    n1218_o2 <= n1218_i2;
    n1219_o2 <= n1219_i2;
    n1220_o2 <= n1220_i2;
    n1221_o2 <= n1221_i2;
    n1222_o2 <= n1222_i2;
    n1223_o2 <= n1223_i2;
    n1224_o2 <= n1224_i2;
    n1225_o2 <= n1225_i2;
    n1226_o2 <= n1226_i2;
    n1227_o2 <= n1227_i2;
    n1228_o2 <= n1228_i2;
    n1229_o2 <= n1229_i2;
    n1230_o2 <= n1230_i2;
    n1231_o2 <= n1231_i2;
    n1232_o2 <= n1232_i2;
    n1233_o2 <= n1233_i2;
    n1234_o2 <= n1234_i2;
    n1235_o2 <= n1235_i2;
    n1236_o2 <= n1236_i2;
    n1237_o2 <= n1237_i2;
    n1238_o2 <= n1238_i2;
    G374_o2 <= G374_i2;
    G376_o2 <= G376_i2;
    G370_o2 <= G370_i2;
    G372_o2 <= G372_i2;
    G373_o2 <= G373_i2;
    G377_o2 <= G377_i2;
    G371_o2 <= G371_i2;
    G375_o2 <= G375_i2;
    G354_o2 <= G354_i2;
    G356_o2 <= G356_i2;
    G350_o2 <= G350_i2;
    G352_o2 <= G352_i2;
    G353_o2 <= G353_i2;
    G357_o2 <= G357_i2;
    G351_o2 <= G351_i2;
    G355_o2 <= G355_i2;
    G386_o2 <= G386_i2;
    G391_o2 <= G391_i2;
    n283_lo_buf_o2 <= n283_lo_buf_i2;
    n295_lo_buf_o2 <= n295_lo_buf_i2;
    n307_lo_buf_o2 <= n307_lo_buf_i2;
    n319_lo_buf_o2 <= n319_lo_buf_i2;
    n331_lo_buf_o2 <= n331_lo_buf_i2;
    n343_lo_buf_o2 <= n343_lo_buf_i2;
    n355_lo_buf_o2 <= n355_lo_buf_i2;
    n367_lo_buf_o2 <= n367_lo_buf_i2;
    n379_lo_buf_o2 <= n379_lo_buf_i2;
    n391_lo_buf_o2 <= n391_lo_buf_i2;
    n403_lo_buf_o2 <= n403_lo_buf_i2;
    n415_lo_buf_o2 <= n415_lo_buf_i2;
    n427_lo_buf_o2 <= n427_lo_buf_i2;
    n439_lo_buf_o2 <= n439_lo_buf_i2;
    n451_lo_buf_o2 <= n451_lo_buf_i2;
    n463_lo_buf_o2 <= n463_lo_buf_i2;
    n475_lo_buf_o2 <= n475_lo_buf_i2;
    n487_lo_buf_o2 <= n487_lo_buf_i2;
    n499_lo_buf_o2 <= n499_lo_buf_i2;
    n511_lo_buf_o2 <= n511_lo_buf_i2;
    n523_lo_buf_o2 <= n523_lo_buf_i2;
    n535_lo_buf_o2 <= n535_lo_buf_i2;
    n547_lo_buf_o2 <= n547_lo_buf_i2;
    n559_lo_buf_o2 <= n559_lo_buf_i2;
    n571_lo_buf_o2 <= n571_lo_buf_i2;
    n583_lo_buf_o2 <= n583_lo_buf_i2;
    n595_lo_buf_o2 <= n595_lo_buf_i2;
    n607_lo_buf_o2 <= n607_lo_buf_i2;
    n619_lo_buf_o2 <= n619_lo_buf_i2;
    n631_lo_buf_o2 <= n631_lo_buf_i2;
    n643_lo_buf_o2 <= n643_lo_buf_i2;
    n655_lo_buf_o2 <= n655_lo_buf_i2;
    G234_o2 <= G234_i2;
    G247_o2 <= G247_i2;
    G260_o2 <= G260_i2;
    G273_o2 <= G273_i2;
    G286_o2 <= G286_i2;
    G299_o2 <= G299_i2;
    G312_o2 <= G312_i2;
    G325_o2 <= G325_i2;
    n667_lo_buf_o2 <= n667_lo_buf_i2;
    n679_lo_buf_o2 <= n679_lo_buf_i2;
    n691_lo_buf_o2 <= n691_lo_buf_i2;
    n703_lo_buf_o2 <= n703_lo_buf_i2;
    n715_lo_buf_o2 <= n715_lo_buf_i2;
    n727_lo_buf_o2 <= n727_lo_buf_i2;
    n739_lo_buf_o2 <= n739_lo_buf_i2;
    n751_lo_buf_o2 <= n751_lo_buf_i2;
    n763_lo_buf_o2 <= n763_lo_buf_i2;
    G186_o2 <= G186_i2;
    G189_o2 <= G189_i2;
    G192_o2 <= G192_i2;
    G195_o2 <= G195_i2;
    G198_o2 <= G198_i2;
    G201_o2 <= G201_i2;
    G204_o2 <= G204_i2;
    G207_o2 <= G207_i2;
    n280_lo_buf_o2 <= n280_lo_buf_i2;
    n292_lo_buf_o2 <= n292_lo_buf_i2;
    n304_lo_buf_o2 <= n304_lo_buf_i2;
    n316_lo_buf_o2 <= n316_lo_buf_i2;
    n328_lo_buf_o2 <= n328_lo_buf_i2;
    n340_lo_buf_o2 <= n340_lo_buf_i2;
    n352_lo_buf_o2 <= n352_lo_buf_i2;
    n364_lo_buf_o2 <= n364_lo_buf_i2;
    n376_lo_buf_o2 <= n376_lo_buf_i2;
    n388_lo_buf_o2 <= n388_lo_buf_i2;
    n400_lo_buf_o2 <= n400_lo_buf_i2;
    n412_lo_buf_o2 <= n412_lo_buf_i2;
    n424_lo_buf_o2 <= n424_lo_buf_i2;
    n436_lo_buf_o2 <= n436_lo_buf_i2;
    n448_lo_buf_o2 <= n448_lo_buf_i2;
    n460_lo_buf_o2 <= n460_lo_buf_i2;
    n472_lo_buf_o2 <= n472_lo_buf_i2;
    n484_lo_buf_o2 <= n484_lo_buf_i2;
    n496_lo_buf_o2 <= n496_lo_buf_i2;
    n508_lo_buf_o2 <= n508_lo_buf_i2;
    n520_lo_buf_o2 <= n520_lo_buf_i2;
    n532_lo_buf_o2 <= n532_lo_buf_i2;
    n544_lo_buf_o2 <= n544_lo_buf_i2;
    n556_lo_buf_o2 <= n556_lo_buf_i2;
    n568_lo_buf_o2 <= n568_lo_buf_i2;
    n580_lo_buf_o2 <= n580_lo_buf_i2;
    n592_lo_buf_o2 <= n592_lo_buf_i2;
    n604_lo_buf_o2 <= n604_lo_buf_i2;
    n616_lo_buf_o2 <= n616_lo_buf_i2;
    n628_lo_buf_o2 <= n628_lo_buf_i2;
    n640_lo_buf_o2 <= n640_lo_buf_i2;
    n652_lo_buf_o2 <= n652_lo_buf_i2;
  end
  initial begin
    n286_lo <= 1'b0;
    n298_lo <= 1'b0;
    n310_lo <= 1'b0;
    n322_lo <= 1'b0;
    n334_lo <= 1'b0;
    n346_lo <= 1'b0;
    n358_lo <= 1'b0;
    n370_lo <= 1'b0;
    n382_lo <= 1'b0;
    n394_lo <= 1'b0;
    n406_lo <= 1'b0;
    n418_lo <= 1'b0;
    n430_lo <= 1'b0;
    n442_lo <= 1'b0;
    n454_lo <= 1'b0;
    n466_lo <= 1'b0;
    n478_lo <= 1'b0;
    n490_lo <= 1'b0;
    n502_lo <= 1'b0;
    n514_lo <= 1'b0;
    n526_lo <= 1'b0;
    n538_lo <= 1'b0;
    n550_lo <= 1'b0;
    n562_lo <= 1'b0;
    n574_lo <= 1'b0;
    n586_lo <= 1'b0;
    n598_lo <= 1'b0;
    n610_lo <= 1'b0;
    n622_lo <= 1'b0;
    n634_lo <= 1'b0;
    n646_lo <= 1'b0;
    n658_lo <= 1'b0;
    n661_lo <= 1'b0;
    n673_lo <= 1'b0;
    n685_lo <= 1'b0;
    n697_lo <= 1'b0;
    n709_lo <= 1'b0;
    n721_lo <= 1'b0;
    n733_lo <= 1'b0;
    n745_lo <= 1'b0;
    n757_lo <= 1'b0;
    n1248_o2 <= 1'b0;
    n1249_o2 <= 1'b0;
    n1250_o2 <= 1'b0;
    n1251_o2 <= 1'b0;
    n1252_o2 <= 1'b0;
    n1253_o2 <= 1'b0;
    n1254_o2 <= 1'b0;
    n1255_o2 <= 1'b0;
    n1207_o2 <= 1'b0;
    n1208_o2 <= 1'b0;
    n1209_o2 <= 1'b0;
    n1210_o2 <= 1'b0;
    n1211_o2 <= 1'b0;
    n1212_o2 <= 1'b0;
    n1213_o2 <= 1'b0;
    n1214_o2 <= 1'b0;
    n1215_o2 <= 1'b0;
    n1216_o2 <= 1'b0;
    n1217_o2 <= 1'b0;
    n1218_o2 <= 1'b0;
    n1219_o2 <= 1'b0;
    n1220_o2 <= 1'b0;
    n1221_o2 <= 1'b0;
    n1222_o2 <= 1'b0;
    n1223_o2 <= 1'b0;
    n1224_o2 <= 1'b0;
    n1225_o2 <= 1'b0;
    n1226_o2 <= 1'b0;
    n1227_o2 <= 1'b0;
    n1228_o2 <= 1'b0;
    n1229_o2 <= 1'b0;
    n1230_o2 <= 1'b0;
    n1231_o2 <= 1'b0;
    n1232_o2 <= 1'b0;
    n1233_o2 <= 1'b0;
    n1234_o2 <= 1'b0;
    n1235_o2 <= 1'b0;
    n1236_o2 <= 1'b0;
    n1237_o2 <= 1'b0;
    n1238_o2 <= 1'b0;
    G374_o2 <= 1'b0;
    G376_o2 <= 1'b0;
    G370_o2 <= 1'b0;
    G372_o2 <= 1'b0;
    G373_o2 <= 1'b0;
    G377_o2 <= 1'b0;
    G371_o2 <= 1'b0;
    G375_o2 <= 1'b0;
    G354_o2 <= 1'b0;
    G356_o2 <= 1'b0;
    G350_o2 <= 1'b0;
    G352_o2 <= 1'b0;
    G353_o2 <= 1'b0;
    G357_o2 <= 1'b0;
    G351_o2 <= 1'b0;
    G355_o2 <= 1'b0;
    G386_o2 <= 1'b0;
    G391_o2 <= 1'b0;
    n283_lo_buf_o2 <= 1'b0;
    n295_lo_buf_o2 <= 1'b0;
    n307_lo_buf_o2 <= 1'b0;
    n319_lo_buf_o2 <= 1'b0;
    n331_lo_buf_o2 <= 1'b0;
    n343_lo_buf_o2 <= 1'b0;
    n355_lo_buf_o2 <= 1'b0;
    n367_lo_buf_o2 <= 1'b0;
    n379_lo_buf_o2 <= 1'b0;
    n391_lo_buf_o2 <= 1'b0;
    n403_lo_buf_o2 <= 1'b0;
    n415_lo_buf_o2 <= 1'b0;
    n427_lo_buf_o2 <= 1'b0;
    n439_lo_buf_o2 <= 1'b0;
    n451_lo_buf_o2 <= 1'b0;
    n463_lo_buf_o2 <= 1'b0;
    n475_lo_buf_o2 <= 1'b0;
    n487_lo_buf_o2 <= 1'b0;
    n499_lo_buf_o2 <= 1'b0;
    n511_lo_buf_o2 <= 1'b0;
    n523_lo_buf_o2 <= 1'b0;
    n535_lo_buf_o2 <= 1'b0;
    n547_lo_buf_o2 <= 1'b0;
    n559_lo_buf_o2 <= 1'b0;
    n571_lo_buf_o2 <= 1'b0;
    n583_lo_buf_o2 <= 1'b0;
    n595_lo_buf_o2 <= 1'b0;
    n607_lo_buf_o2 <= 1'b0;
    n619_lo_buf_o2 <= 1'b0;
    n631_lo_buf_o2 <= 1'b0;
    n643_lo_buf_o2 <= 1'b0;
    n655_lo_buf_o2 <= 1'b0;
    G234_o2 <= 1'b0;
    G247_o2 <= 1'b0;
    G260_o2 <= 1'b0;
    G273_o2 <= 1'b0;
    G286_o2 <= 1'b0;
    G299_o2 <= 1'b0;
    G312_o2 <= 1'b0;
    G325_o2 <= 1'b0;
    n667_lo_buf_o2 <= 1'b0;
    n679_lo_buf_o2 <= 1'b0;
    n691_lo_buf_o2 <= 1'b0;
    n703_lo_buf_o2 <= 1'b0;
    n715_lo_buf_o2 <= 1'b0;
    n727_lo_buf_o2 <= 1'b0;
    n739_lo_buf_o2 <= 1'b0;
    n751_lo_buf_o2 <= 1'b0;
    n763_lo_buf_o2 <= 1'b0;
    G186_o2 <= 1'b0;
    G189_o2 <= 1'b0;
    G192_o2 <= 1'b0;
    G195_o2 <= 1'b0;
    G198_o2 <= 1'b0;
    G201_o2 <= 1'b0;
    G204_o2 <= 1'b0;
    G207_o2 <= 1'b0;
    n280_lo_buf_o2 <= 1'b0;
    n292_lo_buf_o2 <= 1'b0;
    n304_lo_buf_o2 <= 1'b0;
    n316_lo_buf_o2 <= 1'b0;
    n328_lo_buf_o2 <= 1'b0;
    n340_lo_buf_o2 <= 1'b0;
    n352_lo_buf_o2 <= 1'b0;
    n364_lo_buf_o2 <= 1'b0;
    n376_lo_buf_o2 <= 1'b0;
    n388_lo_buf_o2 <= 1'b0;
    n400_lo_buf_o2 <= 1'b0;
    n412_lo_buf_o2 <= 1'b0;
    n424_lo_buf_o2 <= 1'b0;
    n436_lo_buf_o2 <= 1'b0;
    n448_lo_buf_o2 <= 1'b0;
    n460_lo_buf_o2 <= 1'b0;
    n472_lo_buf_o2 <= 1'b0;
    n484_lo_buf_o2 <= 1'b0;
    n496_lo_buf_o2 <= 1'b0;
    n508_lo_buf_o2 <= 1'b0;
    n520_lo_buf_o2 <= 1'b0;
    n532_lo_buf_o2 <= 1'b0;
    n544_lo_buf_o2 <= 1'b0;
    n556_lo_buf_o2 <= 1'b0;
    n568_lo_buf_o2 <= 1'b0;
    n580_lo_buf_o2 <= 1'b0;
    n592_lo_buf_o2 <= 1'b0;
    n604_lo_buf_o2 <= 1'b0;
    n616_lo_buf_o2 <= 1'b0;
    n628_lo_buf_o2 <= 1'b0;
    n640_lo_buf_o2 <= 1'b0;
    n652_lo_buf_o2 <= 1'b0;
  end
endmodule


