// Benchmark "c499" written by ABC on Sun Oct 29 19:31:47 2023

module c499 (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41,
    G468, G469, G470, G471, G472, G473, G474, G475, G476, G477, G478, G479,
    G480, G481, G482, G483, G484, G485, G486, G487, G488, G489, G490, G491,
    G492, G493, G494, G495, G496, G497, G498, G499  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41;
  output G468, G469, G470, G471, G472, G473, G474, G475, G476, G477, G478,
    G479, G480, G481, G482, G483, G484, G485, G486, G487, G488, G489, G490,
    G491, G492, G493, G494, G495, G496, G497, G498, G499;
  reg n277_lo, n280_lo, n283_lo, n286_lo, n289_lo, n292_lo, n295_lo,
    n298_lo, n301_lo, n304_lo, n307_lo, n310_lo, n313_lo, n316_lo, n319_lo,
    n322_lo, n325_lo, n328_lo, n331_lo, n334_lo, n337_lo, n340_lo, n343_lo,
    n346_lo, n349_lo, n352_lo, n355_lo, n358_lo, n361_lo, n364_lo, n367_lo,
    n370_lo, n373_lo, n376_lo, n379_lo, n382_lo, n385_lo, n388_lo, n391_lo,
    n394_lo, n397_lo, n400_lo, n403_lo, n406_lo, n409_lo, n412_lo, n415_lo,
    n418_lo, n421_lo, n424_lo, n427_lo, n430_lo, n433_lo, n436_lo, n439_lo,
    n442_lo, n445_lo, n448_lo, n451_lo, n454_lo, n457_lo, n460_lo, n463_lo,
    n466_lo, n469_lo, n472_lo, n475_lo, n478_lo, n481_lo, n484_lo, n487_lo,
    n490_lo, n493_lo, n496_lo, n499_lo, n502_lo, n505_lo, n508_lo, n511_lo,
    n514_lo, n517_lo, n520_lo, n523_lo, n526_lo, n529_lo, n532_lo, n535_lo,
    n538_lo, n541_lo, n544_lo, n547_lo, n550_lo, n553_lo, n556_lo, n559_lo,
    n562_lo, n565_lo, n568_lo, n571_lo, n574_lo, n577_lo, n580_lo, n583_lo,
    n586_lo, n589_lo, n592_lo, n595_lo, n598_lo, n601_lo, n604_lo, n607_lo,
    n610_lo, n613_lo, n616_lo, n619_lo, n622_lo, n625_lo, n628_lo, n631_lo,
    n634_lo, n637_lo, n640_lo, n643_lo, n646_lo, n649_lo, n652_lo, n655_lo,
    n658_lo, n661_lo, n664_lo, n667_lo, n670_lo, n673_lo, n676_lo, n679_lo,
    n682_lo, n685_lo, n688_lo, n691_lo, n694_lo, n697_lo, n700_lo, n703_lo,
    n706_lo, n709_lo, n712_lo, n715_lo, n718_lo, n721_lo, n724_lo, n727_lo,
    n730_lo, n733_lo, n736_lo, n739_lo, n742_lo, n745_lo, n748_lo, n751_lo,
    n754_lo, n757_lo, n760_lo, n763_lo, n766_lo;
  wire new_G146_, new_G147_, new_G148_, new_G149_, new_G150_, new_G151_,
    new_G152_, new_G153_, new_G154_, new_G155_, new_G156_, new_G157_,
    new_G158_, new_G159_, new_G160_, new_G161_, new_G162_, new_G163_,
    new_G164_, new_G165_, new_G166_, new_G167_, new_G168_, new_G169_,
    new_G170_, new_G171_, new_G172_, new_G173_, new_G174_, new_G175_,
    new_G176_, new_G177_, new_G178_, new_G179_, new_G180_, new_G181_,
    new_G182_, new_G183_, new_G184_, new_G185_, new_G186_, new_G189_,
    new_G192_, new_G195_, new_G198_, new_G201_, new_G204_, new_G207_,
    new_G210_, new_G211_, new_G212_, new_G213_, new_G214_, new_G215_,
    new_G216_, new_G217_, new_G218_, new_G219_, new_G220_, new_G221_,
    new_G222_, new_G223_, new_G224_, new_G225_, new_G226_, new_G227_,
    new_G228_, new_G229_, new_G230_, new_G231_, new_G232_, new_G233_,
    new_G234_, new_G247_, new_G260_, new_G273_, new_G286_, new_G299_,
    new_G312_, new_G325_, new_G338_, new_G339_, new_G340_, new_G341_,
    new_G342_, new_G343_, new_G344_, new_G345_, new_G346_, new_G347_,
    new_G348_, new_G349_, new_G350_, new_G351_, new_G352_, new_G353_,
    new_G354_, new_G355_, new_G356_, new_G357_, new_G358_, new_G359_,
    new_G360_, new_G361_, new_G362_, new_G363_, new_G364_, new_G365_,
    new_G366_, new_G367_, new_G368_, new_G369_, new_G370_, new_G371_,
    new_G372_, new_G373_, new_G374_, new_G375_, new_G376_, new_G377_,
    new_G378_, new_G379_, new_G380_, new_G381_, new_G382_, new_G383_,
    new_G384_, new_G385_, new_G386_, new_G391_, new_G396_, new_G401_,
    new_G406_, new_G411_, new_G416_, new_G421_, new_G426_, new_G431_,
    new_G436_, new_G437_, new_G438_, new_G439_, new_G440_, new_G441_,
    new_G442_, new_G443_, new_G444_, new_G445_, new_G446_, new_G447_,
    new_G448_, new_G449_, new_G450_, new_G451_, new_G452_, new_G453_,
    new_G454_, new_G455_, new_G456_, new_G457_, new_G458_, new_G459_,
    new_G460_, new_G461_, new_G462_, new_G463_, new_G464_, new_G465_,
    new_G466_, new_G467_, n277_li, n280_li, n283_li, n286_li, n289_li,
    n292_li, n295_li, n298_li, n301_li, n304_li, n307_li, n310_li, n313_li,
    n316_li, n319_li, n322_li, n325_li, n328_li, n331_li, n334_li, n337_li,
    n340_li, n343_li, n346_li, n349_li, n352_li, n355_li, n358_li, n361_li,
    n364_li, n367_li, n370_li, n373_li, n376_li, n379_li, n382_li, n385_li,
    n388_li, n391_li, n394_li, n397_li, n400_li, n403_li, n406_li, n409_li,
    n412_li, n415_li, n418_li, n421_li, n424_li, n427_li, n430_li, n433_li,
    n436_li, n439_li, n442_li, n445_li, n448_li, n451_li, n454_li, n457_li,
    n460_li, n463_li, n466_li, n469_li, n472_li, n475_li, n478_li, n481_li,
    n484_li, n487_li, n490_li, n493_li, n496_li, n499_li, n502_li, n505_li,
    n508_li, n511_li, n514_li, n517_li, n520_li, n523_li, n526_li, n529_li,
    n532_li, n535_li, n538_li, n541_li, n544_li, n547_li, n550_li, n553_li,
    n556_li, n559_li, n562_li, n565_li, n568_li, n571_li, n574_li, n577_li,
    n580_li, n583_li, n586_li, n589_li, n592_li, n595_li, n598_li, n601_li,
    n604_li, n607_li, n610_li, n613_li, n616_li, n619_li, n622_li, n625_li,
    n628_li, n631_li, n634_li, n637_li, n640_li, n643_li, n646_li, n649_li,
    n652_li, n655_li, n658_li, n661_li, n664_li, n667_li, n670_li, n673_li,
    n676_li, n679_li, n682_li, n685_li, n688_li, n691_li, n694_li, n697_li,
    n700_li, n703_li, n706_li, n709_li, n712_li, n715_li, n718_li, n721_li,
    n724_li, n727_li, n730_li, n733_li, n736_li, n739_li, n742_li, n745_li,
    n748_li, n751_li, n754_li, n757_li, n760_li, n763_li, n766_li;
  assign new_G146_ = n286_lo ^ n298_lo;
  assign new_G147_ = n310_lo ^ n322_lo;
  assign new_G148_ = n334_lo ^ n346_lo;
  assign new_G149_ = n358_lo ^ n370_lo;
  assign new_G150_ = n382_lo ^ n394_lo;
  assign new_G151_ = n406_lo ^ n418_lo;
  assign new_G152_ = n430_lo ^ n442_lo;
  assign new_G153_ = n454_lo ^ n466_lo;
  assign new_G154_ = n478_lo ^ n490_lo;
  assign new_G155_ = n502_lo ^ n514_lo;
  assign new_G156_ = n526_lo ^ n538_lo;
  assign new_G157_ = n550_lo ^ n562_lo;
  assign new_G158_ = n574_lo ^ n586_lo;
  assign new_G159_ = n598_lo ^ n610_lo;
  assign new_G160_ = n622_lo ^ n634_lo;
  assign new_G161_ = n646_lo ^ n658_lo;
  assign new_G162_ = n670_lo & n766_lo;
  assign new_G163_ = n682_lo & n766_lo;
  assign new_G164_ = n694_lo & n766_lo;
  assign new_G165_ = n706_lo & n766_lo;
  assign new_G166_ = n718_lo & n766_lo;
  assign new_G167_ = n730_lo & n766_lo;
  assign new_G168_ = n742_lo & n766_lo;
  assign new_G169_ = n754_lo & n766_lo;
  assign new_G170_ = n286_lo ^ n334_lo;
  assign new_G171_ = n382_lo ^ n430_lo;
  assign new_G172_ = n298_lo ^ n346_lo;
  assign new_G173_ = n394_lo ^ n442_lo;
  assign new_G174_ = n310_lo ^ n358_lo;
  assign new_G175_ = n406_lo ^ n454_lo;
  assign new_G176_ = n322_lo ^ n370_lo;
  assign new_G177_ = n418_lo ^ n466_lo;
  assign new_G178_ = n478_lo ^ n526_lo;
  assign new_G179_ = n574_lo ^ n622_lo;
  assign new_G180_ = n490_lo ^ n538_lo;
  assign new_G181_ = n586_lo ^ n634_lo;
  assign new_G182_ = n502_lo ^ n550_lo;
  assign new_G183_ = n598_lo ^ n646_lo;
  assign new_G184_ = n514_lo ^ n562_lo;
  assign new_G185_ = n610_lo ^ n658_lo;
  assign new_G186_ = new_G146_ ^ new_G147_;
  assign new_G189_ = new_G148_ ^ new_G149_;
  assign new_G192_ = new_G150_ ^ new_G151_;
  assign new_G195_ = new_G152_ ^ new_G153_;
  assign new_G198_ = new_G154_ ^ new_G155_;
  assign new_G201_ = new_G156_ ^ new_G157_;
  assign new_G204_ = new_G158_ ^ new_G159_;
  assign new_G207_ = new_G160_ ^ new_G161_;
  assign new_G210_ = new_G170_ ^ new_G171_;
  assign new_G211_ = new_G172_ ^ new_G173_;
  assign new_G212_ = new_G174_ ^ new_G175_;
  assign new_G213_ = new_G176_ ^ new_G177_;
  assign new_G214_ = new_G178_ ^ new_G179_;
  assign new_G215_ = new_G180_ ^ new_G181_;
  assign new_G216_ = new_G182_ ^ new_G183_;
  assign new_G217_ = new_G184_ ^ new_G185_;
  assign new_G218_ = new_G186_ ^ new_G189_;
  assign new_G219_ = new_G192_ ^ new_G195_;
  assign new_G220_ = new_G186_ ^ new_G192_;
  assign new_G221_ = new_G189_ ^ new_G195_;
  assign new_G222_ = new_G198_ ^ new_G201_;
  assign new_G223_ = new_G204_ ^ new_G207_;
  assign new_G224_ = new_G198_ ^ new_G204_;
  assign new_G225_ = new_G201_ ^ new_G207_;
  assign new_G226_ = new_G162_ ^ new_G222_;
  assign new_G227_ = new_G163_ ^ new_G223_;
  assign new_G228_ = new_G164_ ^ new_G224_;
  assign new_G229_ = new_G165_ ^ new_G225_;
  assign new_G230_ = new_G166_ ^ new_G218_;
  assign new_G231_ = new_G167_ ^ new_G219_;
  assign new_G232_ = new_G168_ ^ new_G220_;
  assign new_G233_ = new_G169_ ^ new_G221_;
  assign new_G234_ = new_G210_ ^ new_G226_;
  assign new_G247_ = new_G211_ ^ new_G227_;
  assign new_G260_ = new_G212_ ^ new_G228_;
  assign new_G273_ = new_G213_ ^ new_G229_;
  assign new_G286_ = new_G214_ ^ new_G230_;
  assign new_G299_ = new_G215_ ^ new_G231_;
  assign new_G312_ = new_G216_ ^ new_G232_;
  assign new_G325_ = new_G217_ ^ new_G233_;
  assign new_G338_ = ~new_G234_;
  assign new_G339_ = ~new_G247_;
  assign new_G340_ = ~new_G260_;
  assign new_G341_ = ~new_G234_;
  assign new_G342_ = ~new_G247_;
  assign new_G343_ = ~new_G273_;
  assign new_G344_ = ~new_G234_;
  assign new_G345_ = ~new_G260_;
  assign new_G346_ = ~new_G273_;
  assign new_G347_ = ~new_G247_;
  assign new_G348_ = ~new_G260_;
  assign new_G349_ = ~new_G273_;
  assign new_G350_ = ~new_G299_;
  assign new_G351_ = ~new_G325_;
  assign new_G352_ = ~new_G299_;
  assign new_G353_ = ~new_G312_;
  assign new_G354_ = ~new_G286_;
  assign new_G355_ = ~new_G325_;
  assign new_G356_ = ~new_G286_;
  assign new_G357_ = ~new_G312_;
  assign new_G358_ = ~new_G286_;
  assign new_G359_ = ~new_G299_;
  assign new_G360_ = ~new_G312_;
  assign new_G361_ = ~new_G286_;
  assign new_G362_ = ~new_G299_;
  assign new_G363_ = ~new_G325_;
  assign new_G364_ = ~new_G286_;
  assign new_G365_ = ~new_G312_;
  assign new_G366_ = ~new_G325_;
  assign new_G367_ = ~new_G299_;
  assign new_G368_ = ~new_G312_;
  assign new_G369_ = ~new_G325_;
  assign new_G370_ = ~new_G247_;
  assign new_G371_ = ~new_G273_;
  assign new_G372_ = ~new_G247_;
  assign new_G373_ = ~new_G260_;
  assign new_G374_ = ~new_G234_;
  assign new_G375_ = ~new_G273_;
  assign new_G376_ = ~new_G234_;
  assign new_G377_ = ~new_G260_;
  assign new_G378_ = new_G273_ & new_G338_ & new_G339_ & new_G340_;
  assign new_G379_ = new_G343_ & new_G341_ & new_G342_ & new_G260_;
  assign new_G380_ = new_G346_ & new_G344_ & new_G247_ & new_G345_;
  assign new_G381_ = new_G349_ & new_G234_ & new_G347_ & new_G348_;
  assign new_G382_ = new_G325_ & new_G358_ & new_G359_ & new_G360_;
  assign new_G383_ = new_G363_ & new_G361_ & new_G362_ & new_G312_;
  assign new_G384_ = new_G366_ & new_G364_ & new_G299_ & new_G365_;
  assign new_G385_ = new_G369_ & new_G286_ & new_G367_ & new_G368_;
  assign new_G386_ = new_G381_ | new_G380_ | new_G378_ | new_G379_;
  assign new_G391_ = new_G385_ | new_G384_ | new_G382_ | new_G383_;
  assign new_G396_ = new_G351_ & new_G286_ & new_G350_ & new_G312_ & new_G386_;
  assign new_G401_ = new_G325_ & new_G286_ & new_G352_ & new_G353_ & new_G386_;
  assign new_G406_ = new_G355_ & new_G354_ & new_G299_ & new_G312_ & new_G386_;
  assign new_G411_ = new_G325_ & new_G356_ & new_G299_ & new_G357_ & new_G386_;
  assign new_G416_ = new_G371_ & new_G234_ & new_G370_ & new_G260_ & new_G391_;
  assign new_G421_ = new_G273_ & new_G234_ & new_G372_ & new_G373_ & new_G391_;
  assign new_G426_ = new_G375_ & new_G374_ & new_G247_ & new_G260_ & new_G391_;
  assign new_G431_ = new_G273_ & new_G376_ & new_G247_ & new_G377_ & new_G391_;
  assign new_G436_ = new_G234_ & new_G396_;
  assign new_G437_ = new_G247_ & new_G396_;
  assign new_G438_ = new_G260_ & new_G396_;
  assign new_G439_ = new_G273_ & new_G396_;
  assign new_G440_ = new_G234_ & new_G401_;
  assign new_G441_ = new_G247_ & new_G401_;
  assign new_G442_ = new_G260_ & new_G401_;
  assign new_G443_ = new_G273_ & new_G401_;
  assign new_G444_ = new_G234_ & new_G406_;
  assign new_G445_ = new_G247_ & new_G406_;
  assign new_G446_ = new_G260_ & new_G406_;
  assign new_G447_ = new_G273_ & new_G406_;
  assign new_G448_ = new_G234_ & new_G411_;
  assign new_G449_ = new_G247_ & new_G411_;
  assign new_G450_ = new_G260_ & new_G411_;
  assign new_G451_ = new_G273_ & new_G411_;
  assign new_G452_ = new_G286_ & new_G416_;
  assign new_G453_ = new_G299_ & new_G416_;
  assign new_G454_ = new_G312_ & new_G416_;
  assign new_G455_ = new_G325_ & new_G416_;
  assign new_G456_ = new_G286_ & new_G421_;
  assign new_G457_ = new_G299_ & new_G421_;
  assign new_G458_ = new_G312_ & new_G421_;
  assign new_G459_ = new_G325_ & new_G421_;
  assign new_G460_ = new_G286_ & new_G426_;
  assign new_G461_ = new_G299_ & new_G426_;
  assign new_G462_ = new_G312_ & new_G426_;
  assign new_G463_ = new_G325_ & new_G426_;
  assign new_G464_ = new_G286_ & new_G431_;
  assign new_G465_ = new_G299_ & new_G431_;
  assign new_G466_ = new_G312_ & new_G431_;
  assign new_G467_ = new_G325_ & new_G431_;
  assign G468 = n286_lo ^ new_G436_;
  assign G469 = n298_lo ^ new_G437_;
  assign G470 = n310_lo ^ new_G438_;
  assign G471 = n322_lo ^ new_G439_;
  assign G472 = n334_lo ^ new_G440_;
  assign G473 = n346_lo ^ new_G441_;
  assign G474 = n358_lo ^ new_G442_;
  assign G475 = n370_lo ^ new_G443_;
  assign G476 = n382_lo ^ new_G444_;
  assign G477 = n394_lo ^ new_G445_;
  assign G478 = n406_lo ^ new_G446_;
  assign G479 = n418_lo ^ new_G447_;
  assign G480 = n430_lo ^ new_G448_;
  assign G481 = n442_lo ^ new_G449_;
  assign G482 = n454_lo ^ new_G450_;
  assign G483 = n466_lo ^ new_G451_;
  assign G484 = n478_lo ^ new_G452_;
  assign G485 = n490_lo ^ new_G453_;
  assign G486 = n502_lo ^ new_G454_;
  assign G487 = n514_lo ^ new_G455_;
  assign G488 = n526_lo ^ new_G456_;
  assign G489 = n538_lo ^ new_G457_;
  assign G490 = n550_lo ^ new_G458_;
  assign G491 = n562_lo ^ new_G459_;
  assign G492 = n574_lo ^ new_G460_;
  assign G493 = n586_lo ^ new_G461_;
  assign G494 = n598_lo ^ new_G462_;
  assign G495 = n610_lo ^ new_G463_;
  assign G496 = n622_lo ^ new_G464_;
  assign G497 = n634_lo ^ new_G465_;
  assign G498 = n646_lo ^ new_G466_;
  assign G499 = n658_lo ^ new_G467_;
  assign n277_li = G1;
  assign n280_li = n277_lo;
  assign n283_li = n280_lo;
  assign n286_li = n283_lo;
  assign n289_li = G2;
  assign n292_li = n289_lo;
  assign n295_li = n292_lo;
  assign n298_li = n295_lo;
  assign n301_li = G3;
  assign n304_li = n301_lo;
  assign n307_li = n304_lo;
  assign n310_li = n307_lo;
  assign n313_li = G4;
  assign n316_li = n313_lo;
  assign n319_li = n316_lo;
  assign n322_li = n319_lo;
  assign n325_li = G5;
  assign n328_li = n325_lo;
  assign n331_li = n328_lo;
  assign n334_li = n331_lo;
  assign n337_li = G6;
  assign n340_li = n337_lo;
  assign n343_li = n340_lo;
  assign n346_li = n343_lo;
  assign n349_li = G7;
  assign n352_li = n349_lo;
  assign n355_li = n352_lo;
  assign n358_li = n355_lo;
  assign n361_li = G8;
  assign n364_li = n361_lo;
  assign n367_li = n364_lo;
  assign n370_li = n367_lo;
  assign n373_li = G9;
  assign n376_li = n373_lo;
  assign n379_li = n376_lo;
  assign n382_li = n379_lo;
  assign n385_li = G10;
  assign n388_li = n385_lo;
  assign n391_li = n388_lo;
  assign n394_li = n391_lo;
  assign n397_li = G11;
  assign n400_li = n397_lo;
  assign n403_li = n400_lo;
  assign n406_li = n403_lo;
  assign n409_li = G12;
  assign n412_li = n409_lo;
  assign n415_li = n412_lo;
  assign n418_li = n415_lo;
  assign n421_li = G13;
  assign n424_li = n421_lo;
  assign n427_li = n424_lo;
  assign n430_li = n427_lo;
  assign n433_li = G14;
  assign n436_li = n433_lo;
  assign n439_li = n436_lo;
  assign n442_li = n439_lo;
  assign n445_li = G15;
  assign n448_li = n445_lo;
  assign n451_li = n448_lo;
  assign n454_li = n451_lo;
  assign n457_li = G16;
  assign n460_li = n457_lo;
  assign n463_li = n460_lo;
  assign n466_li = n463_lo;
  assign n469_li = G17;
  assign n472_li = n469_lo;
  assign n475_li = n472_lo;
  assign n478_li = n475_lo;
  assign n481_li = G18;
  assign n484_li = n481_lo;
  assign n487_li = n484_lo;
  assign n490_li = n487_lo;
  assign n493_li = G19;
  assign n496_li = n493_lo;
  assign n499_li = n496_lo;
  assign n502_li = n499_lo;
  assign n505_li = G20;
  assign n508_li = n505_lo;
  assign n511_li = n508_lo;
  assign n514_li = n511_lo;
  assign n517_li = G21;
  assign n520_li = n517_lo;
  assign n523_li = n520_lo;
  assign n526_li = n523_lo;
  assign n529_li = G22;
  assign n532_li = n529_lo;
  assign n535_li = n532_lo;
  assign n538_li = n535_lo;
  assign n541_li = G23;
  assign n544_li = n541_lo;
  assign n547_li = n544_lo;
  assign n550_li = n547_lo;
  assign n553_li = G24;
  assign n556_li = n553_lo;
  assign n559_li = n556_lo;
  assign n562_li = n559_lo;
  assign n565_li = G25;
  assign n568_li = n565_lo;
  assign n571_li = n568_lo;
  assign n574_li = n571_lo;
  assign n577_li = G26;
  assign n580_li = n577_lo;
  assign n583_li = n580_lo;
  assign n586_li = n583_lo;
  assign n589_li = G27;
  assign n592_li = n589_lo;
  assign n595_li = n592_lo;
  assign n598_li = n595_lo;
  assign n601_li = G28;
  assign n604_li = n601_lo;
  assign n607_li = n604_lo;
  assign n610_li = n607_lo;
  assign n613_li = G29;
  assign n616_li = n613_lo;
  assign n619_li = n616_lo;
  assign n622_li = n619_lo;
  assign n625_li = G30;
  assign n628_li = n625_lo;
  assign n631_li = n628_lo;
  assign n634_li = n631_lo;
  assign n637_li = G31;
  assign n640_li = n637_lo;
  assign n643_li = n640_lo;
  assign n646_li = n643_lo;
  assign n649_li = G32;
  assign n652_li = n649_lo;
  assign n655_li = n652_lo;
  assign n658_li = n655_lo;
  assign n661_li = G33;
  assign n664_li = n661_lo;
  assign n667_li = n664_lo;
  assign n670_li = n667_lo;
  assign n673_li = G34;
  assign n676_li = n673_lo;
  assign n679_li = n676_lo;
  assign n682_li = n679_lo;
  assign n685_li = G35;
  assign n688_li = n685_lo;
  assign n691_li = n688_lo;
  assign n694_li = n691_lo;
  assign n697_li = G36;
  assign n700_li = n697_lo;
  assign n703_li = n700_lo;
  assign n706_li = n703_lo;
  assign n709_li = G37;
  assign n712_li = n709_lo;
  assign n715_li = n712_lo;
  assign n718_li = n715_lo;
  assign n721_li = G38;
  assign n724_li = n721_lo;
  assign n727_li = n724_lo;
  assign n730_li = n727_lo;
  assign n733_li = G39;
  assign n736_li = n733_lo;
  assign n739_li = n736_lo;
  assign n742_li = n739_lo;
  assign n745_li = G40;
  assign n748_li = n745_lo;
  assign n751_li = n748_lo;
  assign n754_li = n751_lo;
  assign n757_li = G41;
  assign n760_li = n757_lo;
  assign n763_li = n760_lo;
  assign n766_li = n763_lo;
  always @ (posedge clock) begin
    n277_lo <= n277_li;
    n280_lo <= n280_li;
    n283_lo <= n283_li;
    n286_lo <= n286_li;
    n289_lo <= n289_li;
    n292_lo <= n292_li;
    n295_lo <= n295_li;
    n298_lo <= n298_li;
    n301_lo <= n301_li;
    n304_lo <= n304_li;
    n307_lo <= n307_li;
    n310_lo <= n310_li;
    n313_lo <= n313_li;
    n316_lo <= n316_li;
    n319_lo <= n319_li;
    n322_lo <= n322_li;
    n325_lo <= n325_li;
    n328_lo <= n328_li;
    n331_lo <= n331_li;
    n334_lo <= n334_li;
    n337_lo <= n337_li;
    n340_lo <= n340_li;
    n343_lo <= n343_li;
    n346_lo <= n346_li;
    n349_lo <= n349_li;
    n352_lo <= n352_li;
    n355_lo <= n355_li;
    n358_lo <= n358_li;
    n361_lo <= n361_li;
    n364_lo <= n364_li;
    n367_lo <= n367_li;
    n370_lo <= n370_li;
    n373_lo <= n373_li;
    n376_lo <= n376_li;
    n379_lo <= n379_li;
    n382_lo <= n382_li;
    n385_lo <= n385_li;
    n388_lo <= n388_li;
    n391_lo <= n391_li;
    n394_lo <= n394_li;
    n397_lo <= n397_li;
    n400_lo <= n400_li;
    n403_lo <= n403_li;
    n406_lo <= n406_li;
    n409_lo <= n409_li;
    n412_lo <= n412_li;
    n415_lo <= n415_li;
    n418_lo <= n418_li;
    n421_lo <= n421_li;
    n424_lo <= n424_li;
    n427_lo <= n427_li;
    n430_lo <= n430_li;
    n433_lo <= n433_li;
    n436_lo <= n436_li;
    n439_lo <= n439_li;
    n442_lo <= n442_li;
    n445_lo <= n445_li;
    n448_lo <= n448_li;
    n451_lo <= n451_li;
    n454_lo <= n454_li;
    n457_lo <= n457_li;
    n460_lo <= n460_li;
    n463_lo <= n463_li;
    n466_lo <= n466_li;
    n469_lo <= n469_li;
    n472_lo <= n472_li;
    n475_lo <= n475_li;
    n478_lo <= n478_li;
    n481_lo <= n481_li;
    n484_lo <= n484_li;
    n487_lo <= n487_li;
    n490_lo <= n490_li;
    n493_lo <= n493_li;
    n496_lo <= n496_li;
    n499_lo <= n499_li;
    n502_lo <= n502_li;
    n505_lo <= n505_li;
    n508_lo <= n508_li;
    n511_lo <= n511_li;
    n514_lo <= n514_li;
    n517_lo <= n517_li;
    n520_lo <= n520_li;
    n523_lo <= n523_li;
    n526_lo <= n526_li;
    n529_lo <= n529_li;
    n532_lo <= n532_li;
    n535_lo <= n535_li;
    n538_lo <= n538_li;
    n541_lo <= n541_li;
    n544_lo <= n544_li;
    n547_lo <= n547_li;
    n550_lo <= n550_li;
    n553_lo <= n553_li;
    n556_lo <= n556_li;
    n559_lo <= n559_li;
    n562_lo <= n562_li;
    n565_lo <= n565_li;
    n568_lo <= n568_li;
    n571_lo <= n571_li;
    n574_lo <= n574_li;
    n577_lo <= n577_li;
    n580_lo <= n580_li;
    n583_lo <= n583_li;
    n586_lo <= n586_li;
    n589_lo <= n589_li;
    n592_lo <= n592_li;
    n595_lo <= n595_li;
    n598_lo <= n598_li;
    n601_lo <= n601_li;
    n604_lo <= n604_li;
    n607_lo <= n607_li;
    n610_lo <= n610_li;
    n613_lo <= n613_li;
    n616_lo <= n616_li;
    n619_lo <= n619_li;
    n622_lo <= n622_li;
    n625_lo <= n625_li;
    n628_lo <= n628_li;
    n631_lo <= n631_li;
    n634_lo <= n634_li;
    n637_lo <= n637_li;
    n640_lo <= n640_li;
    n643_lo <= n643_li;
    n646_lo <= n646_li;
    n649_lo <= n649_li;
    n652_lo <= n652_li;
    n655_lo <= n655_li;
    n658_lo <= n658_li;
    n661_lo <= n661_li;
    n664_lo <= n664_li;
    n667_lo <= n667_li;
    n670_lo <= n670_li;
    n673_lo <= n673_li;
    n676_lo <= n676_li;
    n679_lo <= n679_li;
    n682_lo <= n682_li;
    n685_lo <= n685_li;
    n688_lo <= n688_li;
    n691_lo <= n691_li;
    n694_lo <= n694_li;
    n697_lo <= n697_li;
    n700_lo <= n700_li;
    n703_lo <= n703_li;
    n706_lo <= n706_li;
    n709_lo <= n709_li;
    n712_lo <= n712_li;
    n715_lo <= n715_li;
    n718_lo <= n718_li;
    n721_lo <= n721_li;
    n724_lo <= n724_li;
    n727_lo <= n727_li;
    n730_lo <= n730_li;
    n733_lo <= n733_li;
    n736_lo <= n736_li;
    n739_lo <= n739_li;
    n742_lo <= n742_li;
    n745_lo <= n745_li;
    n748_lo <= n748_li;
    n751_lo <= n751_li;
    n754_lo <= n754_li;
    n757_lo <= n757_li;
    n760_lo <= n760_li;
    n763_lo <= n763_li;
    n766_lo <= n766_li;
  end
  initial begin
    n277_lo <= 1'b0;
    n280_lo <= 1'b0;
    n283_lo <= 1'b0;
    n286_lo <= 1'b0;
    n289_lo <= 1'b0;
    n292_lo <= 1'b0;
    n295_lo <= 1'b0;
    n298_lo <= 1'b0;
    n301_lo <= 1'b0;
    n304_lo <= 1'b0;
    n307_lo <= 1'b0;
    n310_lo <= 1'b0;
    n313_lo <= 1'b0;
    n316_lo <= 1'b0;
    n319_lo <= 1'b0;
    n322_lo <= 1'b0;
    n325_lo <= 1'b0;
    n328_lo <= 1'b0;
    n331_lo <= 1'b0;
    n334_lo <= 1'b0;
    n337_lo <= 1'b0;
    n340_lo <= 1'b0;
    n343_lo <= 1'b0;
    n346_lo <= 1'b0;
    n349_lo <= 1'b0;
    n352_lo <= 1'b0;
    n355_lo <= 1'b0;
    n358_lo <= 1'b0;
    n361_lo <= 1'b0;
    n364_lo <= 1'b0;
    n367_lo <= 1'b0;
    n370_lo <= 1'b0;
    n373_lo <= 1'b0;
    n376_lo <= 1'b0;
    n379_lo <= 1'b0;
    n382_lo <= 1'b0;
    n385_lo <= 1'b0;
    n388_lo <= 1'b0;
    n391_lo <= 1'b0;
    n394_lo <= 1'b0;
    n397_lo <= 1'b0;
    n400_lo <= 1'b0;
    n403_lo <= 1'b0;
    n406_lo <= 1'b0;
    n409_lo <= 1'b0;
    n412_lo <= 1'b0;
    n415_lo <= 1'b0;
    n418_lo <= 1'b0;
    n421_lo <= 1'b0;
    n424_lo <= 1'b0;
    n427_lo <= 1'b0;
    n430_lo <= 1'b0;
    n433_lo <= 1'b0;
    n436_lo <= 1'b0;
    n439_lo <= 1'b0;
    n442_lo <= 1'b0;
    n445_lo <= 1'b0;
    n448_lo <= 1'b0;
    n451_lo <= 1'b0;
    n454_lo <= 1'b0;
    n457_lo <= 1'b0;
    n460_lo <= 1'b0;
    n463_lo <= 1'b0;
    n466_lo <= 1'b0;
    n469_lo <= 1'b0;
    n472_lo <= 1'b0;
    n475_lo <= 1'b0;
    n478_lo <= 1'b0;
    n481_lo <= 1'b0;
    n484_lo <= 1'b0;
    n487_lo <= 1'b0;
    n490_lo <= 1'b0;
    n493_lo <= 1'b0;
    n496_lo <= 1'b0;
    n499_lo <= 1'b0;
    n502_lo <= 1'b0;
    n505_lo <= 1'b0;
    n508_lo <= 1'b0;
    n511_lo <= 1'b0;
    n514_lo <= 1'b0;
    n517_lo <= 1'b0;
    n520_lo <= 1'b0;
    n523_lo <= 1'b0;
    n526_lo <= 1'b0;
    n529_lo <= 1'b0;
    n532_lo <= 1'b0;
    n535_lo <= 1'b0;
    n538_lo <= 1'b0;
    n541_lo <= 1'b0;
    n544_lo <= 1'b0;
    n547_lo <= 1'b0;
    n550_lo <= 1'b0;
    n553_lo <= 1'b0;
    n556_lo <= 1'b0;
    n559_lo <= 1'b0;
    n562_lo <= 1'b0;
    n565_lo <= 1'b0;
    n568_lo <= 1'b0;
    n571_lo <= 1'b0;
    n574_lo <= 1'b0;
    n577_lo <= 1'b0;
    n580_lo <= 1'b0;
    n583_lo <= 1'b0;
    n586_lo <= 1'b0;
    n589_lo <= 1'b0;
    n592_lo <= 1'b0;
    n595_lo <= 1'b0;
    n598_lo <= 1'b0;
    n601_lo <= 1'b0;
    n604_lo <= 1'b0;
    n607_lo <= 1'b0;
    n610_lo <= 1'b0;
    n613_lo <= 1'b0;
    n616_lo <= 1'b0;
    n619_lo <= 1'b0;
    n622_lo <= 1'b0;
    n625_lo <= 1'b0;
    n628_lo <= 1'b0;
    n631_lo <= 1'b0;
    n634_lo <= 1'b0;
    n637_lo <= 1'b0;
    n640_lo <= 1'b0;
    n643_lo <= 1'b0;
    n646_lo <= 1'b0;
    n649_lo <= 1'b0;
    n652_lo <= 1'b0;
    n655_lo <= 1'b0;
    n658_lo <= 1'b0;
    n661_lo <= 1'b0;
    n664_lo <= 1'b0;
    n667_lo <= 1'b0;
    n670_lo <= 1'b0;
    n673_lo <= 1'b0;
    n676_lo <= 1'b0;
    n679_lo <= 1'b0;
    n682_lo <= 1'b0;
    n685_lo <= 1'b0;
    n688_lo <= 1'b0;
    n691_lo <= 1'b0;
    n694_lo <= 1'b0;
    n697_lo <= 1'b0;
    n700_lo <= 1'b0;
    n703_lo <= 1'b0;
    n706_lo <= 1'b0;
    n709_lo <= 1'b0;
    n712_lo <= 1'b0;
    n715_lo <= 1'b0;
    n718_lo <= 1'b0;
    n721_lo <= 1'b0;
    n724_lo <= 1'b0;
    n727_lo <= 1'b0;
    n730_lo <= 1'b0;
    n733_lo <= 1'b0;
    n736_lo <= 1'b0;
    n739_lo <= 1'b0;
    n742_lo <= 1'b0;
    n745_lo <= 1'b0;
    n748_lo <= 1'b0;
    n751_lo <= 1'b0;
    n754_lo <= 1'b0;
    n757_lo <= 1'b0;
    n760_lo <= 1'b0;
    n763_lo <= 1'b0;
    n766_lo <= 1'b0;
  end
endmodule


