
module mymod
(
  G1_p,
  G1_n,
  G2_p,
  G2_n,
  G3_p,
  G3_n,
  G4_p,
  G4_n,
  G5_p,
  G5_n,
  G6_p,
  G6_n,
  G7_p,
  G7_n,
  G8_p,
  G8_n,
  G9_p,
  G9_n,
  G10_p,
  G10_n,
  G11_p,
  G11_n,
  G12_p,
  G12_n,
  G13_p,
  G13_n,
  G14_p,
  G14_n,
  G15_p,
  G15_n,
  G16_p,
  G16_n,
  G17_p,
  G17_n,
  G18_p,
  G18_n,
  G19_p,
  G19_n,
  G20_p,
  G20_n,
  G21_p,
  G21_n,
  G22_p,
  G22_n,
  G23_p,
  G23_n,
  G24_p,
  G24_n,
  G25_p,
  G25_n,
  G26_p,
  G26_n,
  G27_p,
  G27_n,
  G28_p,
  G28_n,
  G29_p,
  G29_n,
  G30_p,
  G30_n,
  G31_p,
  G31_n,
  G32_p,
  G32_n,
  G6257_p,
  G6258_p,
  G6259_p,
  G6260_p,
  G6261_p,
  G6262_p,
  G6263_p,
  G6264_p,
  G6265_p,
  G6266_p,
  G6267_p,
  G6268_p,
  G6269_p,
  G6270_p,
  G6271_p,
  G6272_p,
  G6273_p,
  G6274_p,
  G6275_p,
  G6276_p,
  G6277_p,
  G6278_p,
  G6279_p,
  G6280_p,
  G6281_p,
  G6282_p,
  G6283_p,
  G6284_p,
  G6285_p,
  G6286_p,
  G6287_p,
  G6288_n
);

  input G1_p;input G1_n;input G2_p;input G2_n;input G3_p;input G3_n;input G4_p;input G4_n;input G5_p;input G5_n;input G6_p;input G6_n;input G7_p;input G7_n;input G8_p;input G8_n;input G9_p;input G9_n;input G10_p;input G10_n;input G11_p;input G11_n;input G12_p;input G12_n;input G13_p;input G13_n;input G14_p;input G14_n;input G15_p;input G15_n;input G16_p;input G16_n;input G17_p;input G17_n;input G18_p;input G18_n;input G19_p;input G19_n;input G20_p;input G20_n;input G21_p;input G21_n;input G22_p;input G22_n;input G23_p;input G23_n;input G24_p;input G24_n;input G25_p;input G25_n;input G26_p;input G26_n;input G27_p;input G27_n;input G28_p;input G28_n;input G29_p;input G29_n;input G30_p;input G30_n;input G31_p;input G31_n;input G32_p;input G32_n;
  output G6257_p;output G6258_p;output G6259_p;output G6260_p;output G6261_p;output G6262_p;output G6263_p;output G6264_p;output G6265_p;output G6266_p;output G6267_p;output G6268_p;output G6269_p;output G6270_p;output G6271_p;output G6272_p;output G6273_p;output G6274_p;output G6275_p;output G6276_p;output G6277_p;output G6278_p;output G6279_p;output G6280_p;output G6281_p;output G6282_p;output G6283_p;output G6284_p;output G6285_p;output G6286_p;output G6287_p;output G6288_n;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire ffc_0_p;
  wire ffc_0_n;
  wire ffc_1_p;
  wire ffc_1_n;
  wire ffc_2_p;
  wire ffc_2_n;
  wire ffc_3_p;
  wire ffc_3_n;
  wire ffc_4_p;
  wire ffc_4_n;
  wire ffc_5_p;
  wire ffc_5_n;
  wire ffc_6_p;
  wire ffc_6_n;
  wire ffc_7_p;
  wire ffc_7_n;
  wire ffc_8_p;
  wire ffc_8_n;
  wire ffc_9_p;
  wire ffc_9_n;
  wire ffc_10_p;
  wire ffc_10_n;
  wire ffc_11_p;
  wire ffc_11_n;
  wire ffc_12_p;
  wire ffc_12_n;
  wire ffc_13_p;
  wire ffc_13_n;
  wire ffc_14_p;
  wire ffc_14_n;
  wire ffc_15_p;
  wire ffc_15_n;
  wire ffc_16_p;
  wire ffc_16_n;
  wire ffc_17_p;
  wire ffc_17_n;
  wire ffc_18_p;
  wire ffc_18_n;
  wire ffc_19_p;
  wire ffc_19_n;
  wire ffc_20_p;
  wire ffc_20_n;
  wire ffc_21_p;
  wire ffc_21_n;
  wire ffc_22_p;
  wire ffc_22_n;
  wire ffc_23_p;
  wire ffc_23_n;
  wire ffc_24_p;
  wire ffc_24_n;
  wire ffc_25_p;
  wire ffc_25_n;
  wire ffc_26_p;
  wire ffc_26_n;
  wire ffc_27_p;
  wire ffc_27_n;
  wire ffc_28_p;
  wire ffc_28_n;
  wire ffc_29_p;
  wire ffc_29_n;
  wire ffc_30_p;
  wire ffc_30_n;
  wire ffc_31_p;
  wire ffc_31_n;
  wire ffc_32_p;
  wire ffc_32_n;
  wire ffc_33_p;
  wire ffc_33_n;
  wire ffc_34_p;
  wire ffc_34_n;
  wire ffc_35_p;
  wire ffc_35_n;
  wire ffc_36_p;
  wire ffc_36_n;
  wire ffc_37_p;
  wire ffc_37_n;
  wire ffc_38_p;
  wire ffc_38_n;
  wire ffc_39_p;
  wire ffc_39_n;
  wire ffc_40_p;
  wire ffc_40_n;
  wire ffc_41_p;
  wire ffc_41_n;
  wire ffc_42_p;
  wire ffc_42_n;
  wire ffc_43_p;
  wire ffc_43_n;
  wire ffc_44_p;
  wire ffc_44_n;
  wire ffc_45_p;
  wire ffc_45_n;
  wire ffc_46_p;
  wire ffc_46_n;
  wire ffc_47_p;
  wire ffc_47_n;
  wire ffc_48_p;
  wire ffc_48_n;
  wire ffc_49_p;
  wire ffc_49_n;
  wire ffc_50_p;
  wire ffc_50_n;
  wire ffc_51_p;
  wire ffc_51_n;
  wire ffc_52_p;
  wire ffc_52_n;
  wire ffc_53_p;
  wire ffc_53_n;
  wire ffc_54_p;
  wire ffc_54_n;
  wire ffc_55_p;
  wire ffc_55_n;
  wire ffc_56_p;
  wire ffc_56_n;
  wire ffc_57_p;
  wire ffc_57_n;
  wire ffc_58_p;
  wire ffc_58_n;
  wire ffc_59_p;
  wire ffc_59_n;
  wire ffc_60_p;
  wire ffc_60_n;
  wire ffc_61_p;
  wire ffc_61_n;
  wire ffc_62_p;
  wire ffc_62_n;
  wire ffc_63_p;
  wire ffc_63_n;
  wire ffc_64_p;
  wire ffc_64_n;
  wire ffc_65_p;
  wire ffc_65_n;
  wire ffc_66_p;
  wire ffc_66_n;
  wire ffc_67_p;
  wire ffc_67_n;
  wire ffc_68_p;
  wire ffc_68_n;
  wire ffc_69_p;
  wire ffc_69_n;
  wire ffc_70_p;
  wire ffc_70_n;
  wire ffc_71_p;
  wire ffc_71_n;
  wire ffc_72_p;
  wire ffc_72_n;
  wire ffc_73_p;
  wire ffc_73_n;
  wire ffc_74_p;
  wire ffc_74_n;
  wire ffc_75_p;
  wire ffc_75_n;
  wire ffc_76_p;
  wire ffc_76_n;
  wire ffc_77_p;
  wire ffc_77_n;
  wire ffc_78_p;
  wire ffc_78_n;
  wire ffc_79_p;
  wire ffc_79_n;
  wire ffc_80_p;
  wire ffc_80_n;
  wire ffc_81_p;
  wire ffc_81_n;
  wire ffc_82_p;
  wire ffc_82_n;
  wire ffc_83_p;
  wire ffc_83_n;
  wire ffc_84_p;
  wire ffc_84_n;
  wire ffc_85_p;
  wire ffc_85_n;
  wire ffc_86_p;
  wire ffc_86_n;
  wire ffc_87_p;
  wire ffc_87_n;
  wire ffc_88_p;
  wire ffc_88_n;
  wire ffc_89_p;
  wire ffc_89_n;
  wire ffc_90_p;
  wire ffc_90_n;
  wire ffc_91_p;
  wire ffc_91_n;
  wire ffc_92_p;
  wire ffc_92_n;
  wire ffc_93_p;
  wire ffc_93_n;
  wire ffc_94_p;
  wire ffc_94_n;
  wire ffc_95_p;
  wire ffc_95_n;
  wire ffc_96_p;
  wire ffc_96_n;
  wire ffc_97_p;
  wire ffc_97_n;
  wire ffc_98_p;
  wire ffc_98_n;
  wire ffc_99_p;
  wire ffc_99_n;
  wire ffc_100_p;
  wire ffc_100_n;
  wire ffc_101_p;
  wire ffc_101_n;
  wire ffc_102_p;
  wire ffc_102_n;
  wire ffc_103_p;
  wire ffc_103_n;
  wire ffc_104_p;
  wire ffc_104_n;
  wire ffc_105_p;
  wire ffc_105_n;
  wire ffc_106_p;
  wire ffc_106_n;
  wire ffc_107_p;
  wire ffc_107_n;
  wire ffc_108_p;
  wire ffc_108_n;
  wire ffc_109_p;
  wire ffc_109_n;
  wire ffc_110_p;
  wire ffc_110_n;
  wire ffc_111_p;
  wire ffc_111_n;
  wire ffc_112_p;
  wire ffc_112_n;
  wire ffc_113_p;
  wire ffc_113_n;
  wire ffc_114_p;
  wire ffc_114_n;
  wire ffc_115_p;
  wire ffc_115_n;
  wire ffc_116_p;
  wire ffc_116_n;
  wire ffc_117_p;
  wire ffc_117_n;
  wire ffc_118_p;
  wire ffc_118_n;
  wire ffc_119_p;
  wire ffc_119_n;
  wire ffc_120_p;
  wire ffc_120_n;
  wire ffc_121_p;
  wire ffc_121_n;
  wire ffc_122_p;
  wire ffc_122_n;
  wire ffc_123_p;
  wire ffc_123_n;
  wire ffc_124_p;
  wire ffc_124_n;
  wire ffc_125_p;
  wire ffc_125_n;
  wire ffc_126_p;
  wire ffc_126_n;
  wire ffc_127_p;
  wire ffc_127_n;
  wire ffc_128_p;
  wire ffc_128_n;
  wire ffc_129_p;
  wire ffc_129_n;
  wire ffc_130_p;
  wire ffc_130_n;
  wire ffc_131_p;
  wire ffc_131_n;
  wire ffc_132_p;
  wire ffc_132_n;
  wire ffc_133_p;
  wire ffc_133_n;
  wire ffc_134_p;
  wire ffc_134_n;
  wire ffc_135_p;
  wire ffc_135_n;
  wire ffc_136_p;
  wire ffc_136_n;
  wire ffc_137_p;
  wire ffc_137_n;
  wire ffc_138_p;
  wire ffc_138_n;
  wire ffc_139_p;
  wire ffc_139_n;
  wire ffc_140_p;
  wire ffc_140_n;
  wire ffc_141_p;
  wire ffc_141_n;
  wire ffc_142_p;
  wire ffc_142_n;
  wire ffc_143_p;
  wire ffc_143_n;
  wire ffc_144_p;
  wire ffc_144_n;
  wire ffc_145_p;
  wire ffc_145_n;
  wire ffc_146_p;
  wire ffc_146_n;
  wire ffc_147_p;
  wire ffc_147_n;
  wire ffc_148_p;
  wire ffc_148_n;
  wire ffc_149_p;
  wire ffc_149_n;
  wire ffc_150_p;
  wire ffc_150_n;
  wire ffc_151_p;
  wire ffc_151_n;
  wire ffc_152_p;
  wire ffc_152_n;
  wire ffc_153_p;
  wire ffc_153_n;
  wire ffc_154_p;
  wire ffc_154_n;
  wire ffc_155_p;
  wire ffc_155_n;
  wire ffc_156_p;
  wire ffc_156_n;
  wire ffc_157_p;
  wire ffc_157_n;
  wire ffc_158_p;
  wire ffc_158_n;
  wire ffc_159_p;
  wire ffc_159_n;
  wire ffc_160_p;
  wire ffc_160_n;
  wire ffc_161_p;
  wire ffc_161_n;
  wire ffc_162_p;
  wire ffc_162_n;
  wire ffc_163_p;
  wire ffc_163_n;
  wire ffc_164_p;
  wire ffc_164_n;
  wire ffc_165_p;
  wire ffc_165_n;
  wire ffc_166_p;
  wire ffc_166_n;
  wire ffc_167_p;
  wire ffc_167_n;
  wire ffc_168_p;
  wire ffc_168_n;
  wire ffc_169_p;
  wire ffc_169_n;
  wire ffc_170_p;
  wire ffc_170_n;
  wire ffc_171_p;
  wire ffc_171_n;
  wire ffc_172_p;
  wire ffc_172_n;
  wire ffc_173_p;
  wire ffc_173_n;
  wire ffc_174_p;
  wire ffc_174_n;
  wire ffc_175_p;
  wire ffc_175_n;
  wire ffc_176_p;
  wire ffc_176_n;
  wire ffc_177_p;
  wire ffc_177_n;
  wire ffc_178_p;
  wire ffc_178_n;
  wire ffc_179_p;
  wire ffc_179_n;
  wire ffc_180_p;
  wire ffc_180_n;
  wire ffc_181_p;
  wire ffc_181_n;
  wire ffc_182_p;
  wire ffc_182_n;
  wire ffc_183_p;
  wire ffc_183_n;
  wire ffc_184_p;
  wire ffc_184_n;
  wire ffc_185_p;
  wire ffc_185_n;
  wire ffc_186_p;
  wire ffc_186_n;
  wire ffc_187_p;
  wire ffc_187_n;
  wire ffc_188_p;
  wire ffc_188_n;
  wire ffc_189_p;
  wire ffc_189_n;
  wire ffc_190_p;
  wire ffc_190_n;
  wire ffc_191_p;
  wire ffc_191_n;
  wire ffc_192_p;
  wire ffc_192_n;
  wire ffc_193_p;
  wire ffc_193_n;
  wire ffc_194_p;
  wire ffc_194_n;
  wire ffc_195_p;
  wire ffc_195_n;
  wire ffc_196_p;
  wire ffc_196_n;
  wire ffc_197_p;
  wire ffc_197_n;
  wire ffc_198_p;
  wire ffc_198_n;
  wire ffc_199_p;
  wire ffc_199_n;
  wire ffc_200_p;
  wire ffc_200_n;
  wire ffc_201_p;
  wire ffc_201_n;
  wire ffc_202_p;
  wire ffc_202_n;
  wire ffc_203_p;
  wire ffc_203_n;
  wire ffc_204_p;
  wire ffc_204_n;
  wire ffc_205_p;
  wire ffc_205_n;
  wire ffc_206_p;
  wire ffc_206_n;
  wire ffc_207_p;
  wire ffc_207_n;
  wire ffc_208_p;
  wire ffc_208_n;
  wire ffc_209_p;
  wire ffc_209_n;
  wire ffc_210_p;
  wire ffc_210_n;
  wire ffc_211_p;
  wire ffc_211_n;
  wire ffc_212_p;
  wire ffc_212_n;
  wire ffc_213_p;
  wire ffc_213_n;
  wire ffc_214_p;
  wire ffc_214_n;
  wire ffc_215_p;
  wire ffc_215_n;
  wire ffc_216_p;
  wire ffc_216_n;
  wire ffc_217_p;
  wire ffc_217_n;
  wire ffc_218_p;
  wire ffc_218_n;
  wire ffc_219_p;
  wire ffc_219_n;
  wire ffc_220_p;
  wire ffc_220_n;
  wire ffc_221_p;
  wire ffc_221_n;
  wire ffc_222_p;
  wire ffc_222_n;
  wire ffc_223_p;
  wire ffc_223_n;
  wire ffc_224_p;
  wire ffc_224_n;
  wire ffc_225_p;
  wire ffc_225_n;
  wire ffc_226_p;
  wire ffc_226_n;
  wire ffc_227_p;
  wire ffc_227_n;
  wire ffc_228_p;
  wire ffc_228_n;
  wire ffc_229_p;
  wire ffc_229_n;
  wire ffc_230_p;
  wire ffc_230_n;
  wire ffc_231_p;
  wire ffc_231_n;
  wire ffc_232_p;
  wire ffc_232_n;
  wire ffc_233_p;
  wire ffc_233_n;
  wire ffc_234_p;
  wire ffc_234_n;
  wire ffc_235_p;
  wire ffc_235_n;
  wire ffc_236_p;
  wire ffc_236_n;
  wire ffc_237_p;
  wire ffc_237_n;
  wire ffc_238_p;
  wire ffc_238_n;
  wire ffc_239_p;
  wire ffc_239_n;
  wire ffc_240_p;
  wire ffc_240_n;
  wire ffc_241_p;
  wire ffc_241_n;
  wire ffc_242_p;
  wire ffc_242_n;
  wire ffc_243_p;
  wire ffc_243_n;
  wire ffc_244_p;
  wire ffc_244_n;
  wire ffc_245_p;
  wire ffc_245_n;
  wire ffc_246_p;
  wire ffc_246_n;
  wire ffc_247_p;
  wire ffc_247_n;
  wire ffc_248_p;
  wire ffc_248_n;
  wire ffc_249_p;
  wire ffc_249_n;
  wire ffc_250_p;
  wire ffc_250_n;
  wire ffc_251_p;
  wire ffc_251_n;
  wire ffc_252_p;
  wire ffc_252_n;
  wire ffc_253_p;
  wire ffc_253_n;
  wire ffc_254_p;
  wire ffc_254_n;
  wire ffc_255_p;
  wire ffc_255_n;
  wire ffc_256_p;
  wire ffc_256_n;
  wire ffc_257_p;
  wire ffc_257_n;
  wire ffc_258_p;
  wire ffc_258_n;
  wire ffc_259_p;
  wire ffc_259_n;
  wire ffc_260_p;
  wire ffc_260_n;
  wire ffc_261_p;
  wire ffc_261_n;
  wire ffc_262_p;
  wire ffc_262_n;
  wire ffc_263_p;
  wire ffc_263_n;
  wire ffc_264_p;
  wire ffc_264_n;
  wire ffc_265_p;
  wire ffc_265_n;
  wire ffc_266_p;
  wire ffc_266_n;
  wire ffc_267_p;
  wire ffc_267_n;
  wire ffc_268_p;
  wire ffc_268_n;
  wire ffc_269_p;
  wire ffc_269_n;
  wire ffc_270_p;
  wire ffc_270_n;
  wire ffc_271_p;
  wire ffc_271_n;
  wire ffc_272_p;
  wire ffc_272_n;
  wire ffc_273_p;
  wire ffc_273_n;
  wire ffc_274_p;
  wire ffc_274_n;
  wire ffc_275_p;
  wire ffc_275_n;
  wire ffc_276_p;
  wire ffc_276_n;
  wire ffc_277_p;
  wire ffc_277_n;
  wire ffc_278_p;
  wire ffc_278_n;
  wire ffc_279_p;
  wire ffc_279_n;
  wire ffc_280_p;
  wire ffc_280_n;
  wire ffc_281_p;
  wire ffc_281_n;
  wire ffc_282_p;
  wire ffc_282_n;
  wire ffc_283_p;
  wire ffc_283_n;
  wire ffc_284_p;
  wire ffc_284_n;
  wire ffc_285_p;
  wire ffc_285_n;
  wire ffc_286_p;
  wire ffc_286_n;
  wire ffc_287_p;
  wire ffc_287_n;
  wire ffc_288_p;
  wire ffc_288_n;
  wire ffc_289_p;
  wire ffc_289_n;
  wire ffc_290_p;
  wire ffc_290_n;
  wire ffc_291_p;
  wire ffc_291_n;
  wire ffc_292_p;
  wire ffc_292_n;
  wire ffc_293_p;
  wire ffc_293_n;
  wire ffc_294_p;
  wire ffc_294_n;
  wire ffc_295_p;
  wire ffc_295_n;
  wire ffc_296_p;
  wire ffc_296_n;
  wire ffc_297_p;
  wire ffc_297_n;
  wire ffc_298_p;
  wire ffc_298_n;
  wire ffc_299_p;
  wire ffc_299_n;
  wire ffc_300_p;
  wire ffc_300_n;
  wire ffc_301_p;
  wire ffc_301_n;
  wire ffc_302_p;
  wire ffc_302_n;
  wire ffc_303_p;
  wire ffc_303_n;
  wire ffc_304_p;
  wire ffc_304_n;
  wire ffc_305_p;
  wire ffc_305_n;
  wire ffc_306_p;
  wire ffc_306_n;
  wire ffc_307_p;
  wire ffc_307_n;
  wire ffc_308_p;
  wire ffc_308_n;
  wire ffc_309_p;
  wire ffc_309_n;
  wire ffc_310_p;
  wire ffc_310_n;
  wire ffc_311_p;
  wire ffc_311_n;
  wire ffc_312_p;
  wire ffc_312_n;
  wire ffc_313_p;
  wire ffc_313_n;
  wire ffc_314_p;
  wire ffc_314_n;
  wire ffc_315_p;
  wire ffc_315_n;
  wire ffc_316_p;
  wire ffc_316_n;
  wire ffc_317_p;
  wire ffc_317_n;
  wire ffc_318_p;
  wire ffc_318_n;
  wire ffc_319_p;
  wire ffc_319_n;
  wire ffc_320_p;
  wire ffc_320_n;
  wire ffc_321_p;
  wire ffc_321_n;
  wire ffc_322_p;
  wire ffc_322_n;
  wire ffc_323_p;
  wire ffc_323_n;
  wire ffc_324_p;
  wire ffc_324_n;
  wire ffc_325_p;
  wire ffc_325_n;
  wire ffc_326_p;
  wire ffc_326_n;
  wire ffc_327_p;
  wire ffc_327_n;
  wire ffc_328_p;
  wire ffc_328_n;
  wire ffc_329_p;
  wire ffc_329_n;
  wire ffc_330_p;
  wire ffc_330_n;
  wire ffc_331_p;
  wire ffc_331_n;
  wire ffc_332_p;
  wire ffc_332_n;
  wire ffc_333_p;
  wire ffc_333_n;
  wire ffc_334_p;
  wire ffc_334_n;
  wire ffc_335_p;
  wire ffc_335_n;
  wire ffc_336_p;
  wire ffc_336_n;
  wire ffc_337_p;
  wire ffc_337_n;
  wire ffc_338_p;
  wire ffc_338_n;
  wire ffc_339_p;
  wire ffc_339_n;
  wire ffc_340_p;
  wire ffc_340_n;
  wire ffc_341_p;
  wire ffc_341_n;
  wire ffc_342_p;
  wire ffc_342_n;
  wire ffc_343_p;
  wire ffc_343_n;
  wire ffc_344_p;
  wire ffc_344_n;
  wire ffc_345_p;
  wire ffc_345_n;
  wire ffc_346_p;
  wire ffc_346_n;
  wire ffc_347_p;
  wire ffc_347_n;
  wire ffc_348_p;
  wire ffc_348_n;
  wire ffc_349_p;
  wire ffc_349_n;
  wire ffc_350_p;
  wire ffc_350_n;
  wire ffc_351_p;
  wire ffc_351_n;
  wire ffc_352_p;
  wire ffc_352_n;
  wire ffc_353_p;
  wire ffc_353_n;
  wire ffc_354_p;
  wire ffc_354_n;
  wire ffc_355_p;
  wire ffc_355_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire g693_p;
  wire g693_n;
  wire g694_p;
  wire g694_n;
  wire g695_p;
  wire g695_n;
  wire g696_p;
  wire g696_n;
  wire g697_p;
  wire g697_n;
  wire g698_p;
  wire g698_n;
  wire g699_p;
  wire g699_n;
  wire g700_p;
  wire g700_n;
  wire g701_p;
  wire g701_n;
  wire g702_p;
  wire g702_n;
  wire g703_p;
  wire g703_n;
  wire g704_p;
  wire g704_n;
  wire g705_p;
  wire g705_n;
  wire g706_p;
  wire g706_n;
  wire g707_p;
  wire g707_n;
  wire g708_p;
  wire g708_n;
  wire g709_p;
  wire g709_n;
  wire g710_p;
  wire g710_n;
  wire g711_p;
  wire g711_n;
  wire g712_p;
  wire g712_n;
  wire g713_p;
  wire g713_n;
  wire g714_p;
  wire g714_n;
  wire g715_p;
  wire g715_n;
  wire g716_p;
  wire g716_n;
  wire g717_p;
  wire g717_n;
  wire g718_p;
  wire g718_n;
  wire g719_p;
  wire g719_n;
  wire g720_p;
  wire g720_n;
  wire g721_p;
  wire g721_n;
  wire g722_p;
  wire g722_n;
  wire g723_p;
  wire g723_n;
  wire g724_p;
  wire g724_n;
  wire g725_p;
  wire g725_n;
  wire g726_p;
  wire g726_n;
  wire g727_p;
  wire g727_n;
  wire g728_p;
  wire g728_n;
  wire g729_p;
  wire g729_n;
  wire g730_p;
  wire g730_n;
  wire g731_p;
  wire g731_n;
  wire g732_p;
  wire g732_n;
  wire g733_p;
  wire g733_n;
  wire g734_p;
  wire g734_n;
  wire g735_p;
  wire g735_n;
  wire g736_p;
  wire g736_n;
  wire g737_p;
  wire g737_n;
  wire g738_p;
  wire g738_n;
  wire g739_p;
  wire g739_n;
  wire g740_p;
  wire g740_n;
  wire g741_p;
  wire g741_n;
  wire g742_p;
  wire g742_n;
  wire g743_p;
  wire g743_n;
  wire g744_p;
  wire g744_n;
  wire g745_p;
  wire g745_n;
  wire g746_p;
  wire g746_n;
  wire g747_p;
  wire g747_n;
  wire g748_p;
  wire g748_n;
  wire g749_p;
  wire g749_n;
  wire g750_p;
  wire g750_n;
  wire g751_p;
  wire g751_n;
  wire g752_p;
  wire g752_n;
  wire g753_p;
  wire g753_n;
  wire g754_p;
  wire g754_n;
  wire g755_p;
  wire g755_n;
  wire g756_p;
  wire g756_n;
  wire g757_p;
  wire g757_n;
  wire g758_p;
  wire g758_n;
  wire g759_p;
  wire g759_n;
  wire g760_p;
  wire g760_n;
  wire g761_p;
  wire g761_n;
  wire g762_p;
  wire g762_n;
  wire g763_p;
  wire g763_n;
  wire g764_p;
  wire g764_n;
  wire g765_p;
  wire g765_n;
  wire g766_p;
  wire g766_n;
  wire g767_p;
  wire g767_n;
  wire g768_p;
  wire g768_n;
  wire g769_p;
  wire g769_n;
  wire g770_p;
  wire g770_n;
  wire g771_p;
  wire g771_n;
  wire g772_p;
  wire g772_n;
  wire g773_p;
  wire g773_n;
  wire g774_p;
  wire g774_n;
  wire g775_p;
  wire g775_n;
  wire g776_p;
  wire g776_n;
  wire g777_p;
  wire g777_n;
  wire g778_p;
  wire g778_n;
  wire g779_p;
  wire g779_n;
  wire g780_p;
  wire g780_n;
  wire g781_p;
  wire g781_n;
  wire g782_p;
  wire g782_n;
  wire g783_p;
  wire g783_n;
  wire g784_p;
  wire g784_n;
  wire g785_p;
  wire g785_n;
  wire g786_p;
  wire g786_n;
  wire g787_p;
  wire g787_n;
  wire g788_p;
  wire g788_n;
  wire g789_p;
  wire g789_n;
  wire g790_p;
  wire g790_n;
  wire g791_p;
  wire g791_n;
  wire g792_p;
  wire g792_n;
  wire g793_p;
  wire g793_n;
  wire g794_p;
  wire g794_n;
  wire g795_p;
  wire g795_n;
  wire g796_p;
  wire g796_n;
  wire g797_p;
  wire g797_n;
  wire g798_p;
  wire g798_n;
  wire g799_p;
  wire g799_n;
  wire g800_p;
  wire g800_n;
  wire g801_p;
  wire g801_n;
  wire g802_p;
  wire g802_n;
  wire g803_p;
  wire g803_n;
  wire g804_p;
  wire g804_n;
  wire g805_p;
  wire g805_n;
  wire g806_p;
  wire g806_n;
  wire g807_p;
  wire g807_n;
  wire g808_p;
  wire g808_n;
  wire g809_p;
  wire g809_n;
  wire g810_p;
  wire g810_n;
  wire g811_p;
  wire g811_n;
  wire g812_p;
  wire g812_n;
  wire g813_p;
  wire g813_n;
  wire g814_p;
  wire g814_n;
  wire g815_p;
  wire g815_n;
  wire g816_p;
  wire g816_n;
  wire g817_p;
  wire g817_n;
  wire g818_p;
  wire g818_n;
  wire g819_p;
  wire g819_n;
  wire g820_p;
  wire g820_n;
  wire g821_p;
  wire g821_n;
  wire g822_p;
  wire g822_n;
  wire g823_p;
  wire g823_n;
  wire g824_p;
  wire g824_n;
  wire g825_p;
  wire g825_n;
  wire g826_p;
  wire g826_n;
  wire g827_p;
  wire g827_n;
  wire g828_p;
  wire g828_n;
  wire g829_p;
  wire g829_n;
  wire g830_p;
  wire g830_n;
  wire g831_p;
  wire g831_n;
  wire g832_p;
  wire g832_n;
  wire g833_p;
  wire g833_n;
  wire g834_p;
  wire g834_n;
  wire g835_p;
  wire g835_n;
  wire g836_p;
  wire g836_n;
  wire g837_p;
  wire g837_n;
  wire g838_p;
  wire g838_n;
  wire g839_p;
  wire g839_n;
  wire g840_p;
  wire g840_n;
  wire g841_p;
  wire g841_n;
  wire g842_p;
  wire g842_n;
  wire g843_p;
  wire g843_n;
  wire g844_p;
  wire g844_n;
  wire g845_p;
  wire g845_n;
  wire g846_p;
  wire g846_n;
  wire g847_p;
  wire g847_n;
  wire g848_p;
  wire g848_n;
  wire g849_p;
  wire g849_n;
  wire g850_p;
  wire g850_n;
  wire g851_p;
  wire g851_n;
  wire g852_p;
  wire g852_n;
  wire g853_p;
  wire g853_n;
  wire g854_p;
  wire g854_n;
  wire g855_p;
  wire g855_n;
  wire g856_p;
  wire g856_n;
  wire g857_p;
  wire g857_n;
  wire g858_p;
  wire g858_n;
  wire g859_p;
  wire g859_n;
  wire g860_p;
  wire g860_n;
  wire g861_p;
  wire g861_n;
  wire g862_p;
  wire g862_n;
  wire g863_p;
  wire g863_n;
  wire g864_p;
  wire g864_n;
  wire g865_p;
  wire g865_n;
  wire g866_p;
  wire g866_n;
  wire g867_p;
  wire g867_n;
  wire g868_p;
  wire g868_n;
  wire g869_p;
  wire g869_n;
  wire g870_p;
  wire g870_n;
  wire g871_p;
  wire g871_n;
  wire g872_p;
  wire g872_n;
  wire g873_p;
  wire g873_n;
  wire g874_p;
  wire g874_n;
  wire g875_p;
  wire g875_n;
  wire g876_p;
  wire g876_n;
  wire g877_p;
  wire g877_n;
  wire g878_p;
  wire g878_n;
  wire g879_p;
  wire g879_n;
  wire g880_p;
  wire g880_n;
  wire g881_p;
  wire g881_n;
  wire g882_p;
  wire g882_n;
  wire g883_p;
  wire g883_n;
  wire g884_p;
  wire g884_n;
  wire g885_p;
  wire g885_n;
  wire g886_p;
  wire g886_n;
  wire g887_p;
  wire g887_n;
  wire g888_p;
  wire g888_n;
  wire g889_p;
  wire g889_n;
  wire g890_p;
  wire g890_n;
  wire g891_p;
  wire g891_n;
  wire g892_p;
  wire g892_n;
  wire g893_p;
  wire g893_n;
  wire g894_p;
  wire g894_n;
  wire g895_p;
  wire g895_n;
  wire g896_p;
  wire g896_n;
  wire g897_p;
  wire g897_n;
  wire g898_p;
  wire g898_n;
  wire g899_p;
  wire g899_n;
  wire g900_p;
  wire g900_n;
  wire g901_p;
  wire g901_n;
  wire g902_p;
  wire g902_n;
  wire g903_p;
  wire g903_n;
  wire g904_p;
  wire g904_n;
  wire g905_p;
  wire g905_n;
  wire g906_p;
  wire g906_n;
  wire g907_p;
  wire g907_n;
  wire g908_p;
  wire g908_n;
  wire g909_p;
  wire g909_n;
  wire g910_p;
  wire g910_n;
  wire g911_p;
  wire g911_n;
  wire g912_p;
  wire g912_n;
  wire g913_p;
  wire g913_n;
  wire g914_p;
  wire g914_n;
  wire g915_p;
  wire g915_n;
  wire g916_p;
  wire g916_n;
  wire g917_p;
  wire g917_n;
  wire g918_p;
  wire g918_n;
  wire g919_p;
  wire g919_n;
  wire g920_p;
  wire g920_n;
  wire g921_p;
  wire g921_n;
  wire g922_p;
  wire g922_n;
  wire g923_p;
  wire g923_n;
  wire g924_p;
  wire g924_n;
  wire g925_p;
  wire g925_n;
  wire g926_p;
  wire g926_n;
  wire g927_p;
  wire g927_n;
  wire g928_p;
  wire g928_n;
  wire g929_p;
  wire g929_n;
  wire g930_p;
  wire g930_n;
  wire g931_p;
  wire g931_n;
  wire g932_p;
  wire g932_n;
  wire g933_p;
  wire g933_n;
  wire g934_p;
  wire g934_n;
  wire g935_p;
  wire g935_n;
  wire g936_p;
  wire g936_n;
  wire g937_p;
  wire g937_n;
  wire g938_p;
  wire g938_n;
  wire g939_p;
  wire g939_n;
  wire g940_p;
  wire g940_n;
  wire g941_p;
  wire g941_n;
  wire g942_p;
  wire g942_n;
  wire g943_p;
  wire g943_n;
  wire g944_p;
  wire g944_n;
  wire g945_p;
  wire g945_n;
  wire g946_p;
  wire g946_n;
  wire g947_p;
  wire g947_n;
  wire g948_p;
  wire g948_n;
  wire g949_p;
  wire g949_n;
  wire g950_p;
  wire g950_n;
  wire g951_p;
  wire g951_n;
  wire g952_p;
  wire g952_n;
  wire g953_p;
  wire g953_n;
  wire g954_p;
  wire g954_n;
  wire g955_p;
  wire g955_n;
  wire g956_p;
  wire g956_n;
  wire g957_p;
  wire g957_n;
  wire g958_p;
  wire g958_n;
  wire g959_p;
  wire g959_n;
  wire g960_p;
  wire g960_n;
  wire g961_p;
  wire g961_n;
  wire g962_p;
  wire g962_n;
  wire g963_p;
  wire g963_n;
  wire g964_p;
  wire g964_n;
  wire g965_p;
  wire g965_n;
  wire g966_p;
  wire g966_n;
  wire g967_p;
  wire g967_n;
  wire g968_p;
  wire g968_n;
  wire g969_p;
  wire g969_n;
  wire g970_p;
  wire g970_n;
  wire g971_p;
  wire g971_n;
  wire g972_p;
  wire g972_n;
  wire g973_p;
  wire g973_n;
  wire g974_p;
  wire g974_n;
  wire g975_p;
  wire g975_n;
  wire g976_p;
  wire g976_n;
  wire g977_p;
  wire g977_n;
  wire g978_p;
  wire g978_n;
  wire g979_p;
  wire g979_n;
  wire g980_p;
  wire g980_n;
  wire g981_p;
  wire g981_n;
  wire g982_p;
  wire g982_n;
  wire g983_p;
  wire g983_n;
  wire g984_p;
  wire g984_n;
  wire g985_p;
  wire g985_n;
  wire g986_p;
  wire g986_n;
  wire g987_p;
  wire g987_n;
  wire g988_p;
  wire g988_n;
  wire g989_p;
  wire g989_n;
  wire g990_p;
  wire g990_n;
  wire g991_p;
  wire g991_n;
  wire g992_p;
  wire g992_n;
  wire g993_p;
  wire g993_n;
  wire g994_p;
  wire g994_n;
  wire g995_p;
  wire g995_n;
  wire g996_p;
  wire g996_n;
  wire g997_p;
  wire g997_n;
  wire g998_p;
  wire g998_n;
  wire g999_p;
  wire g999_n;
  wire g1000_p;
  wire g1000_n;
  wire g1001_p;
  wire g1001_n;
  wire g1002_p;
  wire g1002_n;
  wire g1003_p;
  wire g1003_n;
  wire g1004_p;
  wire g1004_n;
  wire g1005_p;
  wire g1005_n;
  wire g1006_p;
  wire g1006_n;
  wire g1007_p;
  wire g1007_n;
  wire g1008_p;
  wire g1008_n;
  wire g1009_p;
  wire g1009_n;
  wire g1010_p;
  wire g1010_n;
  wire g1011_p;
  wire g1011_n;
  wire g1012_p;
  wire g1012_n;
  wire g1013_p;
  wire g1013_n;
  wire g1014_p;
  wire g1014_n;
  wire g1015_p;
  wire g1015_n;
  wire g1016_p;
  wire g1016_n;
  wire g1017_p;
  wire g1017_n;
  wire g1018_p;
  wire g1018_n;
  wire g1019_p;
  wire g1019_n;
  wire g1020_p;
  wire g1020_n;
  wire g1021_p;
  wire g1021_n;
  wire g1022_p;
  wire g1022_n;
  wire g1023_p;
  wire g1023_n;
  wire g1024_p;
  wire g1024_n;
  wire g1025_p;
  wire g1025_n;
  wire g1026_p;
  wire g1026_n;
  wire g1027_p;
  wire g1027_n;
  wire g1028_p;
  wire g1028_n;
  wire g1029_p;
  wire g1029_n;
  wire g1030_p;
  wire g1030_n;
  wire g1031_p;
  wire g1031_n;
  wire g1032_p;
  wire g1032_n;
  wire g1033_p;
  wire g1033_n;
  wire g1034_p;
  wire g1034_n;
  wire g1035_p;
  wire g1035_n;
  wire g1036_p;
  wire g1036_n;
  wire g1037_p;
  wire g1037_n;
  wire g1038_p;
  wire g1038_n;
  wire g1039_p;
  wire g1039_n;
  wire g1040_p;
  wire g1040_n;
  wire g1041_p;
  wire g1041_n;
  wire g1042_p;
  wire g1042_n;
  wire g1043_p;
  wire g1043_n;
  wire g1044_p;
  wire g1044_n;
  wire g1045_p;
  wire g1045_n;
  wire g1046_p;
  wire g1046_n;
  wire g1047_p;
  wire g1047_n;
  wire g1048_p;
  wire g1048_n;
  wire g1049_p;
  wire g1049_n;
  wire g1050_p;
  wire g1050_n;
  wire g1051_p;
  wire g1051_n;
  wire g1052_p;
  wire g1052_n;
  wire g1053_p;
  wire g1053_n;
  wire g1054_p;
  wire g1054_n;
  wire g1055_p;
  wire g1055_n;
  wire g1056_p;
  wire g1056_n;
  wire g1057_p;
  wire g1057_n;
  wire g1058_p;
  wire g1058_n;
  wire g1059_p;
  wire g1059_n;
  wire g1060_p;
  wire g1060_n;
  wire g1061_p;
  wire g1061_n;
  wire g1062_p;
  wire g1062_n;
  wire g1063_p;
  wire g1063_n;
  wire g1064_p;
  wire g1064_n;
  wire g1065_p;
  wire g1065_n;
  wire g1066_p;
  wire g1066_n;
  wire g1067_p;
  wire g1067_n;
  wire g1068_p;
  wire g1068_n;
  wire g1069_p;
  wire g1069_n;
  wire g1070_p;
  wire g1070_n;
  wire g1071_p;
  wire g1071_n;
  wire g1072_p;
  wire g1072_n;
  wire g1073_p;
  wire g1073_n;
  wire g1074_p;
  wire g1074_n;
  wire g1075_p;
  wire g1075_n;
  wire g1076_p;
  wire g1076_n;
  wire g1077_p;
  wire g1077_n;
  wire g1078_p;
  wire g1078_n;
  wire g1079_p;
  wire g1079_n;
  wire g1080_p;
  wire g1080_n;
  wire g1081_p;
  wire g1081_n;
  wire g1082_p;
  wire g1082_n;
  wire g1083_p;
  wire g1083_n;
  wire g1084_p;
  wire g1084_n;
  wire g1085_p;
  wire g1085_n;
  wire g1086_p;
  wire g1086_n;
  wire g1087_p;
  wire g1087_n;
  wire g1088_p;
  wire g1088_n;
  wire g1089_p;
  wire g1089_n;
  wire g1090_p;
  wire g1090_n;
  wire g1091_p;
  wire g1091_n;
  wire g1092_p;
  wire g1092_n;
  wire g1093_p;
  wire g1093_n;
  wire g1094_p;
  wire g1094_n;
  wire g1095_p;
  wire g1095_n;
  wire g1096_p;
  wire g1096_n;
  wire g1097_p;
  wire g1097_n;
  wire g1098_p;
  wire g1098_n;
  wire g1099_p;
  wire g1099_n;
  wire g1100_p;
  wire g1100_n;
  wire g1101_p;
  wire g1101_n;
  wire g1102_p;
  wire g1102_n;
  wire g1103_p;
  wire g1103_n;
  wire g1104_p;
  wire g1104_n;
  wire g1105_p;
  wire g1105_n;
  wire g1106_p;
  wire g1106_n;
  wire g1107_p;
  wire g1107_n;
  wire g1108_p;
  wire g1108_n;
  wire g1109_p;
  wire g1109_n;
  wire g1110_p;
  wire g1110_n;
  wire g1111_p;
  wire g1111_n;
  wire g1112_p;
  wire g1112_n;
  wire g1113_p;
  wire g1113_n;
  wire g1114_p;
  wire g1114_n;
  wire g1115_p;
  wire g1115_n;
  wire g1116_p;
  wire g1116_n;
  wire g1117_p;
  wire g1117_n;
  wire g1118_p;
  wire g1118_n;
  wire g1119_p;
  wire g1119_n;
  wire g1120_p;
  wire g1120_n;
  wire g1121_p;
  wire g1121_n;
  wire g1122_p;
  wire g1122_n;
  wire g1123_p;
  wire g1123_n;
  wire g1124_p;
  wire g1124_n;
  wire g1125_p;
  wire g1125_n;
  wire g1126_p;
  wire g1126_n;
  wire g1127_p;
  wire g1127_n;
  wire g1128_p;
  wire g1128_n;
  wire g1129_p;
  wire g1129_n;
  wire g1130_p;
  wire g1130_n;
  wire g1131_p;
  wire g1131_n;
  wire g1132_p;
  wire g1132_n;
  wire g1133_p;
  wire g1133_n;
  wire g1134_p;
  wire g1134_n;
  wire g1135_p;
  wire g1135_n;
  wire g1136_p;
  wire g1136_n;
  wire g1137_p;
  wire g1137_n;
  wire g1138_p;
  wire g1138_n;
  wire g1139_p;
  wire g1139_n;
  wire g1140_p;
  wire g1140_n;
  wire g1141_p;
  wire g1141_n;
  wire g1142_p;
  wire g1142_n;
  wire g1143_p;
  wire g1143_n;
  wire g1144_p;
  wire g1144_n;
  wire g1145_p;
  wire g1145_n;
  wire g1146_p;
  wire g1146_n;
  wire g1147_p;
  wire g1147_n;
  wire g1148_p;
  wire g1148_n;
  wire g1149_p;
  wire g1149_n;
  wire g1150_p;
  wire g1150_n;
  wire g1151_p;
  wire g1151_n;
  wire g1152_p;
  wire g1152_n;
  wire g1153_p;
  wire g1153_n;
  wire g1154_p;
  wire g1154_n;
  wire g1155_p;
  wire g1155_n;
  wire g1156_p;
  wire g1156_n;
  wire g1157_p;
  wire g1157_n;
  wire g1158_p;
  wire g1158_n;
  wire g1159_p;
  wire g1159_n;
  wire g1160_p;
  wire g1160_n;
  wire g1161_p;
  wire g1161_n;
  wire g1162_p;
  wire g1162_n;
  wire g1163_p;
  wire g1163_n;
  wire g1164_p;
  wire g1164_n;
  wire g1165_p;
  wire g1165_n;
  wire g1166_p;
  wire g1166_n;
  wire g1167_p;
  wire g1167_n;
  wire g1168_p;
  wire g1168_n;
  wire g1169_p;
  wire g1169_n;
  wire g1170_p;
  wire g1170_n;
  wire g1171_p;
  wire g1171_n;
  wire g1172_p;
  wire g1172_n;
  wire g1173_p;
  wire g1173_n;
  wire g1174_p;
  wire g1174_n;
  wire g1175_p;
  wire g1175_n;
  wire g1176_p;
  wire g1176_n;
  wire g1177_p;
  wire g1177_n;
  wire g1178_p;
  wire g1178_n;
  wire g1179_p;
  wire g1179_n;
  wire g1180_p;
  wire g1180_n;
  wire g1181_p;
  wire g1181_n;
  wire g1182_p;
  wire g1182_n;
  wire g1183_p;
  wire g1183_n;
  wire g1184_p;
  wire g1184_n;
  wire g1185_p;
  wire g1185_n;
  wire g1186_p;
  wire g1186_n;
  wire g1187_p;
  wire g1187_n;
  wire g1188_p;
  wire g1188_n;
  wire g1189_p;
  wire g1189_n;
  wire g1190_p;
  wire g1190_n;
  wire g1191_p;
  wire g1191_n;
  wire g1192_p;
  wire g1192_n;
  wire g1193_p;
  wire g1193_n;
  wire g1194_p;
  wire g1194_n;
  wire g1195_p;
  wire g1195_n;
  wire g1196_p;
  wire g1196_n;
  wire g1197_p;
  wire g1197_n;
  wire g1198_p;
  wire g1198_n;
  wire g1199_p;
  wire g1199_n;
  wire g1200_p;
  wire g1200_n;
  wire g1201_p;
  wire g1201_n;
  wire g1202_p;
  wire g1202_n;
  wire g1203_p;
  wire g1203_n;
  wire g1204_p;
  wire g1204_n;
  wire g1205_p;
  wire g1205_n;
  wire g1206_p;
  wire g1206_n;
  wire g1207_p;
  wire g1207_n;
  wire g1208_p;
  wire g1208_n;
  wire g1209_p;
  wire g1209_n;
  wire g1210_p;
  wire g1210_n;
  wire g1211_p;
  wire g1211_n;
  wire g1212_p;
  wire g1212_n;
  wire g1213_p;
  wire g1213_n;
  wire g1214_p;
  wire g1214_n;
  wire g1215_p;
  wire g1215_n;
  wire g1216_p;
  wire g1216_n;
  wire g1217_p;
  wire g1217_n;
  wire g1218_p;
  wire g1218_n;
  wire g1219_p;
  wire g1219_n;
  wire g1220_p;
  wire g1220_n;
  wire g1221_p;
  wire g1221_n;
  wire g1222_p;
  wire g1222_n;
  wire g1223_p;
  wire g1223_n;
  wire g1224_p;
  wire g1224_n;
  wire g1225_p;
  wire g1225_n;
  wire g1226_p;
  wire g1226_n;
  wire g1227_p;
  wire g1227_n;
  wire g1228_p;
  wire g1228_n;
  wire g1229_p;
  wire g1229_n;
  wire g1230_p;
  wire g1230_n;
  wire g1231_p;
  wire g1231_n;
  wire g1232_p;
  wire g1232_n;
  wire g1233_p;
  wire g1233_n;
  wire g1234_p;
  wire g1234_n;
  wire g1235_p;
  wire g1235_n;
  wire g1236_p;
  wire g1236_n;
  wire g1237_p;
  wire g1237_n;
  wire g1238_p;
  wire g1238_n;
  wire g1239_p;
  wire g1239_n;
  wire g1240_p;
  wire g1240_n;
  wire g1241_p;
  wire g1241_n;
  wire g1242_p;
  wire g1242_n;
  wire g1243_p;
  wire g1243_n;
  wire g1244_p;
  wire g1244_n;
  wire g1245_p;
  wire g1245_n;
  wire g1246_p;
  wire g1246_n;
  wire g1247_p;
  wire g1247_n;
  wire g1248_p;
  wire g1248_n;
  wire g1249_p;
  wire g1249_n;
  wire g1250_p;
  wire g1250_n;
  wire g1251_p;
  wire g1251_n;
  wire g1252_p;
  wire g1252_n;
  wire g1253_p;
  wire g1253_n;
  wire g1254_p;
  wire g1254_n;
  wire g1255_p;
  wire g1255_n;
  wire g1256_p;
  wire g1256_n;
  wire g1257_p;
  wire g1257_n;
  wire g1258_p;
  wire g1258_n;
  wire g1259_p;
  wire g1259_n;
  wire g1260_p;
  wire g1260_n;
  wire g1261_p;
  wire g1261_n;
  wire g1262_p;
  wire g1262_n;
  wire g1263_p;
  wire g1263_n;
  wire g1264_p;
  wire g1264_n;
  wire g1265_p;
  wire g1265_n;
  wire g1266_p;
  wire g1266_n;
  wire g1267_p;
  wire g1267_n;
  wire g1268_p;
  wire g1268_n;
  wire g1269_p;
  wire g1269_n;
  wire g1270_p;
  wire g1270_n;
  wire g1271_p;
  wire g1271_n;
  wire g1272_p;
  wire g1272_n;
  wire g1273_p;
  wire g1273_n;
  wire g1274_p;
  wire g1274_n;
  wire g1275_p;
  wire g1275_n;
  wire g1276_p;
  wire g1276_n;
  wire g1277_p;
  wire g1277_n;
  wire g1278_p;
  wire g1278_n;
  wire g1279_p;
  wire g1279_n;
  wire g1280_p;
  wire g1280_n;
  wire g1281_p;
  wire g1281_n;
  wire g1282_p;
  wire g1282_n;
  wire g1283_p;
  wire g1283_n;
  wire g1284_p;
  wire g1284_n;
  wire g1285_p;
  wire g1285_n;
  wire g1286_p;
  wire g1286_n;
  wire g1287_p;
  wire g1287_n;
  wire g1288_p;
  wire g1288_n;
  wire g1289_p;
  wire g1289_n;
  wire g1290_p;
  wire g1290_n;
  wire g1291_p;
  wire g1291_n;
  wire g1292_p;
  wire g1292_n;
  wire g1293_p;
  wire g1293_n;
  wire g1294_p;
  wire g1294_n;
  wire g1295_p;
  wire g1295_n;
  wire g1296_p;
  wire g1296_n;
  wire g1297_p;
  wire g1297_n;
  wire g1298_p;
  wire g1298_n;
  wire g1299_p;
  wire g1299_n;
  wire g1300_p;
  wire g1300_n;
  wire g1301_p;
  wire g1301_n;
  wire g1302_p;
  wire g1302_n;
  wire g1303_p;
  wire g1303_n;
  wire g1304_p;
  wire g1304_n;
  wire g1305_p;
  wire g1305_n;
  wire g1306_p;
  wire g1306_n;
  wire g1307_p;
  wire g1307_n;
  wire g1308_p;
  wire g1308_n;
  wire g1309_p;
  wire g1309_n;
  wire g1310_p;
  wire g1310_n;
  wire g1311_p;
  wire g1311_n;
  wire g1312_p;
  wire g1312_n;
  wire g1313_p;
  wire g1313_n;
  wire g1314_p;
  wire g1314_n;
  wire g1315_p;
  wire g1315_n;
  wire g1316_p;
  wire g1316_n;
  wire g1317_p;
  wire g1317_n;
  wire g1318_p;
  wire g1318_n;
  wire g1319_p;
  wire g1319_n;
  wire g1320_p;
  wire g1320_n;
  wire g1321_p;
  wire g1321_n;
  wire g1322_p;
  wire g1322_n;
  wire g1323_p;
  wire g1323_n;
  wire g1324_p;
  wire g1324_n;
  wire g1325_p;
  wire g1325_n;
  wire g1326_p;
  wire g1326_n;
  wire g1327_p;
  wire g1327_n;
  wire g1328_p;
  wire g1328_n;
  wire g1329_p;
  wire g1329_n;
  wire g1330_p;
  wire g1330_n;
  wire g1331_p;
  wire g1331_n;
  wire g1332_p;
  wire g1332_n;
  wire g1333_p;
  wire g1333_n;
  wire g1334_p;
  wire g1334_n;
  wire g1335_p;
  wire g1335_n;
  wire g1336_p;
  wire g1336_n;
  wire g1337_p;
  wire g1337_n;
  wire g1338_p;
  wire g1338_n;
  wire g1339_p;
  wire g1339_n;
  wire g1340_p;
  wire g1340_n;
  wire g1341_p;
  wire g1341_n;
  wire g1342_p;
  wire g1342_n;
  wire g1343_p;
  wire g1343_n;
  wire g1344_p;
  wire g1344_n;
  wire g1345_p;
  wire g1345_n;
  wire g1346_p;
  wire g1346_n;
  wire g1347_p;
  wire g1347_n;
  wire g1348_p;
  wire g1348_n;
  wire g1349_p;
  wire g1349_n;
  wire g1350_p;
  wire g1350_n;
  wire g1351_p;
  wire g1351_n;
  wire g1352_p;
  wire g1352_n;
  wire g1353_p;
  wire g1353_n;
  wire g1354_p;
  wire g1354_n;
  wire g1355_p;
  wire g1355_n;
  wire g1356_p;
  wire g1356_n;
  wire g1357_p;
  wire g1357_n;
  wire g1358_p;
  wire g1358_n;
  wire g1359_p;
  wire g1359_n;
  wire g1360_p;
  wire g1360_n;
  wire g1361_p;
  wire g1361_n;
  wire g1362_p;
  wire g1362_n;
  wire g1363_p;
  wire g1363_n;
  wire g1364_p;
  wire g1364_n;
  wire g1365_p;
  wire g1365_n;
  wire g1366_p;
  wire g1366_n;
  wire g1367_p;
  wire g1367_n;
  wire g1368_p;
  wire g1368_n;
  wire g1369_p;
  wire g1369_n;
  wire g1370_p;
  wire g1370_n;
  wire g1371_p;
  wire g1371_n;
  wire g1372_p;
  wire g1372_n;
  wire g1373_p;
  wire g1373_n;
  wire g1374_p;
  wire g1374_n;
  wire g1375_p;
  wire g1375_n;
  wire g1376_p;
  wire g1376_n;
  wire g1377_p;
  wire g1377_n;
  wire g1378_p;
  wire g1378_n;
  wire g1379_p;
  wire g1379_n;
  wire g1380_p;
  wire g1380_n;
  wire g1381_p;
  wire g1381_n;
  wire g1382_p;
  wire g1382_n;
  wire g1383_p;
  wire g1383_n;
  wire g1384_p;
  wire g1384_n;
  wire g1385_p;
  wire g1385_n;
  wire g1386_p;
  wire g1386_n;
  wire g1387_p;
  wire g1387_n;
  wire g1388_p;
  wire g1388_n;
  wire g1389_p;
  wire g1389_n;
  wire g1390_p;
  wire g1390_n;
  wire g1391_p;
  wire g1391_n;
  wire g1392_p;
  wire g1392_n;
  wire g1393_p;
  wire g1393_n;
  wire g1394_p;
  wire g1394_n;
  wire g1395_p;
  wire g1395_n;
  wire g1396_p;
  wire g1396_n;
  wire g1397_p;
  wire g1397_n;
  wire g1398_p;
  wire g1398_n;
  wire g1399_p;
  wire g1399_n;
  wire g1400_p;
  wire g1400_n;
  wire g1401_p;
  wire g1401_n;
  wire g1402_p;
  wire g1402_n;
  wire g1403_p;
  wire g1403_n;
  wire g1404_p;
  wire g1404_n;
  wire g1405_p;
  wire g1405_n;
  wire g1406_p;
  wire g1406_n;
  wire g1407_p;
  wire g1407_n;
  wire g1408_p;
  wire g1408_n;
  wire g1409_p;
  wire g1409_n;
  wire g1410_p;
  wire g1410_n;
  wire g1411_p;
  wire g1411_n;
  wire g1412_p;
  wire g1412_n;
  wire g1413_p;
  wire g1413_n;
  wire g1414_p;
  wire g1414_n;
  wire g1415_p;
  wire g1415_n;
  wire g1416_p;
  wire g1416_n;
  wire g1417_p;
  wire g1417_n;
  wire g1418_p;
  wire g1418_n;
  wire g1419_p;
  wire g1419_n;
  wire g1420_p;
  wire g1420_n;
  wire g1421_p;
  wire g1421_n;
  wire g1422_p;
  wire g1422_n;
  wire g1423_p;
  wire g1423_n;
  wire g1424_p;
  wire g1424_n;
  wire g1425_p;
  wire g1425_n;
  wire g1426_p;
  wire g1426_n;
  wire g1427_p;
  wire g1427_n;
  wire g1428_p;
  wire g1428_n;
  wire g1429_p;
  wire g1429_n;
  wire g1430_p;
  wire g1430_n;
  wire g1431_p;
  wire g1431_n;
  wire g1432_p;
  wire g1432_n;
  wire g1433_p;
  wire g1433_n;
  wire g1434_p;
  wire g1434_n;
  wire g1435_p;
  wire g1435_n;
  wire g1436_p;
  wire g1436_n;
  wire g1437_p;
  wire g1437_n;
  wire g1438_p;
  wire g1438_n;
  wire g1439_p;
  wire g1439_n;
  wire g1440_p;
  wire g1440_n;
  wire g1441_p;
  wire g1441_n;
  wire g1442_p;
  wire g1442_n;
  wire g1443_p;
  wire g1443_n;
  wire g1444_p;
  wire g1444_n;
  wire g1445_p;
  wire g1445_n;
  wire g1446_p;
  wire g1446_n;
  wire g1447_p;
  wire g1447_n;
  wire g1448_p;
  wire g1448_n;
  wire g1449_p;
  wire g1449_n;
  wire g1450_p;
  wire g1450_n;
  wire g1451_p;
  wire g1451_n;
  wire g1452_p;
  wire g1452_n;
  wire g1453_p;
  wire g1453_n;
  wire g1454_p;
  wire g1454_n;
  wire g1455_p;
  wire g1455_n;
  wire g1456_p;
  wire g1456_n;
  wire g1457_p;
  wire g1457_n;
  wire g1458_p;
  wire g1458_n;
  wire g1459_p;
  wire g1459_n;
  wire g1460_p;
  wire g1460_n;
  wire g1461_p;
  wire g1461_n;
  wire g1462_p;
  wire g1462_n;
  wire g1463_p;
  wire g1463_n;
  wire g1464_p;
  wire g1464_n;
  wire g1465_p;
  wire g1465_n;
  wire g1466_p;
  wire g1466_n;
  wire g1467_p;
  wire g1467_n;
  wire g1468_p;
  wire g1468_n;
  wire g1469_p;
  wire g1469_n;
  wire g1470_p;
  wire g1470_n;
  wire g1471_p;
  wire g1471_n;
  wire g1472_p;
  wire g1472_n;
  wire g1473_p;
  wire g1473_n;
  wire g1474_p;
  wire g1474_n;
  wire g1475_p;
  wire g1475_n;
  wire g1476_p;
  wire g1476_n;
  wire g1477_p;
  wire g1477_n;
  wire g1478_p;
  wire g1478_n;
  wire g1479_p;
  wire g1479_n;
  wire g1480_p;
  wire g1480_n;
  wire g1481_p;
  wire g1481_n;
  wire g1482_p;
  wire g1482_n;
  wire g1483_p;
  wire g1483_n;
  wire g1484_p;
  wire g1484_n;
  wire g1485_p;
  wire g1485_n;
  wire g1486_p;
  wire g1486_n;
  wire g1487_p;
  wire g1487_n;
  wire g1488_p;
  wire g1488_n;
  wire g1489_p;
  wire g1489_n;
  wire g1490_p;
  wire g1490_n;
  wire g1491_p;
  wire g1491_n;
  wire g1492_p;
  wire g1492_n;
  wire g1493_p;
  wire g1493_n;
  wire g1494_p;
  wire g1494_n;
  wire g1495_p;
  wire g1495_n;
  wire g1496_p;
  wire g1496_n;
  wire g1497_p;
  wire g1497_n;
  wire g1498_p;
  wire g1498_n;
  wire g1499_p;
  wire g1499_n;
  wire g1500_p;
  wire g1500_n;
  wire g1501_p;
  wire g1501_n;
  wire g1502_p;
  wire g1502_n;
  wire g1503_p;
  wire g1503_n;
  wire g1504_p;
  wire g1504_n;
  wire g1505_p;
  wire g1505_n;
  wire g1506_p;
  wire g1506_n;
  wire g1507_p;
  wire g1507_n;
  wire g1508_p;
  wire g1508_n;
  wire g1509_p;
  wire g1509_n;
  wire g1510_p;
  wire g1510_n;
  wire g1511_p;
  wire g1511_n;
  wire g1512_p;
  wire g1512_n;
  wire g1513_p;
  wire g1513_n;
  wire g1514_p;
  wire g1514_n;
  wire g1515_p;
  wire g1515_n;
  wire g1516_p;
  wire g1516_n;
  wire g1517_p;
  wire g1517_n;
  wire g1518_p;
  wire g1518_n;
  wire g1519_p;
  wire g1519_n;
  wire g1520_p;
  wire g1520_n;
  wire g1521_p;
  wire g1521_n;
  wire g1522_p;
  wire g1522_n;
  wire g1523_p;
  wire g1523_n;
  wire g1524_p;
  wire g1524_n;
  wire g1525_p;
  wire g1525_n;
  wire g1526_p;
  wire g1526_n;
  wire g1527_p;
  wire g1527_n;
  wire g1528_p;
  wire g1528_n;
  wire g1529_p;
  wire g1529_n;
  wire g1530_p;
  wire g1530_n;
  wire g1531_p;
  wire g1531_n;
  wire g1532_p;
  wire g1532_n;
  wire g1533_p;
  wire g1533_n;
  wire g1534_p;
  wire g1534_n;
  wire g1535_p;
  wire g1535_n;
  wire g1536_p;
  wire g1536_n;
  wire g1537_p;
  wire g1537_n;
  wire g1538_p;
  wire g1538_n;
  wire g1539_p;
  wire g1539_n;
  wire g1540_p;
  wire g1540_n;
  wire g1541_p;
  wire g1541_n;
  wire g1542_p;
  wire g1542_n;
  wire g1543_p;
  wire g1543_n;
  wire g1544_p;
  wire g1544_n;
  wire g1545_p;
  wire g1545_n;
  wire g1546_p;
  wire g1546_n;
  wire g1547_p;
  wire g1547_n;
  wire g1548_p;
  wire g1548_n;
  wire g1549_p;
  wire g1549_n;
  wire g1550_p;
  wire g1550_n;
  wire g1551_p;
  wire g1551_n;
  wire g1552_p;
  wire g1552_n;
  wire g1553_p;
  wire g1553_n;
  wire g1554_p;
  wire g1554_n;
  wire g1555_p;
  wire g1555_n;
  wire g1556_p;
  wire g1556_n;
  wire g1557_p;
  wire g1557_n;
  wire g1558_p;
  wire g1558_n;
  wire g1559_p;
  wire g1559_n;
  wire g1560_p;
  wire g1560_n;
  wire g1561_p;
  wire g1561_n;
  wire g1562_p;
  wire g1562_n;
  wire g1563_p;
  wire g1563_n;
  wire g1564_p;
  wire g1564_n;
  wire g1565_p;
  wire g1565_n;
  wire g1566_p;
  wire g1566_n;
  wire g1567_p;
  wire g1567_n;
  wire g1568_p;
  wire g1568_n;
  wire g1569_p;
  wire g1569_n;
  wire g1570_p;
  wire g1570_n;
  wire g1571_p;
  wire g1571_n;
  wire g1572_p;
  wire g1572_n;
  wire g1573_p;
  wire g1573_n;
  wire g1574_p;
  wire g1574_n;
  wire g1575_p;
  wire g1575_n;
  wire g1576_p;
  wire g1576_n;
  wire g1577_p;
  wire g1577_n;
  wire g1578_p;
  wire g1578_n;
  wire g1579_p;
  wire g1579_n;
  wire g1580_p;
  wire g1580_n;
  wire g1581_p;
  wire g1581_n;
  wire g1582_p;
  wire g1582_n;
  wire g1583_p;
  wire g1583_n;
  wire g1584_p;
  wire g1584_n;
  wire g1585_p;
  wire g1585_n;
  wire g1586_p;
  wire g1586_n;
  wire g1587_p;
  wire g1587_n;
  wire g1588_p;
  wire g1588_n;
  wire g1589_p;
  wire g1589_n;
  wire g1590_p;
  wire g1590_n;
  wire g1591_p;
  wire g1591_n;
  wire g1592_p;
  wire g1592_n;
  wire g1593_p;
  wire g1593_n;
  wire g1594_p;
  wire g1594_n;
  wire g1595_p;
  wire g1595_n;
  wire g1596_p;
  wire g1596_n;
  wire g1597_p;
  wire g1597_n;
  wire g1598_p;
  wire g1598_n;
  wire g1599_p;
  wire g1599_n;
  wire g1600_p;
  wire g1600_n;
  wire g1601_p;
  wire g1601_n;
  wire g1602_p;
  wire g1602_n;
  wire g1603_p;
  wire g1603_n;
  wire g1604_p;
  wire g1604_n;
  wire g1605_p;
  wire g1605_n;
  wire g1606_p;
  wire g1606_n;
  wire g1607_p;
  wire g1607_n;
  wire g1608_p;
  wire g1608_n;
  wire g1609_p;
  wire g1609_n;
  wire g1610_p;
  wire g1610_n;
  wire g1611_p;
  wire g1611_n;
  wire g1612_p;
  wire g1612_n;
  wire g1613_p;
  wire g1613_n;
  wire g1614_p;
  wire g1614_n;
  wire g1615_p;
  wire g1615_n;
  wire g1616_p;
  wire g1616_n;
  wire g1617_p;
  wire g1617_n;
  wire g1618_p;
  wire g1618_n;
  wire g1619_p;
  wire g1619_n;
  wire g1620_p;
  wire g1620_n;
  wire g1621_p;
  wire g1621_n;
  wire g1622_p;
  wire g1622_n;
  wire g1623_p;
  wire g1623_n;
  wire g1624_p;
  wire g1624_n;
  wire g1625_p;
  wire g1625_n;
  wire g1626_p;
  wire g1626_n;
  wire g1627_p;
  wire g1627_n;
  wire g1628_p;
  wire g1628_n;
  wire g1629_p;
  wire g1629_n;
  wire g1630_p;
  wire g1630_n;
  wire g1631_p;
  wire g1631_n;
  wire g1632_p;
  wire g1632_n;
  wire g1633_p;
  wire g1633_n;
  wire g1634_p;
  wire g1634_n;
  wire g1635_p;
  wire g1635_n;
  wire g1636_p;
  wire g1636_n;
  wire g1637_p;
  wire g1637_n;
  wire g1638_p;
  wire g1638_n;
  wire g1639_p;
  wire g1639_n;
  wire g1640_p;
  wire g1640_n;
  wire g1641_p;
  wire g1641_n;
  wire g1642_p;
  wire g1642_n;
  wire g1643_p;
  wire g1643_n;
  wire g1644_p;
  wire g1644_n;
  wire g1645_p;
  wire g1645_n;
  wire g1646_p;
  wire g1646_n;
  wire g1647_p;
  wire g1647_n;
  wire g1648_p;
  wire g1648_n;
  wire g1649_p;
  wire g1649_n;
  wire g1650_p;
  wire g1650_n;
  wire g1651_p;
  wire g1651_n;
  wire g1652_p;
  wire g1652_n;
  wire g1653_p;
  wire g1653_n;
  wire g1654_p;
  wire g1654_n;
  wire g1655_p;
  wire g1655_n;
  wire g1656_p;
  wire g1656_n;
  wire g1657_p;
  wire g1657_n;
  wire g1658_p;
  wire g1658_n;
  wire g1659_p;
  wire g1659_n;
  wire g1660_p;
  wire g1660_n;
  wire g1661_p;
  wire g1661_n;
  wire g1662_p;
  wire g1662_n;
  wire g1663_p;
  wire g1663_n;
  wire g1664_p;
  wire g1664_n;
  wire g1665_p;
  wire g1665_n;
  wire g1666_p;
  wire g1666_n;
  wire g1667_p;
  wire g1667_n;
  wire g1668_p;
  wire g1668_n;
  wire g1669_p;
  wire g1669_n;
  wire g1670_p;
  wire g1670_n;
  wire g1671_p;
  wire g1671_n;
  wire g1672_p;
  wire g1672_n;
  wire g1673_p;
  wire g1673_n;
  wire g1674_p;
  wire g1674_n;
  wire g1675_p;
  wire g1675_n;
  wire g1676_p;
  wire g1676_n;
  wire g1677_p;
  wire g1677_n;
  wire g1678_p;
  wire g1678_n;
  wire g1679_p;
  wire g1679_n;
  wire g1680_p;
  wire g1680_n;
  wire g1681_p;
  wire g1681_n;
  wire g1682_p;
  wire g1682_n;
  wire g1683_p;
  wire g1683_n;
  wire g1684_p;
  wire g1684_n;
  wire g1685_p;
  wire g1685_n;
  wire g1686_p;
  wire g1686_n;
  wire g1687_p;
  wire g1687_n;
  wire g1688_p;
  wire g1688_n;
  wire g1689_p;
  wire g1689_n;
  wire g1690_p;
  wire g1690_n;
  wire g1691_p;
  wire g1691_n;
  wire g1692_p;
  wire g1692_n;
  wire g1693_p;
  wire g1693_n;
  wire g1694_p;
  wire g1694_n;
  wire g1695_p;
  wire g1695_n;
  wire g1696_p;
  wire g1696_n;
  wire g1697_p;
  wire g1697_n;
  wire g1698_p;
  wire g1698_n;
  wire g1699_p;
  wire g1699_n;
  wire g1700_p;
  wire g1700_n;
  wire g1701_p;
  wire g1701_n;
  wire g1702_p;
  wire g1702_n;
  wire g1703_p;
  wire g1703_n;
  wire g1704_p;
  wire g1704_n;
  wire g1705_p;
  wire g1705_n;
  wire g1706_p;
  wire g1706_n;
  wire g1707_p;
  wire g1707_n;
  wire g1708_p;
  wire g1708_n;
  wire g1709_p;
  wire g1709_n;
  wire g1710_p;
  wire g1710_n;
  wire g1711_p;
  wire g1711_n;
  wire g1712_p;
  wire g1712_n;
  wire g1713_p;
  wire g1713_n;
  wire g1714_p;
  wire g1714_n;
  wire g1715_p;
  wire g1715_n;
  wire g1716_p;
  wire g1716_n;
  wire g1717_p;
  wire g1717_n;
  wire g1718_p;
  wire g1718_n;
  wire g1719_p;
  wire g1719_n;
  wire g1720_p;
  wire g1720_n;
  wire g1721_p;
  wire g1721_n;
  wire g1722_p;
  wire g1722_n;
  wire g1723_p;
  wire g1723_n;
  wire g1724_p;
  wire g1724_n;
  wire g1725_p;
  wire g1725_n;
  wire g1726_p;
  wire g1726_n;
  wire g1727_p;
  wire g1727_n;
  wire g1728_p;
  wire g1728_n;
  wire g1729_p;
  wire g1729_n;
  wire g1730_p;
  wire g1730_n;
  wire g1731_p;
  wire g1731_n;
  wire g1732_p;
  wire g1732_n;
  wire g1733_p;
  wire g1733_n;
  wire g1734_p;
  wire g1734_n;
  wire g1735_p;
  wire g1735_n;
  wire g1736_p;
  wire g1736_n;
  wire g1737_p;
  wire g1737_n;
  wire g1738_p;
  wire g1738_n;
  wire g1739_p;
  wire g1739_n;
  wire g1740_p;
  wire g1740_n;
  wire g1741_p;
  wire g1741_n;
  wire g1742_p;
  wire g1742_n;
  wire g1743_p;
  wire g1743_n;
  wire g1744_p;
  wire g1744_n;
  wire g1745_p;
  wire g1745_n;
  wire g1746_p;
  wire g1746_n;
  wire g1747_p;
  wire g1747_n;
  wire g1748_p;
  wire g1748_n;
  wire g1749_p;
  wire g1749_n;
  wire g1750_p;
  wire g1750_n;
  wire g1751_p;
  wire g1751_n;
  wire g1752_p;
  wire g1752_n;
  wire g1753_p;
  wire g1753_n;
  wire g1754_p;
  wire g1754_n;
  wire g1755_p;
  wire g1755_n;
  wire g1756_p;
  wire g1756_n;
  wire g1757_p;
  wire g1757_n;
  wire g1758_p;
  wire g1758_n;
  wire g1759_p;
  wire g1759_n;
  wire g1760_p;
  wire g1760_n;
  wire g1761_p;
  wire g1761_n;
  wire g1762_p;
  wire g1762_n;
  wire g1763_p;
  wire g1763_n;
  wire g1764_p;
  wire g1764_n;
  wire g1765_p;
  wire g1765_n;
  wire g1766_p;
  wire g1766_n;
  wire g1767_p;
  wire g1767_n;
  wire g1768_p;
  wire g1768_n;
  wire g1769_p;
  wire g1769_n;
  wire g1770_p;
  wire g1770_n;
  wire g1771_p;
  wire g1771_n;
  wire g1772_p;
  wire g1772_n;
  wire g1773_p;
  wire g1773_n;
  wire g1774_p;
  wire g1774_n;
  wire g1775_p;
  wire g1775_n;
  wire g1776_p;
  wire g1776_n;
  wire g1777_p;
  wire g1777_n;
  wire g1778_p;
  wire g1778_n;
  wire g1779_p;
  wire g1779_n;
  wire g1780_p;
  wire g1780_n;
  wire g1781_p;
  wire g1781_n;
  wire g1782_p;
  wire g1782_n;
  wire g1783_p;
  wire g1783_n;
  wire g1784_p;
  wire g1784_n;
  wire g1785_p;
  wire g1785_n;
  wire g1786_p;
  wire g1786_n;
  wire g1787_p;
  wire g1787_n;
  wire g1788_p;
  wire g1788_n;
  wire g1789_p;
  wire g1789_n;
  wire g1790_p;
  wire g1790_n;
  wire g1791_p;
  wire g1791_n;
  wire g1792_p;
  wire g1792_n;
  wire g1793_p;
  wire g1793_n;
  wire g1794_p;
  wire g1794_n;
  wire g1795_p;
  wire g1795_n;
  wire g1796_p;
  wire g1796_n;
  wire g1797_p;
  wire g1797_n;
  wire g1798_p;
  wire g1798_n;
  wire g1799_p;
  wire g1799_n;
  wire g1800_p;
  wire g1800_n;
  wire g1801_p;
  wire g1801_n;
  wire g1802_p;
  wire g1802_n;
  wire g1803_p;
  wire g1803_n;
  wire g1804_p;
  wire g1804_n;
  wire g1805_p;
  wire g1805_n;
  wire g1806_p;
  wire g1806_n;
  wire g1807_p;
  wire g1807_n;
  wire g1808_p;
  wire g1808_n;
  wire g1809_p;
  wire g1809_n;
  wire g1810_p;
  wire g1810_n;
  wire g1811_p;
  wire g1811_n;
  wire g1812_p;
  wire g1812_n;
  wire g1813_p;
  wire g1813_n;
  wire g1814_p;
  wire g1814_n;
  wire g1815_p;
  wire g1815_n;
  wire g1816_p;
  wire g1816_n;
  wire g1817_p;
  wire g1817_n;
  wire g1818_p;
  wire g1818_n;
  wire g1819_p;
  wire g1819_n;
  wire g1820_p;
  wire g1820_n;
  wire g1821_p;
  wire g1821_n;
  wire g1822_p;
  wire g1822_n;
  wire g1823_p;
  wire g1823_n;
  wire g1824_p;
  wire g1824_n;
  wire g1825_p;
  wire g1825_n;
  wire g1826_p;
  wire g1826_n;
  wire g1827_p;
  wire g1827_n;
  wire g1828_p;
  wire g1828_n;
  wire g1829_p;
  wire g1829_n;
  wire g1830_p;
  wire g1830_n;
  wire g1831_p;
  wire g1831_n;
  wire g1832_p;
  wire g1832_n;
  wire g1833_p;
  wire g1833_n;
  wire g1834_p;
  wire g1834_n;
  wire g1835_p;
  wire g1835_n;
  wire g1836_p;
  wire g1836_n;
  wire g1837_p;
  wire g1837_n;
  wire g1838_p;
  wire g1838_n;
  wire g1839_p;
  wire g1839_n;
  wire g1840_p;
  wire g1840_n;
  wire g1841_p;
  wire g1841_n;
  wire g1842_p;
  wire g1842_n;
  wire g1843_p;
  wire g1843_n;
  wire g1844_p;
  wire g1844_n;
  wire g1845_p;
  wire g1845_n;
  wire g1846_p;
  wire g1846_n;
  wire g1847_p;
  wire g1847_n;
  wire g1848_p;
  wire g1848_n;
  wire g1849_p;
  wire g1849_n;
  wire g1850_p;
  wire g1850_n;
  wire g1851_p;
  wire g1851_n;
  wire g1852_p;
  wire g1852_n;
  wire g1853_p;
  wire g1853_n;
  wire g1854_p;
  wire g1854_n;
  wire g1855_p;
  wire g1855_n;
  wire g1856_p;
  wire g1856_n;
  wire g1857_p;
  wire g1857_n;
  wire g1858_p;
  wire g1858_n;
  wire g1859_p;
  wire g1859_n;
  wire g1860_p;
  wire g1860_n;
  wire g1861_p;
  wire g1861_n;
  wire g1862_p;
  wire g1862_n;
  wire g1863_p;
  wire g1863_n;
  wire g1864_p;
  wire g1864_n;
  wire g1865_p;
  wire g1865_n;
  wire g1866_p;
  wire g1866_n;
  wire g1867_p;
  wire g1867_n;
  wire g1868_p;
  wire g1868_n;
  wire g1869_p;
  wire g1869_n;
  wire g1870_p;
  wire g1870_n;
  wire g1871_p;
  wire g1871_n;
  wire g1872_p;
  wire g1872_n;
  wire g1873_p;
  wire g1873_n;
  wire g1874_p;
  wire g1874_n;
  wire g1875_p;
  wire g1875_n;
  wire g1876_p;
  wire g1876_n;
  wire g1877_p;
  wire g1877_n;
  wire g1878_p;
  wire g1878_n;
  wire g1879_p;
  wire g1879_n;
  wire g1880_p;
  wire g1880_n;
  wire g1881_p;
  wire g1881_n;
  wire g1882_p;
  wire g1882_n;
  wire g1883_p;
  wire g1883_n;
  wire g1884_p;
  wire g1884_n;
  wire g1885_p;
  wire g1885_n;
  wire g1886_p;
  wire g1886_n;
  wire g1887_p;
  wire g1887_n;
  wire g1888_p;
  wire g1888_n;
  wire g1889_p;
  wire g1889_n;
  wire g1890_p;
  wire g1890_n;
  wire g1891_p;
  wire g1891_n;
  wire g1892_p;
  wire g1892_n;
  wire g1893_p;
  wire g1893_n;
  wire g1894_p;
  wire g1894_n;
  wire g1895_p;
  wire g1895_n;
  wire g1896_p;
  wire g1896_n;
  wire g1897_p;
  wire g1897_n;
  wire g1898_p;
  wire g1898_n;
  wire g1899_p;
  wire g1899_n;
  wire g1900_p;
  wire g1900_n;
  wire g1901_p;
  wire g1901_n;
  wire g1902_p;
  wire g1902_n;
  wire g1903_p;
  wire g1903_n;
  wire g1904_p;
  wire g1904_n;
  wire g1905_p;
  wire g1905_n;
  wire g1906_p;
  wire g1906_n;
  wire g1907_p;
  wire g1907_n;
  wire g1908_p;
  wire g1908_n;
  wire g1909_p;
  wire g1909_n;
  wire g1910_p;
  wire g1910_n;
  wire g1911_p;
  wire g1911_n;
  wire g1912_p;
  wire g1912_n;
  wire g1913_p;
  wire g1913_n;
  wire g1914_p;
  wire g1914_n;
  wire g1915_p;
  wire g1915_n;
  wire g1916_p;
  wire g1916_n;
  wire g1917_p;
  wire g1917_n;
  wire g1918_p;
  wire g1918_n;
  wire g1919_p;
  wire g1919_n;
  wire g1920_p;
  wire g1920_n;
  wire g1921_p;
  wire g1921_n;
  wire g1922_p;
  wire g1922_n;
  wire g1923_p;
  wire g1923_n;
  wire g1924_p;
  wire g1924_n;
  wire g1925_p;
  wire g1925_n;
  wire g1926_p;
  wire g1926_n;
  wire g1927_p;
  wire g1927_n;
  wire g1928_p;
  wire g1928_n;
  wire g1929_p;
  wire g1929_n;
  wire g1930_p;
  wire g1930_n;
  wire g1931_p;
  wire g1931_n;
  wire g1932_p;
  wire g1932_n;
  wire g1933_p;
  wire g1933_n;
  wire g1934_p;
  wire g1934_n;
  wire g1935_p;
  wire g1935_n;
  wire g1936_p;
  wire g1936_n;
  wire g1937_p;
  wire g1937_n;
  wire g1938_p;
  wire g1938_n;
  wire g1939_p;
  wire g1939_n;
  wire g1940_p;
  wire g1940_n;
  wire g1941_p;
  wire g1941_n;
  wire g1942_p;
  wire g1942_n;
  wire g1943_p;
  wire g1943_n;
  wire g1944_p;
  wire g1944_n;
  wire g1945_p;
  wire g1945_n;
  wire g1946_p;
  wire g1946_n;
  wire g1947_p;
  wire g1947_n;
  wire g1948_p;
  wire g1948_n;
  wire g1949_p;
  wire g1949_n;
  wire g1950_p;
  wire g1950_n;
  wire g1951_p;
  wire g1951_n;
  wire g1952_p;
  wire g1952_n;
  wire g1953_p;
  wire g1953_n;
  wire g1954_p;
  wire g1954_n;
  wire g1955_p;
  wire g1955_n;
  wire g1956_p;
  wire g1956_n;
  wire g1957_p;
  wire g1957_n;
  wire g1958_p;
  wire g1958_n;
  wire g1959_p;
  wire g1959_n;
  wire g1960_p;
  wire g1960_n;
  wire g1961_p;
  wire g1961_n;
  wire g1962_p;
  wire g1962_n;
  wire g1963_p;
  wire g1963_n;
  wire g1964_p;
  wire g1964_n;
  wire g1965_p;
  wire g1965_n;
  wire g1966_p;
  wire g1966_n;
  wire g1967_p;
  wire g1967_n;
  wire g1968_p;
  wire g1968_n;
  wire g1969_p;
  wire g1969_n;
  wire g1970_p;
  wire g1970_n;
  wire g1971_p;
  wire g1971_n;
  wire g1972_p;
  wire g1972_n;
  wire g1973_p;
  wire g1973_n;
  wire g1974_p;
  wire g1974_n;
  wire g1975_p;
  wire g1975_n;
  wire g1976_p;
  wire g1976_n;
  wire g1977_p;
  wire g1977_n;
  wire g1978_p;
  wire g1978_n;
  wire g1979_p;
  wire g1979_n;
  wire g1980_p;
  wire g1980_n;
  wire g1981_p;
  wire g1981_n;
  wire g1982_p;
  wire g1982_n;
  wire g1983_p;
  wire g1983_n;
  wire g1984_p;
  wire g1984_n;
  wire g1985_p;
  wire g1985_n;
  wire g1986_p;
  wire g1986_n;
  wire g1987_p;
  wire g1987_n;
  wire g1988_p;
  wire g1988_n;
  wire g1989_p;
  wire g1989_n;
  wire g1990_p;
  wire g1990_n;
  wire g1991_p;
  wire g1991_n;
  wire g1992_p;
  wire g1992_n;
  wire g1993_p;
  wire g1993_n;
  wire g1994_p;
  wire g1994_n;
  wire g1995_p;
  wire g1995_n;
  wire g1996_p;
  wire g1996_n;
  wire g1997_p;
  wire g1997_n;
  wire g1998_p;
  wire g1998_n;
  wire g1999_p;
  wire g1999_n;
  wire g2000_p;
  wire g2000_n;
  wire g2001_p;
  wire g2001_n;
  wire g2002_p;
  wire g2002_n;
  wire g2003_p;
  wire g2003_n;
  wire g2004_p;
  wire g2004_n;
  wire g2005_p;
  wire g2005_n;
  wire g2006_p;
  wire g2006_n;
  wire g2007_p;
  wire g2007_n;
  wire g2008_p;
  wire g2008_n;
  wire g2009_p;
  wire g2009_n;
  wire g2010_p;
  wire g2010_n;
  wire g2011_p;
  wire g2011_n;
  wire g2012_p;
  wire g2012_n;
  wire g2013_p;
  wire g2013_n;
  wire g2014_p;
  wire g2014_n;
  wire g2015_p;
  wire g2015_n;
  wire g2016_p;
  wire g2016_n;
  wire g2017_p;
  wire g2017_n;
  wire g2018_p;
  wire g2018_n;
  wire g2019_p;
  wire g2019_n;
  wire g2020_p;
  wire g2020_n;
  wire g2021_p;
  wire g2021_n;
  wire g2022_p;
  wire g2022_n;
  wire g2023_p;
  wire g2023_n;
  wire g2024_p;
  wire g2024_n;
  wire g2025_p;
  wire g2025_n;
  wire g2026_p;
  wire g2026_n;
  wire g2027_p;
  wire g2027_n;
  wire g2028_p;
  wire g2028_n;
  wire g2029_p;
  wire g2029_n;
  wire g2030_p;
  wire g2030_n;
  wire g2031_p;
  wire g2031_n;
  wire g2032_p;
  wire g2032_n;
  wire g2033_p;
  wire g2033_n;
  wire g2034_p;
  wire g2034_n;
  wire g2035_p;
  wire g2035_n;
  wire g2036_p;
  wire g2036_n;
  wire g2037_p;
  wire g2037_n;
  wire g2038_p;
  wire g2038_n;
  wire g2039_p;
  wire g2039_n;
  wire g2040_p;
  wire g2040_n;
  wire g2041_p;
  wire g2041_n;
  wire g2042_p;
  wire g2042_n;
  wire g2043_p;
  wire g2043_n;
  wire g2044_p;
  wire g2044_n;
  wire g2045_p;
  wire g2045_n;
  wire g2046_p;
  wire g2046_n;
  wire g2047_p;
  wire g2047_n;
  wire g2048_p;
  wire g2048_n;
  wire g2049_p;
  wire g2049_n;
  wire g2050_p;
  wire g2050_n;
  wire g2051_p;
  wire g2051_n;
  wire g2052_p;
  wire g2052_n;
  wire g2053_p;
  wire g2053_n;
  wire g2054_p;
  wire g2054_n;
  wire g2055_p;
  wire g2055_n;
  wire g2056_p;
  wire g2056_n;
  wire g2057_p;
  wire g2057_n;
  wire g2058_p;
  wire g2058_n;
  wire g2059_p;
  wire g2059_n;
  wire g2060_p;
  wire g2060_n;
  wire g2061_p;
  wire g2061_n;
  wire g2062_p;
  wire g2062_n;
  wire g2063_p;
  wire g2063_n;
  wire g2064_p;
  wire g2064_n;
  wire g2065_p;
  wire g2065_n;
  wire g2066_p;
  wire g2066_n;
  wire g2067_p;
  wire g2067_n;
  wire g2068_p;
  wire g2068_n;
  wire g2069_p;
  wire g2069_n;
  wire g2070_p;
  wire g2070_n;
  wire g2071_p;
  wire g2071_n;
  wire g2072_p;
  wire g2072_n;
  wire g2073_p;
  wire g2073_n;
  wire g2074_p;
  wire g2074_n;
  wire g2075_p;
  wire g2075_n;
  wire g2076_p;
  wire g2076_n;
  wire g2077_p;
  wire g2077_n;
  wire g2078_p;
  wire g2078_n;
  wire g2079_p;
  wire g2079_n;
  wire g2080_p;
  wire g2080_n;
  wire g2081_p;
  wire g2081_n;
  wire g2082_p;
  wire g2082_n;
  wire g2083_p;
  wire g2083_n;
  wire g2084_p;
  wire g2084_n;
  wire g2085_p;
  wire g2085_n;
  wire g2086_p;
  wire g2086_n;
  wire g2087_p;
  wire g2087_n;
  wire g2088_p;
  wire g2088_n;
  wire g2089_p;
  wire g2089_n;
  wire g2090_p;
  wire g2090_n;
  wire g2091_p;
  wire g2091_n;
  wire g2092_p;
  wire g2092_n;
  wire g2093_p;
  wire g2093_n;
  wire g2094_p;
  wire g2094_n;
  wire g2095_p;
  wire g2095_n;
  wire g2096_p;
  wire g2096_n;
  wire g2097_p;
  wire g2097_n;
  wire g2098_p;
  wire g2098_n;
  wire g2099_p;
  wire g2099_n;
  wire g2100_p;
  wire g2100_n;
  wire g2101_p;
  wire g2101_n;
  wire g2102_p;
  wire g2102_n;
  wire g2103_p;
  wire g2103_n;
  wire g2104_p;
  wire g2104_n;
  wire g2105_p;
  wire g2105_n;
  wire g2106_p;
  wire g2106_n;
  wire g2107_p;
  wire g2107_n;
  wire g2108_p;
  wire g2108_n;
  wire g2109_p;
  wire g2109_n;
  wire g2110_p;
  wire g2110_n;
  wire g2111_p;
  wire g2111_n;
  wire g2112_p;
  wire g2112_n;
  wire g2113_p;
  wire g2113_n;
  wire g2114_p;
  wire g2114_n;
  wire g2115_p;
  wire g2115_n;
  wire g2116_p;
  wire g2116_n;
  wire g2117_p;
  wire g2117_n;
  wire g2118_p;
  wire g2118_n;
  wire g2119_p;
  wire g2119_n;
  wire g2120_p;
  wire g2120_n;
  wire g2121_p;
  wire g2121_n;
  wire g2122_p;
  wire g2122_n;
  wire g2123_p;
  wire g2123_n;
  wire g2124_p;
  wire g2124_n;
  wire g2125_p;
  wire g2125_n;
  wire g2126_p;
  wire g2126_n;
  wire g2127_p;
  wire g2127_n;
  wire g2128_p;
  wire g2128_n;
  wire g2129_p;
  wire g2129_n;
  wire g2130_p;
  wire g2130_n;
  wire g2131_p;
  wire g2131_n;
  wire g2132_p;
  wire g2132_n;
  wire g2133_p;
  wire g2133_n;
  wire g2134_p;
  wire g2134_n;
  wire g2135_p;
  wire g2135_n;
  wire g2136_p;
  wire g2136_n;
  wire g2137_p;
  wire g2137_n;
  wire g2138_p;
  wire g2138_n;
  wire g2139_p;
  wire g2139_n;
  wire g2140_p;
  wire g2140_n;
  wire g2141_p;
  wire g2141_n;
  wire g2142_p;
  wire g2142_n;
  wire g2143_p;
  wire g2143_n;
  wire g2144_p;
  wire g2144_n;
  wire g2145_p;
  wire g2145_n;
  wire g2146_p;
  wire g2146_n;
  wire g2147_p;
  wire g2147_n;
  wire g2148_p;
  wire g2148_n;
  wire g2149_p;
  wire g2149_n;
  wire g2150_p;
  wire g2150_n;
  wire g2151_p;
  wire g2151_n;
  wire g2152_p;
  wire g2152_n;
  wire g2153_p;
  wire g2153_n;
  wire g2154_p;
  wire g2154_n;
  wire g2155_p;
  wire g2155_n;
  wire g2156_p;
  wire g2156_n;
  wire g2157_p;
  wire g2157_n;
  wire g2158_p;
  wire g2158_n;
  wire g2159_p;
  wire g2159_n;
  wire g2160_p;
  wire g2160_n;
  wire g2161_p;
  wire g2161_n;
  wire g2162_p;
  wire g2162_n;
  wire g2163_p;
  wire g2163_n;
  wire g2164_p;
  wire g2164_n;
  wire g2165_p;
  wire g2165_n;
  wire g2166_p;
  wire g2166_n;
  wire g2167_p;
  wire g2167_n;
  wire g2168_p;
  wire g2168_n;
  wire g2169_p;
  wire g2169_n;
  wire g2170_p;
  wire g2170_n;
  wire g2171_p;
  wire g2171_n;
  wire g2172_p;
  wire g2172_n;
  wire g2173_p;
  wire g2173_n;
  wire g2174_p;
  wire g2174_n;
  wire g2175_p;
  wire g2175_n;
  wire g2176_p;
  wire g2176_n;
  wire g2177_p;
  wire g2177_n;
  wire g2178_p;
  wire g2178_n;
  wire g2179_p;
  wire g2179_n;
  wire g2180_p;
  wire g2180_n;
  wire g2181_p;
  wire g2181_n;
  wire g2182_p;
  wire g2182_n;
  wire g2183_p;
  wire g2183_n;
  wire g2184_p;
  wire g2184_n;
  wire g2185_p;
  wire g2185_n;
  wire g2186_p;
  wire g2186_n;
  wire g2187_p;
  wire g2187_n;
  wire g2188_p;
  wire g2188_n;
  wire g2189_p;
  wire g2189_n;
  wire g2190_p;
  wire g2190_n;
  wire g2191_p;
  wire g2191_n;
  wire g2192_p;
  wire g2192_n;
  wire g2193_p;
  wire g2193_n;
  wire g2194_p;
  wire g2194_n;
  wire g2195_p;
  wire g2195_n;
  wire g2196_p;
  wire g2196_n;
  wire g2197_p;
  wire g2197_n;
  wire g2198_p;
  wire g2198_n;
  wire g2199_p;
  wire g2199_n;
  wire g2200_p;
  wire g2200_n;
  wire g2201_p;
  wire g2201_n;
  wire g2202_p;
  wire g2202_n;
  wire g2203_p;
  wire g2203_n;
  wire g2204_p;
  wire g2204_n;
  wire g2205_p;
  wire g2205_n;
  wire g2206_p;
  wire g2206_n;
  wire g2207_p;
  wire g2207_n;
  wire g2208_p;
  wire g2208_n;
  wire g2209_p;
  wire g2209_n;
  wire g2210_p;
  wire g2210_n;
  wire g2211_p;
  wire g2211_n;
  wire g2212_p;
  wire g2212_n;
  wire g2213_p;
  wire g2213_n;
  wire g2214_p;
  wire g2214_n;
  wire g2215_p;
  wire g2215_n;
  wire g2216_p;
  wire g2216_n;
  wire g2217_p;
  wire g2217_n;
  wire g2218_p;
  wire g2218_n;
  wire g2219_p;
  wire g2219_n;
  wire g2220_p;
  wire g2220_n;
  wire g2221_p;
  wire g2221_n;
  wire g2222_p;
  wire g2222_n;
  wire g2223_p;
  wire g2223_n;
  wire g2224_p;
  wire g2224_n;
  wire g2225_p;
  wire g2225_n;
  wire g2226_p;
  wire g2226_n;
  wire g2227_p;
  wire g2227_n;
  wire g2228_p;
  wire g2228_n;
  wire g2229_p;
  wire g2229_n;
  wire g2230_p;
  wire g2230_n;
  wire g2231_p;
  wire g2231_n;
  wire g2232_p;
  wire g2232_n;
  wire g2233_p;
  wire g2233_n;
  wire g2234_p;
  wire g2234_n;
  wire g2235_p;
  wire g2235_n;
  wire g2236_p;
  wire g2236_n;
  wire g2237_p;
  wire g2237_n;
  wire g2238_p;
  wire g2238_n;
  wire g2239_p;
  wire g2239_n;
  wire g2240_p;
  wire g2240_n;
  wire g2241_p;
  wire g2241_n;
  wire g2242_p;
  wire g2242_n;
  wire g2243_p;
  wire g2243_n;
  wire g2244_p;
  wire g2244_n;
  wire g2245_p;
  wire g2245_n;
  wire g2246_p;
  wire g2246_n;
  wire g2247_p;
  wire g2247_n;
  wire g2248_p;
  wire g2248_n;
  wire g2249_p;
  wire g2249_n;
  wire g2250_p;
  wire g2250_n;
  wire g2251_p;
  wire g2251_n;
  wire g2252_p;
  wire g2252_n;
  wire g2253_p;
  wire g2253_n;
  wire g2254_p;
  wire g2254_n;
  wire g2255_p;
  wire g2255_n;
  wire g2256_p;
  wire g2256_n;
  wire g2257_p;
  wire g2257_n;
  wire g2258_p;
  wire g2258_n;
  wire ffc_244_p_spl_;
  wire ffc_242_p_spl_;
  wire ffc_242_n_spl_;
  wire g432_p_spl_;
  wire g433_n_spl_;
  wire g434_p_spl_;
  wire ffc_232_n_spl_;
  wire ffc_232_p_spl_;
  wire g438_n_spl_;
  wire g439_p_spl_;
  wire g438_p_spl_;
  wire g439_n_spl_;
  wire g440_n_spl_;
  wire g440_p_spl_;
  wire g437_p_spl_;
  wire g442_n_spl_;
  wire g443_p_spl_;
  wire ffc_30_p_spl_;
  wire ffc_30_p_spl_0;
  wire ffc_30_p_spl_00;
  wire ffc_30_p_spl_01;
  wire ffc_30_p_spl_1;
  wire ffc_30_p_spl_10;
  wire ffc_30_n_spl_;
  wire ffc_30_n_spl_0;
  wire ffc_30_n_spl_00;
  wire ffc_30_n_spl_01;
  wire ffc_30_n_spl_1;
  wire ffc_30_n_spl_10;
  wire ffc_240_p_spl_;
  wire ffc_240_n_spl_;
  wire g448_n_spl_;
  wire g449_p_spl_;
  wire g448_p_spl_;
  wire g449_n_spl_;
  wire g450_n_spl_;
  wire g450_p_spl_;
  wire g447_n_spl_;
  wire g452_p_spl_;
  wire g447_p_spl_;
  wire g452_n_spl_;
  wire g453_n_spl_;
  wire g453_p_spl_;
  wire g446_p_spl_;
  wire g455_n_spl_;
  wire g456_p_spl_;
  wire ffc_234_n_spl_;
  wire ffc_234_p_spl_;
  wire g462_n_spl_;
  wire g463_p_spl_;
  wire g462_p_spl_;
  wire g463_n_spl_;
  wire g464_n_spl_;
  wire g464_p_spl_;
  wire g461_n_spl_;
  wire g466_p_spl_;
  wire g461_p_spl_;
  wire g466_n_spl_;
  wire g467_n_spl_;
  wire g467_p_spl_;
  wire g460_n_spl_;
  wire g469_p_spl_;
  wire g460_p_spl_;
  wire g469_n_spl_;
  wire g470_n_spl_;
  wire g470_p_spl_;
  wire g459_p_spl_;
  wire g472_n_spl_;
  wire g473_p_spl_;
  wire ffc_4_p_spl_;
  wire ffc_26_p_spl_;
  wire ffc_26_p_spl_0;
  wire ffc_26_p_spl_1;
  wire ffc_4_n_spl_;
  wire ffc_26_n_spl_;
  wire ffc_26_n_spl_0;
  wire ffc_26_n_spl_1;
  wire ffc_238_p_spl_;
  wire ffc_238_n_spl_;
  wire g480_n_spl_;
  wire g481_p_spl_;
  wire g480_p_spl_;
  wire g481_n_spl_;
  wire g482_n_spl_;
  wire g482_p_spl_;
  wire g479_n_spl_;
  wire g484_p_spl_;
  wire g479_p_spl_;
  wire g484_n_spl_;
  wire g485_n_spl_;
  wire g485_p_spl_;
  wire g478_n_spl_;
  wire g487_p_spl_;
  wire g478_p_spl_;
  wire g487_n_spl_;
  wire g488_n_spl_;
  wire g488_p_spl_;
  wire g477_n_spl_;
  wire g490_p_spl_;
  wire g477_p_spl_;
  wire g490_n_spl_;
  wire g491_n_spl_;
  wire g491_p_spl_;
  wire g476_p_spl_;
  wire g493_n_spl_;
  wire g494_p_spl_;
  wire ffc_5_p_spl_;
  wire ffc_5_n_spl_;
  wire ffc_236_n_spl_;
  wire ffc_236_p_spl_;
  wire g502_n_spl_;
  wire g503_p_spl_;
  wire g502_p_spl_;
  wire g503_n_spl_;
  wire g504_n_spl_;
  wire g504_p_spl_;
  wire g501_n_spl_;
  wire g506_p_spl_;
  wire g501_p_spl_;
  wire g506_n_spl_;
  wire g507_n_spl_;
  wire g507_p_spl_;
  wire g500_n_spl_;
  wire g509_p_spl_;
  wire g500_p_spl_;
  wire g509_n_spl_;
  wire g510_n_spl_;
  wire g510_p_spl_;
  wire g499_n_spl_;
  wire g512_p_spl_;
  wire g499_p_spl_;
  wire g512_n_spl_;
  wire g513_n_spl_;
  wire g513_p_spl_;
  wire g498_n_spl_;
  wire g515_p_spl_;
  wire g498_p_spl_;
  wire g515_n_spl_;
  wire g516_n_spl_;
  wire g516_p_spl_;
  wire g497_p_spl_;
  wire g518_n_spl_;
  wire g519_p_spl_;
  wire ffc_6_p_spl_;
  wire ffc_6_n_spl_;
  wire ffc_7_p_spl_;
  wire ffc_7_p_spl_0;
  wire ffc_7_n_spl_;
  wire ffc_7_n_spl_0;
  wire g527_n_spl_;
  wire g528_n_spl_;
  wire g527_p_spl_;
  wire g528_p_spl_;
  wire g529_n_spl_;
  wire g529_p_spl_;
  wire g526_n_spl_;
  wire g531_p_spl_;
  wire g526_p_spl_;
  wire g531_n_spl_;
  wire g532_n_spl_;
  wire g532_p_spl_;
  wire g525_n_spl_;
  wire g534_p_spl_;
  wire g525_p_spl_;
  wire g534_n_spl_;
  wire g535_n_spl_;
  wire g535_p_spl_;
  wire g524_n_spl_;
  wire g537_p_spl_;
  wire g524_p_spl_;
  wire g537_n_spl_;
  wire g538_n_spl_;
  wire g538_p_spl_;
  wire g523_n_spl_;
  wire g540_p_spl_;
  wire g523_p_spl_;
  wire g540_n_spl_;
  wire g541_n_spl_;
  wire g541_p_spl_;
  wire g522_p_spl_;
  wire g543_n_spl_;
  wire g544_p_spl_;
  wire g550_n_spl_;
  wire g551_n_spl_;
  wire g550_p_spl_;
  wire g551_p_spl_;
  wire g552_n_spl_;
  wire g552_p_spl_;
  wire g549_n_spl_;
  wire g554_p_spl_;
  wire g549_p_spl_;
  wire g554_n_spl_;
  wire g555_n_spl_;
  wire g555_p_spl_;
  wire g548_n_spl_;
  wire g557_p_spl_;
  wire g548_p_spl_;
  wire g557_n_spl_;
  wire g558_n_spl_;
  wire g558_p_spl_;
  wire g547_p_spl_;
  wire g560_n_spl_;
  wire g561_p_spl_;
  wire g564_n_spl_;
  wire g565_n_spl_;
  wire g564_p_spl_;
  wire g565_p_spl_;
  wire g566_n_spl_;
  wire g570_n_spl_;
  wire ffc_25_p_spl_;
  wire ffc_25_p_spl_0;
  wire ffc_25_p_spl_00;
  wire ffc_25_p_spl_000;
  wire ffc_25_p_spl_001;
  wire ffc_25_p_spl_01;
  wire ffc_25_p_spl_010;
  wire ffc_25_p_spl_011;
  wire ffc_25_p_spl_1;
  wire ffc_25_p_spl_10;
  wire ffc_25_p_spl_11;
  wire ffc_80_p_spl_;
  wire ffc_25_n_spl_;
  wire ffc_25_n_spl_0;
  wire ffc_25_n_spl_00;
  wire ffc_25_n_spl_000;
  wire ffc_25_n_spl_001;
  wire ffc_25_n_spl_01;
  wire ffc_25_n_spl_010;
  wire ffc_25_n_spl_011;
  wire ffc_25_n_spl_1;
  wire ffc_25_n_spl_10;
  wire ffc_25_n_spl_11;
  wire ffc_80_n_spl_;
  wire ffc_272_p_spl_;
  wire g575_n_spl_;
  wire g576_p_spl_;
  wire g575_p_spl_;
  wire g576_n_spl_;
  wire g577_n_spl_;
  wire g577_p_spl_;
  wire g579_p_spl_;
  wire g574_p_spl_;
  wire ffc_29_n_spl_;
  wire ffc_29_n_spl_0;
  wire ffc_29_n_spl_00;
  wire ffc_29_n_spl_000;
  wire ffc_29_n_spl_01;
  wire ffc_29_n_spl_1;
  wire ffc_29_n_spl_10;
  wire ffc_29_n_spl_11;
  wire g580_p_spl_;
  wire ffc_79_p_spl_;
  wire ffc_79_n_spl_;
  wire ffc_270_n_spl_;
  wire ffc_275_n_spl_;
  wire ffc_270_p_spl_;
  wire ffc_275_p_spl_;
  wire g584_n_spl_;
  wire g584_p_spl_;
  wire g583_n_spl_;
  wire g586_p_spl_;
  wire g583_p_spl_;
  wire g586_n_spl_;
  wire g587_n_spl_;
  wire g587_p_spl_;
  wire g582_n_spl_;
  wire g589_p_spl_;
  wire g581_n_spl_;
  wire g592_p_spl_;
  wire g593_p_spl_;
  wire ffc_29_p_spl_;
  wire ffc_29_p_spl_0;
  wire ffc_29_p_spl_00;
  wire ffc_29_p_spl_01;
  wire ffc_29_p_spl_1;
  wire ffc_29_p_spl_10;
  wire ffc_29_p_spl_11;
  wire ffc_64_p_spl_;
  wire ffc_64_n_spl_;
  wire ffc_268_n_spl_;
  wire ffc_276_n_spl_;
  wire ffc_268_p_spl_;
  wire ffc_276_p_spl_;
  wire g598_n_spl_;
  wire g598_p_spl_;
  wire g597_n_spl_;
  wire g600_p_spl_;
  wire g597_p_spl_;
  wire g600_n_spl_;
  wire g601_n_spl_;
  wire g601_p_spl_;
  wire g596_n_spl_;
  wire g603_p_spl_;
  wire g596_p_spl_;
  wire g603_n_spl_;
  wire g604_n_spl_;
  wire g604_p_spl_;
  wire g595_n_spl_;
  wire g606_p_spl_;
  wire g607_n_spl_;
  wire g594_n_spl_;
  wire g609_p_spl_;
  wire ffc_65_p_spl_;
  wire ffc_65_n_spl_;
  wire ffc_269_n_spl_;
  wire ffc_277_n_spl_;
  wire ffc_269_p_spl_;
  wire ffc_277_p_spl_;
  wire g615_n_spl_;
  wire g615_p_spl_;
  wire g614_n_spl_;
  wire g617_p_spl_;
  wire g614_p_spl_;
  wire g617_n_spl_;
  wire g618_n_spl_;
  wire g618_p_spl_;
  wire g613_n_spl_;
  wire g620_p_spl_;
  wire g613_p_spl_;
  wire g620_n_spl_;
  wire g621_n_spl_;
  wire g621_p_spl_;
  wire g612_n_spl_;
  wire g623_p_spl_;
  wire g612_p_spl_;
  wire g623_n_spl_;
  wire g624_n_spl_;
  wire g624_p_spl_;
  wire g611_n_spl_;
  wire g626_p_spl_;
  wire ffc_135_p_spl_;
  wire ffc_135_p_spl_0;
  wire ffc_135_p_spl_00;
  wire ffc_135_p_spl_1;
  wire ffc_287_p_spl_;
  wire ffc_287_p_spl_0;
  wire ffc_287_p_spl_00;
  wire ffc_287_p_spl_000;
  wire ffc_287_p_spl_001;
  wire ffc_287_p_spl_01;
  wire ffc_287_p_spl_010;
  wire ffc_287_p_spl_011;
  wire ffc_287_p_spl_1;
  wire ffc_287_p_spl_10;
  wire ffc_287_p_spl_100;
  wire ffc_287_p_spl_101;
  wire ffc_287_p_spl_11;
  wire ffc_287_p_spl_110;
  wire ffc_287_p_spl_111;
  wire ffc_135_n_spl_;
  wire ffc_135_n_spl_0;
  wire ffc_135_n_spl_00;
  wire ffc_135_n_spl_1;
  wire ffc_287_n_spl_;
  wire ffc_287_n_spl_0;
  wire ffc_287_n_spl_00;
  wire ffc_287_n_spl_000;
  wire ffc_287_n_spl_001;
  wire ffc_287_n_spl_01;
  wire ffc_287_n_spl_010;
  wire ffc_287_n_spl_011;
  wire ffc_287_n_spl_1;
  wire ffc_287_n_spl_10;
  wire ffc_287_n_spl_100;
  wire ffc_287_n_spl_101;
  wire ffc_287_n_spl_11;
  wire ffc_287_n_spl_110;
  wire ffc_287_n_spl_111;
  wire g610_n_spl_;
  wire g629_p_spl_;
  wire ffc_285_n_spl_;
  wire ffc_286_n_spl_;
  wire ffc_285_p_spl_;
  wire ffc_286_p_spl_;
  wire g632_n_spl_;
  wire g632_p_spl_;
  wire g634_p_spl_;
  wire g630_p_spl_;
  wire g631_p_spl_;
  wire ffc_66_p_spl_;
  wire ffc_66_n_spl_;
  wire ffc_261_n_spl_;
  wire ffc_284_p_spl_;
  wire ffc_261_p_spl_;
  wire ffc_284_n_spl_;
  wire g642_n_spl_;
  wire g642_p_spl_;
  wire g641_n_spl_;
  wire g644_p_spl_;
  wire g641_p_spl_;
  wire g644_n_spl_;
  wire g645_n_spl_;
  wire g645_p_spl_;
  wire g640_n_spl_;
  wire g647_p_spl_;
  wire g640_p_spl_;
  wire g647_n_spl_;
  wire g648_n_spl_;
  wire g648_p_spl_;
  wire g639_n_spl_;
  wire g650_p_spl_;
  wire g639_p_spl_;
  wire g650_n_spl_;
  wire g651_n_spl_;
  wire g651_p_spl_;
  wire g638_n_spl_;
  wire g653_p_spl_;
  wire g638_p_spl_;
  wire g653_n_spl_;
  wire g654_n_spl_;
  wire g654_p_spl_;
  wire g637_n_spl_;
  wire g656_p_spl_;
  wire ffc_15_p_spl_;
  wire ffc_15_p_spl_0;
  wire ffc_15_p_spl_00;
  wire ffc_15_p_spl_000;
  wire ffc_15_p_spl_001;
  wire ffc_15_p_spl_01;
  wire ffc_15_p_spl_010;
  wire ffc_15_p_spl_011;
  wire ffc_15_p_spl_1;
  wire ffc_15_p_spl_10;
  wire ffc_15_p_spl_100;
  wire ffc_15_p_spl_101;
  wire ffc_15_p_spl_11;
  wire ffc_15_p_spl_110;
  wire ffc_15_p_spl_111;
  wire ffc_15_n_spl_;
  wire ffc_15_n_spl_0;
  wire ffc_15_n_spl_00;
  wire ffc_15_n_spl_000;
  wire ffc_15_n_spl_001;
  wire ffc_15_n_spl_01;
  wire ffc_15_n_spl_010;
  wire ffc_15_n_spl_011;
  wire ffc_15_n_spl_1;
  wire ffc_15_n_spl_10;
  wire ffc_15_n_spl_100;
  wire ffc_15_n_spl_101;
  wire ffc_15_n_spl_11;
  wire g636_n_spl_;
  wire g659_p_spl_;
  wire g635_p_spl_;
  wire ffc_133_p_spl_;
  wire ffc_133_p_spl_0;
  wire ffc_133_p_spl_00;
  wire ffc_133_p_spl_1;
  wire ffc_133_n_spl_;
  wire ffc_133_n_spl_0;
  wire ffc_133_n_spl_00;
  wire ffc_133_n_spl_1;
  wire ffc_310_p_spl_;
  wire ffc_310_n_spl_;
  wire g663_n_spl_;
  wire g664_p_spl_;
  wire g663_p_spl_;
  wire g664_n_spl_;
  wire g665_n_spl_;
  wire g665_p_spl_;
  wire g662_n_spl_;
  wire g667_p_spl_;
  wire g662_p_spl_;
  wire g667_n_spl_;
  wire g668_n_spl_;
  wire g668_p_spl_;
  wire g670_p_spl_;
  wire g660_p_spl_;
  wire ffc_207_p_spl_;
  wire ffc_207_p_spl_0;
  wire ffc_207_p_spl_00;
  wire ffc_207_p_spl_1;
  wire ffc_325_p_spl_;
  wire ffc_325_p_spl_0;
  wire ffc_207_n_spl_;
  wire ffc_207_n_spl_0;
  wire ffc_207_n_spl_00;
  wire ffc_207_n_spl_1;
  wire ffc_325_n_spl_;
  wire ffc_325_n_spl_0;
  wire ffc_341_p_spl_;
  wire ffc_341_n_spl_;
  wire g661_p_spl_;
  wire ffc_67_p_spl_;
  wire ffc_67_n_spl_;
  wire ffc_68_p_spl_;
  wire ffc_68_p_spl_0;
  wire ffc_214_p_spl_;
  wire ffc_214_p_spl_0;
  wire ffc_214_p_spl_00;
  wire ffc_214_p_spl_000;
  wire ffc_214_p_spl_01;
  wire ffc_214_p_spl_1;
  wire ffc_214_p_spl_10;
  wire ffc_214_p_spl_11;
  wire ffc_68_n_spl_;
  wire ffc_68_n_spl_0;
  wire ffc_214_n_spl_;
  wire ffc_214_n_spl_0;
  wire ffc_214_n_spl_00;
  wire ffc_214_n_spl_000;
  wire ffc_214_n_spl_01;
  wire ffc_214_n_spl_1;
  wire ffc_214_n_spl_10;
  wire ffc_214_n_spl_11;
  wire ffc_267_n_spl_;
  wire ffc_278_n_spl_;
  wire ffc_267_p_spl_;
  wire ffc_278_p_spl_;
  wire g681_n_spl_;
  wire g681_p_spl_;
  wire g680_n_spl_;
  wire g683_p_spl_;
  wire g680_p_spl_;
  wire g683_n_spl_;
  wire g684_n_spl_;
  wire g684_p_spl_;
  wire g679_n_spl_;
  wire g686_p_spl_;
  wire g679_p_spl_;
  wire g686_n_spl_;
  wire g687_n_spl_;
  wire g687_p_spl_;
  wire g678_n_spl_;
  wire g689_p_spl_;
  wire g678_p_spl_;
  wire g689_n_spl_;
  wire g690_n_spl_;
  wire g690_p_spl_;
  wire g677_n_spl_;
  wire g692_p_spl_;
  wire g677_p_spl_;
  wire g692_n_spl_;
  wire g693_n_spl_;
  wire g693_p_spl_;
  wire g676_n_spl_;
  wire g695_p_spl_;
  wire g676_p_spl_;
  wire g695_n_spl_;
  wire g696_n_spl_;
  wire g696_p_spl_;
  wire g675_n_spl_;
  wire g698_p_spl_;
  wire g673_p_spl_;
  wire g672_p_spl_;
  wire ffc_17_p_spl_;
  wire ffc_17_p_spl_0;
  wire ffc_17_p_spl_00;
  wire ffc_17_p_spl_000;
  wire ffc_17_p_spl_001;
  wire ffc_17_p_spl_01;
  wire ffc_17_p_spl_010;
  wire ffc_17_p_spl_011;
  wire ffc_17_p_spl_1;
  wire ffc_17_p_spl_10;
  wire ffc_17_p_spl_100;
  wire ffc_17_p_spl_11;
  wire ffc_17_n_spl_;
  wire ffc_17_n_spl_0;
  wire ffc_17_n_spl_00;
  wire ffc_17_n_spl_000;
  wire ffc_17_n_spl_001;
  wire ffc_17_n_spl_01;
  wire ffc_17_n_spl_010;
  wire ffc_17_n_spl_1;
  wire ffc_17_n_spl_10;
  wire ffc_17_n_spl_11;
  wire ffc_9_p_spl_;
  wire ffc_9_p_spl_0;
  wire ffc_9_p_spl_00;
  wire ffc_9_p_spl_000;
  wire ffc_9_p_spl_001;
  wire ffc_9_p_spl_01;
  wire ffc_9_p_spl_010;
  wire ffc_9_p_spl_011;
  wire ffc_9_p_spl_1;
  wire ffc_9_p_spl_10;
  wire ffc_9_p_spl_100;
  wire ffc_9_p_spl_101;
  wire ffc_9_p_spl_11;
  wire ffc_9_p_spl_110;
  wire ffc_9_p_spl_111;
  wire ffc_9_n_spl_;
  wire ffc_9_n_spl_0;
  wire ffc_9_n_spl_00;
  wire ffc_9_n_spl_000;
  wire ffc_9_n_spl_001;
  wire ffc_9_n_spl_01;
  wire ffc_9_n_spl_010;
  wire ffc_9_n_spl_011;
  wire ffc_9_n_spl_1;
  wire ffc_9_n_spl_10;
  wire ffc_9_n_spl_100;
  wire ffc_9_n_spl_101;
  wire ffc_9_n_spl_11;
  wire ffc_9_n_spl_110;
  wire ffc_9_n_spl_111;
  wire ffc_264_n_spl_;
  wire ffc_281_p_spl_;
  wire ffc_264_p_spl_;
  wire ffc_281_n_spl_;
  wire g706_n_spl_;
  wire g706_p_spl_;
  wire g705_n_spl_;
  wire g708_p_spl_;
  wire g705_p_spl_;
  wire g708_n_spl_;
  wire ffc_75_p_spl_;
  wire ffc_75_p_spl_0;
  wire ffc_75_p_spl_1;
  wire ffc_160_p_spl_;
  wire ffc_160_p_spl_0;
  wire ffc_160_p_spl_1;
  wire ffc_75_n_spl_;
  wire ffc_75_n_spl_0;
  wire ffc_160_n_spl_;
  wire ffc_160_n_spl_0;
  wire ffc_160_n_spl_1;
  wire g709_n_spl_;
  wire g709_p_spl_;
  wire g710_n_spl_;
  wire g712_p_spl_;
  wire g710_p_spl_;
  wire g712_n_spl_;
  wire g713_n_spl_;
  wire g713_p_spl_;
  wire ffc_76_p_spl_;
  wire ffc_76_p_spl_0;
  wire ffc_76_n_spl_;
  wire ffc_76_n_spl_0;
  wire ffc_77_p_spl_;
  wire ffc_77_p_spl_0;
  wire ffc_77_p_spl_1;
  wire ffc_77_n_spl_;
  wire ffc_77_n_spl_0;
  wire g716_n_spl_;
  wire g717_n_spl_;
  wire g716_p_spl_;
  wire g717_p_spl_;
  wire g718_n_spl_;
  wire g718_p_spl_;
  wire g715_n_spl_;
  wire g720_p_spl_;
  wire g715_p_spl_;
  wire g720_n_spl_;
  wire g721_n_spl_;
  wire g721_p_spl_;
  wire g714_n_spl_;
  wire g723_p_spl_;
  wire g714_p_spl_;
  wire g723_n_spl_;
  wire ffc_174_p_spl_;
  wire ffc_174_p_spl_0;
  wire ffc_174_p_spl_00;
  wire ffc_174_p_spl_01;
  wire ffc_174_p_spl_1;
  wire ffc_174_p_spl_10;
  wire ffc_174_n_spl_;
  wire ffc_174_n_spl_0;
  wire ffc_174_n_spl_00;
  wire ffc_174_n_spl_01;
  wire ffc_174_n_spl_1;
  wire ffc_174_n_spl_10;
  wire g724_n_spl_;
  wire g724_p_spl_;
  wire g725_n_spl_;
  wire g727_p_spl_;
  wire g725_p_spl_;
  wire g727_n_spl_;
  wire g728_n_spl_;
  wire g728_p_spl_;
  wire g731_n_spl_;
  wire g732_n_spl_;
  wire g731_p_spl_;
  wire g732_p_spl_;
  wire g733_n_spl_;
  wire g733_p_spl_;
  wire g730_n_spl_;
  wire g735_p_spl_;
  wire g730_p_spl_;
  wire g735_n_spl_;
  wire g736_n_spl_;
  wire g736_p_spl_;
  wire g729_n_spl_;
  wire g738_p_spl_;
  wire g729_p_spl_;
  wire g738_n_spl_;
  wire ffc_263_n_spl_;
  wire ffc_282_p_spl_;
  wire ffc_263_p_spl_;
  wire ffc_282_n_spl_;
  wire g741_n_spl_;
  wire g741_p_spl_;
  wire g740_n_spl_;
  wire g743_p_spl_;
  wire g740_p_spl_;
  wire g743_n_spl_;
  wire ffc_72_p_spl_;
  wire ffc_72_p_spl_0;
  wire ffc_72_p_spl_1;
  wire ffc_72_n_spl_;
  wire ffc_72_n_spl_0;
  wire g744_n_spl_;
  wire g744_p_spl_;
  wire g745_n_spl_;
  wire g747_p_spl_;
  wire g745_p_spl_;
  wire g747_n_spl_;
  wire g748_n_spl_;
  wire g748_p_spl_;
  wire ffc_73_p_spl_;
  wire ffc_73_p_spl_0;
  wire ffc_73_n_spl_;
  wire ffc_73_n_spl_0;
  wire ffc_74_p_spl_;
  wire ffc_74_p_spl_0;
  wire ffc_74_p_spl_1;
  wire ffc_74_n_spl_;
  wire ffc_74_n_spl_0;
  wire ffc_265_n_spl_;
  wire ffc_280_n_spl_;
  wire ffc_265_p_spl_;
  wire ffc_280_p_spl_;
  wire g753_n_spl_;
  wire g753_p_spl_;
  wire g752_n_spl_;
  wire g755_p_spl_;
  wire g752_p_spl_;
  wire g755_n_spl_;
  wire g756_n_spl_;
  wire g756_p_spl_;
  wire g751_n_spl_;
  wire g758_p_spl_;
  wire g751_p_spl_;
  wire g758_n_spl_;
  wire g759_n_spl_;
  wire g759_p_spl_;
  wire g750_n_spl_;
  wire g761_p_spl_;
  wire g750_p_spl_;
  wire g761_n_spl_;
  wire g762_n_spl_;
  wire g762_p_spl_;
  wire g749_n_spl_;
  wire g764_p_spl_;
  wire g749_p_spl_;
  wire g764_n_spl_;
  wire g765_n_spl_;
  wire g765_p_spl_;
  wire g766_n_spl_;
  wire g768_p_spl_;
  wire g766_p_spl_;
  wire g768_n_spl_;
  wire g769_n_spl_;
  wire g769_p_spl_;
  wire g774_n_spl_;
  wire g776_p_spl_;
  wire g774_p_spl_;
  wire g776_n_spl_;
  wire g777_n_spl_;
  wire g777_p_spl_;
  wire g773_n_spl_;
  wire g779_p_spl_;
  wire g773_p_spl_;
  wire g779_n_spl_;
  wire g780_n_spl_;
  wire g780_p_spl_;
  wire g772_n_spl_;
  wire g782_p_spl_;
  wire g772_p_spl_;
  wire g782_n_spl_;
  wire g783_n_spl_;
  wire g783_p_spl_;
  wire g771_n_spl_;
  wire g785_p_spl_;
  wire g771_p_spl_;
  wire g785_n_spl_;
  wire g786_n_spl_;
  wire g786_p_spl_;
  wire g770_n_spl_;
  wire g788_p_spl_;
  wire g770_p_spl_;
  wire g788_n_spl_;
  wire ffc_262_n_spl_;
  wire ffc_283_p_spl_;
  wire ffc_262_p_spl_;
  wire ffc_283_n_spl_;
  wire g791_n_spl_;
  wire g791_p_spl_;
  wire g790_n_spl_;
  wire g793_p_spl_;
  wire g790_p_spl_;
  wire g793_n_spl_;
  wire ffc_69_p_spl_;
  wire ffc_69_p_spl_0;
  wire ffc_69_n_spl_;
  wire ffc_69_n_spl_0;
  wire g794_n_spl_;
  wire g794_p_spl_;
  wire g795_n_spl_;
  wire g797_p_spl_;
  wire g795_p_spl_;
  wire g797_n_spl_;
  wire g798_n_spl_;
  wire g798_p_spl_;
  wire ffc_70_p_spl_;
  wire ffc_70_n_spl_;
  wire ffc_70_n_spl_0;
  wire ffc_71_p_spl_;
  wire ffc_71_p_spl_0;
  wire ffc_71_p_spl_1;
  wire ffc_71_n_spl_;
  wire ffc_71_n_spl_0;
  wire ffc_266_n_spl_;
  wire ffc_279_n_spl_;
  wire ffc_266_p_spl_;
  wire ffc_279_p_spl_;
  wire g803_n_spl_;
  wire g803_p_spl_;
  wire g802_n_spl_;
  wire g805_p_spl_;
  wire g802_p_spl_;
  wire g805_n_spl_;
  wire g806_n_spl_;
  wire g806_p_spl_;
  wire g801_n_spl_;
  wire g808_p_spl_;
  wire g801_p_spl_;
  wire g808_n_spl_;
  wire g809_n_spl_;
  wire g809_p_spl_;
  wire g800_n_spl_;
  wire g811_p_spl_;
  wire g800_p_spl_;
  wire g811_n_spl_;
  wire g812_n_spl_;
  wire g812_p_spl_;
  wire g799_n_spl_;
  wire g814_p_spl_;
  wire g799_p_spl_;
  wire g814_n_spl_;
  wire g815_n_spl_;
  wire g815_p_spl_;
  wire g816_n_spl_;
  wire g818_p_spl_;
  wire g816_p_spl_;
  wire g818_n_spl_;
  wire g819_n_spl_;
  wire g819_p_spl_;
  wire g824_n_spl_;
  wire g826_p_spl_;
  wire g824_p_spl_;
  wire g826_n_spl_;
  wire g827_n_spl_;
  wire g827_p_spl_;
  wire g823_n_spl_;
  wire g829_p_spl_;
  wire g823_p_spl_;
  wire g829_n_spl_;
  wire g830_n_spl_;
  wire g830_p_spl_;
  wire g822_n_spl_;
  wire g832_p_spl_;
  wire g822_p_spl_;
  wire g832_n_spl_;
  wire g833_n_spl_;
  wire g833_p_spl_;
  wire g821_n_spl_;
  wire g835_p_spl_;
  wire g821_p_spl_;
  wire g835_n_spl_;
  wire g836_n_spl_;
  wire g836_p_spl_;
  wire g820_n_spl_;
  wire g838_p_spl_;
  wire g820_p_spl_;
  wire g838_n_spl_;
  wire g674_n_spl_;
  wire g701_p_spl_;
  wire g671_p_spl_;
  wire ffc_118_p_spl_;
  wire ffc_118_p_spl_0;
  wire ffc_118_p_spl_00;
  wire ffc_118_p_spl_01;
  wire ffc_118_p_spl_1;
  wire ffc_118_n_spl_;
  wire ffc_118_n_spl_0;
  wire ffc_118_n_spl_00;
  wire ffc_118_n_spl_1;
  wire ffc_296_p_spl_;
  wire ffc_296_n_spl_;
  wire g844_n_spl_;
  wire g845_p_spl_;
  wire g844_p_spl_;
  wire g845_n_spl_;
  wire g846_n_spl_;
  wire g846_p_spl_;
  wire g843_n_spl_;
  wire g848_p_spl_;
  wire g843_p_spl_;
  wire g848_n_spl_;
  wire g849_n_spl_;
  wire g849_p_spl_;
  wire g842_n_spl_;
  wire g851_p_spl_;
  wire g842_p_spl_;
  wire g851_n_spl_;
  wire g852_n_spl_;
  wire g852_p_spl_;
  wire g841_n_spl_;
  wire g854_p_spl_;
  wire g841_p_spl_;
  wire g854_n_spl_;
  wire g855_n_spl_;
  wire g855_p_spl_;
  wire g702_p_spl_;
  wire ffc_339_n_spl_;
  wire ffc_355_p_spl_;
  wire ffc_339_p_spl_;
  wire ffc_355_n_spl_;
  wire g859_n_spl_;
  wire g859_p_spl_;
  wire g858_n_spl_;
  wire g861_p_spl_;
  wire g858_p_spl_;
  wire g861_n_spl_;
  wire g862_n_spl_;
  wire g862_p_spl_;
  wire g857_p_spl_;
  wire g703_p_spl_;
  wire g864_p_spl_;
  wire g704_p_spl_;
  wire g840_p_spl_;
  wire g872_n_spl_;
  wire g874_p_spl_;
  wire g872_p_spl_;
  wire g874_n_spl_;
  wire g875_n_spl_;
  wire g875_p_spl_;
  wire g871_n_spl_;
  wire g877_p_spl_;
  wire g871_p_spl_;
  wire g877_n_spl_;
  wire g878_n_spl_;
  wire g878_p_spl_;
  wire g870_n_spl_;
  wire g880_p_spl_;
  wire g870_p_spl_;
  wire g880_n_spl_;
  wire g881_n_spl_;
  wire g881_p_spl_;
  wire g869_n_spl_;
  wire g883_p_spl_;
  wire g869_p_spl_;
  wire g883_n_spl_;
  wire g884_n_spl_;
  wire g884_p_spl_;
  wire g868_n_spl_;
  wire g886_p_spl_;
  wire ffc_10_p_spl_;
  wire ffc_10_p_spl_0;
  wire ffc_10_p_spl_00;
  wire ffc_10_p_spl_000;
  wire ffc_10_p_spl_001;
  wire ffc_10_p_spl_01;
  wire ffc_10_p_spl_010;
  wire ffc_10_p_spl_011;
  wire ffc_10_p_spl_1;
  wire ffc_10_p_spl_10;
  wire ffc_10_p_spl_100;
  wire ffc_10_p_spl_101;
  wire ffc_10_p_spl_11;
  wire ffc_10_p_spl_110;
  wire ffc_10_n_spl_;
  wire ffc_10_n_spl_0;
  wire ffc_10_n_spl_00;
  wire ffc_10_n_spl_000;
  wire ffc_10_n_spl_001;
  wire ffc_10_n_spl_01;
  wire ffc_10_n_spl_010;
  wire ffc_10_n_spl_011;
  wire ffc_10_n_spl_1;
  wire ffc_10_n_spl_10;
  wire ffc_10_n_spl_100;
  wire ffc_10_n_spl_101;
  wire ffc_10_n_spl_11;
  wire ffc_10_n_spl_110;
  wire ffc_10_n_spl_111;
  wire g866_p_spl_;
  wire ffc_195_p_spl_;
  wire ffc_195_p_spl_0;
  wire ffc_195_p_spl_00;
  wire ffc_195_p_spl_1;
  wire ffc_195_n_spl_;
  wire ffc_195_n_spl_0;
  wire ffc_195_n_spl_1;
  wire ffc_326_n_spl_;
  wire ffc_343_p_spl_;
  wire ffc_326_p_spl_;
  wire ffc_343_n_spl_;
  wire g894_n_spl_;
  wire g894_p_spl_;
  wire g893_n_spl_;
  wire g896_p_spl_;
  wire g893_p_spl_;
  wire g896_n_spl_;
  wire g897_n_spl_;
  wire g897_p_spl_;
  wire g892_n_spl_;
  wire g899_p_spl_;
  wire g892_p_spl_;
  wire g899_n_spl_;
  wire g900_n_spl_;
  wire g900_p_spl_;
  wire g891_n_spl_;
  wire g902_p_spl_;
  wire g891_p_spl_;
  wire g902_n_spl_;
  wire g903_n_spl_;
  wire g903_p_spl_;
  wire g905_p_spl_;
  wire g890_p_spl_;
  wire ffc_19_p_spl_;
  wire ffc_19_p_spl_0;
  wire ffc_19_p_spl_00;
  wire ffc_19_p_spl_000;
  wire ffc_19_p_spl_001;
  wire ffc_19_p_spl_01;
  wire ffc_19_p_spl_1;
  wire ffc_19_p_spl_10;
  wire ffc_19_p_spl_11;
  wire ffc_19_n_spl_;
  wire ffc_19_n_spl_0;
  wire ffc_19_n_spl_00;
  wire ffc_19_n_spl_01;
  wire ffc_19_n_spl_1;
  wire ffc_19_n_spl_10;
  wire ffc_19_n_spl_11;
  wire g839_n_spl_;
  wire g789_n_spl_;
  wire g739_n_spl_;
  wire g925_n_spl_;
  wire g927_p_spl_;
  wire g925_p_spl_;
  wire g927_n_spl_;
  wire g928_p_spl_;
  wire g924_n_spl_;
  wire g930_p_spl_;
  wire g924_p_spl_;
  wire g930_n_spl_;
  wire g931_p_spl_;
  wire g937_n_spl_;
  wire g939_p_spl_;
  wire g937_p_spl_;
  wire g939_n_spl_;
  wire g940_p_spl_;
  wire g936_n_spl_;
  wire g942_p_spl_;
  wire g936_p_spl_;
  wire g942_n_spl_;
  wire g943_p_spl_;
  wire g949_n_spl_;
  wire g951_p_spl_;
  wire g949_p_spl_;
  wire g951_n_spl_;
  wire g952_p_spl_;
  wire g948_n_spl_;
  wire g954_p_spl_;
  wire g948_p_spl_;
  wire g954_n_spl_;
  wire g955_p_spl_;
  wire g867_n_spl_;
  wire g889_p_spl_;
  wire g865_p_spl_;
  wire ffc_119_p_spl_;
  wire ffc_119_p_spl_0;
  wire ffc_119_p_spl_00;
  wire ffc_119_p_spl_01;
  wire ffc_119_p_spl_1;
  wire ffc_119_n_spl_;
  wire ffc_119_n_spl_0;
  wire ffc_119_n_spl_00;
  wire ffc_119_n_spl_1;
  wire ffc_298_p_spl_;
  wire ffc_298_n_spl_;
  wire g965_n_spl_;
  wire g966_p_spl_;
  wire g965_p_spl_;
  wire g966_n_spl_;
  wire g967_n_spl_;
  wire g967_p_spl_;
  wire g964_n_spl_;
  wire g969_p_spl_;
  wire g964_p_spl_;
  wire g969_n_spl_;
  wire g970_n_spl_;
  wire g970_p_spl_;
  wire g963_n_spl_;
  wire g972_p_spl_;
  wire g963_p_spl_;
  wire g972_n_spl_;
  wire g973_n_spl_;
  wire g973_p_spl_;
  wire g962_n_spl_;
  wire g975_p_spl_;
  wire g962_p_spl_;
  wire g975_n_spl_;
  wire g976_n_spl_;
  wire g976_p_spl_;
  wire g961_n_spl_;
  wire g978_p_spl_;
  wire g961_p_spl_;
  wire g978_n_spl_;
  wire g979_n_spl_;
  wire g979_p_spl_;
  wire g960_n_spl_;
  wire g981_p_spl_;
  wire g960_p_spl_;
  wire g981_n_spl_;
  wire g982_n_spl_;
  wire g982_p_spl_;
  wire G2_p_spl_;
  wire G2_p_spl_0;
  wire G2_p_spl_00;
  wire G2_p_spl_01;
  wire G2_p_spl_1;
  wire G17_p_spl_;
  wire G17_p_spl_0;
  wire G17_p_spl_00;
  wire G17_p_spl_000;
  wire G17_p_spl_001;
  wire G17_p_spl_01;
  wire G17_p_spl_010;
  wire G17_p_spl_011;
  wire G17_p_spl_1;
  wire G17_p_spl_10;
  wire G17_p_spl_100;
  wire G17_p_spl_101;
  wire G17_p_spl_11;
  wire G17_p_spl_110;
  wire G17_p_spl_111;
  wire G2_n_spl_;
  wire G2_n_spl_0;
  wire G2_n_spl_1;
  wire G17_n_spl_;
  wire G17_n_spl_0;
  wire G17_n_spl_00;
  wire G17_n_spl_000;
  wire G17_n_spl_001;
  wire G17_n_spl_01;
  wire G17_n_spl_010;
  wire G17_n_spl_011;
  wire G17_n_spl_1;
  wire G17_n_spl_10;
  wire G17_n_spl_100;
  wire G17_n_spl_101;
  wire G17_n_spl_11;
  wire G17_n_spl_110;
  wire G1_p_spl_;
  wire G1_p_spl_0;
  wire G18_p_spl_;
  wire G18_p_spl_0;
  wire G18_p_spl_00;
  wire G18_p_spl_000;
  wire G18_p_spl_001;
  wire G18_p_spl_01;
  wire G18_p_spl_010;
  wire G18_p_spl_011;
  wire G18_p_spl_1;
  wire G18_p_spl_10;
  wire G18_p_spl_100;
  wire G18_p_spl_101;
  wire G18_p_spl_11;
  wire G18_p_spl_110;
  wire G18_p_spl_111;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire G18_n_spl_;
  wire G18_n_spl_0;
  wire G18_n_spl_00;
  wire G18_n_spl_000;
  wire G18_n_spl_001;
  wire G18_n_spl_01;
  wire G18_n_spl_010;
  wire G18_n_spl_011;
  wire G18_n_spl_1;
  wire G18_n_spl_10;
  wire G18_n_spl_100;
  wire G18_n_spl_101;
  wire G18_n_spl_11;
  wire G18_n_spl_110;
  wire G18_n_spl_111;
  wire g984_p_spl_;
  wire g907_p_spl_;
  wire ffc_11_p_spl_;
  wire ffc_11_p_spl_0;
  wire ffc_11_p_spl_00;
  wire ffc_11_p_spl_000;
  wire ffc_11_p_spl_001;
  wire ffc_11_p_spl_01;
  wire ffc_11_p_spl_010;
  wire ffc_11_p_spl_011;
  wire ffc_11_p_spl_1;
  wire ffc_11_p_spl_10;
  wire ffc_11_p_spl_100;
  wire ffc_11_p_spl_101;
  wire ffc_11_p_spl_11;
  wire ffc_11_n_spl_;
  wire ffc_11_n_spl_0;
  wire ffc_11_n_spl_00;
  wire ffc_11_n_spl_000;
  wire ffc_11_n_spl_001;
  wire ffc_11_n_spl_01;
  wire ffc_11_n_spl_010;
  wire ffc_11_n_spl_011;
  wire ffc_11_n_spl_1;
  wire ffc_11_n_spl_10;
  wire ffc_11_n_spl_100;
  wire ffc_11_n_spl_101;
  wire ffc_11_n_spl_11;
  wire g985_p_spl_;
  wire g986_p_spl_;
  wire g906_p_spl_;
  wire ffc_180_p_spl_;
  wire ffc_180_p_spl_0;
  wire ffc_180_p_spl_00;
  wire ffc_180_p_spl_1;
  wire ffc_180_n_spl_;
  wire ffc_180_n_spl_0;
  wire ffc_180_n_spl_1;
  wire ffc_327_n_spl_;
  wire ffc_344_p_spl_;
  wire ffc_327_p_spl_;
  wire ffc_344_n_spl_;
  wire g995_n_spl_;
  wire g995_p_spl_;
  wire g994_n_spl_;
  wire g997_p_spl_;
  wire g994_p_spl_;
  wire g997_n_spl_;
  wire g998_n_spl_;
  wire g998_p_spl_;
  wire g993_n_spl_;
  wire g1000_p_spl_;
  wire g993_p_spl_;
  wire g1000_n_spl_;
  wire g1001_n_spl_;
  wire g1001_p_spl_;
  wire g992_n_spl_;
  wire g1003_p_spl_;
  wire g992_p_spl_;
  wire g1003_n_spl_;
  wire g1004_n_spl_;
  wire g1004_p_spl_;
  wire g991_n_spl_;
  wire g1006_p_spl_;
  wire g991_p_spl_;
  wire g1006_n_spl_;
  wire g1007_n_spl_;
  wire g1007_p_spl_;
  wire g990_n_spl_;
  wire g1009_p_spl_;
  wire g990_p_spl_;
  wire g1009_n_spl_;
  wire g1010_n_spl_;
  wire g1010_p_spl_;
  wire g959_p_spl_;
  wire g958_n_spl_;
  wire G19_p_spl_;
  wire G19_p_spl_0;
  wire G19_p_spl_00;
  wire G19_p_spl_000;
  wire G19_p_spl_001;
  wire G19_p_spl_01;
  wire G19_p_spl_010;
  wire G19_p_spl_011;
  wire G19_p_spl_1;
  wire G19_p_spl_10;
  wire G19_p_spl_100;
  wire G19_p_spl_101;
  wire G19_p_spl_11;
  wire G19_p_spl_110;
  wire G19_p_spl_111;
  wire G19_n_spl_;
  wire G19_n_spl_0;
  wire G19_n_spl_00;
  wire G19_n_spl_000;
  wire G19_n_spl_001;
  wire G19_n_spl_01;
  wire G19_n_spl_010;
  wire G19_n_spl_011;
  wire G19_n_spl_1;
  wire G19_n_spl_10;
  wire G19_n_spl_100;
  wire G19_n_spl_101;
  wire G19_n_spl_11;
  wire G19_n_spl_110;
  wire G19_n_spl_111;
  wire ffc_290_n_spl_;
  wire ffc_290_p_spl_;
  wire ffc_130_p_spl_;
  wire ffc_130_p_spl_0;
  wire ffc_130_p_spl_00;
  wire ffc_130_p_spl_1;
  wire ffc_206_p_spl_;
  wire ffc_130_n_spl_;
  wire ffc_130_n_spl_0;
  wire ffc_206_n_spl_;
  wire ffc_292_p_spl_;
  wire ffc_292_n_spl_;
  wire g1018_n_spl_;
  wire g1019_p_spl_;
  wire g1018_p_spl_;
  wire g1019_n_spl_;
  wire g1020_n_spl_;
  wire g1020_p_spl_;
  wire g1017_n_spl_;
  wire g1022_p_spl_;
  wire g1017_p_spl_;
  wire g1022_n_spl_;
  wire ffc_129_p_spl_;
  wire ffc_129_p_spl_0;
  wire ffc_129_p_spl_1;
  wire ffc_224_p_spl_;
  wire ffc_224_p_spl_0;
  wire ffc_224_p_spl_00;
  wire ffc_224_p_spl_1;
  wire ffc_129_n_spl_;
  wire ffc_129_n_spl_0;
  wire ffc_224_n_spl_;
  wire ffc_224_n_spl_0;
  wire ffc_224_n_spl_00;
  wire ffc_224_n_spl_1;
  wire g1023_n_spl_;
  wire g1023_p_spl_;
  wire g1024_n_spl_;
  wire g1026_p_spl_;
  wire g1024_p_spl_;
  wire g1026_n_spl_;
  wire g1027_n_spl_;
  wire g1027_p_spl_;
  wire ffc_131_p_spl_;
  wire ffc_131_p_spl_0;
  wire ffc_131_p_spl_1;
  wire ffc_131_n_spl_;
  wire ffc_131_n_spl_0;
  wire g1030_n_spl_;
  wire g1031_n_spl_;
  wire g1030_p_spl_;
  wire g1031_p_spl_;
  wire g1032_n_spl_;
  wire g1032_p_spl_;
  wire g1029_n_spl_;
  wire g1034_p_spl_;
  wire g1029_p_spl_;
  wire g1034_n_spl_;
  wire g1035_n_spl_;
  wire g1035_p_spl_;
  wire g1028_n_spl_;
  wire g1037_p_spl_;
  wire g1028_p_spl_;
  wire g1037_n_spl_;
  wire g1038_n_spl_;
  wire g1038_p_spl_;
  wire g1039_n_spl_;
  wire g1041_p_spl_;
  wire g1039_p_spl_;
  wire g1041_n_spl_;
  wire g1042_n_spl_;
  wire g1042_p_spl_;
  wire g1045_n_spl_;
  wire g1046_n_spl_;
  wire g1045_p_spl_;
  wire g1046_p_spl_;
  wire g1047_n_spl_;
  wire g1047_p_spl_;
  wire g1044_n_spl_;
  wire g1049_p_spl_;
  wire g1044_p_spl_;
  wire g1049_n_spl_;
  wire g1050_n_spl_;
  wire g1050_p_spl_;
  wire g1043_n_spl_;
  wire g1052_p_spl_;
  wire g1043_p_spl_;
  wire g1052_n_spl_;
  wire ffc_288_n_spl_;
  wire ffc_288_p_spl_;
  wire ffc_127_p_spl_;
  wire ffc_127_p_spl_0;
  wire ffc_127_p_spl_00;
  wire ffc_127_p_spl_1;
  wire ffc_127_n_spl_;
  wire ffc_127_n_spl_0;
  wire ffc_294_p_spl_;
  wire ffc_294_n_spl_;
  wire g1055_n_spl_;
  wire g1056_p_spl_;
  wire g1055_p_spl_;
  wire g1056_n_spl_;
  wire g1057_n_spl_;
  wire g1057_p_spl_;
  wire g1054_n_spl_;
  wire g1059_p_spl_;
  wire g1054_p_spl_;
  wire g1059_n_spl_;
  wire ffc_126_p_spl_;
  wire ffc_126_p_spl_0;
  wire ffc_126_p_spl_1;
  wire ffc_126_n_spl_;
  wire ffc_126_n_spl_0;
  wire g1060_n_spl_;
  wire g1060_p_spl_;
  wire g1061_n_spl_;
  wire g1063_p_spl_;
  wire g1061_p_spl_;
  wire g1063_n_spl_;
  wire g1064_n_spl_;
  wire g1064_p_spl_;
  wire ffc_128_p_spl_;
  wire ffc_128_p_spl_0;
  wire ffc_128_p_spl_1;
  wire ffc_128_n_spl_;
  wire ffc_128_n_spl_0;
  wire g1069_n_spl_;
  wire g1070_p_spl_;
  wire g1069_p_spl_;
  wire g1070_n_spl_;
  wire g1071_n_spl_;
  wire g1071_p_spl_;
  wire g1068_n_spl_;
  wire g1073_p_spl_;
  wire g1068_p_spl_;
  wire g1073_n_spl_;
  wire g1074_n_spl_;
  wire g1074_p_spl_;
  wire g1067_n_spl_;
  wire g1076_p_spl_;
  wire g1067_p_spl_;
  wire g1076_n_spl_;
  wire g1077_n_spl_;
  wire g1077_p_spl_;
  wire g1066_n_spl_;
  wire g1079_p_spl_;
  wire g1066_p_spl_;
  wire g1079_n_spl_;
  wire g1080_n_spl_;
  wire g1080_p_spl_;
  wire g1065_n_spl_;
  wire g1082_p_spl_;
  wire g1065_p_spl_;
  wire g1082_n_spl_;
  wire g1083_n_spl_;
  wire g1083_p_spl_;
  wire g1084_n_spl_;
  wire g1086_p_spl_;
  wire g1084_p_spl_;
  wire g1086_n_spl_;
  wire g1087_n_spl_;
  wire g1087_p_spl_;
  wire g1092_n_spl_;
  wire g1094_p_spl_;
  wire g1092_p_spl_;
  wire g1094_n_spl_;
  wire g1095_n_spl_;
  wire g1095_p_spl_;
  wire g1091_n_spl_;
  wire g1097_p_spl_;
  wire g1091_p_spl_;
  wire g1097_n_spl_;
  wire g1098_n_spl_;
  wire g1098_p_spl_;
  wire g1090_n_spl_;
  wire g1100_p_spl_;
  wire g1090_p_spl_;
  wire g1100_n_spl_;
  wire g1101_n_spl_;
  wire g1101_p_spl_;
  wire g1089_n_spl_;
  wire g1103_p_spl_;
  wire g1089_p_spl_;
  wire g1103_n_spl_;
  wire g1104_n_spl_;
  wire g1104_p_spl_;
  wire g1088_n_spl_;
  wire g1106_p_spl_;
  wire g1088_p_spl_;
  wire g1106_n_spl_;
  wire ffc_123_p_spl_;
  wire ffc_123_p_spl_0;
  wire ffc_123_p_spl_00;
  wire ffc_123_p_spl_1;
  wire ffc_123_n_spl_;
  wire ffc_123_n_spl_0;
  wire ffc_123_n_spl_1;
  wire ffc_306_p_spl_;
  wire ffc_306_n_spl_;
  wire g1108_n_spl_;
  wire g1109_p_spl_;
  wire g1108_p_spl_;
  wire g1109_n_spl_;
  wire g1110_n_spl_;
  wire g1110_p_spl_;
  wire ffc_124_p_spl_;
  wire ffc_124_p_spl_0;
  wire ffc_124_p_spl_00;
  wire ffc_124_p_spl_1;
  wire ffc_124_n_spl_;
  wire ffc_124_n_spl_0;
  wire ffc_308_p_spl_;
  wire ffc_308_n_spl_;
  wire g1112_n_spl_;
  wire g1113_p_spl_;
  wire g1112_p_spl_;
  wire g1113_n_spl_;
  wire g1114_n_spl_;
  wire g1114_p_spl_;
  wire g1111_n_spl_;
  wire g1116_p_spl_;
  wire g1111_p_spl_;
  wire g1116_n_spl_;
  wire g1117_n_spl_;
  wire g1117_p_spl_;
  wire g1118_n_spl_;
  wire g1120_p_spl_;
  wire g1118_p_spl_;
  wire g1120_n_spl_;
  wire g1121_n_spl_;
  wire g1121_p_spl_;
  wire ffc_125_p_spl_;
  wire ffc_125_p_spl_0;
  wire ffc_125_p_spl_1;
  wire ffc_125_n_spl_;
  wire ffc_125_n_spl_0;
  wire g1126_n_spl_;
  wire g1127_p_spl_;
  wire g1126_p_spl_;
  wire g1127_n_spl_;
  wire g1128_n_spl_;
  wire g1128_p_spl_;
  wire g1125_n_spl_;
  wire g1130_p_spl_;
  wire g1125_p_spl_;
  wire g1130_n_spl_;
  wire g1131_n_spl_;
  wire g1131_p_spl_;
  wire g1124_n_spl_;
  wire g1133_p_spl_;
  wire g1124_p_spl_;
  wire g1133_n_spl_;
  wire g1134_n_spl_;
  wire g1134_p_spl_;
  wire g1123_n_spl_;
  wire g1136_p_spl_;
  wire g1123_p_spl_;
  wire g1136_n_spl_;
  wire g1137_n_spl_;
  wire g1137_p_spl_;
  wire g1122_n_spl_;
  wire g1139_p_spl_;
  wire g1122_p_spl_;
  wire g1139_n_spl_;
  wire g1140_n_spl_;
  wire g1140_p_spl_;
  wire g1141_n_spl_;
  wire g1143_p_spl_;
  wire g1141_p_spl_;
  wire g1143_n_spl_;
  wire g1144_n_spl_;
  wire g1144_p_spl_;
  wire g1149_n_spl_;
  wire g1151_p_spl_;
  wire g1149_p_spl_;
  wire g1151_n_spl_;
  wire g1152_n_spl_;
  wire g1152_p_spl_;
  wire g1148_n_spl_;
  wire g1154_p_spl_;
  wire g1148_p_spl_;
  wire g1154_n_spl_;
  wire g1155_n_spl_;
  wire g1155_p_spl_;
  wire g1147_n_spl_;
  wire g1157_p_spl_;
  wire g1147_p_spl_;
  wire g1157_n_spl_;
  wire g1158_n_spl_;
  wire g1158_p_spl_;
  wire g1146_n_spl_;
  wire g1160_p_spl_;
  wire g1146_p_spl_;
  wire g1160_n_spl_;
  wire g1161_n_spl_;
  wire g1161_p_spl_;
  wire g1145_n_spl_;
  wire g1163_p_spl_;
  wire g1145_p_spl_;
  wire g1163_n_spl_;
  wire ffc_120_p_spl_;
  wire ffc_120_p_spl_0;
  wire ffc_120_p_spl_00;
  wire ffc_120_p_spl_01;
  wire ffc_120_p_spl_1;
  wire ffc_120_n_spl_;
  wire ffc_120_n_spl_0;
  wire ffc_120_n_spl_00;
  wire ffc_120_n_spl_1;
  wire ffc_300_p_spl_;
  wire ffc_300_n_spl_;
  wire g1165_n_spl_;
  wire g1166_p_spl_;
  wire g1165_p_spl_;
  wire g1166_n_spl_;
  wire g1167_n_spl_;
  wire g1167_p_spl_;
  wire ffc_121_p_spl_;
  wire ffc_121_p_spl_0;
  wire ffc_121_p_spl_00;
  wire ffc_121_p_spl_01;
  wire ffc_121_p_spl_1;
  wire ffc_121_n_spl_;
  wire ffc_121_n_spl_0;
  wire ffc_121_n_spl_1;
  wire ffc_302_p_spl_;
  wire ffc_302_n_spl_;
  wire g1169_n_spl_;
  wire g1170_p_spl_;
  wire g1169_p_spl_;
  wire g1170_n_spl_;
  wire g1171_n_spl_;
  wire g1171_p_spl_;
  wire g1168_n_spl_;
  wire g1173_p_spl_;
  wire g1168_p_spl_;
  wire g1173_n_spl_;
  wire g1174_n_spl_;
  wire g1174_p_spl_;
  wire g1175_n_spl_;
  wire g1177_p_spl_;
  wire g1175_p_spl_;
  wire g1177_n_spl_;
  wire g1178_n_spl_;
  wire g1178_p_spl_;
  wire ffc_122_p_spl_;
  wire ffc_122_p_spl_0;
  wire ffc_122_p_spl_00;
  wire ffc_122_p_spl_1;
  wire ffc_122_n_spl_;
  wire ffc_122_n_spl_0;
  wire ffc_122_n_spl_1;
  wire ffc_304_p_spl_;
  wire ffc_304_n_spl_;
  wire g1182_n_spl_;
  wire g1183_p_spl_;
  wire g1182_p_spl_;
  wire g1183_n_spl_;
  wire g1184_n_spl_;
  wire g1184_p_spl_;
  wire g1181_n_spl_;
  wire g1186_p_spl_;
  wire g1181_p_spl_;
  wire g1186_n_spl_;
  wire g1187_n_spl_;
  wire g1187_p_spl_;
  wire g1180_n_spl_;
  wire g1189_p_spl_;
  wire g1180_p_spl_;
  wire g1189_n_spl_;
  wire g1190_n_spl_;
  wire g1190_p_spl_;
  wire g1179_n_spl_;
  wire g1192_p_spl_;
  wire g1179_p_spl_;
  wire g1192_n_spl_;
  wire g1193_n_spl_;
  wire g1193_p_spl_;
  wire g1194_n_spl_;
  wire g1196_p_spl_;
  wire g1194_p_spl_;
  wire g1196_n_spl_;
  wire g1197_n_spl_;
  wire g1197_p_spl_;
  wire g1202_n_spl_;
  wire g1204_p_spl_;
  wire g1202_p_spl_;
  wire g1204_n_spl_;
  wire g1205_n_spl_;
  wire g1205_p_spl_;
  wire g1201_n_spl_;
  wire g1207_p_spl_;
  wire g1201_p_spl_;
  wire g1207_n_spl_;
  wire g1208_n_spl_;
  wire g1208_p_spl_;
  wire g1200_n_spl_;
  wire g1210_p_spl_;
  wire g1200_p_spl_;
  wire g1210_n_spl_;
  wire g1211_n_spl_;
  wire g1211_p_spl_;
  wire g1199_n_spl_;
  wire g1213_p_spl_;
  wire g1199_p_spl_;
  wire g1213_n_spl_;
  wire g1214_n_spl_;
  wire g1214_p_spl_;
  wire g1198_n_spl_;
  wire g1216_p_spl_;
  wire g1198_p_spl_;
  wire g1216_n_spl_;
  wire g1217_n_spl_;
  wire g1217_p_spl_;
  wire g1218_n_spl_;
  wire g1220_p_spl_;
  wire g1218_p_spl_;
  wire g1220_n_spl_;
  wire g1221_n_spl_;
  wire g1221_p_spl_;
  wire g1226_n_spl_;
  wire g1228_p_spl_;
  wire g1226_p_spl_;
  wire g1228_n_spl_;
  wire g1229_n_spl_;
  wire g1229_p_spl_;
  wire g1225_n_spl_;
  wire g1231_p_spl_;
  wire g1225_p_spl_;
  wire g1231_n_spl_;
  wire g1232_n_spl_;
  wire g1232_p_spl_;
  wire g1224_n_spl_;
  wire g1234_p_spl_;
  wire g1224_p_spl_;
  wire g1234_n_spl_;
  wire g1235_n_spl_;
  wire g1235_p_spl_;
  wire g1223_n_spl_;
  wire g1237_p_spl_;
  wire g1223_p_spl_;
  wire g1237_n_spl_;
  wire g1238_n_spl_;
  wire g1238_p_spl_;
  wire g1222_n_spl_;
  wire g1240_p_spl_;
  wire g1222_p_spl_;
  wire g1240_n_spl_;
  wire g1012_p_spl_;
  wire g988_p_spl_;
  wire G3_p_spl_;
  wire G3_p_spl_0;
  wire G3_p_spl_00;
  wire G3_p_spl_01;
  wire G3_p_spl_1;
  wire G3_n_spl_;
  wire G3_n_spl_0;
  wire G3_n_spl_1;
  wire g1243_p_spl_;
  wire g1244_p_spl_;
  wire g1243_n_spl_;
  wire g1244_n_spl_;
  wire g1245_n_spl_;
  wire g1245_n_spl_0;
  wire g1245_p_spl_;
  wire g1245_p_spl_0;
  wire g989_n_spl_;
  wire g1247_n_spl_;
  wire g989_p_spl_;
  wire g989_p_spl_0;
  wire g1247_p_spl_;
  wire g1248_n_spl_;
  wire g1248_p_spl_;
  wire g987_p_spl_;
  wire g1257_n_spl_;
  wire g1259_p_spl_;
  wire g1257_p_spl_;
  wire g1259_n_spl_;
  wire g1260_n_spl_;
  wire g1260_p_spl_;
  wire g1256_n_spl_;
  wire g1262_p_spl_;
  wire g1256_p_spl_;
  wire g1262_n_spl_;
  wire g1263_n_spl_;
  wire g1263_p_spl_;
  wire g1255_n_spl_;
  wire g1265_p_spl_;
  wire g1255_p_spl_;
  wire g1265_n_spl_;
  wire g1266_n_spl_;
  wire g1266_p_spl_;
  wire g1254_n_spl_;
  wire g1268_p_spl_;
  wire g1254_p_spl_;
  wire g1268_n_spl_;
  wire g1269_n_spl_;
  wire g1269_p_spl_;
  wire g1253_n_spl_;
  wire g1271_p_spl_;
  wire g1253_p_spl_;
  wire g1271_n_spl_;
  wire g1272_n_spl_;
  wire g1272_p_spl_;
  wire g1252_n_spl_;
  wire g1274_p_spl_;
  wire g1252_p_spl_;
  wire g1274_n_spl_;
  wire g1275_n_spl_;
  wire g1275_p_spl_;
  wire ffc_336_n_spl_;
  wire ffc_353_p_spl_;
  wire ffc_336_p_spl_;
  wire ffc_353_n_spl_;
  wire g1279_n_spl_;
  wire g1279_p_spl_;
  wire ffc_337_n_spl_;
  wire ffc_354_p_spl_;
  wire ffc_337_p_spl_;
  wire ffc_354_n_spl_;
  wire g1281_n_spl_;
  wire g1281_p_spl_;
  wire g1280_n_spl_;
  wire g1283_p_spl_;
  wire g1280_p_spl_;
  wire g1283_n_spl_;
  wire ffc_190_p_spl_;
  wire ffc_190_p_spl_0;
  wire ffc_190_p_spl_1;
  wire ffc_190_n_spl_;
  wire ffc_190_n_spl_0;
  wire g1284_n_spl_;
  wire g1284_p_spl_;
  wire g1285_n_spl_;
  wire g1287_p_spl_;
  wire g1285_p_spl_;
  wire g1287_n_spl_;
  wire g1288_n_spl_;
  wire g1288_p_spl_;
  wire ffc_191_p_spl_;
  wire ffc_191_p_spl_0;
  wire ffc_191_n_spl_;
  wire ffc_191_n_spl_0;
  wire ffc_192_p_spl_;
  wire ffc_192_p_spl_0;
  wire ffc_192_p_spl_1;
  wire ffc_192_n_spl_;
  wire ffc_192_n_spl_0;
  wire ffc_338_n_spl_;
  wire ffc_340_n_spl_;
  wire ffc_338_p_spl_;
  wire ffc_340_p_spl_;
  wire g1293_n_spl_;
  wire g1293_p_spl_;
  wire g1292_n_spl_;
  wire g1295_p_spl_;
  wire g1292_p_spl_;
  wire g1295_n_spl_;
  wire g1296_n_spl_;
  wire g1296_p_spl_;
  wire g1291_n_spl_;
  wire g1298_p_spl_;
  wire g1291_p_spl_;
  wire g1298_n_spl_;
  wire g1299_n_spl_;
  wire g1299_p_spl_;
  wire g1290_n_spl_;
  wire g1301_p_spl_;
  wire g1290_p_spl_;
  wire g1301_n_spl_;
  wire g1302_n_spl_;
  wire g1302_p_spl_;
  wire g1289_n_spl_;
  wire g1304_p_spl_;
  wire g1289_p_spl_;
  wire g1304_n_spl_;
  wire g1305_n_spl_;
  wire g1305_p_spl_;
  wire g1306_n_spl_;
  wire g1308_p_spl_;
  wire g1306_p_spl_;
  wire g1308_n_spl_;
  wire g1309_n_spl_;
  wire g1309_p_spl_;
  wire ffc_193_p_spl_;
  wire ffc_193_p_spl_0;
  wire ffc_193_n_spl_;
  wire ffc_193_n_spl_0;
  wire g1314_n_spl_;
  wire g1315_n_spl_;
  wire g1314_p_spl_;
  wire g1315_p_spl_;
  wire g1316_n_spl_;
  wire g1316_p_spl_;
  wire g1313_n_spl_;
  wire g1318_p_spl_;
  wire g1313_p_spl_;
  wire g1318_n_spl_;
  wire g1319_n_spl_;
  wire g1319_p_spl_;
  wire g1312_n_spl_;
  wire g1321_p_spl_;
  wire g1312_p_spl_;
  wire g1321_n_spl_;
  wire g1322_n_spl_;
  wire g1322_p_spl_;
  wire g1311_n_spl_;
  wire g1324_p_spl_;
  wire g1311_p_spl_;
  wire g1324_n_spl_;
  wire g1325_n_spl_;
  wire g1325_p_spl_;
  wire g1310_n_spl_;
  wire g1327_p_spl_;
  wire g1310_p_spl_;
  wire g1327_n_spl_;
  wire ffc_333_n_spl_;
  wire ffc_350_p_spl_;
  wire ffc_333_p_spl_;
  wire ffc_350_n_spl_;
  wire g1329_n_spl_;
  wire g1329_p_spl_;
  wire ffc_334_n_spl_;
  wire ffc_351_p_spl_;
  wire ffc_334_p_spl_;
  wire ffc_351_n_spl_;
  wire g1331_n_spl_;
  wire g1331_p_spl_;
  wire g1330_n_spl_;
  wire g1333_p_spl_;
  wire g1330_p_spl_;
  wire g1333_n_spl_;
  wire ffc_187_p_spl_;
  wire ffc_187_p_spl_0;
  wire ffc_187_p_spl_00;
  wire ffc_187_p_spl_1;
  wire ffc_187_n_spl_;
  wire ffc_187_n_spl_0;
  wire ffc_187_n_spl_1;
  wire g1334_n_spl_;
  wire g1334_p_spl_;
  wire g1335_n_spl_;
  wire g1337_p_spl_;
  wire g1335_p_spl_;
  wire g1337_n_spl_;
  wire g1338_n_spl_;
  wire g1338_p_spl_;
  wire ffc_188_p_spl_;
  wire ffc_188_p_spl_0;
  wire ffc_188_p_spl_1;
  wire ffc_188_n_spl_;
  wire ffc_188_n_spl_0;
  wire ffc_188_n_spl_1;
  wire ffc_335_n_spl_;
  wire ffc_352_p_spl_;
  wire ffc_335_p_spl_;
  wire ffc_352_n_spl_;
  wire g1342_n_spl_;
  wire g1342_p_spl_;
  wire g1341_n_spl_;
  wire g1344_p_spl_;
  wire g1341_p_spl_;
  wire g1344_n_spl_;
  wire g1345_n_spl_;
  wire g1345_p_spl_;
  wire g1340_n_spl_;
  wire g1347_p_spl_;
  wire g1340_p_spl_;
  wire g1347_n_spl_;
  wire g1348_n_spl_;
  wire g1348_p_spl_;
  wire g1339_n_spl_;
  wire g1350_p_spl_;
  wire g1339_p_spl_;
  wire g1350_n_spl_;
  wire g1351_n_spl_;
  wire g1351_p_spl_;
  wire g1352_n_spl_;
  wire g1354_p_spl_;
  wire g1352_p_spl_;
  wire g1354_n_spl_;
  wire g1355_n_spl_;
  wire g1355_p_spl_;
  wire ffc_189_p_spl_;
  wire ffc_189_p_spl_0;
  wire ffc_189_p_spl_1;
  wire ffc_189_n_spl_;
  wire ffc_189_n_spl_0;
  wire g1360_n_spl_;
  wire g1362_p_spl_;
  wire g1360_p_spl_;
  wire g1362_n_spl_;
  wire g1363_n_spl_;
  wire g1363_p_spl_;
  wire g1359_n_spl_;
  wire g1365_p_spl_;
  wire g1359_p_spl_;
  wire g1365_n_spl_;
  wire g1366_n_spl_;
  wire g1366_p_spl_;
  wire g1358_n_spl_;
  wire g1368_p_spl_;
  wire g1358_p_spl_;
  wire g1368_n_spl_;
  wire g1369_n_spl_;
  wire g1369_p_spl_;
  wire g1357_n_spl_;
  wire g1371_p_spl_;
  wire g1357_p_spl_;
  wire g1371_n_spl_;
  wire g1372_n_spl_;
  wire g1372_p_spl_;
  wire g1356_n_spl_;
  wire g1374_p_spl_;
  wire g1356_p_spl_;
  wire g1374_n_spl_;
  wire g1375_n_spl_;
  wire g1375_p_spl_;
  wire g1376_n_spl_;
  wire g1378_p_spl_;
  wire g1376_p_spl_;
  wire g1378_n_spl_;
  wire g1379_n_spl_;
  wire g1379_p_spl_;
  wire g1384_n_spl_;
  wire g1386_p_spl_;
  wire g1384_p_spl_;
  wire g1386_n_spl_;
  wire g1387_n_spl_;
  wire g1387_p_spl_;
  wire g1383_n_spl_;
  wire g1389_p_spl_;
  wire g1383_p_spl_;
  wire g1389_n_spl_;
  wire g1390_n_spl_;
  wire g1390_p_spl_;
  wire g1382_n_spl_;
  wire g1392_p_spl_;
  wire g1382_p_spl_;
  wire g1392_n_spl_;
  wire g1393_n_spl_;
  wire g1393_p_spl_;
  wire g1381_n_spl_;
  wire g1395_p_spl_;
  wire g1381_p_spl_;
  wire g1395_n_spl_;
  wire g1396_n_spl_;
  wire g1396_p_spl_;
  wire g1380_n_spl_;
  wire g1398_p_spl_;
  wire g1380_p_spl_;
  wire g1398_n_spl_;
  wire g1250_p_spl_;
  wire g1016_p_spl_;
  wire ffc_21_n_spl_;
  wire ffc_21_n_spl_0;
  wire ffc_21_n_spl_00;
  wire ffc_21_n_spl_1;
  wire ffc_12_n_spl_;
  wire ffc_12_n_spl_0;
  wire ffc_12_n_spl_00;
  wire ffc_12_n_spl_000;
  wire ffc_12_n_spl_001;
  wire ffc_12_n_spl_01;
  wire ffc_12_n_spl_010;
  wire ffc_12_n_spl_1;
  wire ffc_12_n_spl_10;
  wire ffc_12_n_spl_11;
  wire G20_n_spl_;
  wire G20_n_spl_0;
  wire G20_n_spl_00;
  wire G20_n_spl_000;
  wire G20_n_spl_001;
  wire G20_n_spl_01;
  wire G20_n_spl_010;
  wire G20_n_spl_011;
  wire G20_n_spl_1;
  wire G20_n_spl_10;
  wire G20_n_spl_100;
  wire G20_n_spl_101;
  wire G20_n_spl_11;
  wire G20_n_spl_110;
  wire g946_n_spl_;
  wire g1404_n_spl_;
  wire g1406_p_spl_;
  wire g934_n_spl_;
  wire g1409_n_spl_;
  wire g1411_p_spl_;
  wire g922_n_spl_;
  wire g1414_n_spl_;
  wire g1416_p_spl_;
  wire g919_n_spl_;
  wire g1419_n_spl_;
  wire g1421_p_spl_;
  wire g915_n_spl_;
  wire g1424_n_spl_;
  wire g1426_p_spl_;
  wire g911_n_spl_;
  wire g1429_n_spl_;
  wire g1431_p_spl_;
  wire g1013_n_spl_;
  wire g1015_p_spl_;
  wire ffc_21_p_spl_;
  wire ffc_21_p_spl_0;
  wire ffc_21_p_spl_00;
  wire ffc_21_p_spl_1;
  wire g1241_n_spl_;
  wire g1164_n_spl_;
  wire g1107_n_spl_;
  wire g1053_n_spl_;
  wire g1459_n_spl_;
  wire g1461_p_spl_;
  wire g1459_p_spl_;
  wire g1461_n_spl_;
  wire g1462_n_spl_;
  wire g1462_p_spl_;
  wire g1458_n_spl_;
  wire g1464_p_spl_;
  wire g1458_p_spl_;
  wire g1464_n_spl_;
  wire g1465_n_spl_;
  wire g1465_p_spl_;
  wire g1457_n_spl_;
  wire g1467_p_spl_;
  wire g1457_p_spl_;
  wire g1467_n_spl_;
  wire g1468_n_spl_;
  wire g1468_p_spl_;
  wire g1456_n_spl_;
  wire g1470_p_spl_;
  wire g1456_p_spl_;
  wire g1470_n_spl_;
  wire g1471_n_spl_;
  wire g1471_p_spl_;
  wire g1455_n_spl_;
  wire g1473_p_spl_;
  wire g1454_n_spl_;
  wire g1476_p_spl_;
  wire g1480_n_spl_;
  wire g1482_p_spl_;
  wire g1480_p_spl_;
  wire g1482_n_spl_;
  wire g1483_n_spl_;
  wire g1479_n_spl_;
  wire g1485_p_spl_;
  wire g1479_p_spl_;
  wire g1485_n_spl_;
  wire g1486_n_spl_;
  wire g1492_n_spl_;
  wire g1494_p_spl_;
  wire g1492_p_spl_;
  wire g1494_n_spl_;
  wire g1495_n_spl_;
  wire g1491_n_spl_;
  wire g1497_p_spl_;
  wire g1491_p_spl_;
  wire g1497_n_spl_;
  wire g1498_n_spl_;
  wire g1504_n_spl_;
  wire g1506_p_spl_;
  wire g1504_p_spl_;
  wire g1506_n_spl_;
  wire g1507_n_spl_;
  wire g1503_n_spl_;
  wire g1509_p_spl_;
  wire g1503_p_spl_;
  wire g1509_n_spl_;
  wire g1510_n_spl_;
  wire g1278_n_spl_;
  wire ffc_12_p_spl_;
  wire ffc_12_p_spl_0;
  wire ffc_12_p_spl_00;
  wire ffc_12_p_spl_000;
  wire ffc_12_p_spl_001;
  wire ffc_12_p_spl_01;
  wire ffc_12_p_spl_1;
  wire ffc_12_p_spl_10;
  wire ffc_12_p_spl_11;
  wire g1399_n_spl_;
  wire g1328_n_spl_;
  wire g1526_n_spl_;
  wire g1527_n_spl_;
  wire g1526_p_spl_;
  wire g1527_p_spl_;
  wire g1528_p_spl_;
  wire g1525_n_spl_;
  wire g1530_p_spl_;
  wire g1525_p_spl_;
  wire g1530_n_spl_;
  wire g1531_p_spl_;
  wire g1537_n_spl_;
  wire g1539_p_spl_;
  wire g1537_p_spl_;
  wire g1539_n_spl_;
  wire g1540_p_spl_;
  wire g1536_n_spl_;
  wire g1542_p_spl_;
  wire g1536_p_spl_;
  wire g1542_n_spl_;
  wire g1543_p_spl_;
  wire g1242_p_spl_;
  wire ffc_181_p_spl_;
  wire ffc_181_p_spl_0;
  wire ffc_181_p_spl_00;
  wire ffc_181_p_spl_1;
  wire ffc_181_n_spl_;
  wire ffc_181_n_spl_0;
  wire ffc_181_n_spl_1;
  wire ffc_328_n_spl_;
  wire ffc_345_p_spl_;
  wire ffc_328_p_spl_;
  wire ffc_345_n_spl_;
  wire g1554_n_spl_;
  wire g1554_p_spl_;
  wire g1553_n_spl_;
  wire g1556_p_spl_;
  wire g1553_p_spl_;
  wire g1556_n_spl_;
  wire g1557_n_spl_;
  wire g1557_p_spl_;
  wire g1552_n_spl_;
  wire g1559_p_spl_;
  wire g1552_p_spl_;
  wire g1559_n_spl_;
  wire g1560_n_spl_;
  wire g1560_p_spl_;
  wire g1551_n_spl_;
  wire g1562_p_spl_;
  wire g1551_p_spl_;
  wire g1562_n_spl_;
  wire g1563_n_spl_;
  wire g1563_p_spl_;
  wire g1550_n_spl_;
  wire g1565_p_spl_;
  wire g1550_p_spl_;
  wire g1565_n_spl_;
  wire g1566_n_spl_;
  wire g1566_p_spl_;
  wire g1549_n_spl_;
  wire g1568_p_spl_;
  wire g1549_p_spl_;
  wire g1568_n_spl_;
  wire g1569_n_spl_;
  wire g1569_p_spl_;
  wire g1548_n_spl_;
  wire g1571_p_spl_;
  wire g1548_p_spl_;
  wire g1571_n_spl_;
  wire g1572_n_spl_;
  wire g1572_p_spl_;
  wire g1547_n_spl_;
  wire g1574_p_spl_;
  wire g1400_p_spl_;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_00;
  wire G4_p_spl_01;
  wire G4_p_spl_1;
  wire G4_n_spl_;
  wire G4_n_spl_0;
  wire G4_n_spl_1;
  wire g1580_p_spl_;
  wire g1581_p_spl_;
  wire g1580_n_spl_;
  wire g1581_n_spl_;
  wire g1582_n_spl_;
  wire g1582_n_spl_0;
  wire g1582_p_spl_;
  wire g1582_p_spl_0;
  wire g1584_n_spl_;
  wire g1584_p_spl_;
  wire g1585_n_spl_;
  wire g1585_p_spl_;
  wire g1579_n_spl_;
  wire g1587_p_spl_;
  wire g1579_p_spl_;
  wire g1587_n_spl_;
  wire g1588_n_spl_;
  wire g1588_p_spl_;
  wire g1578_n_spl_;
  wire g1590_p_spl_;
  wire g1603_n_spl_;
  wire g1605_p_spl_;
  wire g1603_p_spl_;
  wire g1605_n_spl_;
  wire g1606_n_spl_;
  wire g1606_p_spl_;
  wire g1602_n_spl_;
  wire g1608_p_spl_;
  wire g1602_p_spl_;
  wire g1608_n_spl_;
  wire g1609_n_spl_;
  wire g1609_p_spl_;
  wire g1601_n_spl_;
  wire g1611_p_spl_;
  wire g1601_p_spl_;
  wire g1611_n_spl_;
  wire g1612_n_spl_;
  wire g1616_n_spl_;
  wire g1618_n_spl_;
  wire g1620_p_spl_;
  wire g1618_p_spl_;
  wire g1620_n_spl_;
  wire g1621_n_spl_;
  wire g1625_n_spl_;
  wire g1477_p_spl_;
  wire g1401_n_spl_;
  wire g1515_p_spl_;
  wire g1402_n_spl_;
  wire g1577_p_spl_;
  wire g1403_n_spl_;
  wire g1593_p_spl_;
  wire g1438_n_spl_;
  wire g1442_n_spl_;
  wire g1446_n_spl_;
  wire g1450_n_spl_;
  wire g1453_n_spl_;
  wire g1489_n_spl_;
  wire g1501_n_spl_;
  wire g1513_n_spl_;
  wire g1630_p_spl_;
  wire ffc_182_p_spl_;
  wire ffc_182_p_spl_0;
  wire ffc_182_p_spl_00;
  wire ffc_182_p_spl_1;
  wire ffc_182_n_spl_;
  wire ffc_182_n_spl_0;
  wire ffc_182_n_spl_1;
  wire ffc_329_n_spl_;
  wire ffc_346_p_spl_;
  wire ffc_329_p_spl_;
  wire ffc_346_n_spl_;
  wire g1661_n_spl_;
  wire g1661_p_spl_;
  wire g1660_n_spl_;
  wire g1663_p_spl_;
  wire g1660_p_spl_;
  wire g1663_n_spl_;
  wire g1664_n_spl_;
  wire g1664_p_spl_;
  wire g1659_n_spl_;
  wire g1666_p_spl_;
  wire g1659_p_spl_;
  wire g1666_n_spl_;
  wire g1667_n_spl_;
  wire g1667_p_spl_;
  wire g1658_n_spl_;
  wire g1669_p_spl_;
  wire g1658_p_spl_;
  wire g1669_n_spl_;
  wire g1670_n_spl_;
  wire g1670_p_spl_;
  wire g1657_n_spl_;
  wire g1672_p_spl_;
  wire g1657_p_spl_;
  wire g1672_n_spl_;
  wire g1673_n_spl_;
  wire g1673_p_spl_;
  wire g1656_n_spl_;
  wire g1675_p_spl_;
  wire g1656_p_spl_;
  wire g1675_n_spl_;
  wire g1676_n_spl_;
  wire g1676_p_spl_;
  wire g1655_n_spl_;
  wire g1678_p_spl_;
  wire g1655_p_spl_;
  wire g1678_n_spl_;
  wire g1679_n_spl_;
  wire g1679_p_spl_;
  wire g1654_n_spl_;
  wire g1681_p_spl_;
  wire g1654_p_spl_;
  wire g1681_n_spl_;
  wire g1682_n_spl_;
  wire g1685_n_spl_;
  wire g1546_n_spl_;
  wire g1688_n_spl_;
  wire g1690_p_spl_;
  wire g1534_n_spl_;
  wire g1693_n_spl_;
  wire g1695_p_spl_;
  wire g1698_n_spl_;
  wire g1699_n_spl_;
  wire g1523_n_spl_;
  wire g1702_n_spl_;
  wire g1704_p_spl_;
  wire ffc_183_p_spl_;
  wire ffc_183_p_spl_0;
  wire ffc_183_p_spl_00;
  wire ffc_183_p_spl_1;
  wire ffc_183_n_spl_;
  wire ffc_183_n_spl_0;
  wire ffc_183_n_spl_1;
  wire ffc_330_n_spl_;
  wire ffc_347_p_spl_;
  wire ffc_330_p_spl_;
  wire ffc_347_n_spl_;
  wire g1714_n_spl_;
  wire g1714_p_spl_;
  wire g1713_n_spl_;
  wire g1716_p_spl_;
  wire g1713_p_spl_;
  wire g1716_n_spl_;
  wire g1717_n_spl_;
  wire g1717_p_spl_;
  wire g1712_n_spl_;
  wire g1719_p_spl_;
  wire g1712_p_spl_;
  wire g1719_n_spl_;
  wire g1720_n_spl_;
  wire g1720_p_spl_;
  wire g1711_n_spl_;
  wire g1722_p_spl_;
  wire g1711_p_spl_;
  wire g1722_n_spl_;
  wire g1723_n_spl_;
  wire g1723_p_spl_;
  wire g1710_n_spl_;
  wire g1725_p_spl_;
  wire g1710_p_spl_;
  wire g1725_n_spl_;
  wire g1726_n_spl_;
  wire g1726_p_spl_;
  wire g1709_n_spl_;
  wire g1728_p_spl_;
  wire g1709_p_spl_;
  wire g1728_n_spl_;
  wire g1729_n_spl_;
  wire g1729_p_spl_;
  wire g1708_n_spl_;
  wire g1731_p_spl_;
  wire g1708_p_spl_;
  wire g1731_n_spl_;
  wire g1732_n_spl_;
  wire g1732_p_spl_;
  wire g1707_n_spl_;
  wire g1734_p_spl_;
  wire g1707_p_spl_;
  wire g1734_n_spl_;
  wire g1735_p_spl_;
  wire g1739_p_spl_;
  wire ffc_184_p_spl_;
  wire ffc_184_p_spl_0;
  wire ffc_184_p_spl_00;
  wire ffc_184_p_spl_1;
  wire ffc_184_n_spl_;
  wire ffc_184_n_spl_0;
  wire ffc_184_n_spl_1;
  wire ffc_331_n_spl_;
  wire ffc_348_p_spl_;
  wire ffc_331_p_spl_;
  wire ffc_348_n_spl_;
  wire g1749_n_spl_;
  wire g1749_p_spl_;
  wire g1748_n_spl_;
  wire g1751_p_spl_;
  wire g1748_p_spl_;
  wire g1751_n_spl_;
  wire g1752_n_spl_;
  wire g1752_p_spl_;
  wire g1747_n_spl_;
  wire g1754_p_spl_;
  wire g1747_p_spl_;
  wire g1754_n_spl_;
  wire g1755_n_spl_;
  wire g1755_p_spl_;
  wire g1746_n_spl_;
  wire g1757_p_spl_;
  wire g1746_p_spl_;
  wire g1757_n_spl_;
  wire g1758_n_spl_;
  wire g1758_p_spl_;
  wire g1745_n_spl_;
  wire g1760_p_spl_;
  wire g1745_p_spl_;
  wire g1760_n_spl_;
  wire g1761_n_spl_;
  wire g1761_p_spl_;
  wire g1744_n_spl_;
  wire g1763_p_spl_;
  wire g1744_p_spl_;
  wire g1763_n_spl_;
  wire g1764_n_spl_;
  wire g1764_p_spl_;
  wire g1743_n_spl_;
  wire g1766_p_spl_;
  wire g1743_p_spl_;
  wire g1766_n_spl_;
  wire g1767_n_spl_;
  wire g1767_p_spl_;
  wire g1742_n_spl_;
  wire g1769_p_spl_;
  wire g1742_p_spl_;
  wire g1769_n_spl_;
  wire g1770_p_spl_;
  wire g1741_n_spl_;
  wire g1772_p_spl_;
  wire g1740_n_spl_;
  wire g1775_p_spl_;
  wire ffc_185_p_spl_;
  wire ffc_185_p_spl_0;
  wire ffc_185_p_spl_00;
  wire ffc_185_p_spl_1;
  wire ffc_185_n_spl_;
  wire ffc_185_n_spl_0;
  wire ffc_185_n_spl_1;
  wire ffc_332_n_spl_;
  wire ffc_349_p_spl_;
  wire ffc_332_p_spl_;
  wire ffc_349_n_spl_;
  wire g1787_n_spl_;
  wire g1787_p_spl_;
  wire g1786_n_spl_;
  wire g1789_p_spl_;
  wire g1786_p_spl_;
  wire g1789_n_spl_;
  wire g1790_n_spl_;
  wire g1790_p_spl_;
  wire g1785_n_spl_;
  wire g1792_p_spl_;
  wire g1785_p_spl_;
  wire g1792_n_spl_;
  wire g1793_n_spl_;
  wire g1793_p_spl_;
  wire g1784_n_spl_;
  wire g1795_p_spl_;
  wire g1784_p_spl_;
  wire g1795_n_spl_;
  wire g1796_n_spl_;
  wire g1796_p_spl_;
  wire g1783_n_spl_;
  wire g1798_p_spl_;
  wire g1783_p_spl_;
  wire g1798_n_spl_;
  wire g1799_n_spl_;
  wire g1799_p_spl_;
  wire g1782_n_spl_;
  wire g1801_p_spl_;
  wire g1782_p_spl_;
  wire g1801_n_spl_;
  wire g1802_n_spl_;
  wire g1802_p_spl_;
  wire g1781_n_spl_;
  wire g1804_p_spl_;
  wire g1781_p_spl_;
  wire g1804_n_spl_;
  wire g1805_n_spl_;
  wire g1805_p_spl_;
  wire g1780_n_spl_;
  wire g1807_p_spl_;
  wire g1780_p_spl_;
  wire g1807_n_spl_;
  wire g1808_p_spl_;
  wire g1779_n_spl_;
  wire g1810_p_spl_;
  wire g1778_n_spl_;
  wire g1813_p_spl_;
  wire ffc_186_p_spl_;
  wire ffc_186_p_spl_0;
  wire ffc_186_p_spl_00;
  wire ffc_186_p_spl_1;
  wire ffc_186_n_spl_;
  wire ffc_186_n_spl_0;
  wire ffc_186_n_spl_1;
  wire g1824_n_spl_;
  wire g1826_p_spl_;
  wire g1824_p_spl_;
  wire g1826_n_spl_;
  wire g1827_n_spl_;
  wire g1827_p_spl_;
  wire g1823_n_spl_;
  wire g1829_p_spl_;
  wire g1823_p_spl_;
  wire g1829_n_spl_;
  wire g1830_n_spl_;
  wire g1830_p_spl_;
  wire g1822_n_spl_;
  wire g1832_p_spl_;
  wire g1822_p_spl_;
  wire g1832_n_spl_;
  wire g1833_n_spl_;
  wire g1833_p_spl_;
  wire g1821_n_spl_;
  wire g1835_p_spl_;
  wire g1821_p_spl_;
  wire g1835_n_spl_;
  wire g1836_n_spl_;
  wire g1836_p_spl_;
  wire g1820_n_spl_;
  wire g1838_p_spl_;
  wire g1820_p_spl_;
  wire g1838_n_spl_;
  wire g1839_n_spl_;
  wire g1839_p_spl_;
  wire g1819_n_spl_;
  wire g1841_p_spl_;
  wire g1819_p_spl_;
  wire g1841_n_spl_;
  wire g1842_n_spl_;
  wire g1842_p_spl_;
  wire g1818_n_spl_;
  wire g1844_p_spl_;
  wire g1818_p_spl_;
  wire g1844_n_spl_;
  wire g1845_p_spl_;
  wire g1817_n_spl_;
  wire g1847_p_spl_;
  wire g1816_n_spl_;
  wire g1850_p_spl_;
  wire g1859_n_spl_;
  wire g1861_p_spl_;
  wire g1859_p_spl_;
  wire g1861_n_spl_;
  wire g1862_n_spl_;
  wire g1862_p_spl_;
  wire g1858_n_spl_;
  wire g1864_p_spl_;
  wire g1858_p_spl_;
  wire g1864_n_spl_;
  wire g1865_n_spl_;
  wire g1865_p_spl_;
  wire g1857_n_spl_;
  wire g1867_p_spl_;
  wire g1857_p_spl_;
  wire g1867_n_spl_;
  wire g1868_n_spl_;
  wire g1868_p_spl_;
  wire g1856_n_spl_;
  wire g1870_p_spl_;
  wire g1856_p_spl_;
  wire g1870_n_spl_;
  wire g1871_n_spl_;
  wire g1871_p_spl_;
  wire g1855_n_spl_;
  wire g1873_p_spl_;
  wire g1855_p_spl_;
  wire g1873_n_spl_;
  wire g1874_p_spl_;
  wire g1854_n_spl_;
  wire g1876_p_spl_;
  wire g1853_n_spl_;
  wire g1879_p_spl_;
  wire g1886_n_spl_;
  wire g1888_p_spl_;
  wire g1886_p_spl_;
  wire g1888_n_spl_;
  wire g1889_n_spl_;
  wire g1889_p_spl_;
  wire g1885_n_spl_;
  wire g1891_p_spl_;
  wire g1885_p_spl_;
  wire g1891_n_spl_;
  wire g1892_n_spl_;
  wire g1892_p_spl_;
  wire g1884_n_spl_;
  wire g1894_p_spl_;
  wire g1884_p_spl_;
  wire g1894_n_spl_;
  wire g1895_p_spl_;
  wire g1883_n_spl_;
  wire g1897_p_spl_;
  wire g1882_n_spl_;
  wire g1900_p_spl_;
  wire g1905_n_spl_;
  wire g1907_p_spl_;
  wire g1905_p_spl_;
  wire g1907_n_spl_;
  wire g1908_p_spl_;
  wire g1904_n_spl_;
  wire g1910_p_spl_;
  wire g1903_n_spl_;
  wire g1913_p_spl_;
  wire g1519_n_spl_;
  wire g1916_n_spl_;
  wire g1918_p_spl_;
  wire g1921_p_spl_;
  wire g1923_n_spl_;
  wire G5_p_spl_;
  wire G5_p_spl_0;
  wire G5_p_spl_00;
  wire G5_p_spl_01;
  wire G5_p_spl_1;
  wire G5_n_spl_;
  wire G5_n_spl_0;
  wire G5_n_spl_1;
  wire g1926_p_spl_;
  wire g1927_p_spl_;
  wire g1926_n_spl_;
  wire g1927_n_spl_;
  wire g1928_n_spl_;
  wire g1928_n_spl_0;
  wire g1928_p_spl_;
  wire g1928_p_spl_0;
  wire g1930_n_spl_;
  wire g1930_p_spl_;
  wire g1931_n_spl_;
  wire g1931_p_spl_;
  wire g1932_n_spl_;
  wire g1934_p_spl_;
  wire g1932_p_spl_;
  wire g1934_n_spl_;
  wire g1935_n_spl_;
  wire g1935_p_spl_;
  wire G6_p_spl_;
  wire G6_p_spl_0;
  wire G6_p_spl_00;
  wire G6_p_spl_01;
  wire G6_p_spl_1;
  wire G6_n_spl_;
  wire G6_n_spl_0;
  wire G6_n_spl_1;
  wire g1938_p_spl_;
  wire g1939_p_spl_;
  wire g1938_n_spl_;
  wire g1939_n_spl_;
  wire g1940_n_spl_;
  wire g1940_n_spl_0;
  wire g1940_p_spl_;
  wire g1940_p_spl_0;
  wire g1942_n_spl_;
  wire g1942_p_spl_;
  wire g1943_n_spl_;
  wire g1943_p_spl_;
  wire g1937_n_spl_;
  wire g1945_p_spl_;
  wire g1937_p_spl_;
  wire g1945_n_spl_;
  wire g1946_n_spl_;
  wire g1946_p_spl_;
  wire g1936_n_spl_;
  wire g1948_p_spl_;
  wire g1936_p_spl_;
  wire g1948_n_spl_;
  wire G20_p_spl_;
  wire G20_p_spl_0;
  wire G20_p_spl_00;
  wire G20_p_spl_000;
  wire G20_p_spl_001;
  wire G20_p_spl_01;
  wire G20_p_spl_010;
  wire G20_p_spl_011;
  wire G20_p_spl_1;
  wire G20_p_spl_10;
  wire G20_p_spl_100;
  wire G20_p_spl_101;
  wire G20_p_spl_11;
  wire G20_p_spl_110;
  wire g1949_n_spl_;
  wire g1949_p_spl_;
  wire g1950_n_spl_;
  wire g1952_p_spl_;
  wire g1950_p_spl_;
  wire g1952_n_spl_;
  wire g1953_n_spl_;
  wire g1953_p_spl_;
  wire G7_p_spl_;
  wire G7_p_spl_0;
  wire G7_p_spl_00;
  wire G7_p_spl_01;
  wire G7_p_spl_1;
  wire G7_n_spl_;
  wire G7_n_spl_0;
  wire G7_n_spl_1;
  wire g1958_p_spl_;
  wire g1959_p_spl_;
  wire g1958_n_spl_;
  wire g1959_n_spl_;
  wire g1960_n_spl_;
  wire g1960_n_spl_0;
  wire g1960_p_spl_;
  wire g1960_p_spl_0;
  wire g1962_n_spl_;
  wire g1962_p_spl_;
  wire g1963_n_spl_;
  wire g1963_p_spl_;
  wire g1957_n_spl_;
  wire g1965_p_spl_;
  wire g1957_p_spl_;
  wire g1965_n_spl_;
  wire g1966_n_spl_;
  wire g1966_p_spl_;
  wire g1956_n_spl_;
  wire g1968_p_spl_;
  wire g1956_p_spl_;
  wire g1968_n_spl_;
  wire g1969_n_spl_;
  wire g1969_p_spl_;
  wire g1955_n_spl_;
  wire g1971_p_spl_;
  wire g1955_p_spl_;
  wire g1971_n_spl_;
  wire g1972_n_spl_;
  wire g1972_p_spl_;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire G8_p_spl_00;
  wire G8_p_spl_01;
  wire G8_p_spl_1;
  wire G8_n_spl_;
  wire G8_n_spl_0;
  wire G8_n_spl_1;
  wire g1980_p_spl_;
  wire g1981_p_spl_;
  wire g1980_n_spl_;
  wire g1981_n_spl_;
  wire g1982_n_spl_;
  wire g1982_n_spl_0;
  wire g1982_p_spl_;
  wire g1982_p_spl_0;
  wire g1984_n_spl_;
  wire g1984_p_spl_;
  wire g1985_n_spl_;
  wire g1985_p_spl_;
  wire g1979_n_spl_;
  wire g1987_p_spl_;
  wire g1979_p_spl_;
  wire g1987_n_spl_;
  wire g1988_n_spl_;
  wire g1988_p_spl_;
  wire g1978_n_spl_;
  wire g1990_p_spl_;
  wire g1978_p_spl_;
  wire g1990_n_spl_;
  wire g1991_n_spl_;
  wire g1991_p_spl_;
  wire g1977_n_spl_;
  wire g1993_p_spl_;
  wire g1977_p_spl_;
  wire g1993_n_spl_;
  wire g1994_n_spl_;
  wire g1994_p_spl_;
  wire G9_p_spl_;
  wire G9_p_spl_0;
  wire G9_p_spl_00;
  wire G9_p_spl_01;
  wire G9_p_spl_1;
  wire G9_n_spl_;
  wire G9_n_spl_0;
  wire G9_n_spl_1;
  wire g2002_p_spl_;
  wire g2003_p_spl_;
  wire g2002_n_spl_;
  wire g2003_n_spl_;
  wire g2004_n_spl_;
  wire g2004_n_spl_0;
  wire g2004_p_spl_;
  wire g2004_p_spl_0;
  wire g2006_n_spl_;
  wire g2006_p_spl_;
  wire g2007_n_spl_;
  wire g2007_p_spl_;
  wire g2001_n_spl_;
  wire g2009_p_spl_;
  wire g2001_p_spl_;
  wire g2009_n_spl_;
  wire g2010_n_spl_;
  wire g2010_p_spl_;
  wire g2000_n_spl_;
  wire g2012_p_spl_;
  wire g2000_p_spl_;
  wire g2012_n_spl_;
  wire g2013_n_spl_;
  wire g2013_p_spl_;
  wire g1999_n_spl_;
  wire g2015_p_spl_;
  wire g1999_p_spl_;
  wire g2015_n_spl_;
  wire g2016_n_spl_;
  wire g2016_p_spl_;
  wire G10_p_spl_;
  wire G10_p_spl_0;
  wire G10_p_spl_00;
  wire G10_p_spl_01;
  wire G10_p_spl_1;
  wire G10_n_spl_;
  wire G10_n_spl_0;
  wire G10_n_spl_1;
  wire g2024_p_spl_;
  wire g2025_p_spl_;
  wire g2024_n_spl_;
  wire g2025_n_spl_;
  wire g2026_n_spl_;
  wire g2026_n_spl_0;
  wire g2026_p_spl_;
  wire g2026_p_spl_0;
  wire g2028_n_spl_;
  wire g2028_p_spl_;
  wire g2029_n_spl_;
  wire g2029_p_spl_;
  wire g2023_n_spl_;
  wire g2031_p_spl_;
  wire g2023_p_spl_;
  wire g2031_n_spl_;
  wire g2032_n_spl_;
  wire g2032_p_spl_;
  wire g2022_n_spl_;
  wire g2034_p_spl_;
  wire g2022_p_spl_;
  wire g2034_n_spl_;
  wire g2035_n_spl_;
  wire g2035_p_spl_;
  wire g2021_n_spl_;
  wire g2037_p_spl_;
  wire g2021_p_spl_;
  wire g2037_n_spl_;
  wire g2038_n_spl_;
  wire g2038_p_spl_;
  wire G11_p_spl_;
  wire G11_p_spl_0;
  wire G11_p_spl_00;
  wire G11_p_spl_01;
  wire G11_p_spl_1;
  wire G11_n_spl_;
  wire G11_n_spl_0;
  wire G11_n_spl_1;
  wire g2046_p_spl_;
  wire g2047_p_spl_;
  wire g2046_n_spl_;
  wire g2047_n_spl_;
  wire g2048_n_spl_;
  wire g2048_n_spl_0;
  wire g2048_p_spl_;
  wire g2048_p_spl_0;
  wire g2050_n_spl_;
  wire g2050_p_spl_;
  wire g2051_n_spl_;
  wire g2051_p_spl_;
  wire g2045_n_spl_;
  wire g2053_p_spl_;
  wire g2045_p_spl_;
  wire g2053_n_spl_;
  wire g2054_n_spl_;
  wire g2054_p_spl_;
  wire g2044_n_spl_;
  wire g2056_p_spl_;
  wire g2044_p_spl_;
  wire g2056_n_spl_;
  wire g2057_n_spl_;
  wire g2057_p_spl_;
  wire g2043_n_spl_;
  wire g2059_p_spl_;
  wire g2043_p_spl_;
  wire g2059_n_spl_;
  wire g2060_n_spl_;
  wire g2060_p_spl_;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire G12_p_spl_00;
  wire G12_p_spl_01;
  wire G12_p_spl_1;
  wire G12_n_spl_;
  wire G12_n_spl_0;
  wire G12_n_spl_1;
  wire g2068_p_spl_;
  wire g2069_p_spl_;
  wire g2068_n_spl_;
  wire g2069_n_spl_;
  wire g2070_n_spl_;
  wire g2070_n_spl_0;
  wire g2070_p_spl_;
  wire g2070_p_spl_0;
  wire g2072_n_spl_;
  wire g2072_p_spl_;
  wire g2073_n_spl_;
  wire g2073_p_spl_;
  wire g2067_n_spl_;
  wire g2075_p_spl_;
  wire g2067_p_spl_;
  wire g2075_n_spl_;
  wire g2076_n_spl_;
  wire g2076_p_spl_;
  wire g2066_n_spl_;
  wire g2078_p_spl_;
  wire g2066_p_spl_;
  wire g2078_n_spl_;
  wire g2079_n_spl_;
  wire g2079_p_spl_;
  wire g2065_n_spl_;
  wire g2081_p_spl_;
  wire g2065_p_spl_;
  wire g2081_n_spl_;
  wire g2082_n_spl_;
  wire g2082_p_spl_;
  wire G13_p_spl_;
  wire G13_p_spl_0;
  wire G13_p_spl_00;
  wire G13_p_spl_01;
  wire G13_p_spl_1;
  wire G13_n_spl_;
  wire G13_n_spl_0;
  wire G13_n_spl_1;
  wire g2090_p_spl_;
  wire g2091_p_spl_;
  wire g2090_n_spl_;
  wire g2091_n_spl_;
  wire g2092_n_spl_;
  wire g2092_n_spl_0;
  wire g2092_p_spl_;
  wire g2092_p_spl_0;
  wire g2094_n_spl_;
  wire g2094_p_spl_;
  wire g2095_n_spl_;
  wire g2095_p_spl_;
  wire g2089_n_spl_;
  wire g2097_p_spl_;
  wire g2089_p_spl_;
  wire g2097_n_spl_;
  wire g2098_n_spl_;
  wire g2098_p_spl_;
  wire g2088_n_spl_;
  wire g2100_p_spl_;
  wire g2088_p_spl_;
  wire g2100_n_spl_;
  wire g2101_n_spl_;
  wire g2101_p_spl_;
  wire g2087_n_spl_;
  wire g2103_p_spl_;
  wire g2087_p_spl_;
  wire g2103_n_spl_;
  wire g2104_n_spl_;
  wire g2104_p_spl_;
  wire G14_p_spl_;
  wire G14_p_spl_0;
  wire G14_p_spl_00;
  wire G14_p_spl_01;
  wire G14_p_spl_1;
  wire G14_n_spl_;
  wire G14_n_spl_0;
  wire G14_n_spl_1;
  wire g2112_p_spl_;
  wire g2113_p_spl_;
  wire g2112_n_spl_;
  wire g2113_n_spl_;
  wire g2114_n_spl_;
  wire g2114_n_spl_0;
  wire g2114_p_spl_;
  wire g2114_p_spl_0;
  wire g2116_n_spl_;
  wire g2116_p_spl_;
  wire g2117_n_spl_;
  wire g2117_p_spl_;
  wire g2111_n_spl_;
  wire g2119_p_spl_;
  wire g2111_p_spl_;
  wire g2119_n_spl_;
  wire g2120_n_spl_;
  wire g2120_p_spl_;
  wire g2110_n_spl_;
  wire g2122_p_spl_;
  wire g2110_p_spl_;
  wire g2122_n_spl_;
  wire g2123_n_spl_;
  wire g2123_p_spl_;
  wire g2109_n_spl_;
  wire g2125_p_spl_;
  wire g2109_p_spl_;
  wire g2125_n_spl_;
  wire g2126_n_spl_;
  wire g2126_p_spl_;
  wire G15_p_spl_;
  wire G15_p_spl_0;
  wire G15_p_spl_00;
  wire G15_p_spl_1;
  wire G15_n_spl_;
  wire G15_n_spl_0;
  wire G15_n_spl_1;
  wire g2134_p_spl_;
  wire g2135_p_spl_;
  wire g2134_n_spl_;
  wire g2135_n_spl_;
  wire g2136_n_spl_;
  wire g2136_n_spl_0;
  wire g2136_p_spl_;
  wire g2136_p_spl_0;
  wire g2138_n_spl_;
  wire g2138_p_spl_;
  wire g2139_n_spl_;
  wire g2139_p_spl_;
  wire g2133_n_spl_;
  wire g2141_p_spl_;
  wire g2133_p_spl_;
  wire g2141_n_spl_;
  wire g2142_n_spl_;
  wire g2142_p_spl_;
  wire g2132_n_spl_;
  wire g2144_p_spl_;
  wire g2132_p_spl_;
  wire g2144_n_spl_;
  wire g2145_n_spl_;
  wire g2145_p_spl_;
  wire g2131_n_spl_;
  wire g2147_p_spl_;
  wire g2131_p_spl_;
  wire g2147_n_spl_;
  wire g2148_n_spl_;
  wire g2148_p_spl_;
  wire G16_p_spl_;
  wire G16_p_spl_0;
  wire G16_p_spl_00;
  wire G16_p_spl_1;
  wire G16_n_spl_;
  wire G16_n_spl_0;
  wire g2156_p_spl_;
  wire g2157_p_spl_;
  wire g2156_n_spl_;
  wire g2157_n_spl_;
  wire g2158_n_spl_;
  wire g2158_p_spl_;
  wire g2160_n_spl_;
  wire g2160_p_spl_;
  wire g2161_n_spl_;
  wire g2161_p_spl_;
  wire g2155_n_spl_;
  wire g2163_p_spl_;
  wire g2155_p_spl_;
  wire g2163_n_spl_;
  wire g2164_n_spl_;
  wire g2164_p_spl_;
  wire g2154_n_spl_;
  wire g2166_p_spl_;
  wire g2154_p_spl_;
  wire g2166_n_spl_;
  wire g2167_n_spl_;
  wire g2167_p_spl_;
  wire g2153_n_spl_;
  wire g2169_p_spl_;
  wire g2153_p_spl_;
  wire g2169_n_spl_;
  wire g2170_n_spl_;
  wire g2170_p_spl_;
  wire g2177_p_spl_;
  wire g2177_n_spl_;
  wire g2178_p_spl_;
  wire g2179_n_spl_;
  wire g2178_n_spl_;
  wire g2179_p_spl_;
  wire g2180_n_spl_;
  wire g2180_p_spl_;
  wire g2176_n_spl_;
  wire g2182_p_spl_;
  wire g2176_p_spl_;
  wire g2182_n_spl_;
  wire g2183_n_spl_;
  wire g2183_p_spl_;
  wire g2175_n_spl_;
  wire g2185_p_spl_;
  wire g2175_p_spl_;
  wire g2185_n_spl_;
  wire g2186_n_spl_;
  wire g2186_p_spl_;
  wire g2192_n_spl_;
  wire g2193_n_spl_;
  wire g2192_p_spl_;
  wire g2193_p_spl_;
  wire g2194_n_spl_;
  wire g2191_n_spl_;
  wire g2196_p_spl_;
  wire g2191_p_spl_;
  wire g2196_n_spl_;
  wire g2197_n_spl_;
  wire g2201_n_spl_;
  wire g2203_p_spl_;
  wire g2201_p_spl_;
  wire g2203_n_spl_;
  wire g2204_n_spl_;
  wire g2204_p_spl_;
  wire g2205_n_spl_;
  wire g2207_p_spl_;
  wire g2208_n_spl_;
  wire G21_p_spl_;
  wire G21_p_spl_0;
  wire G21_p_spl_00;
  wire G21_p_spl_000;
  wire G21_p_spl_001;
  wire G21_p_spl_01;
  wire G21_p_spl_010;
  wire G21_p_spl_011;
  wire G21_p_spl_1;
  wire G21_p_spl_10;
  wire G21_p_spl_100;
  wire G21_p_spl_101;
  wire G21_p_spl_11;
  wire g1631_p_spl_;
  wire g2228_n_spl_;
  wire g2230_p_spl_;
  wire g1975_n_spl_;
  wire g1997_n_spl_;
  wire g2019_n_spl_;
  wire g2041_n_spl_;
  wire g2063_n_spl_;
  wire g2085_n_spl_;
  wire g2107_n_spl_;
  wire g2129_n_spl_;
  wire g2151_n_spl_;
  wire g2173_n_spl_;
  wire g2189_n_spl_;
  wire g2200_n_spl_;
  wire g2212_n_spl_;

  andX
  g_g389_p
  (
    .dout(g389_p),
    .din1(ffc_0_p),
    .din2(ffc_8_p)
  );


  orX
  g_g390_n
  (
    .dout(g390_n),
    .din1(ffc_31_p),
    .din2(ffc_32_p)
  );


  andX
  g_g391_p
  (
    .dout(g391_p),
    .din1(ffc_33_n),
    .din2(g390_n)
  );


  andX
  g_g392_p
  (
    .dout(g392_p),
    .din1(ffc_34_p),
    .din2(ffc_35_n)
  );


  orX
  g_g393_n
  (
    .dout(g393_n),
    .din1(ffc_36_p),
    .din2(g392_p)
  );


  andX
  g_g394_p
  (
    .dout(g394_p),
    .din1(ffc_37_p),
    .din2(ffc_38_n)
  );


  orX
  g_g395_n
  (
    .dout(g395_n),
    .din1(ffc_39_p),
    .din2(g394_p)
  );


  andX
  g_g396_p
  (
    .dout(g396_p),
    .din1(ffc_40_p),
    .din2(ffc_41_n)
  );


  orX
  g_g397_n
  (
    .dout(g397_n),
    .din1(ffc_42_p),
    .din2(g396_p)
  );


  andX
  g_g398_p
  (
    .dout(g398_p),
    .din1(ffc_43_p),
    .din2(ffc_44_n)
  );


  orX
  g_g399_n
  (
    .dout(g399_n),
    .din1(ffc_45_p),
    .din2(g398_p)
  );


  andX
  g_g400_p
  (
    .dout(g400_p),
    .din1(ffc_46_p),
    .din2(ffc_47_n)
  );


  orX
  g_g401_n
  (
    .dout(g401_n),
    .din1(ffc_48_p),
    .din2(g400_p)
  );


  andX
  g_g402_p
  (
    .dout(g402_p),
    .din1(ffc_49_p),
    .din2(ffc_50_n)
  );


  orX
  g_g403_n
  (
    .dout(g403_n),
    .din1(ffc_51_p),
    .din2(g402_p)
  );


  andX
  g_g404_p
  (
    .dout(g404_p),
    .din1(ffc_52_p),
    .din2(ffc_53_n)
  );


  orX
  g_g405_n
  (
    .dout(g405_n),
    .din1(ffc_54_p),
    .din2(g404_p)
  );


  andX
  g_g406_p
  (
    .dout(g406_p),
    .din1(ffc_55_p),
    .din2(ffc_56_n)
  );


  orX
  g_g407_n
  (
    .dout(g407_n),
    .din1(ffc_57_p),
    .din2(g406_p)
  );


  andX
  g_g408_p
  (
    .dout(g408_p),
    .din1(ffc_58_p),
    .din2(ffc_59_n)
  );


  orX
  g_g409_n
  (
    .dout(g409_n),
    .din1(ffc_60_p),
    .din2(g408_p)
  );


  andX
  g_g410_p
  (
    .dout(g410_p),
    .din1(ffc_61_p),
    .din2(ffc_62_n)
  );


  orX
  g_g411_n
  (
    .dout(g411_n),
    .din1(ffc_63_p),
    .din2(g410_p)
  );


  andX
  g_g412_p
  (
    .dout(g412_p),
    .din1(ffc_81_p),
    .din2(ffc_82_n)
  );


  orX
  g_g413_n
  (
    .dout(g413_n),
    .din1(ffc_85_p),
    .din2(g412_p)
  );


  andX
  g_g414_p
  (
    .dout(g414_p),
    .din1(ffc_90_p),
    .din2(ffc_92_n)
  );


  orX
  g_g415_n
  (
    .dout(g415_n),
    .din1(ffc_95_p),
    .din2(g414_p)
  );


  andX
  g_g416_p
  (
    .dout(g416_p),
    .din1(ffc_99_p),
    .din2(ffc_101_n)
  );


  orX
  g_g417_n
  (
    .dout(g417_n),
    .din1(ffc_104_p),
    .din2(g416_p)
  );


  andX
  g_g418_p
  (
    .dout(g418_p),
    .din1(ffc_108_p),
    .din2(ffc_110_n)
  );


  orX
  g_g419_n
  (
    .dout(g419_n),
    .din1(ffc_113_p),
    .din2(g418_p)
  );


  orX
  g_g420_n
  (
    .dout(g420_n),
    .din1(ffc_115_p),
    .din2(ffc_116_p)
  );


  andX
  g_g421_p
  (
    .dout(g421_p),
    .din1(ffc_136_n),
    .din2(g420_n)
  );


  andX
  g_g422_p
  (
    .dout(g422_p),
    .din1(ffc_136_p),
    .din2(ffc_137_n)
  );


  orX
  g_g423_n
  (
    .dout(g423_n),
    .din1(ffc_143_p),
    .din2(g422_p)
  );


  andX
  g_g424_p
  (
    .dout(g424_p),
    .din1(ffc_149_p),
    .din2(ffc_150_n)
  );


  orX
  g_g425_n
  (
    .dout(g425_n),
    .din1(ffc_155_p),
    .din2(g424_p)
  );


  andX
  g_g426_p
  (
    .dout(g426_p),
    .din1(ffc_161_p),
    .din2(ffc_162_n)
  );


  orX
  g_g427_n
  (
    .dout(g427_n),
    .din1(ffc_169_p),
    .din2(g426_p)
  );


  andX
  g_g428_p
  (
    .dout(g428_p),
    .din1(ffc_175_p),
    .din2(ffc_176_n)
  );


  orX
  g_g429_n
  (
    .dout(g429_n),
    .din1(ffc_204_p),
    .din2(g428_p)
  );


  andX
  g_g430_p
  (
    .dout(g430_p),
    .din1(ffc_215_p),
    .din2(ffc_216_n)
  );


  orX
  g_g431_n
  (
    .dout(g431_n),
    .din1(ffc_244_p_spl_),
    .din2(g430_p)
  );


  andX
  g_g432_p
  (
    .dout(g432_p),
    .din1(ffc_203_p),
    .din2(ffc_244_n)
  );


  orX
  g_g432_n
  (
    .dout(g432_n),
    .din1(ffc_203_n),
    .din2(ffc_244_p_spl_)
  );


  andX
  g_g433_p
  (
    .dout(g433_p),
    .din1(ffc_242_p_spl_),
    .din2(ffc_243_n)
  );


  orX
  g_g433_n
  (
    .dout(g433_n),
    .din1(ffc_242_n_spl_),
    .din2(ffc_243_p)
  );


  andX
  g_g434_p
  (
    .dout(g434_p),
    .din1(g432_n),
    .din2(g433_p)
  );


  orX
  g_g434_n
  (
    .dout(g434_n),
    .din1(g432_p_spl_),
    .din2(g433_n_spl_)
  );


  andX
  g_g435_p
  (
    .dout(g435_p),
    .din1(g432_p_spl_),
    .din2(g433_n_spl_)
  );


  orX
  g_g436_n
  (
    .dout(g436_n),
    .din1(g434_p_spl_),
    .din2(g435_p)
  );


  andX
  g_g437_p
  (
    .dout(g437_p),
    .din1(ffc_242_p_spl_),
    .din2(g434_n)
  );


  orX
  g_g437_n
  (
    .dout(g437_n),
    .din1(ffc_242_n_spl_),
    .din2(g434_p_spl_)
  );


  andX
  g_g438_p
  (
    .dout(g438_p),
    .din1(ffc_168_p),
    .din2(ffc_197_n)
  );


  orX
  g_g438_n
  (
    .dout(g438_n),
    .din1(ffc_168_n),
    .din2(ffc_197_p)
  );


  andX
  g_g439_p
  (
    .dout(g439_p),
    .din1(ffc_232_n_spl_),
    .din2(ffc_233_n)
  );


  orX
  g_g439_n
  (
    .dout(g439_n),
    .din1(ffc_232_p_spl_),
    .din2(ffc_233_p)
  );


  andX
  g_g440_p
  (
    .dout(g440_p),
    .din1(g438_n_spl_),
    .din2(g439_p_spl_)
  );


  orX
  g_g440_n
  (
    .dout(g440_n),
    .din1(g438_p_spl_),
    .din2(g439_n_spl_)
  );


  andX
  g_g441_p
  (
    .dout(g441_p),
    .din1(g438_p_spl_),
    .din2(g439_n_spl_)
  );


  orX
  g_g441_n
  (
    .dout(g441_n),
    .din1(g438_n_spl_),
    .din2(g439_p_spl_)
  );


  andX
  g_g442_p
  (
    .dout(g442_p),
    .din1(g440_n_spl_),
    .din2(g441_n)
  );


  orX
  g_g442_n
  (
    .dout(g442_n),
    .din1(g440_p_spl_),
    .din2(g441_p)
  );


  andX
  g_g443_p
  (
    .dout(g443_p),
    .din1(g437_n),
    .din2(g442_p)
  );


  orX
  g_g443_n
  (
    .dout(g443_n),
    .din1(g437_p_spl_),
    .din2(g442_n_spl_)
  );


  andX
  g_g444_p
  (
    .dout(g444_p),
    .din1(g437_p_spl_),
    .din2(g442_n_spl_)
  );


  orX
  g_g445_n
  (
    .dout(g445_n),
    .din1(g443_p_spl_),
    .din2(g444_p)
  );


  andX
  g_g446_p
  (
    .dout(g446_p),
    .din1(g440_n_spl_),
    .din2(g443_n)
  );


  orX
  g_g446_n
  (
    .dout(g446_n),
    .din1(g440_p_spl_),
    .din2(g443_p_spl_)
  );


  andX
  g_g447_p
  (
    .dout(g447_p),
    .din1(ffc_202_p),
    .din2(ffc_232_n_spl_)
  );


  orX
  g_g447_n
  (
    .dout(g447_n),
    .din1(ffc_202_n),
    .din2(ffc_232_p_spl_)
  );


  andX
  g_g448_p
  (
    .dout(g448_p),
    .din1(ffc_1_p),
    .din2(ffc_30_p_spl_00)
  );


  orX
  g_g448_n
  (
    .dout(g448_n),
    .din1(ffc_1_n),
    .din2(ffc_30_n_spl_00)
  );


  andX
  g_g449_p
  (
    .dout(g449_p),
    .din1(ffc_240_p_spl_),
    .din2(ffc_241_n)
  );


  orX
  g_g449_n
  (
    .dout(g449_n),
    .din1(ffc_240_n_spl_),
    .din2(ffc_241_p)
  );


  andX
  g_g450_p
  (
    .dout(g450_p),
    .din1(g448_n_spl_),
    .din2(g449_p_spl_)
  );


  orX
  g_g450_n
  (
    .dout(g450_n),
    .din1(g448_p_spl_),
    .din2(g449_n_spl_)
  );


  andX
  g_g451_p
  (
    .dout(g451_p),
    .din1(g448_p_spl_),
    .din2(g449_n_spl_)
  );


  orX
  g_g451_n
  (
    .dout(g451_n),
    .din1(g448_n_spl_),
    .din2(g449_p_spl_)
  );


  andX
  g_g452_p
  (
    .dout(g452_p),
    .din1(g450_n_spl_),
    .din2(g451_n)
  );


  orX
  g_g452_n
  (
    .dout(g452_n),
    .din1(g450_p_spl_),
    .din2(g451_p)
  );


  andX
  g_g453_p
  (
    .dout(g453_p),
    .din1(g447_n_spl_),
    .din2(g452_p_spl_)
  );


  orX
  g_g453_n
  (
    .dout(g453_n),
    .din1(g447_p_spl_),
    .din2(g452_n_spl_)
  );


  andX
  g_g454_p
  (
    .dout(g454_p),
    .din1(g447_p_spl_),
    .din2(g452_n_spl_)
  );


  orX
  g_g454_n
  (
    .dout(g454_n),
    .din1(g447_n_spl_),
    .din2(g452_p_spl_)
  );


  andX
  g_g455_p
  (
    .dout(g455_p),
    .din1(g453_n_spl_),
    .din2(g454_n)
  );


  orX
  g_g455_n
  (
    .dout(g455_n),
    .din1(g453_p_spl_),
    .din2(g454_p)
  );


  andX
  g_g456_p
  (
    .dout(g456_p),
    .din1(g446_n),
    .din2(g455_p)
  );


  orX
  g_g456_n
  (
    .dout(g456_n),
    .din1(g446_p_spl_),
    .din2(g455_n_spl_)
  );


  andX
  g_g457_p
  (
    .dout(g457_p),
    .din1(g446_p_spl_),
    .din2(g455_n_spl_)
  );


  orX
  g_g458_n
  (
    .dout(g458_n),
    .din1(g456_p_spl_),
    .din2(g457_p)
  );


  andX
  g_g459_p
  (
    .dout(g459_p),
    .din1(g453_n_spl_),
    .din2(g456_n)
  );


  orX
  g_g459_n
  (
    .dout(g459_n),
    .din1(g453_p_spl_),
    .din2(g456_p_spl_)
  );


  andX
  g_g460_p
  (
    .dout(g460_p),
    .din1(ffc_240_p_spl_),
    .din2(g450_n_spl_)
  );


  orX
  g_g460_n
  (
    .dout(g460_n),
    .din1(ffc_240_n_spl_),
    .din2(g450_p_spl_)
  );


  andX
  g_g461_p
  (
    .dout(g461_p),
    .din1(ffc_2_p),
    .din2(ffc_30_p_spl_00)
  );


  orX
  g_g461_n
  (
    .dout(g461_n),
    .din1(ffc_2_n),
    .din2(ffc_30_n_spl_00)
  );


  andX
  g_g462_p
  (
    .dout(g462_p),
    .din1(ffc_167_p),
    .din2(ffc_198_n)
  );


  orX
  g_g462_n
  (
    .dout(g462_n),
    .din1(ffc_167_n),
    .din2(ffc_198_p)
  );


  andX
  g_g463_p
  (
    .dout(g463_p),
    .din1(ffc_234_n_spl_),
    .din2(ffc_235_n)
  );


  orX
  g_g463_n
  (
    .dout(g463_n),
    .din1(ffc_234_p_spl_),
    .din2(ffc_235_p)
  );


  andX
  g_g464_p
  (
    .dout(g464_p),
    .din1(g462_n_spl_),
    .din2(g463_p_spl_)
  );


  orX
  g_g464_n
  (
    .dout(g464_n),
    .din1(g462_p_spl_),
    .din2(g463_n_spl_)
  );


  andX
  g_g465_p
  (
    .dout(g465_p),
    .din1(g462_p_spl_),
    .din2(g463_n_spl_)
  );


  orX
  g_g465_n
  (
    .dout(g465_n),
    .din1(g462_n_spl_),
    .din2(g463_p_spl_)
  );


  andX
  g_g466_p
  (
    .dout(g466_p),
    .din1(g464_n_spl_),
    .din2(g465_n)
  );


  orX
  g_g466_n
  (
    .dout(g466_n),
    .din1(g464_p_spl_),
    .din2(g465_p)
  );


  andX
  g_g467_p
  (
    .dout(g467_p),
    .din1(g461_n_spl_),
    .din2(g466_p_spl_)
  );


  orX
  g_g467_n
  (
    .dout(g467_n),
    .din1(g461_p_spl_),
    .din2(g466_n_spl_)
  );


  andX
  g_g468_p
  (
    .dout(g468_p),
    .din1(g461_p_spl_),
    .din2(g466_n_spl_)
  );


  orX
  g_g468_n
  (
    .dout(g468_n),
    .din1(g461_n_spl_),
    .din2(g466_p_spl_)
  );


  andX
  g_g469_p
  (
    .dout(g469_p),
    .din1(g467_n_spl_),
    .din2(g468_n)
  );


  orX
  g_g469_n
  (
    .dout(g469_n),
    .din1(g467_p_spl_),
    .din2(g468_p)
  );


  andX
  g_g470_p
  (
    .dout(g470_p),
    .din1(g460_n_spl_),
    .din2(g469_p_spl_)
  );


  orX
  g_g470_n
  (
    .dout(g470_n),
    .din1(g460_p_spl_),
    .din2(g469_n_spl_)
  );


  andX
  g_g471_p
  (
    .dout(g471_p),
    .din1(g460_p_spl_),
    .din2(g469_n_spl_)
  );


  orX
  g_g471_n
  (
    .dout(g471_n),
    .din1(g460_n_spl_),
    .din2(g469_p_spl_)
  );


  andX
  g_g472_p
  (
    .dout(g472_p),
    .din1(g470_n_spl_),
    .din2(g471_n)
  );


  orX
  g_g472_n
  (
    .dout(g472_n),
    .din1(g470_p_spl_),
    .din2(g471_p)
  );


  andX
  g_g473_p
  (
    .dout(g473_p),
    .din1(g459_n),
    .din2(g472_p)
  );


  orX
  g_g473_n
  (
    .dout(g473_n),
    .din1(g459_p_spl_),
    .din2(g472_n_spl_)
  );


  andX
  g_g474_p
  (
    .dout(g474_p),
    .din1(g459_p_spl_),
    .din2(g472_n_spl_)
  );


  orX
  g_g475_n
  (
    .dout(g475_n),
    .din1(g473_p_spl_),
    .din2(g474_p)
  );


  andX
  g_g476_p
  (
    .dout(g476_p),
    .din1(g470_n_spl_),
    .din2(g473_n)
  );


  orX
  g_g476_n
  (
    .dout(g476_n),
    .din1(g470_p_spl_),
    .din2(g473_p_spl_)
  );


  andX
  g_g477_p
  (
    .dout(g477_p),
    .din1(g464_n_spl_),
    .din2(g467_n_spl_)
  );


  orX
  g_g477_n
  (
    .dout(g477_n),
    .din1(g464_p_spl_),
    .din2(g467_p_spl_)
  );


  andX
  g_g478_p
  (
    .dout(g478_p),
    .din1(ffc_3_p),
    .din2(ffc_30_p_spl_01)
  );


  orX
  g_g478_n
  (
    .dout(g478_n),
    .din1(ffc_3_n),
    .din2(ffc_30_n_spl_01)
  );


  andX
  g_g479_p
  (
    .dout(g479_p),
    .din1(ffc_201_p),
    .din2(ffc_234_n_spl_)
  );


  orX
  g_g479_n
  (
    .dout(g479_n),
    .din1(ffc_201_n),
    .din2(ffc_234_p_spl_)
  );


  andX
  g_g480_p
  (
    .dout(g480_p),
    .din1(ffc_4_p_spl_),
    .din2(ffc_26_p_spl_0)
  );


  orX
  g_g480_n
  (
    .dout(g480_n),
    .din1(ffc_4_n_spl_),
    .din2(ffc_26_n_spl_0)
  );


  andX
  g_g481_p
  (
    .dout(g481_p),
    .din1(ffc_238_p_spl_),
    .din2(ffc_239_n)
  );


  orX
  g_g481_n
  (
    .dout(g481_n),
    .din1(ffc_238_n_spl_),
    .din2(ffc_239_p)
  );


  andX
  g_g482_p
  (
    .dout(g482_p),
    .din1(g480_n_spl_),
    .din2(g481_p_spl_)
  );


  orX
  g_g482_n
  (
    .dout(g482_n),
    .din1(g480_p_spl_),
    .din2(g481_n_spl_)
  );


  andX
  g_g483_p
  (
    .dout(g483_p),
    .din1(g480_p_spl_),
    .din2(g481_n_spl_)
  );


  orX
  g_g483_n
  (
    .dout(g483_n),
    .din1(g480_n_spl_),
    .din2(g481_p_spl_)
  );


  andX
  g_g484_p
  (
    .dout(g484_p),
    .din1(g482_n_spl_),
    .din2(g483_n)
  );


  orX
  g_g484_n
  (
    .dout(g484_n),
    .din1(g482_p_spl_),
    .din2(g483_p)
  );


  andX
  g_g485_p
  (
    .dout(g485_p),
    .din1(g479_n_spl_),
    .din2(g484_p_spl_)
  );


  orX
  g_g485_n
  (
    .dout(g485_n),
    .din1(g479_p_spl_),
    .din2(g484_n_spl_)
  );


  andX
  g_g486_p
  (
    .dout(g486_p),
    .din1(g479_p_spl_),
    .din2(g484_n_spl_)
  );


  orX
  g_g486_n
  (
    .dout(g486_n),
    .din1(g479_n_spl_),
    .din2(g484_p_spl_)
  );


  andX
  g_g487_p
  (
    .dout(g487_p),
    .din1(g485_n_spl_),
    .din2(g486_n)
  );


  orX
  g_g487_n
  (
    .dout(g487_n),
    .din1(g485_p_spl_),
    .din2(g486_p)
  );


  andX
  g_g488_p
  (
    .dout(g488_p),
    .din1(g478_n_spl_),
    .din2(g487_p_spl_)
  );


  orX
  g_g488_n
  (
    .dout(g488_n),
    .din1(g478_p_spl_),
    .din2(g487_n_spl_)
  );


  andX
  g_g489_p
  (
    .dout(g489_p),
    .din1(g478_p_spl_),
    .din2(g487_n_spl_)
  );


  orX
  g_g489_n
  (
    .dout(g489_n),
    .din1(g478_n_spl_),
    .din2(g487_p_spl_)
  );


  andX
  g_g490_p
  (
    .dout(g490_p),
    .din1(g488_n_spl_),
    .din2(g489_n)
  );


  orX
  g_g490_n
  (
    .dout(g490_n),
    .din1(g488_p_spl_),
    .din2(g489_p)
  );


  andX
  g_g491_p
  (
    .dout(g491_p),
    .din1(g477_n_spl_),
    .din2(g490_p_spl_)
  );


  orX
  g_g491_n
  (
    .dout(g491_n),
    .din1(g477_p_spl_),
    .din2(g490_n_spl_)
  );


  andX
  g_g492_p
  (
    .dout(g492_p),
    .din1(g477_p_spl_),
    .din2(g490_n_spl_)
  );


  orX
  g_g492_n
  (
    .dout(g492_n),
    .din1(g477_n_spl_),
    .din2(g490_p_spl_)
  );


  andX
  g_g493_p
  (
    .dout(g493_p),
    .din1(g491_n_spl_),
    .din2(g492_n)
  );


  orX
  g_g493_n
  (
    .dout(g493_n),
    .din1(g491_p_spl_),
    .din2(g492_p)
  );


  andX
  g_g494_p
  (
    .dout(g494_p),
    .din1(g476_n),
    .din2(g493_p)
  );


  orX
  g_g494_n
  (
    .dout(g494_n),
    .din1(g476_p_spl_),
    .din2(g493_n_spl_)
  );


  andX
  g_g495_p
  (
    .dout(g495_p),
    .din1(g476_p_spl_),
    .din2(g493_n_spl_)
  );


  orX
  g_g496_n
  (
    .dout(g496_n),
    .din1(g494_p_spl_),
    .din2(g495_p)
  );


  andX
  g_g497_p
  (
    .dout(g497_p),
    .din1(g491_n_spl_),
    .din2(g494_n)
  );


  orX
  g_g497_n
  (
    .dout(g497_n),
    .din1(g491_p_spl_),
    .din2(g494_p_spl_)
  );


  andX
  g_g498_p
  (
    .dout(g498_p),
    .din1(g485_n_spl_),
    .din2(g488_n_spl_)
  );


  orX
  g_g498_n
  (
    .dout(g498_n),
    .din1(g485_p_spl_),
    .din2(g488_p_spl_)
  );


  andX
  g_g499_p
  (
    .dout(g499_p),
    .din1(ffc_4_p_spl_),
    .din2(ffc_30_p_spl_01)
  );


  orX
  g_g499_n
  (
    .dout(g499_n),
    .din1(ffc_4_n_spl_),
    .din2(ffc_30_n_spl_01)
  );


  andX
  g_g500_p
  (
    .dout(g500_p),
    .din1(ffc_238_p_spl_),
    .din2(g482_n_spl_)
  );


  orX
  g_g500_n
  (
    .dout(g500_n),
    .din1(ffc_238_n_spl_),
    .din2(g482_p_spl_)
  );


  andX
  g_g501_p
  (
    .dout(g501_p),
    .din1(ffc_5_p_spl_),
    .din2(ffc_26_p_spl_0)
  );


  orX
  g_g501_n
  (
    .dout(g501_n),
    .din1(ffc_5_n_spl_),
    .din2(ffc_26_n_spl_0)
  );


  andX
  g_g502_p
  (
    .dout(g502_p),
    .din1(ffc_166_p),
    .din2(ffc_199_n)
  );


  orX
  g_g502_n
  (
    .dout(g502_n),
    .din1(ffc_166_n),
    .din2(ffc_199_p)
  );


  andX
  g_g503_p
  (
    .dout(g503_p),
    .din1(ffc_236_n_spl_),
    .din2(ffc_237_n)
  );


  orX
  g_g503_n
  (
    .dout(g503_n),
    .din1(ffc_236_p_spl_),
    .din2(ffc_237_p)
  );


  andX
  g_g504_p
  (
    .dout(g504_p),
    .din1(g502_n_spl_),
    .din2(g503_p_spl_)
  );


  orX
  g_g504_n
  (
    .dout(g504_n),
    .din1(g502_p_spl_),
    .din2(g503_n_spl_)
  );


  andX
  g_g505_p
  (
    .dout(g505_p),
    .din1(g502_p_spl_),
    .din2(g503_n_spl_)
  );


  orX
  g_g505_n
  (
    .dout(g505_n),
    .din1(g502_n_spl_),
    .din2(g503_p_spl_)
  );


  andX
  g_g506_p
  (
    .dout(g506_p),
    .din1(g504_n_spl_),
    .din2(g505_n)
  );


  orX
  g_g506_n
  (
    .dout(g506_n),
    .din1(g504_p_spl_),
    .din2(g505_p)
  );


  andX
  g_g507_p
  (
    .dout(g507_p),
    .din1(g501_n_spl_),
    .din2(g506_p_spl_)
  );


  orX
  g_g507_n
  (
    .dout(g507_n),
    .din1(g501_p_spl_),
    .din2(g506_n_spl_)
  );


  andX
  g_g508_p
  (
    .dout(g508_p),
    .din1(g501_p_spl_),
    .din2(g506_n_spl_)
  );


  orX
  g_g508_n
  (
    .dout(g508_n),
    .din1(g501_n_spl_),
    .din2(g506_p_spl_)
  );


  andX
  g_g509_p
  (
    .dout(g509_p),
    .din1(g507_n_spl_),
    .din2(g508_n)
  );


  orX
  g_g509_n
  (
    .dout(g509_n),
    .din1(g507_p_spl_),
    .din2(g508_p)
  );


  andX
  g_g510_p
  (
    .dout(g510_p),
    .din1(g500_n_spl_),
    .din2(g509_p_spl_)
  );


  orX
  g_g510_n
  (
    .dout(g510_n),
    .din1(g500_p_spl_),
    .din2(g509_n_spl_)
  );


  andX
  g_g511_p
  (
    .dout(g511_p),
    .din1(g500_p_spl_),
    .din2(g509_n_spl_)
  );


  orX
  g_g511_n
  (
    .dout(g511_n),
    .din1(g500_n_spl_),
    .din2(g509_p_spl_)
  );


  andX
  g_g512_p
  (
    .dout(g512_p),
    .din1(g510_n_spl_),
    .din2(g511_n)
  );


  orX
  g_g512_n
  (
    .dout(g512_n),
    .din1(g510_p_spl_),
    .din2(g511_p)
  );


  andX
  g_g513_p
  (
    .dout(g513_p),
    .din1(g499_n_spl_),
    .din2(g512_p_spl_)
  );


  orX
  g_g513_n
  (
    .dout(g513_n),
    .din1(g499_p_spl_),
    .din2(g512_n_spl_)
  );


  andX
  g_g514_p
  (
    .dout(g514_p),
    .din1(g499_p_spl_),
    .din2(g512_n_spl_)
  );


  orX
  g_g514_n
  (
    .dout(g514_n),
    .din1(g499_n_spl_),
    .din2(g512_p_spl_)
  );


  andX
  g_g515_p
  (
    .dout(g515_p),
    .din1(g513_n_spl_),
    .din2(g514_n)
  );


  orX
  g_g515_n
  (
    .dout(g515_n),
    .din1(g513_p_spl_),
    .din2(g514_p)
  );


  andX
  g_g516_p
  (
    .dout(g516_p),
    .din1(g498_n_spl_),
    .din2(g515_p_spl_)
  );


  orX
  g_g516_n
  (
    .dout(g516_n),
    .din1(g498_p_spl_),
    .din2(g515_n_spl_)
  );


  andX
  g_g517_p
  (
    .dout(g517_p),
    .din1(g498_p_spl_),
    .din2(g515_n_spl_)
  );


  orX
  g_g517_n
  (
    .dout(g517_n),
    .din1(g498_n_spl_),
    .din2(g515_p_spl_)
  );


  andX
  g_g518_p
  (
    .dout(g518_p),
    .din1(g516_n_spl_),
    .din2(g517_n)
  );


  orX
  g_g518_n
  (
    .dout(g518_n),
    .din1(g516_p_spl_),
    .din2(g517_p)
  );


  andX
  g_g519_p
  (
    .dout(g519_p),
    .din1(g497_n),
    .din2(g518_p)
  );


  orX
  g_g519_n
  (
    .dout(g519_n),
    .din1(g497_p_spl_),
    .din2(g518_n_spl_)
  );


  andX
  g_g520_p
  (
    .dout(g520_p),
    .din1(g497_p_spl_),
    .din2(g518_n_spl_)
  );


  orX
  g_g521_n
  (
    .dout(g521_n),
    .din1(g519_p_spl_),
    .din2(g520_p)
  );


  andX
  g_g522_p
  (
    .dout(g522_p),
    .din1(g516_n_spl_),
    .din2(g519_n)
  );


  orX
  g_g522_n
  (
    .dout(g522_n),
    .din1(g516_p_spl_),
    .din2(g519_p_spl_)
  );


  andX
  g_g523_p
  (
    .dout(g523_p),
    .din1(g510_n_spl_),
    .din2(g513_n_spl_)
  );


  orX
  g_g523_n
  (
    .dout(g523_n),
    .din1(g510_p_spl_),
    .din2(g513_p_spl_)
  );


  andX
  g_g524_p
  (
    .dout(g524_p),
    .din1(ffc_5_p_spl_),
    .din2(ffc_30_p_spl_10)
  );


  orX
  g_g524_n
  (
    .dout(g524_n),
    .din1(ffc_5_n_spl_),
    .din2(ffc_30_n_spl_10)
  );


  andX
  g_g525_p
  (
    .dout(g525_p),
    .din1(g504_n_spl_),
    .din2(g507_n_spl_)
  );


  orX
  g_g525_n
  (
    .dout(g525_n),
    .din1(g504_p_spl_),
    .din2(g507_p_spl_)
  );


  andX
  g_g526_p
  (
    .dout(g526_p),
    .din1(ffc_6_p_spl_),
    .din2(ffc_26_p_spl_1)
  );


  orX
  g_g526_n
  (
    .dout(g526_n),
    .din1(ffc_6_n_spl_),
    .din2(ffc_26_n_spl_1)
  );


  andX
  g_g527_p
  (
    .dout(g527_p),
    .din1(ffc_7_p_spl_0),
    .din2(ffc_22_p)
  );


  orX
  g_g527_n
  (
    .dout(g527_n),
    .din1(ffc_7_n_spl_0),
    .din2(ffc_22_n)
  );


  andX
  g_g528_p
  (
    .dout(g528_p),
    .din1(ffc_200_p),
    .din2(ffc_236_n_spl_)
  );


  orX
  g_g528_n
  (
    .dout(g528_n),
    .din1(ffc_200_n),
    .din2(ffc_236_p_spl_)
  );


  andX
  g_g529_p
  (
    .dout(g529_p),
    .din1(g527_n_spl_),
    .din2(g528_n_spl_)
  );


  orX
  g_g529_n
  (
    .dout(g529_n),
    .din1(g527_p_spl_),
    .din2(g528_p_spl_)
  );


  andX
  g_g530_p
  (
    .dout(g530_p),
    .din1(g527_p_spl_),
    .din2(g528_p_spl_)
  );


  orX
  g_g530_n
  (
    .dout(g530_n),
    .din1(g527_n_spl_),
    .din2(g528_n_spl_)
  );


  andX
  g_g531_p
  (
    .dout(g531_p),
    .din1(g529_n_spl_),
    .din2(g530_n)
  );


  orX
  g_g531_n
  (
    .dout(g531_n),
    .din1(g529_p_spl_),
    .din2(g530_p)
  );


  andX
  g_g532_p
  (
    .dout(g532_p),
    .din1(g526_n_spl_),
    .din2(g531_p_spl_)
  );


  orX
  g_g532_n
  (
    .dout(g532_n),
    .din1(g526_p_spl_),
    .din2(g531_n_spl_)
  );


  andX
  g_g533_p
  (
    .dout(g533_p),
    .din1(g526_p_spl_),
    .din2(g531_n_spl_)
  );


  orX
  g_g533_n
  (
    .dout(g533_n),
    .din1(g526_n_spl_),
    .din2(g531_p_spl_)
  );


  andX
  g_g534_p
  (
    .dout(g534_p),
    .din1(g532_n_spl_),
    .din2(g533_n)
  );


  orX
  g_g534_n
  (
    .dout(g534_n),
    .din1(g532_p_spl_),
    .din2(g533_p)
  );


  andX
  g_g535_p
  (
    .dout(g535_p),
    .din1(g525_n_spl_),
    .din2(g534_p_spl_)
  );


  orX
  g_g535_n
  (
    .dout(g535_n),
    .din1(g525_p_spl_),
    .din2(g534_n_spl_)
  );


  andX
  g_g536_p
  (
    .dout(g536_p),
    .din1(g525_p_spl_),
    .din2(g534_n_spl_)
  );


  orX
  g_g536_n
  (
    .dout(g536_n),
    .din1(g525_n_spl_),
    .din2(g534_p_spl_)
  );


  andX
  g_g537_p
  (
    .dout(g537_p),
    .din1(g535_n_spl_),
    .din2(g536_n)
  );


  orX
  g_g537_n
  (
    .dout(g537_n),
    .din1(g535_p_spl_),
    .din2(g536_p)
  );


  andX
  g_g538_p
  (
    .dout(g538_p),
    .din1(g524_n_spl_),
    .din2(g537_p_spl_)
  );


  orX
  g_g538_n
  (
    .dout(g538_n),
    .din1(g524_p_spl_),
    .din2(g537_n_spl_)
  );


  andX
  g_g539_p
  (
    .dout(g539_p),
    .din1(g524_p_spl_),
    .din2(g537_n_spl_)
  );


  orX
  g_g539_n
  (
    .dout(g539_n),
    .din1(g524_n_spl_),
    .din2(g537_p_spl_)
  );


  andX
  g_g540_p
  (
    .dout(g540_p),
    .din1(g538_n_spl_),
    .din2(g539_n)
  );


  orX
  g_g540_n
  (
    .dout(g540_n),
    .din1(g538_p_spl_),
    .din2(g539_p)
  );


  andX
  g_g541_p
  (
    .dout(g541_p),
    .din1(g523_n_spl_),
    .din2(g540_p_spl_)
  );


  orX
  g_g541_n
  (
    .dout(g541_n),
    .din1(g523_p_spl_),
    .din2(g540_n_spl_)
  );


  andX
  g_g542_p
  (
    .dout(g542_p),
    .din1(g523_p_spl_),
    .din2(g540_n_spl_)
  );


  orX
  g_g542_n
  (
    .dout(g542_n),
    .din1(g523_n_spl_),
    .din2(g540_p_spl_)
  );


  andX
  g_g543_p
  (
    .dout(g543_p),
    .din1(g541_n_spl_),
    .din2(g542_n)
  );


  orX
  g_g543_n
  (
    .dout(g543_n),
    .din1(g541_p_spl_),
    .din2(g542_p)
  );


  andX
  g_g544_p
  (
    .dout(g544_p),
    .din1(g522_n),
    .din2(g543_p)
  );


  orX
  g_g544_n
  (
    .dout(g544_n),
    .din1(g522_p_spl_),
    .din2(g543_n_spl_)
  );


  andX
  g_g545_p
  (
    .dout(g545_p),
    .din1(g522_p_spl_),
    .din2(g543_n_spl_)
  );


  orX
  g_g546_n
  (
    .dout(g546_n),
    .din1(g544_p_spl_),
    .din2(g545_p)
  );


  andX
  g_g547_p
  (
    .dout(g547_p),
    .din1(g541_n_spl_),
    .din2(g544_n)
  );


  orX
  g_g547_n
  (
    .dout(g547_n),
    .din1(g541_p_spl_),
    .din2(g544_p_spl_)
  );


  andX
  g_g548_p
  (
    .dout(g548_p),
    .din1(g535_n_spl_),
    .din2(g538_n_spl_)
  );


  orX
  g_g548_n
  (
    .dout(g548_n),
    .din1(g535_p_spl_),
    .din2(g538_p_spl_)
  );


  andX
  g_g549_p
  (
    .dout(g549_p),
    .din1(ffc_6_p_spl_),
    .din2(ffc_30_p_spl_10)
  );


  orX
  g_g549_n
  (
    .dout(g549_n),
    .din1(ffc_6_n_spl_),
    .din2(ffc_30_n_spl_10)
  );


  andX
  g_g550_p
  (
    .dout(g550_p),
    .din1(ffc_7_p_spl_0),
    .din2(ffc_26_p_spl_1)
  );


  orX
  g_g550_n
  (
    .dout(g550_n),
    .din1(ffc_7_n_spl_0),
    .din2(ffc_26_n_spl_1)
  );


  andX
  g_g551_p
  (
    .dout(g551_p),
    .din1(g529_n_spl_),
    .din2(g532_n_spl_)
  );


  orX
  g_g551_n
  (
    .dout(g551_n),
    .din1(g529_p_spl_),
    .din2(g532_p_spl_)
  );


  andX
  g_g552_p
  (
    .dout(g552_p),
    .din1(g550_n_spl_),
    .din2(g551_n_spl_)
  );


  orX
  g_g552_n
  (
    .dout(g552_n),
    .din1(g550_p_spl_),
    .din2(g551_p_spl_)
  );


  andX
  g_g553_p
  (
    .dout(g553_p),
    .din1(g550_p_spl_),
    .din2(g551_p_spl_)
  );


  orX
  g_g553_n
  (
    .dout(g553_n),
    .din1(g550_n_spl_),
    .din2(g551_n_spl_)
  );


  andX
  g_g554_p
  (
    .dout(g554_p),
    .din1(g552_n_spl_),
    .din2(g553_n)
  );


  orX
  g_g554_n
  (
    .dout(g554_n),
    .din1(g552_p_spl_),
    .din2(g553_p)
  );


  andX
  g_g555_p
  (
    .dout(g555_p),
    .din1(g549_n_spl_),
    .din2(g554_p_spl_)
  );


  orX
  g_g555_n
  (
    .dout(g555_n),
    .din1(g549_p_spl_),
    .din2(g554_n_spl_)
  );


  andX
  g_g556_p
  (
    .dout(g556_p),
    .din1(g549_p_spl_),
    .din2(g554_n_spl_)
  );


  orX
  g_g556_n
  (
    .dout(g556_n),
    .din1(g549_n_spl_),
    .din2(g554_p_spl_)
  );


  andX
  g_g557_p
  (
    .dout(g557_p),
    .din1(g555_n_spl_),
    .din2(g556_n)
  );


  orX
  g_g557_n
  (
    .dout(g557_n),
    .din1(g555_p_spl_),
    .din2(g556_p)
  );


  andX
  g_g558_p
  (
    .dout(g558_p),
    .din1(g548_n_spl_),
    .din2(g557_p_spl_)
  );


  orX
  g_g558_n
  (
    .dout(g558_n),
    .din1(g548_p_spl_),
    .din2(g557_n_spl_)
  );


  andX
  g_g559_p
  (
    .dout(g559_p),
    .din1(g548_p_spl_),
    .din2(g557_n_spl_)
  );


  orX
  g_g559_n
  (
    .dout(g559_n),
    .din1(g548_n_spl_),
    .din2(g557_p_spl_)
  );


  andX
  g_g560_p
  (
    .dout(g560_p),
    .din1(g558_n_spl_),
    .din2(g559_n)
  );


  orX
  g_g560_n
  (
    .dout(g560_n),
    .din1(g558_p_spl_),
    .din2(g559_p)
  );


  andX
  g_g561_p
  (
    .dout(g561_p),
    .din1(g547_n),
    .din2(g560_p)
  );


  orX
  g_g561_n
  (
    .dout(g561_n),
    .din1(g547_p_spl_),
    .din2(g560_n_spl_)
  );


  andX
  g_g562_p
  (
    .dout(g562_p),
    .din1(g547_p_spl_),
    .din2(g560_n_spl_)
  );


  orX
  g_g563_n
  (
    .dout(g563_n),
    .din1(g561_p_spl_),
    .din2(g562_p)
  );


  andX
  g_g564_p
  (
    .dout(g564_p),
    .din1(ffc_7_p_spl_),
    .din2(ffc_30_p_spl_1)
  );


  orX
  g_g564_n
  (
    .dout(g564_n),
    .din1(ffc_7_n_spl_),
    .din2(ffc_30_n_spl_1)
  );


  andX
  g_g565_p
  (
    .dout(g565_p),
    .din1(g552_n_spl_),
    .din2(g555_n_spl_)
  );


  orX
  g_g565_n
  (
    .dout(g565_n),
    .din1(g552_p_spl_),
    .din2(g555_p_spl_)
  );


  andX
  g_g566_p
  (
    .dout(g566_p),
    .din1(g564_n_spl_),
    .din2(g565_n_spl_)
  );


  orX
  g_g566_n
  (
    .dout(g566_n),
    .din1(g564_p_spl_),
    .din2(g565_p_spl_)
  );


  andX
  g_g567_p
  (
    .dout(g567_p),
    .din1(g558_n_spl_),
    .din2(g561_n)
  );


  orX
  g_g567_n
  (
    .dout(g567_n),
    .din1(g558_p_spl_),
    .din2(g561_p_spl_)
  );


  andX
  g_g568_p
  (
    .dout(g568_p),
    .din1(g564_p_spl_),
    .din2(g565_p_spl_)
  );


  orX
  g_g568_n
  (
    .dout(g568_n),
    .din1(g564_n_spl_),
    .din2(g565_n_spl_)
  );


  andX
  g_g569_p
  (
    .dout(g569_p),
    .din1(g566_n_spl_),
    .din2(g568_n)
  );


  orX
  g_g569_n
  (
    .dout(g569_n),
    .din1(g566_p),
    .din2(g568_p)
  );


  orX
  g_g570_n
  (
    .dout(g570_n),
    .din1(g567_p),
    .din2(g569_n)
  );


  andX
  g_g571_p
  (
    .dout(g571_p),
    .din1(g566_n_spl_),
    .din2(g570_n_spl_)
  );


  orX
  g_g572_n
  (
    .dout(g572_n),
    .din1(g567_n),
    .din2(g569_p)
  );


  andX
  g_g573_p
  (
    .dout(g573_p),
    .din1(g570_n_spl_),
    .din2(g572_n)
  );


  andX
  g_g574_p
  (
    .dout(g574_p),
    .din1(ffc_25_p_spl_000),
    .din2(ffc_80_p_spl_)
  );


  orX
  g_g574_n
  (
    .dout(g574_n),
    .din1(ffc_25_n_spl_000),
    .din2(ffc_80_n_spl_)
  );


  andX
  g_g575_p
  (
    .dout(g575_p),
    .din1(ffc_225_p),
    .din2(ffc_272_n)
  );


  orX
  g_g575_n
  (
    .dout(g575_n),
    .din1(ffc_225_n),
    .din2(ffc_272_p_spl_)
  );


  andX
  g_g576_p
  (
    .dout(g576_p),
    .din1(ffc_250_n),
    .din2(ffc_271_n)
  );


  orX
  g_g576_n
  (
    .dout(g576_n),
    .din1(ffc_250_p),
    .din2(ffc_271_p)
  );


  andX
  g_g577_p
  (
    .dout(g577_p),
    .din1(g575_n_spl_),
    .din2(g576_p_spl_)
  );


  orX
  g_g577_n
  (
    .dout(g577_n),
    .din1(g575_p_spl_),
    .din2(g576_n_spl_)
  );


  andX
  g_g578_p
  (
    .dout(g578_p),
    .din1(g575_p_spl_),
    .din2(g576_n_spl_)
  );


  orX
  g_g578_n
  (
    .dout(g578_n),
    .din1(g575_n_spl_),
    .din2(g576_p_spl_)
  );


  andX
  g_g579_p
  (
    .dout(g579_p),
    .din1(g577_n_spl_),
    .din2(g578_n)
  );


  orX
  g_g579_n
  (
    .dout(g579_n),
    .din1(g577_p_spl_),
    .din2(g578_p)
  );


  andX
  g_g580_p
  (
    .dout(g580_p),
    .din1(g574_n),
    .din2(g579_p_spl_)
  );


  orX
  g_g580_n
  (
    .dout(g580_n),
    .din1(g574_p_spl_),
    .din2(g579_n)
  );


  orX
  g_g581_n
  (
    .dout(g581_n),
    .din1(ffc_29_n_spl_000),
    .din2(ffc_80_n_spl_)
  );


  andX
  g_g582_p
  (
    .dout(g582_p),
    .din1(g577_n_spl_),
    .din2(g580_n)
  );


  orX
  g_g582_n
  (
    .dout(g582_n),
    .din1(g577_p_spl_),
    .din2(g580_p_spl_)
  );


  andX
  g_g583_p
  (
    .dout(g583_p),
    .din1(ffc_25_p_spl_000),
    .din2(ffc_79_p_spl_)
  );


  orX
  g_g583_n
  (
    .dout(g583_n),
    .din1(ffc_25_n_spl_000),
    .din2(ffc_79_n_spl_)
  );


  andX
  g_g584_p
  (
    .dout(g584_p),
    .din1(ffc_270_n_spl_),
    .din2(ffc_275_n_spl_)
  );


  orX
  g_g584_n
  (
    .dout(g584_n),
    .din1(ffc_270_p_spl_),
    .din2(ffc_275_p_spl_)
  );


  andX
  g_g585_p
  (
    .dout(g585_p),
    .din1(ffc_270_p_spl_),
    .din2(ffc_275_p_spl_)
  );


  orX
  g_g585_n
  (
    .dout(g585_n),
    .din1(ffc_270_n_spl_),
    .din2(ffc_275_n_spl_)
  );


  andX
  g_g586_p
  (
    .dout(g586_p),
    .din1(g584_n_spl_),
    .din2(g585_n)
  );


  orX
  g_g586_n
  (
    .dout(g586_n),
    .din1(g584_p_spl_),
    .din2(g585_p)
  );


  andX
  g_g587_p
  (
    .dout(g587_p),
    .din1(g583_n_spl_),
    .din2(g586_p_spl_)
  );


  orX
  g_g587_n
  (
    .dout(g587_n),
    .din1(g583_p_spl_),
    .din2(g586_n_spl_)
  );


  andX
  g_g588_p
  (
    .dout(g588_p),
    .din1(g583_p_spl_),
    .din2(g586_n_spl_)
  );


  orX
  g_g588_n
  (
    .dout(g588_n),
    .din1(g583_n_spl_),
    .din2(g586_p_spl_)
  );


  andX
  g_g589_p
  (
    .dout(g589_p),
    .din1(g587_n_spl_),
    .din2(g588_n)
  );


  orX
  g_g589_n
  (
    .dout(g589_n),
    .din1(g587_p_spl_),
    .din2(g588_p)
  );


  andX
  g_g590_p
  (
    .dout(g590_p),
    .din1(g582_n_spl_),
    .din2(g589_p_spl_)
  );


  orX
  g_g590_n
  (
    .dout(g590_n),
    .din1(g582_p),
    .din2(g589_n)
  );


  orX
  g_g591_n
  (
    .dout(g591_n),
    .din1(g582_n_spl_),
    .din2(g589_p_spl_)
  );


  andX
  g_g592_p
  (
    .dout(g592_p),
    .din1(g590_n),
    .din2(g591_n)
  );


  andX
  g_g593_p
  (
    .dout(g593_p),
    .din1(g581_n_spl_),
    .din2(g592_p_spl_)
  );


  orX
  g_g594_n
  (
    .dout(g594_n),
    .din1(g590_p),
    .din2(g593_p_spl_)
  );


  andX
  g_g595_p
  (
    .dout(g595_p),
    .din1(ffc_29_p_spl_00),
    .din2(ffc_79_p_spl_)
  );


  orX
  g_g595_n
  (
    .dout(g595_n),
    .din1(ffc_29_n_spl_000),
    .din2(ffc_79_n_spl_)
  );


  andX
  g_g596_p
  (
    .dout(g596_p),
    .din1(g584_n_spl_),
    .din2(g587_n_spl_)
  );


  orX
  g_g596_n
  (
    .dout(g596_n),
    .din1(g584_p_spl_),
    .din2(g587_p_spl_)
  );


  andX
  g_g597_p
  (
    .dout(g597_p),
    .din1(ffc_25_p_spl_001),
    .din2(ffc_64_p_spl_)
  );


  orX
  g_g597_n
  (
    .dout(g597_n),
    .din1(ffc_25_n_spl_001),
    .din2(ffc_64_n_spl_)
  );


  andX
  g_g598_p
  (
    .dout(g598_p),
    .din1(ffc_268_n_spl_),
    .din2(ffc_276_n_spl_)
  );


  orX
  g_g598_n
  (
    .dout(g598_n),
    .din1(ffc_268_p_spl_),
    .din2(ffc_276_p_spl_)
  );


  andX
  g_g599_p
  (
    .dout(g599_p),
    .din1(ffc_268_p_spl_),
    .din2(ffc_276_p_spl_)
  );


  orX
  g_g599_n
  (
    .dout(g599_n),
    .din1(ffc_268_n_spl_),
    .din2(ffc_276_n_spl_)
  );


  andX
  g_g600_p
  (
    .dout(g600_p),
    .din1(g598_n_spl_),
    .din2(g599_n)
  );


  orX
  g_g600_n
  (
    .dout(g600_n),
    .din1(g598_p_spl_),
    .din2(g599_p)
  );


  andX
  g_g601_p
  (
    .dout(g601_p),
    .din1(g597_n_spl_),
    .din2(g600_p_spl_)
  );


  orX
  g_g601_n
  (
    .dout(g601_n),
    .din1(g597_p_spl_),
    .din2(g600_n_spl_)
  );


  andX
  g_g602_p
  (
    .dout(g602_p),
    .din1(g597_p_spl_),
    .din2(g600_n_spl_)
  );


  orX
  g_g602_n
  (
    .dout(g602_n),
    .din1(g597_n_spl_),
    .din2(g600_p_spl_)
  );


  andX
  g_g603_p
  (
    .dout(g603_p),
    .din1(g601_n_spl_),
    .din2(g602_n)
  );


  orX
  g_g603_n
  (
    .dout(g603_n),
    .din1(g601_p_spl_),
    .din2(g602_p)
  );


  andX
  g_g604_p
  (
    .dout(g604_p),
    .din1(g596_n_spl_),
    .din2(g603_p_spl_)
  );


  orX
  g_g604_n
  (
    .dout(g604_n),
    .din1(g596_p_spl_),
    .din2(g603_n_spl_)
  );


  andX
  g_g605_p
  (
    .dout(g605_p),
    .din1(g596_p_spl_),
    .din2(g603_n_spl_)
  );


  orX
  g_g605_n
  (
    .dout(g605_n),
    .din1(g596_n_spl_),
    .din2(g603_p_spl_)
  );


  andX
  g_g606_p
  (
    .dout(g606_p),
    .din1(g604_n_spl_),
    .din2(g605_n)
  );


  orX
  g_g606_n
  (
    .dout(g606_n),
    .din1(g604_p_spl_),
    .din2(g605_p)
  );


  andX
  g_g607_p
  (
    .dout(g607_p),
    .din1(g595_n_spl_),
    .din2(g606_p_spl_)
  );


  orX
  g_g607_n
  (
    .dout(g607_n),
    .din1(g595_p),
    .din2(g606_n)
  );


  orX
  g_g608_n
  (
    .dout(g608_n),
    .din1(g595_n_spl_),
    .din2(g606_p_spl_)
  );


  andX
  g_g609_p
  (
    .dout(g609_p),
    .din1(g607_n_spl_),
    .din2(g608_n)
  );


  orX
  g_g610_n
  (
    .dout(g610_n),
    .din1(g594_n_spl_),
    .din2(g609_p_spl_)
  );


  andX
  g_g611_p
  (
    .dout(g611_p),
    .din1(g604_n_spl_),
    .din2(g607_n_spl_)
  );


  orX
  g_g611_n
  (
    .dout(g611_n),
    .din1(g604_p_spl_),
    .din2(g607_p)
  );


  andX
  g_g612_p
  (
    .dout(g612_p),
    .din1(ffc_29_p_spl_00),
    .din2(ffc_64_p_spl_)
  );


  orX
  g_g612_n
  (
    .dout(g612_n),
    .din1(ffc_29_n_spl_00),
    .din2(ffc_64_n_spl_)
  );


  andX
  g_g613_p
  (
    .dout(g613_p),
    .din1(g598_n_spl_),
    .din2(g601_n_spl_)
  );


  orX
  g_g613_n
  (
    .dout(g613_n),
    .din1(g598_p_spl_),
    .din2(g601_p_spl_)
  );


  andX
  g_g614_p
  (
    .dout(g614_p),
    .din1(ffc_25_p_spl_001),
    .din2(ffc_65_p_spl_)
  );


  orX
  g_g614_n
  (
    .dout(g614_n),
    .din1(ffc_25_n_spl_001),
    .din2(ffc_65_n_spl_)
  );


  andX
  g_g615_p
  (
    .dout(g615_p),
    .din1(ffc_269_n_spl_),
    .din2(ffc_277_n_spl_)
  );


  orX
  g_g615_n
  (
    .dout(g615_n),
    .din1(ffc_269_p_spl_),
    .din2(ffc_277_p_spl_)
  );


  andX
  g_g616_p
  (
    .dout(g616_p),
    .din1(ffc_269_p_spl_),
    .din2(ffc_277_p_spl_)
  );


  orX
  g_g616_n
  (
    .dout(g616_n),
    .din1(ffc_269_n_spl_),
    .din2(ffc_277_n_spl_)
  );


  andX
  g_g617_p
  (
    .dout(g617_p),
    .din1(g615_n_spl_),
    .din2(g616_n)
  );


  orX
  g_g617_n
  (
    .dout(g617_n),
    .din1(g615_p_spl_),
    .din2(g616_p)
  );


  andX
  g_g618_p
  (
    .dout(g618_p),
    .din1(g614_n_spl_),
    .din2(g617_p_spl_)
  );


  orX
  g_g618_n
  (
    .dout(g618_n),
    .din1(g614_p_spl_),
    .din2(g617_n_spl_)
  );


  andX
  g_g619_p
  (
    .dout(g619_p),
    .din1(g614_p_spl_),
    .din2(g617_n_spl_)
  );


  orX
  g_g619_n
  (
    .dout(g619_n),
    .din1(g614_n_spl_),
    .din2(g617_p_spl_)
  );


  andX
  g_g620_p
  (
    .dout(g620_p),
    .din1(g618_n_spl_),
    .din2(g619_n)
  );


  orX
  g_g620_n
  (
    .dout(g620_n),
    .din1(g618_p_spl_),
    .din2(g619_p)
  );


  andX
  g_g621_p
  (
    .dout(g621_p),
    .din1(g613_n_spl_),
    .din2(g620_p_spl_)
  );


  orX
  g_g621_n
  (
    .dout(g621_n),
    .din1(g613_p_spl_),
    .din2(g620_n_spl_)
  );


  andX
  g_g622_p
  (
    .dout(g622_p),
    .din1(g613_p_spl_),
    .din2(g620_n_spl_)
  );


  orX
  g_g622_n
  (
    .dout(g622_n),
    .din1(g613_n_spl_),
    .din2(g620_p_spl_)
  );


  andX
  g_g623_p
  (
    .dout(g623_p),
    .din1(g621_n_spl_),
    .din2(g622_n)
  );


  orX
  g_g623_n
  (
    .dout(g623_n),
    .din1(g621_p_spl_),
    .din2(g622_p)
  );


  andX
  g_g624_p
  (
    .dout(g624_p),
    .din1(g612_n_spl_),
    .din2(g623_p_spl_)
  );


  orX
  g_g624_n
  (
    .dout(g624_n),
    .din1(g612_p_spl_),
    .din2(g623_n_spl_)
  );


  andX
  g_g625_p
  (
    .dout(g625_p),
    .din1(g612_p_spl_),
    .din2(g623_n_spl_)
  );


  orX
  g_g625_n
  (
    .dout(g625_n),
    .din1(g612_n_spl_),
    .din2(g623_p_spl_)
  );


  andX
  g_g626_p
  (
    .dout(g626_p),
    .din1(g624_n_spl_),
    .din2(g625_n)
  );


  orX
  g_g626_n
  (
    .dout(g626_n),
    .din1(g624_p_spl_),
    .din2(g625_p)
  );


  andX
  g_g627_p
  (
    .dout(g627_p),
    .din1(g611_n_spl_),
    .din2(g626_p_spl_)
  );


  orX
  g_g627_n
  (
    .dout(g627_n),
    .din1(g611_p),
    .din2(g626_n)
  );


  orX
  g_g628_n
  (
    .dout(g628_n),
    .din1(g611_n_spl_),
    .din2(g626_p_spl_)
  );


  andX
  g_g629_p
  (
    .dout(g629_p),
    .din1(g627_n),
    .din2(g628_n)
  );


  andX
  g_g630_p
  (
    .dout(g630_p),
    .din1(ffc_135_p_spl_00),
    .din2(ffc_287_p_spl_000)
  );


  orX
  g_g630_n
  (
    .dout(g630_n),
    .din1(ffc_135_n_spl_00),
    .din2(ffc_287_n_spl_000)
  );


  andX
  g_g631_p
  (
    .dout(g631_p),
    .din1(g610_n_spl_),
    .din2(g629_p_spl_)
  );


  andX
  g_g632_p
  (
    .dout(g632_p),
    .din1(ffc_285_n_spl_),
    .din2(ffc_286_n_spl_)
  );


  orX
  g_g632_n
  (
    .dout(g632_n),
    .din1(ffc_285_p_spl_),
    .din2(ffc_286_p_spl_)
  );


  andX
  g_g633_p
  (
    .dout(g633_p),
    .din1(ffc_285_p_spl_),
    .din2(ffc_286_p_spl_)
  );


  orX
  g_g633_n
  (
    .dout(g633_n),
    .din1(ffc_285_n_spl_),
    .din2(ffc_286_n_spl_)
  );


  andX
  g_g634_p
  (
    .dout(g634_p),
    .din1(g632_n_spl_),
    .din2(g633_n)
  );


  orX
  g_g634_n
  (
    .dout(g634_n),
    .din1(g632_p_spl_),
    .din2(g633_p)
  );


  andX
  g_g635_p
  (
    .dout(g635_p),
    .din1(g630_n),
    .din2(g634_p_spl_)
  );


  orX
  g_g635_n
  (
    .dout(g635_n),
    .din1(g630_p_spl_),
    .din2(g634_n)
  );


  orX
  g_g636_n
  (
    .dout(g636_n),
    .din1(g627_p),
    .din2(g631_p_spl_)
  );


  andX
  g_g637_p
  (
    .dout(g637_p),
    .din1(g621_n_spl_),
    .din2(g624_n_spl_)
  );


  orX
  g_g637_n
  (
    .dout(g637_n),
    .din1(g621_p_spl_),
    .din2(g624_p_spl_)
  );


  andX
  g_g638_p
  (
    .dout(g638_p),
    .din1(ffc_29_p_spl_01),
    .din2(ffc_65_p_spl_)
  );


  orX
  g_g638_n
  (
    .dout(g638_n),
    .din1(ffc_29_n_spl_01),
    .din2(ffc_65_n_spl_)
  );


  andX
  g_g639_p
  (
    .dout(g639_p),
    .din1(g615_n_spl_),
    .din2(g618_n_spl_)
  );


  orX
  g_g639_n
  (
    .dout(g639_n),
    .din1(g615_p_spl_),
    .din2(g618_p_spl_)
  );


  andX
  g_g640_p
  (
    .dout(g640_p),
    .din1(ffc_25_p_spl_010),
    .din2(ffc_66_p_spl_)
  );


  orX
  g_g640_n
  (
    .dout(g640_n),
    .din1(ffc_25_n_spl_010),
    .din2(ffc_66_n_spl_)
  );


  andX
  g_g641_p
  (
    .dout(g641_p),
    .din1(ffc_221_p),
    .din2(ffc_245_n)
  );


  orX
  g_g641_n
  (
    .dout(g641_n),
    .din1(ffc_221_n),
    .din2(ffc_245_p)
  );


  andX
  g_g642_p
  (
    .dout(g642_p),
    .din1(ffc_261_n_spl_),
    .din2(ffc_284_p_spl_)
  );


  orX
  g_g642_n
  (
    .dout(g642_n),
    .din1(ffc_261_p_spl_),
    .din2(ffc_284_n_spl_)
  );


  andX
  g_g643_p
  (
    .dout(g643_p),
    .din1(ffc_261_p_spl_),
    .din2(ffc_284_n_spl_)
  );


  orX
  g_g643_n
  (
    .dout(g643_n),
    .din1(ffc_261_n_spl_),
    .din2(ffc_284_p_spl_)
  );


  andX
  g_g644_p
  (
    .dout(g644_p),
    .din1(g642_n_spl_),
    .din2(g643_n)
  );


  orX
  g_g644_n
  (
    .dout(g644_n),
    .din1(g642_p_spl_),
    .din2(g643_p)
  );


  andX
  g_g645_p
  (
    .dout(g645_p),
    .din1(g641_n_spl_),
    .din2(g644_p_spl_)
  );


  orX
  g_g645_n
  (
    .dout(g645_n),
    .din1(g641_p_spl_),
    .din2(g644_n_spl_)
  );


  andX
  g_g646_p
  (
    .dout(g646_p),
    .din1(g641_p_spl_),
    .din2(g644_n_spl_)
  );


  orX
  g_g646_n
  (
    .dout(g646_n),
    .din1(g641_n_spl_),
    .din2(g644_p_spl_)
  );


  andX
  g_g647_p
  (
    .dout(g647_p),
    .din1(g645_n_spl_),
    .din2(g646_n)
  );


  orX
  g_g647_n
  (
    .dout(g647_n),
    .din1(g645_p_spl_),
    .din2(g646_p)
  );


  andX
  g_g648_p
  (
    .dout(g648_p),
    .din1(g640_n_spl_),
    .din2(g647_p_spl_)
  );


  orX
  g_g648_n
  (
    .dout(g648_n),
    .din1(g640_p_spl_),
    .din2(g647_n_spl_)
  );


  andX
  g_g649_p
  (
    .dout(g649_p),
    .din1(g640_p_spl_),
    .din2(g647_n_spl_)
  );


  orX
  g_g649_n
  (
    .dout(g649_n),
    .din1(g640_n_spl_),
    .din2(g647_p_spl_)
  );


  andX
  g_g650_p
  (
    .dout(g650_p),
    .din1(g648_n_spl_),
    .din2(g649_n)
  );


  orX
  g_g650_n
  (
    .dout(g650_n),
    .din1(g648_p_spl_),
    .din2(g649_p)
  );


  andX
  g_g651_p
  (
    .dout(g651_p),
    .din1(g639_n_spl_),
    .din2(g650_p_spl_)
  );


  orX
  g_g651_n
  (
    .dout(g651_n),
    .din1(g639_p_spl_),
    .din2(g650_n_spl_)
  );


  andX
  g_g652_p
  (
    .dout(g652_p),
    .din1(g639_p_spl_),
    .din2(g650_n_spl_)
  );


  orX
  g_g652_n
  (
    .dout(g652_n),
    .din1(g639_n_spl_),
    .din2(g650_p_spl_)
  );


  andX
  g_g653_p
  (
    .dout(g653_p),
    .din1(g651_n_spl_),
    .din2(g652_n)
  );


  orX
  g_g653_n
  (
    .dout(g653_n),
    .din1(g651_p_spl_),
    .din2(g652_p)
  );


  andX
  g_g654_p
  (
    .dout(g654_p),
    .din1(g638_n_spl_),
    .din2(g653_p_spl_)
  );


  orX
  g_g654_n
  (
    .dout(g654_n),
    .din1(g638_p_spl_),
    .din2(g653_n_spl_)
  );


  andX
  g_g655_p
  (
    .dout(g655_p),
    .din1(g638_p_spl_),
    .din2(g653_n_spl_)
  );


  orX
  g_g655_n
  (
    .dout(g655_n),
    .din1(g638_n_spl_),
    .din2(g653_p_spl_)
  );


  andX
  g_g656_p
  (
    .dout(g656_p),
    .din1(g654_n_spl_),
    .din2(g655_n)
  );


  orX
  g_g656_n
  (
    .dout(g656_n),
    .din1(g654_p_spl_),
    .din2(g655_p)
  );


  andX
  g_g657_p
  (
    .dout(g657_p),
    .din1(g637_n_spl_),
    .din2(g656_p_spl_)
  );


  orX
  g_g657_n
  (
    .dout(g657_n),
    .din1(g637_p),
    .din2(g656_n)
  );


  orX
  g_g658_n
  (
    .dout(g658_n),
    .din1(g637_n_spl_),
    .din2(g656_p_spl_)
  );


  andX
  g_g659_p
  (
    .dout(g659_p),
    .din1(g657_n),
    .din2(g658_n)
  );


  andX
  g_g660_p
  (
    .dout(g660_p),
    .din1(ffc_15_p_spl_000),
    .din2(ffc_135_p_spl_00)
  );


  orX
  g_g660_n
  (
    .dout(g660_n),
    .din1(ffc_15_n_spl_000),
    .din2(ffc_135_n_spl_00)
  );


  andX
  g_g661_p
  (
    .dout(g661_p),
    .din1(g636_n_spl_),
    .din2(g659_p_spl_)
  );


  andX
  g_g662_p
  (
    .dout(g662_p),
    .din1(g632_n_spl_),
    .din2(g635_n)
  );


  orX
  g_g662_n
  (
    .dout(g662_n),
    .din1(g632_p_spl_),
    .din2(g635_p_spl_)
  );


  andX
  g_g663_p
  (
    .dout(g663_p),
    .din1(ffc_133_p_spl_00),
    .din2(ffc_287_p_spl_000)
  );


  orX
  g_g663_n
  (
    .dout(g663_n),
    .din1(ffc_133_n_spl_00),
    .din2(ffc_287_n_spl_000)
  );


  andX
  g_g664_p
  (
    .dout(g664_p),
    .din1(ffc_310_p_spl_),
    .din2(ffc_311_n)
  );


  orX
  g_g664_n
  (
    .dout(g664_n),
    .din1(ffc_310_n_spl_),
    .din2(ffc_311_p)
  );


  andX
  g_g665_p
  (
    .dout(g665_p),
    .din1(g663_n_spl_),
    .din2(g664_p_spl_)
  );


  orX
  g_g665_n
  (
    .dout(g665_n),
    .din1(g663_p_spl_),
    .din2(g664_n_spl_)
  );


  andX
  g_g666_p
  (
    .dout(g666_p),
    .din1(g663_p_spl_),
    .din2(g664_n_spl_)
  );


  orX
  g_g666_n
  (
    .dout(g666_n),
    .din1(g663_n_spl_),
    .din2(g664_p_spl_)
  );


  andX
  g_g667_p
  (
    .dout(g667_p),
    .din1(g665_n_spl_),
    .din2(g666_n)
  );


  orX
  g_g667_n
  (
    .dout(g667_n),
    .din1(g665_p_spl_),
    .din2(g666_p)
  );


  andX
  g_g668_p
  (
    .dout(g668_p),
    .din1(g662_n_spl_),
    .din2(g667_p_spl_)
  );


  orX
  g_g668_n
  (
    .dout(g668_n),
    .din1(g662_p_spl_),
    .din2(g667_n_spl_)
  );


  andX
  g_g669_p
  (
    .dout(g669_p),
    .din1(g662_p_spl_),
    .din2(g667_n_spl_)
  );


  orX
  g_g669_n
  (
    .dout(g669_n),
    .din1(g662_n_spl_),
    .din2(g667_p_spl_)
  );


  andX
  g_g670_p
  (
    .dout(g670_p),
    .din1(g668_n_spl_),
    .din2(g669_n)
  );


  orX
  g_g670_n
  (
    .dout(g670_n),
    .din1(g668_p_spl_),
    .din2(g669_p)
  );


  andX
  g_g671_p
  (
    .dout(g671_p),
    .din1(g660_n),
    .din2(g670_p_spl_)
  );


  orX
  g_g671_n
  (
    .dout(g671_n),
    .din1(g660_p_spl_),
    .din2(g670_n)
  );


  andX
  g_g672_p
  (
    .dout(g672_p),
    .din1(ffc_207_p_spl_00),
    .din2(ffc_325_p_spl_0)
  );


  orX
  g_g672_n
  (
    .dout(g672_n),
    .din1(ffc_207_n_spl_00),
    .din2(ffc_325_n_spl_0)
  );


  andX
  g_g673_p
  (
    .dout(g673_p),
    .din1(ffc_341_p_spl_),
    .din2(ffc_342_n)
  );


  orX
  g_g673_n
  (
    .dout(g673_n),
    .din1(ffc_341_n_spl_),
    .din2(ffc_342_p)
  );


  orX
  g_g674_n
  (
    .dout(g674_n),
    .din1(g657_p),
    .din2(g661_p_spl_)
  );


  andX
  g_g675_p
  (
    .dout(g675_p),
    .din1(g651_n_spl_),
    .din2(g654_n_spl_)
  );


  orX
  g_g675_n
  (
    .dout(g675_n),
    .din1(g651_p_spl_),
    .din2(g654_p_spl_)
  );


  andX
  g_g676_p
  (
    .dout(g676_p),
    .din1(ffc_29_p_spl_01),
    .din2(ffc_66_p_spl_)
  );


  orX
  g_g676_n
  (
    .dout(g676_n),
    .din1(ffc_29_n_spl_01),
    .din2(ffc_66_n_spl_)
  );


  andX
  g_g677_p
  (
    .dout(g677_p),
    .din1(g645_n_spl_),
    .din2(g648_n_spl_)
  );


  orX
  g_g677_n
  (
    .dout(g677_n),
    .din1(g645_p_spl_),
    .din2(g648_p_spl_)
  );


  andX
  g_g678_p
  (
    .dout(g678_p),
    .din1(ffc_25_p_spl_010),
    .din2(ffc_67_p_spl_)
  );


  orX
  g_g678_n
  (
    .dout(g678_n),
    .din1(ffc_25_n_spl_010),
    .din2(ffc_67_n_spl_)
  );


  andX
  g_g679_p
  (
    .dout(g679_p),
    .din1(ffc_253_p),
    .din2(g642_n_spl_)
  );


  orX
  g_g679_n
  (
    .dout(g679_n),
    .din1(ffc_253_n),
    .din2(g642_p_spl_)
  );


  andX
  g_g680_p
  (
    .dout(g680_p),
    .din1(ffc_68_p_spl_0),
    .din2(ffc_214_p_spl_000)
  );


  orX
  g_g680_n
  (
    .dout(g680_n),
    .din1(ffc_68_n_spl_0),
    .din2(ffc_214_n_spl_000)
  );


  andX
  g_g681_p
  (
    .dout(g681_p),
    .din1(ffc_267_n_spl_),
    .din2(ffc_278_n_spl_)
  );


  orX
  g_g681_n
  (
    .dout(g681_n),
    .din1(ffc_267_p_spl_),
    .din2(ffc_278_p_spl_)
  );


  andX
  g_g682_p
  (
    .dout(g682_p),
    .din1(ffc_267_p_spl_),
    .din2(ffc_278_p_spl_)
  );


  orX
  g_g682_n
  (
    .dout(g682_n),
    .din1(ffc_267_n_spl_),
    .din2(ffc_278_n_spl_)
  );


  andX
  g_g683_p
  (
    .dout(g683_p),
    .din1(g681_n_spl_),
    .din2(g682_n)
  );


  orX
  g_g683_n
  (
    .dout(g683_n),
    .din1(g681_p_spl_),
    .din2(g682_p)
  );


  andX
  g_g684_p
  (
    .dout(g684_p),
    .din1(g680_n_spl_),
    .din2(g683_p_spl_)
  );


  orX
  g_g684_n
  (
    .dout(g684_n),
    .din1(g680_p_spl_),
    .din2(g683_n_spl_)
  );


  andX
  g_g685_p
  (
    .dout(g685_p),
    .din1(g680_p_spl_),
    .din2(g683_n_spl_)
  );


  orX
  g_g685_n
  (
    .dout(g685_n),
    .din1(g680_n_spl_),
    .din2(g683_p_spl_)
  );


  andX
  g_g686_p
  (
    .dout(g686_p),
    .din1(g684_n_spl_),
    .din2(g685_n)
  );


  orX
  g_g686_n
  (
    .dout(g686_n),
    .din1(g684_p_spl_),
    .din2(g685_p)
  );


  andX
  g_g687_p
  (
    .dout(g687_p),
    .din1(g679_n_spl_),
    .din2(g686_p_spl_)
  );


  orX
  g_g687_n
  (
    .dout(g687_n),
    .din1(g679_p_spl_),
    .din2(g686_n_spl_)
  );


  andX
  g_g688_p
  (
    .dout(g688_p),
    .din1(g679_p_spl_),
    .din2(g686_n_spl_)
  );


  orX
  g_g688_n
  (
    .dout(g688_n),
    .din1(g679_n_spl_),
    .din2(g686_p_spl_)
  );


  andX
  g_g689_p
  (
    .dout(g689_p),
    .din1(g687_n_spl_),
    .din2(g688_n)
  );


  orX
  g_g689_n
  (
    .dout(g689_n),
    .din1(g687_p_spl_),
    .din2(g688_p)
  );


  andX
  g_g690_p
  (
    .dout(g690_p),
    .din1(g678_n_spl_),
    .din2(g689_p_spl_)
  );


  orX
  g_g690_n
  (
    .dout(g690_n),
    .din1(g678_p_spl_),
    .din2(g689_n_spl_)
  );


  andX
  g_g691_p
  (
    .dout(g691_p),
    .din1(g678_p_spl_),
    .din2(g689_n_spl_)
  );


  orX
  g_g691_n
  (
    .dout(g691_n),
    .din1(g678_n_spl_),
    .din2(g689_p_spl_)
  );


  andX
  g_g692_p
  (
    .dout(g692_p),
    .din1(g690_n_spl_),
    .din2(g691_n)
  );


  orX
  g_g692_n
  (
    .dout(g692_n),
    .din1(g690_p_spl_),
    .din2(g691_p)
  );


  andX
  g_g693_p
  (
    .dout(g693_p),
    .din1(g677_n_spl_),
    .din2(g692_p_spl_)
  );


  orX
  g_g693_n
  (
    .dout(g693_n),
    .din1(g677_p_spl_),
    .din2(g692_n_spl_)
  );


  andX
  g_g694_p
  (
    .dout(g694_p),
    .din1(g677_p_spl_),
    .din2(g692_n_spl_)
  );


  orX
  g_g694_n
  (
    .dout(g694_n),
    .din1(g677_n_spl_),
    .din2(g692_p_spl_)
  );


  andX
  g_g695_p
  (
    .dout(g695_p),
    .din1(g693_n_spl_),
    .din2(g694_n)
  );


  orX
  g_g695_n
  (
    .dout(g695_n),
    .din1(g693_p_spl_),
    .din2(g694_p)
  );


  andX
  g_g696_p
  (
    .dout(g696_p),
    .din1(g676_n_spl_),
    .din2(g695_p_spl_)
  );


  orX
  g_g696_n
  (
    .dout(g696_n),
    .din1(g676_p_spl_),
    .din2(g695_n_spl_)
  );


  andX
  g_g697_p
  (
    .dout(g697_p),
    .din1(g676_p_spl_),
    .din2(g695_n_spl_)
  );


  orX
  g_g697_n
  (
    .dout(g697_n),
    .din1(g676_n_spl_),
    .din2(g695_p_spl_)
  );


  andX
  g_g698_p
  (
    .dout(g698_p),
    .din1(g696_n_spl_),
    .din2(g697_n)
  );


  orX
  g_g698_n
  (
    .dout(g698_n),
    .din1(g696_p_spl_),
    .din2(g697_p)
  );


  andX
  g_g699_p
  (
    .dout(g699_p),
    .din1(g675_n_spl_),
    .din2(g698_p_spl_)
  );


  orX
  g_g699_n
  (
    .dout(g699_n),
    .din1(g675_p),
    .din2(g698_n)
  );


  orX
  g_g700_n
  (
    .dout(g700_n),
    .din1(g675_n_spl_),
    .din2(g698_p_spl_)
  );


  andX
  g_g701_p
  (
    .dout(g701_p),
    .din1(g699_n),
    .din2(g700_n)
  );


  andX
  g_g702_p
  (
    .dout(g702_p),
    .din1(g672_n),
    .din2(g673_p_spl_)
  );


  orX
  g_g702_n
  (
    .dout(g702_n),
    .din1(g672_p_spl_),
    .din2(g673_n)
  );


  andX
  g_g703_p
  (
    .dout(g703_p),
    .din1(ffc_17_p_spl_000),
    .din2(ffc_135_p_spl_0)
  );


  orX
  g_g703_n
  (
    .dout(g703_n),
    .din1(ffc_17_n_spl_000),
    .din2(ffc_135_n_spl_0)
  );


  andX
  g_g704_p
  (
    .dout(g704_p),
    .din1(ffc_9_p_spl_000),
    .din2(ffc_207_p_spl_00)
  );


  orX
  g_g704_n
  (
    .dout(g704_n),
    .din1(ffc_9_n_spl_000),
    .din2(ffc_207_n_spl_00)
  );


  andX
  g_g705_p
  (
    .dout(g705_p),
    .din1(ffc_218_p),
    .din2(ffc_248_n)
  );


  orX
  g_g705_n
  (
    .dout(g705_n),
    .din1(ffc_218_n),
    .din2(ffc_248_p)
  );


  andX
  g_g706_p
  (
    .dout(g706_p),
    .din1(ffc_264_n_spl_),
    .din2(ffc_281_p_spl_)
  );


  orX
  g_g706_n
  (
    .dout(g706_n),
    .din1(ffc_264_p_spl_),
    .din2(ffc_281_n_spl_)
  );


  andX
  g_g707_p
  (
    .dout(g707_p),
    .din1(ffc_264_p_spl_),
    .din2(ffc_281_n_spl_)
  );


  orX
  g_g707_n
  (
    .dout(g707_n),
    .din1(ffc_264_n_spl_),
    .din2(ffc_281_p_spl_)
  );


  andX
  g_g708_p
  (
    .dout(g708_p),
    .din1(g706_n_spl_),
    .din2(g707_n)
  );


  orX
  g_g708_n
  (
    .dout(g708_n),
    .din1(g706_p_spl_),
    .din2(g707_p)
  );


  andX
  g_g709_p
  (
    .dout(g709_p),
    .din1(g705_n_spl_),
    .din2(g708_p_spl_)
  );


  orX
  g_g709_n
  (
    .dout(g709_n),
    .din1(g705_p_spl_),
    .din2(g708_n_spl_)
  );


  andX
  g_g710_p
  (
    .dout(g710_p),
    .din1(ffc_75_p_spl_0),
    .din2(ffc_160_p_spl_0)
  );


  orX
  g_g710_n
  (
    .dout(g710_n),
    .din1(ffc_75_n_spl_0),
    .din2(ffc_160_n_spl_0)
  );


  andX
  g_g711_p
  (
    .dout(g711_p),
    .din1(g705_p_spl_),
    .din2(g708_n_spl_)
  );


  orX
  g_g711_n
  (
    .dout(g711_n),
    .din1(g705_n_spl_),
    .din2(g708_p_spl_)
  );


  andX
  g_g712_p
  (
    .dout(g712_p),
    .din1(g709_n_spl_),
    .din2(g711_n)
  );


  orX
  g_g712_n
  (
    .dout(g712_n),
    .din1(g709_p_spl_),
    .din2(g711_p)
  );


  andX
  g_g713_p
  (
    .dout(g713_p),
    .din1(g710_n_spl_),
    .din2(g712_p_spl_)
  );


  orX
  g_g713_n
  (
    .dout(g713_n),
    .din1(g710_p_spl_),
    .din2(g712_n_spl_)
  );


  andX
  g_g714_p
  (
    .dout(g714_p),
    .din1(g709_n_spl_),
    .din2(g713_n_spl_)
  );


  orX
  g_g714_n
  (
    .dout(g714_n),
    .din1(g709_p_spl_),
    .din2(g713_p_spl_)
  );


  andX
  g_g715_p
  (
    .dout(g715_p),
    .din1(ffc_76_p_spl_0),
    .din2(ffc_160_p_spl_0)
  );


  orX
  g_g715_n
  (
    .dout(g715_n),
    .din1(ffc_76_n_spl_0),
    .din2(ffc_160_n_spl_0)
  );


  andX
  g_g716_p
  (
    .dout(g716_p),
    .din1(ffc_77_p_spl_0),
    .din2(ffc_148_p)
  );


  orX
  g_g716_n
  (
    .dout(g716_n),
    .din1(ffc_77_n_spl_0),
    .din2(ffc_148_n)
  );


  andX
  g_g717_p
  (
    .dout(g717_p),
    .din1(ffc_249_p),
    .din2(g706_n_spl_)
  );


  orX
  g_g717_n
  (
    .dout(g717_n),
    .din1(ffc_249_n),
    .din2(g706_p_spl_)
  );


  andX
  g_g718_p
  (
    .dout(g718_p),
    .din1(g716_n_spl_),
    .din2(g717_n_spl_)
  );


  orX
  g_g718_n
  (
    .dout(g718_n),
    .din1(g716_p_spl_),
    .din2(g717_p_spl_)
  );


  andX
  g_g719_p
  (
    .dout(g719_p),
    .din1(g716_p_spl_),
    .din2(g717_p_spl_)
  );


  orX
  g_g719_n
  (
    .dout(g719_n),
    .din1(g716_n_spl_),
    .din2(g717_n_spl_)
  );


  andX
  g_g720_p
  (
    .dout(g720_p),
    .din1(g718_n_spl_),
    .din2(g719_n)
  );


  orX
  g_g720_n
  (
    .dout(g720_n),
    .din1(g718_p_spl_),
    .din2(g719_p)
  );


  andX
  g_g721_p
  (
    .dout(g721_p),
    .din1(g715_n_spl_),
    .din2(g720_p_spl_)
  );


  orX
  g_g721_n
  (
    .dout(g721_n),
    .din1(g715_p_spl_),
    .din2(g720_n_spl_)
  );


  andX
  g_g722_p
  (
    .dout(g722_p),
    .din1(g715_p_spl_),
    .din2(g720_n_spl_)
  );


  orX
  g_g722_n
  (
    .dout(g722_n),
    .din1(g715_n_spl_),
    .din2(g720_p_spl_)
  );


  andX
  g_g723_p
  (
    .dout(g723_p),
    .din1(g721_n_spl_),
    .din2(g722_n)
  );


  orX
  g_g723_n
  (
    .dout(g723_n),
    .din1(g721_p_spl_),
    .din2(g722_p)
  );


  andX
  g_g724_p
  (
    .dout(g724_p),
    .din1(g714_n_spl_),
    .din2(g723_p_spl_)
  );


  orX
  g_g724_n
  (
    .dout(g724_n),
    .din1(g714_p_spl_),
    .din2(g723_n_spl_)
  );


  andX
  g_g725_p
  (
    .dout(g725_p),
    .din1(ffc_75_p_spl_0),
    .din2(ffc_174_p_spl_00)
  );


  orX
  g_g725_n
  (
    .dout(g725_n),
    .din1(ffc_75_n_spl_0),
    .din2(ffc_174_n_spl_00)
  );


  andX
  g_g726_p
  (
    .dout(g726_p),
    .din1(g714_p_spl_),
    .din2(g723_n_spl_)
  );


  orX
  g_g726_n
  (
    .dout(g726_n),
    .din1(g714_n_spl_),
    .din2(g723_p_spl_)
  );


  andX
  g_g727_p
  (
    .dout(g727_p),
    .din1(g724_n_spl_),
    .din2(g726_n)
  );


  orX
  g_g727_n
  (
    .dout(g727_n),
    .din1(g724_p_spl_),
    .din2(g726_p)
  );


  andX
  g_g728_p
  (
    .dout(g728_p),
    .din1(g725_n_spl_),
    .din2(g727_p_spl_)
  );


  orX
  g_g728_n
  (
    .dout(g728_n),
    .din1(g725_p_spl_),
    .din2(g727_n_spl_)
  );


  andX
  g_g729_p
  (
    .dout(g729_p),
    .din1(g724_n_spl_),
    .din2(g728_n_spl_)
  );


  orX
  g_g729_n
  (
    .dout(g729_n),
    .din1(g724_p_spl_),
    .din2(g728_p_spl_)
  );


  andX
  g_g730_p
  (
    .dout(g730_p),
    .din1(ffc_76_p_spl_0),
    .din2(ffc_174_p_spl_00)
  );


  orX
  g_g730_n
  (
    .dout(g730_n),
    .din1(ffc_76_n_spl_0),
    .din2(ffc_174_n_spl_00)
  );


  andX
  g_g731_p
  (
    .dout(g731_p),
    .din1(ffc_77_p_spl_0),
    .din2(ffc_160_p_spl_1)
  );


  orX
  g_g731_n
  (
    .dout(g731_n),
    .din1(ffc_77_n_spl_0),
    .din2(ffc_160_n_spl_1)
  );


  andX
  g_g732_p
  (
    .dout(g732_p),
    .din1(g718_n_spl_),
    .din2(g721_n_spl_)
  );


  orX
  g_g732_n
  (
    .dout(g732_n),
    .din1(g718_p_spl_),
    .din2(g721_p_spl_)
  );


  andX
  g_g733_p
  (
    .dout(g733_p),
    .din1(g731_n_spl_),
    .din2(g732_n_spl_)
  );


  orX
  g_g733_n
  (
    .dout(g733_n),
    .din1(g731_p_spl_),
    .din2(g732_p_spl_)
  );


  andX
  g_g734_p
  (
    .dout(g734_p),
    .din1(g731_p_spl_),
    .din2(g732_p_spl_)
  );


  orX
  g_g734_n
  (
    .dout(g734_n),
    .din1(g731_n_spl_),
    .din2(g732_n_spl_)
  );


  andX
  g_g735_p
  (
    .dout(g735_p),
    .din1(g733_n_spl_),
    .din2(g734_n)
  );


  orX
  g_g735_n
  (
    .dout(g735_n),
    .din1(g733_p_spl_),
    .din2(g734_p)
  );


  andX
  g_g736_p
  (
    .dout(g736_p),
    .din1(g730_n_spl_),
    .din2(g735_p_spl_)
  );


  orX
  g_g736_n
  (
    .dout(g736_n),
    .din1(g730_p_spl_),
    .din2(g735_n_spl_)
  );


  andX
  g_g737_p
  (
    .dout(g737_p),
    .din1(g730_p_spl_),
    .din2(g735_n_spl_)
  );


  orX
  g_g737_n
  (
    .dout(g737_n),
    .din1(g730_n_spl_),
    .din2(g735_p_spl_)
  );


  andX
  g_g738_p
  (
    .dout(g738_p),
    .din1(g736_n_spl_),
    .din2(g737_n)
  );


  orX
  g_g738_n
  (
    .dout(g738_n),
    .din1(g736_p_spl_),
    .din2(g737_p)
  );


  andX
  g_g739_p
  (
    .dout(g739_p),
    .din1(g729_n_spl_),
    .din2(g738_p_spl_)
  );


  orX
  g_g739_n
  (
    .dout(g739_n),
    .din1(g729_p_spl_),
    .din2(g738_n_spl_)
  );


  andX
  g_g740_p
  (
    .dout(g740_p),
    .din1(ffc_219_p),
    .din2(ffc_247_n)
  );


  orX
  g_g740_n
  (
    .dout(g740_n),
    .din1(ffc_219_n),
    .din2(ffc_247_p)
  );


  andX
  g_g741_p
  (
    .dout(g741_p),
    .din1(ffc_263_n_spl_),
    .din2(ffc_282_p_spl_)
  );


  orX
  g_g741_n
  (
    .dout(g741_n),
    .din1(ffc_263_p_spl_),
    .din2(ffc_282_n_spl_)
  );


  andX
  g_g742_p
  (
    .dout(g742_p),
    .din1(ffc_263_p_spl_),
    .din2(ffc_282_n_spl_)
  );


  orX
  g_g742_n
  (
    .dout(g742_n),
    .din1(ffc_263_n_spl_),
    .din2(ffc_282_p_spl_)
  );


  andX
  g_g743_p
  (
    .dout(g743_p),
    .din1(g741_n_spl_),
    .din2(g742_n)
  );


  orX
  g_g743_n
  (
    .dout(g743_n),
    .din1(g741_p_spl_),
    .din2(g742_p)
  );


  andX
  g_g744_p
  (
    .dout(g744_p),
    .din1(g740_n_spl_),
    .din2(g743_p_spl_)
  );


  orX
  g_g744_n
  (
    .dout(g744_n),
    .din1(g740_p_spl_),
    .din2(g743_n_spl_)
  );


  andX
  g_g745_p
  (
    .dout(g745_p),
    .din1(ffc_72_p_spl_0),
    .din2(ffc_174_p_spl_01)
  );


  orX
  g_g745_n
  (
    .dout(g745_n),
    .din1(ffc_72_n_spl_0),
    .din2(ffc_174_n_spl_01)
  );


  andX
  g_g746_p
  (
    .dout(g746_p),
    .din1(g740_p_spl_),
    .din2(g743_n_spl_)
  );


  orX
  g_g746_n
  (
    .dout(g746_n),
    .din1(g740_n_spl_),
    .din2(g743_p_spl_)
  );


  andX
  g_g747_p
  (
    .dout(g747_p),
    .din1(g744_n_spl_),
    .din2(g746_n)
  );


  orX
  g_g747_n
  (
    .dout(g747_n),
    .din1(g744_p_spl_),
    .din2(g746_p)
  );


  andX
  g_g748_p
  (
    .dout(g748_p),
    .din1(g745_n_spl_),
    .din2(g747_p_spl_)
  );


  orX
  g_g748_n
  (
    .dout(g748_n),
    .din1(g745_p_spl_),
    .din2(g747_n_spl_)
  );


  andX
  g_g749_p
  (
    .dout(g749_p),
    .din1(g744_n_spl_),
    .din2(g748_n_spl_)
  );


  orX
  g_g749_n
  (
    .dout(g749_n),
    .din1(g744_p_spl_),
    .din2(g748_p_spl_)
  );


  andX
  g_g750_p
  (
    .dout(g750_p),
    .din1(ffc_73_p_spl_0),
    .din2(ffc_174_p_spl_01)
  );


  orX
  g_g750_n
  (
    .dout(g750_n),
    .din1(ffc_73_n_spl_0),
    .din2(ffc_174_n_spl_01)
  );


  andX
  g_g751_p
  (
    .dout(g751_p),
    .din1(ffc_251_p),
    .din2(g741_n_spl_)
  );


  orX
  g_g751_n
  (
    .dout(g751_n),
    .din1(ffc_251_n),
    .din2(g741_p_spl_)
  );


  andX
  g_g752_p
  (
    .dout(g752_p),
    .din1(ffc_74_p_spl_0),
    .din2(ffc_160_p_spl_1)
  );


  orX
  g_g752_n
  (
    .dout(g752_n),
    .din1(ffc_74_n_spl_0),
    .din2(ffc_160_n_spl_1)
  );


  andX
  g_g753_p
  (
    .dout(g753_p),
    .din1(ffc_265_n_spl_),
    .din2(ffc_280_n_spl_)
  );


  orX
  g_g753_n
  (
    .dout(g753_n),
    .din1(ffc_265_p_spl_),
    .din2(ffc_280_p_spl_)
  );


  andX
  g_g754_p
  (
    .dout(g754_p),
    .din1(ffc_265_p_spl_),
    .din2(ffc_280_p_spl_)
  );


  orX
  g_g754_n
  (
    .dout(g754_n),
    .din1(ffc_265_n_spl_),
    .din2(ffc_280_n_spl_)
  );


  andX
  g_g755_p
  (
    .dout(g755_p),
    .din1(g753_n_spl_),
    .din2(g754_n)
  );


  orX
  g_g755_n
  (
    .dout(g755_n),
    .din1(g753_p_spl_),
    .din2(g754_p)
  );


  andX
  g_g756_p
  (
    .dout(g756_p),
    .din1(g752_n_spl_),
    .din2(g755_p_spl_)
  );


  orX
  g_g756_n
  (
    .dout(g756_n),
    .din1(g752_p_spl_),
    .din2(g755_n_spl_)
  );


  andX
  g_g757_p
  (
    .dout(g757_p),
    .din1(g752_p_spl_),
    .din2(g755_n_spl_)
  );


  orX
  g_g757_n
  (
    .dout(g757_n),
    .din1(g752_n_spl_),
    .din2(g755_p_spl_)
  );


  andX
  g_g758_p
  (
    .dout(g758_p),
    .din1(g756_n_spl_),
    .din2(g757_n)
  );


  orX
  g_g758_n
  (
    .dout(g758_n),
    .din1(g756_p_spl_),
    .din2(g757_p)
  );


  andX
  g_g759_p
  (
    .dout(g759_p),
    .din1(g751_n_spl_),
    .din2(g758_p_spl_)
  );


  orX
  g_g759_n
  (
    .dout(g759_n),
    .din1(g751_p_spl_),
    .din2(g758_n_spl_)
  );


  andX
  g_g760_p
  (
    .dout(g760_p),
    .din1(g751_p_spl_),
    .din2(g758_n_spl_)
  );


  orX
  g_g760_n
  (
    .dout(g760_n),
    .din1(g751_n_spl_),
    .din2(g758_p_spl_)
  );


  andX
  g_g761_p
  (
    .dout(g761_p),
    .din1(g759_n_spl_),
    .din2(g760_n)
  );


  orX
  g_g761_n
  (
    .dout(g761_n),
    .din1(g759_p_spl_),
    .din2(g760_p)
  );


  andX
  g_g762_p
  (
    .dout(g762_p),
    .din1(g750_n_spl_),
    .din2(g761_p_spl_)
  );


  orX
  g_g762_n
  (
    .dout(g762_n),
    .din1(g750_p_spl_),
    .din2(g761_n_spl_)
  );


  andX
  g_g763_p
  (
    .dout(g763_p),
    .din1(g750_p_spl_),
    .din2(g761_n_spl_)
  );


  orX
  g_g763_n
  (
    .dout(g763_n),
    .din1(g750_n_spl_),
    .din2(g761_p_spl_)
  );


  andX
  g_g764_p
  (
    .dout(g764_p),
    .din1(g762_n_spl_),
    .din2(g763_n)
  );


  orX
  g_g764_n
  (
    .dout(g764_n),
    .din1(g762_p_spl_),
    .din2(g763_p)
  );


  andX
  g_g765_p
  (
    .dout(g765_p),
    .din1(g749_n_spl_),
    .din2(g764_p_spl_)
  );


  orX
  g_g765_n
  (
    .dout(g765_n),
    .din1(g749_p_spl_),
    .din2(g764_n_spl_)
  );


  andX
  g_g766_p
  (
    .dout(g766_p),
    .din1(ffc_72_p_spl_0),
    .din2(ffc_214_p_spl_000)
  );


  orX
  g_g766_n
  (
    .dout(g766_n),
    .din1(ffc_72_n_spl_0),
    .din2(ffc_214_n_spl_000)
  );


  andX
  g_g767_p
  (
    .dout(g767_p),
    .din1(g749_p_spl_),
    .din2(g764_n_spl_)
  );


  orX
  g_g767_n
  (
    .dout(g767_n),
    .din1(g749_n_spl_),
    .din2(g764_p_spl_)
  );


  andX
  g_g768_p
  (
    .dout(g768_p),
    .din1(g765_n_spl_),
    .din2(g767_n)
  );


  orX
  g_g768_n
  (
    .dout(g768_n),
    .din1(g765_p_spl_),
    .din2(g767_p)
  );


  andX
  g_g769_p
  (
    .dout(g769_p),
    .din1(g766_n_spl_),
    .din2(g768_p_spl_)
  );


  orX
  g_g769_n
  (
    .dout(g769_n),
    .din1(g766_p_spl_),
    .din2(g768_n_spl_)
  );


  andX
  g_g770_p
  (
    .dout(g770_p),
    .din1(g765_n_spl_),
    .din2(g769_n_spl_)
  );


  orX
  g_g770_n
  (
    .dout(g770_n),
    .din1(g765_p_spl_),
    .din2(g769_p_spl_)
  );


  andX
  g_g771_p
  (
    .dout(g771_p),
    .din1(ffc_73_p_spl_0),
    .din2(ffc_214_p_spl_00)
  );


  orX
  g_g771_n
  (
    .dout(g771_n),
    .din1(ffc_73_n_spl_0),
    .din2(ffc_214_n_spl_00)
  );


  andX
  g_g772_p
  (
    .dout(g772_p),
    .din1(g759_n_spl_),
    .din2(g762_n_spl_)
  );


  orX
  g_g772_n
  (
    .dout(g772_n),
    .din1(g759_p_spl_),
    .din2(g762_p_spl_)
  );


  andX
  g_g773_p
  (
    .dout(g773_p),
    .din1(ffc_74_p_spl_0),
    .din2(ffc_174_p_spl_10)
  );


  orX
  g_g773_n
  (
    .dout(g773_n),
    .din1(ffc_74_n_spl_0),
    .din2(ffc_174_n_spl_10)
  );


  andX
  g_g774_p
  (
    .dout(g774_p),
    .din1(g753_n_spl_),
    .din2(g756_n_spl_)
  );


  orX
  g_g774_n
  (
    .dout(g774_n),
    .din1(g753_p_spl_),
    .din2(g756_p_spl_)
  );


  andX
  g_g775_p
  (
    .dout(g775_p),
    .din1(g710_p_spl_),
    .din2(g712_n_spl_)
  );


  orX
  g_g775_n
  (
    .dout(g775_n),
    .din1(g710_n_spl_),
    .din2(g712_p_spl_)
  );


  andX
  g_g776_p
  (
    .dout(g776_p),
    .din1(g713_n_spl_),
    .din2(g775_n)
  );


  orX
  g_g776_n
  (
    .dout(g776_n),
    .din1(g713_p_spl_),
    .din2(g775_p)
  );


  andX
  g_g777_p
  (
    .dout(g777_p),
    .din1(g774_n_spl_),
    .din2(g776_p_spl_)
  );


  orX
  g_g777_n
  (
    .dout(g777_n),
    .din1(g774_p_spl_),
    .din2(g776_n_spl_)
  );


  andX
  g_g778_p
  (
    .dout(g778_p),
    .din1(g774_p_spl_),
    .din2(g776_n_spl_)
  );


  orX
  g_g778_n
  (
    .dout(g778_n),
    .din1(g774_n_spl_),
    .din2(g776_p_spl_)
  );


  andX
  g_g779_p
  (
    .dout(g779_p),
    .din1(g777_n_spl_),
    .din2(g778_n)
  );


  orX
  g_g779_n
  (
    .dout(g779_n),
    .din1(g777_p_spl_),
    .din2(g778_p)
  );


  andX
  g_g780_p
  (
    .dout(g780_p),
    .din1(g773_n_spl_),
    .din2(g779_p_spl_)
  );


  orX
  g_g780_n
  (
    .dout(g780_n),
    .din1(g773_p_spl_),
    .din2(g779_n_spl_)
  );


  andX
  g_g781_p
  (
    .dout(g781_p),
    .din1(g773_p_spl_),
    .din2(g779_n_spl_)
  );


  orX
  g_g781_n
  (
    .dout(g781_n),
    .din1(g773_n_spl_),
    .din2(g779_p_spl_)
  );


  andX
  g_g782_p
  (
    .dout(g782_p),
    .din1(g780_n_spl_),
    .din2(g781_n)
  );


  orX
  g_g782_n
  (
    .dout(g782_n),
    .din1(g780_p_spl_),
    .din2(g781_p)
  );


  andX
  g_g783_p
  (
    .dout(g783_p),
    .din1(g772_n_spl_),
    .din2(g782_p_spl_)
  );


  orX
  g_g783_n
  (
    .dout(g783_n),
    .din1(g772_p_spl_),
    .din2(g782_n_spl_)
  );


  andX
  g_g784_p
  (
    .dout(g784_p),
    .din1(g772_p_spl_),
    .din2(g782_n_spl_)
  );


  orX
  g_g784_n
  (
    .dout(g784_n),
    .din1(g772_n_spl_),
    .din2(g782_p_spl_)
  );


  andX
  g_g785_p
  (
    .dout(g785_p),
    .din1(g783_n_spl_),
    .din2(g784_n)
  );


  orX
  g_g785_n
  (
    .dout(g785_n),
    .din1(g783_p_spl_),
    .din2(g784_p)
  );


  andX
  g_g786_p
  (
    .dout(g786_p),
    .din1(g771_n_spl_),
    .din2(g785_p_spl_)
  );


  orX
  g_g786_n
  (
    .dout(g786_n),
    .din1(g771_p_spl_),
    .din2(g785_n_spl_)
  );


  andX
  g_g787_p
  (
    .dout(g787_p),
    .din1(g771_p_spl_),
    .din2(g785_n_spl_)
  );


  orX
  g_g787_n
  (
    .dout(g787_n),
    .din1(g771_n_spl_),
    .din2(g785_p_spl_)
  );


  andX
  g_g788_p
  (
    .dout(g788_p),
    .din1(g786_n_spl_),
    .din2(g787_n)
  );


  orX
  g_g788_n
  (
    .dout(g788_n),
    .din1(g786_p_spl_),
    .din2(g787_p)
  );


  andX
  g_g789_p
  (
    .dout(g789_p),
    .din1(g770_n_spl_),
    .din2(g788_p_spl_)
  );


  orX
  g_g789_n
  (
    .dout(g789_n),
    .din1(g770_p_spl_),
    .din2(g788_n_spl_)
  );


  andX
  g_g790_p
  (
    .dout(g790_p),
    .din1(ffc_220_p),
    .din2(ffc_246_n)
  );


  orX
  g_g790_n
  (
    .dout(g790_n),
    .din1(ffc_220_n),
    .din2(ffc_246_p)
  );


  andX
  g_g791_p
  (
    .dout(g791_p),
    .din1(ffc_262_n_spl_),
    .din2(ffc_283_p_spl_)
  );


  orX
  g_g791_n
  (
    .dout(g791_n),
    .din1(ffc_262_p_spl_),
    .din2(ffc_283_n_spl_)
  );


  andX
  g_g792_p
  (
    .dout(g792_p),
    .din1(ffc_262_p_spl_),
    .din2(ffc_283_n_spl_)
  );


  orX
  g_g792_n
  (
    .dout(g792_n),
    .din1(ffc_262_n_spl_),
    .din2(ffc_283_p_spl_)
  );


  andX
  g_g793_p
  (
    .dout(g793_p),
    .din1(g791_n_spl_),
    .din2(g792_n)
  );


  orX
  g_g793_n
  (
    .dout(g793_n),
    .din1(g791_p_spl_),
    .din2(g792_p)
  );


  andX
  g_g794_p
  (
    .dout(g794_p),
    .din1(g790_n_spl_),
    .din2(g793_p_spl_)
  );


  orX
  g_g794_n
  (
    .dout(g794_n),
    .din1(g790_p_spl_),
    .din2(g793_n_spl_)
  );


  andX
  g_g795_p
  (
    .dout(g795_p),
    .din1(ffc_69_p_spl_0),
    .din2(ffc_214_p_spl_01)
  );


  orX
  g_g795_n
  (
    .dout(g795_n),
    .din1(ffc_69_n_spl_0),
    .din2(ffc_214_n_spl_01)
  );


  andX
  g_g796_p
  (
    .dout(g796_p),
    .din1(g790_p_spl_),
    .din2(g793_n_spl_)
  );


  orX
  g_g796_n
  (
    .dout(g796_n),
    .din1(g790_n_spl_),
    .din2(g793_p_spl_)
  );


  andX
  g_g797_p
  (
    .dout(g797_p),
    .din1(g794_n_spl_),
    .din2(g796_n)
  );


  orX
  g_g797_n
  (
    .dout(g797_n),
    .din1(g794_p_spl_),
    .din2(g796_p)
  );


  andX
  g_g798_p
  (
    .dout(g798_p),
    .din1(g795_n_spl_),
    .din2(g797_p_spl_)
  );


  orX
  g_g798_n
  (
    .dout(g798_n),
    .din1(g795_p_spl_),
    .din2(g797_n_spl_)
  );


  andX
  g_g799_p
  (
    .dout(g799_p),
    .din1(g794_n_spl_),
    .din2(g798_n_spl_)
  );


  orX
  g_g799_n
  (
    .dout(g799_n),
    .din1(g794_p_spl_),
    .din2(g798_p_spl_)
  );


  andX
  g_g800_p
  (
    .dout(g800_p),
    .din1(ffc_70_p_spl_),
    .din2(ffc_214_p_spl_01)
  );


  orX
  g_g800_n
  (
    .dout(g800_n),
    .din1(ffc_70_n_spl_0),
    .din2(ffc_214_n_spl_01)
  );


  andX
  g_g801_p
  (
    .dout(g801_p),
    .din1(ffc_252_p),
    .din2(g791_n_spl_)
  );


  orX
  g_g801_n
  (
    .dout(g801_n),
    .din1(ffc_252_n),
    .din2(g791_p_spl_)
  );


  andX
  g_g802_p
  (
    .dout(g802_p),
    .din1(ffc_71_p_spl_0),
    .din2(ffc_174_p_spl_10)
  );


  orX
  g_g802_n
  (
    .dout(g802_n),
    .din1(ffc_71_n_spl_0),
    .din2(ffc_174_n_spl_10)
  );


  andX
  g_g803_p
  (
    .dout(g803_p),
    .din1(ffc_266_n_spl_),
    .din2(ffc_279_n_spl_)
  );


  orX
  g_g803_n
  (
    .dout(g803_n),
    .din1(ffc_266_p_spl_),
    .din2(ffc_279_p_spl_)
  );


  andX
  g_g804_p
  (
    .dout(g804_p),
    .din1(ffc_266_p_spl_),
    .din2(ffc_279_p_spl_)
  );


  orX
  g_g804_n
  (
    .dout(g804_n),
    .din1(ffc_266_n_spl_),
    .din2(ffc_279_n_spl_)
  );


  andX
  g_g805_p
  (
    .dout(g805_p),
    .din1(g803_n_spl_),
    .din2(g804_n)
  );


  orX
  g_g805_n
  (
    .dout(g805_n),
    .din1(g803_p_spl_),
    .din2(g804_p)
  );


  andX
  g_g806_p
  (
    .dout(g806_p),
    .din1(g802_n_spl_),
    .din2(g805_p_spl_)
  );


  orX
  g_g806_n
  (
    .dout(g806_n),
    .din1(g802_p_spl_),
    .din2(g805_n_spl_)
  );


  andX
  g_g807_p
  (
    .dout(g807_p),
    .din1(g802_p_spl_),
    .din2(g805_n_spl_)
  );


  orX
  g_g807_n
  (
    .dout(g807_n),
    .din1(g802_n_spl_),
    .din2(g805_p_spl_)
  );


  andX
  g_g808_p
  (
    .dout(g808_p),
    .din1(g806_n_spl_),
    .din2(g807_n)
  );


  orX
  g_g808_n
  (
    .dout(g808_n),
    .din1(g806_p_spl_),
    .din2(g807_p)
  );


  andX
  g_g809_p
  (
    .dout(g809_p),
    .din1(g801_n_spl_),
    .din2(g808_p_spl_)
  );


  orX
  g_g809_n
  (
    .dout(g809_n),
    .din1(g801_p_spl_),
    .din2(g808_n_spl_)
  );


  andX
  g_g810_p
  (
    .dout(g810_p),
    .din1(g801_p_spl_),
    .din2(g808_n_spl_)
  );


  orX
  g_g810_n
  (
    .dout(g810_n),
    .din1(g801_n_spl_),
    .din2(g808_p_spl_)
  );


  andX
  g_g811_p
  (
    .dout(g811_p),
    .din1(g809_n_spl_),
    .din2(g810_n)
  );


  orX
  g_g811_n
  (
    .dout(g811_n),
    .din1(g809_p_spl_),
    .din2(g810_p)
  );


  andX
  g_g812_p
  (
    .dout(g812_p),
    .din1(g800_n_spl_),
    .din2(g811_p_spl_)
  );


  orX
  g_g812_n
  (
    .dout(g812_n),
    .din1(g800_p_spl_),
    .din2(g811_n_spl_)
  );


  andX
  g_g813_p
  (
    .dout(g813_p),
    .din1(g800_p_spl_),
    .din2(g811_n_spl_)
  );


  orX
  g_g813_n
  (
    .dout(g813_n),
    .din1(g800_n_spl_),
    .din2(g811_p_spl_)
  );


  andX
  g_g814_p
  (
    .dout(g814_p),
    .din1(g812_n_spl_),
    .din2(g813_n)
  );


  orX
  g_g814_n
  (
    .dout(g814_n),
    .din1(g812_p_spl_),
    .din2(g813_p)
  );


  andX
  g_g815_p
  (
    .dout(g815_p),
    .din1(g799_n_spl_),
    .din2(g814_p_spl_)
  );


  orX
  g_g815_n
  (
    .dout(g815_n),
    .din1(g799_p_spl_),
    .din2(g814_n_spl_)
  );


  andX
  g_g816_p
  (
    .dout(g816_p),
    .din1(ffc_25_p_spl_011),
    .din2(ffc_69_p_spl_0)
  );


  orX
  g_g816_n
  (
    .dout(g816_n),
    .din1(ffc_25_n_spl_011),
    .din2(ffc_69_n_spl_0)
  );


  andX
  g_g817_p
  (
    .dout(g817_p),
    .din1(g799_p_spl_),
    .din2(g814_n_spl_)
  );


  orX
  g_g817_n
  (
    .dout(g817_n),
    .din1(g799_n_spl_),
    .din2(g814_p_spl_)
  );


  andX
  g_g818_p
  (
    .dout(g818_p),
    .din1(g815_n_spl_),
    .din2(g817_n)
  );


  orX
  g_g818_n
  (
    .dout(g818_n),
    .din1(g815_p_spl_),
    .din2(g817_p)
  );


  andX
  g_g819_p
  (
    .dout(g819_p),
    .din1(g816_n_spl_),
    .din2(g818_p_spl_)
  );


  orX
  g_g819_n
  (
    .dout(g819_n),
    .din1(g816_p_spl_),
    .din2(g818_n_spl_)
  );


  andX
  g_g820_p
  (
    .dout(g820_p),
    .din1(g815_n_spl_),
    .din2(g819_n_spl_)
  );


  orX
  g_g820_n
  (
    .dout(g820_n),
    .din1(g815_p_spl_),
    .din2(g819_p_spl_)
  );


  andX
  g_g821_p
  (
    .dout(g821_p),
    .din1(ffc_25_p_spl_011),
    .din2(ffc_70_p_spl_)
  );


  orX
  g_g821_n
  (
    .dout(g821_n),
    .din1(ffc_25_n_spl_011),
    .din2(ffc_70_n_spl_0)
  );


  andX
  g_g822_p
  (
    .dout(g822_p),
    .din1(g809_n_spl_),
    .din2(g812_n_spl_)
  );


  orX
  g_g822_n
  (
    .dout(g822_n),
    .din1(g809_p_spl_),
    .din2(g812_p_spl_)
  );


  andX
  g_g823_p
  (
    .dout(g823_p),
    .din1(ffc_71_p_spl_0),
    .din2(ffc_214_p_spl_10)
  );


  orX
  g_g823_n
  (
    .dout(g823_n),
    .din1(ffc_71_n_spl_0),
    .din2(ffc_214_n_spl_10)
  );


  andX
  g_g824_p
  (
    .dout(g824_p),
    .din1(g803_n_spl_),
    .din2(g806_n_spl_)
  );


  orX
  g_g824_n
  (
    .dout(g824_n),
    .din1(g803_p_spl_),
    .din2(g806_p_spl_)
  );


  andX
  g_g825_p
  (
    .dout(g825_p),
    .din1(g745_p_spl_),
    .din2(g747_n_spl_)
  );


  orX
  g_g825_n
  (
    .dout(g825_n),
    .din1(g745_n_spl_),
    .din2(g747_p_spl_)
  );


  andX
  g_g826_p
  (
    .dout(g826_p),
    .din1(g748_n_spl_),
    .din2(g825_n)
  );


  orX
  g_g826_n
  (
    .dout(g826_n),
    .din1(g748_p_spl_),
    .din2(g825_p)
  );


  andX
  g_g827_p
  (
    .dout(g827_p),
    .din1(g824_n_spl_),
    .din2(g826_p_spl_)
  );


  orX
  g_g827_n
  (
    .dout(g827_n),
    .din1(g824_p_spl_),
    .din2(g826_n_spl_)
  );


  andX
  g_g828_p
  (
    .dout(g828_p),
    .din1(g824_p_spl_),
    .din2(g826_n_spl_)
  );


  orX
  g_g828_n
  (
    .dout(g828_n),
    .din1(g824_n_spl_),
    .din2(g826_p_spl_)
  );


  andX
  g_g829_p
  (
    .dout(g829_p),
    .din1(g827_n_spl_),
    .din2(g828_n)
  );


  orX
  g_g829_n
  (
    .dout(g829_n),
    .din1(g827_p_spl_),
    .din2(g828_p)
  );


  andX
  g_g830_p
  (
    .dout(g830_p),
    .din1(g823_n_spl_),
    .din2(g829_p_spl_)
  );


  orX
  g_g830_n
  (
    .dout(g830_n),
    .din1(g823_p_spl_),
    .din2(g829_n_spl_)
  );


  andX
  g_g831_p
  (
    .dout(g831_p),
    .din1(g823_p_spl_),
    .din2(g829_n_spl_)
  );


  orX
  g_g831_n
  (
    .dout(g831_n),
    .din1(g823_n_spl_),
    .din2(g829_p_spl_)
  );


  andX
  g_g832_p
  (
    .dout(g832_p),
    .din1(g830_n_spl_),
    .din2(g831_n)
  );


  orX
  g_g832_n
  (
    .dout(g832_n),
    .din1(g830_p_spl_),
    .din2(g831_p)
  );


  andX
  g_g833_p
  (
    .dout(g833_p),
    .din1(g822_n_spl_),
    .din2(g832_p_spl_)
  );


  orX
  g_g833_n
  (
    .dout(g833_n),
    .din1(g822_p_spl_),
    .din2(g832_n_spl_)
  );


  andX
  g_g834_p
  (
    .dout(g834_p),
    .din1(g822_p_spl_),
    .din2(g832_n_spl_)
  );


  orX
  g_g834_n
  (
    .dout(g834_n),
    .din1(g822_n_spl_),
    .din2(g832_p_spl_)
  );


  andX
  g_g835_p
  (
    .dout(g835_p),
    .din1(g833_n_spl_),
    .din2(g834_n)
  );


  orX
  g_g835_n
  (
    .dout(g835_n),
    .din1(g833_p_spl_),
    .din2(g834_p)
  );


  andX
  g_g836_p
  (
    .dout(g836_p),
    .din1(g821_n_spl_),
    .din2(g835_p_spl_)
  );


  orX
  g_g836_n
  (
    .dout(g836_n),
    .din1(g821_p_spl_),
    .din2(g835_n_spl_)
  );


  andX
  g_g837_p
  (
    .dout(g837_p),
    .din1(g821_p_spl_),
    .din2(g835_n_spl_)
  );


  orX
  g_g837_n
  (
    .dout(g837_n),
    .din1(g821_n_spl_),
    .din2(g835_p_spl_)
  );


  andX
  g_g838_p
  (
    .dout(g838_p),
    .din1(g836_n_spl_),
    .din2(g837_n)
  );


  orX
  g_g838_n
  (
    .dout(g838_n),
    .din1(g836_p_spl_),
    .din2(g837_p)
  );


  andX
  g_g839_p
  (
    .dout(g839_p),
    .din1(g820_n_spl_),
    .din2(g838_p_spl_)
  );


  orX
  g_g839_n
  (
    .dout(g839_n),
    .din1(g820_p_spl_),
    .din2(g838_n_spl_)
  );


  andX
  g_g840_p
  (
    .dout(g840_p),
    .din1(g674_n_spl_),
    .din2(g701_p_spl_)
  );


  andX
  g_g841_p
  (
    .dout(g841_p),
    .din1(g668_n_spl_),
    .din2(g671_n)
  );


  orX
  g_g841_n
  (
    .dout(g841_n),
    .din1(g668_p_spl_),
    .din2(g671_p_spl_)
  );


  andX
  g_g842_p
  (
    .dout(g842_p),
    .din1(ffc_15_p_spl_000),
    .din2(ffc_133_p_spl_00)
  );


  orX
  g_g842_n
  (
    .dout(g842_n),
    .din1(ffc_15_n_spl_000),
    .din2(ffc_133_n_spl_00)
  );


  andX
  g_g843_p
  (
    .dout(g843_p),
    .din1(ffc_310_p_spl_),
    .din2(g665_n_spl_)
  );


  orX
  g_g843_n
  (
    .dout(g843_n),
    .din1(ffc_310_n_spl_),
    .din2(g665_p_spl_)
  );


  andX
  g_g844_p
  (
    .dout(g844_p),
    .din1(ffc_118_p_spl_00),
    .din2(ffc_287_p_spl_001)
  );


  orX
  g_g844_n
  (
    .dout(g844_n),
    .din1(ffc_118_n_spl_00),
    .din2(ffc_287_n_spl_001)
  );


  andX
  g_g845_p
  (
    .dout(g845_p),
    .din1(ffc_296_p_spl_),
    .din2(ffc_297_n)
  );


  orX
  g_g845_n
  (
    .dout(g845_n),
    .din1(ffc_296_n_spl_),
    .din2(ffc_297_p)
  );


  andX
  g_g846_p
  (
    .dout(g846_p),
    .din1(g844_n_spl_),
    .din2(g845_p_spl_)
  );


  orX
  g_g846_n
  (
    .dout(g846_n),
    .din1(g844_p_spl_),
    .din2(g845_n_spl_)
  );


  andX
  g_g847_p
  (
    .dout(g847_p),
    .din1(g844_p_spl_),
    .din2(g845_n_spl_)
  );


  orX
  g_g847_n
  (
    .dout(g847_n),
    .din1(g844_n_spl_),
    .din2(g845_p_spl_)
  );


  andX
  g_g848_p
  (
    .dout(g848_p),
    .din1(g846_n_spl_),
    .din2(g847_n)
  );


  orX
  g_g848_n
  (
    .dout(g848_n),
    .din1(g846_p_spl_),
    .din2(g847_p)
  );


  andX
  g_g849_p
  (
    .dout(g849_p),
    .din1(g843_n_spl_),
    .din2(g848_p_spl_)
  );


  orX
  g_g849_n
  (
    .dout(g849_n),
    .din1(g843_p_spl_),
    .din2(g848_n_spl_)
  );


  andX
  g_g850_p
  (
    .dout(g850_p),
    .din1(g843_p_spl_),
    .din2(g848_n_spl_)
  );


  orX
  g_g850_n
  (
    .dout(g850_n),
    .din1(g843_n_spl_),
    .din2(g848_p_spl_)
  );


  andX
  g_g851_p
  (
    .dout(g851_p),
    .din1(g849_n_spl_),
    .din2(g850_n)
  );


  orX
  g_g851_n
  (
    .dout(g851_n),
    .din1(g849_p_spl_),
    .din2(g850_p)
  );


  andX
  g_g852_p
  (
    .dout(g852_p),
    .din1(g842_n_spl_),
    .din2(g851_p_spl_)
  );


  orX
  g_g852_n
  (
    .dout(g852_n),
    .din1(g842_p_spl_),
    .din2(g851_n_spl_)
  );


  andX
  g_g853_p
  (
    .dout(g853_p),
    .din1(g842_p_spl_),
    .din2(g851_n_spl_)
  );


  orX
  g_g853_n
  (
    .dout(g853_n),
    .din1(g842_n_spl_),
    .din2(g851_p_spl_)
  );


  andX
  g_g854_p
  (
    .dout(g854_p),
    .din1(g852_n_spl_),
    .din2(g853_n)
  );


  orX
  g_g854_n
  (
    .dout(g854_n),
    .din1(g852_p_spl_),
    .din2(g853_p)
  );


  andX
  g_g855_p
  (
    .dout(g855_p),
    .din1(g841_n_spl_),
    .din2(g854_p_spl_)
  );


  orX
  g_g855_n
  (
    .dout(g855_n),
    .din1(g841_p_spl_),
    .din2(g854_n_spl_)
  );


  andX
  g_g856_p
  (
    .dout(g856_p),
    .din1(g841_p_spl_),
    .din2(g854_n_spl_)
  );


  orX
  g_g856_n
  (
    .dout(g856_n),
    .din1(g841_n_spl_),
    .din2(g854_p_spl_)
  );


  andX
  g_g857_p
  (
    .dout(g857_p),
    .din1(g855_n_spl_),
    .din2(g856_n)
  );


  orX
  g_g857_n
  (
    .dout(g857_n),
    .din1(g855_p_spl_),
    .din2(g856_p)
  );


  andX
  g_g858_p
  (
    .dout(g858_p),
    .din1(ffc_341_p_spl_),
    .din2(g702_n)
  );


  orX
  g_g858_n
  (
    .dout(g858_n),
    .din1(ffc_341_n_spl_),
    .din2(g702_p_spl_)
  );


  andX
  g_g859_p
  (
    .dout(g859_p),
    .din1(ffc_339_n_spl_),
    .din2(ffc_355_p_spl_)
  );


  orX
  g_g859_n
  (
    .dout(g859_n),
    .din1(ffc_339_p_spl_),
    .din2(ffc_355_n_spl_)
  );


  andX
  g_g860_p
  (
    .dout(g860_p),
    .din1(ffc_339_p_spl_),
    .din2(ffc_355_n_spl_)
  );


  orX
  g_g860_n
  (
    .dout(g860_n),
    .din1(ffc_339_n_spl_),
    .din2(ffc_355_p_spl_)
  );


  andX
  g_g861_p
  (
    .dout(g861_p),
    .din1(g859_n_spl_),
    .din2(g860_n)
  );


  orX
  g_g861_n
  (
    .dout(g861_n),
    .din1(g859_p_spl_),
    .din2(g860_p)
  );


  andX
  g_g862_p
  (
    .dout(g862_p),
    .din1(g858_n_spl_),
    .din2(g861_p_spl_)
  );


  orX
  g_g862_n
  (
    .dout(g862_n),
    .din1(g858_p_spl_),
    .din2(g861_n_spl_)
  );


  andX
  g_g863_p
  (
    .dout(g863_p),
    .din1(g858_p_spl_),
    .din2(g861_n_spl_)
  );


  orX
  g_g863_n
  (
    .dout(g863_n),
    .din1(g858_n_spl_),
    .din2(g861_p_spl_)
  );


  andX
  g_g864_p
  (
    .dout(g864_p),
    .din1(g862_n_spl_),
    .din2(g863_n)
  );


  orX
  g_g864_n
  (
    .dout(g864_n),
    .din1(g862_p_spl_),
    .din2(g863_p)
  );


  andX
  g_g865_p
  (
    .dout(g865_p),
    .din1(g703_n),
    .din2(g857_p_spl_)
  );


  orX
  g_g865_n
  (
    .dout(g865_n),
    .din1(g703_p_spl_),
    .din2(g857_n)
  );


  andX
  g_g866_p
  (
    .dout(g866_p),
    .din1(g704_n),
    .din2(g864_p_spl_)
  );


  orX
  g_g866_n
  (
    .dout(g866_n),
    .din1(g704_p_spl_),
    .din2(g864_n)
  );


  orX
  g_g867_n
  (
    .dout(g867_n),
    .din1(g699_p),
    .din2(g840_p_spl_)
  );


  andX
  g_g868_p
  (
    .dout(g868_p),
    .din1(g693_n_spl_),
    .din2(g696_n_spl_)
  );


  orX
  g_g868_n
  (
    .dout(g868_n),
    .din1(g693_p_spl_),
    .din2(g696_p_spl_)
  );


  andX
  g_g869_p
  (
    .dout(g869_p),
    .din1(ffc_29_p_spl_10),
    .din2(ffc_67_p_spl_)
  );


  orX
  g_g869_n
  (
    .dout(g869_n),
    .din1(ffc_29_n_spl_10),
    .din2(ffc_67_n_spl_)
  );


  andX
  g_g870_p
  (
    .dout(g870_p),
    .din1(g687_n_spl_),
    .din2(g690_n_spl_)
  );


  orX
  g_g870_n
  (
    .dout(g870_n),
    .din1(g687_p_spl_),
    .din2(g690_p_spl_)
  );


  andX
  g_g871_p
  (
    .dout(g871_p),
    .din1(ffc_25_p_spl_10),
    .din2(ffc_68_p_spl_0)
  );


  orX
  g_g871_n
  (
    .dout(g871_n),
    .din1(ffc_25_n_spl_10),
    .din2(ffc_68_n_spl_0)
  );


  andX
  g_g872_p
  (
    .dout(g872_p),
    .din1(g681_n_spl_),
    .din2(g684_n_spl_)
  );


  orX
  g_g872_n
  (
    .dout(g872_n),
    .din1(g681_p_spl_),
    .din2(g684_p_spl_)
  );


  andX
  g_g873_p
  (
    .dout(g873_p),
    .din1(g795_p_spl_),
    .din2(g797_n_spl_)
  );


  orX
  g_g873_n
  (
    .dout(g873_n),
    .din1(g795_n_spl_),
    .din2(g797_p_spl_)
  );


  andX
  g_g874_p
  (
    .dout(g874_p),
    .din1(g798_n_spl_),
    .din2(g873_n)
  );


  orX
  g_g874_n
  (
    .dout(g874_n),
    .din1(g798_p_spl_),
    .din2(g873_p)
  );


  andX
  g_g875_p
  (
    .dout(g875_p),
    .din1(g872_n_spl_),
    .din2(g874_p_spl_)
  );


  orX
  g_g875_n
  (
    .dout(g875_n),
    .din1(g872_p_spl_),
    .din2(g874_n_spl_)
  );


  andX
  g_g876_p
  (
    .dout(g876_p),
    .din1(g872_p_spl_),
    .din2(g874_n_spl_)
  );


  orX
  g_g876_n
  (
    .dout(g876_n),
    .din1(g872_n_spl_),
    .din2(g874_p_spl_)
  );


  andX
  g_g877_p
  (
    .dout(g877_p),
    .din1(g875_n_spl_),
    .din2(g876_n)
  );


  orX
  g_g877_n
  (
    .dout(g877_n),
    .din1(g875_p_spl_),
    .din2(g876_p)
  );


  andX
  g_g878_p
  (
    .dout(g878_p),
    .din1(g871_n_spl_),
    .din2(g877_p_spl_)
  );


  orX
  g_g878_n
  (
    .dout(g878_n),
    .din1(g871_p_spl_),
    .din2(g877_n_spl_)
  );


  andX
  g_g879_p
  (
    .dout(g879_p),
    .din1(g871_p_spl_),
    .din2(g877_n_spl_)
  );


  orX
  g_g879_n
  (
    .dout(g879_n),
    .din1(g871_n_spl_),
    .din2(g877_p_spl_)
  );


  andX
  g_g880_p
  (
    .dout(g880_p),
    .din1(g878_n_spl_),
    .din2(g879_n)
  );


  orX
  g_g880_n
  (
    .dout(g880_n),
    .din1(g878_p_spl_),
    .din2(g879_p)
  );


  andX
  g_g881_p
  (
    .dout(g881_p),
    .din1(g870_n_spl_),
    .din2(g880_p_spl_)
  );


  orX
  g_g881_n
  (
    .dout(g881_n),
    .din1(g870_p_spl_),
    .din2(g880_n_spl_)
  );


  andX
  g_g882_p
  (
    .dout(g882_p),
    .din1(g870_p_spl_),
    .din2(g880_n_spl_)
  );


  orX
  g_g882_n
  (
    .dout(g882_n),
    .din1(g870_n_spl_),
    .din2(g880_p_spl_)
  );


  andX
  g_g883_p
  (
    .dout(g883_p),
    .din1(g881_n_spl_),
    .din2(g882_n)
  );


  orX
  g_g883_n
  (
    .dout(g883_n),
    .din1(g881_p_spl_),
    .din2(g882_p)
  );


  andX
  g_g884_p
  (
    .dout(g884_p),
    .din1(g869_n_spl_),
    .din2(g883_p_spl_)
  );


  orX
  g_g884_n
  (
    .dout(g884_n),
    .din1(g869_p_spl_),
    .din2(g883_n_spl_)
  );


  andX
  g_g885_p
  (
    .dout(g885_p),
    .din1(g869_p_spl_),
    .din2(g883_n_spl_)
  );


  orX
  g_g885_n
  (
    .dout(g885_n),
    .din1(g869_n_spl_),
    .din2(g883_p_spl_)
  );


  andX
  g_g886_p
  (
    .dout(g886_p),
    .din1(g884_n_spl_),
    .din2(g885_n)
  );


  orX
  g_g886_n
  (
    .dout(g886_n),
    .din1(g884_p_spl_),
    .din2(g885_p)
  );


  andX
  g_g887_p
  (
    .dout(g887_p),
    .din1(g868_n_spl_),
    .din2(g886_p_spl_)
  );


  orX
  g_g887_n
  (
    .dout(g887_n),
    .din1(g868_p),
    .din2(g886_n)
  );


  orX
  g_g888_n
  (
    .dout(g888_n),
    .din1(g868_n_spl_),
    .din2(g886_p_spl_)
  );


  andX
  g_g889_p
  (
    .dout(g889_p),
    .din1(g887_n),
    .din2(g888_n)
  );


  andX
  g_g890_p
  (
    .dout(g890_p),
    .din1(ffc_10_p_spl_000),
    .din2(ffc_207_p_spl_0)
  );


  orX
  g_g890_n
  (
    .dout(g890_n),
    .din1(ffc_10_n_spl_000),
    .din2(ffc_207_n_spl_0)
  );


  andX
  g_g891_p
  (
    .dout(g891_p),
    .din1(g862_n_spl_),
    .din2(g866_n)
  );


  orX
  g_g891_n
  (
    .dout(g891_n),
    .din1(g862_p_spl_),
    .din2(g866_p_spl_)
  );


  andX
  g_g892_p
  (
    .dout(g892_p),
    .din1(ffc_9_p_spl_000),
    .din2(ffc_195_p_spl_00)
  );


  orX
  g_g892_n
  (
    .dout(g892_n),
    .din1(ffc_9_n_spl_000),
    .din2(ffc_195_n_spl_0)
  );


  andX
  g_g893_p
  (
    .dout(g893_p),
    .din1(ffc_324_p),
    .din2(g859_n_spl_)
  );


  orX
  g_g893_n
  (
    .dout(g893_n),
    .din1(ffc_324_n),
    .din2(g859_p_spl_)
  );


  andX
  g_g894_p
  (
    .dout(g894_p),
    .din1(ffc_326_n_spl_),
    .din2(ffc_343_p_spl_)
  );


  orX
  g_g894_n
  (
    .dout(g894_n),
    .din1(ffc_326_p_spl_),
    .din2(ffc_343_n_spl_)
  );


  andX
  g_g895_p
  (
    .dout(g895_p),
    .din1(ffc_326_p_spl_),
    .din2(ffc_343_n_spl_)
  );


  orX
  g_g895_n
  (
    .dout(g895_n),
    .din1(ffc_326_n_spl_),
    .din2(ffc_343_p_spl_)
  );


  andX
  g_g896_p
  (
    .dout(g896_p),
    .din1(g894_n_spl_),
    .din2(g895_n)
  );


  orX
  g_g896_n
  (
    .dout(g896_n),
    .din1(g894_p_spl_),
    .din2(g895_p)
  );


  andX
  g_g897_p
  (
    .dout(g897_p),
    .din1(g893_n_spl_),
    .din2(g896_p_spl_)
  );


  orX
  g_g897_n
  (
    .dout(g897_n),
    .din1(g893_p_spl_),
    .din2(g896_n_spl_)
  );


  andX
  g_g898_p
  (
    .dout(g898_p),
    .din1(g893_p_spl_),
    .din2(g896_n_spl_)
  );


  orX
  g_g898_n
  (
    .dout(g898_n),
    .din1(g893_n_spl_),
    .din2(g896_p_spl_)
  );


  andX
  g_g899_p
  (
    .dout(g899_p),
    .din1(g897_n_spl_),
    .din2(g898_n)
  );


  orX
  g_g899_n
  (
    .dout(g899_n),
    .din1(g897_p_spl_),
    .din2(g898_p)
  );


  andX
  g_g900_p
  (
    .dout(g900_p),
    .din1(g892_n_spl_),
    .din2(g899_p_spl_)
  );


  orX
  g_g900_n
  (
    .dout(g900_n),
    .din1(g892_p_spl_),
    .din2(g899_n_spl_)
  );


  andX
  g_g901_p
  (
    .dout(g901_p),
    .din1(g892_p_spl_),
    .din2(g899_n_spl_)
  );


  orX
  g_g901_n
  (
    .dout(g901_n),
    .din1(g892_n_spl_),
    .din2(g899_p_spl_)
  );


  andX
  g_g902_p
  (
    .dout(g902_p),
    .din1(g900_n_spl_),
    .din2(g901_n)
  );


  orX
  g_g902_n
  (
    .dout(g902_n),
    .din1(g900_p_spl_),
    .din2(g901_p)
  );


  andX
  g_g903_p
  (
    .dout(g903_p),
    .din1(g891_n_spl_),
    .din2(g902_p_spl_)
  );


  orX
  g_g903_n
  (
    .dout(g903_n),
    .din1(g891_p_spl_),
    .din2(g902_n_spl_)
  );


  andX
  g_g904_p
  (
    .dout(g904_p),
    .din1(g891_p_spl_),
    .din2(g902_n_spl_)
  );


  orX
  g_g904_n
  (
    .dout(g904_n),
    .din1(g891_n_spl_),
    .din2(g902_p_spl_)
  );


  andX
  g_g905_p
  (
    .dout(g905_p),
    .din1(g903_n_spl_),
    .din2(g904_n)
  );


  orX
  g_g905_n
  (
    .dout(g905_n),
    .din1(g903_p_spl_),
    .din2(g904_p)
  );


  andX
  g_g906_p
  (
    .dout(g906_p),
    .din1(g890_n),
    .din2(g905_p_spl_)
  );


  orX
  g_g906_n
  (
    .dout(g906_n),
    .din1(g890_p_spl_),
    .din2(g905_n)
  );


  andX
  g_g907_p
  (
    .dout(g907_p),
    .din1(ffc_19_p_spl_000),
    .din2(ffc_135_p_spl_1)
  );


  orX
  g_g907_n
  (
    .dout(g907_n),
    .din1(ffc_19_n_spl_00),
    .din2(ffc_135_n_spl_1)
  );


  andX
  g_g908_p
  (
    .dout(g908_p),
    .din1(ffc_29_p_spl_10),
    .din2(ffc_69_p_spl_)
  );


  orX
  g_g908_n
  (
    .dout(g908_n),
    .din1(ffc_29_n_spl_10),
    .din2(ffc_69_n_spl_)
  );


  andX
  g_g909_p
  (
    .dout(g909_p),
    .din1(g820_p_spl_),
    .din2(g838_n_spl_)
  );


  orX
  g_g909_n
  (
    .dout(g909_n),
    .din1(g820_n_spl_),
    .din2(g838_p_spl_)
  );


  andX
  g_g910_p
  (
    .dout(g910_p),
    .din1(g839_n_spl_),
    .din2(g909_n)
  );


  orX
  g_g910_n
  (
    .dout(g910_n),
    .din1(g839_p),
    .din2(g909_p)
  );


  orX
  g_g911_n
  (
    .dout(g911_n),
    .din1(g908_p),
    .din2(g910_n)
  );


  andX
  g_g912_p
  (
    .dout(g912_p),
    .din1(ffc_25_p_spl_10),
    .din2(ffc_72_p_spl_1)
  );


  orX
  g_g912_n
  (
    .dout(g912_n),
    .din1(ffc_25_n_spl_10),
    .din2(ffc_72_n_spl_)
  );


  andX
  g_g913_p
  (
    .dout(g913_p),
    .din1(g770_p_spl_),
    .din2(g788_n_spl_)
  );


  orX
  g_g913_n
  (
    .dout(g913_n),
    .din1(g770_n_spl_),
    .din2(g788_p_spl_)
  );


  andX
  g_g914_p
  (
    .dout(g914_p),
    .din1(g789_n_spl_),
    .din2(g913_n)
  );


  orX
  g_g914_n
  (
    .dout(g914_n),
    .din1(g789_p),
    .din2(g913_p)
  );


  orX
  g_g915_n
  (
    .dout(g915_n),
    .din1(g912_p),
    .din2(g914_n)
  );


  andX
  g_g916_p
  (
    .dout(g916_p),
    .din1(ffc_75_p_spl_1),
    .din2(ffc_214_p_spl_10)
  );


  orX
  g_g916_n
  (
    .dout(g916_n),
    .din1(ffc_75_n_spl_),
    .din2(ffc_214_n_spl_10)
  );


  andX
  g_g917_p
  (
    .dout(g917_p),
    .din1(g729_p_spl_),
    .din2(g738_n_spl_)
  );


  orX
  g_g917_n
  (
    .dout(g917_n),
    .din1(g729_n_spl_),
    .din2(g738_p_spl_)
  );


  andX
  g_g918_p
  (
    .dout(g918_p),
    .din1(g739_n_spl_),
    .din2(g917_n)
  );


  orX
  g_g918_n
  (
    .dout(g918_n),
    .din1(g739_p),
    .din2(g917_p)
  );


  orX
  g_g919_n
  (
    .dout(g919_n),
    .din1(g916_p),
    .din2(g918_n)
  );


  andX
  g_g920_p
  (
    .dout(g920_p),
    .din1(ffc_77_p_spl_1),
    .din2(ffc_174_p_spl_1)
  );


  orX
  g_g920_n
  (
    .dout(g920_n),
    .din1(ffc_77_n_spl_),
    .din2(ffc_174_n_spl_1)
  );


  andX
  g_g921_p
  (
    .dout(g921_p),
    .din1(g733_n_spl_),
    .din2(g736_n_spl_)
  );


  orX
  g_g921_n
  (
    .dout(g921_n),
    .din1(g733_p_spl_),
    .din2(g736_p_spl_)
  );


  orX
  g_g922_n
  (
    .dout(g922_n),
    .din1(g920_p),
    .din2(g921_p)
  );


  andX
  g_g923_p
  (
    .dout(g923_p),
    .din1(g783_n_spl_),
    .din2(g786_n_spl_)
  );


  orX
  g_g923_n
  (
    .dout(g923_n),
    .din1(g783_p_spl_),
    .din2(g786_p_spl_)
  );


  andX
  g_g924_p
  (
    .dout(g924_p),
    .din1(ffc_74_p_spl_1),
    .din2(ffc_214_p_spl_11)
  );


  orX
  g_g924_n
  (
    .dout(g924_n),
    .din1(ffc_74_n_spl_),
    .din2(ffc_214_n_spl_11)
  );


  andX
  g_g925_p
  (
    .dout(g925_p),
    .din1(g777_n_spl_),
    .din2(g780_n_spl_)
  );


  orX
  g_g925_n
  (
    .dout(g925_n),
    .din1(g777_p_spl_),
    .din2(g780_p_spl_)
  );


  andX
  g_g926_p
  (
    .dout(g926_p),
    .din1(g725_p_spl_),
    .din2(g727_n_spl_)
  );


  orX
  g_g926_n
  (
    .dout(g926_n),
    .din1(g725_n_spl_),
    .din2(g727_p_spl_)
  );


  andX
  g_g927_p
  (
    .dout(g927_p),
    .din1(g728_n_spl_),
    .din2(g926_n)
  );


  orX
  g_g927_n
  (
    .dout(g927_n),
    .din1(g728_p_spl_),
    .din2(g926_p)
  );


  andX
  g_g928_p
  (
    .dout(g928_p),
    .din1(g925_n_spl_),
    .din2(g927_p_spl_)
  );


  orX
  g_g928_n
  (
    .dout(g928_n),
    .din1(g925_p_spl_),
    .din2(g927_n_spl_)
  );


  andX
  g_g929_p
  (
    .dout(g929_p),
    .din1(g925_p_spl_),
    .din2(g927_n_spl_)
  );


  orX
  g_g929_n
  (
    .dout(g929_n),
    .din1(g925_n_spl_),
    .din2(g927_p_spl_)
  );


  andX
  g_g930_p
  (
    .dout(g930_p),
    .din1(g928_n),
    .din2(g929_n)
  );


  orX
  g_g930_n
  (
    .dout(g930_n),
    .din1(g928_p_spl_),
    .din2(g929_p)
  );


  andX
  g_g931_p
  (
    .dout(g931_p),
    .din1(g924_n_spl_),
    .din2(g930_p_spl_)
  );


  orX
  g_g931_n
  (
    .dout(g931_n),
    .din1(g924_p_spl_),
    .din2(g930_n_spl_)
  );


  andX
  g_g932_p
  (
    .dout(g932_p),
    .din1(g924_p_spl_),
    .din2(g930_n_spl_)
  );


  orX
  g_g932_n
  (
    .dout(g932_n),
    .din1(g924_n_spl_),
    .din2(g930_p_spl_)
  );


  andX
  g_g933_p
  (
    .dout(g933_p),
    .din1(g931_n),
    .din2(g932_n)
  );


  orX
  g_g933_n
  (
    .dout(g933_n),
    .din1(g931_p_spl_),
    .din2(g932_p)
  );


  orX
  g_g934_n
  (
    .dout(g934_n),
    .din1(g923_p),
    .din2(g933_n)
  );


  andX
  g_g935_p
  (
    .dout(g935_p),
    .din1(g833_n_spl_),
    .din2(g836_n_spl_)
  );


  orX
  g_g935_n
  (
    .dout(g935_n),
    .din1(g833_p_spl_),
    .din2(g836_p_spl_)
  );


  andX
  g_g936_p
  (
    .dout(g936_p),
    .din1(ffc_25_p_spl_11),
    .din2(ffc_71_p_spl_1)
  );


  orX
  g_g936_n
  (
    .dout(g936_n),
    .din1(ffc_25_n_spl_11),
    .din2(ffc_71_n_spl_)
  );


  andX
  g_g937_p
  (
    .dout(g937_p),
    .din1(g827_n_spl_),
    .din2(g830_n_spl_)
  );


  orX
  g_g937_n
  (
    .dout(g937_n),
    .din1(g827_p_spl_),
    .din2(g830_p_spl_)
  );


  andX
  g_g938_p
  (
    .dout(g938_p),
    .din1(g766_p_spl_),
    .din2(g768_n_spl_)
  );


  orX
  g_g938_n
  (
    .dout(g938_n),
    .din1(g766_n_spl_),
    .din2(g768_p_spl_)
  );


  andX
  g_g939_p
  (
    .dout(g939_p),
    .din1(g769_n_spl_),
    .din2(g938_n)
  );


  orX
  g_g939_n
  (
    .dout(g939_n),
    .din1(g769_p_spl_),
    .din2(g938_p)
  );


  andX
  g_g940_p
  (
    .dout(g940_p),
    .din1(g937_n_spl_),
    .din2(g939_p_spl_)
  );


  orX
  g_g940_n
  (
    .dout(g940_n),
    .din1(g937_p_spl_),
    .din2(g939_n_spl_)
  );


  andX
  g_g941_p
  (
    .dout(g941_p),
    .din1(g937_p_spl_),
    .din2(g939_n_spl_)
  );


  orX
  g_g941_n
  (
    .dout(g941_n),
    .din1(g937_n_spl_),
    .din2(g939_p_spl_)
  );


  andX
  g_g942_p
  (
    .dout(g942_p),
    .din1(g940_n),
    .din2(g941_n)
  );


  orX
  g_g942_n
  (
    .dout(g942_n),
    .din1(g940_p_spl_),
    .din2(g941_p)
  );


  andX
  g_g943_p
  (
    .dout(g943_p),
    .din1(g936_n_spl_),
    .din2(g942_p_spl_)
  );


  orX
  g_g943_n
  (
    .dout(g943_n),
    .din1(g936_p_spl_),
    .din2(g942_n_spl_)
  );


  andX
  g_g944_p
  (
    .dout(g944_p),
    .din1(g936_p_spl_),
    .din2(g942_n_spl_)
  );


  orX
  g_g944_n
  (
    .dout(g944_n),
    .din1(g936_n_spl_),
    .din2(g942_p_spl_)
  );


  andX
  g_g945_p
  (
    .dout(g945_p),
    .din1(g943_n),
    .din2(g944_n)
  );


  orX
  g_g945_n
  (
    .dout(g945_n),
    .din1(g943_p_spl_),
    .din2(g944_p)
  );


  orX
  g_g946_n
  (
    .dout(g946_n),
    .din1(g935_p),
    .din2(g945_n)
  );


  andX
  g_g947_p
  (
    .dout(g947_p),
    .din1(g881_n_spl_),
    .din2(g884_n_spl_)
  );


  orX
  g_g947_n
  (
    .dout(g947_n),
    .din1(g881_p_spl_),
    .din2(g884_p_spl_)
  );


  andX
  g_g948_p
  (
    .dout(g948_p),
    .din1(ffc_29_p_spl_11),
    .din2(ffc_68_p_spl_)
  );


  orX
  g_g948_n
  (
    .dout(g948_n),
    .din1(ffc_29_n_spl_11),
    .din2(ffc_68_n_spl_)
  );


  andX
  g_g949_p
  (
    .dout(g949_p),
    .din1(g875_n_spl_),
    .din2(g878_n_spl_)
  );


  orX
  g_g949_n
  (
    .dout(g949_n),
    .din1(g875_p_spl_),
    .din2(g878_p_spl_)
  );


  andX
  g_g950_p
  (
    .dout(g950_p),
    .din1(g816_p_spl_),
    .din2(g818_n_spl_)
  );


  orX
  g_g950_n
  (
    .dout(g950_n),
    .din1(g816_n_spl_),
    .din2(g818_p_spl_)
  );


  andX
  g_g951_p
  (
    .dout(g951_p),
    .din1(g819_n_spl_),
    .din2(g950_n)
  );


  orX
  g_g951_n
  (
    .dout(g951_n),
    .din1(g819_p_spl_),
    .din2(g950_p)
  );


  andX
  g_g952_p
  (
    .dout(g952_p),
    .din1(g949_n_spl_),
    .din2(g951_p_spl_)
  );


  orX
  g_g952_n
  (
    .dout(g952_n),
    .din1(g949_p_spl_),
    .din2(g951_n_spl_)
  );


  andX
  g_g953_p
  (
    .dout(g953_p),
    .din1(g949_p_spl_),
    .din2(g951_n_spl_)
  );


  orX
  g_g953_n
  (
    .dout(g953_n),
    .din1(g949_n_spl_),
    .din2(g951_p_spl_)
  );


  andX
  g_g954_p
  (
    .dout(g954_p),
    .din1(g952_n),
    .din2(g953_n)
  );


  orX
  g_g954_n
  (
    .dout(g954_n),
    .din1(g952_p_spl_),
    .din2(g953_p)
  );


  andX
  g_g955_p
  (
    .dout(g955_p),
    .din1(g948_n_spl_),
    .din2(g954_p_spl_)
  );


  orX
  g_g955_n
  (
    .dout(g955_n),
    .din1(g948_p_spl_),
    .din2(g954_n_spl_)
  );


  andX
  g_g956_p
  (
    .dout(g956_p),
    .din1(g948_p_spl_),
    .din2(g954_n_spl_)
  );


  orX
  g_g956_n
  (
    .dout(g956_n),
    .din1(g948_n_spl_),
    .din2(g954_p_spl_)
  );


  andX
  g_g957_p
  (
    .dout(g957_p),
    .din1(g955_n),
    .din2(g956_n)
  );


  orX
  g_g957_n
  (
    .dout(g957_n),
    .din1(g955_p_spl_),
    .din2(g956_p)
  );


  orX
  g_g958_n
  (
    .dout(g958_n),
    .din1(g947_p),
    .din2(g957_n)
  );


  andX
  g_g959_p
  (
    .dout(g959_p),
    .din1(g867_n_spl_),
    .din2(g889_p_spl_)
  );


  andX
  g_g960_p
  (
    .dout(g960_p),
    .din1(g855_n_spl_),
    .din2(g865_n)
  );


  orX
  g_g960_n
  (
    .dout(g960_n),
    .din1(g855_p_spl_),
    .din2(g865_p_spl_)
  );


  andX
  g_g961_p
  (
    .dout(g961_p),
    .din1(ffc_17_p_spl_000),
    .din2(ffc_133_p_spl_0)
  );


  orX
  g_g961_n
  (
    .dout(g961_n),
    .din1(ffc_17_n_spl_000),
    .din2(ffc_133_n_spl_0)
  );


  andX
  g_g962_p
  (
    .dout(g962_p),
    .din1(g849_n_spl_),
    .din2(g852_n_spl_)
  );


  orX
  g_g962_n
  (
    .dout(g962_n),
    .din1(g849_p_spl_),
    .din2(g852_p_spl_)
  );


  andX
  g_g963_p
  (
    .dout(g963_p),
    .din1(ffc_15_p_spl_001),
    .din2(ffc_118_p_spl_00)
  );


  orX
  g_g963_n
  (
    .dout(g963_n),
    .din1(ffc_15_n_spl_001),
    .din2(ffc_118_n_spl_00)
  );


  andX
  g_g964_p
  (
    .dout(g964_p),
    .din1(ffc_296_p_spl_),
    .din2(g846_n_spl_)
  );


  orX
  g_g964_n
  (
    .dout(g964_n),
    .din1(ffc_296_n_spl_),
    .din2(g846_p_spl_)
  );


  andX
  g_g965_p
  (
    .dout(g965_p),
    .din1(ffc_119_p_spl_00),
    .din2(ffc_287_p_spl_001)
  );


  orX
  g_g965_n
  (
    .dout(g965_n),
    .din1(ffc_119_n_spl_00),
    .din2(ffc_287_n_spl_001)
  );


  andX
  g_g966_p
  (
    .dout(g966_p),
    .din1(ffc_298_p_spl_),
    .din2(ffc_299_n)
  );


  orX
  g_g966_n
  (
    .dout(g966_n),
    .din1(ffc_298_n_spl_),
    .din2(ffc_299_p)
  );


  andX
  g_g967_p
  (
    .dout(g967_p),
    .din1(g965_n_spl_),
    .din2(g966_p_spl_)
  );


  orX
  g_g967_n
  (
    .dout(g967_n),
    .din1(g965_p_spl_),
    .din2(g966_n_spl_)
  );


  andX
  g_g968_p
  (
    .dout(g968_p),
    .din1(g965_p_spl_),
    .din2(g966_n_spl_)
  );


  orX
  g_g968_n
  (
    .dout(g968_n),
    .din1(g965_n_spl_),
    .din2(g966_p_spl_)
  );


  andX
  g_g969_p
  (
    .dout(g969_p),
    .din1(g967_n_spl_),
    .din2(g968_n)
  );


  orX
  g_g969_n
  (
    .dout(g969_n),
    .din1(g967_p_spl_),
    .din2(g968_p)
  );


  andX
  g_g970_p
  (
    .dout(g970_p),
    .din1(g964_n_spl_),
    .din2(g969_p_spl_)
  );


  orX
  g_g970_n
  (
    .dout(g970_n),
    .din1(g964_p_spl_),
    .din2(g969_n_spl_)
  );


  andX
  g_g971_p
  (
    .dout(g971_p),
    .din1(g964_p_spl_),
    .din2(g969_n_spl_)
  );


  orX
  g_g971_n
  (
    .dout(g971_n),
    .din1(g964_n_spl_),
    .din2(g969_p_spl_)
  );


  andX
  g_g972_p
  (
    .dout(g972_p),
    .din1(g970_n_spl_),
    .din2(g971_n)
  );


  orX
  g_g972_n
  (
    .dout(g972_n),
    .din1(g970_p_spl_),
    .din2(g971_p)
  );


  andX
  g_g973_p
  (
    .dout(g973_p),
    .din1(g963_n_spl_),
    .din2(g972_p_spl_)
  );


  orX
  g_g973_n
  (
    .dout(g973_n),
    .din1(g963_p_spl_),
    .din2(g972_n_spl_)
  );


  andX
  g_g974_p
  (
    .dout(g974_p),
    .din1(g963_p_spl_),
    .din2(g972_n_spl_)
  );


  orX
  g_g974_n
  (
    .dout(g974_n),
    .din1(g963_n_spl_),
    .din2(g972_p_spl_)
  );


  andX
  g_g975_p
  (
    .dout(g975_p),
    .din1(g973_n_spl_),
    .din2(g974_n)
  );


  orX
  g_g975_n
  (
    .dout(g975_n),
    .din1(g973_p_spl_),
    .din2(g974_p)
  );


  andX
  g_g976_p
  (
    .dout(g976_p),
    .din1(g962_n_spl_),
    .din2(g975_p_spl_)
  );


  orX
  g_g976_n
  (
    .dout(g976_n),
    .din1(g962_p_spl_),
    .din2(g975_n_spl_)
  );


  andX
  g_g977_p
  (
    .dout(g977_p),
    .din1(g962_p_spl_),
    .din2(g975_n_spl_)
  );


  orX
  g_g977_n
  (
    .dout(g977_n),
    .din1(g962_n_spl_),
    .din2(g975_p_spl_)
  );


  andX
  g_g978_p
  (
    .dout(g978_p),
    .din1(g976_n_spl_),
    .din2(g977_n)
  );


  orX
  g_g978_n
  (
    .dout(g978_n),
    .din1(g976_p_spl_),
    .din2(g977_p)
  );


  andX
  g_g979_p
  (
    .dout(g979_p),
    .din1(g961_n_spl_),
    .din2(g978_p_spl_)
  );


  orX
  g_g979_n
  (
    .dout(g979_n),
    .din1(g961_p_spl_),
    .din2(g978_n_spl_)
  );


  andX
  g_g980_p
  (
    .dout(g980_p),
    .din1(g961_p_spl_),
    .din2(g978_n_spl_)
  );


  orX
  g_g980_n
  (
    .dout(g980_n),
    .din1(g961_n_spl_),
    .din2(g978_p_spl_)
  );


  andX
  g_g981_p
  (
    .dout(g981_p),
    .din1(g979_n_spl_),
    .din2(g980_n)
  );


  orX
  g_g981_n
  (
    .dout(g981_n),
    .din1(g979_p_spl_),
    .din2(g980_p)
  );


  andX
  g_g982_p
  (
    .dout(g982_p),
    .din1(g960_n_spl_),
    .din2(g981_p_spl_)
  );


  orX
  g_g982_n
  (
    .dout(g982_n),
    .din1(g960_p_spl_),
    .din2(g981_n_spl_)
  );


  andX
  g_g983_p
  (
    .dout(g983_p),
    .din1(g960_p_spl_),
    .din2(g981_n_spl_)
  );


  orX
  g_g983_n
  (
    .dout(g983_n),
    .din1(g960_n_spl_),
    .din2(g981_p_spl_)
  );


  andX
  g_g984_p
  (
    .dout(g984_p),
    .din1(g982_n_spl_),
    .din2(g983_n)
  );


  orX
  g_g984_n
  (
    .dout(g984_n),
    .din1(g982_p_spl_),
    .din2(g983_p)
  );


  andX
  g_g985_p
  (
    .dout(g985_p),
    .din1(G2_p_spl_00),
    .din2(G17_p_spl_000)
  );


  orX
  g_g985_n
  (
    .dout(g985_n),
    .din1(G2_n_spl_0),
    .din2(G17_n_spl_000)
  );


  andX
  g_g986_p
  (
    .dout(g986_p),
    .din1(G1_p_spl_0),
    .din2(G18_p_spl_000)
  );


  orX
  g_g986_n
  (
    .dout(g986_n),
    .din1(G1_n_spl_0),
    .din2(G18_n_spl_000)
  );


  andX
  g_g987_p
  (
    .dout(g987_p),
    .din1(g907_n),
    .din2(g984_p_spl_)
  );


  orX
  g_g987_n
  (
    .dout(g987_n),
    .din1(g907_p_spl_),
    .din2(g984_n)
  );


  andX
  g_g988_p
  (
    .dout(g988_p),
    .din1(ffc_11_p_spl_000),
    .din2(ffc_207_p_spl_1)
  );


  orX
  g_g988_n
  (
    .dout(g988_n),
    .din1(ffc_11_n_spl_000),
    .din2(ffc_207_n_spl_1)
  );


  andX
  g_g989_p
  (
    .dout(g989_p),
    .din1(g985_p_spl_),
    .din2(g986_p_spl_)
  );


  orX
  g_g989_n
  (
    .dout(g989_n),
    .din1(g985_n),
    .din2(g986_n)
  );


  andX
  g_g990_p
  (
    .dout(g990_p),
    .din1(g903_n_spl_),
    .din2(g906_n)
  );


  orX
  g_g990_n
  (
    .dout(g990_n),
    .din1(g903_p_spl_),
    .din2(g906_p_spl_)
  );


  andX
  g_g991_p
  (
    .dout(g991_p),
    .din1(ffc_10_p_spl_000),
    .din2(ffc_195_p_spl_00)
  );


  orX
  g_g991_n
  (
    .dout(g991_n),
    .din1(ffc_10_n_spl_000),
    .din2(ffc_195_n_spl_0)
  );


  andX
  g_g992_p
  (
    .dout(g992_p),
    .din1(g897_n_spl_),
    .din2(g900_n_spl_)
  );


  orX
  g_g992_n
  (
    .dout(g992_n),
    .din1(g897_p_spl_),
    .din2(g900_p_spl_)
  );


  andX
  g_g993_p
  (
    .dout(g993_p),
    .din1(ffc_9_p_spl_001),
    .din2(ffc_180_p_spl_00)
  );


  orX
  g_g993_n
  (
    .dout(g993_n),
    .din1(ffc_9_n_spl_001),
    .din2(ffc_180_n_spl_0)
  );


  andX
  g_g994_p
  (
    .dout(g994_p),
    .din1(ffc_312_p),
    .din2(g894_n_spl_)
  );


  orX
  g_g994_n
  (
    .dout(g994_n),
    .din1(ffc_312_n),
    .din2(g894_p_spl_)
  );


  andX
  g_g995_p
  (
    .dout(g995_p),
    .din1(ffc_327_n_spl_),
    .din2(ffc_344_p_spl_)
  );


  orX
  g_g995_n
  (
    .dout(g995_n),
    .din1(ffc_327_p_spl_),
    .din2(ffc_344_n_spl_)
  );


  andX
  g_g996_p
  (
    .dout(g996_p),
    .din1(ffc_327_p_spl_),
    .din2(ffc_344_n_spl_)
  );


  orX
  g_g996_n
  (
    .dout(g996_n),
    .din1(ffc_327_n_spl_),
    .din2(ffc_344_p_spl_)
  );


  andX
  g_g997_p
  (
    .dout(g997_p),
    .din1(g995_n_spl_),
    .din2(g996_n)
  );


  orX
  g_g997_n
  (
    .dout(g997_n),
    .din1(g995_p_spl_),
    .din2(g996_p)
  );


  andX
  g_g998_p
  (
    .dout(g998_p),
    .din1(g994_n_spl_),
    .din2(g997_p_spl_)
  );


  orX
  g_g998_n
  (
    .dout(g998_n),
    .din1(g994_p_spl_),
    .din2(g997_n_spl_)
  );


  andX
  g_g999_p
  (
    .dout(g999_p),
    .din1(g994_p_spl_),
    .din2(g997_n_spl_)
  );


  orX
  g_g999_n
  (
    .dout(g999_n),
    .din1(g994_n_spl_),
    .din2(g997_p_spl_)
  );


  andX
  g_g1000_p
  (
    .dout(g1000_p),
    .din1(g998_n_spl_),
    .din2(g999_n)
  );


  orX
  g_g1000_n
  (
    .dout(g1000_n),
    .din1(g998_p_spl_),
    .din2(g999_p)
  );


  andX
  g_g1001_p
  (
    .dout(g1001_p),
    .din1(g993_n_spl_),
    .din2(g1000_p_spl_)
  );


  orX
  g_g1001_n
  (
    .dout(g1001_n),
    .din1(g993_p_spl_),
    .din2(g1000_n_spl_)
  );


  andX
  g_g1002_p
  (
    .dout(g1002_p),
    .din1(g993_p_spl_),
    .din2(g1000_n_spl_)
  );


  orX
  g_g1002_n
  (
    .dout(g1002_n),
    .din1(g993_n_spl_),
    .din2(g1000_p_spl_)
  );


  andX
  g_g1003_p
  (
    .dout(g1003_p),
    .din1(g1001_n_spl_),
    .din2(g1002_n)
  );


  orX
  g_g1003_n
  (
    .dout(g1003_n),
    .din1(g1001_p_spl_),
    .din2(g1002_p)
  );


  andX
  g_g1004_p
  (
    .dout(g1004_p),
    .din1(g992_n_spl_),
    .din2(g1003_p_spl_)
  );


  orX
  g_g1004_n
  (
    .dout(g1004_n),
    .din1(g992_p_spl_),
    .din2(g1003_n_spl_)
  );


  andX
  g_g1005_p
  (
    .dout(g1005_p),
    .din1(g992_p_spl_),
    .din2(g1003_n_spl_)
  );


  orX
  g_g1005_n
  (
    .dout(g1005_n),
    .din1(g992_n_spl_),
    .din2(g1003_p_spl_)
  );


  andX
  g_g1006_p
  (
    .dout(g1006_p),
    .din1(g1004_n_spl_),
    .din2(g1005_n)
  );


  orX
  g_g1006_n
  (
    .dout(g1006_n),
    .din1(g1004_p_spl_),
    .din2(g1005_p)
  );


  andX
  g_g1007_p
  (
    .dout(g1007_p),
    .din1(g991_n_spl_),
    .din2(g1006_p_spl_)
  );


  orX
  g_g1007_n
  (
    .dout(g1007_n),
    .din1(g991_p_spl_),
    .din2(g1006_n_spl_)
  );


  andX
  g_g1008_p
  (
    .dout(g1008_p),
    .din1(g991_p_spl_),
    .din2(g1006_n_spl_)
  );


  orX
  g_g1008_n
  (
    .dout(g1008_n),
    .din1(g991_n_spl_),
    .din2(g1006_p_spl_)
  );


  andX
  g_g1009_p
  (
    .dout(g1009_p),
    .din1(g1007_n_spl_),
    .din2(g1008_n)
  );


  orX
  g_g1009_n
  (
    .dout(g1009_n),
    .din1(g1007_p_spl_),
    .din2(g1008_p)
  );


  andX
  g_g1010_p
  (
    .dout(g1010_p),
    .din1(g990_n_spl_),
    .din2(g1009_p_spl_)
  );


  orX
  g_g1010_n
  (
    .dout(g1010_n),
    .din1(g990_p_spl_),
    .din2(g1009_n_spl_)
  );


  andX
  g_g1011_p
  (
    .dout(g1011_p),
    .din1(g990_p_spl_),
    .din2(g1009_n_spl_)
  );


  orX
  g_g1011_n
  (
    .dout(g1011_n),
    .din1(g990_n_spl_),
    .din2(g1009_p_spl_)
  );


  andX
  g_g1012_p
  (
    .dout(g1012_p),
    .din1(g1010_n_spl_),
    .din2(g1011_n)
  );


  orX
  g_g1012_n
  (
    .dout(g1012_n),
    .din1(g1010_p_spl_),
    .din2(g1011_p)
  );


  orX
  g_g1013_n
  (
    .dout(g1013_n),
    .din1(g887_p),
    .din2(g959_p_spl_)
  );


  orX
  g_g1014_n
  (
    .dout(g1014_n),
    .din1(g947_n),
    .din2(g957_p)
  );


  andX
  g_g1015_p
  (
    .dout(g1015_p),
    .din1(g958_n_spl_),
    .din2(g1014_n)
  );


  andX
  g_g1016_p
  (
    .dout(g1016_p),
    .din1(G1_p_spl_0),
    .din2(G19_p_spl_000)
  );


  orX
  g_g1016_n
  (
    .dout(g1016_n),
    .din1(G1_n_spl_0),
    .din2(G19_n_spl_000)
  );


  andX
  g_g1017_p
  (
    .dout(g1017_p),
    .din1(ffc_257_p),
    .din2(ffc_290_n_spl_)
  );


  orX
  g_g1017_n
  (
    .dout(g1017_n),
    .din1(ffc_257_n),
    .din2(ffc_290_p_spl_)
  );


  andX
  g_g1018_p
  (
    .dout(g1018_p),
    .din1(ffc_130_p_spl_00),
    .din2(ffc_206_p_spl_)
  );


  orX
  g_g1018_n
  (
    .dout(g1018_n),
    .din1(ffc_130_n_spl_0),
    .din2(ffc_206_n_spl_)
  );


  andX
  g_g1019_p
  (
    .dout(g1019_p),
    .din1(ffc_292_p_spl_),
    .din2(ffc_293_n)
  );


  orX
  g_g1019_n
  (
    .dout(g1019_n),
    .din1(ffc_292_n_spl_),
    .din2(ffc_293_p)
  );


  andX
  g_g1020_p
  (
    .dout(g1020_p),
    .din1(g1018_n_spl_),
    .din2(g1019_p_spl_)
  );


  orX
  g_g1020_n
  (
    .dout(g1020_n),
    .din1(g1018_p_spl_),
    .din2(g1019_n_spl_)
  );


  andX
  g_g1021_p
  (
    .dout(g1021_p),
    .din1(g1018_p_spl_),
    .din2(g1019_n_spl_)
  );


  orX
  g_g1021_n
  (
    .dout(g1021_n),
    .din1(g1018_n_spl_),
    .din2(g1019_p_spl_)
  );


  andX
  g_g1022_p
  (
    .dout(g1022_p),
    .din1(g1020_n_spl_),
    .din2(g1021_n)
  );


  orX
  g_g1022_n
  (
    .dout(g1022_n),
    .din1(g1020_p_spl_),
    .din2(g1021_p)
  );


  andX
  g_g1023_p
  (
    .dout(g1023_p),
    .din1(g1017_n_spl_),
    .din2(g1022_p_spl_)
  );


  orX
  g_g1023_n
  (
    .dout(g1023_n),
    .din1(g1017_p_spl_),
    .din2(g1022_n_spl_)
  );


  andX
  g_g1024_p
  (
    .dout(g1024_p),
    .din1(ffc_129_p_spl_0),
    .din2(ffc_224_p_spl_00)
  );


  orX
  g_g1024_n
  (
    .dout(g1024_n),
    .din1(ffc_129_n_spl_0),
    .din2(ffc_224_n_spl_00)
  );


  andX
  g_g1025_p
  (
    .dout(g1025_p),
    .din1(g1017_p_spl_),
    .din2(g1022_n_spl_)
  );


  orX
  g_g1025_n
  (
    .dout(g1025_n),
    .din1(g1017_n_spl_),
    .din2(g1022_p_spl_)
  );


  andX
  g_g1026_p
  (
    .dout(g1026_p),
    .din1(g1023_n_spl_),
    .din2(g1025_n)
  );


  orX
  g_g1026_n
  (
    .dout(g1026_n),
    .din1(g1023_p_spl_),
    .din2(g1025_p)
  );


  andX
  g_g1027_p
  (
    .dout(g1027_p),
    .din1(g1024_n_spl_),
    .din2(g1026_p_spl_)
  );


  orX
  g_g1027_n
  (
    .dout(g1027_n),
    .din1(g1024_p_spl_),
    .din2(g1026_n_spl_)
  );


  andX
  g_g1028_p
  (
    .dout(g1028_p),
    .din1(g1023_n_spl_),
    .din2(g1027_n_spl_)
  );


  orX
  g_g1028_n
  (
    .dout(g1028_n),
    .din1(g1023_p_spl_),
    .din2(g1027_p_spl_)
  );


  andX
  g_g1029_p
  (
    .dout(g1029_p),
    .din1(ffc_130_p_spl_00),
    .din2(ffc_224_p_spl_00)
  );


  orX
  g_g1029_n
  (
    .dout(g1029_n),
    .din1(ffc_130_n_spl_0),
    .din2(ffc_224_n_spl_00)
  );


  andX
  g_g1030_p
  (
    .dout(g1030_p),
    .din1(ffc_131_p_spl_0),
    .din2(ffc_206_p_spl_)
  );


  orX
  g_g1030_n
  (
    .dout(g1030_n),
    .din1(ffc_131_n_spl_0),
    .din2(ffc_206_n_spl_)
  );


  andX
  g_g1031_p
  (
    .dout(g1031_p),
    .din1(ffc_292_p_spl_),
    .din2(g1020_n_spl_)
  );


  orX
  g_g1031_n
  (
    .dout(g1031_n),
    .din1(ffc_292_n_spl_),
    .din2(g1020_p_spl_)
  );


  andX
  g_g1032_p
  (
    .dout(g1032_p),
    .din1(g1030_n_spl_),
    .din2(g1031_n_spl_)
  );


  orX
  g_g1032_n
  (
    .dout(g1032_n),
    .din1(g1030_p_spl_),
    .din2(g1031_p_spl_)
  );


  andX
  g_g1033_p
  (
    .dout(g1033_p),
    .din1(g1030_p_spl_),
    .din2(g1031_p_spl_)
  );


  orX
  g_g1033_n
  (
    .dout(g1033_n),
    .din1(g1030_n_spl_),
    .din2(g1031_n_spl_)
  );


  andX
  g_g1034_p
  (
    .dout(g1034_p),
    .din1(g1032_n_spl_),
    .din2(g1033_n)
  );


  orX
  g_g1034_n
  (
    .dout(g1034_n),
    .din1(g1032_p_spl_),
    .din2(g1033_p)
  );


  andX
  g_g1035_p
  (
    .dout(g1035_p),
    .din1(g1029_n_spl_),
    .din2(g1034_p_spl_)
  );


  orX
  g_g1035_n
  (
    .dout(g1035_n),
    .din1(g1029_p_spl_),
    .din2(g1034_n_spl_)
  );


  andX
  g_g1036_p
  (
    .dout(g1036_p),
    .din1(g1029_p_spl_),
    .din2(g1034_n_spl_)
  );


  orX
  g_g1036_n
  (
    .dout(g1036_n),
    .din1(g1029_n_spl_),
    .din2(g1034_p_spl_)
  );


  andX
  g_g1037_p
  (
    .dout(g1037_p),
    .din1(g1035_n_spl_),
    .din2(g1036_n)
  );


  orX
  g_g1037_n
  (
    .dout(g1037_n),
    .din1(g1035_p_spl_),
    .din2(g1036_p)
  );


  andX
  g_g1038_p
  (
    .dout(g1038_p),
    .din1(g1028_n_spl_),
    .din2(g1037_p_spl_)
  );


  orX
  g_g1038_n
  (
    .dout(g1038_n),
    .din1(g1028_p_spl_),
    .din2(g1037_n_spl_)
  );


  andX
  g_g1039_p
  (
    .dout(g1039_p),
    .din1(ffc_129_p_spl_0),
    .din2(ffc_287_p_spl_010)
  );


  orX
  g_g1039_n
  (
    .dout(g1039_n),
    .din1(ffc_129_n_spl_0),
    .din2(ffc_287_n_spl_010)
  );


  andX
  g_g1040_p
  (
    .dout(g1040_p),
    .din1(g1028_p_spl_),
    .din2(g1037_n_spl_)
  );


  orX
  g_g1040_n
  (
    .dout(g1040_n),
    .din1(g1028_n_spl_),
    .din2(g1037_p_spl_)
  );


  andX
  g_g1041_p
  (
    .dout(g1041_p),
    .din1(g1038_n_spl_),
    .din2(g1040_n)
  );


  orX
  g_g1041_n
  (
    .dout(g1041_n),
    .din1(g1038_p_spl_),
    .din2(g1040_p)
  );


  andX
  g_g1042_p
  (
    .dout(g1042_p),
    .din1(g1039_n_spl_),
    .din2(g1041_p_spl_)
  );


  orX
  g_g1042_n
  (
    .dout(g1042_n),
    .din1(g1039_p_spl_),
    .din2(g1041_n_spl_)
  );


  andX
  g_g1043_p
  (
    .dout(g1043_p),
    .din1(g1038_n_spl_),
    .din2(g1042_n_spl_)
  );


  orX
  g_g1043_n
  (
    .dout(g1043_n),
    .din1(g1038_p_spl_),
    .din2(g1042_p_spl_)
  );


  andX
  g_g1044_p
  (
    .dout(g1044_p),
    .din1(ffc_130_p_spl_0),
    .din2(ffc_287_p_spl_010)
  );


  orX
  g_g1044_n
  (
    .dout(g1044_n),
    .din1(ffc_130_n_spl_),
    .din2(ffc_287_n_spl_010)
  );


  andX
  g_g1045_p
  (
    .dout(g1045_p),
    .din1(ffc_131_p_spl_0),
    .din2(ffc_224_p_spl_0)
  );


  orX
  g_g1045_n
  (
    .dout(g1045_n),
    .din1(ffc_131_n_spl_0),
    .din2(ffc_224_n_spl_0)
  );


  andX
  g_g1046_p
  (
    .dout(g1046_p),
    .din1(g1032_n_spl_),
    .din2(g1035_n_spl_)
  );


  orX
  g_g1046_n
  (
    .dout(g1046_n),
    .din1(g1032_p_spl_),
    .din2(g1035_p_spl_)
  );


  andX
  g_g1047_p
  (
    .dout(g1047_p),
    .din1(g1045_n_spl_),
    .din2(g1046_n_spl_)
  );


  orX
  g_g1047_n
  (
    .dout(g1047_n),
    .din1(g1045_p_spl_),
    .din2(g1046_p_spl_)
  );


  andX
  g_g1048_p
  (
    .dout(g1048_p),
    .din1(g1045_p_spl_),
    .din2(g1046_p_spl_)
  );


  orX
  g_g1048_n
  (
    .dout(g1048_n),
    .din1(g1045_n_spl_),
    .din2(g1046_n_spl_)
  );


  andX
  g_g1049_p
  (
    .dout(g1049_p),
    .din1(g1047_n_spl_),
    .din2(g1048_n)
  );


  orX
  g_g1049_n
  (
    .dout(g1049_n),
    .din1(g1047_p_spl_),
    .din2(g1048_p)
  );


  andX
  g_g1050_p
  (
    .dout(g1050_p),
    .din1(g1044_n_spl_),
    .din2(g1049_p_spl_)
  );


  orX
  g_g1050_n
  (
    .dout(g1050_n),
    .din1(g1044_p_spl_),
    .din2(g1049_n_spl_)
  );


  andX
  g_g1051_p
  (
    .dout(g1051_p),
    .din1(g1044_p_spl_),
    .din2(g1049_n_spl_)
  );


  orX
  g_g1051_n
  (
    .dout(g1051_n),
    .din1(g1044_n_spl_),
    .din2(g1049_p_spl_)
  );


  andX
  g_g1052_p
  (
    .dout(g1052_p),
    .din1(g1050_n_spl_),
    .din2(g1051_n)
  );


  orX
  g_g1052_n
  (
    .dout(g1052_n),
    .din1(g1050_p_spl_),
    .din2(g1051_p)
  );


  andX
  g_g1053_p
  (
    .dout(g1053_p),
    .din1(g1043_n_spl_),
    .din2(g1052_p_spl_)
  );


  orX
  g_g1053_n
  (
    .dout(g1053_n),
    .din1(g1043_p_spl_),
    .din2(g1052_n_spl_)
  );


  andX
  g_g1054_p
  (
    .dout(g1054_p),
    .din1(ffc_258_p),
    .din2(ffc_288_n_spl_)
  );


  orX
  g_g1054_n
  (
    .dout(g1054_n),
    .din1(ffc_258_n),
    .din2(ffc_288_p_spl_)
  );


  andX
  g_g1055_p
  (
    .dout(g1055_p),
    .din1(ffc_127_p_spl_00),
    .din2(ffc_224_p_spl_1)
  );


  orX
  g_g1055_n
  (
    .dout(g1055_n),
    .din1(ffc_127_n_spl_0),
    .din2(ffc_224_n_spl_1)
  );


  andX
  g_g1056_p
  (
    .dout(g1056_p),
    .din1(ffc_294_p_spl_),
    .din2(ffc_295_n)
  );


  orX
  g_g1056_n
  (
    .dout(g1056_n),
    .din1(ffc_294_n_spl_),
    .din2(ffc_295_p)
  );


  andX
  g_g1057_p
  (
    .dout(g1057_p),
    .din1(g1055_n_spl_),
    .din2(g1056_p_spl_)
  );


  orX
  g_g1057_n
  (
    .dout(g1057_n),
    .din1(g1055_p_spl_),
    .din2(g1056_n_spl_)
  );


  andX
  g_g1058_p
  (
    .dout(g1058_p),
    .din1(g1055_p_spl_),
    .din2(g1056_n_spl_)
  );


  orX
  g_g1058_n
  (
    .dout(g1058_n),
    .din1(g1055_n_spl_),
    .din2(g1056_p_spl_)
  );


  andX
  g_g1059_p
  (
    .dout(g1059_p),
    .din1(g1057_n_spl_),
    .din2(g1058_n)
  );


  orX
  g_g1059_n
  (
    .dout(g1059_n),
    .din1(g1057_p_spl_),
    .din2(g1058_p)
  );


  andX
  g_g1060_p
  (
    .dout(g1060_p),
    .din1(g1054_n_spl_),
    .din2(g1059_p_spl_)
  );


  orX
  g_g1060_n
  (
    .dout(g1060_n),
    .din1(g1054_p_spl_),
    .din2(g1059_n_spl_)
  );


  andX
  g_g1061_p
  (
    .dout(g1061_p),
    .din1(ffc_126_p_spl_0),
    .din2(ffc_287_p_spl_011)
  );


  orX
  g_g1061_n
  (
    .dout(g1061_n),
    .din1(ffc_126_n_spl_0),
    .din2(ffc_287_n_spl_011)
  );


  andX
  g_g1062_p
  (
    .dout(g1062_p),
    .din1(g1054_p_spl_),
    .din2(g1059_n_spl_)
  );


  orX
  g_g1062_n
  (
    .dout(g1062_n),
    .din1(g1054_n_spl_),
    .din2(g1059_p_spl_)
  );


  andX
  g_g1063_p
  (
    .dout(g1063_p),
    .din1(g1060_n_spl_),
    .din2(g1062_n)
  );


  orX
  g_g1063_n
  (
    .dout(g1063_n),
    .din1(g1060_p_spl_),
    .din2(g1062_p)
  );


  andX
  g_g1064_p
  (
    .dout(g1064_p),
    .din1(g1061_n_spl_),
    .din2(g1063_p_spl_)
  );


  orX
  g_g1064_n
  (
    .dout(g1064_n),
    .din1(g1061_p_spl_),
    .din2(g1063_n_spl_)
  );


  andX
  g_g1065_p
  (
    .dout(g1065_p),
    .din1(g1060_n_spl_),
    .din2(g1064_n_spl_)
  );


  orX
  g_g1065_n
  (
    .dout(g1065_n),
    .din1(g1060_p_spl_),
    .din2(g1064_p_spl_)
  );


  andX
  g_g1066_p
  (
    .dout(g1066_p),
    .din1(ffc_127_p_spl_00),
    .din2(ffc_287_p_spl_011)
  );


  orX
  g_g1066_n
  (
    .dout(g1066_n),
    .din1(ffc_127_n_spl_0),
    .din2(ffc_287_n_spl_011)
  );


  andX
  g_g1067_p
  (
    .dout(g1067_p),
    .din1(ffc_294_p_spl_),
    .din2(g1057_n_spl_)
  );


  orX
  g_g1067_n
  (
    .dout(g1067_n),
    .din1(ffc_294_n_spl_),
    .din2(g1057_p_spl_)
  );


  andX
  g_g1068_p
  (
    .dout(g1068_p),
    .din1(ffc_128_p_spl_0),
    .din2(ffc_224_p_spl_1)
  );


  orX
  g_g1068_n
  (
    .dout(g1068_n),
    .din1(ffc_128_n_spl_0),
    .din2(ffc_224_n_spl_1)
  );


  andX
  g_g1069_p
  (
    .dout(g1069_p),
    .din1(ffc_226_p),
    .din2(ffc_256_n)
  );


  orX
  g_g1069_n
  (
    .dout(g1069_n),
    .din1(ffc_226_n),
    .din2(ffc_256_p)
  );


  andX
  g_g1070_p
  (
    .dout(g1070_p),
    .din1(ffc_290_n_spl_),
    .din2(ffc_291_n)
  );


  orX
  g_g1070_n
  (
    .dout(g1070_n),
    .din1(ffc_290_p_spl_),
    .din2(ffc_291_p)
  );


  andX
  g_g1071_p
  (
    .dout(g1071_p),
    .din1(g1069_n_spl_),
    .din2(g1070_p_spl_)
  );


  orX
  g_g1071_n
  (
    .dout(g1071_n),
    .din1(g1069_p_spl_),
    .din2(g1070_n_spl_)
  );


  andX
  g_g1072_p
  (
    .dout(g1072_p),
    .din1(g1069_p_spl_),
    .din2(g1070_n_spl_)
  );


  orX
  g_g1072_n
  (
    .dout(g1072_n),
    .din1(g1069_n_spl_),
    .din2(g1070_p_spl_)
  );


  andX
  g_g1073_p
  (
    .dout(g1073_p),
    .din1(g1071_n_spl_),
    .din2(g1072_n)
  );


  orX
  g_g1073_n
  (
    .dout(g1073_n),
    .din1(g1071_p_spl_),
    .din2(g1072_p)
  );


  andX
  g_g1074_p
  (
    .dout(g1074_p),
    .din1(g1068_n_spl_),
    .din2(g1073_p_spl_)
  );


  orX
  g_g1074_n
  (
    .dout(g1074_n),
    .din1(g1068_p_spl_),
    .din2(g1073_n_spl_)
  );


  andX
  g_g1075_p
  (
    .dout(g1075_p),
    .din1(g1068_p_spl_),
    .din2(g1073_n_spl_)
  );


  orX
  g_g1075_n
  (
    .dout(g1075_n),
    .din1(g1068_n_spl_),
    .din2(g1073_p_spl_)
  );


  andX
  g_g1076_p
  (
    .dout(g1076_p),
    .din1(g1074_n_spl_),
    .din2(g1075_n)
  );


  orX
  g_g1076_n
  (
    .dout(g1076_n),
    .din1(g1074_p_spl_),
    .din2(g1075_p)
  );


  andX
  g_g1077_p
  (
    .dout(g1077_p),
    .din1(g1067_n_spl_),
    .din2(g1076_p_spl_)
  );


  orX
  g_g1077_n
  (
    .dout(g1077_n),
    .din1(g1067_p_spl_),
    .din2(g1076_n_spl_)
  );


  andX
  g_g1078_p
  (
    .dout(g1078_p),
    .din1(g1067_p_spl_),
    .din2(g1076_n_spl_)
  );


  orX
  g_g1078_n
  (
    .dout(g1078_n),
    .din1(g1067_n_spl_),
    .din2(g1076_p_spl_)
  );


  andX
  g_g1079_p
  (
    .dout(g1079_p),
    .din1(g1077_n_spl_),
    .din2(g1078_n)
  );


  orX
  g_g1079_n
  (
    .dout(g1079_n),
    .din1(g1077_p_spl_),
    .din2(g1078_p)
  );


  andX
  g_g1080_p
  (
    .dout(g1080_p),
    .din1(g1066_n_spl_),
    .din2(g1079_p_spl_)
  );


  orX
  g_g1080_n
  (
    .dout(g1080_n),
    .din1(g1066_p_spl_),
    .din2(g1079_n_spl_)
  );


  andX
  g_g1081_p
  (
    .dout(g1081_p),
    .din1(g1066_p_spl_),
    .din2(g1079_n_spl_)
  );


  orX
  g_g1081_n
  (
    .dout(g1081_n),
    .din1(g1066_n_spl_),
    .din2(g1079_p_spl_)
  );


  andX
  g_g1082_p
  (
    .dout(g1082_p),
    .din1(g1080_n_spl_),
    .din2(g1081_n)
  );


  orX
  g_g1082_n
  (
    .dout(g1082_n),
    .din1(g1080_p_spl_),
    .din2(g1081_p)
  );


  andX
  g_g1083_p
  (
    .dout(g1083_p),
    .din1(g1065_n_spl_),
    .din2(g1082_p_spl_)
  );


  orX
  g_g1083_n
  (
    .dout(g1083_n),
    .din1(g1065_p_spl_),
    .din2(g1082_n_spl_)
  );


  andX
  g_g1084_p
  (
    .dout(g1084_p),
    .din1(ffc_15_p_spl_001),
    .din2(ffc_126_p_spl_0)
  );


  orX
  g_g1084_n
  (
    .dout(g1084_n),
    .din1(ffc_15_n_spl_001),
    .din2(ffc_126_n_spl_0)
  );


  andX
  g_g1085_p
  (
    .dout(g1085_p),
    .din1(g1065_p_spl_),
    .din2(g1082_n_spl_)
  );


  orX
  g_g1085_n
  (
    .dout(g1085_n),
    .din1(g1065_n_spl_),
    .din2(g1082_p_spl_)
  );


  andX
  g_g1086_p
  (
    .dout(g1086_p),
    .din1(g1083_n_spl_),
    .din2(g1085_n)
  );


  orX
  g_g1086_n
  (
    .dout(g1086_n),
    .din1(g1083_p_spl_),
    .din2(g1085_p)
  );


  andX
  g_g1087_p
  (
    .dout(g1087_p),
    .din1(g1084_n_spl_),
    .din2(g1086_p_spl_)
  );


  orX
  g_g1087_n
  (
    .dout(g1087_n),
    .din1(g1084_p_spl_),
    .din2(g1086_n_spl_)
  );


  andX
  g_g1088_p
  (
    .dout(g1088_p),
    .din1(g1083_n_spl_),
    .din2(g1087_n_spl_)
  );


  orX
  g_g1088_n
  (
    .dout(g1088_n),
    .din1(g1083_p_spl_),
    .din2(g1087_p_spl_)
  );


  andX
  g_g1089_p
  (
    .dout(g1089_p),
    .din1(ffc_15_p_spl_010),
    .din2(ffc_127_p_spl_0)
  );


  orX
  g_g1089_n
  (
    .dout(g1089_n),
    .din1(ffc_15_n_spl_010),
    .din2(ffc_127_n_spl_)
  );


  andX
  g_g1090_p
  (
    .dout(g1090_p),
    .din1(g1077_n_spl_),
    .din2(g1080_n_spl_)
  );


  orX
  g_g1090_n
  (
    .dout(g1090_n),
    .din1(g1077_p_spl_),
    .din2(g1080_p_spl_)
  );


  andX
  g_g1091_p
  (
    .dout(g1091_p),
    .din1(ffc_128_p_spl_0),
    .din2(ffc_287_p_spl_100)
  );


  orX
  g_g1091_n
  (
    .dout(g1091_n),
    .din1(ffc_128_n_spl_0),
    .din2(ffc_287_n_spl_100)
  );


  andX
  g_g1092_p
  (
    .dout(g1092_p),
    .din1(g1071_n_spl_),
    .din2(g1074_n_spl_)
  );


  orX
  g_g1092_n
  (
    .dout(g1092_n),
    .din1(g1071_p_spl_),
    .din2(g1074_p_spl_)
  );


  andX
  g_g1093_p
  (
    .dout(g1093_p),
    .din1(g1024_p_spl_),
    .din2(g1026_n_spl_)
  );


  orX
  g_g1093_n
  (
    .dout(g1093_n),
    .din1(g1024_n_spl_),
    .din2(g1026_p_spl_)
  );


  andX
  g_g1094_p
  (
    .dout(g1094_p),
    .din1(g1027_n_spl_),
    .din2(g1093_n)
  );


  orX
  g_g1094_n
  (
    .dout(g1094_n),
    .din1(g1027_p_spl_),
    .din2(g1093_p)
  );


  andX
  g_g1095_p
  (
    .dout(g1095_p),
    .din1(g1092_n_spl_),
    .din2(g1094_p_spl_)
  );


  orX
  g_g1095_n
  (
    .dout(g1095_n),
    .din1(g1092_p_spl_),
    .din2(g1094_n_spl_)
  );


  andX
  g_g1096_p
  (
    .dout(g1096_p),
    .din1(g1092_p_spl_),
    .din2(g1094_n_spl_)
  );


  orX
  g_g1096_n
  (
    .dout(g1096_n),
    .din1(g1092_n_spl_),
    .din2(g1094_p_spl_)
  );


  andX
  g_g1097_p
  (
    .dout(g1097_p),
    .din1(g1095_n_spl_),
    .din2(g1096_n)
  );


  orX
  g_g1097_n
  (
    .dout(g1097_n),
    .din1(g1095_p_spl_),
    .din2(g1096_p)
  );


  andX
  g_g1098_p
  (
    .dout(g1098_p),
    .din1(g1091_n_spl_),
    .din2(g1097_p_spl_)
  );


  orX
  g_g1098_n
  (
    .dout(g1098_n),
    .din1(g1091_p_spl_),
    .din2(g1097_n_spl_)
  );


  andX
  g_g1099_p
  (
    .dout(g1099_p),
    .din1(g1091_p_spl_),
    .din2(g1097_n_spl_)
  );


  orX
  g_g1099_n
  (
    .dout(g1099_n),
    .din1(g1091_n_spl_),
    .din2(g1097_p_spl_)
  );


  andX
  g_g1100_p
  (
    .dout(g1100_p),
    .din1(g1098_n_spl_),
    .din2(g1099_n)
  );


  orX
  g_g1100_n
  (
    .dout(g1100_n),
    .din1(g1098_p_spl_),
    .din2(g1099_p)
  );


  andX
  g_g1101_p
  (
    .dout(g1101_p),
    .din1(g1090_n_spl_),
    .din2(g1100_p_spl_)
  );


  orX
  g_g1101_n
  (
    .dout(g1101_n),
    .din1(g1090_p_spl_),
    .din2(g1100_n_spl_)
  );


  andX
  g_g1102_p
  (
    .dout(g1102_p),
    .din1(g1090_p_spl_),
    .din2(g1100_n_spl_)
  );


  orX
  g_g1102_n
  (
    .dout(g1102_n),
    .din1(g1090_n_spl_),
    .din2(g1100_p_spl_)
  );


  andX
  g_g1103_p
  (
    .dout(g1103_p),
    .din1(g1101_n_spl_),
    .din2(g1102_n)
  );


  orX
  g_g1103_n
  (
    .dout(g1103_n),
    .din1(g1101_p_spl_),
    .din2(g1102_p)
  );


  andX
  g_g1104_p
  (
    .dout(g1104_p),
    .din1(g1089_n_spl_),
    .din2(g1103_p_spl_)
  );


  orX
  g_g1104_n
  (
    .dout(g1104_n),
    .din1(g1089_p_spl_),
    .din2(g1103_n_spl_)
  );


  andX
  g_g1105_p
  (
    .dout(g1105_p),
    .din1(g1089_p_spl_),
    .din2(g1103_n_spl_)
  );


  orX
  g_g1105_n
  (
    .dout(g1105_n),
    .din1(g1089_n_spl_),
    .din2(g1103_p_spl_)
  );


  andX
  g_g1106_p
  (
    .dout(g1106_p),
    .din1(g1104_n_spl_),
    .din2(g1105_n)
  );


  orX
  g_g1106_n
  (
    .dout(g1106_n),
    .din1(g1104_p_spl_),
    .din2(g1105_p)
  );


  andX
  g_g1107_p
  (
    .dout(g1107_p),
    .din1(g1088_n_spl_),
    .din2(g1106_p_spl_)
  );


  orX
  g_g1107_n
  (
    .dout(g1107_n),
    .din1(g1088_p_spl_),
    .din2(g1106_n_spl_)
  );


  andX
  g_g1108_p
  (
    .dout(g1108_p),
    .din1(ffc_123_p_spl_00),
    .din2(ffc_287_p_spl_100)
  );


  orX
  g_g1108_n
  (
    .dout(g1108_n),
    .din1(ffc_123_n_spl_0),
    .din2(ffc_287_n_spl_100)
  );


  andX
  g_g1109_p
  (
    .dout(g1109_p),
    .din1(ffc_306_p_spl_),
    .din2(ffc_307_n)
  );


  orX
  g_g1109_n
  (
    .dout(g1109_n),
    .din1(ffc_306_n_spl_),
    .din2(ffc_307_p)
  );


  andX
  g_g1110_p
  (
    .dout(g1110_p),
    .din1(g1108_n_spl_),
    .din2(g1109_p_spl_)
  );


  orX
  g_g1110_n
  (
    .dout(g1110_n),
    .din1(g1108_p_spl_),
    .din2(g1109_n_spl_)
  );


  andX
  g_g1111_p
  (
    .dout(g1111_p),
    .din1(ffc_306_p_spl_),
    .din2(g1110_n_spl_)
  );


  orX
  g_g1111_n
  (
    .dout(g1111_n),
    .din1(ffc_306_n_spl_),
    .din2(g1110_p_spl_)
  );


  andX
  g_g1112_p
  (
    .dout(g1112_p),
    .din1(ffc_124_p_spl_00),
    .din2(ffc_287_p_spl_101)
  );


  orX
  g_g1112_n
  (
    .dout(g1112_n),
    .din1(ffc_124_n_spl_0),
    .din2(ffc_287_n_spl_101)
  );


  andX
  g_g1113_p
  (
    .dout(g1113_p),
    .din1(ffc_308_p_spl_),
    .din2(ffc_309_n)
  );


  orX
  g_g1113_n
  (
    .dout(g1113_n),
    .din1(ffc_308_n_spl_),
    .din2(ffc_309_p)
  );


  andX
  g_g1114_p
  (
    .dout(g1114_p),
    .din1(g1112_n_spl_),
    .din2(g1113_p_spl_)
  );


  orX
  g_g1114_n
  (
    .dout(g1114_n),
    .din1(g1112_p_spl_),
    .din2(g1113_n_spl_)
  );


  andX
  g_g1115_p
  (
    .dout(g1115_p),
    .din1(g1112_p_spl_),
    .din2(g1113_n_spl_)
  );


  orX
  g_g1115_n
  (
    .dout(g1115_n),
    .din1(g1112_n_spl_),
    .din2(g1113_p_spl_)
  );


  andX
  g_g1116_p
  (
    .dout(g1116_p),
    .din1(g1114_n_spl_),
    .din2(g1115_n)
  );


  orX
  g_g1116_n
  (
    .dout(g1116_n),
    .din1(g1114_p_spl_),
    .din2(g1115_p)
  );


  andX
  g_g1117_p
  (
    .dout(g1117_p),
    .din1(g1111_n_spl_),
    .din2(g1116_p_spl_)
  );


  orX
  g_g1117_n
  (
    .dout(g1117_n),
    .din1(g1111_p_spl_),
    .din2(g1116_n_spl_)
  );


  andX
  g_g1118_p
  (
    .dout(g1118_p),
    .din1(ffc_15_p_spl_010),
    .din2(ffc_123_p_spl_00)
  );


  orX
  g_g1118_n
  (
    .dout(g1118_n),
    .din1(ffc_15_n_spl_010),
    .din2(ffc_123_n_spl_0)
  );


  andX
  g_g1119_p
  (
    .dout(g1119_p),
    .din1(g1111_p_spl_),
    .din2(g1116_n_spl_)
  );


  orX
  g_g1119_n
  (
    .dout(g1119_n),
    .din1(g1111_n_spl_),
    .din2(g1116_p_spl_)
  );


  andX
  g_g1120_p
  (
    .dout(g1120_p),
    .din1(g1117_n_spl_),
    .din2(g1119_n)
  );


  orX
  g_g1120_n
  (
    .dout(g1120_n),
    .din1(g1117_p_spl_),
    .din2(g1119_p)
  );


  andX
  g_g1121_p
  (
    .dout(g1121_p),
    .din1(g1118_n_spl_),
    .din2(g1120_p_spl_)
  );


  orX
  g_g1121_n
  (
    .dout(g1121_n),
    .din1(g1118_p_spl_),
    .din2(g1120_n_spl_)
  );


  andX
  g_g1122_p
  (
    .dout(g1122_p),
    .din1(g1117_n_spl_),
    .din2(g1121_n_spl_)
  );


  orX
  g_g1122_n
  (
    .dout(g1122_n),
    .din1(g1117_p_spl_),
    .din2(g1121_p_spl_)
  );


  andX
  g_g1123_p
  (
    .dout(g1123_p),
    .din1(ffc_15_p_spl_011),
    .din2(ffc_124_p_spl_00)
  );


  orX
  g_g1123_n
  (
    .dout(g1123_n),
    .din1(ffc_15_n_spl_011),
    .din2(ffc_124_n_spl_0)
  );


  andX
  g_g1124_p
  (
    .dout(g1124_p),
    .din1(ffc_308_p_spl_),
    .din2(g1114_n_spl_)
  );


  orX
  g_g1124_n
  (
    .dout(g1124_n),
    .din1(ffc_308_n_spl_),
    .din2(g1114_p_spl_)
  );


  andX
  g_g1125_p
  (
    .dout(g1125_p),
    .din1(ffc_125_p_spl_0),
    .din2(ffc_287_p_spl_101)
  );


  orX
  g_g1125_n
  (
    .dout(g1125_n),
    .din1(ffc_125_n_spl_0),
    .din2(ffc_287_n_spl_101)
  );


  andX
  g_g1126_p
  (
    .dout(g1126_p),
    .din1(ffc_227_p),
    .din2(ffc_255_n)
  );


  orX
  g_g1126_n
  (
    .dout(g1126_n),
    .din1(ffc_227_n),
    .din2(ffc_255_p)
  );


  andX
  g_g1127_p
  (
    .dout(g1127_p),
    .din1(ffc_288_n_spl_),
    .din2(ffc_289_n)
  );


  orX
  g_g1127_n
  (
    .dout(g1127_n),
    .din1(ffc_288_p_spl_),
    .din2(ffc_289_p)
  );


  andX
  g_g1128_p
  (
    .dout(g1128_p),
    .din1(g1126_n_spl_),
    .din2(g1127_p_spl_)
  );


  orX
  g_g1128_n
  (
    .dout(g1128_n),
    .din1(g1126_p_spl_),
    .din2(g1127_n_spl_)
  );


  andX
  g_g1129_p
  (
    .dout(g1129_p),
    .din1(g1126_p_spl_),
    .din2(g1127_n_spl_)
  );


  orX
  g_g1129_n
  (
    .dout(g1129_n),
    .din1(g1126_n_spl_),
    .din2(g1127_p_spl_)
  );


  andX
  g_g1130_p
  (
    .dout(g1130_p),
    .din1(g1128_n_spl_),
    .din2(g1129_n)
  );


  orX
  g_g1130_n
  (
    .dout(g1130_n),
    .din1(g1128_p_spl_),
    .din2(g1129_p)
  );


  andX
  g_g1131_p
  (
    .dout(g1131_p),
    .din1(g1125_n_spl_),
    .din2(g1130_p_spl_)
  );


  orX
  g_g1131_n
  (
    .dout(g1131_n),
    .din1(g1125_p_spl_),
    .din2(g1130_n_spl_)
  );


  andX
  g_g1132_p
  (
    .dout(g1132_p),
    .din1(g1125_p_spl_),
    .din2(g1130_n_spl_)
  );


  orX
  g_g1132_n
  (
    .dout(g1132_n),
    .din1(g1125_n_spl_),
    .din2(g1130_p_spl_)
  );


  andX
  g_g1133_p
  (
    .dout(g1133_p),
    .din1(g1131_n_spl_),
    .din2(g1132_n)
  );


  orX
  g_g1133_n
  (
    .dout(g1133_n),
    .din1(g1131_p_spl_),
    .din2(g1132_p)
  );


  andX
  g_g1134_p
  (
    .dout(g1134_p),
    .din1(g1124_n_spl_),
    .din2(g1133_p_spl_)
  );


  orX
  g_g1134_n
  (
    .dout(g1134_n),
    .din1(g1124_p_spl_),
    .din2(g1133_n_spl_)
  );


  andX
  g_g1135_p
  (
    .dout(g1135_p),
    .din1(g1124_p_spl_),
    .din2(g1133_n_spl_)
  );


  orX
  g_g1135_n
  (
    .dout(g1135_n),
    .din1(g1124_n_spl_),
    .din2(g1133_p_spl_)
  );


  andX
  g_g1136_p
  (
    .dout(g1136_p),
    .din1(g1134_n_spl_),
    .din2(g1135_n)
  );


  orX
  g_g1136_n
  (
    .dout(g1136_n),
    .din1(g1134_p_spl_),
    .din2(g1135_p)
  );


  andX
  g_g1137_p
  (
    .dout(g1137_p),
    .din1(g1123_n_spl_),
    .din2(g1136_p_spl_)
  );


  orX
  g_g1137_n
  (
    .dout(g1137_n),
    .din1(g1123_p_spl_),
    .din2(g1136_n_spl_)
  );


  andX
  g_g1138_p
  (
    .dout(g1138_p),
    .din1(g1123_p_spl_),
    .din2(g1136_n_spl_)
  );


  orX
  g_g1138_n
  (
    .dout(g1138_n),
    .din1(g1123_n_spl_),
    .din2(g1136_p_spl_)
  );


  andX
  g_g1139_p
  (
    .dout(g1139_p),
    .din1(g1137_n_spl_),
    .din2(g1138_n)
  );


  orX
  g_g1139_n
  (
    .dout(g1139_n),
    .din1(g1137_p_spl_),
    .din2(g1138_p)
  );


  andX
  g_g1140_p
  (
    .dout(g1140_p),
    .din1(g1122_n_spl_),
    .din2(g1139_p_spl_)
  );


  orX
  g_g1140_n
  (
    .dout(g1140_n),
    .din1(g1122_p_spl_),
    .din2(g1139_n_spl_)
  );


  andX
  g_g1141_p
  (
    .dout(g1141_p),
    .din1(ffc_17_p_spl_001),
    .din2(ffc_123_p_spl_0)
  );


  orX
  g_g1141_n
  (
    .dout(g1141_n),
    .din1(ffc_17_n_spl_001),
    .din2(ffc_123_n_spl_1)
  );


  andX
  g_g1142_p
  (
    .dout(g1142_p),
    .din1(g1122_p_spl_),
    .din2(g1139_n_spl_)
  );


  orX
  g_g1142_n
  (
    .dout(g1142_n),
    .din1(g1122_n_spl_),
    .din2(g1139_p_spl_)
  );


  andX
  g_g1143_p
  (
    .dout(g1143_p),
    .din1(g1140_n_spl_),
    .din2(g1142_n)
  );


  orX
  g_g1143_n
  (
    .dout(g1143_n),
    .din1(g1140_p_spl_),
    .din2(g1142_p)
  );


  andX
  g_g1144_p
  (
    .dout(g1144_p),
    .din1(g1141_n_spl_),
    .din2(g1143_p_spl_)
  );


  orX
  g_g1144_n
  (
    .dout(g1144_n),
    .din1(g1141_p_spl_),
    .din2(g1143_n_spl_)
  );


  andX
  g_g1145_p
  (
    .dout(g1145_p),
    .din1(g1140_n_spl_),
    .din2(g1144_n_spl_)
  );


  orX
  g_g1145_n
  (
    .dout(g1145_n),
    .din1(g1140_p_spl_),
    .din2(g1144_p_spl_)
  );


  andX
  g_g1146_p
  (
    .dout(g1146_p),
    .din1(ffc_17_p_spl_001),
    .din2(ffc_124_p_spl_0)
  );


  orX
  g_g1146_n
  (
    .dout(g1146_n),
    .din1(ffc_17_n_spl_001),
    .din2(ffc_124_n_spl_)
  );


  andX
  g_g1147_p
  (
    .dout(g1147_p),
    .din1(g1134_n_spl_),
    .din2(g1137_n_spl_)
  );


  orX
  g_g1147_n
  (
    .dout(g1147_n),
    .din1(g1134_p_spl_),
    .din2(g1137_p_spl_)
  );


  andX
  g_g1148_p
  (
    .dout(g1148_p),
    .din1(ffc_15_p_spl_011),
    .din2(ffc_125_p_spl_0)
  );


  orX
  g_g1148_n
  (
    .dout(g1148_n),
    .din1(ffc_15_n_spl_011),
    .din2(ffc_125_n_spl_0)
  );


  andX
  g_g1149_p
  (
    .dout(g1149_p),
    .din1(g1128_n_spl_),
    .din2(g1131_n_spl_)
  );


  orX
  g_g1149_n
  (
    .dout(g1149_n),
    .din1(g1128_p_spl_),
    .din2(g1131_p_spl_)
  );


  andX
  g_g1150_p
  (
    .dout(g1150_p),
    .din1(g1061_p_spl_),
    .din2(g1063_n_spl_)
  );


  orX
  g_g1150_n
  (
    .dout(g1150_n),
    .din1(g1061_n_spl_),
    .din2(g1063_p_spl_)
  );


  andX
  g_g1151_p
  (
    .dout(g1151_p),
    .din1(g1064_n_spl_),
    .din2(g1150_n)
  );


  orX
  g_g1151_n
  (
    .dout(g1151_n),
    .din1(g1064_p_spl_),
    .din2(g1150_p)
  );


  andX
  g_g1152_p
  (
    .dout(g1152_p),
    .din1(g1149_n_spl_),
    .din2(g1151_p_spl_)
  );


  orX
  g_g1152_n
  (
    .dout(g1152_n),
    .din1(g1149_p_spl_),
    .din2(g1151_n_spl_)
  );


  andX
  g_g1153_p
  (
    .dout(g1153_p),
    .din1(g1149_p_spl_),
    .din2(g1151_n_spl_)
  );


  orX
  g_g1153_n
  (
    .dout(g1153_n),
    .din1(g1149_n_spl_),
    .din2(g1151_p_spl_)
  );


  andX
  g_g1154_p
  (
    .dout(g1154_p),
    .din1(g1152_n_spl_),
    .din2(g1153_n)
  );


  orX
  g_g1154_n
  (
    .dout(g1154_n),
    .din1(g1152_p_spl_),
    .din2(g1153_p)
  );


  andX
  g_g1155_p
  (
    .dout(g1155_p),
    .din1(g1148_n_spl_),
    .din2(g1154_p_spl_)
  );


  orX
  g_g1155_n
  (
    .dout(g1155_n),
    .din1(g1148_p_spl_),
    .din2(g1154_n_spl_)
  );


  andX
  g_g1156_p
  (
    .dout(g1156_p),
    .din1(g1148_p_spl_),
    .din2(g1154_n_spl_)
  );


  orX
  g_g1156_n
  (
    .dout(g1156_n),
    .din1(g1148_n_spl_),
    .din2(g1154_p_spl_)
  );


  andX
  g_g1157_p
  (
    .dout(g1157_p),
    .din1(g1155_n_spl_),
    .din2(g1156_n)
  );


  orX
  g_g1157_n
  (
    .dout(g1157_n),
    .din1(g1155_p_spl_),
    .din2(g1156_p)
  );


  andX
  g_g1158_p
  (
    .dout(g1158_p),
    .din1(g1147_n_spl_),
    .din2(g1157_p_spl_)
  );


  orX
  g_g1158_n
  (
    .dout(g1158_n),
    .din1(g1147_p_spl_),
    .din2(g1157_n_spl_)
  );


  andX
  g_g1159_p
  (
    .dout(g1159_p),
    .din1(g1147_p_spl_),
    .din2(g1157_n_spl_)
  );


  orX
  g_g1159_n
  (
    .dout(g1159_n),
    .din1(g1147_n_spl_),
    .din2(g1157_p_spl_)
  );


  andX
  g_g1160_p
  (
    .dout(g1160_p),
    .din1(g1158_n_spl_),
    .din2(g1159_n)
  );


  orX
  g_g1160_n
  (
    .dout(g1160_n),
    .din1(g1158_p_spl_),
    .din2(g1159_p)
  );


  andX
  g_g1161_p
  (
    .dout(g1161_p),
    .din1(g1146_n_spl_),
    .din2(g1160_p_spl_)
  );


  orX
  g_g1161_n
  (
    .dout(g1161_n),
    .din1(g1146_p_spl_),
    .din2(g1160_n_spl_)
  );


  andX
  g_g1162_p
  (
    .dout(g1162_p),
    .din1(g1146_p_spl_),
    .din2(g1160_n_spl_)
  );


  orX
  g_g1162_n
  (
    .dout(g1162_n),
    .din1(g1146_n_spl_),
    .din2(g1160_p_spl_)
  );


  andX
  g_g1163_p
  (
    .dout(g1163_p),
    .din1(g1161_n_spl_),
    .din2(g1162_n)
  );


  orX
  g_g1163_n
  (
    .dout(g1163_n),
    .din1(g1161_p_spl_),
    .din2(g1162_p)
  );


  andX
  g_g1164_p
  (
    .dout(g1164_p),
    .din1(g1145_n_spl_),
    .din2(g1163_p_spl_)
  );


  orX
  g_g1164_n
  (
    .dout(g1164_n),
    .din1(g1145_p_spl_),
    .din2(g1163_n_spl_)
  );


  andX
  g_g1165_p
  (
    .dout(g1165_p),
    .din1(ffc_120_p_spl_00),
    .din2(ffc_287_p_spl_110)
  );


  orX
  g_g1165_n
  (
    .dout(g1165_n),
    .din1(ffc_120_n_spl_00),
    .din2(ffc_287_n_spl_110)
  );


  andX
  g_g1166_p
  (
    .dout(g1166_p),
    .din1(ffc_300_p_spl_),
    .din2(ffc_301_n)
  );


  orX
  g_g1166_n
  (
    .dout(g1166_n),
    .din1(ffc_300_n_spl_),
    .din2(ffc_301_p)
  );


  andX
  g_g1167_p
  (
    .dout(g1167_p),
    .din1(g1165_n_spl_),
    .din2(g1166_p_spl_)
  );


  orX
  g_g1167_n
  (
    .dout(g1167_n),
    .din1(g1165_p_spl_),
    .din2(g1166_n_spl_)
  );


  andX
  g_g1168_p
  (
    .dout(g1168_p),
    .din1(ffc_300_p_spl_),
    .din2(g1167_n_spl_)
  );


  orX
  g_g1168_n
  (
    .dout(g1168_n),
    .din1(ffc_300_n_spl_),
    .din2(g1167_p_spl_)
  );


  andX
  g_g1169_p
  (
    .dout(g1169_p),
    .din1(ffc_121_p_spl_00),
    .din2(ffc_287_p_spl_110)
  );


  orX
  g_g1169_n
  (
    .dout(g1169_n),
    .din1(ffc_121_n_spl_0),
    .din2(ffc_287_n_spl_110)
  );


  andX
  g_g1170_p
  (
    .dout(g1170_p),
    .din1(ffc_302_p_spl_),
    .din2(ffc_303_n)
  );


  orX
  g_g1170_n
  (
    .dout(g1170_n),
    .din1(ffc_302_n_spl_),
    .din2(ffc_303_p)
  );


  andX
  g_g1171_p
  (
    .dout(g1171_p),
    .din1(g1169_n_spl_),
    .din2(g1170_p_spl_)
  );


  orX
  g_g1171_n
  (
    .dout(g1171_n),
    .din1(g1169_p_spl_),
    .din2(g1170_n_spl_)
  );


  andX
  g_g1172_p
  (
    .dout(g1172_p),
    .din1(g1169_p_spl_),
    .din2(g1170_n_spl_)
  );


  orX
  g_g1172_n
  (
    .dout(g1172_n),
    .din1(g1169_n_spl_),
    .din2(g1170_p_spl_)
  );


  andX
  g_g1173_p
  (
    .dout(g1173_p),
    .din1(g1171_n_spl_),
    .din2(g1172_n)
  );


  orX
  g_g1173_n
  (
    .dout(g1173_n),
    .din1(g1171_p_spl_),
    .din2(g1172_p)
  );


  andX
  g_g1174_p
  (
    .dout(g1174_p),
    .din1(g1168_n_spl_),
    .din2(g1173_p_spl_)
  );


  orX
  g_g1174_n
  (
    .dout(g1174_n),
    .din1(g1168_p_spl_),
    .din2(g1173_n_spl_)
  );


  andX
  g_g1175_p
  (
    .dout(g1175_p),
    .din1(ffc_15_p_spl_100),
    .din2(ffc_120_p_spl_00)
  );


  orX
  g_g1175_n
  (
    .dout(g1175_n),
    .din1(ffc_15_n_spl_100),
    .din2(ffc_120_n_spl_00)
  );


  andX
  g_g1176_p
  (
    .dout(g1176_p),
    .din1(g1168_p_spl_),
    .din2(g1173_n_spl_)
  );


  orX
  g_g1176_n
  (
    .dout(g1176_n),
    .din1(g1168_n_spl_),
    .din2(g1173_p_spl_)
  );


  andX
  g_g1177_p
  (
    .dout(g1177_p),
    .din1(g1174_n_spl_),
    .din2(g1176_n)
  );


  orX
  g_g1177_n
  (
    .dout(g1177_n),
    .din1(g1174_p_spl_),
    .din2(g1176_p)
  );


  andX
  g_g1178_p
  (
    .dout(g1178_p),
    .din1(g1175_n_spl_),
    .din2(g1177_p_spl_)
  );


  orX
  g_g1178_n
  (
    .dout(g1178_n),
    .din1(g1175_p_spl_),
    .din2(g1177_n_spl_)
  );


  andX
  g_g1179_p
  (
    .dout(g1179_p),
    .din1(g1174_n_spl_),
    .din2(g1178_n_spl_)
  );


  orX
  g_g1179_n
  (
    .dout(g1179_n),
    .din1(g1174_p_spl_),
    .din2(g1178_p_spl_)
  );


  andX
  g_g1180_p
  (
    .dout(g1180_p),
    .din1(ffc_15_p_spl_100),
    .din2(ffc_121_p_spl_00)
  );


  orX
  g_g1180_n
  (
    .dout(g1180_n),
    .din1(ffc_15_n_spl_100),
    .din2(ffc_121_n_spl_0)
  );


  andX
  g_g1181_p
  (
    .dout(g1181_p),
    .din1(ffc_302_p_spl_),
    .din2(g1171_n_spl_)
  );


  orX
  g_g1181_n
  (
    .dout(g1181_n),
    .din1(ffc_302_n_spl_),
    .din2(g1171_p_spl_)
  );


  andX
  g_g1182_p
  (
    .dout(g1182_p),
    .din1(ffc_122_p_spl_00),
    .din2(ffc_287_p_spl_111)
  );


  orX
  g_g1182_n
  (
    .dout(g1182_n),
    .din1(ffc_122_n_spl_0),
    .din2(ffc_287_n_spl_111)
  );


  andX
  g_g1183_p
  (
    .dout(g1183_p),
    .din1(ffc_304_p_spl_),
    .din2(ffc_305_n)
  );


  orX
  g_g1183_n
  (
    .dout(g1183_n),
    .din1(ffc_304_n_spl_),
    .din2(ffc_305_p)
  );


  andX
  g_g1184_p
  (
    .dout(g1184_p),
    .din1(g1182_n_spl_),
    .din2(g1183_p_spl_)
  );


  orX
  g_g1184_n
  (
    .dout(g1184_n),
    .din1(g1182_p_spl_),
    .din2(g1183_n_spl_)
  );


  andX
  g_g1185_p
  (
    .dout(g1185_p),
    .din1(g1182_p_spl_),
    .din2(g1183_n_spl_)
  );


  orX
  g_g1185_n
  (
    .dout(g1185_n),
    .din1(g1182_n_spl_),
    .din2(g1183_p_spl_)
  );


  andX
  g_g1186_p
  (
    .dout(g1186_p),
    .din1(g1184_n_spl_),
    .din2(g1185_n)
  );


  orX
  g_g1186_n
  (
    .dout(g1186_n),
    .din1(g1184_p_spl_),
    .din2(g1185_p)
  );


  andX
  g_g1187_p
  (
    .dout(g1187_p),
    .din1(g1181_n_spl_),
    .din2(g1186_p_spl_)
  );


  orX
  g_g1187_n
  (
    .dout(g1187_n),
    .din1(g1181_p_spl_),
    .din2(g1186_n_spl_)
  );


  andX
  g_g1188_p
  (
    .dout(g1188_p),
    .din1(g1181_p_spl_),
    .din2(g1186_n_spl_)
  );


  orX
  g_g1188_n
  (
    .dout(g1188_n),
    .din1(g1181_n_spl_),
    .din2(g1186_p_spl_)
  );


  andX
  g_g1189_p
  (
    .dout(g1189_p),
    .din1(g1187_n_spl_),
    .din2(g1188_n)
  );


  orX
  g_g1189_n
  (
    .dout(g1189_n),
    .din1(g1187_p_spl_),
    .din2(g1188_p)
  );


  andX
  g_g1190_p
  (
    .dout(g1190_p),
    .din1(g1180_n_spl_),
    .din2(g1189_p_spl_)
  );


  orX
  g_g1190_n
  (
    .dout(g1190_n),
    .din1(g1180_p_spl_),
    .din2(g1189_n_spl_)
  );


  andX
  g_g1191_p
  (
    .dout(g1191_p),
    .din1(g1180_p_spl_),
    .din2(g1189_n_spl_)
  );


  orX
  g_g1191_n
  (
    .dout(g1191_n),
    .din1(g1180_n_spl_),
    .din2(g1189_p_spl_)
  );


  andX
  g_g1192_p
  (
    .dout(g1192_p),
    .din1(g1190_n_spl_),
    .din2(g1191_n)
  );


  orX
  g_g1192_n
  (
    .dout(g1192_n),
    .din1(g1190_p_spl_),
    .din2(g1191_p)
  );


  andX
  g_g1193_p
  (
    .dout(g1193_p),
    .din1(g1179_n_spl_),
    .din2(g1192_p_spl_)
  );


  orX
  g_g1193_n
  (
    .dout(g1193_n),
    .din1(g1179_p_spl_),
    .din2(g1192_n_spl_)
  );


  andX
  g_g1194_p
  (
    .dout(g1194_p),
    .din1(ffc_17_p_spl_010),
    .din2(ffc_120_p_spl_01)
  );


  orX
  g_g1194_n
  (
    .dout(g1194_n),
    .din1(ffc_17_n_spl_010),
    .din2(ffc_120_n_spl_0)
  );


  andX
  g_g1195_p
  (
    .dout(g1195_p),
    .din1(g1179_p_spl_),
    .din2(g1192_n_spl_)
  );


  orX
  g_g1195_n
  (
    .dout(g1195_n),
    .din1(g1179_n_spl_),
    .din2(g1192_p_spl_)
  );


  andX
  g_g1196_p
  (
    .dout(g1196_p),
    .din1(g1193_n_spl_),
    .din2(g1195_n)
  );


  orX
  g_g1196_n
  (
    .dout(g1196_n),
    .din1(g1193_p_spl_),
    .din2(g1195_p)
  );


  andX
  g_g1197_p
  (
    .dout(g1197_p),
    .din1(g1194_n_spl_),
    .din2(g1196_p_spl_)
  );


  orX
  g_g1197_n
  (
    .dout(g1197_n),
    .din1(g1194_p_spl_),
    .din2(g1196_n_spl_)
  );


  andX
  g_g1198_p
  (
    .dout(g1198_p),
    .din1(g1193_n_spl_),
    .din2(g1197_n_spl_)
  );


  orX
  g_g1198_n
  (
    .dout(g1198_n),
    .din1(g1193_p_spl_),
    .din2(g1197_p_spl_)
  );


  andX
  g_g1199_p
  (
    .dout(g1199_p),
    .din1(ffc_17_p_spl_010),
    .din2(ffc_121_p_spl_01)
  );


  orX
  g_g1199_n
  (
    .dout(g1199_n),
    .din1(ffc_17_n_spl_010),
    .din2(ffc_121_n_spl_1)
  );


  andX
  g_g1200_p
  (
    .dout(g1200_p),
    .din1(g1187_n_spl_),
    .din2(g1190_n_spl_)
  );


  orX
  g_g1200_n
  (
    .dout(g1200_n),
    .din1(g1187_p_spl_),
    .din2(g1190_p_spl_)
  );


  andX
  g_g1201_p
  (
    .dout(g1201_p),
    .din1(ffc_15_p_spl_101),
    .din2(ffc_122_p_spl_00)
  );


  orX
  g_g1201_n
  (
    .dout(g1201_n),
    .din1(ffc_15_n_spl_101),
    .din2(ffc_122_n_spl_0)
  );


  andX
  g_g1202_p
  (
    .dout(g1202_p),
    .din1(ffc_304_p_spl_),
    .din2(g1184_n_spl_)
  );


  orX
  g_g1202_n
  (
    .dout(g1202_n),
    .din1(ffc_304_n_spl_),
    .din2(g1184_p_spl_)
  );


  andX
  g_g1203_p
  (
    .dout(g1203_p),
    .din1(g1108_p_spl_),
    .din2(g1109_n_spl_)
  );


  orX
  g_g1203_n
  (
    .dout(g1203_n),
    .din1(g1108_n_spl_),
    .din2(g1109_p_spl_)
  );


  andX
  g_g1204_p
  (
    .dout(g1204_p),
    .din1(g1110_n_spl_),
    .din2(g1203_n)
  );


  orX
  g_g1204_n
  (
    .dout(g1204_n),
    .din1(g1110_p_spl_),
    .din2(g1203_p)
  );


  andX
  g_g1205_p
  (
    .dout(g1205_p),
    .din1(g1202_n_spl_),
    .din2(g1204_p_spl_)
  );


  orX
  g_g1205_n
  (
    .dout(g1205_n),
    .din1(g1202_p_spl_),
    .din2(g1204_n_spl_)
  );


  andX
  g_g1206_p
  (
    .dout(g1206_p),
    .din1(g1202_p_spl_),
    .din2(g1204_n_spl_)
  );


  orX
  g_g1206_n
  (
    .dout(g1206_n),
    .din1(g1202_n_spl_),
    .din2(g1204_p_spl_)
  );


  andX
  g_g1207_p
  (
    .dout(g1207_p),
    .din1(g1205_n_spl_),
    .din2(g1206_n)
  );


  orX
  g_g1207_n
  (
    .dout(g1207_n),
    .din1(g1205_p_spl_),
    .din2(g1206_p)
  );


  andX
  g_g1208_p
  (
    .dout(g1208_p),
    .din1(g1201_n_spl_),
    .din2(g1207_p_spl_)
  );


  orX
  g_g1208_n
  (
    .dout(g1208_n),
    .din1(g1201_p_spl_),
    .din2(g1207_n_spl_)
  );


  andX
  g_g1209_p
  (
    .dout(g1209_p),
    .din1(g1201_p_spl_),
    .din2(g1207_n_spl_)
  );


  orX
  g_g1209_n
  (
    .dout(g1209_n),
    .din1(g1201_n_spl_),
    .din2(g1207_p_spl_)
  );


  andX
  g_g1210_p
  (
    .dout(g1210_p),
    .din1(g1208_n_spl_),
    .din2(g1209_n)
  );


  orX
  g_g1210_n
  (
    .dout(g1210_n),
    .din1(g1208_p_spl_),
    .din2(g1209_p)
  );


  andX
  g_g1211_p
  (
    .dout(g1211_p),
    .din1(g1200_n_spl_),
    .din2(g1210_p_spl_)
  );


  orX
  g_g1211_n
  (
    .dout(g1211_n),
    .din1(g1200_p_spl_),
    .din2(g1210_n_spl_)
  );


  andX
  g_g1212_p
  (
    .dout(g1212_p),
    .din1(g1200_p_spl_),
    .din2(g1210_n_spl_)
  );


  orX
  g_g1212_n
  (
    .dout(g1212_n),
    .din1(g1200_n_spl_),
    .din2(g1210_p_spl_)
  );


  andX
  g_g1213_p
  (
    .dout(g1213_p),
    .din1(g1211_n_spl_),
    .din2(g1212_n)
  );


  orX
  g_g1213_n
  (
    .dout(g1213_n),
    .din1(g1211_p_spl_),
    .din2(g1212_p)
  );


  andX
  g_g1214_p
  (
    .dout(g1214_p),
    .din1(g1199_n_spl_),
    .din2(g1213_p_spl_)
  );


  orX
  g_g1214_n
  (
    .dout(g1214_n),
    .din1(g1199_p_spl_),
    .din2(g1213_n_spl_)
  );


  andX
  g_g1215_p
  (
    .dout(g1215_p),
    .din1(g1199_p_spl_),
    .din2(g1213_n_spl_)
  );


  orX
  g_g1215_n
  (
    .dout(g1215_n),
    .din1(g1199_n_spl_),
    .din2(g1213_p_spl_)
  );


  andX
  g_g1216_p
  (
    .dout(g1216_p),
    .din1(g1214_n_spl_),
    .din2(g1215_n)
  );


  orX
  g_g1216_n
  (
    .dout(g1216_n),
    .din1(g1214_p_spl_),
    .din2(g1215_p)
  );


  andX
  g_g1217_p
  (
    .dout(g1217_p),
    .din1(g1198_n_spl_),
    .din2(g1216_p_spl_)
  );


  orX
  g_g1217_n
  (
    .dout(g1217_n),
    .din1(g1198_p_spl_),
    .din2(g1216_n_spl_)
  );


  andX
  g_g1218_p
  (
    .dout(g1218_p),
    .din1(ffc_19_p_spl_000),
    .din2(ffc_120_p_spl_01)
  );


  orX
  g_g1218_n
  (
    .dout(g1218_n),
    .din1(ffc_19_n_spl_00),
    .din2(ffc_120_n_spl_1)
  );


  andX
  g_g1219_p
  (
    .dout(g1219_p),
    .din1(g1198_p_spl_),
    .din2(g1216_n_spl_)
  );


  orX
  g_g1219_n
  (
    .dout(g1219_n),
    .din1(g1198_n_spl_),
    .din2(g1216_p_spl_)
  );


  andX
  g_g1220_p
  (
    .dout(g1220_p),
    .din1(g1217_n_spl_),
    .din2(g1219_n)
  );


  orX
  g_g1220_n
  (
    .dout(g1220_n),
    .din1(g1217_p_spl_),
    .din2(g1219_p)
  );


  andX
  g_g1221_p
  (
    .dout(g1221_p),
    .din1(g1218_n_spl_),
    .din2(g1220_p_spl_)
  );


  orX
  g_g1221_n
  (
    .dout(g1221_n),
    .din1(g1218_p_spl_),
    .din2(g1220_n_spl_)
  );


  andX
  g_g1222_p
  (
    .dout(g1222_p),
    .din1(g1217_n_spl_),
    .din2(g1221_n_spl_)
  );


  orX
  g_g1222_n
  (
    .dout(g1222_n),
    .din1(g1217_p_spl_),
    .din2(g1221_p_spl_)
  );


  andX
  g_g1223_p
  (
    .dout(g1223_p),
    .din1(ffc_19_p_spl_001),
    .din2(ffc_121_p_spl_01)
  );


  orX
  g_g1223_n
  (
    .dout(g1223_n),
    .din1(ffc_19_n_spl_01),
    .din2(ffc_121_n_spl_1)
  );


  andX
  g_g1224_p
  (
    .dout(g1224_p),
    .din1(g1211_n_spl_),
    .din2(g1214_n_spl_)
  );


  orX
  g_g1224_n
  (
    .dout(g1224_n),
    .din1(g1211_p_spl_),
    .din2(g1214_p_spl_)
  );


  andX
  g_g1225_p
  (
    .dout(g1225_p),
    .din1(ffc_17_p_spl_011),
    .din2(ffc_122_p_spl_0)
  );


  orX
  g_g1225_n
  (
    .dout(g1225_n),
    .din1(ffc_17_n_spl_01),
    .din2(ffc_122_n_spl_1)
  );


  andX
  g_g1226_p
  (
    .dout(g1226_p),
    .din1(g1205_n_spl_),
    .din2(g1208_n_spl_)
  );


  orX
  g_g1226_n
  (
    .dout(g1226_n),
    .din1(g1205_p_spl_),
    .din2(g1208_p_spl_)
  );


  andX
  g_g1227_p
  (
    .dout(g1227_p),
    .din1(g1118_p_spl_),
    .din2(g1120_n_spl_)
  );


  orX
  g_g1227_n
  (
    .dout(g1227_n),
    .din1(g1118_n_spl_),
    .din2(g1120_p_spl_)
  );


  andX
  g_g1228_p
  (
    .dout(g1228_p),
    .din1(g1121_n_spl_),
    .din2(g1227_n)
  );


  orX
  g_g1228_n
  (
    .dout(g1228_n),
    .din1(g1121_p_spl_),
    .din2(g1227_p)
  );


  andX
  g_g1229_p
  (
    .dout(g1229_p),
    .din1(g1226_n_spl_),
    .din2(g1228_p_spl_)
  );


  orX
  g_g1229_n
  (
    .dout(g1229_n),
    .din1(g1226_p_spl_),
    .din2(g1228_n_spl_)
  );


  andX
  g_g1230_p
  (
    .dout(g1230_p),
    .din1(g1226_p_spl_),
    .din2(g1228_n_spl_)
  );


  orX
  g_g1230_n
  (
    .dout(g1230_n),
    .din1(g1226_n_spl_),
    .din2(g1228_p_spl_)
  );


  andX
  g_g1231_p
  (
    .dout(g1231_p),
    .din1(g1229_n_spl_),
    .din2(g1230_n)
  );


  orX
  g_g1231_n
  (
    .dout(g1231_n),
    .din1(g1229_p_spl_),
    .din2(g1230_p)
  );


  andX
  g_g1232_p
  (
    .dout(g1232_p),
    .din1(g1225_n_spl_),
    .din2(g1231_p_spl_)
  );


  orX
  g_g1232_n
  (
    .dout(g1232_n),
    .din1(g1225_p_spl_),
    .din2(g1231_n_spl_)
  );


  andX
  g_g1233_p
  (
    .dout(g1233_p),
    .din1(g1225_p_spl_),
    .din2(g1231_n_spl_)
  );


  orX
  g_g1233_n
  (
    .dout(g1233_n),
    .din1(g1225_n_spl_),
    .din2(g1231_p_spl_)
  );


  andX
  g_g1234_p
  (
    .dout(g1234_p),
    .din1(g1232_n_spl_),
    .din2(g1233_n)
  );


  orX
  g_g1234_n
  (
    .dout(g1234_n),
    .din1(g1232_p_spl_),
    .din2(g1233_p)
  );


  andX
  g_g1235_p
  (
    .dout(g1235_p),
    .din1(g1224_n_spl_),
    .din2(g1234_p_spl_)
  );


  orX
  g_g1235_n
  (
    .dout(g1235_n),
    .din1(g1224_p_spl_),
    .din2(g1234_n_spl_)
  );


  andX
  g_g1236_p
  (
    .dout(g1236_p),
    .din1(g1224_p_spl_),
    .din2(g1234_n_spl_)
  );


  orX
  g_g1236_n
  (
    .dout(g1236_n),
    .din1(g1224_n_spl_),
    .din2(g1234_p_spl_)
  );


  andX
  g_g1237_p
  (
    .dout(g1237_p),
    .din1(g1235_n_spl_),
    .din2(g1236_n)
  );


  orX
  g_g1237_n
  (
    .dout(g1237_n),
    .din1(g1235_p_spl_),
    .din2(g1236_p)
  );


  andX
  g_g1238_p
  (
    .dout(g1238_p),
    .din1(g1223_n_spl_),
    .din2(g1237_p_spl_)
  );


  orX
  g_g1238_n
  (
    .dout(g1238_n),
    .din1(g1223_p_spl_),
    .din2(g1237_n_spl_)
  );


  andX
  g_g1239_p
  (
    .dout(g1239_p),
    .din1(g1223_p_spl_),
    .din2(g1237_n_spl_)
  );


  orX
  g_g1239_n
  (
    .dout(g1239_n),
    .din1(g1223_n_spl_),
    .din2(g1237_p_spl_)
  );


  andX
  g_g1240_p
  (
    .dout(g1240_p),
    .din1(g1238_n_spl_),
    .din2(g1239_n)
  );


  orX
  g_g1240_n
  (
    .dout(g1240_n),
    .din1(g1238_p_spl_),
    .din2(g1239_p)
  );


  andX
  g_g1241_p
  (
    .dout(g1241_p),
    .din1(g1222_n_spl_),
    .din2(g1240_p_spl_)
  );


  orX
  g_g1241_n
  (
    .dout(g1241_n),
    .din1(g1222_p_spl_),
    .din2(g1240_n_spl_)
  );


  andX
  g_g1242_p
  (
    .dout(g1242_p),
    .din1(g988_n),
    .din2(g1012_p_spl_)
  );


  orX
  g_g1242_n
  (
    .dout(g1242_n),
    .din1(g988_p_spl_),
    .din2(g1012_n)
  );


  andX
  g_g1243_p
  (
    .dout(g1243_p),
    .din1(G3_p_spl_00),
    .din2(G17_p_spl_000)
  );


  orX
  g_g1243_n
  (
    .dout(g1243_n),
    .din1(G3_n_spl_0),
    .din2(G17_n_spl_000)
  );


  andX
  g_g1244_p
  (
    .dout(g1244_p),
    .din1(G2_p_spl_00),
    .din2(G18_p_spl_000)
  );


  orX
  g_g1244_n
  (
    .dout(g1244_n),
    .din1(G2_n_spl_0),
    .din2(G18_n_spl_000)
  );


  andX
  g_g1245_p
  (
    .dout(g1245_p),
    .din1(g1243_p_spl_),
    .din2(g1244_p_spl_)
  );


  orX
  g_g1245_n
  (
    .dout(g1245_n),
    .din1(g1243_n_spl_),
    .din2(g1244_n_spl_)
  );


  andX
  g_g1246_p
  (
    .dout(g1246_p),
    .din1(g1243_n_spl_),
    .din2(g1244_n_spl_)
  );


  orX
  g_g1246_n
  (
    .dout(g1246_n),
    .din1(g1243_p_spl_),
    .din2(g1244_p_spl_)
  );


  andX
  g_g1247_p
  (
    .dout(g1247_p),
    .din1(g1245_n_spl_0),
    .din2(g1246_n)
  );


  orX
  g_g1247_n
  (
    .dout(g1247_n),
    .din1(g1245_p_spl_0),
    .din2(g1246_p)
  );


  andX
  g_g1248_p
  (
    .dout(g1248_p),
    .din1(g989_n_spl_),
    .din2(g1247_n_spl_)
  );


  orX
  g_g1248_n
  (
    .dout(g1248_n),
    .din1(g989_p_spl_0),
    .din2(g1247_p_spl_)
  );


  andX
  g_g1249_p
  (
    .dout(g1249_p),
    .din1(g989_p_spl_0),
    .din2(g1247_p_spl_)
  );


  orX
  g_g1249_n
  (
    .dout(g1249_n),
    .din1(g989_n_spl_),
    .din2(g1247_n_spl_)
  );


  andX
  g_g1250_p
  (
    .dout(g1250_p),
    .din1(g1248_n_spl_),
    .din2(g1249_n)
  );


  orX
  g_g1250_n
  (
    .dout(g1250_n),
    .din1(g1248_p_spl_),
    .din2(g1249_p)
  );


  andX
  g_g1251_p
  (
    .dout(g1251_p),
    .din1(g982_n_spl_),
    .din2(g987_n)
  );


  orX
  g_g1251_n
  (
    .dout(g1251_n),
    .din1(g982_p_spl_),
    .din2(g987_p_spl_)
  );


  andX
  g_g1252_p
  (
    .dout(g1252_p),
    .din1(ffc_19_p_spl_001),
    .din2(ffc_133_p_spl_1)
  );


  orX
  g_g1252_n
  (
    .dout(g1252_n),
    .din1(ffc_19_n_spl_01),
    .din2(ffc_133_n_spl_1)
  );


  andX
  g_g1253_p
  (
    .dout(g1253_p),
    .din1(g976_n_spl_),
    .din2(g979_n_spl_)
  );


  orX
  g_g1253_n
  (
    .dout(g1253_n),
    .din1(g976_p_spl_),
    .din2(g979_p_spl_)
  );


  andX
  g_g1254_p
  (
    .dout(g1254_p),
    .din1(ffc_17_p_spl_011),
    .din2(ffc_118_p_spl_01)
  );


  orX
  g_g1254_n
  (
    .dout(g1254_n),
    .din1(ffc_17_n_spl_10),
    .din2(ffc_118_n_spl_0)
  );


  andX
  g_g1255_p
  (
    .dout(g1255_p),
    .din1(g970_n_spl_),
    .din2(g973_n_spl_)
  );


  orX
  g_g1255_n
  (
    .dout(g1255_n),
    .din1(g970_p_spl_),
    .din2(g973_p_spl_)
  );


  andX
  g_g1256_p
  (
    .dout(g1256_p),
    .din1(ffc_15_p_spl_101),
    .din2(ffc_119_p_spl_00)
  );


  orX
  g_g1256_n
  (
    .dout(g1256_n),
    .din1(ffc_15_n_spl_101),
    .din2(ffc_119_n_spl_00)
  );


  andX
  g_g1257_p
  (
    .dout(g1257_p),
    .din1(ffc_298_p_spl_),
    .din2(g967_n_spl_)
  );


  orX
  g_g1257_n
  (
    .dout(g1257_n),
    .din1(ffc_298_n_spl_),
    .din2(g967_p_spl_)
  );


  andX
  g_g1258_p
  (
    .dout(g1258_p),
    .din1(g1165_p_spl_),
    .din2(g1166_n_spl_)
  );


  orX
  g_g1258_n
  (
    .dout(g1258_n),
    .din1(g1165_n_spl_),
    .din2(g1166_p_spl_)
  );


  andX
  g_g1259_p
  (
    .dout(g1259_p),
    .din1(g1167_n_spl_),
    .din2(g1258_n)
  );


  orX
  g_g1259_n
  (
    .dout(g1259_n),
    .din1(g1167_p_spl_),
    .din2(g1258_p)
  );


  andX
  g_g1260_p
  (
    .dout(g1260_p),
    .din1(g1257_n_spl_),
    .din2(g1259_p_spl_)
  );


  orX
  g_g1260_n
  (
    .dout(g1260_n),
    .din1(g1257_p_spl_),
    .din2(g1259_n_spl_)
  );


  andX
  g_g1261_p
  (
    .dout(g1261_p),
    .din1(g1257_p_spl_),
    .din2(g1259_n_spl_)
  );


  orX
  g_g1261_n
  (
    .dout(g1261_n),
    .din1(g1257_n_spl_),
    .din2(g1259_p_spl_)
  );


  andX
  g_g1262_p
  (
    .dout(g1262_p),
    .din1(g1260_n_spl_),
    .din2(g1261_n)
  );


  orX
  g_g1262_n
  (
    .dout(g1262_n),
    .din1(g1260_p_spl_),
    .din2(g1261_p)
  );


  andX
  g_g1263_p
  (
    .dout(g1263_p),
    .din1(g1256_n_spl_),
    .din2(g1262_p_spl_)
  );


  orX
  g_g1263_n
  (
    .dout(g1263_n),
    .din1(g1256_p_spl_),
    .din2(g1262_n_spl_)
  );


  andX
  g_g1264_p
  (
    .dout(g1264_p),
    .din1(g1256_p_spl_),
    .din2(g1262_n_spl_)
  );


  orX
  g_g1264_n
  (
    .dout(g1264_n),
    .din1(g1256_n_spl_),
    .din2(g1262_p_spl_)
  );


  andX
  g_g1265_p
  (
    .dout(g1265_p),
    .din1(g1263_n_spl_),
    .din2(g1264_n)
  );


  orX
  g_g1265_n
  (
    .dout(g1265_n),
    .din1(g1263_p_spl_),
    .din2(g1264_p)
  );


  andX
  g_g1266_p
  (
    .dout(g1266_p),
    .din1(g1255_n_spl_),
    .din2(g1265_p_spl_)
  );


  orX
  g_g1266_n
  (
    .dout(g1266_n),
    .din1(g1255_p_spl_),
    .din2(g1265_n_spl_)
  );


  andX
  g_g1267_p
  (
    .dout(g1267_p),
    .din1(g1255_p_spl_),
    .din2(g1265_n_spl_)
  );


  orX
  g_g1267_n
  (
    .dout(g1267_n),
    .din1(g1255_n_spl_),
    .din2(g1265_p_spl_)
  );


  andX
  g_g1268_p
  (
    .dout(g1268_p),
    .din1(g1266_n_spl_),
    .din2(g1267_n)
  );


  orX
  g_g1268_n
  (
    .dout(g1268_n),
    .din1(g1266_p_spl_),
    .din2(g1267_p)
  );


  andX
  g_g1269_p
  (
    .dout(g1269_p),
    .din1(g1254_n_spl_),
    .din2(g1268_p_spl_)
  );


  orX
  g_g1269_n
  (
    .dout(g1269_n),
    .din1(g1254_p_spl_),
    .din2(g1268_n_spl_)
  );


  andX
  g_g1270_p
  (
    .dout(g1270_p),
    .din1(g1254_p_spl_),
    .din2(g1268_n_spl_)
  );


  orX
  g_g1270_n
  (
    .dout(g1270_n),
    .din1(g1254_n_spl_),
    .din2(g1268_p_spl_)
  );


  andX
  g_g1271_p
  (
    .dout(g1271_p),
    .din1(g1269_n_spl_),
    .din2(g1270_n)
  );


  orX
  g_g1271_n
  (
    .dout(g1271_n),
    .din1(g1269_p_spl_),
    .din2(g1270_p)
  );


  andX
  g_g1272_p
  (
    .dout(g1272_p),
    .din1(g1253_n_spl_),
    .din2(g1271_p_spl_)
  );


  orX
  g_g1272_n
  (
    .dout(g1272_n),
    .din1(g1253_p_spl_),
    .din2(g1271_n_spl_)
  );


  andX
  g_g1273_p
  (
    .dout(g1273_p),
    .din1(g1253_p_spl_),
    .din2(g1271_n_spl_)
  );


  orX
  g_g1273_n
  (
    .dout(g1273_n),
    .din1(g1253_n_spl_),
    .din2(g1271_p_spl_)
  );


  andX
  g_g1274_p
  (
    .dout(g1274_p),
    .din1(g1272_n_spl_),
    .din2(g1273_n)
  );


  orX
  g_g1274_n
  (
    .dout(g1274_n),
    .din1(g1272_p_spl_),
    .din2(g1273_p)
  );


  andX
  g_g1275_p
  (
    .dout(g1275_p),
    .din1(g1252_n_spl_),
    .din2(g1274_p_spl_)
  );


  orX
  g_g1275_n
  (
    .dout(g1275_n),
    .din1(g1252_p_spl_),
    .din2(g1274_n_spl_)
  );


  andX
  g_g1276_p
  (
    .dout(g1276_p),
    .din1(g1252_p_spl_),
    .din2(g1274_n_spl_)
  );


  orX
  g_g1276_n
  (
    .dout(g1276_n),
    .din1(g1252_n_spl_),
    .din2(g1274_p_spl_)
  );


  andX
  g_g1277_p
  (
    .dout(g1277_p),
    .din1(g1275_n_spl_),
    .din2(g1276_n)
  );


  orX
  g_g1277_n
  (
    .dout(g1277_n),
    .din1(g1275_p_spl_),
    .din2(g1276_p)
  );


  orX
  g_g1278_n
  (
    .dout(g1278_n),
    .din1(g1251_p),
    .din2(g1277_n)
  );


  andX
  g_g1279_p
  (
    .dout(g1279_p),
    .din1(ffc_336_n_spl_),
    .din2(ffc_353_p_spl_)
  );


  orX
  g_g1279_n
  (
    .dout(g1279_n),
    .din1(ffc_336_p_spl_),
    .din2(ffc_353_n_spl_)
  );


  andX
  g_g1280_p
  (
    .dout(g1280_p),
    .din1(ffc_322_p),
    .din2(g1279_n_spl_)
  );


  orX
  g_g1280_n
  (
    .dout(g1280_n),
    .din1(ffc_322_n),
    .din2(g1279_p_spl_)
  );


  andX
  g_g1281_p
  (
    .dout(g1281_p),
    .din1(ffc_337_n_spl_),
    .din2(ffc_354_p_spl_)
  );


  orX
  g_g1281_n
  (
    .dout(g1281_n),
    .din1(ffc_337_p_spl_),
    .din2(ffc_354_n_spl_)
  );


  andX
  g_g1282_p
  (
    .dout(g1282_p),
    .din1(ffc_337_p_spl_),
    .din2(ffc_354_n_spl_)
  );


  orX
  g_g1282_n
  (
    .dout(g1282_n),
    .din1(ffc_337_n_spl_),
    .din2(ffc_354_p_spl_)
  );


  andX
  g_g1283_p
  (
    .dout(g1283_p),
    .din1(g1281_n_spl_),
    .din2(g1282_n)
  );


  orX
  g_g1283_n
  (
    .dout(g1283_n),
    .din1(g1281_p_spl_),
    .din2(g1282_p)
  );


  andX
  g_g1284_p
  (
    .dout(g1284_p),
    .din1(g1280_n_spl_),
    .din2(g1283_p_spl_)
  );


  orX
  g_g1284_n
  (
    .dout(g1284_n),
    .din1(g1280_p_spl_),
    .din2(g1283_n_spl_)
  );


  andX
  g_g1285_p
  (
    .dout(g1285_p),
    .din1(ffc_9_p_spl_001),
    .din2(ffc_190_p_spl_0)
  );


  orX
  g_g1285_n
  (
    .dout(g1285_n),
    .din1(ffc_9_n_spl_001),
    .din2(ffc_190_n_spl_0)
  );


  andX
  g_g1286_p
  (
    .dout(g1286_p),
    .din1(g1280_p_spl_),
    .din2(g1283_n_spl_)
  );


  orX
  g_g1286_n
  (
    .dout(g1286_n),
    .din1(g1280_n_spl_),
    .din2(g1283_p_spl_)
  );


  andX
  g_g1287_p
  (
    .dout(g1287_p),
    .din1(g1284_n_spl_),
    .din2(g1286_n)
  );


  orX
  g_g1287_n
  (
    .dout(g1287_n),
    .din1(g1284_p_spl_),
    .din2(g1286_p)
  );


  andX
  g_g1288_p
  (
    .dout(g1288_p),
    .din1(g1285_n_spl_),
    .din2(g1287_p_spl_)
  );


  orX
  g_g1288_n
  (
    .dout(g1288_n),
    .din1(g1285_p_spl_),
    .din2(g1287_n_spl_)
  );


  andX
  g_g1289_p
  (
    .dout(g1289_p),
    .din1(g1284_n_spl_),
    .din2(g1288_n_spl_)
  );


  orX
  g_g1289_n
  (
    .dout(g1289_n),
    .din1(g1284_p_spl_),
    .din2(g1288_p_spl_)
  );


  andX
  g_g1290_p
  (
    .dout(g1290_p),
    .din1(ffc_9_p_spl_010),
    .din2(ffc_191_p_spl_0)
  );


  orX
  g_g1290_n
  (
    .dout(g1290_n),
    .din1(ffc_9_n_spl_010),
    .din2(ffc_191_n_spl_0)
  );


  andX
  g_g1291_p
  (
    .dout(g1291_p),
    .din1(ffc_323_p),
    .din2(g1281_n_spl_)
  );


  orX
  g_g1291_n
  (
    .dout(g1291_n),
    .din1(ffc_323_n),
    .din2(g1281_p_spl_)
  );


  andX
  g_g1292_p
  (
    .dout(g1292_p),
    .din1(ffc_192_p_spl_0),
    .din2(ffc_325_p_spl_0)
  );


  orX
  g_g1292_n
  (
    .dout(g1292_n),
    .din1(ffc_192_n_spl_0),
    .din2(ffc_325_n_spl_0)
  );


  andX
  g_g1293_p
  (
    .dout(g1293_p),
    .din1(ffc_338_n_spl_),
    .din2(ffc_340_n_spl_)
  );


  orX
  g_g1293_n
  (
    .dout(g1293_n),
    .din1(ffc_338_p_spl_),
    .din2(ffc_340_p_spl_)
  );


  andX
  g_g1294_p
  (
    .dout(g1294_p),
    .din1(ffc_338_p_spl_),
    .din2(ffc_340_p_spl_)
  );


  orX
  g_g1294_n
  (
    .dout(g1294_n),
    .din1(ffc_338_n_spl_),
    .din2(ffc_340_n_spl_)
  );


  andX
  g_g1295_p
  (
    .dout(g1295_p),
    .din1(g1293_n_spl_),
    .din2(g1294_n)
  );


  orX
  g_g1295_n
  (
    .dout(g1295_n),
    .din1(g1293_p_spl_),
    .din2(g1294_p)
  );


  andX
  g_g1296_p
  (
    .dout(g1296_p),
    .din1(g1292_n_spl_),
    .din2(g1295_p_spl_)
  );


  orX
  g_g1296_n
  (
    .dout(g1296_n),
    .din1(g1292_p_spl_),
    .din2(g1295_n_spl_)
  );


  andX
  g_g1297_p
  (
    .dout(g1297_p),
    .din1(g1292_p_spl_),
    .din2(g1295_n_spl_)
  );


  orX
  g_g1297_n
  (
    .dout(g1297_n),
    .din1(g1292_n_spl_),
    .din2(g1295_p_spl_)
  );


  andX
  g_g1298_p
  (
    .dout(g1298_p),
    .din1(g1296_n_spl_),
    .din2(g1297_n)
  );


  orX
  g_g1298_n
  (
    .dout(g1298_n),
    .din1(g1296_p_spl_),
    .din2(g1297_p)
  );


  andX
  g_g1299_p
  (
    .dout(g1299_p),
    .din1(g1291_n_spl_),
    .din2(g1298_p_spl_)
  );


  orX
  g_g1299_n
  (
    .dout(g1299_n),
    .din1(g1291_p_spl_),
    .din2(g1298_n_spl_)
  );


  andX
  g_g1300_p
  (
    .dout(g1300_p),
    .din1(g1291_p_spl_),
    .din2(g1298_n_spl_)
  );


  orX
  g_g1300_n
  (
    .dout(g1300_n),
    .din1(g1291_n_spl_),
    .din2(g1298_p_spl_)
  );


  andX
  g_g1301_p
  (
    .dout(g1301_p),
    .din1(g1299_n_spl_),
    .din2(g1300_n)
  );


  orX
  g_g1301_n
  (
    .dout(g1301_n),
    .din1(g1299_p_spl_),
    .din2(g1300_p)
  );


  andX
  g_g1302_p
  (
    .dout(g1302_p),
    .din1(g1290_n_spl_),
    .din2(g1301_p_spl_)
  );


  orX
  g_g1302_n
  (
    .dout(g1302_n),
    .din1(g1290_p_spl_),
    .din2(g1301_n_spl_)
  );


  andX
  g_g1303_p
  (
    .dout(g1303_p),
    .din1(g1290_p_spl_),
    .din2(g1301_n_spl_)
  );


  orX
  g_g1303_n
  (
    .dout(g1303_n),
    .din1(g1290_n_spl_),
    .din2(g1301_p_spl_)
  );


  andX
  g_g1304_p
  (
    .dout(g1304_p),
    .din1(g1302_n_spl_),
    .din2(g1303_n)
  );


  orX
  g_g1304_n
  (
    .dout(g1304_n),
    .din1(g1302_p_spl_),
    .din2(g1303_p)
  );


  andX
  g_g1305_p
  (
    .dout(g1305_p),
    .din1(g1289_n_spl_),
    .din2(g1304_p_spl_)
  );


  orX
  g_g1305_n
  (
    .dout(g1305_n),
    .din1(g1289_p_spl_),
    .din2(g1304_n_spl_)
  );


  andX
  g_g1306_p
  (
    .dout(g1306_p),
    .din1(ffc_10_p_spl_001),
    .din2(ffc_190_p_spl_0)
  );


  orX
  g_g1306_n
  (
    .dout(g1306_n),
    .din1(ffc_10_n_spl_001),
    .din2(ffc_190_n_spl_0)
  );


  andX
  g_g1307_p
  (
    .dout(g1307_p),
    .din1(g1289_p_spl_),
    .din2(g1304_n_spl_)
  );


  orX
  g_g1307_n
  (
    .dout(g1307_n),
    .din1(g1289_n_spl_),
    .din2(g1304_p_spl_)
  );


  andX
  g_g1308_p
  (
    .dout(g1308_p),
    .din1(g1305_n_spl_),
    .din2(g1307_n)
  );


  orX
  g_g1308_n
  (
    .dout(g1308_n),
    .din1(g1305_p_spl_),
    .din2(g1307_p)
  );


  andX
  g_g1309_p
  (
    .dout(g1309_p),
    .din1(g1306_n_spl_),
    .din2(g1308_p_spl_)
  );


  orX
  g_g1309_n
  (
    .dout(g1309_n),
    .din1(g1306_p_spl_),
    .din2(g1308_n_spl_)
  );


  andX
  g_g1310_p
  (
    .dout(g1310_p),
    .din1(g1305_n_spl_),
    .din2(g1309_n_spl_)
  );


  orX
  g_g1310_n
  (
    .dout(g1310_n),
    .din1(g1305_p_spl_),
    .din2(g1309_p_spl_)
  );


  andX
  g_g1311_p
  (
    .dout(g1311_p),
    .din1(ffc_10_p_spl_001),
    .din2(ffc_191_p_spl_0)
  );


  orX
  g_g1311_n
  (
    .dout(g1311_n),
    .din1(ffc_10_n_spl_001),
    .din2(ffc_191_n_spl_0)
  );


  andX
  g_g1312_p
  (
    .dout(g1312_p),
    .din1(g1299_n_spl_),
    .din2(g1302_n_spl_)
  );


  orX
  g_g1312_n
  (
    .dout(g1312_n),
    .din1(g1299_p_spl_),
    .din2(g1302_p_spl_)
  );


  andX
  g_g1313_p
  (
    .dout(g1313_p),
    .din1(ffc_9_p_spl_010),
    .din2(ffc_192_p_spl_0)
  );


  orX
  g_g1313_n
  (
    .dout(g1313_n),
    .din1(ffc_9_n_spl_010),
    .din2(ffc_192_n_spl_0)
  );


  andX
  g_g1314_p
  (
    .dout(g1314_p),
    .din1(ffc_193_p_spl_0),
    .din2(ffc_325_p_spl_)
  );


  orX
  g_g1314_n
  (
    .dout(g1314_n),
    .din1(ffc_193_n_spl_0),
    .din2(ffc_325_n_spl_)
  );


  andX
  g_g1315_p
  (
    .dout(g1315_p),
    .din1(g1293_n_spl_),
    .din2(g1296_n_spl_)
  );


  orX
  g_g1315_n
  (
    .dout(g1315_n),
    .din1(g1293_p_spl_),
    .din2(g1296_p_spl_)
  );


  andX
  g_g1316_p
  (
    .dout(g1316_p),
    .din1(g1314_n_spl_),
    .din2(g1315_n_spl_)
  );


  orX
  g_g1316_n
  (
    .dout(g1316_n),
    .din1(g1314_p_spl_),
    .din2(g1315_p_spl_)
  );


  andX
  g_g1317_p
  (
    .dout(g1317_p),
    .din1(g1314_p_spl_),
    .din2(g1315_p_spl_)
  );


  orX
  g_g1317_n
  (
    .dout(g1317_n),
    .din1(g1314_n_spl_),
    .din2(g1315_n_spl_)
  );


  andX
  g_g1318_p
  (
    .dout(g1318_p),
    .din1(g1316_n_spl_),
    .din2(g1317_n)
  );


  orX
  g_g1318_n
  (
    .dout(g1318_n),
    .din1(g1316_p_spl_),
    .din2(g1317_p)
  );


  andX
  g_g1319_p
  (
    .dout(g1319_p),
    .din1(g1313_n_spl_),
    .din2(g1318_p_spl_)
  );


  orX
  g_g1319_n
  (
    .dout(g1319_n),
    .din1(g1313_p_spl_),
    .din2(g1318_n_spl_)
  );


  andX
  g_g1320_p
  (
    .dout(g1320_p),
    .din1(g1313_p_spl_),
    .din2(g1318_n_spl_)
  );


  orX
  g_g1320_n
  (
    .dout(g1320_n),
    .din1(g1313_n_spl_),
    .din2(g1318_p_spl_)
  );


  andX
  g_g1321_p
  (
    .dout(g1321_p),
    .din1(g1319_n_spl_),
    .din2(g1320_n)
  );


  orX
  g_g1321_n
  (
    .dout(g1321_n),
    .din1(g1319_p_spl_),
    .din2(g1320_p)
  );


  andX
  g_g1322_p
  (
    .dout(g1322_p),
    .din1(g1312_n_spl_),
    .din2(g1321_p_spl_)
  );


  orX
  g_g1322_n
  (
    .dout(g1322_n),
    .din1(g1312_p_spl_),
    .din2(g1321_n_spl_)
  );


  andX
  g_g1323_p
  (
    .dout(g1323_p),
    .din1(g1312_p_spl_),
    .din2(g1321_n_spl_)
  );


  orX
  g_g1323_n
  (
    .dout(g1323_n),
    .din1(g1312_n_spl_),
    .din2(g1321_p_spl_)
  );


  andX
  g_g1324_p
  (
    .dout(g1324_p),
    .din1(g1322_n_spl_),
    .din2(g1323_n)
  );


  orX
  g_g1324_n
  (
    .dout(g1324_n),
    .din1(g1322_p_spl_),
    .din2(g1323_p)
  );


  andX
  g_g1325_p
  (
    .dout(g1325_p),
    .din1(g1311_n_spl_),
    .din2(g1324_p_spl_)
  );


  orX
  g_g1325_n
  (
    .dout(g1325_n),
    .din1(g1311_p_spl_),
    .din2(g1324_n_spl_)
  );


  andX
  g_g1326_p
  (
    .dout(g1326_p),
    .din1(g1311_p_spl_),
    .din2(g1324_n_spl_)
  );


  orX
  g_g1326_n
  (
    .dout(g1326_n),
    .din1(g1311_n_spl_),
    .din2(g1324_p_spl_)
  );


  andX
  g_g1327_p
  (
    .dout(g1327_p),
    .din1(g1325_n_spl_),
    .din2(g1326_n)
  );


  orX
  g_g1327_n
  (
    .dout(g1327_n),
    .din1(g1325_p_spl_),
    .din2(g1326_p)
  );


  andX
  g_g1328_p
  (
    .dout(g1328_p),
    .din1(g1310_n_spl_),
    .din2(g1327_p_spl_)
  );


  orX
  g_g1328_n
  (
    .dout(g1328_n),
    .din1(g1310_p_spl_),
    .din2(g1327_n_spl_)
  );


  andX
  g_g1329_p
  (
    .dout(g1329_p),
    .din1(ffc_333_n_spl_),
    .din2(ffc_350_p_spl_)
  );


  orX
  g_g1329_n
  (
    .dout(g1329_n),
    .din1(ffc_333_p_spl_),
    .din2(ffc_350_n_spl_)
  );


  andX
  g_g1330_p
  (
    .dout(g1330_p),
    .din1(ffc_319_p),
    .din2(g1329_n_spl_)
  );


  orX
  g_g1330_n
  (
    .dout(g1330_n),
    .din1(ffc_319_n),
    .din2(g1329_p_spl_)
  );


  andX
  g_g1331_p
  (
    .dout(g1331_p),
    .din1(ffc_334_n_spl_),
    .din2(ffc_351_p_spl_)
  );


  orX
  g_g1331_n
  (
    .dout(g1331_n),
    .din1(ffc_334_p_spl_),
    .din2(ffc_351_n_spl_)
  );


  andX
  g_g1332_p
  (
    .dout(g1332_p),
    .din1(ffc_334_p_spl_),
    .din2(ffc_351_n_spl_)
  );


  orX
  g_g1332_n
  (
    .dout(g1332_n),
    .din1(ffc_334_n_spl_),
    .din2(ffc_351_p_spl_)
  );


  andX
  g_g1333_p
  (
    .dout(g1333_p),
    .din1(g1331_n_spl_),
    .din2(g1332_n)
  );


  orX
  g_g1333_n
  (
    .dout(g1333_n),
    .din1(g1331_p_spl_),
    .din2(g1332_p)
  );


  andX
  g_g1334_p
  (
    .dout(g1334_p),
    .din1(g1330_n_spl_),
    .din2(g1333_p_spl_)
  );


  orX
  g_g1334_n
  (
    .dout(g1334_n),
    .din1(g1330_p_spl_),
    .din2(g1333_n_spl_)
  );


  andX
  g_g1335_p
  (
    .dout(g1335_p),
    .din1(ffc_9_p_spl_011),
    .din2(ffc_187_p_spl_00)
  );


  orX
  g_g1335_n
  (
    .dout(g1335_n),
    .din1(ffc_9_n_spl_011),
    .din2(ffc_187_n_spl_0)
  );


  andX
  g_g1336_p
  (
    .dout(g1336_p),
    .din1(g1330_p_spl_),
    .din2(g1333_n_spl_)
  );


  orX
  g_g1336_n
  (
    .dout(g1336_n),
    .din1(g1330_n_spl_),
    .din2(g1333_p_spl_)
  );


  andX
  g_g1337_p
  (
    .dout(g1337_p),
    .din1(g1334_n_spl_),
    .din2(g1336_n)
  );


  orX
  g_g1337_n
  (
    .dout(g1337_n),
    .din1(g1334_p_spl_),
    .din2(g1336_p)
  );


  andX
  g_g1338_p
  (
    .dout(g1338_p),
    .din1(g1335_n_spl_),
    .din2(g1337_p_spl_)
  );


  orX
  g_g1338_n
  (
    .dout(g1338_n),
    .din1(g1335_p_spl_),
    .din2(g1337_n_spl_)
  );


  andX
  g_g1339_p
  (
    .dout(g1339_p),
    .din1(g1334_n_spl_),
    .din2(g1338_n_spl_)
  );


  orX
  g_g1339_n
  (
    .dout(g1339_n),
    .din1(g1334_p_spl_),
    .din2(g1338_p_spl_)
  );


  andX
  g_g1340_p
  (
    .dout(g1340_p),
    .din1(ffc_9_p_spl_011),
    .din2(ffc_188_p_spl_0)
  );


  orX
  g_g1340_n
  (
    .dout(g1340_n),
    .din1(ffc_9_n_spl_011),
    .din2(ffc_188_n_spl_0)
  );


  andX
  g_g1341_p
  (
    .dout(g1341_p),
    .din1(ffc_320_p),
    .din2(g1331_n_spl_)
  );


  orX
  g_g1341_n
  (
    .dout(g1341_n),
    .din1(ffc_320_n),
    .din2(g1331_p_spl_)
  );


  andX
  g_g1342_p
  (
    .dout(g1342_p),
    .din1(ffc_335_n_spl_),
    .din2(ffc_352_p_spl_)
  );


  orX
  g_g1342_n
  (
    .dout(g1342_n),
    .din1(ffc_335_p_spl_),
    .din2(ffc_352_n_spl_)
  );


  andX
  g_g1343_p
  (
    .dout(g1343_p),
    .din1(ffc_335_p_spl_),
    .din2(ffc_352_n_spl_)
  );


  orX
  g_g1343_n
  (
    .dout(g1343_n),
    .din1(ffc_335_n_spl_),
    .din2(ffc_352_p_spl_)
  );


  andX
  g_g1344_p
  (
    .dout(g1344_p),
    .din1(g1342_n_spl_),
    .din2(g1343_n)
  );


  orX
  g_g1344_n
  (
    .dout(g1344_n),
    .din1(g1342_p_spl_),
    .din2(g1343_p)
  );


  andX
  g_g1345_p
  (
    .dout(g1345_p),
    .din1(g1341_n_spl_),
    .din2(g1344_p_spl_)
  );


  orX
  g_g1345_n
  (
    .dout(g1345_n),
    .din1(g1341_p_spl_),
    .din2(g1344_n_spl_)
  );


  andX
  g_g1346_p
  (
    .dout(g1346_p),
    .din1(g1341_p_spl_),
    .din2(g1344_n_spl_)
  );


  orX
  g_g1346_n
  (
    .dout(g1346_n),
    .din1(g1341_n_spl_),
    .din2(g1344_p_spl_)
  );


  andX
  g_g1347_p
  (
    .dout(g1347_p),
    .din1(g1345_n_spl_),
    .din2(g1346_n)
  );


  orX
  g_g1347_n
  (
    .dout(g1347_n),
    .din1(g1345_p_spl_),
    .din2(g1346_p)
  );


  andX
  g_g1348_p
  (
    .dout(g1348_p),
    .din1(g1340_n_spl_),
    .din2(g1347_p_spl_)
  );


  orX
  g_g1348_n
  (
    .dout(g1348_n),
    .din1(g1340_p_spl_),
    .din2(g1347_n_spl_)
  );


  andX
  g_g1349_p
  (
    .dout(g1349_p),
    .din1(g1340_p_spl_),
    .din2(g1347_n_spl_)
  );


  orX
  g_g1349_n
  (
    .dout(g1349_n),
    .din1(g1340_n_spl_),
    .din2(g1347_p_spl_)
  );


  andX
  g_g1350_p
  (
    .dout(g1350_p),
    .din1(g1348_n_spl_),
    .din2(g1349_n)
  );


  orX
  g_g1350_n
  (
    .dout(g1350_n),
    .din1(g1348_p_spl_),
    .din2(g1349_p)
  );


  andX
  g_g1351_p
  (
    .dout(g1351_p),
    .din1(g1339_n_spl_),
    .din2(g1350_p_spl_)
  );


  orX
  g_g1351_n
  (
    .dout(g1351_n),
    .din1(g1339_p_spl_),
    .din2(g1350_n_spl_)
  );


  andX
  g_g1352_p
  (
    .dout(g1352_p),
    .din1(ffc_10_p_spl_010),
    .din2(ffc_187_p_spl_00)
  );


  orX
  g_g1352_n
  (
    .dout(g1352_n),
    .din1(ffc_10_n_spl_010),
    .din2(ffc_187_n_spl_0)
  );


  andX
  g_g1353_p
  (
    .dout(g1353_p),
    .din1(g1339_p_spl_),
    .din2(g1350_n_spl_)
  );


  orX
  g_g1353_n
  (
    .dout(g1353_n),
    .din1(g1339_n_spl_),
    .din2(g1350_p_spl_)
  );


  andX
  g_g1354_p
  (
    .dout(g1354_p),
    .din1(g1351_n_spl_),
    .din2(g1353_n)
  );


  orX
  g_g1354_n
  (
    .dout(g1354_n),
    .din1(g1351_p_spl_),
    .din2(g1353_p)
  );


  andX
  g_g1355_p
  (
    .dout(g1355_p),
    .din1(g1352_n_spl_),
    .din2(g1354_p_spl_)
  );


  orX
  g_g1355_n
  (
    .dout(g1355_n),
    .din1(g1352_p_spl_),
    .din2(g1354_n_spl_)
  );


  andX
  g_g1356_p
  (
    .dout(g1356_p),
    .din1(g1351_n_spl_),
    .din2(g1355_n_spl_)
  );


  orX
  g_g1356_n
  (
    .dout(g1356_n),
    .din1(g1351_p_spl_),
    .din2(g1355_p_spl_)
  );


  andX
  g_g1357_p
  (
    .dout(g1357_p),
    .din1(ffc_10_p_spl_010),
    .din2(ffc_188_p_spl_0)
  );


  orX
  g_g1357_n
  (
    .dout(g1357_n),
    .din1(ffc_10_n_spl_010),
    .din2(ffc_188_n_spl_0)
  );


  andX
  g_g1358_p
  (
    .dout(g1358_p),
    .din1(g1345_n_spl_),
    .din2(g1348_n_spl_)
  );


  orX
  g_g1358_n
  (
    .dout(g1358_n),
    .din1(g1345_p_spl_),
    .din2(g1348_p_spl_)
  );


  andX
  g_g1359_p
  (
    .dout(g1359_p),
    .din1(ffc_9_p_spl_100),
    .din2(ffc_189_p_spl_0)
  );


  orX
  g_g1359_n
  (
    .dout(g1359_n),
    .din1(ffc_9_n_spl_100),
    .din2(ffc_189_n_spl_0)
  );


  andX
  g_g1360_p
  (
    .dout(g1360_p),
    .din1(ffc_321_p),
    .din2(g1342_n_spl_)
  );


  orX
  g_g1360_n
  (
    .dout(g1360_n),
    .din1(ffc_321_n),
    .din2(g1342_p_spl_)
  );


  andX
  g_g1361_p
  (
    .dout(g1361_p),
    .din1(ffc_336_p_spl_),
    .din2(ffc_353_n_spl_)
  );


  orX
  g_g1361_n
  (
    .dout(g1361_n),
    .din1(ffc_336_n_spl_),
    .din2(ffc_353_p_spl_)
  );


  andX
  g_g1362_p
  (
    .dout(g1362_p),
    .din1(g1279_n_spl_),
    .din2(g1361_n)
  );


  orX
  g_g1362_n
  (
    .dout(g1362_n),
    .din1(g1279_p_spl_),
    .din2(g1361_p)
  );


  andX
  g_g1363_p
  (
    .dout(g1363_p),
    .din1(g1360_n_spl_),
    .din2(g1362_p_spl_)
  );


  orX
  g_g1363_n
  (
    .dout(g1363_n),
    .din1(g1360_p_spl_),
    .din2(g1362_n_spl_)
  );


  andX
  g_g1364_p
  (
    .dout(g1364_p),
    .din1(g1360_p_spl_),
    .din2(g1362_n_spl_)
  );


  orX
  g_g1364_n
  (
    .dout(g1364_n),
    .din1(g1360_n_spl_),
    .din2(g1362_p_spl_)
  );


  andX
  g_g1365_p
  (
    .dout(g1365_p),
    .din1(g1363_n_spl_),
    .din2(g1364_n)
  );


  orX
  g_g1365_n
  (
    .dout(g1365_n),
    .din1(g1363_p_spl_),
    .din2(g1364_p)
  );


  andX
  g_g1366_p
  (
    .dout(g1366_p),
    .din1(g1359_n_spl_),
    .din2(g1365_p_spl_)
  );


  orX
  g_g1366_n
  (
    .dout(g1366_n),
    .din1(g1359_p_spl_),
    .din2(g1365_n_spl_)
  );


  andX
  g_g1367_p
  (
    .dout(g1367_p),
    .din1(g1359_p_spl_),
    .din2(g1365_n_spl_)
  );


  orX
  g_g1367_n
  (
    .dout(g1367_n),
    .din1(g1359_n_spl_),
    .din2(g1365_p_spl_)
  );


  andX
  g_g1368_p
  (
    .dout(g1368_p),
    .din1(g1366_n_spl_),
    .din2(g1367_n)
  );


  orX
  g_g1368_n
  (
    .dout(g1368_n),
    .din1(g1366_p_spl_),
    .din2(g1367_p)
  );


  andX
  g_g1369_p
  (
    .dout(g1369_p),
    .din1(g1358_n_spl_),
    .din2(g1368_p_spl_)
  );


  orX
  g_g1369_n
  (
    .dout(g1369_n),
    .din1(g1358_p_spl_),
    .din2(g1368_n_spl_)
  );


  andX
  g_g1370_p
  (
    .dout(g1370_p),
    .din1(g1358_p_spl_),
    .din2(g1368_n_spl_)
  );


  orX
  g_g1370_n
  (
    .dout(g1370_n),
    .din1(g1358_n_spl_),
    .din2(g1368_p_spl_)
  );


  andX
  g_g1371_p
  (
    .dout(g1371_p),
    .din1(g1369_n_spl_),
    .din2(g1370_n)
  );


  orX
  g_g1371_n
  (
    .dout(g1371_n),
    .din1(g1369_p_spl_),
    .din2(g1370_p)
  );


  andX
  g_g1372_p
  (
    .dout(g1372_p),
    .din1(g1357_n_spl_),
    .din2(g1371_p_spl_)
  );


  orX
  g_g1372_n
  (
    .dout(g1372_n),
    .din1(g1357_p_spl_),
    .din2(g1371_n_spl_)
  );


  andX
  g_g1373_p
  (
    .dout(g1373_p),
    .din1(g1357_p_spl_),
    .din2(g1371_n_spl_)
  );


  orX
  g_g1373_n
  (
    .dout(g1373_n),
    .din1(g1357_n_spl_),
    .din2(g1371_p_spl_)
  );


  andX
  g_g1374_p
  (
    .dout(g1374_p),
    .din1(g1372_n_spl_),
    .din2(g1373_n)
  );


  orX
  g_g1374_n
  (
    .dout(g1374_n),
    .din1(g1372_p_spl_),
    .din2(g1373_p)
  );


  andX
  g_g1375_p
  (
    .dout(g1375_p),
    .din1(g1356_n_spl_),
    .din2(g1374_p_spl_)
  );


  orX
  g_g1375_n
  (
    .dout(g1375_n),
    .din1(g1356_p_spl_),
    .din2(g1374_n_spl_)
  );


  andX
  g_g1376_p
  (
    .dout(g1376_p),
    .din1(ffc_11_p_spl_000),
    .din2(ffc_187_p_spl_0)
  );


  orX
  g_g1376_n
  (
    .dout(g1376_n),
    .din1(ffc_11_n_spl_000),
    .din2(ffc_187_n_spl_1)
  );


  andX
  g_g1377_p
  (
    .dout(g1377_p),
    .din1(g1356_p_spl_),
    .din2(g1374_n_spl_)
  );


  orX
  g_g1377_n
  (
    .dout(g1377_n),
    .din1(g1356_n_spl_),
    .din2(g1374_p_spl_)
  );


  andX
  g_g1378_p
  (
    .dout(g1378_p),
    .din1(g1375_n_spl_),
    .din2(g1377_n)
  );


  orX
  g_g1378_n
  (
    .dout(g1378_n),
    .din1(g1375_p_spl_),
    .din2(g1377_p)
  );


  andX
  g_g1379_p
  (
    .dout(g1379_p),
    .din1(g1376_n_spl_),
    .din2(g1378_p_spl_)
  );


  orX
  g_g1379_n
  (
    .dout(g1379_n),
    .din1(g1376_p_spl_),
    .din2(g1378_n_spl_)
  );


  andX
  g_g1380_p
  (
    .dout(g1380_p),
    .din1(g1375_n_spl_),
    .din2(g1379_n_spl_)
  );


  orX
  g_g1380_n
  (
    .dout(g1380_n),
    .din1(g1375_p_spl_),
    .din2(g1379_p_spl_)
  );


  andX
  g_g1381_p
  (
    .dout(g1381_p),
    .din1(ffc_11_p_spl_001),
    .din2(ffc_188_p_spl_1)
  );


  orX
  g_g1381_n
  (
    .dout(g1381_n),
    .din1(ffc_11_n_spl_001),
    .din2(ffc_188_n_spl_1)
  );


  andX
  g_g1382_p
  (
    .dout(g1382_p),
    .din1(g1369_n_spl_),
    .din2(g1372_n_spl_)
  );


  orX
  g_g1382_n
  (
    .dout(g1382_n),
    .din1(g1369_p_spl_),
    .din2(g1372_p_spl_)
  );


  andX
  g_g1383_p
  (
    .dout(g1383_p),
    .din1(ffc_10_p_spl_011),
    .din2(ffc_189_p_spl_0)
  );


  orX
  g_g1383_n
  (
    .dout(g1383_n),
    .din1(ffc_10_n_spl_011),
    .din2(ffc_189_n_spl_0)
  );


  andX
  g_g1384_p
  (
    .dout(g1384_p),
    .din1(g1363_n_spl_),
    .din2(g1366_n_spl_)
  );


  orX
  g_g1384_n
  (
    .dout(g1384_n),
    .din1(g1363_p_spl_),
    .din2(g1366_p_spl_)
  );


  andX
  g_g1385_p
  (
    .dout(g1385_p),
    .din1(g1285_p_spl_),
    .din2(g1287_n_spl_)
  );


  orX
  g_g1385_n
  (
    .dout(g1385_n),
    .din1(g1285_n_spl_),
    .din2(g1287_p_spl_)
  );


  andX
  g_g1386_p
  (
    .dout(g1386_p),
    .din1(g1288_n_spl_),
    .din2(g1385_n)
  );


  orX
  g_g1386_n
  (
    .dout(g1386_n),
    .din1(g1288_p_spl_),
    .din2(g1385_p)
  );


  andX
  g_g1387_p
  (
    .dout(g1387_p),
    .din1(g1384_n_spl_),
    .din2(g1386_p_spl_)
  );


  orX
  g_g1387_n
  (
    .dout(g1387_n),
    .din1(g1384_p_spl_),
    .din2(g1386_n_spl_)
  );


  andX
  g_g1388_p
  (
    .dout(g1388_p),
    .din1(g1384_p_spl_),
    .din2(g1386_n_spl_)
  );


  orX
  g_g1388_n
  (
    .dout(g1388_n),
    .din1(g1384_n_spl_),
    .din2(g1386_p_spl_)
  );


  andX
  g_g1389_p
  (
    .dout(g1389_p),
    .din1(g1387_n_spl_),
    .din2(g1388_n)
  );


  orX
  g_g1389_n
  (
    .dout(g1389_n),
    .din1(g1387_p_spl_),
    .din2(g1388_p)
  );


  andX
  g_g1390_p
  (
    .dout(g1390_p),
    .din1(g1383_n_spl_),
    .din2(g1389_p_spl_)
  );


  orX
  g_g1390_n
  (
    .dout(g1390_n),
    .din1(g1383_p_spl_),
    .din2(g1389_n_spl_)
  );


  andX
  g_g1391_p
  (
    .dout(g1391_p),
    .din1(g1383_p_spl_),
    .din2(g1389_n_spl_)
  );


  orX
  g_g1391_n
  (
    .dout(g1391_n),
    .din1(g1383_n_spl_),
    .din2(g1389_p_spl_)
  );


  andX
  g_g1392_p
  (
    .dout(g1392_p),
    .din1(g1390_n_spl_),
    .din2(g1391_n)
  );


  orX
  g_g1392_n
  (
    .dout(g1392_n),
    .din1(g1390_p_spl_),
    .din2(g1391_p)
  );


  andX
  g_g1393_p
  (
    .dout(g1393_p),
    .din1(g1382_n_spl_),
    .din2(g1392_p_spl_)
  );


  orX
  g_g1393_n
  (
    .dout(g1393_n),
    .din1(g1382_p_spl_),
    .din2(g1392_n_spl_)
  );


  andX
  g_g1394_p
  (
    .dout(g1394_p),
    .din1(g1382_p_spl_),
    .din2(g1392_n_spl_)
  );


  orX
  g_g1394_n
  (
    .dout(g1394_n),
    .din1(g1382_n_spl_),
    .din2(g1392_p_spl_)
  );


  andX
  g_g1395_p
  (
    .dout(g1395_p),
    .din1(g1393_n_spl_),
    .din2(g1394_n)
  );


  orX
  g_g1395_n
  (
    .dout(g1395_n),
    .din1(g1393_p_spl_),
    .din2(g1394_p)
  );


  andX
  g_g1396_p
  (
    .dout(g1396_p),
    .din1(g1381_n_spl_),
    .din2(g1395_p_spl_)
  );


  orX
  g_g1396_n
  (
    .dout(g1396_n),
    .din1(g1381_p_spl_),
    .din2(g1395_n_spl_)
  );


  andX
  g_g1397_p
  (
    .dout(g1397_p),
    .din1(g1381_p_spl_),
    .din2(g1395_n_spl_)
  );


  orX
  g_g1397_n
  (
    .dout(g1397_n),
    .din1(g1381_n_spl_),
    .din2(g1395_p_spl_)
  );


  andX
  g_g1398_p
  (
    .dout(g1398_p),
    .din1(g1396_n_spl_),
    .din2(g1397_n)
  );


  orX
  g_g1398_n
  (
    .dout(g1398_n),
    .din1(g1396_p_spl_),
    .din2(g1397_p)
  );


  andX
  g_g1399_p
  (
    .dout(g1399_p),
    .din1(g1380_n_spl_),
    .din2(g1398_p_spl_)
  );


  orX
  g_g1399_n
  (
    .dout(g1399_n),
    .din1(g1380_p_spl_),
    .din2(g1398_n_spl_)
  );


  andX
  g_g1400_p
  (
    .dout(g1400_p),
    .din1(g1016_n),
    .din2(g1250_p_spl_)
  );


  orX
  g_g1400_n
  (
    .dout(g1400_n),
    .din1(g1016_p_spl_),
    .din2(g1250_n)
  );


  orX
  g_g1401_n
  (
    .dout(g1401_n),
    .din1(ffc_21_n_spl_00),
    .din2(ffc_135_n_spl_1)
  );


  orX
  g_g1402_n
  (
    .dout(g1402_n),
    .din1(ffc_12_n_spl_000),
    .din2(ffc_207_n_spl_1)
  );


  orX
  g_g1403_n
  (
    .dout(g1403_n),
    .din1(G1_n_spl_),
    .din2(G20_n_spl_000)
  );


  orX
  g_g1404_n
  (
    .dout(g1404_n),
    .din1(ffc_29_n_spl_11),
    .din2(ffc_70_n_spl_)
  );


  orX
  g_g1405_n
  (
    .dout(g1405_n),
    .din1(g935_n),
    .din2(g945_p)
  );


  andX
  g_g1406_p
  (
    .dout(g1406_p),
    .din1(g946_n_spl_),
    .din2(g1405_n)
  );


  andX
  g_g1407_p
  (
    .dout(g1407_p),
    .din1(g1404_n_spl_),
    .din2(g1406_p_spl_)
  );


  orX
  g_g1408_n
  (
    .dout(g1408_n),
    .din1(g1404_n_spl_),
    .din2(g1406_p_spl_)
  );


  orX
  g_g1409_n
  (
    .dout(g1409_n),
    .din1(ffc_25_n_spl_11),
    .din2(ffc_73_n_spl_)
  );


  orX
  g_g1410_n
  (
    .dout(g1410_n),
    .din1(g923_n),
    .din2(g933_p)
  );


  andX
  g_g1411_p
  (
    .dout(g1411_p),
    .din1(g934_n_spl_),
    .din2(g1410_n)
  );


  andX
  g_g1412_p
  (
    .dout(g1412_p),
    .din1(g1409_n_spl_),
    .din2(g1411_p_spl_)
  );


  orX
  g_g1413_n
  (
    .dout(g1413_n),
    .din1(g1409_n_spl_),
    .din2(g1411_p_spl_)
  );


  orX
  g_g1414_n
  (
    .dout(g1414_n),
    .din1(ffc_76_n_spl_),
    .din2(ffc_214_n_spl_11)
  );


  orX
  g_g1415_n
  (
    .dout(g1415_n),
    .din1(g920_n),
    .din2(g921_n)
  );


  andX
  g_g1416_p
  (
    .dout(g1416_p),
    .din1(g922_n_spl_),
    .din2(g1415_n)
  );


  andX
  g_g1417_p
  (
    .dout(g1417_p),
    .din1(g1414_n_spl_),
    .din2(g1416_p_spl_)
  );


  orX
  g_g1418_n
  (
    .dout(g1418_n),
    .din1(g1414_n_spl_),
    .din2(g1416_p_spl_)
  );


  orX
  g_g1419_n
  (
    .dout(g1419_n),
    .din1(g928_p_spl_),
    .din2(g931_p_spl_)
  );


  orX
  g_g1420_n
  (
    .dout(g1420_n),
    .din1(g916_n),
    .din2(g918_p)
  );


  andX
  g_g1421_p
  (
    .dout(g1421_p),
    .din1(g919_n_spl_),
    .din2(g1420_n)
  );


  andX
  g_g1422_p
  (
    .dout(g1422_p),
    .din1(g1419_n_spl_),
    .din2(g1421_p_spl_)
  );


  orX
  g_g1423_n
  (
    .dout(g1423_n),
    .din1(g1419_n_spl_),
    .din2(g1421_p_spl_)
  );


  orX
  g_g1424_n
  (
    .dout(g1424_n),
    .din1(g940_p_spl_),
    .din2(g943_p_spl_)
  );


  orX
  g_g1425_n
  (
    .dout(g1425_n),
    .din1(g912_n),
    .din2(g914_p)
  );


  andX
  g_g1426_p
  (
    .dout(g1426_p),
    .din1(g915_n_spl_),
    .din2(g1425_n)
  );


  andX
  g_g1427_p
  (
    .dout(g1427_p),
    .din1(g1424_n_spl_),
    .din2(g1426_p_spl_)
  );


  orX
  g_g1428_n
  (
    .dout(g1428_n),
    .din1(g1424_n_spl_),
    .din2(g1426_p_spl_)
  );


  orX
  g_g1429_n
  (
    .dout(g1429_n),
    .din1(g952_p_spl_),
    .din2(g955_p_spl_)
  );


  orX
  g_g1430_n
  (
    .dout(g1430_n),
    .din1(g908_n),
    .din2(g910_p)
  );


  andX
  g_g1431_p
  (
    .dout(g1431_p),
    .din1(g911_n_spl_),
    .din2(g1430_n)
  );


  andX
  g_g1432_p
  (
    .dout(g1432_p),
    .din1(g1429_n_spl_),
    .din2(g1431_p_spl_)
  );


  orX
  g_g1433_n
  (
    .dout(g1433_n),
    .din1(g1429_n_spl_),
    .din2(g1431_p_spl_)
  );


  andX
  g_g1434_p
  (
    .dout(g1434_p),
    .din1(g1013_n_spl_),
    .din2(g1015_p_spl_)
  );


  andX
  g_g1435_p
  (
    .dout(g1435_p),
    .din1(ffc_21_p_spl_00),
    .din2(ffc_120_p_spl_1)
  );


  orX
  g_g1435_n
  (
    .dout(g1435_n),
    .din1(ffc_21_n_spl_00),
    .din2(ffc_120_n_spl_1)
  );


  andX
  g_g1436_p
  (
    .dout(g1436_p),
    .din1(g1222_p_spl_),
    .din2(g1240_n_spl_)
  );


  orX
  g_g1436_n
  (
    .dout(g1436_n),
    .din1(g1222_n_spl_),
    .din2(g1240_p_spl_)
  );


  andX
  g_g1437_p
  (
    .dout(g1437_p),
    .din1(g1241_n_spl_),
    .din2(g1436_n)
  );


  orX
  g_g1437_n
  (
    .dout(g1437_n),
    .din1(g1241_p),
    .din2(g1436_p)
  );


  orX
  g_g1438_n
  (
    .dout(g1438_n),
    .din1(g1435_p),
    .din2(g1437_n)
  );


  andX
  g_g1439_p
  (
    .dout(g1439_p),
    .din1(ffc_19_p_spl_01),
    .din2(ffc_123_p_spl_1)
  );


  orX
  g_g1439_n
  (
    .dout(g1439_n),
    .din1(ffc_19_n_spl_10),
    .din2(ffc_123_n_spl_1)
  );


  andX
  g_g1440_p
  (
    .dout(g1440_p),
    .din1(g1145_p_spl_),
    .din2(g1163_n_spl_)
  );


  orX
  g_g1440_n
  (
    .dout(g1440_n),
    .din1(g1145_n_spl_),
    .din2(g1163_p_spl_)
  );


  andX
  g_g1441_p
  (
    .dout(g1441_p),
    .din1(g1164_n_spl_),
    .din2(g1440_n)
  );


  orX
  g_g1441_n
  (
    .dout(g1441_n),
    .din1(g1164_p),
    .din2(g1440_p)
  );


  orX
  g_g1442_n
  (
    .dout(g1442_n),
    .din1(g1439_p),
    .din2(g1441_n)
  );


  andX
  g_g1443_p
  (
    .dout(g1443_p),
    .din1(ffc_17_p_spl_100),
    .din2(ffc_126_p_spl_1)
  );


  orX
  g_g1443_n
  (
    .dout(g1443_n),
    .din1(ffc_17_n_spl_10),
    .din2(ffc_126_n_spl_)
  );


  andX
  g_g1444_p
  (
    .dout(g1444_p),
    .din1(g1088_p_spl_),
    .din2(g1106_n_spl_)
  );


  orX
  g_g1444_n
  (
    .dout(g1444_n),
    .din1(g1088_n_spl_),
    .din2(g1106_p_spl_)
  );


  andX
  g_g1445_p
  (
    .dout(g1445_p),
    .din1(g1107_n_spl_),
    .din2(g1444_n)
  );


  orX
  g_g1445_n
  (
    .dout(g1445_n),
    .din1(g1107_p),
    .din2(g1444_p)
  );


  orX
  g_g1446_n
  (
    .dout(g1446_n),
    .din1(g1443_p),
    .din2(g1445_n)
  );


  andX
  g_g1447_p
  (
    .dout(g1447_p),
    .din1(ffc_15_p_spl_110),
    .din2(ffc_129_p_spl_1)
  );


  orX
  g_g1447_n
  (
    .dout(g1447_n),
    .din1(ffc_15_n_spl_11),
    .din2(ffc_129_n_spl_)
  );


  andX
  g_g1448_p
  (
    .dout(g1448_p),
    .din1(g1043_p_spl_),
    .din2(g1052_n_spl_)
  );


  orX
  g_g1448_n
  (
    .dout(g1448_n),
    .din1(g1043_n_spl_),
    .din2(g1052_p_spl_)
  );


  andX
  g_g1449_p
  (
    .dout(g1449_p),
    .din1(g1053_n_spl_),
    .din2(g1448_n)
  );


  orX
  g_g1449_n
  (
    .dout(g1449_n),
    .din1(g1053_p),
    .din2(g1448_p)
  );


  orX
  g_g1450_n
  (
    .dout(g1450_n),
    .din1(g1447_p),
    .din2(g1449_n)
  );


  andX
  g_g1451_p
  (
    .dout(g1451_p),
    .din1(ffc_131_p_spl_1),
    .din2(ffc_287_p_spl_111)
  );


  orX
  g_g1451_n
  (
    .dout(g1451_n),
    .din1(ffc_131_n_spl_),
    .din2(ffc_287_n_spl_111)
  );


  andX
  g_g1452_p
  (
    .dout(g1452_p),
    .din1(g1047_n_spl_),
    .din2(g1050_n_spl_)
  );


  orX
  g_g1452_n
  (
    .dout(g1452_n),
    .din1(g1047_p_spl_),
    .din2(g1050_p_spl_)
  );


  orX
  g_g1453_n
  (
    .dout(g1453_n),
    .din1(g1451_p),
    .din2(g1452_p)
  );


  orX
  g_g1454_n
  (
    .dout(g1454_n),
    .din1(ffc_21_n_spl_0),
    .din2(ffc_133_n_spl_1)
  );


  andX
  g_g1455_p
  (
    .dout(g1455_p),
    .din1(g1272_n_spl_),
    .din2(g1275_n_spl_)
  );


  orX
  g_g1455_n
  (
    .dout(g1455_n),
    .din1(g1272_p_spl_),
    .din2(g1275_p_spl_)
  );


  andX
  g_g1456_p
  (
    .dout(g1456_p),
    .din1(ffc_19_p_spl_01),
    .din2(ffc_118_p_spl_01)
  );


  orX
  g_g1456_n
  (
    .dout(g1456_n),
    .din1(ffc_19_n_spl_10),
    .din2(ffc_118_n_spl_1)
  );


  andX
  g_g1457_p
  (
    .dout(g1457_p),
    .din1(g1266_n_spl_),
    .din2(g1269_n_spl_)
  );


  orX
  g_g1457_n
  (
    .dout(g1457_n),
    .din1(g1266_p_spl_),
    .din2(g1269_p_spl_)
  );


  andX
  g_g1458_p
  (
    .dout(g1458_p),
    .din1(ffc_17_p_spl_100),
    .din2(ffc_119_p_spl_01)
  );


  orX
  g_g1458_n
  (
    .dout(g1458_n),
    .din1(ffc_17_n_spl_11),
    .din2(ffc_119_n_spl_0)
  );


  andX
  g_g1459_p
  (
    .dout(g1459_p),
    .din1(g1260_n_spl_),
    .din2(g1263_n_spl_)
  );


  orX
  g_g1459_n
  (
    .dout(g1459_n),
    .din1(g1260_p_spl_),
    .din2(g1263_p_spl_)
  );


  andX
  g_g1460_p
  (
    .dout(g1460_p),
    .din1(g1175_p_spl_),
    .din2(g1177_n_spl_)
  );


  orX
  g_g1460_n
  (
    .dout(g1460_n),
    .din1(g1175_n_spl_),
    .din2(g1177_p_spl_)
  );


  andX
  g_g1461_p
  (
    .dout(g1461_p),
    .din1(g1178_n_spl_),
    .din2(g1460_n)
  );


  orX
  g_g1461_n
  (
    .dout(g1461_n),
    .din1(g1178_p_spl_),
    .din2(g1460_p)
  );


  andX
  g_g1462_p
  (
    .dout(g1462_p),
    .din1(g1459_n_spl_),
    .din2(g1461_p_spl_)
  );


  orX
  g_g1462_n
  (
    .dout(g1462_n),
    .din1(g1459_p_spl_),
    .din2(g1461_n_spl_)
  );


  andX
  g_g1463_p
  (
    .dout(g1463_p),
    .din1(g1459_p_spl_),
    .din2(g1461_n_spl_)
  );


  orX
  g_g1463_n
  (
    .dout(g1463_n),
    .din1(g1459_n_spl_),
    .din2(g1461_p_spl_)
  );


  andX
  g_g1464_p
  (
    .dout(g1464_p),
    .din1(g1462_n_spl_),
    .din2(g1463_n)
  );


  orX
  g_g1464_n
  (
    .dout(g1464_n),
    .din1(g1462_p_spl_),
    .din2(g1463_p)
  );


  andX
  g_g1465_p
  (
    .dout(g1465_p),
    .din1(g1458_n_spl_),
    .din2(g1464_p_spl_)
  );


  orX
  g_g1465_n
  (
    .dout(g1465_n),
    .din1(g1458_p_spl_),
    .din2(g1464_n_spl_)
  );


  andX
  g_g1466_p
  (
    .dout(g1466_p),
    .din1(g1458_p_spl_),
    .din2(g1464_n_spl_)
  );


  orX
  g_g1466_n
  (
    .dout(g1466_n),
    .din1(g1458_n_spl_),
    .din2(g1464_p_spl_)
  );


  andX
  g_g1467_p
  (
    .dout(g1467_p),
    .din1(g1465_n_spl_),
    .din2(g1466_n)
  );


  orX
  g_g1467_n
  (
    .dout(g1467_n),
    .din1(g1465_p_spl_),
    .din2(g1466_p)
  );


  andX
  g_g1468_p
  (
    .dout(g1468_p),
    .din1(g1457_n_spl_),
    .din2(g1467_p_spl_)
  );


  orX
  g_g1468_n
  (
    .dout(g1468_n),
    .din1(g1457_p_spl_),
    .din2(g1467_n_spl_)
  );


  andX
  g_g1469_p
  (
    .dout(g1469_p),
    .din1(g1457_p_spl_),
    .din2(g1467_n_spl_)
  );


  orX
  g_g1469_n
  (
    .dout(g1469_n),
    .din1(g1457_n_spl_),
    .din2(g1467_p_spl_)
  );


  andX
  g_g1470_p
  (
    .dout(g1470_p),
    .din1(g1468_n_spl_),
    .din2(g1469_n)
  );


  orX
  g_g1470_n
  (
    .dout(g1470_n),
    .din1(g1468_p_spl_),
    .din2(g1469_p)
  );


  andX
  g_g1471_p
  (
    .dout(g1471_p),
    .din1(g1456_n_spl_),
    .din2(g1470_p_spl_)
  );


  orX
  g_g1471_n
  (
    .dout(g1471_n),
    .din1(g1456_p_spl_),
    .din2(g1470_n_spl_)
  );


  andX
  g_g1472_p
  (
    .dout(g1472_p),
    .din1(g1456_p_spl_),
    .din2(g1470_n_spl_)
  );


  orX
  g_g1472_n
  (
    .dout(g1472_n),
    .din1(g1456_n_spl_),
    .din2(g1470_p_spl_)
  );


  andX
  g_g1473_p
  (
    .dout(g1473_p),
    .din1(g1471_n_spl_),
    .din2(g1472_n)
  );


  orX
  g_g1473_n
  (
    .dout(g1473_n),
    .din1(g1471_p_spl_),
    .din2(g1472_p)
  );


  andX
  g_g1474_p
  (
    .dout(g1474_p),
    .din1(g1455_n_spl_),
    .din2(g1473_p_spl_)
  );


  orX
  g_g1474_n
  (
    .dout(g1474_n),
    .din1(g1455_p),
    .din2(g1473_n)
  );


  orX
  g_g1475_n
  (
    .dout(g1475_n),
    .din1(g1455_n_spl_),
    .din2(g1473_p_spl_)
  );


  andX
  g_g1476_p
  (
    .dout(g1476_p),
    .din1(g1474_n),
    .din2(g1475_n)
  );


  andX
  g_g1477_p
  (
    .dout(g1477_p),
    .din1(g1454_n_spl_),
    .din2(g1476_p_spl_)
  );


  andX
  g_g1478_p
  (
    .dout(g1478_p),
    .din1(g1101_n_spl_),
    .din2(g1104_n_spl_)
  );


  orX
  g_g1478_n
  (
    .dout(g1478_n),
    .din1(g1101_p_spl_),
    .din2(g1104_p_spl_)
  );


  andX
  g_g1479_p
  (
    .dout(g1479_p),
    .din1(ffc_15_p_spl_110),
    .din2(ffc_128_p_spl_1)
  );


  orX
  g_g1479_n
  (
    .dout(g1479_n),
    .din1(ffc_15_n_spl_11),
    .din2(ffc_128_n_spl_)
  );


  andX
  g_g1480_p
  (
    .dout(g1480_p),
    .din1(g1095_n_spl_),
    .din2(g1098_n_spl_)
  );


  orX
  g_g1480_n
  (
    .dout(g1480_n),
    .din1(g1095_p_spl_),
    .din2(g1098_p_spl_)
  );


  andX
  g_g1481_p
  (
    .dout(g1481_p),
    .din1(g1039_p_spl_),
    .din2(g1041_n_spl_)
  );


  orX
  g_g1481_n
  (
    .dout(g1481_n),
    .din1(g1039_n_spl_),
    .din2(g1041_p_spl_)
  );


  andX
  g_g1482_p
  (
    .dout(g1482_p),
    .din1(g1042_n_spl_),
    .din2(g1481_n)
  );


  orX
  g_g1482_n
  (
    .dout(g1482_n),
    .din1(g1042_p_spl_),
    .din2(g1481_p)
  );


  andX
  g_g1483_p
  (
    .dout(g1483_p),
    .din1(g1480_n_spl_),
    .din2(g1482_p_spl_)
  );


  orX
  g_g1483_n
  (
    .dout(g1483_n),
    .din1(g1480_p_spl_),
    .din2(g1482_n_spl_)
  );


  andX
  g_g1484_p
  (
    .dout(g1484_p),
    .din1(g1480_p_spl_),
    .din2(g1482_n_spl_)
  );


  orX
  g_g1484_n
  (
    .dout(g1484_n),
    .din1(g1480_n_spl_),
    .din2(g1482_p_spl_)
  );


  andX
  g_g1485_p
  (
    .dout(g1485_p),
    .din1(g1483_n_spl_),
    .din2(g1484_n)
  );


  orX
  g_g1485_n
  (
    .dout(g1485_n),
    .din1(g1483_p),
    .din2(g1484_p)
  );


  andX
  g_g1486_p
  (
    .dout(g1486_p),
    .din1(g1479_n_spl_),
    .din2(g1485_p_spl_)
  );


  orX
  g_g1486_n
  (
    .dout(g1486_n),
    .din1(g1479_p_spl_),
    .din2(g1485_n_spl_)
  );


  andX
  g_g1487_p
  (
    .dout(g1487_p),
    .din1(g1479_p_spl_),
    .din2(g1485_n_spl_)
  );


  orX
  g_g1487_n
  (
    .dout(g1487_n),
    .din1(g1479_n_spl_),
    .din2(g1485_p_spl_)
  );


  andX
  g_g1488_p
  (
    .dout(g1488_p),
    .din1(g1486_n_spl_),
    .din2(g1487_n)
  );


  orX
  g_g1488_n
  (
    .dout(g1488_n),
    .din1(g1486_p),
    .din2(g1487_p)
  );


  orX
  g_g1489_n
  (
    .dout(g1489_n),
    .din1(g1478_p),
    .din2(g1488_n)
  );


  andX
  g_g1490_p
  (
    .dout(g1490_p),
    .din1(g1158_n_spl_),
    .din2(g1161_n_spl_)
  );


  orX
  g_g1490_n
  (
    .dout(g1490_n),
    .din1(g1158_p_spl_),
    .din2(g1161_p_spl_)
  );


  andX
  g_g1491_p
  (
    .dout(g1491_p),
    .din1(ffc_17_p_spl_10),
    .din2(ffc_125_p_spl_1)
  );


  orX
  g_g1491_n
  (
    .dout(g1491_n),
    .din1(ffc_17_n_spl_11),
    .din2(ffc_125_n_spl_)
  );


  andX
  g_g1492_p
  (
    .dout(g1492_p),
    .din1(g1152_n_spl_),
    .din2(g1155_n_spl_)
  );


  orX
  g_g1492_n
  (
    .dout(g1492_n),
    .din1(g1152_p_spl_),
    .din2(g1155_p_spl_)
  );


  andX
  g_g1493_p
  (
    .dout(g1493_p),
    .din1(g1084_p_spl_),
    .din2(g1086_n_spl_)
  );


  orX
  g_g1493_n
  (
    .dout(g1493_n),
    .din1(g1084_n_spl_),
    .din2(g1086_p_spl_)
  );


  andX
  g_g1494_p
  (
    .dout(g1494_p),
    .din1(g1087_n_spl_),
    .din2(g1493_n)
  );


  orX
  g_g1494_n
  (
    .dout(g1494_n),
    .din1(g1087_p_spl_),
    .din2(g1493_p)
  );


  andX
  g_g1495_p
  (
    .dout(g1495_p),
    .din1(g1492_n_spl_),
    .din2(g1494_p_spl_)
  );


  orX
  g_g1495_n
  (
    .dout(g1495_n),
    .din1(g1492_p_spl_),
    .din2(g1494_n_spl_)
  );


  andX
  g_g1496_p
  (
    .dout(g1496_p),
    .din1(g1492_p_spl_),
    .din2(g1494_n_spl_)
  );


  orX
  g_g1496_n
  (
    .dout(g1496_n),
    .din1(g1492_n_spl_),
    .din2(g1494_p_spl_)
  );


  andX
  g_g1497_p
  (
    .dout(g1497_p),
    .din1(g1495_n_spl_),
    .din2(g1496_n)
  );


  orX
  g_g1497_n
  (
    .dout(g1497_n),
    .din1(g1495_p),
    .din2(g1496_p)
  );


  andX
  g_g1498_p
  (
    .dout(g1498_p),
    .din1(g1491_n_spl_),
    .din2(g1497_p_spl_)
  );


  orX
  g_g1498_n
  (
    .dout(g1498_n),
    .din1(g1491_p_spl_),
    .din2(g1497_n_spl_)
  );


  andX
  g_g1499_p
  (
    .dout(g1499_p),
    .din1(g1491_p_spl_),
    .din2(g1497_n_spl_)
  );


  orX
  g_g1499_n
  (
    .dout(g1499_n),
    .din1(g1491_n_spl_),
    .din2(g1497_p_spl_)
  );


  andX
  g_g1500_p
  (
    .dout(g1500_p),
    .din1(g1498_n_spl_),
    .din2(g1499_n)
  );


  orX
  g_g1500_n
  (
    .dout(g1500_n),
    .din1(g1498_p),
    .din2(g1499_p)
  );


  orX
  g_g1501_n
  (
    .dout(g1501_n),
    .din1(g1490_p),
    .din2(g1500_n)
  );


  andX
  g_g1502_p
  (
    .dout(g1502_p),
    .din1(g1235_n_spl_),
    .din2(g1238_n_spl_)
  );


  orX
  g_g1502_n
  (
    .dout(g1502_n),
    .din1(g1235_p_spl_),
    .din2(g1238_p_spl_)
  );


  andX
  g_g1503_p
  (
    .dout(g1503_p),
    .din1(ffc_19_p_spl_10),
    .din2(ffc_122_p_spl_1)
  );


  orX
  g_g1503_n
  (
    .dout(g1503_n),
    .din1(ffc_19_n_spl_11),
    .din2(ffc_122_n_spl_1)
  );


  andX
  g_g1504_p
  (
    .dout(g1504_p),
    .din1(g1229_n_spl_),
    .din2(g1232_n_spl_)
  );


  orX
  g_g1504_n
  (
    .dout(g1504_n),
    .din1(g1229_p_spl_),
    .din2(g1232_p_spl_)
  );


  andX
  g_g1505_p
  (
    .dout(g1505_p),
    .din1(g1141_p_spl_),
    .din2(g1143_n_spl_)
  );


  orX
  g_g1505_n
  (
    .dout(g1505_n),
    .din1(g1141_n_spl_),
    .din2(g1143_p_spl_)
  );


  andX
  g_g1506_p
  (
    .dout(g1506_p),
    .din1(g1144_n_spl_),
    .din2(g1505_n)
  );


  orX
  g_g1506_n
  (
    .dout(g1506_n),
    .din1(g1144_p_spl_),
    .din2(g1505_p)
  );


  andX
  g_g1507_p
  (
    .dout(g1507_p),
    .din1(g1504_n_spl_),
    .din2(g1506_p_spl_)
  );


  orX
  g_g1507_n
  (
    .dout(g1507_n),
    .din1(g1504_p_spl_),
    .din2(g1506_n_spl_)
  );


  andX
  g_g1508_p
  (
    .dout(g1508_p),
    .din1(g1504_p_spl_),
    .din2(g1506_n_spl_)
  );


  orX
  g_g1508_n
  (
    .dout(g1508_n),
    .din1(g1504_n_spl_),
    .din2(g1506_p_spl_)
  );


  andX
  g_g1509_p
  (
    .dout(g1509_p),
    .din1(g1507_n_spl_),
    .din2(g1508_n)
  );


  orX
  g_g1509_n
  (
    .dout(g1509_n),
    .din1(g1507_p),
    .din2(g1508_p)
  );


  andX
  g_g1510_p
  (
    .dout(g1510_p),
    .din1(g1503_n_spl_),
    .din2(g1509_p_spl_)
  );


  orX
  g_g1510_n
  (
    .dout(g1510_n),
    .din1(g1503_p_spl_),
    .din2(g1509_n_spl_)
  );


  andX
  g_g1511_p
  (
    .dout(g1511_p),
    .din1(g1503_p_spl_),
    .din2(g1509_n_spl_)
  );


  orX
  g_g1511_n
  (
    .dout(g1511_n),
    .din1(g1503_n_spl_),
    .din2(g1509_p_spl_)
  );


  andX
  g_g1512_p
  (
    .dout(g1512_p),
    .din1(g1510_n_spl_),
    .din2(g1511_n)
  );


  orX
  g_g1512_n
  (
    .dout(g1512_n),
    .din1(g1510_p),
    .din2(g1511_p)
  );


  orX
  g_g1513_n
  (
    .dout(g1513_n),
    .din1(g1502_p),
    .din2(g1512_n)
  );


  orX
  g_g1514_n
  (
    .dout(g1514_n),
    .din1(g1251_n),
    .din2(g1277_p)
  );


  andX
  g_g1515_p
  (
    .dout(g1515_p),
    .din1(g1278_n_spl_),
    .din2(g1514_n)
  );


  andX
  g_g1516_p
  (
    .dout(g1516_p),
    .din1(ffc_12_p_spl_000),
    .din2(ffc_187_p_spl_1)
  );


  orX
  g_g1516_n
  (
    .dout(g1516_n),
    .din1(ffc_12_n_spl_000),
    .din2(ffc_187_n_spl_1)
  );


  andX
  g_g1517_p
  (
    .dout(g1517_p),
    .din1(g1380_p_spl_),
    .din2(g1398_n_spl_)
  );


  orX
  g_g1517_n
  (
    .dout(g1517_n),
    .din1(g1380_n_spl_),
    .din2(g1398_p_spl_)
  );


  andX
  g_g1518_p
  (
    .dout(g1518_p),
    .din1(g1399_n_spl_),
    .din2(g1517_n)
  );


  orX
  g_g1518_n
  (
    .dout(g1518_n),
    .din1(g1399_p),
    .din2(g1517_p)
  );


  orX
  g_g1519_n
  (
    .dout(g1519_n),
    .din1(g1516_p),
    .din2(g1518_n)
  );


  andX
  g_g1520_p
  (
    .dout(g1520_p),
    .din1(ffc_11_p_spl_001),
    .din2(ffc_190_p_spl_1)
  );


  orX
  g_g1520_n
  (
    .dout(g1520_n),
    .din1(ffc_11_n_spl_001),
    .din2(ffc_190_n_spl_)
  );


  andX
  g_g1521_p
  (
    .dout(g1521_p),
    .din1(g1310_p_spl_),
    .din2(g1327_n_spl_)
  );


  orX
  g_g1521_n
  (
    .dout(g1521_n),
    .din1(g1310_n_spl_),
    .din2(g1327_p_spl_)
  );


  andX
  g_g1522_p
  (
    .dout(g1522_p),
    .din1(g1328_n_spl_),
    .din2(g1521_n)
  );


  orX
  g_g1522_n
  (
    .dout(g1522_n),
    .din1(g1328_p),
    .din2(g1521_p)
  );


  orX
  g_g1523_n
  (
    .dout(g1523_n),
    .din1(g1520_p),
    .din2(g1522_n)
  );


  andX
  g_g1524_p
  (
    .dout(g1524_p),
    .din1(g1322_n_spl_),
    .din2(g1325_n_spl_)
  );


  orX
  g_g1524_n
  (
    .dout(g1524_n),
    .din1(g1322_p_spl_),
    .din2(g1325_p_spl_)
  );


  andX
  g_g1525_p
  (
    .dout(g1525_p),
    .din1(ffc_10_p_spl_011),
    .din2(ffc_192_p_spl_1)
  );


  orX
  g_g1525_n
  (
    .dout(g1525_n),
    .din1(ffc_10_n_spl_011),
    .din2(ffc_192_n_spl_)
  );


  andX
  g_g1526_p
  (
    .dout(g1526_p),
    .din1(ffc_9_p_spl_100),
    .din2(ffc_193_p_spl_0)
  );


  orX
  g_g1526_n
  (
    .dout(g1526_n),
    .din1(ffc_9_n_spl_100),
    .din2(ffc_193_n_spl_0)
  );


  andX
  g_g1527_p
  (
    .dout(g1527_p),
    .din1(g1316_n_spl_),
    .din2(g1319_n_spl_)
  );


  orX
  g_g1527_n
  (
    .dout(g1527_n),
    .din1(g1316_p_spl_),
    .din2(g1319_p_spl_)
  );


  andX
  g_g1528_p
  (
    .dout(g1528_p),
    .din1(g1526_n_spl_),
    .din2(g1527_n_spl_)
  );


  orX
  g_g1528_n
  (
    .dout(g1528_n),
    .din1(g1526_p_spl_),
    .din2(g1527_p_spl_)
  );


  andX
  g_g1529_p
  (
    .dout(g1529_p),
    .din1(g1526_p_spl_),
    .din2(g1527_p_spl_)
  );


  orX
  g_g1529_n
  (
    .dout(g1529_n),
    .din1(g1526_n_spl_),
    .din2(g1527_n_spl_)
  );


  andX
  g_g1530_p
  (
    .dout(g1530_p),
    .din1(g1528_n),
    .din2(g1529_n)
  );


  orX
  g_g1530_n
  (
    .dout(g1530_n),
    .din1(g1528_p_spl_),
    .din2(g1529_p)
  );


  andX
  g_g1531_p
  (
    .dout(g1531_p),
    .din1(g1525_n_spl_),
    .din2(g1530_p_spl_)
  );


  orX
  g_g1531_n
  (
    .dout(g1531_n),
    .din1(g1525_p_spl_),
    .din2(g1530_n_spl_)
  );


  andX
  g_g1532_p
  (
    .dout(g1532_p),
    .din1(g1525_p_spl_),
    .din2(g1530_n_spl_)
  );


  orX
  g_g1532_n
  (
    .dout(g1532_n),
    .din1(g1525_n_spl_),
    .din2(g1530_p_spl_)
  );


  andX
  g_g1533_p
  (
    .dout(g1533_p),
    .din1(g1531_n),
    .din2(g1532_n)
  );


  orX
  g_g1533_n
  (
    .dout(g1533_n),
    .din1(g1531_p_spl_),
    .din2(g1532_p)
  );


  orX
  g_g1534_n
  (
    .dout(g1534_n),
    .din1(g1524_p),
    .din2(g1533_n)
  );


  andX
  g_g1535_p
  (
    .dout(g1535_p),
    .din1(g1393_n_spl_),
    .din2(g1396_n_spl_)
  );


  orX
  g_g1535_n
  (
    .dout(g1535_n),
    .din1(g1393_p_spl_),
    .din2(g1396_p_spl_)
  );


  andX
  g_g1536_p
  (
    .dout(g1536_p),
    .din1(ffc_11_p_spl_010),
    .din2(ffc_189_p_spl_1)
  );


  orX
  g_g1536_n
  (
    .dout(g1536_n),
    .din1(ffc_11_n_spl_010),
    .din2(ffc_189_n_spl_)
  );


  andX
  g_g1537_p
  (
    .dout(g1537_p),
    .din1(g1387_n_spl_),
    .din2(g1390_n_spl_)
  );


  orX
  g_g1537_n
  (
    .dout(g1537_n),
    .din1(g1387_p_spl_),
    .din2(g1390_p_spl_)
  );


  andX
  g_g1538_p
  (
    .dout(g1538_p),
    .din1(g1306_p_spl_),
    .din2(g1308_n_spl_)
  );


  orX
  g_g1538_n
  (
    .dout(g1538_n),
    .din1(g1306_n_spl_),
    .din2(g1308_p_spl_)
  );


  andX
  g_g1539_p
  (
    .dout(g1539_p),
    .din1(g1309_n_spl_),
    .din2(g1538_n)
  );


  orX
  g_g1539_n
  (
    .dout(g1539_n),
    .din1(g1309_p_spl_),
    .din2(g1538_p)
  );


  andX
  g_g1540_p
  (
    .dout(g1540_p),
    .din1(g1537_n_spl_),
    .din2(g1539_p_spl_)
  );


  orX
  g_g1540_n
  (
    .dout(g1540_n),
    .din1(g1537_p_spl_),
    .din2(g1539_n_spl_)
  );


  andX
  g_g1541_p
  (
    .dout(g1541_p),
    .din1(g1537_p_spl_),
    .din2(g1539_n_spl_)
  );


  orX
  g_g1541_n
  (
    .dout(g1541_n),
    .din1(g1537_n_spl_),
    .din2(g1539_p_spl_)
  );


  andX
  g_g1542_p
  (
    .dout(g1542_p),
    .din1(g1540_n),
    .din2(g1541_n)
  );


  orX
  g_g1542_n
  (
    .dout(g1542_n),
    .din1(g1540_p_spl_),
    .din2(g1541_p)
  );


  andX
  g_g1543_p
  (
    .dout(g1543_p),
    .din1(g1536_n_spl_),
    .din2(g1542_p_spl_)
  );


  orX
  g_g1543_n
  (
    .dout(g1543_n),
    .din1(g1536_p_spl_),
    .din2(g1542_n_spl_)
  );


  andX
  g_g1544_p
  (
    .dout(g1544_p),
    .din1(g1536_p_spl_),
    .din2(g1542_n_spl_)
  );


  orX
  g_g1544_n
  (
    .dout(g1544_n),
    .din1(g1536_n_spl_),
    .din2(g1542_p_spl_)
  );


  andX
  g_g1545_p
  (
    .dout(g1545_p),
    .din1(g1543_n),
    .din2(g1544_n)
  );


  orX
  g_g1545_n
  (
    .dout(g1545_n),
    .din1(g1543_p_spl_),
    .din2(g1544_p)
  );


  orX
  g_g1546_n
  (
    .dout(g1546_n),
    .din1(g1535_p),
    .din2(g1545_n)
  );


  andX
  g_g1547_p
  (
    .dout(g1547_p),
    .din1(g1010_n_spl_),
    .din2(g1242_n)
  );


  orX
  g_g1547_n
  (
    .dout(g1547_n),
    .din1(g1010_p_spl_),
    .din2(g1242_p_spl_)
  );


  andX
  g_g1548_p
  (
    .dout(g1548_p),
    .din1(ffc_11_p_spl_010),
    .din2(ffc_195_p_spl_0)
  );


  orX
  g_g1548_n
  (
    .dout(g1548_n),
    .din1(ffc_11_n_spl_010),
    .din2(ffc_195_n_spl_1)
  );


  andX
  g_g1549_p
  (
    .dout(g1549_p),
    .din1(g1004_n_spl_),
    .din2(g1007_n_spl_)
  );


  orX
  g_g1549_n
  (
    .dout(g1549_n),
    .din1(g1004_p_spl_),
    .din2(g1007_p_spl_)
  );


  andX
  g_g1550_p
  (
    .dout(g1550_p),
    .din1(ffc_10_p_spl_100),
    .din2(ffc_180_p_spl_00)
  );


  orX
  g_g1550_n
  (
    .dout(g1550_n),
    .din1(ffc_10_n_spl_100),
    .din2(ffc_180_n_spl_0)
  );


  andX
  g_g1551_p
  (
    .dout(g1551_p),
    .din1(g998_n_spl_),
    .din2(g1001_n_spl_)
  );


  orX
  g_g1551_n
  (
    .dout(g1551_n),
    .din1(g998_p_spl_),
    .din2(g1001_p_spl_)
  );


  andX
  g_g1552_p
  (
    .dout(g1552_p),
    .din1(ffc_9_p_spl_101),
    .din2(ffc_181_p_spl_00)
  );


  orX
  g_g1552_n
  (
    .dout(g1552_n),
    .din1(ffc_9_n_spl_101),
    .din2(ffc_181_n_spl_0)
  );


  andX
  g_g1553_p
  (
    .dout(g1553_p),
    .din1(ffc_313_p),
    .din2(g995_n_spl_)
  );


  orX
  g_g1553_n
  (
    .dout(g1553_n),
    .din1(ffc_313_n),
    .din2(g995_p_spl_)
  );


  andX
  g_g1554_p
  (
    .dout(g1554_p),
    .din1(ffc_328_n_spl_),
    .din2(ffc_345_p_spl_)
  );


  orX
  g_g1554_n
  (
    .dout(g1554_n),
    .din1(ffc_328_p_spl_),
    .din2(ffc_345_n_spl_)
  );


  andX
  g_g1555_p
  (
    .dout(g1555_p),
    .din1(ffc_328_p_spl_),
    .din2(ffc_345_n_spl_)
  );


  orX
  g_g1555_n
  (
    .dout(g1555_n),
    .din1(ffc_328_n_spl_),
    .din2(ffc_345_p_spl_)
  );


  andX
  g_g1556_p
  (
    .dout(g1556_p),
    .din1(g1554_n_spl_),
    .din2(g1555_n)
  );


  orX
  g_g1556_n
  (
    .dout(g1556_n),
    .din1(g1554_p_spl_),
    .din2(g1555_p)
  );


  andX
  g_g1557_p
  (
    .dout(g1557_p),
    .din1(g1553_n_spl_),
    .din2(g1556_p_spl_)
  );


  orX
  g_g1557_n
  (
    .dout(g1557_n),
    .din1(g1553_p_spl_),
    .din2(g1556_n_spl_)
  );


  andX
  g_g1558_p
  (
    .dout(g1558_p),
    .din1(g1553_p_spl_),
    .din2(g1556_n_spl_)
  );


  orX
  g_g1558_n
  (
    .dout(g1558_n),
    .din1(g1553_n_spl_),
    .din2(g1556_p_spl_)
  );


  andX
  g_g1559_p
  (
    .dout(g1559_p),
    .din1(g1557_n_spl_),
    .din2(g1558_n)
  );


  orX
  g_g1559_n
  (
    .dout(g1559_n),
    .din1(g1557_p_spl_),
    .din2(g1558_p)
  );


  andX
  g_g1560_p
  (
    .dout(g1560_p),
    .din1(g1552_n_spl_),
    .din2(g1559_p_spl_)
  );


  orX
  g_g1560_n
  (
    .dout(g1560_n),
    .din1(g1552_p_spl_),
    .din2(g1559_n_spl_)
  );


  andX
  g_g1561_p
  (
    .dout(g1561_p),
    .din1(g1552_p_spl_),
    .din2(g1559_n_spl_)
  );


  orX
  g_g1561_n
  (
    .dout(g1561_n),
    .din1(g1552_n_spl_),
    .din2(g1559_p_spl_)
  );


  andX
  g_g1562_p
  (
    .dout(g1562_p),
    .din1(g1560_n_spl_),
    .din2(g1561_n)
  );


  orX
  g_g1562_n
  (
    .dout(g1562_n),
    .din1(g1560_p_spl_),
    .din2(g1561_p)
  );


  andX
  g_g1563_p
  (
    .dout(g1563_p),
    .din1(g1551_n_spl_),
    .din2(g1562_p_spl_)
  );


  orX
  g_g1563_n
  (
    .dout(g1563_n),
    .din1(g1551_p_spl_),
    .din2(g1562_n_spl_)
  );


  andX
  g_g1564_p
  (
    .dout(g1564_p),
    .din1(g1551_p_spl_),
    .din2(g1562_n_spl_)
  );


  orX
  g_g1564_n
  (
    .dout(g1564_n),
    .din1(g1551_n_spl_),
    .din2(g1562_p_spl_)
  );


  andX
  g_g1565_p
  (
    .dout(g1565_p),
    .din1(g1563_n_spl_),
    .din2(g1564_n)
  );


  orX
  g_g1565_n
  (
    .dout(g1565_n),
    .din1(g1563_p_spl_),
    .din2(g1564_p)
  );


  andX
  g_g1566_p
  (
    .dout(g1566_p),
    .din1(g1550_n_spl_),
    .din2(g1565_p_spl_)
  );


  orX
  g_g1566_n
  (
    .dout(g1566_n),
    .din1(g1550_p_spl_),
    .din2(g1565_n_spl_)
  );


  andX
  g_g1567_p
  (
    .dout(g1567_p),
    .din1(g1550_p_spl_),
    .din2(g1565_n_spl_)
  );


  orX
  g_g1567_n
  (
    .dout(g1567_n),
    .din1(g1550_n_spl_),
    .din2(g1565_p_spl_)
  );


  andX
  g_g1568_p
  (
    .dout(g1568_p),
    .din1(g1566_n_spl_),
    .din2(g1567_n)
  );


  orX
  g_g1568_n
  (
    .dout(g1568_n),
    .din1(g1566_p_spl_),
    .din2(g1567_p)
  );


  andX
  g_g1569_p
  (
    .dout(g1569_p),
    .din1(g1549_n_spl_),
    .din2(g1568_p_spl_)
  );


  orX
  g_g1569_n
  (
    .dout(g1569_n),
    .din1(g1549_p_spl_),
    .din2(g1568_n_spl_)
  );


  andX
  g_g1570_p
  (
    .dout(g1570_p),
    .din1(g1549_p_spl_),
    .din2(g1568_n_spl_)
  );


  orX
  g_g1570_n
  (
    .dout(g1570_n),
    .din1(g1549_n_spl_),
    .din2(g1568_p_spl_)
  );


  andX
  g_g1571_p
  (
    .dout(g1571_p),
    .din1(g1569_n_spl_),
    .din2(g1570_n)
  );


  orX
  g_g1571_n
  (
    .dout(g1571_n),
    .din1(g1569_p_spl_),
    .din2(g1570_p)
  );


  andX
  g_g1572_p
  (
    .dout(g1572_p),
    .din1(g1548_n_spl_),
    .din2(g1571_p_spl_)
  );


  orX
  g_g1572_n
  (
    .dout(g1572_n),
    .din1(g1548_p_spl_),
    .din2(g1571_n_spl_)
  );


  andX
  g_g1573_p
  (
    .dout(g1573_p),
    .din1(g1548_p_spl_),
    .din2(g1571_n_spl_)
  );


  orX
  g_g1573_n
  (
    .dout(g1573_n),
    .din1(g1548_n_spl_),
    .din2(g1571_p_spl_)
  );


  andX
  g_g1574_p
  (
    .dout(g1574_p),
    .din1(g1572_n_spl_),
    .din2(g1573_n)
  );


  orX
  g_g1574_n
  (
    .dout(g1574_n),
    .din1(g1572_p_spl_),
    .din2(g1573_p)
  );


  andX
  g_g1575_p
  (
    .dout(g1575_p),
    .din1(g1547_n_spl_),
    .din2(g1574_p_spl_)
  );


  orX
  g_g1575_n
  (
    .dout(g1575_n),
    .din1(g1547_p),
    .din2(g1574_n)
  );


  orX
  g_g1576_n
  (
    .dout(g1576_n),
    .din1(g1547_n_spl_),
    .din2(g1574_p_spl_)
  );


  andX
  g_g1577_p
  (
    .dout(g1577_p),
    .din1(g1575_n),
    .din2(g1576_n)
  );


  andX
  g_g1578_p
  (
    .dout(g1578_p),
    .din1(g1248_n_spl_),
    .din2(g1400_n)
  );


  orX
  g_g1578_n
  (
    .dout(g1578_n),
    .din1(g1248_p_spl_),
    .din2(g1400_p_spl_)
  );


  andX
  g_g1579_p
  (
    .dout(g1579_p),
    .din1(G2_p_spl_01),
    .din2(G19_p_spl_000)
  );


  orX
  g_g1579_n
  (
    .dout(g1579_n),
    .din1(G2_n_spl_1),
    .din2(G19_n_spl_000)
  );


  andX
  g_g1580_p
  (
    .dout(g1580_p),
    .din1(G4_p_spl_00),
    .din2(G17_p_spl_001)
  );


  orX
  g_g1580_n
  (
    .dout(g1580_n),
    .din1(G4_n_spl_0),
    .din2(G17_n_spl_001)
  );


  andX
  g_g1581_p
  (
    .dout(g1581_p),
    .din1(G3_p_spl_00),
    .din2(G18_p_spl_001)
  );


  orX
  g_g1581_n
  (
    .dout(g1581_n),
    .din1(G3_n_spl_0),
    .din2(G18_n_spl_001)
  );


  andX
  g_g1582_p
  (
    .dout(g1582_p),
    .din1(g1580_p_spl_),
    .din2(g1581_p_spl_)
  );


  orX
  g_g1582_n
  (
    .dout(g1582_n),
    .din1(g1580_n_spl_),
    .din2(g1581_n_spl_)
  );


  andX
  g_g1583_p
  (
    .dout(g1583_p),
    .din1(g1580_n_spl_),
    .din2(g1581_n_spl_)
  );


  orX
  g_g1583_n
  (
    .dout(g1583_n),
    .din1(g1580_p_spl_),
    .din2(g1581_p_spl_)
  );


  andX
  g_g1584_p
  (
    .dout(g1584_p),
    .din1(g1582_n_spl_0),
    .din2(g1583_n)
  );


  orX
  g_g1584_n
  (
    .dout(g1584_n),
    .din1(g1582_p_spl_0),
    .din2(g1583_p)
  );


  andX
  g_g1585_p
  (
    .dout(g1585_p),
    .din1(g1245_n_spl_0),
    .din2(g1584_n_spl_)
  );


  orX
  g_g1585_n
  (
    .dout(g1585_n),
    .din1(g1245_p_spl_0),
    .din2(g1584_p_spl_)
  );


  andX
  g_g1586_p
  (
    .dout(g1586_p),
    .din1(g1245_p_spl_),
    .din2(g1584_p_spl_)
  );


  orX
  g_g1586_n
  (
    .dout(g1586_n),
    .din1(g1245_n_spl_),
    .din2(g1584_n_spl_)
  );


  andX
  g_g1587_p
  (
    .dout(g1587_p),
    .din1(g1585_n_spl_),
    .din2(g1586_n)
  );


  orX
  g_g1587_n
  (
    .dout(g1587_n),
    .din1(g1585_p_spl_),
    .din2(g1586_p)
  );


  andX
  g_g1588_p
  (
    .dout(g1588_p),
    .din1(g1579_n_spl_),
    .din2(g1587_p_spl_)
  );


  orX
  g_g1588_n
  (
    .dout(g1588_n),
    .din1(g1579_p_spl_),
    .din2(g1587_n_spl_)
  );


  andX
  g_g1589_p
  (
    .dout(g1589_p),
    .din1(g1579_p_spl_),
    .din2(g1587_n_spl_)
  );


  orX
  g_g1589_n
  (
    .dout(g1589_n),
    .din1(g1579_n_spl_),
    .din2(g1587_p_spl_)
  );


  andX
  g_g1590_p
  (
    .dout(g1590_p),
    .din1(g1588_n_spl_),
    .din2(g1589_n)
  );


  orX
  g_g1590_n
  (
    .dout(g1590_n),
    .din1(g1588_p_spl_),
    .din2(g1589_p)
  );


  andX
  g_g1591_p
  (
    .dout(g1591_p),
    .din1(g1578_n_spl_),
    .din2(g1590_p_spl_)
  );


  orX
  g_g1591_n
  (
    .dout(g1591_n),
    .din1(g1578_p),
    .din2(g1590_n)
  );


  orX
  g_g1592_n
  (
    .dout(g1592_n),
    .din1(g1578_n_spl_),
    .din2(g1590_p_spl_)
  );


  andX
  g_g1593_p
  (
    .dout(g1593_p),
    .din1(g1591_n),
    .din2(g1592_n)
  );


  andX
  g_g1594_p
  (
    .dout(g1594_p),
    .din1(ffc_21_p_spl_00),
    .din2(ffc_121_p_spl_1)
  );


  andX
  g_g1595_p
  (
    .dout(g1595_p),
    .din1(ffc_19_p_spl_10),
    .din2(ffc_124_p_spl_1)
  );


  andX
  g_g1596_p
  (
    .dout(g1596_p),
    .din1(ffc_17_p_spl_11),
    .din2(ffc_127_p_spl_1)
  );


  andX
  g_g1597_p
  (
    .dout(g1597_p),
    .din1(ffc_15_p_spl_111),
    .din2(ffc_130_p_spl_1)
  );


  andX
  g_g1598_p
  (
    .dout(g1598_p),
    .din1(g1483_n_spl_),
    .din2(g1486_n_spl_)
  );


  andX
  g_g1599_p
  (
    .dout(g1599_p),
    .din1(g1495_n_spl_),
    .din2(g1498_n_spl_)
  );


  andX
  g_g1600_p
  (
    .dout(g1600_p),
    .din1(g1507_n_spl_),
    .din2(g1510_n_spl_)
  );


  andX
  g_g1601_p
  (
    .dout(g1601_p),
    .din1(g1468_n_spl_),
    .din2(g1471_n_spl_)
  );


  orX
  g_g1601_n
  (
    .dout(g1601_n),
    .din1(g1468_p_spl_),
    .din2(g1471_p_spl_)
  );


  andX
  g_g1602_p
  (
    .dout(g1602_p),
    .din1(ffc_19_p_spl_11),
    .din2(ffc_119_p_spl_01)
  );


  orX
  g_g1602_n
  (
    .dout(g1602_n),
    .din1(ffc_19_n_spl_11),
    .din2(ffc_119_n_spl_1)
  );


  andX
  g_g1603_p
  (
    .dout(g1603_p),
    .din1(g1462_n_spl_),
    .din2(g1465_n_spl_)
  );


  orX
  g_g1603_n
  (
    .dout(g1603_n),
    .din1(g1462_p_spl_),
    .din2(g1465_p_spl_)
  );


  andX
  g_g1604_p
  (
    .dout(g1604_p),
    .din1(g1194_p_spl_),
    .din2(g1196_n_spl_)
  );


  orX
  g_g1604_n
  (
    .dout(g1604_n),
    .din1(g1194_n_spl_),
    .din2(g1196_p_spl_)
  );


  andX
  g_g1605_p
  (
    .dout(g1605_p),
    .din1(g1197_n_spl_),
    .din2(g1604_n)
  );


  orX
  g_g1605_n
  (
    .dout(g1605_n),
    .din1(g1197_p_spl_),
    .din2(g1604_p)
  );


  andX
  g_g1606_p
  (
    .dout(g1606_p),
    .din1(g1603_n_spl_),
    .din2(g1605_p_spl_)
  );


  orX
  g_g1606_n
  (
    .dout(g1606_n),
    .din1(g1603_p_spl_),
    .din2(g1605_n_spl_)
  );


  andX
  g_g1607_p
  (
    .dout(g1607_p),
    .din1(g1603_p_spl_),
    .din2(g1605_n_spl_)
  );


  orX
  g_g1607_n
  (
    .dout(g1607_n),
    .din1(g1603_n_spl_),
    .din2(g1605_p_spl_)
  );


  andX
  g_g1608_p
  (
    .dout(g1608_p),
    .din1(g1606_n_spl_),
    .din2(g1607_n)
  );


  orX
  g_g1608_n
  (
    .dout(g1608_n),
    .din1(g1606_p_spl_),
    .din2(g1607_p)
  );


  andX
  g_g1609_p
  (
    .dout(g1609_p),
    .din1(g1602_n_spl_),
    .din2(g1608_p_spl_)
  );


  orX
  g_g1609_n
  (
    .dout(g1609_n),
    .din1(g1602_p_spl_),
    .din2(g1608_n_spl_)
  );


  andX
  g_g1610_p
  (
    .dout(g1610_p),
    .din1(g1602_p_spl_),
    .din2(g1608_n_spl_)
  );


  orX
  g_g1610_n
  (
    .dout(g1610_n),
    .din1(g1602_n_spl_),
    .din2(g1608_p_spl_)
  );


  andX
  g_g1611_p
  (
    .dout(g1611_p),
    .din1(g1609_n_spl_),
    .din2(g1610_n)
  );


  orX
  g_g1611_n
  (
    .dout(g1611_n),
    .din1(g1609_p_spl_),
    .din2(g1610_p)
  );


  andX
  g_g1612_p
  (
    .dout(g1612_p),
    .din1(g1601_n_spl_),
    .din2(g1611_p_spl_)
  );


  orX
  g_g1612_n
  (
    .dout(g1612_n),
    .din1(g1601_p_spl_),
    .din2(g1611_n_spl_)
  );


  andX
  g_g1613_p
  (
    .dout(g1613_p),
    .din1(ffc_21_p_spl_0),
    .din2(ffc_118_p_spl_1)
  );


  orX
  g_g1613_n
  (
    .dout(g1613_n),
    .din1(ffc_21_n_spl_1),
    .din2(ffc_118_n_spl_1)
  );


  andX
  g_g1614_p
  (
    .dout(g1614_p),
    .din1(g1601_p_spl_),
    .din2(g1611_n_spl_)
  );


  orX
  g_g1614_n
  (
    .dout(g1614_n),
    .din1(g1601_n_spl_),
    .din2(g1611_p_spl_)
  );


  andX
  g_g1615_p
  (
    .dout(g1615_p),
    .din1(g1612_n_spl_),
    .din2(g1614_n)
  );


  orX
  g_g1615_n
  (
    .dout(g1615_n),
    .din1(g1612_p),
    .din2(g1614_p)
  );


  orX
  g_g1616_n
  (
    .dout(g1616_n),
    .din1(g1613_p),
    .din2(g1615_n)
  );


  andX
  g_g1617_p
  (
    .dout(g1617_p),
    .din1(g1612_n_spl_),
    .din2(g1616_n_spl_)
  );


  andX
  g_g1618_p
  (
    .dout(g1618_p),
    .din1(g1606_n_spl_),
    .din2(g1609_n_spl_)
  );


  orX
  g_g1618_n
  (
    .dout(g1618_n),
    .din1(g1606_p_spl_),
    .din2(g1609_p_spl_)
  );


  andX
  g_g1619_p
  (
    .dout(g1619_p),
    .din1(g1218_p_spl_),
    .din2(g1220_n_spl_)
  );


  orX
  g_g1619_n
  (
    .dout(g1619_n),
    .din1(g1218_n_spl_),
    .din2(g1220_p_spl_)
  );


  andX
  g_g1620_p
  (
    .dout(g1620_p),
    .din1(g1221_n_spl_),
    .din2(g1619_n)
  );


  orX
  g_g1620_n
  (
    .dout(g1620_n),
    .din1(g1221_p_spl_),
    .din2(g1619_p)
  );


  andX
  g_g1621_p
  (
    .dout(g1621_p),
    .din1(g1618_n_spl_),
    .din2(g1620_p_spl_)
  );


  orX
  g_g1621_n
  (
    .dout(g1621_n),
    .din1(g1618_p_spl_),
    .din2(g1620_n_spl_)
  );


  andX
  g_g1622_p
  (
    .dout(g1622_p),
    .din1(ffc_21_p_spl_1),
    .din2(ffc_119_p_spl_1)
  );


  orX
  g_g1622_n
  (
    .dout(g1622_n),
    .din1(ffc_21_n_spl_1),
    .din2(ffc_119_n_spl_1)
  );


  andX
  g_g1623_p
  (
    .dout(g1623_p),
    .din1(g1618_p_spl_),
    .din2(g1620_n_spl_)
  );


  orX
  g_g1623_n
  (
    .dout(g1623_n),
    .din1(g1618_n_spl_),
    .din2(g1620_p_spl_)
  );


  andX
  g_g1624_p
  (
    .dout(g1624_p),
    .din1(g1621_n_spl_),
    .din2(g1623_n)
  );


  orX
  g_g1624_n
  (
    .dout(g1624_n),
    .din1(g1621_p),
    .din2(g1623_p)
  );


  orX
  g_g1625_n
  (
    .dout(g1625_n),
    .din1(g1622_p),
    .din2(g1624_n)
  );


  andX
  g_g1626_p
  (
    .dout(g1626_p),
    .din1(g1621_n_spl_),
    .din2(g1625_n_spl_)
  );


  orX
  g_g1627_n
  (
    .dout(g1627_n),
    .din1(g1474_p),
    .din2(g1477_p_spl_)
  );


  orX
  g_g1628_n
  (
    .dout(g1628_n),
    .din1(g1454_n_spl_),
    .din2(g1476_p_spl_)
  );


  andX
  g_g1629_p
  (
    .dout(g1629_p),
    .din1(g1401_n_spl_),
    .din2(g1515_p_spl_)
  );


  andX
  g_g1630_p
  (
    .dout(g1630_p),
    .din1(g1402_n_spl_),
    .din2(g1577_p_spl_)
  );


  andX
  g_g1631_p
  (
    .dout(g1631_p),
    .din1(g1403_n_spl_),
    .din2(g1593_p_spl_)
  );


  orX
  g_g1632_n
  (
    .dout(g1632_n),
    .din1(g1613_n),
    .din2(g1615_p)
  );


  andX
  g_g1633_p
  (
    .dout(g1633_p),
    .din1(g1616_n_spl_),
    .din2(g1632_n)
  );


  orX
  g_g1634_n
  (
    .dout(g1634_n),
    .din1(g1622_n),
    .din2(g1624_p)
  );


  andX
  g_g1635_p
  (
    .dout(g1635_p),
    .din1(g1625_n_spl_),
    .din2(g1634_n)
  );


  orX
  g_g1636_n
  (
    .dout(g1636_n),
    .din1(g1435_n),
    .din2(g1437_p)
  );


  andX
  g_g1637_p
  (
    .dout(g1637_p),
    .din1(g1438_n_spl_),
    .din2(g1636_n)
  );


  orX
  g_g1638_n
  (
    .dout(g1638_n),
    .din1(g1439_n),
    .din2(g1441_p)
  );


  andX
  g_g1639_p
  (
    .dout(g1639_p),
    .din1(g1442_n_spl_),
    .din2(g1638_n)
  );


  orX
  g_g1640_n
  (
    .dout(g1640_n),
    .din1(g1443_n),
    .din2(g1445_p)
  );


  andX
  g_g1641_p
  (
    .dout(g1641_p),
    .din1(g1446_n_spl_),
    .din2(g1640_n)
  );


  orX
  g_g1642_n
  (
    .dout(g1642_n),
    .din1(g1447_n),
    .din2(g1449_p)
  );


  andX
  g_g1643_p
  (
    .dout(g1643_p),
    .din1(g1450_n_spl_),
    .din2(g1642_n)
  );


  orX
  g_g1644_n
  (
    .dout(g1644_n),
    .din1(g1451_n),
    .din2(g1452_n)
  );


  andX
  g_g1645_p
  (
    .dout(g1645_p),
    .din1(g1453_n_spl_),
    .din2(g1644_n)
  );


  orX
  g_g1646_n
  (
    .dout(g1646_n),
    .din1(g1478_n),
    .din2(g1488_p)
  );


  andX
  g_g1647_p
  (
    .dout(g1647_p),
    .din1(g1489_n_spl_),
    .din2(g1646_n)
  );


  orX
  g_g1648_n
  (
    .dout(g1648_n),
    .din1(g1490_n),
    .din2(g1500_p)
  );


  andX
  g_g1649_p
  (
    .dout(g1649_p),
    .din1(g1501_n_spl_),
    .din2(g1648_n)
  );


  orX
  g_g1650_n
  (
    .dout(g1650_n),
    .din1(g1502_n),
    .din2(g1512_p)
  );


  andX
  g_g1651_p
  (
    .dout(g1651_p),
    .din1(g1513_n_spl_),
    .din2(g1650_n)
  );


  orX
  g_g1652_n
  (
    .dout(g1652_n),
    .din1(g1575_p),
    .din2(g1630_p_spl_)
  );


  andX
  g_g1653_p
  (
    .dout(g1653_p),
    .din1(ffc_12_p_spl_000),
    .din2(ffc_195_p_spl_1)
  );


  orX
  g_g1653_n
  (
    .dout(g1653_n),
    .din1(ffc_12_n_spl_001),
    .din2(ffc_195_n_spl_1)
  );


  andX
  g_g1654_p
  (
    .dout(g1654_p),
    .din1(g1569_n_spl_),
    .din2(g1572_n_spl_)
  );


  orX
  g_g1654_n
  (
    .dout(g1654_n),
    .din1(g1569_p_spl_),
    .din2(g1572_p_spl_)
  );


  andX
  g_g1655_p
  (
    .dout(g1655_p),
    .din1(ffc_11_p_spl_011),
    .din2(ffc_180_p_spl_0)
  );


  orX
  g_g1655_n
  (
    .dout(g1655_n),
    .din1(ffc_11_n_spl_011),
    .din2(ffc_180_n_spl_1)
  );


  andX
  g_g1656_p
  (
    .dout(g1656_p),
    .din1(g1563_n_spl_),
    .din2(g1566_n_spl_)
  );


  orX
  g_g1656_n
  (
    .dout(g1656_n),
    .din1(g1563_p_spl_),
    .din2(g1566_p_spl_)
  );


  andX
  g_g1657_p
  (
    .dout(g1657_p),
    .din1(ffc_10_p_spl_100),
    .din2(ffc_181_p_spl_00)
  );


  orX
  g_g1657_n
  (
    .dout(g1657_n),
    .din1(ffc_10_n_spl_100),
    .din2(ffc_181_n_spl_0)
  );


  andX
  g_g1658_p
  (
    .dout(g1658_p),
    .din1(g1557_n_spl_),
    .din2(g1560_n_spl_)
  );


  orX
  g_g1658_n
  (
    .dout(g1658_n),
    .din1(g1557_p_spl_),
    .din2(g1560_p_spl_)
  );


  andX
  g_g1659_p
  (
    .dout(g1659_p),
    .din1(ffc_9_p_spl_101),
    .din2(ffc_182_p_spl_00)
  );


  orX
  g_g1659_n
  (
    .dout(g1659_n),
    .din1(ffc_9_n_spl_101),
    .din2(ffc_182_n_spl_0)
  );


  andX
  g_g1660_p
  (
    .dout(g1660_p),
    .din1(ffc_314_p),
    .din2(g1554_n_spl_)
  );


  orX
  g_g1660_n
  (
    .dout(g1660_n),
    .din1(ffc_314_n),
    .din2(g1554_p_spl_)
  );


  andX
  g_g1661_p
  (
    .dout(g1661_p),
    .din1(ffc_329_n_spl_),
    .din2(ffc_346_p_spl_)
  );


  orX
  g_g1661_n
  (
    .dout(g1661_n),
    .din1(ffc_329_p_spl_),
    .din2(ffc_346_n_spl_)
  );


  andX
  g_g1662_p
  (
    .dout(g1662_p),
    .din1(ffc_329_p_spl_),
    .din2(ffc_346_n_spl_)
  );


  orX
  g_g1662_n
  (
    .dout(g1662_n),
    .din1(ffc_329_n_spl_),
    .din2(ffc_346_p_spl_)
  );


  andX
  g_g1663_p
  (
    .dout(g1663_p),
    .din1(g1661_n_spl_),
    .din2(g1662_n)
  );


  orX
  g_g1663_n
  (
    .dout(g1663_n),
    .din1(g1661_p_spl_),
    .din2(g1662_p)
  );


  andX
  g_g1664_p
  (
    .dout(g1664_p),
    .din1(g1660_n_spl_),
    .din2(g1663_p_spl_)
  );


  orX
  g_g1664_n
  (
    .dout(g1664_n),
    .din1(g1660_p_spl_),
    .din2(g1663_n_spl_)
  );


  andX
  g_g1665_p
  (
    .dout(g1665_p),
    .din1(g1660_p_spl_),
    .din2(g1663_n_spl_)
  );


  orX
  g_g1665_n
  (
    .dout(g1665_n),
    .din1(g1660_n_spl_),
    .din2(g1663_p_spl_)
  );


  andX
  g_g1666_p
  (
    .dout(g1666_p),
    .din1(g1664_n_spl_),
    .din2(g1665_n)
  );


  orX
  g_g1666_n
  (
    .dout(g1666_n),
    .din1(g1664_p_spl_),
    .din2(g1665_p)
  );


  andX
  g_g1667_p
  (
    .dout(g1667_p),
    .din1(g1659_n_spl_),
    .din2(g1666_p_spl_)
  );


  orX
  g_g1667_n
  (
    .dout(g1667_n),
    .din1(g1659_p_spl_),
    .din2(g1666_n_spl_)
  );


  andX
  g_g1668_p
  (
    .dout(g1668_p),
    .din1(g1659_p_spl_),
    .din2(g1666_n_spl_)
  );


  orX
  g_g1668_n
  (
    .dout(g1668_n),
    .din1(g1659_n_spl_),
    .din2(g1666_p_spl_)
  );


  andX
  g_g1669_p
  (
    .dout(g1669_p),
    .din1(g1667_n_spl_),
    .din2(g1668_n)
  );


  orX
  g_g1669_n
  (
    .dout(g1669_n),
    .din1(g1667_p_spl_),
    .din2(g1668_p)
  );


  andX
  g_g1670_p
  (
    .dout(g1670_p),
    .din1(g1658_n_spl_),
    .din2(g1669_p_spl_)
  );


  orX
  g_g1670_n
  (
    .dout(g1670_n),
    .din1(g1658_p_spl_),
    .din2(g1669_n_spl_)
  );


  andX
  g_g1671_p
  (
    .dout(g1671_p),
    .din1(g1658_p_spl_),
    .din2(g1669_n_spl_)
  );


  orX
  g_g1671_n
  (
    .dout(g1671_n),
    .din1(g1658_n_spl_),
    .din2(g1669_p_spl_)
  );


  andX
  g_g1672_p
  (
    .dout(g1672_p),
    .din1(g1670_n_spl_),
    .din2(g1671_n)
  );


  orX
  g_g1672_n
  (
    .dout(g1672_n),
    .din1(g1670_p_spl_),
    .din2(g1671_p)
  );


  andX
  g_g1673_p
  (
    .dout(g1673_p),
    .din1(g1657_n_spl_),
    .din2(g1672_p_spl_)
  );


  orX
  g_g1673_n
  (
    .dout(g1673_n),
    .din1(g1657_p_spl_),
    .din2(g1672_n_spl_)
  );


  andX
  g_g1674_p
  (
    .dout(g1674_p),
    .din1(g1657_p_spl_),
    .din2(g1672_n_spl_)
  );


  orX
  g_g1674_n
  (
    .dout(g1674_n),
    .din1(g1657_n_spl_),
    .din2(g1672_p_spl_)
  );


  andX
  g_g1675_p
  (
    .dout(g1675_p),
    .din1(g1673_n_spl_),
    .din2(g1674_n)
  );


  orX
  g_g1675_n
  (
    .dout(g1675_n),
    .din1(g1673_p_spl_),
    .din2(g1674_p)
  );


  andX
  g_g1676_p
  (
    .dout(g1676_p),
    .din1(g1656_n_spl_),
    .din2(g1675_p_spl_)
  );


  orX
  g_g1676_n
  (
    .dout(g1676_n),
    .din1(g1656_p_spl_),
    .din2(g1675_n_spl_)
  );


  andX
  g_g1677_p
  (
    .dout(g1677_p),
    .din1(g1656_p_spl_),
    .din2(g1675_n_spl_)
  );


  orX
  g_g1677_n
  (
    .dout(g1677_n),
    .din1(g1656_n_spl_),
    .din2(g1675_p_spl_)
  );


  andX
  g_g1678_p
  (
    .dout(g1678_p),
    .din1(g1676_n_spl_),
    .din2(g1677_n)
  );


  orX
  g_g1678_n
  (
    .dout(g1678_n),
    .din1(g1676_p_spl_),
    .din2(g1677_p)
  );


  andX
  g_g1679_p
  (
    .dout(g1679_p),
    .din1(g1655_n_spl_),
    .din2(g1678_p_spl_)
  );


  orX
  g_g1679_n
  (
    .dout(g1679_n),
    .din1(g1655_p_spl_),
    .din2(g1678_n_spl_)
  );


  andX
  g_g1680_p
  (
    .dout(g1680_p),
    .din1(g1655_p_spl_),
    .din2(g1678_n_spl_)
  );


  orX
  g_g1680_n
  (
    .dout(g1680_n),
    .din1(g1655_n_spl_),
    .din2(g1678_p_spl_)
  );


  andX
  g_g1681_p
  (
    .dout(g1681_p),
    .din1(g1679_n_spl_),
    .din2(g1680_n)
  );


  orX
  g_g1681_n
  (
    .dout(g1681_n),
    .din1(g1679_p_spl_),
    .din2(g1680_p)
  );


  andX
  g_g1682_p
  (
    .dout(g1682_p),
    .din1(g1654_n_spl_),
    .din2(g1681_p_spl_)
  );


  orX
  g_g1682_n
  (
    .dout(g1682_n),
    .din1(g1654_p_spl_),
    .din2(g1681_n_spl_)
  );


  andX
  g_g1683_p
  (
    .dout(g1683_p),
    .din1(g1654_p_spl_),
    .din2(g1681_n_spl_)
  );


  orX
  g_g1683_n
  (
    .dout(g1683_n),
    .din1(g1654_n_spl_),
    .din2(g1681_p_spl_)
  );


  andX
  g_g1684_p
  (
    .dout(g1684_p),
    .din1(g1682_n_spl_),
    .din2(g1683_n)
  );


  orX
  g_g1684_n
  (
    .dout(g1684_n),
    .din1(g1682_p),
    .din2(g1683_p)
  );


  orX
  g_g1685_n
  (
    .dout(g1685_n),
    .din1(g1653_p),
    .din2(g1684_n)
  );


  orX
  g_g1686_n
  (
    .dout(g1686_n),
    .din1(g1653_n),
    .din2(g1684_p)
  );


  andX
  g_g1687_p
  (
    .dout(g1687_p),
    .din1(g1685_n_spl_),
    .din2(g1686_n)
  );


  orX
  g_g1688_n
  (
    .dout(g1688_n),
    .din1(ffc_12_n_spl_001),
    .din2(ffc_188_n_spl_1)
  );


  orX
  g_g1689_n
  (
    .dout(g1689_n),
    .din1(g1535_n),
    .din2(g1545_p)
  );


  andX
  g_g1690_p
  (
    .dout(g1690_p),
    .din1(g1546_n_spl_),
    .din2(g1689_n)
  );


  andX
  g_g1691_p
  (
    .dout(g1691_p),
    .din1(g1688_n_spl_),
    .din2(g1690_p_spl_)
  );


  orX
  g_g1692_n
  (
    .dout(g1692_n),
    .din1(g1688_n_spl_),
    .din2(g1690_p_spl_)
  );


  orX
  g_g1693_n
  (
    .dout(g1693_n),
    .din1(ffc_11_n_spl_011),
    .din2(ffc_191_n_spl_)
  );


  orX
  g_g1694_n
  (
    .dout(g1694_n),
    .din1(g1524_n),
    .din2(g1533_p)
  );


  andX
  g_g1695_p
  (
    .dout(g1695_p),
    .din1(g1534_n_spl_),
    .din2(g1694_n)
  );


  andX
  g_g1696_p
  (
    .dout(g1696_p),
    .din1(g1693_n_spl_),
    .din2(g1695_p_spl_)
  );


  orX
  g_g1697_n
  (
    .dout(g1697_n),
    .din1(g1693_n_spl_),
    .din2(g1695_p_spl_)
  );


  orX
  g_g1698_n
  (
    .dout(g1698_n),
    .din1(ffc_10_n_spl_101),
    .din2(ffc_193_n_spl_)
  );


  orX
  g_g1699_n
  (
    .dout(g1699_n),
    .din1(g1528_p_spl_),
    .din2(g1531_p_spl_)
  );


  andX
  g_g1700_p
  (
    .dout(g1700_p),
    .din1(g1698_n_spl_),
    .din2(g1699_n_spl_)
  );


  orX
  g_g1701_n
  (
    .dout(g1701_n),
    .din1(g1698_n_spl_),
    .din2(g1699_n_spl_)
  );


  orX
  g_g1702_n
  (
    .dout(g1702_n),
    .din1(g1540_p_spl_),
    .din2(g1543_p_spl_)
  );


  orX
  g_g1703_n
  (
    .dout(g1703_n),
    .din1(g1520_n),
    .din2(g1522_p)
  );


  andX
  g_g1704_p
  (
    .dout(g1704_p),
    .din1(g1523_n_spl_),
    .din2(g1703_n)
  );


  andX
  g_g1705_p
  (
    .dout(g1705_p),
    .din1(g1702_n_spl_),
    .din2(g1704_p_spl_)
  );


  orX
  g_g1706_n
  (
    .dout(g1706_n),
    .din1(g1702_n_spl_),
    .din2(g1704_p_spl_)
  );


  andX
  g_g1707_p
  (
    .dout(g1707_p),
    .din1(g1676_n_spl_),
    .din2(g1679_n_spl_)
  );


  orX
  g_g1707_n
  (
    .dout(g1707_n),
    .din1(g1676_p_spl_),
    .din2(g1679_p_spl_)
  );


  andX
  g_g1708_p
  (
    .dout(g1708_p),
    .din1(ffc_11_p_spl_011),
    .din2(ffc_181_p_spl_0)
  );


  orX
  g_g1708_n
  (
    .dout(g1708_n),
    .din1(ffc_11_n_spl_100),
    .din2(ffc_181_n_spl_1)
  );


  andX
  g_g1709_p
  (
    .dout(g1709_p),
    .din1(g1670_n_spl_),
    .din2(g1673_n_spl_)
  );


  orX
  g_g1709_n
  (
    .dout(g1709_n),
    .din1(g1670_p_spl_),
    .din2(g1673_p_spl_)
  );


  andX
  g_g1710_p
  (
    .dout(g1710_p),
    .din1(ffc_10_p_spl_101),
    .din2(ffc_182_p_spl_00)
  );


  orX
  g_g1710_n
  (
    .dout(g1710_n),
    .din1(ffc_10_n_spl_101),
    .din2(ffc_182_n_spl_0)
  );


  andX
  g_g1711_p
  (
    .dout(g1711_p),
    .din1(g1664_n_spl_),
    .din2(g1667_n_spl_)
  );


  orX
  g_g1711_n
  (
    .dout(g1711_n),
    .din1(g1664_p_spl_),
    .din2(g1667_p_spl_)
  );


  andX
  g_g1712_p
  (
    .dout(g1712_p),
    .din1(ffc_9_p_spl_110),
    .din2(ffc_183_p_spl_00)
  );


  orX
  g_g1712_n
  (
    .dout(g1712_n),
    .din1(ffc_9_n_spl_110),
    .din2(ffc_183_n_spl_0)
  );


  andX
  g_g1713_p
  (
    .dout(g1713_p),
    .din1(ffc_315_p),
    .din2(g1661_n_spl_)
  );


  orX
  g_g1713_n
  (
    .dout(g1713_n),
    .din1(ffc_315_n),
    .din2(g1661_p_spl_)
  );


  andX
  g_g1714_p
  (
    .dout(g1714_p),
    .din1(ffc_330_n_spl_),
    .din2(ffc_347_p_spl_)
  );


  orX
  g_g1714_n
  (
    .dout(g1714_n),
    .din1(ffc_330_p_spl_),
    .din2(ffc_347_n_spl_)
  );


  andX
  g_g1715_p
  (
    .dout(g1715_p),
    .din1(ffc_330_p_spl_),
    .din2(ffc_347_n_spl_)
  );


  orX
  g_g1715_n
  (
    .dout(g1715_n),
    .din1(ffc_330_n_spl_),
    .din2(ffc_347_p_spl_)
  );


  andX
  g_g1716_p
  (
    .dout(g1716_p),
    .din1(g1714_n_spl_),
    .din2(g1715_n)
  );


  orX
  g_g1716_n
  (
    .dout(g1716_n),
    .din1(g1714_p_spl_),
    .din2(g1715_p)
  );


  andX
  g_g1717_p
  (
    .dout(g1717_p),
    .din1(g1713_n_spl_),
    .din2(g1716_p_spl_)
  );


  orX
  g_g1717_n
  (
    .dout(g1717_n),
    .din1(g1713_p_spl_),
    .din2(g1716_n_spl_)
  );


  andX
  g_g1718_p
  (
    .dout(g1718_p),
    .din1(g1713_p_spl_),
    .din2(g1716_n_spl_)
  );


  orX
  g_g1718_n
  (
    .dout(g1718_n),
    .din1(g1713_n_spl_),
    .din2(g1716_p_spl_)
  );


  andX
  g_g1719_p
  (
    .dout(g1719_p),
    .din1(g1717_n_spl_),
    .din2(g1718_n)
  );


  orX
  g_g1719_n
  (
    .dout(g1719_n),
    .din1(g1717_p_spl_),
    .din2(g1718_p)
  );


  andX
  g_g1720_p
  (
    .dout(g1720_p),
    .din1(g1712_n_spl_),
    .din2(g1719_p_spl_)
  );


  orX
  g_g1720_n
  (
    .dout(g1720_n),
    .din1(g1712_p_spl_),
    .din2(g1719_n_spl_)
  );


  andX
  g_g1721_p
  (
    .dout(g1721_p),
    .din1(g1712_p_spl_),
    .din2(g1719_n_spl_)
  );


  orX
  g_g1721_n
  (
    .dout(g1721_n),
    .din1(g1712_n_spl_),
    .din2(g1719_p_spl_)
  );


  andX
  g_g1722_p
  (
    .dout(g1722_p),
    .din1(g1720_n_spl_),
    .din2(g1721_n)
  );


  orX
  g_g1722_n
  (
    .dout(g1722_n),
    .din1(g1720_p_spl_),
    .din2(g1721_p)
  );


  andX
  g_g1723_p
  (
    .dout(g1723_p),
    .din1(g1711_n_spl_),
    .din2(g1722_p_spl_)
  );


  orX
  g_g1723_n
  (
    .dout(g1723_n),
    .din1(g1711_p_spl_),
    .din2(g1722_n_spl_)
  );


  andX
  g_g1724_p
  (
    .dout(g1724_p),
    .din1(g1711_p_spl_),
    .din2(g1722_n_spl_)
  );


  orX
  g_g1724_n
  (
    .dout(g1724_n),
    .din1(g1711_n_spl_),
    .din2(g1722_p_spl_)
  );


  andX
  g_g1725_p
  (
    .dout(g1725_p),
    .din1(g1723_n_spl_),
    .din2(g1724_n)
  );


  orX
  g_g1725_n
  (
    .dout(g1725_n),
    .din1(g1723_p_spl_),
    .din2(g1724_p)
  );


  andX
  g_g1726_p
  (
    .dout(g1726_p),
    .din1(g1710_n_spl_),
    .din2(g1725_p_spl_)
  );


  orX
  g_g1726_n
  (
    .dout(g1726_n),
    .din1(g1710_p_spl_),
    .din2(g1725_n_spl_)
  );


  andX
  g_g1727_p
  (
    .dout(g1727_p),
    .din1(g1710_p_spl_),
    .din2(g1725_n_spl_)
  );


  orX
  g_g1727_n
  (
    .dout(g1727_n),
    .din1(g1710_n_spl_),
    .din2(g1725_p_spl_)
  );


  andX
  g_g1728_p
  (
    .dout(g1728_p),
    .din1(g1726_n_spl_),
    .din2(g1727_n)
  );


  orX
  g_g1728_n
  (
    .dout(g1728_n),
    .din1(g1726_p_spl_),
    .din2(g1727_p)
  );


  andX
  g_g1729_p
  (
    .dout(g1729_p),
    .din1(g1709_n_spl_),
    .din2(g1728_p_spl_)
  );


  orX
  g_g1729_n
  (
    .dout(g1729_n),
    .din1(g1709_p_spl_),
    .din2(g1728_n_spl_)
  );


  andX
  g_g1730_p
  (
    .dout(g1730_p),
    .din1(g1709_p_spl_),
    .din2(g1728_n_spl_)
  );


  orX
  g_g1730_n
  (
    .dout(g1730_n),
    .din1(g1709_n_spl_),
    .din2(g1728_p_spl_)
  );


  andX
  g_g1731_p
  (
    .dout(g1731_p),
    .din1(g1729_n_spl_),
    .din2(g1730_n)
  );


  orX
  g_g1731_n
  (
    .dout(g1731_n),
    .din1(g1729_p_spl_),
    .din2(g1730_p)
  );


  andX
  g_g1732_p
  (
    .dout(g1732_p),
    .din1(g1708_n_spl_),
    .din2(g1731_p_spl_)
  );


  orX
  g_g1732_n
  (
    .dout(g1732_n),
    .din1(g1708_p_spl_),
    .din2(g1731_n_spl_)
  );


  andX
  g_g1733_p
  (
    .dout(g1733_p),
    .din1(g1708_p_spl_),
    .din2(g1731_n_spl_)
  );


  orX
  g_g1733_n
  (
    .dout(g1733_n),
    .din1(g1708_n_spl_),
    .din2(g1731_p_spl_)
  );


  andX
  g_g1734_p
  (
    .dout(g1734_p),
    .din1(g1732_n_spl_),
    .din2(g1733_n)
  );


  orX
  g_g1734_n
  (
    .dout(g1734_n),
    .din1(g1732_p_spl_),
    .din2(g1733_p)
  );


  andX
  g_g1735_p
  (
    .dout(g1735_p),
    .din1(g1707_n_spl_),
    .din2(g1734_p_spl_)
  );


  orX
  g_g1735_n
  (
    .dout(g1735_n),
    .din1(g1707_p_spl_),
    .din2(g1734_n_spl_)
  );


  andX
  g_g1736_p
  (
    .dout(g1736_p),
    .din1(ffc_12_p_spl_001),
    .din2(ffc_180_p_spl_1)
  );


  orX
  g_g1736_n
  (
    .dout(g1736_n),
    .din1(ffc_12_n_spl_010),
    .din2(ffc_180_n_spl_1)
  );


  andX
  g_g1737_p
  (
    .dout(g1737_p),
    .din1(g1707_p_spl_),
    .din2(g1734_n_spl_)
  );


  orX
  g_g1737_n
  (
    .dout(g1737_n),
    .din1(g1707_n_spl_),
    .din2(g1734_p_spl_)
  );


  andX
  g_g1738_p
  (
    .dout(g1738_p),
    .din1(g1735_n),
    .din2(g1737_n)
  );


  orX
  g_g1738_n
  (
    .dout(g1738_n),
    .din1(g1735_p_spl_),
    .din2(g1737_p)
  );


  andX
  g_g1739_p
  (
    .dout(g1739_p),
    .din1(g1736_n),
    .din2(g1738_p)
  );


  orX
  g_g1740_n
  (
    .dout(g1740_n),
    .din1(g1735_p_spl_),
    .din2(g1739_p_spl_)
  );


  andX
  g_g1741_p
  (
    .dout(g1741_p),
    .din1(ffc_12_p_spl_001),
    .din2(ffc_181_p_spl_1)
  );


  orX
  g_g1741_n
  (
    .dout(g1741_n),
    .din1(ffc_12_n_spl_010),
    .din2(ffc_181_n_spl_1)
  );


  andX
  g_g1742_p
  (
    .dout(g1742_p),
    .din1(g1729_n_spl_),
    .din2(g1732_n_spl_)
  );


  orX
  g_g1742_n
  (
    .dout(g1742_n),
    .din1(g1729_p_spl_),
    .din2(g1732_p_spl_)
  );


  andX
  g_g1743_p
  (
    .dout(g1743_p),
    .din1(ffc_11_p_spl_100),
    .din2(ffc_182_p_spl_0)
  );


  orX
  g_g1743_n
  (
    .dout(g1743_n),
    .din1(ffc_11_n_spl_100),
    .din2(ffc_182_n_spl_1)
  );


  andX
  g_g1744_p
  (
    .dout(g1744_p),
    .din1(g1723_n_spl_),
    .din2(g1726_n_spl_)
  );


  orX
  g_g1744_n
  (
    .dout(g1744_n),
    .din1(g1723_p_spl_),
    .din2(g1726_p_spl_)
  );


  andX
  g_g1745_p
  (
    .dout(g1745_p),
    .din1(ffc_10_p_spl_101),
    .din2(ffc_183_p_spl_00)
  );


  orX
  g_g1745_n
  (
    .dout(g1745_n),
    .din1(ffc_10_n_spl_110),
    .din2(ffc_183_n_spl_0)
  );


  andX
  g_g1746_p
  (
    .dout(g1746_p),
    .din1(g1717_n_spl_),
    .din2(g1720_n_spl_)
  );


  orX
  g_g1746_n
  (
    .dout(g1746_n),
    .din1(g1717_p_spl_),
    .din2(g1720_p_spl_)
  );


  andX
  g_g1747_p
  (
    .dout(g1747_p),
    .din1(ffc_9_p_spl_110),
    .din2(ffc_184_p_spl_00)
  );


  orX
  g_g1747_n
  (
    .dout(g1747_n),
    .din1(ffc_9_n_spl_110),
    .din2(ffc_184_n_spl_0)
  );


  andX
  g_g1748_p
  (
    .dout(g1748_p),
    .din1(ffc_316_p),
    .din2(g1714_n_spl_)
  );


  orX
  g_g1748_n
  (
    .dout(g1748_n),
    .din1(ffc_316_n),
    .din2(g1714_p_spl_)
  );


  andX
  g_g1749_p
  (
    .dout(g1749_p),
    .din1(ffc_331_n_spl_),
    .din2(ffc_348_p_spl_)
  );


  orX
  g_g1749_n
  (
    .dout(g1749_n),
    .din1(ffc_331_p_spl_),
    .din2(ffc_348_n_spl_)
  );


  andX
  g_g1750_p
  (
    .dout(g1750_p),
    .din1(ffc_331_p_spl_),
    .din2(ffc_348_n_spl_)
  );


  orX
  g_g1750_n
  (
    .dout(g1750_n),
    .din1(ffc_331_n_spl_),
    .din2(ffc_348_p_spl_)
  );


  andX
  g_g1751_p
  (
    .dout(g1751_p),
    .din1(g1749_n_spl_),
    .din2(g1750_n)
  );


  orX
  g_g1751_n
  (
    .dout(g1751_n),
    .din1(g1749_p_spl_),
    .din2(g1750_p)
  );


  andX
  g_g1752_p
  (
    .dout(g1752_p),
    .din1(g1748_n_spl_),
    .din2(g1751_p_spl_)
  );


  orX
  g_g1752_n
  (
    .dout(g1752_n),
    .din1(g1748_p_spl_),
    .din2(g1751_n_spl_)
  );


  andX
  g_g1753_p
  (
    .dout(g1753_p),
    .din1(g1748_p_spl_),
    .din2(g1751_n_spl_)
  );


  orX
  g_g1753_n
  (
    .dout(g1753_n),
    .din1(g1748_n_spl_),
    .din2(g1751_p_spl_)
  );


  andX
  g_g1754_p
  (
    .dout(g1754_p),
    .din1(g1752_n_spl_),
    .din2(g1753_n)
  );


  orX
  g_g1754_n
  (
    .dout(g1754_n),
    .din1(g1752_p_spl_),
    .din2(g1753_p)
  );


  andX
  g_g1755_p
  (
    .dout(g1755_p),
    .din1(g1747_n_spl_),
    .din2(g1754_p_spl_)
  );


  orX
  g_g1755_n
  (
    .dout(g1755_n),
    .din1(g1747_p_spl_),
    .din2(g1754_n_spl_)
  );


  andX
  g_g1756_p
  (
    .dout(g1756_p),
    .din1(g1747_p_spl_),
    .din2(g1754_n_spl_)
  );


  orX
  g_g1756_n
  (
    .dout(g1756_n),
    .din1(g1747_n_spl_),
    .din2(g1754_p_spl_)
  );


  andX
  g_g1757_p
  (
    .dout(g1757_p),
    .din1(g1755_n_spl_),
    .din2(g1756_n)
  );


  orX
  g_g1757_n
  (
    .dout(g1757_n),
    .din1(g1755_p_spl_),
    .din2(g1756_p)
  );


  andX
  g_g1758_p
  (
    .dout(g1758_p),
    .din1(g1746_n_spl_),
    .din2(g1757_p_spl_)
  );


  orX
  g_g1758_n
  (
    .dout(g1758_n),
    .din1(g1746_p_spl_),
    .din2(g1757_n_spl_)
  );


  andX
  g_g1759_p
  (
    .dout(g1759_p),
    .din1(g1746_p_spl_),
    .din2(g1757_n_spl_)
  );


  orX
  g_g1759_n
  (
    .dout(g1759_n),
    .din1(g1746_n_spl_),
    .din2(g1757_p_spl_)
  );


  andX
  g_g1760_p
  (
    .dout(g1760_p),
    .din1(g1758_n_spl_),
    .din2(g1759_n)
  );


  orX
  g_g1760_n
  (
    .dout(g1760_n),
    .din1(g1758_p_spl_),
    .din2(g1759_p)
  );


  andX
  g_g1761_p
  (
    .dout(g1761_p),
    .din1(g1745_n_spl_),
    .din2(g1760_p_spl_)
  );


  orX
  g_g1761_n
  (
    .dout(g1761_n),
    .din1(g1745_p_spl_),
    .din2(g1760_n_spl_)
  );


  andX
  g_g1762_p
  (
    .dout(g1762_p),
    .din1(g1745_p_spl_),
    .din2(g1760_n_spl_)
  );


  orX
  g_g1762_n
  (
    .dout(g1762_n),
    .din1(g1745_n_spl_),
    .din2(g1760_p_spl_)
  );


  andX
  g_g1763_p
  (
    .dout(g1763_p),
    .din1(g1761_n_spl_),
    .din2(g1762_n)
  );


  orX
  g_g1763_n
  (
    .dout(g1763_n),
    .din1(g1761_p_spl_),
    .din2(g1762_p)
  );


  andX
  g_g1764_p
  (
    .dout(g1764_p),
    .din1(g1744_n_spl_),
    .din2(g1763_p_spl_)
  );


  orX
  g_g1764_n
  (
    .dout(g1764_n),
    .din1(g1744_p_spl_),
    .din2(g1763_n_spl_)
  );


  andX
  g_g1765_p
  (
    .dout(g1765_p),
    .din1(g1744_p_spl_),
    .din2(g1763_n_spl_)
  );


  orX
  g_g1765_n
  (
    .dout(g1765_n),
    .din1(g1744_n_spl_),
    .din2(g1763_p_spl_)
  );


  andX
  g_g1766_p
  (
    .dout(g1766_p),
    .din1(g1764_n_spl_),
    .din2(g1765_n)
  );


  orX
  g_g1766_n
  (
    .dout(g1766_n),
    .din1(g1764_p_spl_),
    .din2(g1765_p)
  );


  andX
  g_g1767_p
  (
    .dout(g1767_p),
    .din1(g1743_n_spl_),
    .din2(g1766_p_spl_)
  );


  orX
  g_g1767_n
  (
    .dout(g1767_n),
    .din1(g1743_p_spl_),
    .din2(g1766_n_spl_)
  );


  andX
  g_g1768_p
  (
    .dout(g1768_p),
    .din1(g1743_p_spl_),
    .din2(g1766_n_spl_)
  );


  orX
  g_g1768_n
  (
    .dout(g1768_n),
    .din1(g1743_n_spl_),
    .din2(g1766_p_spl_)
  );


  andX
  g_g1769_p
  (
    .dout(g1769_p),
    .din1(g1767_n_spl_),
    .din2(g1768_n)
  );


  orX
  g_g1769_n
  (
    .dout(g1769_n),
    .din1(g1767_p_spl_),
    .din2(g1768_p)
  );


  andX
  g_g1770_p
  (
    .dout(g1770_p),
    .din1(g1742_n_spl_),
    .din2(g1769_p_spl_)
  );


  orX
  g_g1770_n
  (
    .dout(g1770_n),
    .din1(g1742_p_spl_),
    .din2(g1769_n_spl_)
  );


  andX
  g_g1771_p
  (
    .dout(g1771_p),
    .din1(g1742_p_spl_),
    .din2(g1769_n_spl_)
  );


  orX
  g_g1771_n
  (
    .dout(g1771_n),
    .din1(g1742_n_spl_),
    .din2(g1769_p_spl_)
  );


  andX
  g_g1772_p
  (
    .dout(g1772_p),
    .din1(g1770_n),
    .din2(g1771_n)
  );


  orX
  g_g1772_n
  (
    .dout(g1772_n),
    .din1(g1770_p_spl_),
    .din2(g1771_p)
  );


  andX
  g_g1773_p
  (
    .dout(g1773_p),
    .din1(g1741_n_spl_),
    .din2(g1772_p_spl_)
  );


  orX
  g_g1773_n
  (
    .dout(g1773_n),
    .din1(g1741_p),
    .din2(g1772_n)
  );


  orX
  g_g1774_n
  (
    .dout(g1774_n),
    .din1(g1741_n_spl_),
    .din2(g1772_p_spl_)
  );


  andX
  g_g1775_p
  (
    .dout(g1775_p),
    .din1(g1773_n),
    .din2(g1774_n)
  );


  andX
  g_g1776_p
  (
    .dout(g1776_p),
    .din1(g1740_n_spl_),
    .din2(g1775_p_spl_)
  );


  orX
  g_g1777_n
  (
    .dout(g1777_n),
    .din1(g1740_n_spl_),
    .din2(g1775_p_spl_)
  );


  orX
  g_g1778_n
  (
    .dout(g1778_n),
    .din1(g1770_p_spl_),
    .din2(g1773_p)
  );


  andX
  g_g1779_p
  (
    .dout(g1779_p),
    .din1(ffc_12_p_spl_01),
    .din2(ffc_182_p_spl_1)
  );


  orX
  g_g1779_n
  (
    .dout(g1779_n),
    .din1(ffc_12_n_spl_01),
    .din2(ffc_182_n_spl_1)
  );


  andX
  g_g1780_p
  (
    .dout(g1780_p),
    .din1(g1764_n_spl_),
    .din2(g1767_n_spl_)
  );


  orX
  g_g1780_n
  (
    .dout(g1780_n),
    .din1(g1764_p_spl_),
    .din2(g1767_p_spl_)
  );


  andX
  g_g1781_p
  (
    .dout(g1781_p),
    .din1(ffc_11_p_spl_100),
    .din2(ffc_183_p_spl_0)
  );


  orX
  g_g1781_n
  (
    .dout(g1781_n),
    .din1(ffc_11_n_spl_101),
    .din2(ffc_183_n_spl_1)
  );


  andX
  g_g1782_p
  (
    .dout(g1782_p),
    .din1(g1758_n_spl_),
    .din2(g1761_n_spl_)
  );


  orX
  g_g1782_n
  (
    .dout(g1782_n),
    .din1(g1758_p_spl_),
    .din2(g1761_p_spl_)
  );


  andX
  g_g1783_p
  (
    .dout(g1783_p),
    .din1(ffc_10_p_spl_110),
    .din2(ffc_184_p_spl_00)
  );


  orX
  g_g1783_n
  (
    .dout(g1783_n),
    .din1(ffc_10_n_spl_110),
    .din2(ffc_184_n_spl_0)
  );


  andX
  g_g1784_p
  (
    .dout(g1784_p),
    .din1(g1752_n_spl_),
    .din2(g1755_n_spl_)
  );


  orX
  g_g1784_n
  (
    .dout(g1784_n),
    .din1(g1752_p_spl_),
    .din2(g1755_p_spl_)
  );


  andX
  g_g1785_p
  (
    .dout(g1785_p),
    .din1(ffc_9_p_spl_111),
    .din2(ffc_185_p_spl_00)
  );


  orX
  g_g1785_n
  (
    .dout(g1785_n),
    .din1(ffc_9_n_spl_111),
    .din2(ffc_185_n_spl_0)
  );


  andX
  g_g1786_p
  (
    .dout(g1786_p),
    .din1(ffc_317_p),
    .din2(g1749_n_spl_)
  );


  orX
  g_g1786_n
  (
    .dout(g1786_n),
    .din1(ffc_317_n),
    .din2(g1749_p_spl_)
  );


  andX
  g_g1787_p
  (
    .dout(g1787_p),
    .din1(ffc_332_n_spl_),
    .din2(ffc_349_p_spl_)
  );


  orX
  g_g1787_n
  (
    .dout(g1787_n),
    .din1(ffc_332_p_spl_),
    .din2(ffc_349_n_spl_)
  );


  andX
  g_g1788_p
  (
    .dout(g1788_p),
    .din1(ffc_332_p_spl_),
    .din2(ffc_349_n_spl_)
  );


  orX
  g_g1788_n
  (
    .dout(g1788_n),
    .din1(ffc_332_n_spl_),
    .din2(ffc_349_p_spl_)
  );


  andX
  g_g1789_p
  (
    .dout(g1789_p),
    .din1(g1787_n_spl_),
    .din2(g1788_n)
  );


  orX
  g_g1789_n
  (
    .dout(g1789_n),
    .din1(g1787_p_spl_),
    .din2(g1788_p)
  );


  andX
  g_g1790_p
  (
    .dout(g1790_p),
    .din1(g1786_n_spl_),
    .din2(g1789_p_spl_)
  );


  orX
  g_g1790_n
  (
    .dout(g1790_n),
    .din1(g1786_p_spl_),
    .din2(g1789_n_spl_)
  );


  andX
  g_g1791_p
  (
    .dout(g1791_p),
    .din1(g1786_p_spl_),
    .din2(g1789_n_spl_)
  );


  orX
  g_g1791_n
  (
    .dout(g1791_n),
    .din1(g1786_n_spl_),
    .din2(g1789_p_spl_)
  );


  andX
  g_g1792_p
  (
    .dout(g1792_p),
    .din1(g1790_n_spl_),
    .din2(g1791_n)
  );


  orX
  g_g1792_n
  (
    .dout(g1792_n),
    .din1(g1790_p_spl_),
    .din2(g1791_p)
  );


  andX
  g_g1793_p
  (
    .dout(g1793_p),
    .din1(g1785_n_spl_),
    .din2(g1792_p_spl_)
  );


  orX
  g_g1793_n
  (
    .dout(g1793_n),
    .din1(g1785_p_spl_),
    .din2(g1792_n_spl_)
  );


  andX
  g_g1794_p
  (
    .dout(g1794_p),
    .din1(g1785_p_spl_),
    .din2(g1792_n_spl_)
  );


  orX
  g_g1794_n
  (
    .dout(g1794_n),
    .din1(g1785_n_spl_),
    .din2(g1792_p_spl_)
  );


  andX
  g_g1795_p
  (
    .dout(g1795_p),
    .din1(g1793_n_spl_),
    .din2(g1794_n)
  );


  orX
  g_g1795_n
  (
    .dout(g1795_n),
    .din1(g1793_p_spl_),
    .din2(g1794_p)
  );


  andX
  g_g1796_p
  (
    .dout(g1796_p),
    .din1(g1784_n_spl_),
    .din2(g1795_p_spl_)
  );


  orX
  g_g1796_n
  (
    .dout(g1796_n),
    .din1(g1784_p_spl_),
    .din2(g1795_n_spl_)
  );


  andX
  g_g1797_p
  (
    .dout(g1797_p),
    .din1(g1784_p_spl_),
    .din2(g1795_n_spl_)
  );


  orX
  g_g1797_n
  (
    .dout(g1797_n),
    .din1(g1784_n_spl_),
    .din2(g1795_p_spl_)
  );


  andX
  g_g1798_p
  (
    .dout(g1798_p),
    .din1(g1796_n_spl_),
    .din2(g1797_n)
  );


  orX
  g_g1798_n
  (
    .dout(g1798_n),
    .din1(g1796_p_spl_),
    .din2(g1797_p)
  );


  andX
  g_g1799_p
  (
    .dout(g1799_p),
    .din1(g1783_n_spl_),
    .din2(g1798_p_spl_)
  );


  orX
  g_g1799_n
  (
    .dout(g1799_n),
    .din1(g1783_p_spl_),
    .din2(g1798_n_spl_)
  );


  andX
  g_g1800_p
  (
    .dout(g1800_p),
    .din1(g1783_p_spl_),
    .din2(g1798_n_spl_)
  );


  orX
  g_g1800_n
  (
    .dout(g1800_n),
    .din1(g1783_n_spl_),
    .din2(g1798_p_spl_)
  );


  andX
  g_g1801_p
  (
    .dout(g1801_p),
    .din1(g1799_n_spl_),
    .din2(g1800_n)
  );


  orX
  g_g1801_n
  (
    .dout(g1801_n),
    .din1(g1799_p_spl_),
    .din2(g1800_p)
  );


  andX
  g_g1802_p
  (
    .dout(g1802_p),
    .din1(g1782_n_spl_),
    .din2(g1801_p_spl_)
  );


  orX
  g_g1802_n
  (
    .dout(g1802_n),
    .din1(g1782_p_spl_),
    .din2(g1801_n_spl_)
  );


  andX
  g_g1803_p
  (
    .dout(g1803_p),
    .din1(g1782_p_spl_),
    .din2(g1801_n_spl_)
  );


  orX
  g_g1803_n
  (
    .dout(g1803_n),
    .din1(g1782_n_spl_),
    .din2(g1801_p_spl_)
  );


  andX
  g_g1804_p
  (
    .dout(g1804_p),
    .din1(g1802_n_spl_),
    .din2(g1803_n)
  );


  orX
  g_g1804_n
  (
    .dout(g1804_n),
    .din1(g1802_p_spl_),
    .din2(g1803_p)
  );


  andX
  g_g1805_p
  (
    .dout(g1805_p),
    .din1(g1781_n_spl_),
    .din2(g1804_p_spl_)
  );


  orX
  g_g1805_n
  (
    .dout(g1805_n),
    .din1(g1781_p_spl_),
    .din2(g1804_n_spl_)
  );


  andX
  g_g1806_p
  (
    .dout(g1806_p),
    .din1(g1781_p_spl_),
    .din2(g1804_n_spl_)
  );


  orX
  g_g1806_n
  (
    .dout(g1806_n),
    .din1(g1781_n_spl_),
    .din2(g1804_p_spl_)
  );


  andX
  g_g1807_p
  (
    .dout(g1807_p),
    .din1(g1805_n_spl_),
    .din2(g1806_n)
  );


  orX
  g_g1807_n
  (
    .dout(g1807_n),
    .din1(g1805_p_spl_),
    .din2(g1806_p)
  );


  andX
  g_g1808_p
  (
    .dout(g1808_p),
    .din1(g1780_n_spl_),
    .din2(g1807_p_spl_)
  );


  orX
  g_g1808_n
  (
    .dout(g1808_n),
    .din1(g1780_p_spl_),
    .din2(g1807_n_spl_)
  );


  andX
  g_g1809_p
  (
    .dout(g1809_p),
    .din1(g1780_p_spl_),
    .din2(g1807_n_spl_)
  );


  orX
  g_g1809_n
  (
    .dout(g1809_n),
    .din1(g1780_n_spl_),
    .din2(g1807_p_spl_)
  );


  andX
  g_g1810_p
  (
    .dout(g1810_p),
    .din1(g1808_n),
    .din2(g1809_n)
  );


  orX
  g_g1810_n
  (
    .dout(g1810_n),
    .din1(g1808_p_spl_),
    .din2(g1809_p)
  );


  andX
  g_g1811_p
  (
    .dout(g1811_p),
    .din1(g1779_n_spl_),
    .din2(g1810_p_spl_)
  );


  orX
  g_g1811_n
  (
    .dout(g1811_n),
    .din1(g1779_p),
    .din2(g1810_n)
  );


  orX
  g_g1812_n
  (
    .dout(g1812_n),
    .din1(g1779_n_spl_),
    .din2(g1810_p_spl_)
  );


  andX
  g_g1813_p
  (
    .dout(g1813_p),
    .din1(g1811_n),
    .din2(g1812_n)
  );


  andX
  g_g1814_p
  (
    .dout(g1814_p),
    .din1(g1778_n_spl_),
    .din2(g1813_p_spl_)
  );


  orX
  g_g1815_n
  (
    .dout(g1815_n),
    .din1(g1778_n_spl_),
    .din2(g1813_p_spl_)
  );


  orX
  g_g1816_n
  (
    .dout(g1816_n),
    .din1(g1808_p_spl_),
    .din2(g1811_p)
  );


  andX
  g_g1817_p
  (
    .dout(g1817_p),
    .din1(ffc_12_p_spl_01),
    .din2(ffc_183_p_spl_1)
  );


  orX
  g_g1817_n
  (
    .dout(g1817_n),
    .din1(ffc_12_n_spl_10),
    .din2(ffc_183_n_spl_1)
  );


  andX
  g_g1818_p
  (
    .dout(g1818_p),
    .din1(g1802_n_spl_),
    .din2(g1805_n_spl_)
  );


  orX
  g_g1818_n
  (
    .dout(g1818_n),
    .din1(g1802_p_spl_),
    .din2(g1805_p_spl_)
  );


  andX
  g_g1819_p
  (
    .dout(g1819_p),
    .din1(ffc_11_p_spl_101),
    .din2(ffc_184_p_spl_0)
  );


  orX
  g_g1819_n
  (
    .dout(g1819_n),
    .din1(ffc_11_n_spl_101),
    .din2(ffc_184_n_spl_1)
  );


  andX
  g_g1820_p
  (
    .dout(g1820_p),
    .din1(g1796_n_spl_),
    .din2(g1799_n_spl_)
  );


  orX
  g_g1820_n
  (
    .dout(g1820_n),
    .din1(g1796_p_spl_),
    .din2(g1799_p_spl_)
  );


  andX
  g_g1821_p
  (
    .dout(g1821_p),
    .din1(ffc_10_p_spl_110),
    .din2(ffc_185_p_spl_00)
  );


  orX
  g_g1821_n
  (
    .dout(g1821_n),
    .din1(ffc_10_n_spl_111),
    .din2(ffc_185_n_spl_0)
  );


  andX
  g_g1822_p
  (
    .dout(g1822_p),
    .din1(g1790_n_spl_),
    .din2(g1793_n_spl_)
  );


  orX
  g_g1822_n
  (
    .dout(g1822_n),
    .din1(g1790_p_spl_),
    .din2(g1793_p_spl_)
  );


  andX
  g_g1823_p
  (
    .dout(g1823_p),
    .din1(ffc_9_p_spl_111),
    .din2(ffc_186_p_spl_00)
  );


  orX
  g_g1823_n
  (
    .dout(g1823_n),
    .din1(ffc_9_n_spl_111),
    .din2(ffc_186_n_spl_0)
  );


  andX
  g_g1824_p
  (
    .dout(g1824_p),
    .din1(ffc_318_p),
    .din2(g1787_n_spl_)
  );


  orX
  g_g1824_n
  (
    .dout(g1824_n),
    .din1(ffc_318_n),
    .din2(g1787_p_spl_)
  );


  andX
  g_g1825_p
  (
    .dout(g1825_p),
    .din1(ffc_333_p_spl_),
    .din2(ffc_350_n_spl_)
  );


  orX
  g_g1825_n
  (
    .dout(g1825_n),
    .din1(ffc_333_n_spl_),
    .din2(ffc_350_p_spl_)
  );


  andX
  g_g1826_p
  (
    .dout(g1826_p),
    .din1(g1329_n_spl_),
    .din2(g1825_n)
  );


  orX
  g_g1826_n
  (
    .dout(g1826_n),
    .din1(g1329_p_spl_),
    .din2(g1825_p)
  );


  andX
  g_g1827_p
  (
    .dout(g1827_p),
    .din1(g1824_n_spl_),
    .din2(g1826_p_spl_)
  );


  orX
  g_g1827_n
  (
    .dout(g1827_n),
    .din1(g1824_p_spl_),
    .din2(g1826_n_spl_)
  );


  andX
  g_g1828_p
  (
    .dout(g1828_p),
    .din1(g1824_p_spl_),
    .din2(g1826_n_spl_)
  );


  orX
  g_g1828_n
  (
    .dout(g1828_n),
    .din1(g1824_n_spl_),
    .din2(g1826_p_spl_)
  );


  andX
  g_g1829_p
  (
    .dout(g1829_p),
    .din1(g1827_n_spl_),
    .din2(g1828_n)
  );


  orX
  g_g1829_n
  (
    .dout(g1829_n),
    .din1(g1827_p_spl_),
    .din2(g1828_p)
  );


  andX
  g_g1830_p
  (
    .dout(g1830_p),
    .din1(g1823_n_spl_),
    .din2(g1829_p_spl_)
  );


  orX
  g_g1830_n
  (
    .dout(g1830_n),
    .din1(g1823_p_spl_),
    .din2(g1829_n_spl_)
  );


  andX
  g_g1831_p
  (
    .dout(g1831_p),
    .din1(g1823_p_spl_),
    .din2(g1829_n_spl_)
  );


  orX
  g_g1831_n
  (
    .dout(g1831_n),
    .din1(g1823_n_spl_),
    .din2(g1829_p_spl_)
  );


  andX
  g_g1832_p
  (
    .dout(g1832_p),
    .din1(g1830_n_spl_),
    .din2(g1831_n)
  );


  orX
  g_g1832_n
  (
    .dout(g1832_n),
    .din1(g1830_p_spl_),
    .din2(g1831_p)
  );


  andX
  g_g1833_p
  (
    .dout(g1833_p),
    .din1(g1822_n_spl_),
    .din2(g1832_p_spl_)
  );


  orX
  g_g1833_n
  (
    .dout(g1833_n),
    .din1(g1822_p_spl_),
    .din2(g1832_n_spl_)
  );


  andX
  g_g1834_p
  (
    .dout(g1834_p),
    .din1(g1822_p_spl_),
    .din2(g1832_n_spl_)
  );


  orX
  g_g1834_n
  (
    .dout(g1834_n),
    .din1(g1822_n_spl_),
    .din2(g1832_p_spl_)
  );


  andX
  g_g1835_p
  (
    .dout(g1835_p),
    .din1(g1833_n_spl_),
    .din2(g1834_n)
  );


  orX
  g_g1835_n
  (
    .dout(g1835_n),
    .din1(g1833_p_spl_),
    .din2(g1834_p)
  );


  andX
  g_g1836_p
  (
    .dout(g1836_p),
    .din1(g1821_n_spl_),
    .din2(g1835_p_spl_)
  );


  orX
  g_g1836_n
  (
    .dout(g1836_n),
    .din1(g1821_p_spl_),
    .din2(g1835_n_spl_)
  );


  andX
  g_g1837_p
  (
    .dout(g1837_p),
    .din1(g1821_p_spl_),
    .din2(g1835_n_spl_)
  );


  orX
  g_g1837_n
  (
    .dout(g1837_n),
    .din1(g1821_n_spl_),
    .din2(g1835_p_spl_)
  );


  andX
  g_g1838_p
  (
    .dout(g1838_p),
    .din1(g1836_n_spl_),
    .din2(g1837_n)
  );


  orX
  g_g1838_n
  (
    .dout(g1838_n),
    .din1(g1836_p_spl_),
    .din2(g1837_p)
  );


  andX
  g_g1839_p
  (
    .dout(g1839_p),
    .din1(g1820_n_spl_),
    .din2(g1838_p_spl_)
  );


  orX
  g_g1839_n
  (
    .dout(g1839_n),
    .din1(g1820_p_spl_),
    .din2(g1838_n_spl_)
  );


  andX
  g_g1840_p
  (
    .dout(g1840_p),
    .din1(g1820_p_spl_),
    .din2(g1838_n_spl_)
  );


  orX
  g_g1840_n
  (
    .dout(g1840_n),
    .din1(g1820_n_spl_),
    .din2(g1838_p_spl_)
  );


  andX
  g_g1841_p
  (
    .dout(g1841_p),
    .din1(g1839_n_spl_),
    .din2(g1840_n)
  );


  orX
  g_g1841_n
  (
    .dout(g1841_n),
    .din1(g1839_p_spl_),
    .din2(g1840_p)
  );


  andX
  g_g1842_p
  (
    .dout(g1842_p),
    .din1(g1819_n_spl_),
    .din2(g1841_p_spl_)
  );


  orX
  g_g1842_n
  (
    .dout(g1842_n),
    .din1(g1819_p_spl_),
    .din2(g1841_n_spl_)
  );


  andX
  g_g1843_p
  (
    .dout(g1843_p),
    .din1(g1819_p_spl_),
    .din2(g1841_n_spl_)
  );


  orX
  g_g1843_n
  (
    .dout(g1843_n),
    .din1(g1819_n_spl_),
    .din2(g1841_p_spl_)
  );


  andX
  g_g1844_p
  (
    .dout(g1844_p),
    .din1(g1842_n_spl_),
    .din2(g1843_n)
  );


  orX
  g_g1844_n
  (
    .dout(g1844_n),
    .din1(g1842_p_spl_),
    .din2(g1843_p)
  );


  andX
  g_g1845_p
  (
    .dout(g1845_p),
    .din1(g1818_n_spl_),
    .din2(g1844_p_spl_)
  );


  orX
  g_g1845_n
  (
    .dout(g1845_n),
    .din1(g1818_p_spl_),
    .din2(g1844_n_spl_)
  );


  andX
  g_g1846_p
  (
    .dout(g1846_p),
    .din1(g1818_p_spl_),
    .din2(g1844_n_spl_)
  );


  orX
  g_g1846_n
  (
    .dout(g1846_n),
    .din1(g1818_n_spl_),
    .din2(g1844_p_spl_)
  );


  andX
  g_g1847_p
  (
    .dout(g1847_p),
    .din1(g1845_n),
    .din2(g1846_n)
  );


  orX
  g_g1847_n
  (
    .dout(g1847_n),
    .din1(g1845_p_spl_),
    .din2(g1846_p)
  );


  andX
  g_g1848_p
  (
    .dout(g1848_p),
    .din1(g1817_n_spl_),
    .din2(g1847_p_spl_)
  );


  orX
  g_g1848_n
  (
    .dout(g1848_n),
    .din1(g1817_p),
    .din2(g1847_n)
  );


  orX
  g_g1849_n
  (
    .dout(g1849_n),
    .din1(g1817_n_spl_),
    .din2(g1847_p_spl_)
  );


  andX
  g_g1850_p
  (
    .dout(g1850_p),
    .din1(g1848_n),
    .din2(g1849_n)
  );


  andX
  g_g1851_p
  (
    .dout(g1851_p),
    .din1(g1816_n_spl_),
    .din2(g1850_p_spl_)
  );


  orX
  g_g1852_n
  (
    .dout(g1852_n),
    .din1(g1816_n_spl_),
    .din2(g1850_p_spl_)
  );


  orX
  g_g1853_n
  (
    .dout(g1853_n),
    .din1(g1845_p_spl_),
    .din2(g1848_p)
  );


  andX
  g_g1854_p
  (
    .dout(g1854_p),
    .din1(ffc_12_p_spl_10),
    .din2(ffc_184_p_spl_1)
  );


  orX
  g_g1854_n
  (
    .dout(g1854_n),
    .din1(ffc_12_n_spl_10),
    .din2(ffc_184_n_spl_1)
  );


  andX
  g_g1855_p
  (
    .dout(g1855_p),
    .din1(g1839_n_spl_),
    .din2(g1842_n_spl_)
  );


  orX
  g_g1855_n
  (
    .dout(g1855_n),
    .din1(g1839_p_spl_),
    .din2(g1842_p_spl_)
  );


  andX
  g_g1856_p
  (
    .dout(g1856_p),
    .din1(ffc_11_p_spl_101),
    .din2(ffc_185_p_spl_0)
  );


  orX
  g_g1856_n
  (
    .dout(g1856_n),
    .din1(ffc_11_n_spl_11),
    .din2(ffc_185_n_spl_1)
  );


  andX
  g_g1857_p
  (
    .dout(g1857_p),
    .din1(g1833_n_spl_),
    .din2(g1836_n_spl_)
  );


  orX
  g_g1857_n
  (
    .dout(g1857_n),
    .din1(g1833_p_spl_),
    .din2(g1836_p_spl_)
  );


  andX
  g_g1858_p
  (
    .dout(g1858_p),
    .din1(ffc_10_p_spl_11),
    .din2(ffc_186_p_spl_00)
  );


  orX
  g_g1858_n
  (
    .dout(g1858_n),
    .din1(ffc_10_n_spl_111),
    .din2(ffc_186_n_spl_0)
  );


  andX
  g_g1859_p
  (
    .dout(g1859_p),
    .din1(g1827_n_spl_),
    .din2(g1830_n_spl_)
  );


  orX
  g_g1859_n
  (
    .dout(g1859_n),
    .din1(g1827_p_spl_),
    .din2(g1830_p_spl_)
  );


  andX
  g_g1860_p
  (
    .dout(g1860_p),
    .din1(g1335_p_spl_),
    .din2(g1337_n_spl_)
  );


  orX
  g_g1860_n
  (
    .dout(g1860_n),
    .din1(g1335_n_spl_),
    .din2(g1337_p_spl_)
  );


  andX
  g_g1861_p
  (
    .dout(g1861_p),
    .din1(g1338_n_spl_),
    .din2(g1860_n)
  );


  orX
  g_g1861_n
  (
    .dout(g1861_n),
    .din1(g1338_p_spl_),
    .din2(g1860_p)
  );


  andX
  g_g1862_p
  (
    .dout(g1862_p),
    .din1(g1859_n_spl_),
    .din2(g1861_p_spl_)
  );


  orX
  g_g1862_n
  (
    .dout(g1862_n),
    .din1(g1859_p_spl_),
    .din2(g1861_n_spl_)
  );


  andX
  g_g1863_p
  (
    .dout(g1863_p),
    .din1(g1859_p_spl_),
    .din2(g1861_n_spl_)
  );


  orX
  g_g1863_n
  (
    .dout(g1863_n),
    .din1(g1859_n_spl_),
    .din2(g1861_p_spl_)
  );


  andX
  g_g1864_p
  (
    .dout(g1864_p),
    .din1(g1862_n_spl_),
    .din2(g1863_n)
  );


  orX
  g_g1864_n
  (
    .dout(g1864_n),
    .din1(g1862_p_spl_),
    .din2(g1863_p)
  );


  andX
  g_g1865_p
  (
    .dout(g1865_p),
    .din1(g1858_n_spl_),
    .din2(g1864_p_spl_)
  );


  orX
  g_g1865_n
  (
    .dout(g1865_n),
    .din1(g1858_p_spl_),
    .din2(g1864_n_spl_)
  );


  andX
  g_g1866_p
  (
    .dout(g1866_p),
    .din1(g1858_p_spl_),
    .din2(g1864_n_spl_)
  );


  orX
  g_g1866_n
  (
    .dout(g1866_n),
    .din1(g1858_n_spl_),
    .din2(g1864_p_spl_)
  );


  andX
  g_g1867_p
  (
    .dout(g1867_p),
    .din1(g1865_n_spl_),
    .din2(g1866_n)
  );


  orX
  g_g1867_n
  (
    .dout(g1867_n),
    .din1(g1865_p_spl_),
    .din2(g1866_p)
  );


  andX
  g_g1868_p
  (
    .dout(g1868_p),
    .din1(g1857_n_spl_),
    .din2(g1867_p_spl_)
  );


  orX
  g_g1868_n
  (
    .dout(g1868_n),
    .din1(g1857_p_spl_),
    .din2(g1867_n_spl_)
  );


  andX
  g_g1869_p
  (
    .dout(g1869_p),
    .din1(g1857_p_spl_),
    .din2(g1867_n_spl_)
  );


  orX
  g_g1869_n
  (
    .dout(g1869_n),
    .din1(g1857_n_spl_),
    .din2(g1867_p_spl_)
  );


  andX
  g_g1870_p
  (
    .dout(g1870_p),
    .din1(g1868_n_spl_),
    .din2(g1869_n)
  );


  orX
  g_g1870_n
  (
    .dout(g1870_n),
    .din1(g1868_p_spl_),
    .din2(g1869_p)
  );


  andX
  g_g1871_p
  (
    .dout(g1871_p),
    .din1(g1856_n_spl_),
    .din2(g1870_p_spl_)
  );


  orX
  g_g1871_n
  (
    .dout(g1871_n),
    .din1(g1856_p_spl_),
    .din2(g1870_n_spl_)
  );


  andX
  g_g1872_p
  (
    .dout(g1872_p),
    .din1(g1856_p_spl_),
    .din2(g1870_n_spl_)
  );


  orX
  g_g1872_n
  (
    .dout(g1872_n),
    .din1(g1856_n_spl_),
    .din2(g1870_p_spl_)
  );


  andX
  g_g1873_p
  (
    .dout(g1873_p),
    .din1(g1871_n_spl_),
    .din2(g1872_n)
  );


  orX
  g_g1873_n
  (
    .dout(g1873_n),
    .din1(g1871_p_spl_),
    .din2(g1872_p)
  );


  andX
  g_g1874_p
  (
    .dout(g1874_p),
    .din1(g1855_n_spl_),
    .din2(g1873_p_spl_)
  );


  orX
  g_g1874_n
  (
    .dout(g1874_n),
    .din1(g1855_p_spl_),
    .din2(g1873_n_spl_)
  );


  andX
  g_g1875_p
  (
    .dout(g1875_p),
    .din1(g1855_p_spl_),
    .din2(g1873_n_spl_)
  );


  orX
  g_g1875_n
  (
    .dout(g1875_n),
    .din1(g1855_n_spl_),
    .din2(g1873_p_spl_)
  );


  andX
  g_g1876_p
  (
    .dout(g1876_p),
    .din1(g1874_n),
    .din2(g1875_n)
  );


  orX
  g_g1876_n
  (
    .dout(g1876_n),
    .din1(g1874_p_spl_),
    .din2(g1875_p)
  );


  andX
  g_g1877_p
  (
    .dout(g1877_p),
    .din1(g1854_n_spl_),
    .din2(g1876_p_spl_)
  );


  orX
  g_g1877_n
  (
    .dout(g1877_n),
    .din1(g1854_p),
    .din2(g1876_n)
  );


  orX
  g_g1878_n
  (
    .dout(g1878_n),
    .din1(g1854_n_spl_),
    .din2(g1876_p_spl_)
  );


  andX
  g_g1879_p
  (
    .dout(g1879_p),
    .din1(g1877_n),
    .din2(g1878_n)
  );


  andX
  g_g1880_p
  (
    .dout(g1880_p),
    .din1(g1853_n_spl_),
    .din2(g1879_p_spl_)
  );


  orX
  g_g1881_n
  (
    .dout(g1881_n),
    .din1(g1853_n_spl_),
    .din2(g1879_p_spl_)
  );


  orX
  g_g1882_n
  (
    .dout(g1882_n),
    .din1(g1874_p_spl_),
    .din2(g1877_p)
  );


  andX
  g_g1883_p
  (
    .dout(g1883_p),
    .din1(ffc_12_p_spl_10),
    .din2(ffc_185_p_spl_1)
  );


  orX
  g_g1883_n
  (
    .dout(g1883_n),
    .din1(ffc_12_n_spl_11),
    .din2(ffc_185_n_spl_1)
  );


  andX
  g_g1884_p
  (
    .dout(g1884_p),
    .din1(g1868_n_spl_),
    .din2(g1871_n_spl_)
  );


  orX
  g_g1884_n
  (
    .dout(g1884_n),
    .din1(g1868_p_spl_),
    .din2(g1871_p_spl_)
  );


  andX
  g_g1885_p
  (
    .dout(g1885_p),
    .din1(ffc_11_p_spl_11),
    .din2(ffc_186_p_spl_0)
  );


  orX
  g_g1885_n
  (
    .dout(g1885_n),
    .din1(ffc_11_n_spl_11),
    .din2(ffc_186_n_spl_1)
  );


  andX
  g_g1886_p
  (
    .dout(g1886_p),
    .din1(g1862_n_spl_),
    .din2(g1865_n_spl_)
  );


  orX
  g_g1886_n
  (
    .dout(g1886_n),
    .din1(g1862_p_spl_),
    .din2(g1865_p_spl_)
  );


  andX
  g_g1887_p
  (
    .dout(g1887_p),
    .din1(g1352_p_spl_),
    .din2(g1354_n_spl_)
  );


  orX
  g_g1887_n
  (
    .dout(g1887_n),
    .din1(g1352_n_spl_),
    .din2(g1354_p_spl_)
  );


  andX
  g_g1888_p
  (
    .dout(g1888_p),
    .din1(g1355_n_spl_),
    .din2(g1887_n)
  );


  orX
  g_g1888_n
  (
    .dout(g1888_n),
    .din1(g1355_p_spl_),
    .din2(g1887_p)
  );


  andX
  g_g1889_p
  (
    .dout(g1889_p),
    .din1(g1886_n_spl_),
    .din2(g1888_p_spl_)
  );


  orX
  g_g1889_n
  (
    .dout(g1889_n),
    .din1(g1886_p_spl_),
    .din2(g1888_n_spl_)
  );


  andX
  g_g1890_p
  (
    .dout(g1890_p),
    .din1(g1886_p_spl_),
    .din2(g1888_n_spl_)
  );


  orX
  g_g1890_n
  (
    .dout(g1890_n),
    .din1(g1886_n_spl_),
    .din2(g1888_p_spl_)
  );


  andX
  g_g1891_p
  (
    .dout(g1891_p),
    .din1(g1889_n_spl_),
    .din2(g1890_n)
  );


  orX
  g_g1891_n
  (
    .dout(g1891_n),
    .din1(g1889_p_spl_),
    .din2(g1890_p)
  );


  andX
  g_g1892_p
  (
    .dout(g1892_p),
    .din1(g1885_n_spl_),
    .din2(g1891_p_spl_)
  );


  orX
  g_g1892_n
  (
    .dout(g1892_n),
    .din1(g1885_p_spl_),
    .din2(g1891_n_spl_)
  );


  andX
  g_g1893_p
  (
    .dout(g1893_p),
    .din1(g1885_p_spl_),
    .din2(g1891_n_spl_)
  );


  orX
  g_g1893_n
  (
    .dout(g1893_n),
    .din1(g1885_n_spl_),
    .din2(g1891_p_spl_)
  );


  andX
  g_g1894_p
  (
    .dout(g1894_p),
    .din1(g1892_n_spl_),
    .din2(g1893_n)
  );


  orX
  g_g1894_n
  (
    .dout(g1894_n),
    .din1(g1892_p_spl_),
    .din2(g1893_p)
  );


  andX
  g_g1895_p
  (
    .dout(g1895_p),
    .din1(g1884_n_spl_),
    .din2(g1894_p_spl_)
  );


  orX
  g_g1895_n
  (
    .dout(g1895_n),
    .din1(g1884_p_spl_),
    .din2(g1894_n_spl_)
  );


  andX
  g_g1896_p
  (
    .dout(g1896_p),
    .din1(g1884_p_spl_),
    .din2(g1894_n_spl_)
  );


  orX
  g_g1896_n
  (
    .dout(g1896_n),
    .din1(g1884_n_spl_),
    .din2(g1894_p_spl_)
  );


  andX
  g_g1897_p
  (
    .dout(g1897_p),
    .din1(g1895_n),
    .din2(g1896_n)
  );


  orX
  g_g1897_n
  (
    .dout(g1897_n),
    .din1(g1895_p_spl_),
    .din2(g1896_p)
  );


  andX
  g_g1898_p
  (
    .dout(g1898_p),
    .din1(g1883_n_spl_),
    .din2(g1897_p_spl_)
  );


  orX
  g_g1898_n
  (
    .dout(g1898_n),
    .din1(g1883_p),
    .din2(g1897_n)
  );


  orX
  g_g1899_n
  (
    .dout(g1899_n),
    .din1(g1883_n_spl_),
    .din2(g1897_p_spl_)
  );


  andX
  g_g1900_p
  (
    .dout(g1900_p),
    .din1(g1898_n),
    .din2(g1899_n)
  );


  andX
  g_g1901_p
  (
    .dout(g1901_p),
    .din1(g1882_n_spl_),
    .din2(g1900_p_spl_)
  );


  orX
  g_g1902_n
  (
    .dout(g1902_n),
    .din1(g1882_n_spl_),
    .din2(g1900_p_spl_)
  );


  orX
  g_g1903_n
  (
    .dout(g1903_n),
    .din1(g1895_p_spl_),
    .din2(g1898_p)
  );


  andX
  g_g1904_p
  (
    .dout(g1904_p),
    .din1(ffc_12_p_spl_11),
    .din2(ffc_186_p_spl_1)
  );


  orX
  g_g1904_n
  (
    .dout(g1904_n),
    .din1(ffc_12_n_spl_11),
    .din2(ffc_186_n_spl_1)
  );


  andX
  g_g1905_p
  (
    .dout(g1905_p),
    .din1(g1889_n_spl_),
    .din2(g1892_n_spl_)
  );


  orX
  g_g1905_n
  (
    .dout(g1905_n),
    .din1(g1889_p_spl_),
    .din2(g1892_p_spl_)
  );


  andX
  g_g1906_p
  (
    .dout(g1906_p),
    .din1(g1376_p_spl_),
    .din2(g1378_n_spl_)
  );


  orX
  g_g1906_n
  (
    .dout(g1906_n),
    .din1(g1376_n_spl_),
    .din2(g1378_p_spl_)
  );


  andX
  g_g1907_p
  (
    .dout(g1907_p),
    .din1(g1379_n_spl_),
    .din2(g1906_n)
  );


  orX
  g_g1907_n
  (
    .dout(g1907_n),
    .din1(g1379_p_spl_),
    .din2(g1906_p)
  );


  andX
  g_g1908_p
  (
    .dout(g1908_p),
    .din1(g1905_n_spl_),
    .din2(g1907_p_spl_)
  );


  orX
  g_g1908_n
  (
    .dout(g1908_n),
    .din1(g1905_p_spl_),
    .din2(g1907_n_spl_)
  );


  andX
  g_g1909_p
  (
    .dout(g1909_p),
    .din1(g1905_p_spl_),
    .din2(g1907_n_spl_)
  );


  orX
  g_g1909_n
  (
    .dout(g1909_n),
    .din1(g1905_n_spl_),
    .din2(g1907_p_spl_)
  );


  andX
  g_g1910_p
  (
    .dout(g1910_p),
    .din1(g1908_n),
    .din2(g1909_n)
  );


  orX
  g_g1910_n
  (
    .dout(g1910_n),
    .din1(g1908_p_spl_),
    .din2(g1909_p)
  );


  andX
  g_g1911_p
  (
    .dout(g1911_p),
    .din1(g1904_n_spl_),
    .din2(g1910_p_spl_)
  );


  orX
  g_g1911_n
  (
    .dout(g1911_n),
    .din1(g1904_p),
    .din2(g1910_n)
  );


  orX
  g_g1912_n
  (
    .dout(g1912_n),
    .din1(g1904_n_spl_),
    .din2(g1910_p_spl_)
  );


  andX
  g_g1913_p
  (
    .dout(g1913_p),
    .din1(g1911_n),
    .din2(g1912_n)
  );


  andX
  g_g1914_p
  (
    .dout(g1914_p),
    .din1(g1903_n_spl_),
    .din2(g1913_p_spl_)
  );


  orX
  g_g1915_n
  (
    .dout(g1915_n),
    .din1(g1903_n_spl_),
    .din2(g1913_p_spl_)
  );


  orX
  g_g1916_n
  (
    .dout(g1916_n),
    .din1(g1908_p_spl_),
    .din2(g1911_p)
  );


  orX
  g_g1917_n
  (
    .dout(g1917_n),
    .din1(g1516_n),
    .din2(g1518_p)
  );


  andX
  g_g1918_p
  (
    .dout(g1918_p),
    .din1(g1519_n_spl_),
    .din2(g1917_n)
  );


  andX
  g_g1919_p
  (
    .dout(g1919_p),
    .din1(g1916_n_spl_),
    .din2(g1918_p_spl_)
  );


  orX
  g_g1920_n
  (
    .dout(g1920_n),
    .din1(g1916_n_spl_),
    .din2(g1918_p_spl_)
  );


  andX
  g_g1921_p
  (
    .dout(g1921_p),
    .din1(g1682_n_spl_),
    .din2(g1685_n_spl_)
  );


  andX
  g_g1922_p
  (
    .dout(g1922_p),
    .din1(g1736_p),
    .din2(g1738_n)
  );


  orX
  g_g1923_n
  (
    .dout(g1923_n),
    .din1(g1739_p_spl_),
    .din2(g1922_p)
  );


  orX
  g_g1924_n
  (
    .dout(g1924_n),
    .din1(g1921_p_spl_),
    .din2(g1923_n_spl_)
  );


  andX
  g_g1925_p
  (
    .dout(g1925_p),
    .din1(g1921_p_spl_),
    .din2(g1923_n_spl_)
  );


  andX
  g_g1926_p
  (
    .dout(g1926_p),
    .din1(G5_p_spl_00),
    .din2(G17_p_spl_001)
  );


  orX
  g_g1926_n
  (
    .dout(g1926_n),
    .din1(G5_n_spl_0),
    .din2(G17_n_spl_001)
  );


  andX
  g_g1927_p
  (
    .dout(g1927_p),
    .din1(G4_p_spl_00),
    .din2(G18_p_spl_001)
  );


  orX
  g_g1927_n
  (
    .dout(g1927_n),
    .din1(G4_n_spl_0),
    .din2(G18_n_spl_001)
  );


  andX
  g_g1928_p
  (
    .dout(g1928_p),
    .din1(g1926_p_spl_),
    .din2(g1927_p_spl_)
  );


  orX
  g_g1928_n
  (
    .dout(g1928_n),
    .din1(g1926_n_spl_),
    .din2(g1927_n_spl_)
  );


  andX
  g_g1929_p
  (
    .dout(g1929_p),
    .din1(g1926_n_spl_),
    .din2(g1927_n_spl_)
  );


  orX
  g_g1929_n
  (
    .dout(g1929_n),
    .din1(g1926_p_spl_),
    .din2(g1927_p_spl_)
  );


  andX
  g_g1930_p
  (
    .dout(g1930_p),
    .din1(g1928_n_spl_0),
    .din2(g1929_n)
  );


  orX
  g_g1930_n
  (
    .dout(g1930_n),
    .din1(g1928_p_spl_0),
    .din2(g1929_p)
  );


  andX
  g_g1931_p
  (
    .dout(g1931_p),
    .din1(g1582_n_spl_0),
    .din2(g1930_n_spl_)
  );


  orX
  g_g1931_n
  (
    .dout(g1931_n),
    .din1(g1582_p_spl_0),
    .din2(g1930_p_spl_)
  );


  andX
  g_g1932_p
  (
    .dout(g1932_p),
    .din1(G3_p_spl_01),
    .din2(G19_p_spl_001)
  );


  orX
  g_g1932_n
  (
    .dout(g1932_n),
    .din1(G3_n_spl_1),
    .din2(G19_n_spl_001)
  );


  andX
  g_g1933_p
  (
    .dout(g1933_p),
    .din1(g1582_p_spl_),
    .din2(g1930_p_spl_)
  );


  orX
  g_g1933_n
  (
    .dout(g1933_n),
    .din1(g1582_n_spl_),
    .din2(g1930_n_spl_)
  );


  andX
  g_g1934_p
  (
    .dout(g1934_p),
    .din1(g1931_n_spl_),
    .din2(g1933_n)
  );


  orX
  g_g1934_n
  (
    .dout(g1934_n),
    .din1(g1931_p_spl_),
    .din2(g1933_p)
  );


  andX
  g_g1935_p
  (
    .dout(g1935_p),
    .din1(g1932_n_spl_),
    .din2(g1934_p_spl_)
  );


  orX
  g_g1935_n
  (
    .dout(g1935_n),
    .din1(g1932_p_spl_),
    .din2(g1934_n_spl_)
  );


  andX
  g_g1936_p
  (
    .dout(g1936_p),
    .din1(g1931_n_spl_),
    .din2(g1935_n_spl_)
  );


  orX
  g_g1936_n
  (
    .dout(g1936_n),
    .din1(g1931_p_spl_),
    .din2(g1935_p_spl_)
  );


  andX
  g_g1937_p
  (
    .dout(g1937_p),
    .din1(G4_p_spl_01),
    .din2(G19_p_spl_001)
  );


  orX
  g_g1937_n
  (
    .dout(g1937_n),
    .din1(G4_n_spl_1),
    .din2(G19_n_spl_001)
  );


  andX
  g_g1938_p
  (
    .dout(g1938_p),
    .din1(G6_p_spl_00),
    .din2(G17_p_spl_010)
  );


  orX
  g_g1938_n
  (
    .dout(g1938_n),
    .din1(G6_n_spl_0),
    .din2(G17_n_spl_010)
  );


  andX
  g_g1939_p
  (
    .dout(g1939_p),
    .din1(G5_p_spl_00),
    .din2(G18_p_spl_010)
  );


  orX
  g_g1939_n
  (
    .dout(g1939_n),
    .din1(G5_n_spl_0),
    .din2(G18_n_spl_010)
  );


  andX
  g_g1940_p
  (
    .dout(g1940_p),
    .din1(g1938_p_spl_),
    .din2(g1939_p_spl_)
  );


  orX
  g_g1940_n
  (
    .dout(g1940_n),
    .din1(g1938_n_spl_),
    .din2(g1939_n_spl_)
  );


  andX
  g_g1941_p
  (
    .dout(g1941_p),
    .din1(g1938_n_spl_),
    .din2(g1939_n_spl_)
  );


  orX
  g_g1941_n
  (
    .dout(g1941_n),
    .din1(g1938_p_spl_),
    .din2(g1939_p_spl_)
  );


  andX
  g_g1942_p
  (
    .dout(g1942_p),
    .din1(g1940_n_spl_0),
    .din2(g1941_n)
  );


  orX
  g_g1942_n
  (
    .dout(g1942_n),
    .din1(g1940_p_spl_0),
    .din2(g1941_p)
  );


  andX
  g_g1943_p
  (
    .dout(g1943_p),
    .din1(g1928_n_spl_0),
    .din2(g1942_n_spl_)
  );


  orX
  g_g1943_n
  (
    .dout(g1943_n),
    .din1(g1928_p_spl_0),
    .din2(g1942_p_spl_)
  );


  andX
  g_g1944_p
  (
    .dout(g1944_p),
    .din1(g1928_p_spl_),
    .din2(g1942_p_spl_)
  );


  orX
  g_g1944_n
  (
    .dout(g1944_n),
    .din1(g1928_n_spl_),
    .din2(g1942_n_spl_)
  );


  andX
  g_g1945_p
  (
    .dout(g1945_p),
    .din1(g1943_n_spl_),
    .din2(g1944_n)
  );


  orX
  g_g1945_n
  (
    .dout(g1945_n),
    .din1(g1943_p_spl_),
    .din2(g1944_p)
  );


  andX
  g_g1946_p
  (
    .dout(g1946_p),
    .din1(g1937_n_spl_),
    .din2(g1945_p_spl_)
  );


  orX
  g_g1946_n
  (
    .dout(g1946_n),
    .din1(g1937_p_spl_),
    .din2(g1945_n_spl_)
  );


  andX
  g_g1947_p
  (
    .dout(g1947_p),
    .din1(g1937_p_spl_),
    .din2(g1945_n_spl_)
  );


  orX
  g_g1947_n
  (
    .dout(g1947_n),
    .din1(g1937_n_spl_),
    .din2(g1945_p_spl_)
  );


  andX
  g_g1948_p
  (
    .dout(g1948_p),
    .din1(g1946_n_spl_),
    .din2(g1947_n)
  );


  orX
  g_g1948_n
  (
    .dout(g1948_n),
    .din1(g1946_p_spl_),
    .din2(g1947_p)
  );


  andX
  g_g1949_p
  (
    .dout(g1949_p),
    .din1(g1936_n_spl_),
    .din2(g1948_p_spl_)
  );


  orX
  g_g1949_n
  (
    .dout(g1949_n),
    .din1(g1936_p_spl_),
    .din2(g1948_n_spl_)
  );


  andX
  g_g1950_p
  (
    .dout(g1950_p),
    .din1(G3_p_spl_01),
    .din2(G20_p_spl_000)
  );


  orX
  g_g1950_n
  (
    .dout(g1950_n),
    .din1(G3_n_spl_1),
    .din2(G20_n_spl_000)
  );


  andX
  g_g1951_p
  (
    .dout(g1951_p),
    .din1(g1936_p_spl_),
    .din2(g1948_n_spl_)
  );


  orX
  g_g1951_n
  (
    .dout(g1951_n),
    .din1(g1936_n_spl_),
    .din2(g1948_p_spl_)
  );


  andX
  g_g1952_p
  (
    .dout(g1952_p),
    .din1(g1949_n_spl_),
    .din2(g1951_n)
  );


  orX
  g_g1952_n
  (
    .dout(g1952_n),
    .din1(g1949_p_spl_),
    .din2(g1951_p)
  );


  andX
  g_g1953_p
  (
    .dout(g1953_p),
    .din1(g1950_n_spl_),
    .din2(g1952_p_spl_)
  );


  orX
  g_g1953_n
  (
    .dout(g1953_n),
    .din1(g1950_p_spl_),
    .din2(g1952_n_spl_)
  );


  andX
  g_g1954_p
  (
    .dout(g1954_p),
    .din1(g1949_n_spl_),
    .din2(g1953_n_spl_)
  );


  orX
  g_g1954_n
  (
    .dout(g1954_n),
    .din1(g1949_p_spl_),
    .din2(g1953_p_spl_)
  );


  andX
  g_g1955_p
  (
    .dout(g1955_p),
    .din1(G4_p_spl_01),
    .din2(G20_p_spl_000)
  );


  orX
  g_g1955_n
  (
    .dout(g1955_n),
    .din1(G4_n_spl_1),
    .din2(G20_n_spl_001)
  );


  andX
  g_g1956_p
  (
    .dout(g1956_p),
    .din1(g1943_n_spl_),
    .din2(g1946_n_spl_)
  );


  orX
  g_g1956_n
  (
    .dout(g1956_n),
    .din1(g1943_p_spl_),
    .din2(g1946_p_spl_)
  );


  andX
  g_g1957_p
  (
    .dout(g1957_p),
    .din1(G5_p_spl_01),
    .din2(G19_p_spl_010)
  );


  orX
  g_g1957_n
  (
    .dout(g1957_n),
    .din1(G5_n_spl_1),
    .din2(G19_n_spl_010)
  );


  andX
  g_g1958_p
  (
    .dout(g1958_p),
    .din1(G7_p_spl_00),
    .din2(G17_p_spl_010)
  );


  orX
  g_g1958_n
  (
    .dout(g1958_n),
    .din1(G7_n_spl_0),
    .din2(G17_n_spl_010)
  );


  andX
  g_g1959_p
  (
    .dout(g1959_p),
    .din1(G6_p_spl_00),
    .din2(G18_p_spl_010)
  );


  orX
  g_g1959_n
  (
    .dout(g1959_n),
    .din1(G6_n_spl_0),
    .din2(G18_n_spl_010)
  );


  andX
  g_g1960_p
  (
    .dout(g1960_p),
    .din1(g1958_p_spl_),
    .din2(g1959_p_spl_)
  );


  orX
  g_g1960_n
  (
    .dout(g1960_n),
    .din1(g1958_n_spl_),
    .din2(g1959_n_spl_)
  );


  andX
  g_g1961_p
  (
    .dout(g1961_p),
    .din1(g1958_n_spl_),
    .din2(g1959_n_spl_)
  );


  orX
  g_g1961_n
  (
    .dout(g1961_n),
    .din1(g1958_p_spl_),
    .din2(g1959_p_spl_)
  );


  andX
  g_g1962_p
  (
    .dout(g1962_p),
    .din1(g1960_n_spl_0),
    .din2(g1961_n)
  );


  orX
  g_g1962_n
  (
    .dout(g1962_n),
    .din1(g1960_p_spl_0),
    .din2(g1961_p)
  );


  andX
  g_g1963_p
  (
    .dout(g1963_p),
    .din1(g1940_n_spl_0),
    .din2(g1962_n_spl_)
  );


  orX
  g_g1963_n
  (
    .dout(g1963_n),
    .din1(g1940_p_spl_0),
    .din2(g1962_p_spl_)
  );


  andX
  g_g1964_p
  (
    .dout(g1964_p),
    .din1(g1940_p_spl_),
    .din2(g1962_p_spl_)
  );


  orX
  g_g1964_n
  (
    .dout(g1964_n),
    .din1(g1940_n_spl_),
    .din2(g1962_n_spl_)
  );


  andX
  g_g1965_p
  (
    .dout(g1965_p),
    .din1(g1963_n_spl_),
    .din2(g1964_n)
  );


  orX
  g_g1965_n
  (
    .dout(g1965_n),
    .din1(g1963_p_spl_),
    .din2(g1964_p)
  );


  andX
  g_g1966_p
  (
    .dout(g1966_p),
    .din1(g1957_n_spl_),
    .din2(g1965_p_spl_)
  );


  orX
  g_g1966_n
  (
    .dout(g1966_n),
    .din1(g1957_p_spl_),
    .din2(g1965_n_spl_)
  );


  andX
  g_g1967_p
  (
    .dout(g1967_p),
    .din1(g1957_p_spl_),
    .din2(g1965_n_spl_)
  );


  orX
  g_g1967_n
  (
    .dout(g1967_n),
    .din1(g1957_n_spl_),
    .din2(g1965_p_spl_)
  );


  andX
  g_g1968_p
  (
    .dout(g1968_p),
    .din1(g1966_n_spl_),
    .din2(g1967_n)
  );


  orX
  g_g1968_n
  (
    .dout(g1968_n),
    .din1(g1966_p_spl_),
    .din2(g1967_p)
  );


  andX
  g_g1969_p
  (
    .dout(g1969_p),
    .din1(g1956_n_spl_),
    .din2(g1968_p_spl_)
  );


  orX
  g_g1969_n
  (
    .dout(g1969_n),
    .din1(g1956_p_spl_),
    .din2(g1968_n_spl_)
  );


  andX
  g_g1970_p
  (
    .dout(g1970_p),
    .din1(g1956_p_spl_),
    .din2(g1968_n_spl_)
  );


  orX
  g_g1970_n
  (
    .dout(g1970_n),
    .din1(g1956_n_spl_),
    .din2(g1968_p_spl_)
  );


  andX
  g_g1971_p
  (
    .dout(g1971_p),
    .din1(g1969_n_spl_),
    .din2(g1970_n)
  );


  orX
  g_g1971_n
  (
    .dout(g1971_n),
    .din1(g1969_p_spl_),
    .din2(g1970_p)
  );


  andX
  g_g1972_p
  (
    .dout(g1972_p),
    .din1(g1955_n_spl_),
    .din2(g1971_p_spl_)
  );


  orX
  g_g1972_n
  (
    .dout(g1972_n),
    .din1(g1955_p_spl_),
    .din2(g1971_n_spl_)
  );


  andX
  g_g1973_p
  (
    .dout(g1973_p),
    .din1(g1955_p_spl_),
    .din2(g1971_n_spl_)
  );


  orX
  g_g1973_n
  (
    .dout(g1973_n),
    .din1(g1955_n_spl_),
    .din2(g1971_p_spl_)
  );


  andX
  g_g1974_p
  (
    .dout(g1974_p),
    .din1(g1972_n_spl_),
    .din2(g1973_n)
  );


  orX
  g_g1974_n
  (
    .dout(g1974_n),
    .din1(g1972_p_spl_),
    .din2(g1973_p)
  );


  orX
  g_g1975_n
  (
    .dout(g1975_n),
    .din1(g1954_p),
    .din2(g1974_n)
  );


  andX
  g_g1976_p
  (
    .dout(g1976_p),
    .din1(g1969_n_spl_),
    .din2(g1972_n_spl_)
  );


  orX
  g_g1976_n
  (
    .dout(g1976_n),
    .din1(g1969_p_spl_),
    .din2(g1972_p_spl_)
  );


  andX
  g_g1977_p
  (
    .dout(g1977_p),
    .din1(G5_p_spl_01),
    .din2(G20_p_spl_001)
  );


  orX
  g_g1977_n
  (
    .dout(g1977_n),
    .din1(G5_n_spl_1),
    .din2(G20_n_spl_001)
  );


  andX
  g_g1978_p
  (
    .dout(g1978_p),
    .din1(g1963_n_spl_),
    .din2(g1966_n_spl_)
  );


  orX
  g_g1978_n
  (
    .dout(g1978_n),
    .din1(g1963_p_spl_),
    .din2(g1966_p_spl_)
  );


  andX
  g_g1979_p
  (
    .dout(g1979_p),
    .din1(G6_p_spl_01),
    .din2(G19_p_spl_010)
  );


  orX
  g_g1979_n
  (
    .dout(g1979_n),
    .din1(G6_n_spl_1),
    .din2(G19_n_spl_010)
  );


  andX
  g_g1980_p
  (
    .dout(g1980_p),
    .din1(G8_p_spl_00),
    .din2(G17_p_spl_011)
  );


  orX
  g_g1980_n
  (
    .dout(g1980_n),
    .din1(G8_n_spl_0),
    .din2(G17_n_spl_011)
  );


  andX
  g_g1981_p
  (
    .dout(g1981_p),
    .din1(G7_p_spl_00),
    .din2(G18_p_spl_011)
  );


  orX
  g_g1981_n
  (
    .dout(g1981_n),
    .din1(G7_n_spl_0),
    .din2(G18_n_spl_011)
  );


  andX
  g_g1982_p
  (
    .dout(g1982_p),
    .din1(g1980_p_spl_),
    .din2(g1981_p_spl_)
  );


  orX
  g_g1982_n
  (
    .dout(g1982_n),
    .din1(g1980_n_spl_),
    .din2(g1981_n_spl_)
  );


  andX
  g_g1983_p
  (
    .dout(g1983_p),
    .din1(g1980_n_spl_),
    .din2(g1981_n_spl_)
  );


  orX
  g_g1983_n
  (
    .dout(g1983_n),
    .din1(g1980_p_spl_),
    .din2(g1981_p_spl_)
  );


  andX
  g_g1984_p
  (
    .dout(g1984_p),
    .din1(g1982_n_spl_0),
    .din2(g1983_n)
  );


  orX
  g_g1984_n
  (
    .dout(g1984_n),
    .din1(g1982_p_spl_0),
    .din2(g1983_p)
  );


  andX
  g_g1985_p
  (
    .dout(g1985_p),
    .din1(g1960_n_spl_0),
    .din2(g1984_n_spl_)
  );


  orX
  g_g1985_n
  (
    .dout(g1985_n),
    .din1(g1960_p_spl_0),
    .din2(g1984_p_spl_)
  );


  andX
  g_g1986_p
  (
    .dout(g1986_p),
    .din1(g1960_p_spl_),
    .din2(g1984_p_spl_)
  );


  orX
  g_g1986_n
  (
    .dout(g1986_n),
    .din1(g1960_n_spl_),
    .din2(g1984_n_spl_)
  );


  andX
  g_g1987_p
  (
    .dout(g1987_p),
    .din1(g1985_n_spl_),
    .din2(g1986_n)
  );


  orX
  g_g1987_n
  (
    .dout(g1987_n),
    .din1(g1985_p_spl_),
    .din2(g1986_p)
  );


  andX
  g_g1988_p
  (
    .dout(g1988_p),
    .din1(g1979_n_spl_),
    .din2(g1987_p_spl_)
  );


  orX
  g_g1988_n
  (
    .dout(g1988_n),
    .din1(g1979_p_spl_),
    .din2(g1987_n_spl_)
  );


  andX
  g_g1989_p
  (
    .dout(g1989_p),
    .din1(g1979_p_spl_),
    .din2(g1987_n_spl_)
  );


  orX
  g_g1989_n
  (
    .dout(g1989_n),
    .din1(g1979_n_spl_),
    .din2(g1987_p_spl_)
  );


  andX
  g_g1990_p
  (
    .dout(g1990_p),
    .din1(g1988_n_spl_),
    .din2(g1989_n)
  );


  orX
  g_g1990_n
  (
    .dout(g1990_n),
    .din1(g1988_p_spl_),
    .din2(g1989_p)
  );


  andX
  g_g1991_p
  (
    .dout(g1991_p),
    .din1(g1978_n_spl_),
    .din2(g1990_p_spl_)
  );


  orX
  g_g1991_n
  (
    .dout(g1991_n),
    .din1(g1978_p_spl_),
    .din2(g1990_n_spl_)
  );


  andX
  g_g1992_p
  (
    .dout(g1992_p),
    .din1(g1978_p_spl_),
    .din2(g1990_n_spl_)
  );


  orX
  g_g1992_n
  (
    .dout(g1992_n),
    .din1(g1978_n_spl_),
    .din2(g1990_p_spl_)
  );


  andX
  g_g1993_p
  (
    .dout(g1993_p),
    .din1(g1991_n_spl_),
    .din2(g1992_n)
  );


  orX
  g_g1993_n
  (
    .dout(g1993_n),
    .din1(g1991_p_spl_),
    .din2(g1992_p)
  );


  andX
  g_g1994_p
  (
    .dout(g1994_p),
    .din1(g1977_n_spl_),
    .din2(g1993_p_spl_)
  );


  orX
  g_g1994_n
  (
    .dout(g1994_n),
    .din1(g1977_p_spl_),
    .din2(g1993_n_spl_)
  );


  andX
  g_g1995_p
  (
    .dout(g1995_p),
    .din1(g1977_p_spl_),
    .din2(g1993_n_spl_)
  );


  orX
  g_g1995_n
  (
    .dout(g1995_n),
    .din1(g1977_n_spl_),
    .din2(g1993_p_spl_)
  );


  andX
  g_g1996_p
  (
    .dout(g1996_p),
    .din1(g1994_n_spl_),
    .din2(g1995_n)
  );


  orX
  g_g1996_n
  (
    .dout(g1996_n),
    .din1(g1994_p_spl_),
    .din2(g1995_p)
  );


  orX
  g_g1997_n
  (
    .dout(g1997_n),
    .din1(g1976_p),
    .din2(g1996_n)
  );


  andX
  g_g1998_p
  (
    .dout(g1998_p),
    .din1(g1991_n_spl_),
    .din2(g1994_n_spl_)
  );


  orX
  g_g1998_n
  (
    .dout(g1998_n),
    .din1(g1991_p_spl_),
    .din2(g1994_p_spl_)
  );


  andX
  g_g1999_p
  (
    .dout(g1999_p),
    .din1(G6_p_spl_01),
    .din2(G20_p_spl_001)
  );


  orX
  g_g1999_n
  (
    .dout(g1999_n),
    .din1(G6_n_spl_1),
    .din2(G20_n_spl_010)
  );


  andX
  g_g2000_p
  (
    .dout(g2000_p),
    .din1(g1985_n_spl_),
    .din2(g1988_n_spl_)
  );


  orX
  g_g2000_n
  (
    .dout(g2000_n),
    .din1(g1985_p_spl_),
    .din2(g1988_p_spl_)
  );


  andX
  g_g2001_p
  (
    .dout(g2001_p),
    .din1(G7_p_spl_01),
    .din2(G19_p_spl_011)
  );


  orX
  g_g2001_n
  (
    .dout(g2001_n),
    .din1(G7_n_spl_1),
    .din2(G19_n_spl_011)
  );


  andX
  g_g2002_p
  (
    .dout(g2002_p),
    .din1(G9_p_spl_00),
    .din2(G17_p_spl_011)
  );


  orX
  g_g2002_n
  (
    .dout(g2002_n),
    .din1(G9_n_spl_0),
    .din2(G17_n_spl_011)
  );


  andX
  g_g2003_p
  (
    .dout(g2003_p),
    .din1(G8_p_spl_00),
    .din2(G18_p_spl_011)
  );


  orX
  g_g2003_n
  (
    .dout(g2003_n),
    .din1(G8_n_spl_0),
    .din2(G18_n_spl_011)
  );


  andX
  g_g2004_p
  (
    .dout(g2004_p),
    .din1(g2002_p_spl_),
    .din2(g2003_p_spl_)
  );


  orX
  g_g2004_n
  (
    .dout(g2004_n),
    .din1(g2002_n_spl_),
    .din2(g2003_n_spl_)
  );


  andX
  g_g2005_p
  (
    .dout(g2005_p),
    .din1(g2002_n_spl_),
    .din2(g2003_n_spl_)
  );


  orX
  g_g2005_n
  (
    .dout(g2005_n),
    .din1(g2002_p_spl_),
    .din2(g2003_p_spl_)
  );


  andX
  g_g2006_p
  (
    .dout(g2006_p),
    .din1(g2004_n_spl_0),
    .din2(g2005_n)
  );


  orX
  g_g2006_n
  (
    .dout(g2006_n),
    .din1(g2004_p_spl_0),
    .din2(g2005_p)
  );


  andX
  g_g2007_p
  (
    .dout(g2007_p),
    .din1(g1982_n_spl_0),
    .din2(g2006_n_spl_)
  );


  orX
  g_g2007_n
  (
    .dout(g2007_n),
    .din1(g1982_p_spl_0),
    .din2(g2006_p_spl_)
  );


  andX
  g_g2008_p
  (
    .dout(g2008_p),
    .din1(g1982_p_spl_),
    .din2(g2006_p_spl_)
  );


  orX
  g_g2008_n
  (
    .dout(g2008_n),
    .din1(g1982_n_spl_),
    .din2(g2006_n_spl_)
  );


  andX
  g_g2009_p
  (
    .dout(g2009_p),
    .din1(g2007_n_spl_),
    .din2(g2008_n)
  );


  orX
  g_g2009_n
  (
    .dout(g2009_n),
    .din1(g2007_p_spl_),
    .din2(g2008_p)
  );


  andX
  g_g2010_p
  (
    .dout(g2010_p),
    .din1(g2001_n_spl_),
    .din2(g2009_p_spl_)
  );


  orX
  g_g2010_n
  (
    .dout(g2010_n),
    .din1(g2001_p_spl_),
    .din2(g2009_n_spl_)
  );


  andX
  g_g2011_p
  (
    .dout(g2011_p),
    .din1(g2001_p_spl_),
    .din2(g2009_n_spl_)
  );


  orX
  g_g2011_n
  (
    .dout(g2011_n),
    .din1(g2001_n_spl_),
    .din2(g2009_p_spl_)
  );


  andX
  g_g2012_p
  (
    .dout(g2012_p),
    .din1(g2010_n_spl_),
    .din2(g2011_n)
  );


  orX
  g_g2012_n
  (
    .dout(g2012_n),
    .din1(g2010_p_spl_),
    .din2(g2011_p)
  );


  andX
  g_g2013_p
  (
    .dout(g2013_p),
    .din1(g2000_n_spl_),
    .din2(g2012_p_spl_)
  );


  orX
  g_g2013_n
  (
    .dout(g2013_n),
    .din1(g2000_p_spl_),
    .din2(g2012_n_spl_)
  );


  andX
  g_g2014_p
  (
    .dout(g2014_p),
    .din1(g2000_p_spl_),
    .din2(g2012_n_spl_)
  );


  orX
  g_g2014_n
  (
    .dout(g2014_n),
    .din1(g2000_n_spl_),
    .din2(g2012_p_spl_)
  );


  andX
  g_g2015_p
  (
    .dout(g2015_p),
    .din1(g2013_n_spl_),
    .din2(g2014_n)
  );


  orX
  g_g2015_n
  (
    .dout(g2015_n),
    .din1(g2013_p_spl_),
    .din2(g2014_p)
  );


  andX
  g_g2016_p
  (
    .dout(g2016_p),
    .din1(g1999_n_spl_),
    .din2(g2015_p_spl_)
  );


  orX
  g_g2016_n
  (
    .dout(g2016_n),
    .din1(g1999_p_spl_),
    .din2(g2015_n_spl_)
  );


  andX
  g_g2017_p
  (
    .dout(g2017_p),
    .din1(g1999_p_spl_),
    .din2(g2015_n_spl_)
  );


  orX
  g_g2017_n
  (
    .dout(g2017_n),
    .din1(g1999_n_spl_),
    .din2(g2015_p_spl_)
  );


  andX
  g_g2018_p
  (
    .dout(g2018_p),
    .din1(g2016_n_spl_),
    .din2(g2017_n)
  );


  orX
  g_g2018_n
  (
    .dout(g2018_n),
    .din1(g2016_p_spl_),
    .din2(g2017_p)
  );


  orX
  g_g2019_n
  (
    .dout(g2019_n),
    .din1(g1998_p),
    .din2(g2018_n)
  );


  andX
  g_g2020_p
  (
    .dout(g2020_p),
    .din1(g2013_n_spl_),
    .din2(g2016_n_spl_)
  );


  orX
  g_g2020_n
  (
    .dout(g2020_n),
    .din1(g2013_p_spl_),
    .din2(g2016_p_spl_)
  );


  andX
  g_g2021_p
  (
    .dout(g2021_p),
    .din1(G7_p_spl_01),
    .din2(G20_p_spl_010)
  );


  orX
  g_g2021_n
  (
    .dout(g2021_n),
    .din1(G7_n_spl_1),
    .din2(G20_n_spl_010)
  );


  andX
  g_g2022_p
  (
    .dout(g2022_p),
    .din1(g2007_n_spl_),
    .din2(g2010_n_spl_)
  );


  orX
  g_g2022_n
  (
    .dout(g2022_n),
    .din1(g2007_p_spl_),
    .din2(g2010_p_spl_)
  );


  andX
  g_g2023_p
  (
    .dout(g2023_p),
    .din1(G8_p_spl_01),
    .din2(G19_p_spl_011)
  );


  orX
  g_g2023_n
  (
    .dout(g2023_n),
    .din1(G8_n_spl_1),
    .din2(G19_n_spl_011)
  );


  andX
  g_g2024_p
  (
    .dout(g2024_p),
    .din1(G10_p_spl_00),
    .din2(G17_p_spl_100)
  );


  orX
  g_g2024_n
  (
    .dout(g2024_n),
    .din1(G10_n_spl_0),
    .din2(G17_n_spl_100)
  );


  andX
  g_g2025_p
  (
    .dout(g2025_p),
    .din1(G9_p_spl_00),
    .din2(G18_p_spl_100)
  );


  orX
  g_g2025_n
  (
    .dout(g2025_n),
    .din1(G9_n_spl_0),
    .din2(G18_n_spl_100)
  );


  andX
  g_g2026_p
  (
    .dout(g2026_p),
    .din1(g2024_p_spl_),
    .din2(g2025_p_spl_)
  );


  orX
  g_g2026_n
  (
    .dout(g2026_n),
    .din1(g2024_n_spl_),
    .din2(g2025_n_spl_)
  );


  andX
  g_g2027_p
  (
    .dout(g2027_p),
    .din1(g2024_n_spl_),
    .din2(g2025_n_spl_)
  );


  orX
  g_g2027_n
  (
    .dout(g2027_n),
    .din1(g2024_p_spl_),
    .din2(g2025_p_spl_)
  );


  andX
  g_g2028_p
  (
    .dout(g2028_p),
    .din1(g2026_n_spl_0),
    .din2(g2027_n)
  );


  orX
  g_g2028_n
  (
    .dout(g2028_n),
    .din1(g2026_p_spl_0),
    .din2(g2027_p)
  );


  andX
  g_g2029_p
  (
    .dout(g2029_p),
    .din1(g2004_n_spl_0),
    .din2(g2028_n_spl_)
  );


  orX
  g_g2029_n
  (
    .dout(g2029_n),
    .din1(g2004_p_spl_0),
    .din2(g2028_p_spl_)
  );


  andX
  g_g2030_p
  (
    .dout(g2030_p),
    .din1(g2004_p_spl_),
    .din2(g2028_p_spl_)
  );


  orX
  g_g2030_n
  (
    .dout(g2030_n),
    .din1(g2004_n_spl_),
    .din2(g2028_n_spl_)
  );


  andX
  g_g2031_p
  (
    .dout(g2031_p),
    .din1(g2029_n_spl_),
    .din2(g2030_n)
  );


  orX
  g_g2031_n
  (
    .dout(g2031_n),
    .din1(g2029_p_spl_),
    .din2(g2030_p)
  );


  andX
  g_g2032_p
  (
    .dout(g2032_p),
    .din1(g2023_n_spl_),
    .din2(g2031_p_spl_)
  );


  orX
  g_g2032_n
  (
    .dout(g2032_n),
    .din1(g2023_p_spl_),
    .din2(g2031_n_spl_)
  );


  andX
  g_g2033_p
  (
    .dout(g2033_p),
    .din1(g2023_p_spl_),
    .din2(g2031_n_spl_)
  );


  orX
  g_g2033_n
  (
    .dout(g2033_n),
    .din1(g2023_n_spl_),
    .din2(g2031_p_spl_)
  );


  andX
  g_g2034_p
  (
    .dout(g2034_p),
    .din1(g2032_n_spl_),
    .din2(g2033_n)
  );


  orX
  g_g2034_n
  (
    .dout(g2034_n),
    .din1(g2032_p_spl_),
    .din2(g2033_p)
  );


  andX
  g_g2035_p
  (
    .dout(g2035_p),
    .din1(g2022_n_spl_),
    .din2(g2034_p_spl_)
  );


  orX
  g_g2035_n
  (
    .dout(g2035_n),
    .din1(g2022_p_spl_),
    .din2(g2034_n_spl_)
  );


  andX
  g_g2036_p
  (
    .dout(g2036_p),
    .din1(g2022_p_spl_),
    .din2(g2034_n_spl_)
  );


  orX
  g_g2036_n
  (
    .dout(g2036_n),
    .din1(g2022_n_spl_),
    .din2(g2034_p_spl_)
  );


  andX
  g_g2037_p
  (
    .dout(g2037_p),
    .din1(g2035_n_spl_),
    .din2(g2036_n)
  );


  orX
  g_g2037_n
  (
    .dout(g2037_n),
    .din1(g2035_p_spl_),
    .din2(g2036_p)
  );


  andX
  g_g2038_p
  (
    .dout(g2038_p),
    .din1(g2021_n_spl_),
    .din2(g2037_p_spl_)
  );


  orX
  g_g2038_n
  (
    .dout(g2038_n),
    .din1(g2021_p_spl_),
    .din2(g2037_n_spl_)
  );


  andX
  g_g2039_p
  (
    .dout(g2039_p),
    .din1(g2021_p_spl_),
    .din2(g2037_n_spl_)
  );


  orX
  g_g2039_n
  (
    .dout(g2039_n),
    .din1(g2021_n_spl_),
    .din2(g2037_p_spl_)
  );


  andX
  g_g2040_p
  (
    .dout(g2040_p),
    .din1(g2038_n_spl_),
    .din2(g2039_n)
  );


  orX
  g_g2040_n
  (
    .dout(g2040_n),
    .din1(g2038_p_spl_),
    .din2(g2039_p)
  );


  orX
  g_g2041_n
  (
    .dout(g2041_n),
    .din1(g2020_p),
    .din2(g2040_n)
  );


  andX
  g_g2042_p
  (
    .dout(g2042_p),
    .din1(g2035_n_spl_),
    .din2(g2038_n_spl_)
  );


  orX
  g_g2042_n
  (
    .dout(g2042_n),
    .din1(g2035_p_spl_),
    .din2(g2038_p_spl_)
  );


  andX
  g_g2043_p
  (
    .dout(g2043_p),
    .din1(G8_p_spl_01),
    .din2(G20_p_spl_010)
  );


  orX
  g_g2043_n
  (
    .dout(g2043_n),
    .din1(G8_n_spl_1),
    .din2(G20_n_spl_011)
  );


  andX
  g_g2044_p
  (
    .dout(g2044_p),
    .din1(g2029_n_spl_),
    .din2(g2032_n_spl_)
  );


  orX
  g_g2044_n
  (
    .dout(g2044_n),
    .din1(g2029_p_spl_),
    .din2(g2032_p_spl_)
  );


  andX
  g_g2045_p
  (
    .dout(g2045_p),
    .din1(G9_p_spl_01),
    .din2(G19_p_spl_100)
  );


  orX
  g_g2045_n
  (
    .dout(g2045_n),
    .din1(G9_n_spl_1),
    .din2(G19_n_spl_100)
  );


  andX
  g_g2046_p
  (
    .dout(g2046_p),
    .din1(G11_p_spl_00),
    .din2(G17_p_spl_100)
  );


  orX
  g_g2046_n
  (
    .dout(g2046_n),
    .din1(G11_n_spl_0),
    .din2(G17_n_spl_100)
  );


  andX
  g_g2047_p
  (
    .dout(g2047_p),
    .din1(G10_p_spl_00),
    .din2(G18_p_spl_100)
  );


  orX
  g_g2047_n
  (
    .dout(g2047_n),
    .din1(G10_n_spl_0),
    .din2(G18_n_spl_100)
  );


  andX
  g_g2048_p
  (
    .dout(g2048_p),
    .din1(g2046_p_spl_),
    .din2(g2047_p_spl_)
  );


  orX
  g_g2048_n
  (
    .dout(g2048_n),
    .din1(g2046_n_spl_),
    .din2(g2047_n_spl_)
  );


  andX
  g_g2049_p
  (
    .dout(g2049_p),
    .din1(g2046_n_spl_),
    .din2(g2047_n_spl_)
  );


  orX
  g_g2049_n
  (
    .dout(g2049_n),
    .din1(g2046_p_spl_),
    .din2(g2047_p_spl_)
  );


  andX
  g_g2050_p
  (
    .dout(g2050_p),
    .din1(g2048_n_spl_0),
    .din2(g2049_n)
  );


  orX
  g_g2050_n
  (
    .dout(g2050_n),
    .din1(g2048_p_spl_0),
    .din2(g2049_p)
  );


  andX
  g_g2051_p
  (
    .dout(g2051_p),
    .din1(g2026_n_spl_0),
    .din2(g2050_n_spl_)
  );


  orX
  g_g2051_n
  (
    .dout(g2051_n),
    .din1(g2026_p_spl_0),
    .din2(g2050_p_spl_)
  );


  andX
  g_g2052_p
  (
    .dout(g2052_p),
    .din1(g2026_p_spl_),
    .din2(g2050_p_spl_)
  );


  orX
  g_g2052_n
  (
    .dout(g2052_n),
    .din1(g2026_n_spl_),
    .din2(g2050_n_spl_)
  );


  andX
  g_g2053_p
  (
    .dout(g2053_p),
    .din1(g2051_n_spl_),
    .din2(g2052_n)
  );


  orX
  g_g2053_n
  (
    .dout(g2053_n),
    .din1(g2051_p_spl_),
    .din2(g2052_p)
  );


  andX
  g_g2054_p
  (
    .dout(g2054_p),
    .din1(g2045_n_spl_),
    .din2(g2053_p_spl_)
  );


  orX
  g_g2054_n
  (
    .dout(g2054_n),
    .din1(g2045_p_spl_),
    .din2(g2053_n_spl_)
  );


  andX
  g_g2055_p
  (
    .dout(g2055_p),
    .din1(g2045_p_spl_),
    .din2(g2053_n_spl_)
  );


  orX
  g_g2055_n
  (
    .dout(g2055_n),
    .din1(g2045_n_spl_),
    .din2(g2053_p_spl_)
  );


  andX
  g_g2056_p
  (
    .dout(g2056_p),
    .din1(g2054_n_spl_),
    .din2(g2055_n)
  );


  orX
  g_g2056_n
  (
    .dout(g2056_n),
    .din1(g2054_p_spl_),
    .din2(g2055_p)
  );


  andX
  g_g2057_p
  (
    .dout(g2057_p),
    .din1(g2044_n_spl_),
    .din2(g2056_p_spl_)
  );


  orX
  g_g2057_n
  (
    .dout(g2057_n),
    .din1(g2044_p_spl_),
    .din2(g2056_n_spl_)
  );


  andX
  g_g2058_p
  (
    .dout(g2058_p),
    .din1(g2044_p_spl_),
    .din2(g2056_n_spl_)
  );


  orX
  g_g2058_n
  (
    .dout(g2058_n),
    .din1(g2044_n_spl_),
    .din2(g2056_p_spl_)
  );


  andX
  g_g2059_p
  (
    .dout(g2059_p),
    .din1(g2057_n_spl_),
    .din2(g2058_n)
  );


  orX
  g_g2059_n
  (
    .dout(g2059_n),
    .din1(g2057_p_spl_),
    .din2(g2058_p)
  );


  andX
  g_g2060_p
  (
    .dout(g2060_p),
    .din1(g2043_n_spl_),
    .din2(g2059_p_spl_)
  );


  orX
  g_g2060_n
  (
    .dout(g2060_n),
    .din1(g2043_p_spl_),
    .din2(g2059_n_spl_)
  );


  andX
  g_g2061_p
  (
    .dout(g2061_p),
    .din1(g2043_p_spl_),
    .din2(g2059_n_spl_)
  );


  orX
  g_g2061_n
  (
    .dout(g2061_n),
    .din1(g2043_n_spl_),
    .din2(g2059_p_spl_)
  );


  andX
  g_g2062_p
  (
    .dout(g2062_p),
    .din1(g2060_n_spl_),
    .din2(g2061_n)
  );


  orX
  g_g2062_n
  (
    .dout(g2062_n),
    .din1(g2060_p_spl_),
    .din2(g2061_p)
  );


  orX
  g_g2063_n
  (
    .dout(g2063_n),
    .din1(g2042_p),
    .din2(g2062_n)
  );


  andX
  g_g2064_p
  (
    .dout(g2064_p),
    .din1(g2057_n_spl_),
    .din2(g2060_n_spl_)
  );


  orX
  g_g2064_n
  (
    .dout(g2064_n),
    .din1(g2057_p_spl_),
    .din2(g2060_p_spl_)
  );


  andX
  g_g2065_p
  (
    .dout(g2065_p),
    .din1(G9_p_spl_01),
    .din2(G20_p_spl_011)
  );


  orX
  g_g2065_n
  (
    .dout(g2065_n),
    .din1(G9_n_spl_1),
    .din2(G20_n_spl_011)
  );


  andX
  g_g2066_p
  (
    .dout(g2066_p),
    .din1(g2051_n_spl_),
    .din2(g2054_n_spl_)
  );


  orX
  g_g2066_n
  (
    .dout(g2066_n),
    .din1(g2051_p_spl_),
    .din2(g2054_p_spl_)
  );


  andX
  g_g2067_p
  (
    .dout(g2067_p),
    .din1(G10_p_spl_01),
    .din2(G19_p_spl_100)
  );


  orX
  g_g2067_n
  (
    .dout(g2067_n),
    .din1(G10_n_spl_1),
    .din2(G19_n_spl_100)
  );


  andX
  g_g2068_p
  (
    .dout(g2068_p),
    .din1(G12_p_spl_00),
    .din2(G17_p_spl_101)
  );


  orX
  g_g2068_n
  (
    .dout(g2068_n),
    .din1(G12_n_spl_0),
    .din2(G17_n_spl_101)
  );


  andX
  g_g2069_p
  (
    .dout(g2069_p),
    .din1(G11_p_spl_00),
    .din2(G18_p_spl_101)
  );


  orX
  g_g2069_n
  (
    .dout(g2069_n),
    .din1(G11_n_spl_0),
    .din2(G18_n_spl_101)
  );


  andX
  g_g2070_p
  (
    .dout(g2070_p),
    .din1(g2068_p_spl_),
    .din2(g2069_p_spl_)
  );


  orX
  g_g2070_n
  (
    .dout(g2070_n),
    .din1(g2068_n_spl_),
    .din2(g2069_n_spl_)
  );


  andX
  g_g2071_p
  (
    .dout(g2071_p),
    .din1(g2068_n_spl_),
    .din2(g2069_n_spl_)
  );


  orX
  g_g2071_n
  (
    .dout(g2071_n),
    .din1(g2068_p_spl_),
    .din2(g2069_p_spl_)
  );


  andX
  g_g2072_p
  (
    .dout(g2072_p),
    .din1(g2070_n_spl_0),
    .din2(g2071_n)
  );


  orX
  g_g2072_n
  (
    .dout(g2072_n),
    .din1(g2070_p_spl_0),
    .din2(g2071_p)
  );


  andX
  g_g2073_p
  (
    .dout(g2073_p),
    .din1(g2048_n_spl_0),
    .din2(g2072_n_spl_)
  );


  orX
  g_g2073_n
  (
    .dout(g2073_n),
    .din1(g2048_p_spl_0),
    .din2(g2072_p_spl_)
  );


  andX
  g_g2074_p
  (
    .dout(g2074_p),
    .din1(g2048_p_spl_),
    .din2(g2072_p_spl_)
  );


  orX
  g_g2074_n
  (
    .dout(g2074_n),
    .din1(g2048_n_spl_),
    .din2(g2072_n_spl_)
  );


  andX
  g_g2075_p
  (
    .dout(g2075_p),
    .din1(g2073_n_spl_),
    .din2(g2074_n)
  );


  orX
  g_g2075_n
  (
    .dout(g2075_n),
    .din1(g2073_p_spl_),
    .din2(g2074_p)
  );


  andX
  g_g2076_p
  (
    .dout(g2076_p),
    .din1(g2067_n_spl_),
    .din2(g2075_p_spl_)
  );


  orX
  g_g2076_n
  (
    .dout(g2076_n),
    .din1(g2067_p_spl_),
    .din2(g2075_n_spl_)
  );


  andX
  g_g2077_p
  (
    .dout(g2077_p),
    .din1(g2067_p_spl_),
    .din2(g2075_n_spl_)
  );


  orX
  g_g2077_n
  (
    .dout(g2077_n),
    .din1(g2067_n_spl_),
    .din2(g2075_p_spl_)
  );


  andX
  g_g2078_p
  (
    .dout(g2078_p),
    .din1(g2076_n_spl_),
    .din2(g2077_n)
  );


  orX
  g_g2078_n
  (
    .dout(g2078_n),
    .din1(g2076_p_spl_),
    .din2(g2077_p)
  );


  andX
  g_g2079_p
  (
    .dout(g2079_p),
    .din1(g2066_n_spl_),
    .din2(g2078_p_spl_)
  );


  orX
  g_g2079_n
  (
    .dout(g2079_n),
    .din1(g2066_p_spl_),
    .din2(g2078_n_spl_)
  );


  andX
  g_g2080_p
  (
    .dout(g2080_p),
    .din1(g2066_p_spl_),
    .din2(g2078_n_spl_)
  );


  orX
  g_g2080_n
  (
    .dout(g2080_n),
    .din1(g2066_n_spl_),
    .din2(g2078_p_spl_)
  );


  andX
  g_g2081_p
  (
    .dout(g2081_p),
    .din1(g2079_n_spl_),
    .din2(g2080_n)
  );


  orX
  g_g2081_n
  (
    .dout(g2081_n),
    .din1(g2079_p_spl_),
    .din2(g2080_p)
  );


  andX
  g_g2082_p
  (
    .dout(g2082_p),
    .din1(g2065_n_spl_),
    .din2(g2081_p_spl_)
  );


  orX
  g_g2082_n
  (
    .dout(g2082_n),
    .din1(g2065_p_spl_),
    .din2(g2081_n_spl_)
  );


  andX
  g_g2083_p
  (
    .dout(g2083_p),
    .din1(g2065_p_spl_),
    .din2(g2081_n_spl_)
  );


  orX
  g_g2083_n
  (
    .dout(g2083_n),
    .din1(g2065_n_spl_),
    .din2(g2081_p_spl_)
  );


  andX
  g_g2084_p
  (
    .dout(g2084_p),
    .din1(g2082_n_spl_),
    .din2(g2083_n)
  );


  orX
  g_g2084_n
  (
    .dout(g2084_n),
    .din1(g2082_p_spl_),
    .din2(g2083_p)
  );


  orX
  g_g2085_n
  (
    .dout(g2085_n),
    .din1(g2064_p),
    .din2(g2084_n)
  );


  andX
  g_g2086_p
  (
    .dout(g2086_p),
    .din1(g2079_n_spl_),
    .din2(g2082_n_spl_)
  );


  orX
  g_g2086_n
  (
    .dout(g2086_n),
    .din1(g2079_p_spl_),
    .din2(g2082_p_spl_)
  );


  andX
  g_g2087_p
  (
    .dout(g2087_p),
    .din1(G10_p_spl_01),
    .din2(G20_p_spl_011)
  );


  orX
  g_g2087_n
  (
    .dout(g2087_n),
    .din1(G10_n_spl_1),
    .din2(G20_n_spl_100)
  );


  andX
  g_g2088_p
  (
    .dout(g2088_p),
    .din1(g2073_n_spl_),
    .din2(g2076_n_spl_)
  );


  orX
  g_g2088_n
  (
    .dout(g2088_n),
    .din1(g2073_p_spl_),
    .din2(g2076_p_spl_)
  );


  andX
  g_g2089_p
  (
    .dout(g2089_p),
    .din1(G11_p_spl_01),
    .din2(G19_p_spl_101)
  );


  orX
  g_g2089_n
  (
    .dout(g2089_n),
    .din1(G11_n_spl_1),
    .din2(G19_n_spl_101)
  );


  andX
  g_g2090_p
  (
    .dout(g2090_p),
    .din1(G13_p_spl_00),
    .din2(G17_p_spl_101)
  );


  orX
  g_g2090_n
  (
    .dout(g2090_n),
    .din1(G13_n_spl_0),
    .din2(G17_n_spl_101)
  );


  andX
  g_g2091_p
  (
    .dout(g2091_p),
    .din1(G12_p_spl_00),
    .din2(G18_p_spl_101)
  );


  orX
  g_g2091_n
  (
    .dout(g2091_n),
    .din1(G12_n_spl_0),
    .din2(G18_n_spl_101)
  );


  andX
  g_g2092_p
  (
    .dout(g2092_p),
    .din1(g2090_p_spl_),
    .din2(g2091_p_spl_)
  );


  orX
  g_g2092_n
  (
    .dout(g2092_n),
    .din1(g2090_n_spl_),
    .din2(g2091_n_spl_)
  );


  andX
  g_g2093_p
  (
    .dout(g2093_p),
    .din1(g2090_n_spl_),
    .din2(g2091_n_spl_)
  );


  orX
  g_g2093_n
  (
    .dout(g2093_n),
    .din1(g2090_p_spl_),
    .din2(g2091_p_spl_)
  );


  andX
  g_g2094_p
  (
    .dout(g2094_p),
    .din1(g2092_n_spl_0),
    .din2(g2093_n)
  );


  orX
  g_g2094_n
  (
    .dout(g2094_n),
    .din1(g2092_p_spl_0),
    .din2(g2093_p)
  );


  andX
  g_g2095_p
  (
    .dout(g2095_p),
    .din1(g2070_n_spl_0),
    .din2(g2094_n_spl_)
  );


  orX
  g_g2095_n
  (
    .dout(g2095_n),
    .din1(g2070_p_spl_0),
    .din2(g2094_p_spl_)
  );


  andX
  g_g2096_p
  (
    .dout(g2096_p),
    .din1(g2070_p_spl_),
    .din2(g2094_p_spl_)
  );


  orX
  g_g2096_n
  (
    .dout(g2096_n),
    .din1(g2070_n_spl_),
    .din2(g2094_n_spl_)
  );


  andX
  g_g2097_p
  (
    .dout(g2097_p),
    .din1(g2095_n_spl_),
    .din2(g2096_n)
  );


  orX
  g_g2097_n
  (
    .dout(g2097_n),
    .din1(g2095_p_spl_),
    .din2(g2096_p)
  );


  andX
  g_g2098_p
  (
    .dout(g2098_p),
    .din1(g2089_n_spl_),
    .din2(g2097_p_spl_)
  );


  orX
  g_g2098_n
  (
    .dout(g2098_n),
    .din1(g2089_p_spl_),
    .din2(g2097_n_spl_)
  );


  andX
  g_g2099_p
  (
    .dout(g2099_p),
    .din1(g2089_p_spl_),
    .din2(g2097_n_spl_)
  );


  orX
  g_g2099_n
  (
    .dout(g2099_n),
    .din1(g2089_n_spl_),
    .din2(g2097_p_spl_)
  );


  andX
  g_g2100_p
  (
    .dout(g2100_p),
    .din1(g2098_n_spl_),
    .din2(g2099_n)
  );


  orX
  g_g2100_n
  (
    .dout(g2100_n),
    .din1(g2098_p_spl_),
    .din2(g2099_p)
  );


  andX
  g_g2101_p
  (
    .dout(g2101_p),
    .din1(g2088_n_spl_),
    .din2(g2100_p_spl_)
  );


  orX
  g_g2101_n
  (
    .dout(g2101_n),
    .din1(g2088_p_spl_),
    .din2(g2100_n_spl_)
  );


  andX
  g_g2102_p
  (
    .dout(g2102_p),
    .din1(g2088_p_spl_),
    .din2(g2100_n_spl_)
  );


  orX
  g_g2102_n
  (
    .dout(g2102_n),
    .din1(g2088_n_spl_),
    .din2(g2100_p_spl_)
  );


  andX
  g_g2103_p
  (
    .dout(g2103_p),
    .din1(g2101_n_spl_),
    .din2(g2102_n)
  );


  orX
  g_g2103_n
  (
    .dout(g2103_n),
    .din1(g2101_p_spl_),
    .din2(g2102_p)
  );


  andX
  g_g2104_p
  (
    .dout(g2104_p),
    .din1(g2087_n_spl_),
    .din2(g2103_p_spl_)
  );


  orX
  g_g2104_n
  (
    .dout(g2104_n),
    .din1(g2087_p_spl_),
    .din2(g2103_n_spl_)
  );


  andX
  g_g2105_p
  (
    .dout(g2105_p),
    .din1(g2087_p_spl_),
    .din2(g2103_n_spl_)
  );


  orX
  g_g2105_n
  (
    .dout(g2105_n),
    .din1(g2087_n_spl_),
    .din2(g2103_p_spl_)
  );


  andX
  g_g2106_p
  (
    .dout(g2106_p),
    .din1(g2104_n_spl_),
    .din2(g2105_n)
  );


  orX
  g_g2106_n
  (
    .dout(g2106_n),
    .din1(g2104_p_spl_),
    .din2(g2105_p)
  );


  orX
  g_g2107_n
  (
    .dout(g2107_n),
    .din1(g2086_p),
    .din2(g2106_n)
  );


  andX
  g_g2108_p
  (
    .dout(g2108_p),
    .din1(g2101_n_spl_),
    .din2(g2104_n_spl_)
  );


  orX
  g_g2108_n
  (
    .dout(g2108_n),
    .din1(g2101_p_spl_),
    .din2(g2104_p_spl_)
  );


  andX
  g_g2109_p
  (
    .dout(g2109_p),
    .din1(G11_p_spl_01),
    .din2(G20_p_spl_100)
  );


  orX
  g_g2109_n
  (
    .dout(g2109_n),
    .din1(G11_n_spl_1),
    .din2(G20_n_spl_100)
  );


  andX
  g_g2110_p
  (
    .dout(g2110_p),
    .din1(g2095_n_spl_),
    .din2(g2098_n_spl_)
  );


  orX
  g_g2110_n
  (
    .dout(g2110_n),
    .din1(g2095_p_spl_),
    .din2(g2098_p_spl_)
  );


  andX
  g_g2111_p
  (
    .dout(g2111_p),
    .din1(G12_p_spl_01),
    .din2(G19_p_spl_101)
  );


  orX
  g_g2111_n
  (
    .dout(g2111_n),
    .din1(G12_n_spl_1),
    .din2(G19_n_spl_101)
  );


  andX
  g_g2112_p
  (
    .dout(g2112_p),
    .din1(G14_p_spl_00),
    .din2(G17_p_spl_110)
  );


  orX
  g_g2112_n
  (
    .dout(g2112_n),
    .din1(G14_n_spl_0),
    .din2(G17_n_spl_110)
  );


  andX
  g_g2113_p
  (
    .dout(g2113_p),
    .din1(G13_p_spl_00),
    .din2(G18_p_spl_110)
  );


  orX
  g_g2113_n
  (
    .dout(g2113_n),
    .din1(G13_n_spl_0),
    .din2(G18_n_spl_110)
  );


  andX
  g_g2114_p
  (
    .dout(g2114_p),
    .din1(g2112_p_spl_),
    .din2(g2113_p_spl_)
  );


  orX
  g_g2114_n
  (
    .dout(g2114_n),
    .din1(g2112_n_spl_),
    .din2(g2113_n_spl_)
  );


  andX
  g_g2115_p
  (
    .dout(g2115_p),
    .din1(g2112_n_spl_),
    .din2(g2113_n_spl_)
  );


  orX
  g_g2115_n
  (
    .dout(g2115_n),
    .din1(g2112_p_spl_),
    .din2(g2113_p_spl_)
  );


  andX
  g_g2116_p
  (
    .dout(g2116_p),
    .din1(g2114_n_spl_0),
    .din2(g2115_n)
  );


  orX
  g_g2116_n
  (
    .dout(g2116_n),
    .din1(g2114_p_spl_0),
    .din2(g2115_p)
  );


  andX
  g_g2117_p
  (
    .dout(g2117_p),
    .din1(g2092_n_spl_0),
    .din2(g2116_n_spl_)
  );


  orX
  g_g2117_n
  (
    .dout(g2117_n),
    .din1(g2092_p_spl_0),
    .din2(g2116_p_spl_)
  );


  andX
  g_g2118_p
  (
    .dout(g2118_p),
    .din1(g2092_p_spl_),
    .din2(g2116_p_spl_)
  );


  orX
  g_g2118_n
  (
    .dout(g2118_n),
    .din1(g2092_n_spl_),
    .din2(g2116_n_spl_)
  );


  andX
  g_g2119_p
  (
    .dout(g2119_p),
    .din1(g2117_n_spl_),
    .din2(g2118_n)
  );


  orX
  g_g2119_n
  (
    .dout(g2119_n),
    .din1(g2117_p_spl_),
    .din2(g2118_p)
  );


  andX
  g_g2120_p
  (
    .dout(g2120_p),
    .din1(g2111_n_spl_),
    .din2(g2119_p_spl_)
  );


  orX
  g_g2120_n
  (
    .dout(g2120_n),
    .din1(g2111_p_spl_),
    .din2(g2119_n_spl_)
  );


  andX
  g_g2121_p
  (
    .dout(g2121_p),
    .din1(g2111_p_spl_),
    .din2(g2119_n_spl_)
  );


  orX
  g_g2121_n
  (
    .dout(g2121_n),
    .din1(g2111_n_spl_),
    .din2(g2119_p_spl_)
  );


  andX
  g_g2122_p
  (
    .dout(g2122_p),
    .din1(g2120_n_spl_),
    .din2(g2121_n)
  );


  orX
  g_g2122_n
  (
    .dout(g2122_n),
    .din1(g2120_p_spl_),
    .din2(g2121_p)
  );


  andX
  g_g2123_p
  (
    .dout(g2123_p),
    .din1(g2110_n_spl_),
    .din2(g2122_p_spl_)
  );


  orX
  g_g2123_n
  (
    .dout(g2123_n),
    .din1(g2110_p_spl_),
    .din2(g2122_n_spl_)
  );


  andX
  g_g2124_p
  (
    .dout(g2124_p),
    .din1(g2110_p_spl_),
    .din2(g2122_n_spl_)
  );


  orX
  g_g2124_n
  (
    .dout(g2124_n),
    .din1(g2110_n_spl_),
    .din2(g2122_p_spl_)
  );


  andX
  g_g2125_p
  (
    .dout(g2125_p),
    .din1(g2123_n_spl_),
    .din2(g2124_n)
  );


  orX
  g_g2125_n
  (
    .dout(g2125_n),
    .din1(g2123_p_spl_),
    .din2(g2124_p)
  );


  andX
  g_g2126_p
  (
    .dout(g2126_p),
    .din1(g2109_n_spl_),
    .din2(g2125_p_spl_)
  );


  orX
  g_g2126_n
  (
    .dout(g2126_n),
    .din1(g2109_p_spl_),
    .din2(g2125_n_spl_)
  );


  andX
  g_g2127_p
  (
    .dout(g2127_p),
    .din1(g2109_p_spl_),
    .din2(g2125_n_spl_)
  );


  orX
  g_g2127_n
  (
    .dout(g2127_n),
    .din1(g2109_n_spl_),
    .din2(g2125_p_spl_)
  );


  andX
  g_g2128_p
  (
    .dout(g2128_p),
    .din1(g2126_n_spl_),
    .din2(g2127_n)
  );


  orX
  g_g2128_n
  (
    .dout(g2128_n),
    .din1(g2126_p_spl_),
    .din2(g2127_p)
  );


  orX
  g_g2129_n
  (
    .dout(g2129_n),
    .din1(g2108_p),
    .din2(g2128_n)
  );


  andX
  g_g2130_p
  (
    .dout(g2130_p),
    .din1(g2123_n_spl_),
    .din2(g2126_n_spl_)
  );


  orX
  g_g2130_n
  (
    .dout(g2130_n),
    .din1(g2123_p_spl_),
    .din2(g2126_p_spl_)
  );


  andX
  g_g2131_p
  (
    .dout(g2131_p),
    .din1(G12_p_spl_01),
    .din2(G20_p_spl_100)
  );


  orX
  g_g2131_n
  (
    .dout(g2131_n),
    .din1(G12_n_spl_1),
    .din2(G20_n_spl_101)
  );


  andX
  g_g2132_p
  (
    .dout(g2132_p),
    .din1(g2117_n_spl_),
    .din2(g2120_n_spl_)
  );


  orX
  g_g2132_n
  (
    .dout(g2132_n),
    .din1(g2117_p_spl_),
    .din2(g2120_p_spl_)
  );


  andX
  g_g2133_p
  (
    .dout(g2133_p),
    .din1(G13_p_spl_01),
    .din2(G19_p_spl_110)
  );


  orX
  g_g2133_n
  (
    .dout(g2133_n),
    .din1(G13_n_spl_1),
    .din2(G19_n_spl_110)
  );


  andX
  g_g2134_p
  (
    .dout(g2134_p),
    .din1(G15_p_spl_00),
    .din2(G17_p_spl_110)
  );


  orX
  g_g2134_n
  (
    .dout(g2134_n),
    .din1(G15_n_spl_0),
    .din2(G17_n_spl_110)
  );


  andX
  g_g2135_p
  (
    .dout(g2135_p),
    .din1(G14_p_spl_00),
    .din2(G18_p_spl_110)
  );


  orX
  g_g2135_n
  (
    .dout(g2135_n),
    .din1(G14_n_spl_0),
    .din2(G18_n_spl_110)
  );


  andX
  g_g2136_p
  (
    .dout(g2136_p),
    .din1(g2134_p_spl_),
    .din2(g2135_p_spl_)
  );


  orX
  g_g2136_n
  (
    .dout(g2136_n),
    .din1(g2134_n_spl_),
    .din2(g2135_n_spl_)
  );


  andX
  g_g2137_p
  (
    .dout(g2137_p),
    .din1(g2134_n_spl_),
    .din2(g2135_n_spl_)
  );


  orX
  g_g2137_n
  (
    .dout(g2137_n),
    .din1(g2134_p_spl_),
    .din2(g2135_p_spl_)
  );


  andX
  g_g2138_p
  (
    .dout(g2138_p),
    .din1(g2136_n_spl_0),
    .din2(g2137_n)
  );


  orX
  g_g2138_n
  (
    .dout(g2138_n),
    .din1(g2136_p_spl_0),
    .din2(g2137_p)
  );


  andX
  g_g2139_p
  (
    .dout(g2139_p),
    .din1(g2114_n_spl_0),
    .din2(g2138_n_spl_)
  );


  orX
  g_g2139_n
  (
    .dout(g2139_n),
    .din1(g2114_p_spl_0),
    .din2(g2138_p_spl_)
  );


  andX
  g_g2140_p
  (
    .dout(g2140_p),
    .din1(g2114_p_spl_),
    .din2(g2138_p_spl_)
  );


  orX
  g_g2140_n
  (
    .dout(g2140_n),
    .din1(g2114_n_spl_),
    .din2(g2138_n_spl_)
  );


  andX
  g_g2141_p
  (
    .dout(g2141_p),
    .din1(g2139_n_spl_),
    .din2(g2140_n)
  );


  orX
  g_g2141_n
  (
    .dout(g2141_n),
    .din1(g2139_p_spl_),
    .din2(g2140_p)
  );


  andX
  g_g2142_p
  (
    .dout(g2142_p),
    .din1(g2133_n_spl_),
    .din2(g2141_p_spl_)
  );


  orX
  g_g2142_n
  (
    .dout(g2142_n),
    .din1(g2133_p_spl_),
    .din2(g2141_n_spl_)
  );


  andX
  g_g2143_p
  (
    .dout(g2143_p),
    .din1(g2133_p_spl_),
    .din2(g2141_n_spl_)
  );


  orX
  g_g2143_n
  (
    .dout(g2143_n),
    .din1(g2133_n_spl_),
    .din2(g2141_p_spl_)
  );


  andX
  g_g2144_p
  (
    .dout(g2144_p),
    .din1(g2142_n_spl_),
    .din2(g2143_n)
  );


  orX
  g_g2144_n
  (
    .dout(g2144_n),
    .din1(g2142_p_spl_),
    .din2(g2143_p)
  );


  andX
  g_g2145_p
  (
    .dout(g2145_p),
    .din1(g2132_n_spl_),
    .din2(g2144_p_spl_)
  );


  orX
  g_g2145_n
  (
    .dout(g2145_n),
    .din1(g2132_p_spl_),
    .din2(g2144_n_spl_)
  );


  andX
  g_g2146_p
  (
    .dout(g2146_p),
    .din1(g2132_p_spl_),
    .din2(g2144_n_spl_)
  );


  orX
  g_g2146_n
  (
    .dout(g2146_n),
    .din1(g2132_n_spl_),
    .din2(g2144_p_spl_)
  );


  andX
  g_g2147_p
  (
    .dout(g2147_p),
    .din1(g2145_n_spl_),
    .din2(g2146_n)
  );


  orX
  g_g2147_n
  (
    .dout(g2147_n),
    .din1(g2145_p_spl_),
    .din2(g2146_p)
  );


  andX
  g_g2148_p
  (
    .dout(g2148_p),
    .din1(g2131_n_spl_),
    .din2(g2147_p_spl_)
  );


  orX
  g_g2148_n
  (
    .dout(g2148_n),
    .din1(g2131_p_spl_),
    .din2(g2147_n_spl_)
  );


  andX
  g_g2149_p
  (
    .dout(g2149_p),
    .din1(g2131_p_spl_),
    .din2(g2147_n_spl_)
  );


  orX
  g_g2149_n
  (
    .dout(g2149_n),
    .din1(g2131_n_spl_),
    .din2(g2147_p_spl_)
  );


  andX
  g_g2150_p
  (
    .dout(g2150_p),
    .din1(g2148_n_spl_),
    .din2(g2149_n)
  );


  orX
  g_g2150_n
  (
    .dout(g2150_n),
    .din1(g2148_p_spl_),
    .din2(g2149_p)
  );


  orX
  g_g2151_n
  (
    .dout(g2151_n),
    .din1(g2130_p),
    .din2(g2150_n)
  );


  andX
  g_g2152_p
  (
    .dout(g2152_p),
    .din1(g2145_n_spl_),
    .din2(g2148_n_spl_)
  );


  orX
  g_g2152_n
  (
    .dout(g2152_n),
    .din1(g2145_p_spl_),
    .din2(g2148_p_spl_)
  );


  andX
  g_g2153_p
  (
    .dout(g2153_p),
    .din1(G13_p_spl_01),
    .din2(G20_p_spl_101)
  );


  orX
  g_g2153_n
  (
    .dout(g2153_n),
    .din1(G13_n_spl_1),
    .din2(G20_n_spl_101)
  );


  andX
  g_g2154_p
  (
    .dout(g2154_p),
    .din1(g2139_n_spl_),
    .din2(g2142_n_spl_)
  );


  orX
  g_g2154_n
  (
    .dout(g2154_n),
    .din1(g2139_p_spl_),
    .din2(g2142_p_spl_)
  );


  andX
  g_g2155_p
  (
    .dout(g2155_p),
    .din1(G14_p_spl_01),
    .din2(G19_p_spl_110)
  );


  orX
  g_g2155_n
  (
    .dout(g2155_n),
    .din1(G14_n_spl_1),
    .din2(G19_n_spl_110)
  );


  andX
  g_g2156_p
  (
    .dout(g2156_p),
    .din1(G16_p_spl_00),
    .din2(G17_p_spl_111)
  );


  orX
  g_g2156_n
  (
    .dout(g2156_n),
    .din1(G16_n_spl_0),
    .din2(G17_n_spl_11)
  );


  andX
  g_g2157_p
  (
    .dout(g2157_p),
    .din1(G15_p_spl_00),
    .din2(G18_p_spl_111)
  );


  orX
  g_g2157_n
  (
    .dout(g2157_n),
    .din1(G15_n_spl_0),
    .din2(G18_n_spl_111)
  );


  andX
  g_g2158_p
  (
    .dout(g2158_p),
    .din1(g2156_p_spl_),
    .din2(g2157_p_spl_)
  );


  orX
  g_g2158_n
  (
    .dout(g2158_n),
    .din1(g2156_n_spl_),
    .din2(g2157_n_spl_)
  );


  andX
  g_g2159_p
  (
    .dout(g2159_p),
    .din1(g2156_n_spl_),
    .din2(g2157_n_spl_)
  );


  orX
  g_g2159_n
  (
    .dout(g2159_n),
    .din1(g2156_p_spl_),
    .din2(g2157_p_spl_)
  );


  andX
  g_g2160_p
  (
    .dout(g2160_p),
    .din1(g2158_n_spl_),
    .din2(g2159_n)
  );


  orX
  g_g2160_n
  (
    .dout(g2160_n),
    .din1(g2158_p_spl_),
    .din2(g2159_p)
  );


  andX
  g_g2161_p
  (
    .dout(g2161_p),
    .din1(g2136_n_spl_0),
    .din2(g2160_n_spl_)
  );


  orX
  g_g2161_n
  (
    .dout(g2161_n),
    .din1(g2136_p_spl_0),
    .din2(g2160_p_spl_)
  );


  andX
  g_g2162_p
  (
    .dout(g2162_p),
    .din1(g2136_p_spl_),
    .din2(g2160_p_spl_)
  );


  orX
  g_g2162_n
  (
    .dout(g2162_n),
    .din1(g2136_n_spl_),
    .din2(g2160_n_spl_)
  );


  andX
  g_g2163_p
  (
    .dout(g2163_p),
    .din1(g2161_n_spl_),
    .din2(g2162_n)
  );


  orX
  g_g2163_n
  (
    .dout(g2163_n),
    .din1(g2161_p_spl_),
    .din2(g2162_p)
  );


  andX
  g_g2164_p
  (
    .dout(g2164_p),
    .din1(g2155_n_spl_),
    .din2(g2163_p_spl_)
  );


  orX
  g_g2164_n
  (
    .dout(g2164_n),
    .din1(g2155_p_spl_),
    .din2(g2163_n_spl_)
  );


  andX
  g_g2165_p
  (
    .dout(g2165_p),
    .din1(g2155_p_spl_),
    .din2(g2163_n_spl_)
  );


  orX
  g_g2165_n
  (
    .dout(g2165_n),
    .din1(g2155_n_spl_),
    .din2(g2163_p_spl_)
  );


  andX
  g_g2166_p
  (
    .dout(g2166_p),
    .din1(g2164_n_spl_),
    .din2(g2165_n)
  );


  orX
  g_g2166_n
  (
    .dout(g2166_n),
    .din1(g2164_p_spl_),
    .din2(g2165_p)
  );


  andX
  g_g2167_p
  (
    .dout(g2167_p),
    .din1(g2154_n_spl_),
    .din2(g2166_p_spl_)
  );


  orX
  g_g2167_n
  (
    .dout(g2167_n),
    .din1(g2154_p_spl_),
    .din2(g2166_n_spl_)
  );


  andX
  g_g2168_p
  (
    .dout(g2168_p),
    .din1(g2154_p_spl_),
    .din2(g2166_n_spl_)
  );


  orX
  g_g2168_n
  (
    .dout(g2168_n),
    .din1(g2154_n_spl_),
    .din2(g2166_p_spl_)
  );


  andX
  g_g2169_p
  (
    .dout(g2169_p),
    .din1(g2167_n_spl_),
    .din2(g2168_n)
  );


  orX
  g_g2169_n
  (
    .dout(g2169_n),
    .din1(g2167_p_spl_),
    .din2(g2168_p)
  );


  andX
  g_g2170_p
  (
    .dout(g2170_p),
    .din1(g2153_n_spl_),
    .din2(g2169_p_spl_)
  );


  orX
  g_g2170_n
  (
    .dout(g2170_n),
    .din1(g2153_p_spl_),
    .din2(g2169_n_spl_)
  );


  andX
  g_g2171_p
  (
    .dout(g2171_p),
    .din1(g2153_p_spl_),
    .din2(g2169_n_spl_)
  );


  orX
  g_g2171_n
  (
    .dout(g2171_n),
    .din1(g2153_n_spl_),
    .din2(g2169_p_spl_)
  );


  andX
  g_g2172_p
  (
    .dout(g2172_p),
    .din1(g2170_n_spl_),
    .din2(g2171_n)
  );


  orX
  g_g2172_n
  (
    .dout(g2172_n),
    .din1(g2170_p_spl_),
    .din2(g2171_p)
  );


  orX
  g_g2173_n
  (
    .dout(g2173_n),
    .din1(g2152_p),
    .din2(g2172_n)
  );


  andX
  g_g2174_p
  (
    .dout(g2174_p),
    .din1(g2167_n_spl_),
    .din2(g2170_n_spl_)
  );


  orX
  g_g2174_n
  (
    .dout(g2174_n),
    .din1(g2167_p_spl_),
    .din2(g2170_p_spl_)
  );


  andX
  g_g2175_p
  (
    .dout(g2175_p),
    .din1(G14_p_spl_01),
    .din2(G20_p_spl_101)
  );


  orX
  g_g2175_n
  (
    .dout(g2175_n),
    .din1(G14_n_spl_1),
    .din2(G20_n_spl_110)
  );


  andX
  g_g2176_p
  (
    .dout(g2176_p),
    .din1(g2161_n_spl_),
    .din2(g2164_n_spl_)
  );


  orX
  g_g2176_n
  (
    .dout(g2176_n),
    .din1(g2161_p_spl_),
    .din2(g2164_p_spl_)
  );


  andX
  g_g2177_p
  (
    .dout(g2177_p),
    .din1(G16_p_spl_00),
    .din2(G18_p_spl_111)
  );


  orX
  g_g2177_n
  (
    .dout(g2177_n),
    .din1(G16_n_spl_0),
    .din2(G18_n_spl_111)
  );


  andX
  g_g2178_p
  (
    .dout(g2178_p),
    .din1(g2158_n_spl_),
    .din2(g2177_p_spl_)
  );


  orX
  g_g2178_n
  (
    .dout(g2178_n),
    .din1(g2158_p_spl_),
    .din2(g2177_n_spl_)
  );


  andX
  g_g2179_p
  (
    .dout(g2179_p),
    .din1(G15_p_spl_0),
    .din2(G19_p_spl_111)
  );


  orX
  g_g2179_n
  (
    .dout(g2179_n),
    .din1(G15_n_spl_1),
    .din2(G19_n_spl_111)
  );


  andX
  g_g2180_p
  (
    .dout(g2180_p),
    .din1(g2178_p_spl_),
    .din2(g2179_n_spl_)
  );


  orX
  g_g2180_n
  (
    .dout(g2180_n),
    .din1(g2178_n_spl_),
    .din2(g2179_p_spl_)
  );


  andX
  g_g2181_p
  (
    .dout(g2181_p),
    .din1(g2178_n_spl_),
    .din2(g2179_p_spl_)
  );


  orX
  g_g2181_n
  (
    .dout(g2181_n),
    .din1(g2178_p_spl_),
    .din2(g2179_n_spl_)
  );


  andX
  g_g2182_p
  (
    .dout(g2182_p),
    .din1(g2180_n_spl_),
    .din2(g2181_n)
  );


  orX
  g_g2182_n
  (
    .dout(g2182_n),
    .din1(g2180_p_spl_),
    .din2(g2181_p)
  );


  andX
  g_g2183_p
  (
    .dout(g2183_p),
    .din1(g2176_n_spl_),
    .din2(g2182_p_spl_)
  );


  orX
  g_g2183_n
  (
    .dout(g2183_n),
    .din1(g2176_p_spl_),
    .din2(g2182_n_spl_)
  );


  andX
  g_g2184_p
  (
    .dout(g2184_p),
    .din1(g2176_p_spl_),
    .din2(g2182_n_spl_)
  );


  orX
  g_g2184_n
  (
    .dout(g2184_n),
    .din1(g2176_n_spl_),
    .din2(g2182_p_spl_)
  );


  andX
  g_g2185_p
  (
    .dout(g2185_p),
    .din1(g2183_n_spl_),
    .din2(g2184_n)
  );


  orX
  g_g2185_n
  (
    .dout(g2185_n),
    .din1(g2183_p_spl_),
    .din2(g2184_p)
  );


  andX
  g_g2186_p
  (
    .dout(g2186_p),
    .din1(g2175_n_spl_),
    .din2(g2185_p_spl_)
  );


  orX
  g_g2186_n
  (
    .dout(g2186_n),
    .din1(g2175_p_spl_),
    .din2(g2185_n_spl_)
  );


  andX
  g_g2187_p
  (
    .dout(g2187_p),
    .din1(g2175_p_spl_),
    .din2(g2185_n_spl_)
  );


  orX
  g_g2187_n
  (
    .dout(g2187_n),
    .din1(g2175_n_spl_),
    .din2(g2185_p_spl_)
  );


  andX
  g_g2188_p
  (
    .dout(g2188_p),
    .din1(g2186_n_spl_),
    .din2(g2187_n)
  );


  orX
  g_g2188_n
  (
    .dout(g2188_n),
    .din1(g2186_p_spl_),
    .din2(g2187_p)
  );


  orX
  g_g2189_n
  (
    .dout(g2189_n),
    .din1(g2174_p),
    .din2(g2188_n)
  );


  andX
  g_g2190_p
  (
    .dout(g2190_p),
    .din1(g2183_n_spl_),
    .din2(g2186_n_spl_)
  );


  orX
  g_g2190_n
  (
    .dout(g2190_n),
    .din1(g2183_p_spl_),
    .din2(g2186_p_spl_)
  );


  andX
  g_g2191_p
  (
    .dout(g2191_p),
    .din1(G15_p_spl_1),
    .din2(G20_p_spl_110)
  );


  orX
  g_g2191_n
  (
    .dout(g2191_n),
    .din1(G15_n_spl_1),
    .din2(G20_n_spl_110)
  );


  andX
  g_g2192_p
  (
    .dout(g2192_p),
    .din1(G16_p_spl_0),
    .din2(G19_p_spl_111)
  );


  orX
  g_g2192_n
  (
    .dout(g2192_n),
    .din1(G16_n_spl_),
    .din2(G19_n_spl_111)
  );


  andX
  g_g2193_p
  (
    .dout(g2193_p),
    .din1(g2177_p_spl_),
    .din2(g2180_n_spl_)
  );


  orX
  g_g2193_n
  (
    .dout(g2193_n),
    .din1(g2177_n_spl_),
    .din2(g2180_p_spl_)
  );


  andX
  g_g2194_p
  (
    .dout(g2194_p),
    .din1(g2192_n_spl_),
    .din2(g2193_n_spl_)
  );


  orX
  g_g2194_n
  (
    .dout(g2194_n),
    .din1(g2192_p_spl_),
    .din2(g2193_p_spl_)
  );


  andX
  g_g2195_p
  (
    .dout(g2195_p),
    .din1(g2192_p_spl_),
    .din2(g2193_p_spl_)
  );


  orX
  g_g2195_n
  (
    .dout(g2195_n),
    .din1(g2192_n_spl_),
    .din2(g2193_n_spl_)
  );


  andX
  g_g2196_p
  (
    .dout(g2196_p),
    .din1(g2194_n_spl_),
    .din2(g2195_n)
  );


  orX
  g_g2196_n
  (
    .dout(g2196_n),
    .din1(g2194_p),
    .din2(g2195_p)
  );


  andX
  g_g2197_p
  (
    .dout(g2197_p),
    .din1(g2191_n_spl_),
    .din2(g2196_p_spl_)
  );


  orX
  g_g2197_n
  (
    .dout(g2197_n),
    .din1(g2191_p_spl_),
    .din2(g2196_n_spl_)
  );


  andX
  g_g2198_p
  (
    .dout(g2198_p),
    .din1(g2191_p_spl_),
    .din2(g2196_n_spl_)
  );


  orX
  g_g2198_n
  (
    .dout(g2198_n),
    .din1(g2191_n_spl_),
    .din2(g2196_p_spl_)
  );


  andX
  g_g2199_p
  (
    .dout(g2199_p),
    .din1(g2197_n_spl_),
    .din2(g2198_n)
  );


  orX
  g_g2199_n
  (
    .dout(g2199_n),
    .din1(g2197_p),
    .din2(g2198_p)
  );


  orX
  g_g2200_n
  (
    .dout(g2200_n),
    .din1(g2190_p),
    .din2(g2199_n)
  );


  andX
  g_g2201_p
  (
    .dout(g2201_p),
    .din1(g1585_n_spl_),
    .din2(g1588_n_spl_)
  );


  orX
  g_g2201_n
  (
    .dout(g2201_n),
    .din1(g1585_p_spl_),
    .din2(g1588_p_spl_)
  );


  andX
  g_g2202_p
  (
    .dout(g2202_p),
    .din1(g1932_p_spl_),
    .din2(g1934_n_spl_)
  );


  orX
  g_g2202_n
  (
    .dout(g2202_n),
    .din1(g1932_n_spl_),
    .din2(g1934_p_spl_)
  );


  andX
  g_g2203_p
  (
    .dout(g2203_p),
    .din1(g1935_n_spl_),
    .din2(g2202_n)
  );


  orX
  g_g2203_n
  (
    .dout(g2203_n),
    .din1(g1935_p_spl_),
    .din2(g2202_p)
  );


  andX
  g_g2204_p
  (
    .dout(g2204_p),
    .din1(g2201_n_spl_),
    .din2(g2203_p_spl_)
  );


  orX
  g_g2204_n
  (
    .dout(g2204_n),
    .din1(g2201_p_spl_),
    .din2(g2203_n_spl_)
  );


  andX
  g_g2205_p
  (
    .dout(g2205_p),
    .din1(G2_p_spl_01),
    .din2(G20_p_spl_110)
  );


  orX
  g_g2205_n
  (
    .dout(g2205_n),
    .din1(G2_n_spl_1),
    .din2(G20_n_spl_11)
  );


  andX
  g_g2206_p
  (
    .dout(g2206_p),
    .din1(g2201_p_spl_),
    .din2(g2203_n_spl_)
  );


  orX
  g_g2206_n
  (
    .dout(g2206_n),
    .din1(g2201_n_spl_),
    .din2(g2203_p_spl_)
  );


  andX
  g_g2207_p
  (
    .dout(g2207_p),
    .din1(g2204_n_spl_),
    .din2(g2206_n)
  );


  orX
  g_g2207_n
  (
    .dout(g2207_n),
    .din1(g2204_p_spl_),
    .din2(g2206_p)
  );


  andX
  g_g2208_p
  (
    .dout(g2208_p),
    .din1(g2205_n_spl_),
    .din2(g2207_p_spl_)
  );


  orX
  g_g2208_n
  (
    .dout(g2208_n),
    .din1(g2205_p),
    .din2(g2207_n)
  );


  andX
  g_g2209_p
  (
    .dout(g2209_p),
    .din1(g2204_n_spl_),
    .din2(g2208_n_spl_)
  );


  orX
  g_g2209_n
  (
    .dout(g2209_n),
    .din1(g2204_p_spl_),
    .din2(g2208_p)
  );


  andX
  g_g2210_p
  (
    .dout(g2210_p),
    .din1(g1950_p_spl_),
    .din2(g1952_n_spl_)
  );


  orX
  g_g2210_n
  (
    .dout(g2210_n),
    .din1(g1950_n_spl_),
    .din2(g1952_p_spl_)
  );


  andX
  g_g2211_p
  (
    .dout(g2211_p),
    .din1(g1953_n_spl_),
    .din2(g2210_n)
  );


  orX
  g_g2211_n
  (
    .dout(g2211_n),
    .din1(g1953_p_spl_),
    .din2(g2210_p)
  );


  orX
  g_g2212_n
  (
    .dout(g2212_n),
    .din1(g2209_p),
    .din2(g2211_n)
  );


  andX
  g_g2213_p
  (
    .dout(g2213_p),
    .din1(G3_p_spl_1),
    .din2(G21_p_spl_000)
  );


  andX
  g_g2214_p
  (
    .dout(g2214_p),
    .din1(G4_p_spl_1),
    .din2(G21_p_spl_000)
  );


  andX
  g_g2215_p
  (
    .dout(g2215_p),
    .din1(G5_p_spl_1),
    .din2(G21_p_spl_001)
  );


  andX
  g_g2216_p
  (
    .dout(g2216_p),
    .din1(G6_p_spl_1),
    .din2(G21_p_spl_001)
  );


  andX
  g_g2217_p
  (
    .dout(g2217_p),
    .din1(G7_p_spl_1),
    .din2(G21_p_spl_010)
  );


  andX
  g_g2218_p
  (
    .dout(g2218_p),
    .din1(G8_p_spl_1),
    .din2(G21_p_spl_010)
  );


  andX
  g_g2219_p
  (
    .dout(g2219_p),
    .din1(G9_p_spl_1),
    .din2(G21_p_spl_011)
  );


  andX
  g_g2220_p
  (
    .dout(g2220_p),
    .din1(G10_p_spl_1),
    .din2(G21_p_spl_011)
  );


  andX
  g_g2221_p
  (
    .dout(g2221_p),
    .din1(G11_p_spl_1),
    .din2(G21_p_spl_100)
  );


  andX
  g_g2222_p
  (
    .dout(g2222_p),
    .din1(G12_p_spl_1),
    .din2(G21_p_spl_100)
  );


  andX
  g_g2223_p
  (
    .dout(g2223_p),
    .din1(G13_p_spl_1),
    .din2(G21_p_spl_101)
  );


  andX
  g_g2224_p
  (
    .dout(g2224_p),
    .din1(G14_p_spl_1),
    .din2(G21_p_spl_101)
  );


  andX
  g_g2225_p
  (
    .dout(g2225_p),
    .din1(G16_p_spl_1),
    .din2(G20_p_spl_11)
  );


  andX
  g_g2226_p
  (
    .dout(g2226_p),
    .din1(G2_p_spl_1),
    .din2(G21_p_spl_11)
  );


  andX
  g_g2227_p
  (
    .dout(g2227_p),
    .din1(g2194_n_spl_),
    .din2(g2197_n_spl_)
  );


  orX
  g_g2228_n
  (
    .dout(g2228_n),
    .din1(g1591_p),
    .din2(g1631_p_spl_)
  );


  orX
  g_g2229_n
  (
    .dout(g2229_n),
    .din1(g2205_n_spl_),
    .din2(g2207_p_spl_)
  );


  andX
  g_g2230_p
  (
    .dout(g2230_p),
    .din1(g2208_n_spl_),
    .din2(g2229_n)
  );


  andX
  g_g2231_p
  (
    .dout(g2231_p),
    .din1(g2228_n_spl_),
    .din2(g2230_p_spl_)
  );


  orX
  g_g2232_n
  (
    .dout(g2232_n),
    .din1(g2228_n_spl_),
    .din2(g2230_p_spl_)
  );


  orX
  g_g2233_n
  (
    .dout(g2233_n),
    .din1(g1954_n),
    .din2(g1974_p)
  );


  andX
  g_g2234_p
  (
    .dout(g2234_p),
    .din1(g1975_n_spl_),
    .din2(g2233_n)
  );


  orX
  g_g2235_n
  (
    .dout(g2235_n),
    .din1(g1976_n),
    .din2(g1996_p)
  );


  andX
  g_g2236_p
  (
    .dout(g2236_p),
    .din1(g1997_n_spl_),
    .din2(g2235_n)
  );


  orX
  g_g2237_n
  (
    .dout(g2237_n),
    .din1(g1998_n),
    .din2(g2018_p)
  );


  andX
  g_g2238_p
  (
    .dout(g2238_p),
    .din1(g2019_n_spl_),
    .din2(g2237_n)
  );


  orX
  g_g2239_n
  (
    .dout(g2239_n),
    .din1(g2020_n),
    .din2(g2040_p)
  );


  andX
  g_g2240_p
  (
    .dout(g2240_p),
    .din1(g2041_n_spl_),
    .din2(g2239_n)
  );


  orX
  g_g2241_n
  (
    .dout(g2241_n),
    .din1(g2042_n),
    .din2(g2062_p)
  );


  andX
  g_g2242_p
  (
    .dout(g2242_p),
    .din1(g2063_n_spl_),
    .din2(g2241_n)
  );


  orX
  g_g2243_n
  (
    .dout(g2243_n),
    .din1(g2064_n),
    .din2(g2084_p)
  );


  andX
  g_g2244_p
  (
    .dout(g2244_p),
    .din1(g2085_n_spl_),
    .din2(g2243_n)
  );


  orX
  g_g2245_n
  (
    .dout(g2245_n),
    .din1(g2086_n),
    .din2(g2106_p)
  );


  andX
  g_g2246_p
  (
    .dout(g2246_p),
    .din1(g2107_n_spl_),
    .din2(g2245_n)
  );


  orX
  g_g2247_n
  (
    .dout(g2247_n),
    .din1(g2108_n),
    .din2(g2128_p)
  );


  andX
  g_g2248_p
  (
    .dout(g2248_p),
    .din1(g2129_n_spl_),
    .din2(g2247_n)
  );


  orX
  g_g2249_n
  (
    .dout(g2249_n),
    .din1(g2130_n),
    .din2(g2150_p)
  );


  andX
  g_g2250_p
  (
    .dout(g2250_p),
    .din1(g2151_n_spl_),
    .din2(g2249_n)
  );


  orX
  g_g2251_n
  (
    .dout(g2251_n),
    .din1(g2152_n),
    .din2(g2172_p)
  );


  andX
  g_g2252_p
  (
    .dout(g2252_p),
    .din1(g2173_n_spl_),
    .din2(g2251_n)
  );


  orX
  g_g2253_n
  (
    .dout(g2253_n),
    .din1(g2174_n),
    .din2(g2188_p)
  );


  andX
  g_g2254_p
  (
    .dout(g2254_p),
    .din1(g2189_n_spl_),
    .din2(g2253_n)
  );


  orX
  g_g2255_n
  (
    .dout(g2255_n),
    .din1(g2190_n),
    .din2(g2199_p)
  );


  andX
  g_g2256_p
  (
    .dout(g2256_p),
    .din1(g2200_n_spl_),
    .din2(g2255_n)
  );


  orX
  g_g2257_n
  (
    .dout(g2257_n),
    .din1(g2209_n),
    .din2(g2211_p)
  );


  andX
  g_g2258_p
  (
    .dout(g2258_p),
    .din1(g2212_n_spl_),
    .din2(g2257_n)
  );


  buf

  (
    G6257_p,
    g389_p
  );


  buf

  (
    G6258_p,
    g391_p
  );


  buf

  (
    G6259_p,
    g393_n
  );


  buf

  (
    G6260_p,
    g395_n
  );


  buf

  (
    G6261_p,
    g397_n
  );


  buf

  (
    G6262_p,
    g399_n
  );


  buf

  (
    G6263_p,
    g401_n
  );


  buf

  (
    G6264_p,
    g403_n
  );


  buf

  (
    G6265_p,
    g405_n
  );


  buf

  (
    G6266_p,
    g407_n
  );


  buf

  (
    G6267_p,
    g409_n
  );


  buf

  (
    G6268_p,
    g411_n
  );


  buf

  (
    G6269_p,
    g413_n
  );


  buf

  (
    G6270_p,
    g415_n
  );


  buf

  (
    G6271_p,
    g417_n
  );


  buf

  (
    G6272_p,
    g419_n
  );


  buf

  (
    G6273_p,
    g421_p
  );


  buf

  (
    G6274_p,
    g423_n
  );


  buf

  (
    G6275_p,
    g425_n
  );


  buf

  (
    G6276_p,
    g427_n
  );


  buf

  (
    G6277_p,
    g429_n
  );


  buf

  (
    G6278_p,
    g431_n
  );


  buf

  (
    G6279_p,
    g436_n
  );


  buf

  (
    G6280_p,
    g445_n
  );


  buf

  (
    G6281_p,
    g458_n
  );


  buf

  (
    G6282_p,
    g475_n
  );


  buf

  (
    G6283_p,
    g496_n
  );


  buf

  (
    G6284_p,
    g521_n
  );


  buf

  (
    G6285_p,
    g546_n
  );


  buf

  (
    G6286_p,
    g563_n
  );


  buf

  (
    G6287_p,
    g571_p
  );


  buf

  (
    G6288_n,
    g573_p
  );


  DROC
  ffc_0
  (
    .doutp(ffc_0_p),
    .doutn(ffc_0_n),
    .din(ffc_80_p_spl_)
  );


  DROC
  ffc_1
  (
    .doutp(ffc_1_p),
    .doutn(ffc_1_n),
    .din(ffc_71_p_spl_1)
  );


  DROC
  ffc_2
  (
    .doutp(ffc_2_p),
    .doutn(ffc_2_n),
    .din(ffc_72_p_spl_1)
  );


  DROC
  ffc_3
  (
    .doutp(ffc_3_p),
    .doutn(ffc_3_n),
    .din(ffc_73_p_spl_)
  );


  DROC
  ffc_4
  (
    .doutp(ffc_4_p),
    .doutn(ffc_4_n),
    .din(ffc_74_p_spl_1)
  );


  DROC
  ffc_5
  (
    .doutp(ffc_5_p),
    .doutn(ffc_5_n),
    .din(ffc_75_p_spl_1)
  );


  DROC
  ffc_6
  (
    .doutp(ffc_6_p),
    .doutn(ffc_6_n),
    .din(ffc_76_p_spl_)
  );


  DROC
  ffc_7
  (
    .doutp(ffc_7_p),
    .doutn(ffc_7_n),
    .din(ffc_77_p_spl_1)
  );


  DROC
  ffc_8
  (
    .doutp(ffc_8_p),
    .doutn(ffc_8_n),
    .din(ffc_78_p)
  );


  DROC
  ffc_9
  (
    .doutp(ffc_9_p),
    .doutn(ffc_9_n),
    .din(G22_p)
  );


  DROC
  ffc_10
  (
    .doutp(ffc_10_p),
    .doutn(ffc_10_n),
    .din(G23_p)
  );


  DROC
  ffc_11
  (
    .doutp(ffc_11_p),
    .doutn(ffc_11_n),
    .din(G24_p)
  );


  DROC
  ffc_12
  (
    .doutp(ffc_12_p),
    .doutn(ffc_12_n),
    .din(G25_p)
  );


  DROC
  ffc_13
  (
    .doutp(ffc_13_p),
    .doutn(ffc_13_n),
    .din(G26_p)
  );


  DROC
  ffc_14
  (
    .doutp(ffc_14_p),
    .doutn(ffc_14_n),
    .din(G27_p)
  );


  DROC
  ffc_15
  (
    .doutp(ffc_15_p),
    .doutn(ffc_15_n),
    .din(ffc_14_p)
  );


  DROC
  ffc_16
  (
    .doutp(ffc_16_p),
    .doutn(ffc_16_n),
    .din(G28_p)
  );


  DROC
  ffc_17
  (
    .doutp(ffc_17_p),
    .doutn(ffc_17_n),
    .din(ffc_16_p)
  );


  DROC
  ffc_18
  (
    .doutp(ffc_18_p),
    .doutn(ffc_18_n),
    .din(G29_p)
  );


  DROC
  ffc_19
  (
    .doutp(ffc_19_p),
    .doutn(ffc_19_n),
    .din(ffc_18_p)
  );


  DROC
  ffc_20
  (
    .doutp(ffc_20_p),
    .doutn(ffc_20_n),
    .din(G30_p)
  );


  DROC
  ffc_21
  (
    .doutp(ffc_21_p),
    .doutn(ffc_21_n),
    .din(ffc_20_p)
  );


  DROC
  ffc_22
  (
    .doutp(ffc_22_p),
    .doutn(ffc_22_n),
    .din(ffc_214_p_spl_11)
  );


  DROC
  ffc_23
  (
    .doutp(ffc_23_p),
    .doutn(ffc_23_n),
    .din(G31_p)
  );


  DROC
  ffc_24
  (
    .doutp(ffc_24_p),
    .doutn(ffc_24_n),
    .din(ffc_23_p)
  );


  DROC
  ffc_25
  (
    .doutp(ffc_25_p),
    .doutn(ffc_25_n),
    .din(ffc_24_p)
  );


  DROC
  ffc_26
  (
    .doutp(ffc_26_p),
    .doutn(ffc_26_n),
    .din(ffc_25_p_spl_11)
  );


  DROC
  ffc_27
  (
    .doutp(ffc_27_p),
    .doutn(ffc_27_n),
    .din(G32_p)
  );


  DROC
  ffc_28
  (
    .doutp(ffc_28_p),
    .doutn(ffc_28_n),
    .din(ffc_27_p)
  );


  DROC
  ffc_29
  (
    .doutp(ffc_29_p),
    .doutn(ffc_29_n),
    .din(ffc_28_p)
  );


  DROC
  ffc_30
  (
    .doutp(ffc_30_p),
    .doutn(ffc_30_n),
    .din(ffc_29_p_spl_11)
  );


  DROC
  ffc_31
  (
    .doutp(ffc_31_p),
    .doutn(ffc_31_n),
    .din(ffc_84_p)
  );


  DROC
  ffc_32
  (
    .doutp(ffc_32_p),
    .doutn(ffc_32_n),
    .din(ffc_83_p)
  );


  DROC
  ffc_33
  (
    .doutp(ffc_33_p),
    .doutn(ffc_33_n),
    .din(ffc_86_p)
  );


  DROC
  ffc_34
  (
    .doutp(ffc_34_p),
    .doutn(ffc_34_n),
    .din(ffc_87_p)
  );


  DROC
  ffc_35
  (
    .doutp(ffc_35_p),
    .doutn(ffc_35_n),
    .din(ffc_88_p)
  );


  DROC
  ffc_36
  (
    .doutp(ffc_36_p),
    .doutn(ffc_36_n),
    .din(ffc_89_p)
  );


  DROC
  ffc_37
  (
    .doutp(ffc_37_p),
    .doutn(ffc_37_n),
    .din(ffc_91_p)
  );


  DROC
  ffc_38
  (
    .doutp(ffc_38_p),
    .doutn(ffc_38_n),
    .din(ffc_93_p)
  );


  DROC
  ffc_39
  (
    .doutp(ffc_39_p),
    .doutn(ffc_39_n),
    .din(ffc_94_p)
  );


  DROC
  ffc_40
  (
    .doutp(ffc_40_p),
    .doutn(ffc_40_n),
    .din(ffc_96_p)
  );


  DROC
  ffc_41
  (
    .doutp(ffc_41_p),
    .doutn(ffc_41_n),
    .din(ffc_97_p)
  );


  DROC
  ffc_42
  (
    .doutp(ffc_42_p),
    .doutn(ffc_42_n),
    .din(ffc_98_p)
  );


  DROC
  ffc_43
  (
    .doutp(ffc_43_p),
    .doutn(ffc_43_n),
    .din(ffc_100_p)
  );


  DROC
  ffc_44
  (
    .doutp(ffc_44_p),
    .doutn(ffc_44_n),
    .din(ffc_102_p)
  );


  DROC
  ffc_45
  (
    .doutp(ffc_45_p),
    .doutn(ffc_45_n),
    .din(ffc_103_p)
  );


  DROC
  ffc_46
  (
    .doutp(ffc_46_p),
    .doutn(ffc_46_n),
    .din(ffc_105_p)
  );


  DROC
  ffc_47
  (
    .doutp(ffc_47_p),
    .doutn(ffc_47_n),
    .din(ffc_106_p)
  );


  DROC
  ffc_48
  (
    .doutp(ffc_48_p),
    .doutn(ffc_48_n),
    .din(ffc_107_p)
  );


  DROC
  ffc_49
  (
    .doutp(ffc_49_p),
    .doutn(ffc_49_n),
    .din(ffc_109_p)
  );


  DROC
  ffc_50
  (
    .doutp(ffc_50_p),
    .doutn(ffc_50_n),
    .din(ffc_111_p)
  );


  DROC
  ffc_51
  (
    .doutp(ffc_51_p),
    .doutn(ffc_51_n),
    .din(ffc_112_p)
  );


  DROC
  ffc_52
  (
    .doutp(ffc_52_p),
    .doutn(ffc_52_n),
    .din(ffc_114_p)
  );


  DROC
  ffc_53
  (
    .doutp(ffc_53_p),
    .doutn(ffc_53_n),
    .din(ffc_117_p)
  );


  DROC
  ffc_54
  (
    .doutp(ffc_54_p),
    .doutn(ffc_54_n),
    .din(ffc_134_p)
  );


  DROC
  ffc_55
  (
    .doutp(ffc_55_p),
    .doutn(ffc_55_n),
    .din(ffc_141_p)
  );


  DROC
  ffc_56
  (
    .doutp(ffc_56_p),
    .doutn(ffc_56_n),
    .din(ffc_144_p)
  );


  DROC
  ffc_57
  (
    .doutp(ffc_57_p),
    .doutn(ffc_57_n),
    .din(ffc_146_p)
  );


  DROC
  ffc_58
  (
    .doutp(ffc_58_p),
    .doutn(ffc_58_n),
    .din(ffc_154_p)
  );


  DROC
  ffc_59
  (
    .doutp(ffc_59_p),
    .doutn(ffc_59_n),
    .din(ffc_156_p)
  );


  DROC
  ffc_60
  (
    .doutp(ffc_60_p),
    .doutn(ffc_60_n),
    .din(ffc_157_p)
  );


  DROC
  ffc_61
  (
    .doutp(ffc_61_p),
    .doutn(ffc_61_n),
    .din(ffc_164_p)
  );


  DROC
  ffc_62
  (
    .doutp(ffc_62_p),
    .doutn(ffc_62_n),
    .din(ffc_170_p)
  );


  DROC
  ffc_63
  (
    .doutp(ffc_63_p),
    .doutn(ffc_63_n),
    .din(ffc_172_p)
  );


  DROC
  ffc_64
  (
    .doutp(ffc_64_p),
    .doutn(ffc_64_n),
    .din(ffc_118_p_spl_1)
  );


  DROC
  ffc_65
  (
    .doutp(ffc_65_p),
    .doutn(ffc_65_n),
    .din(ffc_119_p_spl_1)
  );


  DROC
  ffc_66
  (
    .doutp(ffc_66_p),
    .doutn(ffc_66_n),
    .din(ffc_120_p_spl_1)
  );


  DROC
  ffc_67
  (
    .doutp(ffc_67_p),
    .doutn(ffc_67_n),
    .din(ffc_121_p_spl_1)
  );


  DROC
  ffc_68
  (
    .doutp(ffc_68_p),
    .doutn(ffc_68_n),
    .din(ffc_122_p_spl_1)
  );


  DROC
  ffc_69
  (
    .doutp(ffc_69_p),
    .doutn(ffc_69_n),
    .din(ffc_123_p_spl_1)
  );


  DROC
  ffc_70
  (
    .doutp(ffc_70_p),
    .doutn(ffc_70_n),
    .din(ffc_124_p_spl_1)
  );


  DROC
  ffc_71
  (
    .doutp(ffc_71_p),
    .doutn(ffc_71_n),
    .din(ffc_125_p_spl_1)
  );


  DROC
  ffc_72
  (
    .doutp(ffc_72_p),
    .doutn(ffc_72_n),
    .din(ffc_126_p_spl_1)
  );


  DROC
  ffc_73
  (
    .doutp(ffc_73_p),
    .doutn(ffc_73_n),
    .din(ffc_127_p_spl_1)
  );


  DROC
  ffc_74
  (
    .doutp(ffc_74_p),
    .doutn(ffc_74_n),
    .din(ffc_128_p_spl_1)
  );


  DROC
  ffc_75
  (
    .doutp(ffc_75_p),
    .doutn(ffc_75_n),
    .din(ffc_129_p_spl_1)
  );


  DROC
  ffc_76
  (
    .doutp(ffc_76_p),
    .doutn(ffc_76_n),
    .din(ffc_130_p_spl_1)
  );


  DROC
  ffc_77
  (
    .doutp(ffc_77_p),
    .doutn(ffc_77_n),
    .din(ffc_131_p_spl_1)
  );


  DROC
  ffc_78
  (
    .doutp(ffc_78_p),
    .doutn(ffc_78_n),
    .din(ffc_132_p)
  );


  DROC
  ffc_79
  (
    .doutp(ffc_79_p),
    .doutn(ffc_79_n),
    .din(ffc_133_p_spl_1)
  );


  DROC
  ffc_80
  (
    .doutp(ffc_80_p),
    .doutn(ffc_80_n),
    .din(ffc_135_p_spl_1)
  );


  DROC
  ffc_81
  (
    .doutp(ffc_81_p),
    .doutn(ffc_81_n),
    .din(ffc_196_p)
  );


  DROC
  ffc_82
  (
    .doutp(ffc_82_p),
    .doutn(ffc_82_n),
    .din(ffc_205_p)
  );


  DROC
  ffc_83
  (
    .doutp(ffc_83_p),
    .doutn(ffc_83_n),
    .din(ffc_138_p)
  );


  DROC
  ffc_84
  (
    .doutp(ffc_84_p),
    .doutn(ffc_84_n),
    .din(ffc_139_p)
  );


  DROC
  ffc_85
  (
    .doutp(ffc_85_p),
    .doutn(ffc_85_n),
    .din(ffc_210_p)
  );


  DROC
  ffc_86
  (
    .doutp(ffc_86_p),
    .doutn(ffc_86_n),
    .din(ffc_140_p)
  );


  DROC
  ffc_87
  (
    .doutp(ffc_87_p),
    .doutn(ffc_87_n),
    .din(ffc_142_p)
  );


  DROC
  ffc_88
  (
    .doutp(ffc_88_p),
    .doutn(ffc_88_n),
    .din(ffc_145_p)
  );


  DROC
  ffc_89
  (
    .doutp(ffc_89_p),
    .doutn(ffc_89_n),
    .din(ffc_147_p)
  );


  DROC
  ffc_90
  (
    .doutp(ffc_90_p),
    .doutn(ffc_90_n),
    .din(ffc_229_p)
  );


  DROC
  ffc_91
  (
    .doutp(ffc_91_p),
    .doutn(ffc_91_n),
    .din(ffc_151_p)
  );


  DROC
  ffc_92
  (
    .doutp(ffc_92_p),
    .doutn(ffc_92_n),
    .din(ffc_254_p)
  );


  DROC
  ffc_93
  (
    .doutp(ffc_93_p),
    .doutn(ffc_93_n),
    .din(ffc_152_p)
  );


  DROC
  ffc_94
  (
    .doutp(ffc_94_p),
    .doutn(ffc_94_n),
    .din(ffc_153_p)
  );


  DROC
  ffc_95
  (
    .doutp(ffc_95_p),
    .doutn(ffc_95_n),
    .din(ffc_272_p_spl_)
  );


  DROC
  ffc_96
  (
    .doutp(ffc_96_p),
    .doutn(ffc_96_n),
    .din(ffc_158_p)
  );


  DROC
  ffc_97
  (
    .doutp(ffc_97_p),
    .doutn(ffc_97_n),
    .din(ffc_159_p)
  );


  DROC
  ffc_98
  (
    .doutp(ffc_98_p),
    .doutn(ffc_98_n),
    .din(ffc_163_p)
  );


  DROC
  ffc_99
  (
    .doutp(ffc_99_p),
    .doutn(ffc_99_n),
    .din(g574_p_spl_)
  );


  DROC
  ffc_100
  (
    .doutp(ffc_100_p),
    .doutn(ffc_100_n),
    .din(ffc_165_p)
  );


  DROC
  ffc_101
  (
    .doutp(ffc_101_p),
    .doutn(ffc_101_n),
    .din(g579_p_spl_)
  );


  DROC
  ffc_102
  (
    .doutp(ffc_102_p),
    .doutn(ffc_102_n),
    .din(ffc_171_p)
  );


  DROC
  ffc_103
  (
    .doutp(ffc_103_p),
    .doutn(ffc_103_n),
    .din(ffc_173_p)
  );


  DROC
  ffc_104
  (
    .doutp(ffc_104_p),
    .doutn(ffc_104_n),
    .din(g580_p_spl_)
  );


  DROC
  ffc_105
  (
    .doutp(ffc_105_p),
    .doutn(ffc_105_n),
    .din(ffc_177_p)
  );


  DROC
  ffc_106
  (
    .doutp(ffc_106_p),
    .doutn(ffc_106_n),
    .din(ffc_178_p)
  );


  DROC
  ffc_107
  (
    .doutp(ffc_107_p),
    .doutn(ffc_107_n),
    .din(ffc_179_p)
  );


  DROC
  ffc_108
  (
    .doutp(ffc_108_n),
    .doutn(ffc_108_p),
    .din(g581_n_spl_)
  );


  DROC
  ffc_109
  (
    .doutp(ffc_109_p),
    .doutn(ffc_109_n),
    .din(ffc_211_p)
  );


  DROC
  ffc_110
  (
    .doutp(ffc_110_p),
    .doutn(ffc_110_n),
    .din(g592_p_spl_)
  );


  DROC
  ffc_111
  (
    .doutp(ffc_111_p),
    .doutn(ffc_111_n),
    .din(ffc_213_p)
  );


  DROC
  ffc_112
  (
    .doutp(ffc_112_p),
    .doutn(ffc_112_n),
    .din(ffc_222_p)
  );


  DROC
  ffc_113
  (
    .doutp(ffc_113_p),
    .doutn(ffc_113_n),
    .din(g593_p_spl_)
  );


  DROC
  ffc_114
  (
    .doutp(ffc_114_p),
    .doutn(ffc_114_n),
    .din(ffc_230_p)
  );


  DROC
  ffc_115
  (
    .doutp(ffc_115_n),
    .doutn(ffc_115_p),
    .din(g594_n_spl_)
  );


  DROC
  ffc_116
  (
    .doutp(ffc_116_n),
    .doutn(ffc_116_p),
    .din(g609_p_spl_)
  );


  DROC
  ffc_117
  (
    .doutp(ffc_117_p),
    .doutn(ffc_117_n),
    .din(ffc_259_p)
  );


  DROC
  ffc_118
  (
    .doutp(ffc_118_p),
    .doutn(ffc_118_n),
    .din(ffc_180_p_spl_1)
  );


  DROC
  ffc_119
  (
    .doutp(ffc_119_p),
    .doutn(ffc_119_n),
    .din(ffc_181_p_spl_1)
  );


  DROC
  ffc_120
  (
    .doutp(ffc_120_p),
    .doutn(ffc_120_n),
    .din(ffc_182_p_spl_1)
  );


  DROC
  ffc_121
  (
    .doutp(ffc_121_p),
    .doutn(ffc_121_n),
    .din(ffc_183_p_spl_1)
  );


  DROC
  ffc_122
  (
    .doutp(ffc_122_p),
    .doutn(ffc_122_n),
    .din(ffc_184_p_spl_1)
  );


  DROC
  ffc_123
  (
    .doutp(ffc_123_p),
    .doutn(ffc_123_n),
    .din(ffc_185_p_spl_1)
  );


  DROC
  ffc_124
  (
    .doutp(ffc_124_p),
    .doutn(ffc_124_n),
    .din(ffc_186_p_spl_1)
  );


  DROC
  ffc_125
  (
    .doutp(ffc_125_p),
    .doutn(ffc_125_n),
    .din(ffc_187_p_spl_1)
  );


  DROC
  ffc_126
  (
    .doutp(ffc_126_p),
    .doutn(ffc_126_n),
    .din(ffc_188_p_spl_1)
  );


  DROC
  ffc_127
  (
    .doutp(ffc_127_p),
    .doutn(ffc_127_n),
    .din(ffc_189_p_spl_1)
  );


  DROC
  ffc_128
  (
    .doutp(ffc_128_p),
    .doutn(ffc_128_n),
    .din(ffc_190_p_spl_1)
  );


  DROC
  ffc_129
  (
    .doutp(ffc_129_p),
    .doutn(ffc_129_n),
    .din(ffc_191_p_spl_)
  );


  DROC
  ffc_130
  (
    .doutp(ffc_130_p),
    .doutn(ffc_130_n),
    .din(ffc_192_p_spl_1)
  );


  DROC
  ffc_131
  (
    .doutp(ffc_131_p),
    .doutn(ffc_131_n),
    .din(ffc_193_p_spl_)
  );


  DROC
  ffc_132
  (
    .doutp(ffc_132_p),
    .doutn(ffc_132_n),
    .din(ffc_194_p)
  );


  DROC
  ffc_133
  (
    .doutp(ffc_133_p),
    .doutn(ffc_133_n),
    .din(ffc_195_p_spl_1)
  );


  DROC
  ffc_134
  (
    .doutp(ffc_134_p),
    .doutn(ffc_134_n),
    .din(ffc_273_p)
  );


  DROC
  ffc_135
  (
    .doutp(ffc_135_p),
    .doutn(ffc_135_n),
    .din(ffc_207_p_spl_1)
  );


  DROC
  ffc_136
  (
    .doutp(ffc_136_n),
    .doutn(ffc_136_p),
    .din(g610_n_spl_)
  );


  DROC
  ffc_137
  (
    .doutp(ffc_137_p),
    .doutn(ffc_137_n),
    .din(g629_p_spl_)
  );


  DROC
  ffc_138
  (
    .doutp(ffc_138_p),
    .doutn(ffc_138_n),
    .din(ffc_208_p)
  );


  DROC
  ffc_139
  (
    .doutp(ffc_139_p),
    .doutn(ffc_139_n),
    .din(ffc_209_p)
  );


  DROC
  ffc_140
  (
    .doutp(ffc_140_p),
    .doutn(ffc_140_n),
    .din(ffc_212_p)
  );


  DROC
  ffc_141
  (
    .doutp(ffc_141_p),
    .doutn(ffc_141_n),
    .din(g630_p_spl_)
  );


  DROC
  ffc_142
  (
    .doutp(ffc_142_p),
    .doutn(ffc_142_n),
    .din(ffc_217_p)
  );


  DROC
  ffc_143
  (
    .doutp(ffc_143_p),
    .doutn(ffc_143_n),
    .din(g631_p_spl_)
  );


  DROC
  ffc_144
  (
    .doutp(ffc_144_p),
    .doutn(ffc_144_n),
    .din(g634_p_spl_)
  );


  DROC
  ffc_145
  (
    .doutp(ffc_145_p),
    .doutn(ffc_145_n),
    .din(ffc_223_p)
  );


  DROC
  ffc_146
  (
    .doutp(ffc_146_p),
    .doutn(ffc_146_n),
    .din(g635_p_spl_)
  );


  DROC
  ffc_147
  (
    .doutp(ffc_147_p),
    .doutn(ffc_147_n),
    .din(ffc_228_p)
  );


  DROC
  ffc_148
  (
    .doutp(ffc_148_p),
    .doutn(ffc_148_n),
    .din(ffc_15_p_spl_111)
  );


  DROC
  ffc_149
  (
    .doutp(ffc_149_n),
    .doutn(ffc_149_p),
    .din(g636_n_spl_)
  );


  DROC
  ffc_150
  (
    .doutp(ffc_150_p),
    .doutn(ffc_150_n),
    .din(g659_p_spl_)
  );


  DROC
  ffc_151
  (
    .doutp(ffc_151_p),
    .doutn(ffc_151_n),
    .din(ffc_231_p)
  );


  DROC
  ffc_152
  (
    .doutp(ffc_152_p),
    .doutn(ffc_152_n),
    .din(ffc_260_p)
  );


  DROC
  ffc_153
  (
    .doutp(ffc_153_p),
    .doutn(ffc_153_n),
    .din(ffc_274_p)
  );


  DROC
  ffc_154
  (
    .doutp(ffc_154_p),
    .doutn(ffc_154_n),
    .din(g660_p_spl_)
  );


  DROC
  ffc_155
  (
    .doutp(ffc_155_p),
    .doutn(ffc_155_n),
    .din(g661_p_spl_)
  );


  DROC
  ffc_156
  (
    .doutp(ffc_156_p),
    .doutn(ffc_156_n),
    .din(g670_p_spl_)
  );


  DROC
  ffc_157
  (
    .doutp(ffc_157_p),
    .doutn(ffc_157_n),
    .din(g671_p_spl_)
  );


  DROC
  ffc_158
  (
    .doutp(ffc_158_p),
    .doutn(ffc_158_n),
    .din(g672_p_spl_)
  );


  DROC
  ffc_159
  (
    .doutp(ffc_159_p),
    .doutn(ffc_159_n),
    .din(g673_p_spl_)
  );


  DROC
  ffc_160
  (
    .doutp(ffc_160_p),
    .doutn(ffc_160_n),
    .din(ffc_17_p_spl_11)
  );


  DROC
  ffc_161
  (
    .doutp(ffc_161_n),
    .doutn(ffc_161_p),
    .din(g674_n_spl_)
  );


  DROC
  ffc_162
  (
    .doutp(ffc_162_p),
    .doutn(ffc_162_n),
    .din(g701_p_spl_)
  );


  DROC
  ffc_163
  (
    .doutp(ffc_163_p),
    .doutn(ffc_163_n),
    .din(g702_p_spl_)
  );


  DROC
  ffc_164
  (
    .doutp(ffc_164_p),
    .doutn(ffc_164_n),
    .din(g703_p_spl_)
  );


  DROC
  ffc_165
  (
    .doutp(ffc_165_p),
    .doutn(ffc_165_n),
    .din(g704_p_spl_)
  );


  DROC
  ffc_166
  (
    .doutp(ffc_166_p),
    .doutn(ffc_166_n),
    .din(g739_n_spl_)
  );


  DROC
  ffc_167
  (
    .doutp(ffc_167_p),
    .doutn(ffc_167_n),
    .din(g789_n_spl_)
  );


  DROC
  ffc_168
  (
    .doutp(ffc_168_p),
    .doutn(ffc_168_n),
    .din(g839_n_spl_)
  );


  DROC
  ffc_169
  (
    .doutp(ffc_169_p),
    .doutn(ffc_169_n),
    .din(g840_p_spl_)
  );


  DROC
  ffc_170
  (
    .doutp(ffc_170_p),
    .doutn(ffc_170_n),
    .din(g857_p_spl_)
  );


  DROC
  ffc_171
  (
    .doutp(ffc_171_p),
    .doutn(ffc_171_n),
    .din(g864_p_spl_)
  );


  DROC
  ffc_172
  (
    .doutp(ffc_172_p),
    .doutn(ffc_172_n),
    .din(g865_p_spl_)
  );


  DROC
  ffc_173
  (
    .doutp(ffc_173_p),
    .doutn(ffc_173_n),
    .din(g866_p_spl_)
  );


  DROC
  ffc_174
  (
    .doutp(ffc_174_p),
    .doutn(ffc_174_n),
    .din(ffc_19_p_spl_11)
  );


  DROC
  ffc_175
  (
    .doutp(ffc_175_n),
    .doutn(ffc_175_p),
    .din(g867_n_spl_)
  );


  DROC
  ffc_176
  (
    .doutp(ffc_176_p),
    .doutn(ffc_176_n),
    .din(g889_p_spl_)
  );


  DROC
  ffc_177
  (
    .doutp(ffc_177_p),
    .doutn(ffc_177_n),
    .din(g890_p_spl_)
  );


  DROC
  ffc_178
  (
    .doutp(ffc_178_p),
    .doutn(ffc_178_n),
    .din(g905_p_spl_)
  );


  DROC
  ffc_179
  (
    .doutp(ffc_179_p),
    .doutn(ffc_179_n),
    .din(g906_p_spl_)
  );


  DROC
  ffc_180
  (
    .doutp(ffc_180_p),
    .doutn(ffc_180_n),
    .din(G3_p_spl_1)
  );


  DROC
  ffc_181
  (
    .doutp(ffc_181_p),
    .doutn(ffc_181_n),
    .din(G4_p_spl_1)
  );


  DROC
  ffc_182
  (
    .doutp(ffc_182_p),
    .doutn(ffc_182_n),
    .din(G5_p_spl_1)
  );


  DROC
  ffc_183
  (
    .doutp(ffc_183_p),
    .doutn(ffc_183_n),
    .din(G6_p_spl_1)
  );


  DROC
  ffc_184
  (
    .doutp(ffc_184_p),
    .doutn(ffc_184_n),
    .din(G7_p_spl_1)
  );


  DROC
  ffc_185
  (
    .doutp(ffc_185_p),
    .doutn(ffc_185_n),
    .din(G8_p_spl_1)
  );


  DROC
  ffc_186
  (
    .doutp(ffc_186_p),
    .doutn(ffc_186_n),
    .din(G9_p_spl_1)
  );


  DROC
  ffc_187
  (
    .doutp(ffc_187_p),
    .doutn(ffc_187_n),
    .din(G10_p_spl_1)
  );


  DROC
  ffc_188
  (
    .doutp(ffc_188_p),
    .doutn(ffc_188_n),
    .din(G11_p_spl_1)
  );


  DROC
  ffc_189
  (
    .doutp(ffc_189_p),
    .doutn(ffc_189_n),
    .din(G12_p_spl_1)
  );


  DROC
  ffc_190
  (
    .doutp(ffc_190_p),
    .doutn(ffc_190_n),
    .din(G13_p_spl_1)
  );


  DROC
  ffc_191
  (
    .doutp(ffc_191_p),
    .doutn(ffc_191_n),
    .din(G14_p_spl_1)
  );


  DROC
  ffc_192
  (
    .doutp(ffc_192_p),
    .doutn(ffc_192_n),
    .din(G15_p_spl_1)
  );


  DROC
  ffc_193
  (
    .doutp(ffc_193_p),
    .doutn(ffc_193_n),
    .din(G16_p_spl_1)
  );


  DROC
  ffc_194
  (
    .doutp(ffc_194_p),
    .doutn(ffc_194_n),
    .din(G17_p_spl_111)
  );


  DROC
  ffc_195
  (
    .doutp(ffc_195_p),
    .doutn(ffc_195_n),
    .din(G2_p_spl_1)
  );


  DROC
  ffc_196
  (
    .doutp(ffc_196_p),
    .doutn(ffc_196_n),
    .din(g907_p_spl_)
  );


  DROC
  ffc_197
  (
    .doutp(ffc_197_n),
    .doutn(ffc_197_p),
    .din(g911_n_spl_)
  );


  DROC
  ffc_198
  (
    .doutp(ffc_198_n),
    .doutn(ffc_198_p),
    .din(g915_n_spl_)
  );


  DROC
  ffc_199
  (
    .doutp(ffc_199_n),
    .doutn(ffc_199_p),
    .din(g919_n_spl_)
  );


  DROC
  ffc_200
  (
    .doutp(ffc_200_p),
    .doutn(ffc_200_n),
    .din(g922_n_spl_)
  );


  DROC
  ffc_201
  (
    .doutp(ffc_201_p),
    .doutn(ffc_201_n),
    .din(g934_n_spl_)
  );


  DROC
  ffc_202
  (
    .doutp(ffc_202_p),
    .doutn(ffc_202_n),
    .din(g946_n_spl_)
  );


  DROC
  ffc_203
  (
    .doutp(ffc_203_p),
    .doutn(ffc_203_n),
    .din(g958_n_spl_)
  );


  DROC
  ffc_204
  (
    .doutp(ffc_204_p),
    .doutn(ffc_204_n),
    .din(g959_p_spl_)
  );


  DROC
  ffc_205
  (
    .doutp(ffc_205_p),
    .doutn(ffc_205_n),
    .din(g984_p_spl_)
  );


  DROC
  ffc_206
  (
    .doutp(ffc_206_p),
    .doutn(ffc_206_n),
    .din(ffc_11_p_spl_11)
  );


  DROC
  ffc_207
  (
    .doutp(ffc_207_p),
    .doutn(ffc_207_n),
    .din(G1_p_spl_)
  );


  DROC
  ffc_208
  (
    .doutp(ffc_208_p),
    .doutn(ffc_208_n),
    .din(g985_p_spl_)
  );


  DROC
  ffc_209
  (
    .doutp(ffc_209_p),
    .doutn(ffc_209_n),
    .din(g986_p_spl_)
  );


  DROC
  ffc_210
  (
    .doutp(ffc_210_p),
    .doutn(ffc_210_n),
    .din(g987_p_spl_)
  );


  DROC
  ffc_211
  (
    .doutp(ffc_211_p),
    .doutn(ffc_211_n),
    .din(g988_p_spl_)
  );


  DROC
  ffc_212
  (
    .doutp(ffc_212_p),
    .doutn(ffc_212_n),
    .din(g989_p_spl_)
  );


  DROC
  ffc_213
  (
    .doutp(ffc_213_p),
    .doutn(ffc_213_n),
    .din(g1012_p_spl_)
  );


  DROC
  ffc_214
  (
    .doutp(ffc_214_p),
    .doutn(ffc_214_n),
    .din(ffc_21_p_spl_1)
  );


  DROC
  ffc_215
  (
    .doutp(ffc_215_n),
    .doutn(ffc_215_p),
    .din(g1013_n_spl_)
  );


  DROC
  ffc_216
  (
    .doutp(ffc_216_p),
    .doutn(ffc_216_n),
    .din(g1015_p_spl_)
  );


  DROC
  ffc_217
  (
    .doutp(ffc_217_p),
    .doutn(ffc_217_n),
    .din(g1016_p_spl_)
  );


  DROC
  ffc_218
  (
    .doutp(ffc_218_p),
    .doutn(ffc_218_n),
    .din(g1053_n_spl_)
  );


  DROC
  ffc_219
  (
    .doutp(ffc_219_p),
    .doutn(ffc_219_n),
    .din(g1107_n_spl_)
  );


  DROC
  ffc_220
  (
    .doutp(ffc_220_p),
    .doutn(ffc_220_n),
    .din(g1164_n_spl_)
  );


  DROC
  ffc_221
  (
    .doutp(ffc_221_p),
    .doutn(ffc_221_n),
    .din(g1241_n_spl_)
  );


  DROC
  ffc_222
  (
    .doutp(ffc_222_p),
    .doutn(ffc_222_n),
    .din(g1242_p_spl_)
  );


  DROC
  ffc_223
  (
    .doutp(ffc_223_p),
    .doutn(ffc_223_n),
    .din(g1250_p_spl_)
  );


  DROC
  ffc_224
  (
    .doutp(ffc_224_p),
    .doutn(ffc_224_n),
    .din(ffc_12_p_spl_11)
  );


  DROC
  ffc_225
  (
    .doutp(ffc_225_p),
    .doutn(ffc_225_n),
    .din(g1278_n_spl_)
  );


  DROC
  ffc_226
  (
    .doutp(ffc_226_p),
    .doutn(ffc_226_n),
    .din(g1328_n_spl_)
  );


  DROC
  ffc_227
  (
    .doutp(ffc_227_p),
    .doutn(ffc_227_n),
    .din(g1399_n_spl_)
  );


  DROC
  ffc_228
  (
    .doutp(ffc_228_p),
    .doutn(ffc_228_n),
    .din(g1400_p_spl_)
  );


  DROC
  ffc_229
  (
    .doutp(ffc_229_n),
    .doutn(ffc_229_p),
    .din(g1401_n_spl_)
  );


  DROC
  ffc_230
  (
    .doutp(ffc_230_n),
    .doutn(ffc_230_p),
    .din(g1402_n_spl_)
  );


  DROC
  ffc_231
  (
    .doutp(ffc_231_n),
    .doutn(ffc_231_p),
    .din(g1403_n_spl_)
  );


  DROC
  ffc_232
  (
    .doutp(ffc_232_p),
    .doutn(ffc_232_n),
    .din(g1407_p)
  );


  DROC
  ffc_233
  (
    .doutp(ffc_233_n),
    .doutn(ffc_233_p),
    .din(g1408_n)
  );


  DROC
  ffc_234
  (
    .doutp(ffc_234_p),
    .doutn(ffc_234_n),
    .din(g1412_p)
  );


  DROC
  ffc_235
  (
    .doutp(ffc_235_n),
    .doutn(ffc_235_p),
    .din(g1413_n)
  );


  DROC
  ffc_236
  (
    .doutp(ffc_236_p),
    .doutn(ffc_236_n),
    .din(g1417_p)
  );


  DROC
  ffc_237
  (
    .doutp(ffc_237_n),
    .doutn(ffc_237_p),
    .din(g1418_n)
  );


  DROC
  ffc_238
  (
    .doutp(ffc_238_n),
    .doutn(ffc_238_p),
    .din(g1422_p)
  );


  DROC
  ffc_239
  (
    .doutp(ffc_239_n),
    .doutn(ffc_239_p),
    .din(g1423_n)
  );


  DROC
  ffc_240
  (
    .doutp(ffc_240_n),
    .doutn(ffc_240_p),
    .din(g1427_p)
  );


  DROC
  ffc_241
  (
    .doutp(ffc_241_n),
    .doutn(ffc_241_p),
    .din(g1428_n)
  );


  DROC
  ffc_242
  (
    .doutp(ffc_242_n),
    .doutn(ffc_242_p),
    .din(g1432_p)
  );


  DROC
  ffc_243
  (
    .doutp(ffc_243_n),
    .doutn(ffc_243_p),
    .din(g1433_n)
  );


  DROC
  ffc_244
  (
    .doutp(ffc_244_p),
    .doutn(ffc_244_n),
    .din(g1434_p)
  );


  DROC
  ffc_245
  (
    .doutp(ffc_245_n),
    .doutn(ffc_245_p),
    .din(g1438_n_spl_)
  );


  DROC
  ffc_246
  (
    .doutp(ffc_246_n),
    .doutn(ffc_246_p),
    .din(g1442_n_spl_)
  );


  DROC
  ffc_247
  (
    .doutp(ffc_247_n),
    .doutn(ffc_247_p),
    .din(g1446_n_spl_)
  );


  DROC
  ffc_248
  (
    .doutp(ffc_248_n),
    .doutn(ffc_248_p),
    .din(g1450_n_spl_)
  );


  DROC
  ffc_249
  (
    .doutp(ffc_249_p),
    .doutn(ffc_249_n),
    .din(g1453_n_spl_)
  );


  DROC
  ffc_250
  (
    .doutp(ffc_250_p),
    .doutn(ffc_250_n),
    .din(g1477_p_spl_)
  );


  DROC
  ffc_251
  (
    .doutp(ffc_251_p),
    .doutn(ffc_251_n),
    .din(g1489_n_spl_)
  );


  DROC
  ffc_252
  (
    .doutp(ffc_252_p),
    .doutn(ffc_252_n),
    .din(g1501_n_spl_)
  );


  DROC
  ffc_253
  (
    .doutp(ffc_253_p),
    .doutn(ffc_253_n),
    .din(g1513_n_spl_)
  );


  DROC
  ffc_254
  (
    .doutp(ffc_254_p),
    .doutn(ffc_254_n),
    .din(g1515_p_spl_)
  );


  DROC
  ffc_255
  (
    .doutp(ffc_255_n),
    .doutn(ffc_255_p),
    .din(g1519_n_spl_)
  );


  DROC
  ffc_256
  (
    .doutp(ffc_256_n),
    .doutn(ffc_256_p),
    .din(g1523_n_spl_)
  );


  DROC
  ffc_257
  (
    .doutp(ffc_257_p),
    .doutn(ffc_257_n),
    .din(g1534_n_spl_)
  );


  DROC
  ffc_258
  (
    .doutp(ffc_258_p),
    .doutn(ffc_258_n),
    .din(g1546_n_spl_)
  );


  DROC
  ffc_259
  (
    .doutp(ffc_259_p),
    .doutn(ffc_259_n),
    .din(g1577_p_spl_)
  );


  DROC
  ffc_260
  (
    .doutp(ffc_260_p),
    .doutn(ffc_260_n),
    .din(g1593_p_spl_)
  );


  DROC
  ffc_261
  (
    .doutp(ffc_261_p),
    .doutn(ffc_261_n),
    .din(g1594_p)
  );


  DROC
  ffc_262
  (
    .doutp(ffc_262_p),
    .doutn(ffc_262_n),
    .din(g1595_p)
  );


  DROC
  ffc_263
  (
    .doutp(ffc_263_p),
    .doutn(ffc_263_n),
    .din(g1596_p)
  );


  DROC
  ffc_264
  (
    .doutp(ffc_264_p),
    .doutn(ffc_264_n),
    .din(g1597_p)
  );


  DROC
  ffc_265
  (
    .doutp(ffc_265_p),
    .doutn(ffc_265_n),
    .din(g1598_p)
  );


  DROC
  ffc_266
  (
    .doutp(ffc_266_p),
    .doutn(ffc_266_n),
    .din(g1599_p)
  );


  DROC
  ffc_267
  (
    .doutp(ffc_267_p),
    .doutn(ffc_267_n),
    .din(g1600_p)
  );


  DROC
  ffc_268
  (
    .doutp(ffc_268_p),
    .doutn(ffc_268_n),
    .din(g1617_p)
  );


  DROC
  ffc_269
  (
    .doutp(ffc_269_p),
    .doutn(ffc_269_n),
    .din(g1626_p)
  );


  DROC
  ffc_270
  (
    .doutp(ffc_270_n),
    .doutn(ffc_270_p),
    .din(g1627_n)
  );


  DROC
  ffc_271
  (
    .doutp(ffc_271_n),
    .doutn(ffc_271_p),
    .din(g1628_n)
  );


  DROC
  ffc_272
  (
    .doutp(ffc_272_p),
    .doutn(ffc_272_n),
    .din(g1629_p)
  );


  DROC
  ffc_273
  (
    .doutp(ffc_273_p),
    .doutn(ffc_273_n),
    .din(g1630_p_spl_)
  );


  DROC
  ffc_274
  (
    .doutp(ffc_274_p),
    .doutn(ffc_274_n),
    .din(g1631_p_spl_)
  );


  DROC
  ffc_275
  (
    .doutp(ffc_275_n),
    .doutn(ffc_275_p),
    .din(g1633_p)
  );


  DROC
  ffc_276
  (
    .doutp(ffc_276_n),
    .doutn(ffc_276_p),
    .din(g1635_p)
  );


  DROC
  ffc_277
  (
    .doutp(ffc_277_n),
    .doutn(ffc_277_p),
    .din(g1637_p)
  );


  DROC
  ffc_278
  (
    .doutp(ffc_278_n),
    .doutn(ffc_278_p),
    .din(g1639_p)
  );


  DROC
  ffc_279
  (
    .doutp(ffc_279_n),
    .doutn(ffc_279_p),
    .din(g1641_p)
  );


  DROC
  ffc_280
  (
    .doutp(ffc_280_n),
    .doutn(ffc_280_p),
    .din(g1643_p)
  );


  DROC
  ffc_281
  (
    .doutp(ffc_281_p),
    .doutn(ffc_281_n),
    .din(g1645_p)
  );


  DROC
  ffc_282
  (
    .doutp(ffc_282_p),
    .doutn(ffc_282_n),
    .din(g1647_p)
  );


  DROC
  ffc_283
  (
    .doutp(ffc_283_p),
    .doutn(ffc_283_n),
    .din(g1649_p)
  );


  DROC
  ffc_284
  (
    .doutp(ffc_284_p),
    .doutn(ffc_284_n),
    .din(g1651_p)
  );


  DROC
  ffc_285
  (
    .doutp(ffc_285_n),
    .doutn(ffc_285_p),
    .din(g1652_n)
  );


  DROC
  ffc_286
  (
    .doutp(ffc_286_n),
    .doutn(ffc_286_p),
    .din(g1687_p)
  );


  DROC
  ffc_287
  (
    .doutp(ffc_287_p),
    .doutn(ffc_287_n),
    .din(ffc_13_p)
  );


  DROC
  ffc_288
  (
    .doutp(ffc_288_p),
    .doutn(ffc_288_n),
    .din(g1691_p)
  );


  DROC
  ffc_289
  (
    .doutp(ffc_289_n),
    .doutn(ffc_289_p),
    .din(g1692_n)
  );


  DROC
  ffc_290
  (
    .doutp(ffc_290_p),
    .doutn(ffc_290_n),
    .din(g1696_p)
  );


  DROC
  ffc_291
  (
    .doutp(ffc_291_n),
    .doutn(ffc_291_p),
    .din(g1697_n)
  );


  DROC
  ffc_292
  (
    .doutp(ffc_292_n),
    .doutn(ffc_292_p),
    .din(g1700_p)
  );


  DROC
  ffc_293
  (
    .doutp(ffc_293_n),
    .doutn(ffc_293_p),
    .din(g1701_n)
  );


  DROC
  ffc_294
  (
    .doutp(ffc_294_n),
    .doutn(ffc_294_p),
    .din(g1705_p)
  );


  DROC
  ffc_295
  (
    .doutp(ffc_295_n),
    .doutn(ffc_295_p),
    .din(g1706_n)
  );


  DROC
  ffc_296
  (
    .doutp(ffc_296_n),
    .doutn(ffc_296_p),
    .din(g1776_p)
  );


  DROC
  ffc_297
  (
    .doutp(ffc_297_n),
    .doutn(ffc_297_p),
    .din(g1777_n)
  );


  DROC
  ffc_298
  (
    .doutp(ffc_298_n),
    .doutn(ffc_298_p),
    .din(g1814_p)
  );


  DROC
  ffc_299
  (
    .doutp(ffc_299_n),
    .doutn(ffc_299_p),
    .din(g1815_n)
  );


  DROC
  ffc_300
  (
    .doutp(ffc_300_n),
    .doutn(ffc_300_p),
    .din(g1851_p)
  );


  DROC
  ffc_301
  (
    .doutp(ffc_301_n),
    .doutn(ffc_301_p),
    .din(g1852_n)
  );


  DROC
  ffc_302
  (
    .doutp(ffc_302_n),
    .doutn(ffc_302_p),
    .din(g1880_p)
  );


  DROC
  ffc_303
  (
    .doutp(ffc_303_n),
    .doutn(ffc_303_p),
    .din(g1881_n)
  );


  DROC
  ffc_304
  (
    .doutp(ffc_304_n),
    .doutn(ffc_304_p),
    .din(g1901_p)
  );


  DROC
  ffc_305
  (
    .doutp(ffc_305_n),
    .doutn(ffc_305_p),
    .din(g1902_n)
  );


  DROC
  ffc_306
  (
    .doutp(ffc_306_n),
    .doutn(ffc_306_p),
    .din(g1914_p)
  );


  DROC
  ffc_307
  (
    .doutp(ffc_307_n),
    .doutn(ffc_307_p),
    .din(g1915_n)
  );


  DROC
  ffc_308
  (
    .doutp(ffc_308_n),
    .doutn(ffc_308_p),
    .din(g1919_p)
  );


  DROC
  ffc_309
  (
    .doutp(ffc_309_n),
    .doutn(ffc_309_p),
    .din(g1920_n)
  );


  DROC
  ffc_310
  (
    .doutp(ffc_310_p),
    .doutn(ffc_310_n),
    .din(g1924_n)
  );


  DROC
  ffc_311
  (
    .doutp(ffc_311_p),
    .doutn(ffc_311_n),
    .din(g1925_p)
  );


  DROC
  ffc_312
  (
    .doutp(ffc_312_p),
    .doutn(ffc_312_n),
    .din(g1975_n_spl_)
  );


  DROC
  ffc_313
  (
    .doutp(ffc_313_p),
    .doutn(ffc_313_n),
    .din(g1997_n_spl_)
  );


  DROC
  ffc_314
  (
    .doutp(ffc_314_p),
    .doutn(ffc_314_n),
    .din(g2019_n_spl_)
  );


  DROC
  ffc_315
  (
    .doutp(ffc_315_p),
    .doutn(ffc_315_n),
    .din(g2041_n_spl_)
  );


  DROC
  ffc_316
  (
    .doutp(ffc_316_p),
    .doutn(ffc_316_n),
    .din(g2063_n_spl_)
  );


  DROC
  ffc_317
  (
    .doutp(ffc_317_p),
    .doutn(ffc_317_n),
    .din(g2085_n_spl_)
  );


  DROC
  ffc_318
  (
    .doutp(ffc_318_p),
    .doutn(ffc_318_n),
    .din(g2107_n_spl_)
  );


  DROC
  ffc_319
  (
    .doutp(ffc_319_p),
    .doutn(ffc_319_n),
    .din(g2129_n_spl_)
  );


  DROC
  ffc_320
  (
    .doutp(ffc_320_p),
    .doutn(ffc_320_n),
    .din(g2151_n_spl_)
  );


  DROC
  ffc_321
  (
    .doutp(ffc_321_p),
    .doutn(ffc_321_n),
    .din(g2173_n_spl_)
  );


  DROC
  ffc_322
  (
    .doutp(ffc_322_p),
    .doutn(ffc_322_n),
    .din(g2189_n_spl_)
  );


  DROC
  ffc_323
  (
    .doutp(ffc_323_p),
    .doutn(ffc_323_n),
    .din(g2200_n_spl_)
  );


  DROC
  ffc_324
  (
    .doutp(ffc_324_p),
    .doutn(ffc_324_n),
    .din(g2212_n_spl_)
  );


  DROC
  ffc_325
  (
    .doutp(ffc_325_p),
    .doutn(ffc_325_n),
    .din(G21_p_spl_11)
  );


  DROC
  ffc_326
  (
    .doutp(ffc_326_p),
    .doutn(ffc_326_n),
    .din(g2213_p)
  );


  DROC
  ffc_327
  (
    .doutp(ffc_327_p),
    .doutn(ffc_327_n),
    .din(g2214_p)
  );


  DROC
  ffc_328
  (
    .doutp(ffc_328_p),
    .doutn(ffc_328_n),
    .din(g2215_p)
  );


  DROC
  ffc_329
  (
    .doutp(ffc_329_p),
    .doutn(ffc_329_n),
    .din(g2216_p)
  );


  DROC
  ffc_330
  (
    .doutp(ffc_330_p),
    .doutn(ffc_330_n),
    .din(g2217_p)
  );


  DROC
  ffc_331
  (
    .doutp(ffc_331_p),
    .doutn(ffc_331_n),
    .din(g2218_p)
  );


  DROC
  ffc_332
  (
    .doutp(ffc_332_p),
    .doutn(ffc_332_n),
    .din(g2219_p)
  );


  DROC
  ffc_333
  (
    .doutp(ffc_333_p),
    .doutn(ffc_333_n),
    .din(g2220_p)
  );


  DROC
  ffc_334
  (
    .doutp(ffc_334_p),
    .doutn(ffc_334_n),
    .din(g2221_p)
  );


  DROC
  ffc_335
  (
    .doutp(ffc_335_p),
    .doutn(ffc_335_n),
    .din(g2222_p)
  );


  DROC
  ffc_336
  (
    .doutp(ffc_336_p),
    .doutn(ffc_336_n),
    .din(g2223_p)
  );


  DROC
  ffc_337
  (
    .doutp(ffc_337_p),
    .doutn(ffc_337_n),
    .din(g2224_p)
  );


  DROC
  ffc_338
  (
    .doutp(ffc_338_p),
    .doutn(ffc_338_n),
    .din(g2225_p)
  );


  DROC
  ffc_339
  (
    .doutp(ffc_339_p),
    .doutn(ffc_339_n),
    .din(g2226_p)
  );


  DROC
  ffc_340
  (
    .doutp(ffc_340_p),
    .doutn(ffc_340_n),
    .din(g2227_p)
  );


  DROC
  ffc_341
  (
    .doutp(ffc_341_n),
    .doutn(ffc_341_p),
    .din(g2231_p)
  );


  DROC
  ffc_342
  (
    .doutp(ffc_342_n),
    .doutn(ffc_342_p),
    .din(g2232_n)
  );


  DROC
  ffc_343
  (
    .doutp(ffc_343_p),
    .doutn(ffc_343_n),
    .din(g2234_p)
  );


  DROC
  ffc_344
  (
    .doutp(ffc_344_p),
    .doutn(ffc_344_n),
    .din(g2236_p)
  );


  DROC
  ffc_345
  (
    .doutp(ffc_345_p),
    .doutn(ffc_345_n),
    .din(g2238_p)
  );


  DROC
  ffc_346
  (
    .doutp(ffc_346_p),
    .doutn(ffc_346_n),
    .din(g2240_p)
  );


  DROC
  ffc_347
  (
    .doutp(ffc_347_p),
    .doutn(ffc_347_n),
    .din(g2242_p)
  );


  DROC
  ffc_348
  (
    .doutp(ffc_348_p),
    .doutn(ffc_348_n),
    .din(g2244_p)
  );


  DROC
  ffc_349
  (
    .doutp(ffc_349_p),
    .doutn(ffc_349_n),
    .din(g2246_p)
  );


  DROC
  ffc_350
  (
    .doutp(ffc_350_p),
    .doutn(ffc_350_n),
    .din(g2248_p)
  );


  DROC
  ffc_351
  (
    .doutp(ffc_351_p),
    .doutn(ffc_351_n),
    .din(g2250_p)
  );


  DROC
  ffc_352
  (
    .doutp(ffc_352_p),
    .doutn(ffc_352_n),
    .din(g2252_p)
  );


  DROC
  ffc_353
  (
    .doutp(ffc_353_p),
    .doutn(ffc_353_n),
    .din(g2254_p)
  );


  DROC
  ffc_354
  (
    .doutp(ffc_354_p),
    .doutn(ffc_354_n),
    .din(g2256_p)
  );


  DROC
  ffc_355
  (
    .doutp(ffc_355_p),
    .doutn(ffc_355_n),
    .din(g2258_p)
  );


  buf

  (
    ffc_244_p_spl_,
    ffc_244_p
  );


  buf

  (
    ffc_242_p_spl_,
    ffc_242_p
  );


  buf

  (
    ffc_242_n_spl_,
    ffc_242_n
  );


  buf

  (
    g432_p_spl_,
    g432_p
  );


  buf

  (
    g433_n_spl_,
    g433_n
  );


  buf

  (
    g434_p_spl_,
    g434_p
  );


  buf

  (
    ffc_232_n_spl_,
    ffc_232_n
  );


  buf

  (
    ffc_232_p_spl_,
    ffc_232_p
  );


  buf

  (
    g438_n_spl_,
    g438_n
  );


  buf

  (
    g439_p_spl_,
    g439_p
  );


  buf

  (
    g438_p_spl_,
    g438_p
  );


  buf

  (
    g439_n_spl_,
    g439_n
  );


  buf

  (
    g440_n_spl_,
    g440_n
  );


  buf

  (
    g440_p_spl_,
    g440_p
  );


  buf

  (
    g437_p_spl_,
    g437_p
  );


  buf

  (
    g442_n_spl_,
    g442_n
  );


  buf

  (
    g443_p_spl_,
    g443_p
  );


  buf

  (
    ffc_30_p_spl_,
    ffc_30_p
  );


  buf

  (
    ffc_30_p_spl_0,
    ffc_30_p_spl_
  );


  buf

  (
    ffc_30_p_spl_00,
    ffc_30_p_spl_0
  );


  buf

  (
    ffc_30_p_spl_01,
    ffc_30_p_spl_0
  );


  buf

  (
    ffc_30_p_spl_1,
    ffc_30_p_spl_
  );


  buf

  (
    ffc_30_p_spl_10,
    ffc_30_p_spl_1
  );


  buf

  (
    ffc_30_n_spl_,
    ffc_30_n
  );


  buf

  (
    ffc_30_n_spl_0,
    ffc_30_n_spl_
  );


  buf

  (
    ffc_30_n_spl_00,
    ffc_30_n_spl_0
  );


  buf

  (
    ffc_30_n_spl_01,
    ffc_30_n_spl_0
  );


  buf

  (
    ffc_30_n_spl_1,
    ffc_30_n_spl_
  );


  buf

  (
    ffc_30_n_spl_10,
    ffc_30_n_spl_1
  );


  buf

  (
    ffc_240_p_spl_,
    ffc_240_p
  );


  buf

  (
    ffc_240_n_spl_,
    ffc_240_n
  );


  buf

  (
    g448_n_spl_,
    g448_n
  );


  buf

  (
    g449_p_spl_,
    g449_p
  );


  buf

  (
    g448_p_spl_,
    g448_p
  );


  buf

  (
    g449_n_spl_,
    g449_n
  );


  buf

  (
    g450_n_spl_,
    g450_n
  );


  buf

  (
    g450_p_spl_,
    g450_p
  );


  buf

  (
    g447_n_spl_,
    g447_n
  );


  buf

  (
    g452_p_spl_,
    g452_p
  );


  buf

  (
    g447_p_spl_,
    g447_p
  );


  buf

  (
    g452_n_spl_,
    g452_n
  );


  buf

  (
    g453_n_spl_,
    g453_n
  );


  buf

  (
    g453_p_spl_,
    g453_p
  );


  buf

  (
    g446_p_spl_,
    g446_p
  );


  buf

  (
    g455_n_spl_,
    g455_n
  );


  buf

  (
    g456_p_spl_,
    g456_p
  );


  buf

  (
    ffc_234_n_spl_,
    ffc_234_n
  );


  buf

  (
    ffc_234_p_spl_,
    ffc_234_p
  );


  buf

  (
    g462_n_spl_,
    g462_n
  );


  buf

  (
    g463_p_spl_,
    g463_p
  );


  buf

  (
    g462_p_spl_,
    g462_p
  );


  buf

  (
    g463_n_spl_,
    g463_n
  );


  buf

  (
    g464_n_spl_,
    g464_n
  );


  buf

  (
    g464_p_spl_,
    g464_p
  );


  buf

  (
    g461_n_spl_,
    g461_n
  );


  buf

  (
    g466_p_spl_,
    g466_p
  );


  buf

  (
    g461_p_spl_,
    g461_p
  );


  buf

  (
    g466_n_spl_,
    g466_n
  );


  buf

  (
    g467_n_spl_,
    g467_n
  );


  buf

  (
    g467_p_spl_,
    g467_p
  );


  buf

  (
    g460_n_spl_,
    g460_n
  );


  buf

  (
    g469_p_spl_,
    g469_p
  );


  buf

  (
    g460_p_spl_,
    g460_p
  );


  buf

  (
    g469_n_spl_,
    g469_n
  );


  buf

  (
    g470_n_spl_,
    g470_n
  );


  buf

  (
    g470_p_spl_,
    g470_p
  );


  buf

  (
    g459_p_spl_,
    g459_p
  );


  buf

  (
    g472_n_spl_,
    g472_n
  );


  buf

  (
    g473_p_spl_,
    g473_p
  );


  buf

  (
    ffc_4_p_spl_,
    ffc_4_p
  );


  buf

  (
    ffc_26_p_spl_,
    ffc_26_p
  );


  buf

  (
    ffc_26_p_spl_0,
    ffc_26_p_spl_
  );


  buf

  (
    ffc_26_p_spl_1,
    ffc_26_p_spl_
  );


  buf

  (
    ffc_4_n_spl_,
    ffc_4_n
  );


  buf

  (
    ffc_26_n_spl_,
    ffc_26_n
  );


  buf

  (
    ffc_26_n_spl_0,
    ffc_26_n_spl_
  );


  buf

  (
    ffc_26_n_spl_1,
    ffc_26_n_spl_
  );


  buf

  (
    ffc_238_p_spl_,
    ffc_238_p
  );


  buf

  (
    ffc_238_n_spl_,
    ffc_238_n
  );


  buf

  (
    g480_n_spl_,
    g480_n
  );


  buf

  (
    g481_p_spl_,
    g481_p
  );


  buf

  (
    g480_p_spl_,
    g480_p
  );


  buf

  (
    g481_n_spl_,
    g481_n
  );


  buf

  (
    g482_n_spl_,
    g482_n
  );


  buf

  (
    g482_p_spl_,
    g482_p
  );


  buf

  (
    g479_n_spl_,
    g479_n
  );


  buf

  (
    g484_p_spl_,
    g484_p
  );


  buf

  (
    g479_p_spl_,
    g479_p
  );


  buf

  (
    g484_n_spl_,
    g484_n
  );


  buf

  (
    g485_n_spl_,
    g485_n
  );


  buf

  (
    g485_p_spl_,
    g485_p
  );


  buf

  (
    g478_n_spl_,
    g478_n
  );


  buf

  (
    g487_p_spl_,
    g487_p
  );


  buf

  (
    g478_p_spl_,
    g478_p
  );


  buf

  (
    g487_n_spl_,
    g487_n
  );


  buf

  (
    g488_n_spl_,
    g488_n
  );


  buf

  (
    g488_p_spl_,
    g488_p
  );


  buf

  (
    g477_n_spl_,
    g477_n
  );


  buf

  (
    g490_p_spl_,
    g490_p
  );


  buf

  (
    g477_p_spl_,
    g477_p
  );


  buf

  (
    g490_n_spl_,
    g490_n
  );


  buf

  (
    g491_n_spl_,
    g491_n
  );


  buf

  (
    g491_p_spl_,
    g491_p
  );


  buf

  (
    g476_p_spl_,
    g476_p
  );


  buf

  (
    g493_n_spl_,
    g493_n
  );


  buf

  (
    g494_p_spl_,
    g494_p
  );


  buf

  (
    ffc_5_p_spl_,
    ffc_5_p
  );


  buf

  (
    ffc_5_n_spl_,
    ffc_5_n
  );


  buf

  (
    ffc_236_n_spl_,
    ffc_236_n
  );


  buf

  (
    ffc_236_p_spl_,
    ffc_236_p
  );


  buf

  (
    g502_n_spl_,
    g502_n
  );


  buf

  (
    g503_p_spl_,
    g503_p
  );


  buf

  (
    g502_p_spl_,
    g502_p
  );


  buf

  (
    g503_n_spl_,
    g503_n
  );


  buf

  (
    g504_n_spl_,
    g504_n
  );


  buf

  (
    g504_p_spl_,
    g504_p
  );


  buf

  (
    g501_n_spl_,
    g501_n
  );


  buf

  (
    g506_p_spl_,
    g506_p
  );


  buf

  (
    g501_p_spl_,
    g501_p
  );


  buf

  (
    g506_n_spl_,
    g506_n
  );


  buf

  (
    g507_n_spl_,
    g507_n
  );


  buf

  (
    g507_p_spl_,
    g507_p
  );


  buf

  (
    g500_n_spl_,
    g500_n
  );


  buf

  (
    g509_p_spl_,
    g509_p
  );


  buf

  (
    g500_p_spl_,
    g500_p
  );


  buf

  (
    g509_n_spl_,
    g509_n
  );


  buf

  (
    g510_n_spl_,
    g510_n
  );


  buf

  (
    g510_p_spl_,
    g510_p
  );


  buf

  (
    g499_n_spl_,
    g499_n
  );


  buf

  (
    g512_p_spl_,
    g512_p
  );


  buf

  (
    g499_p_spl_,
    g499_p
  );


  buf

  (
    g512_n_spl_,
    g512_n
  );


  buf

  (
    g513_n_spl_,
    g513_n
  );


  buf

  (
    g513_p_spl_,
    g513_p
  );


  buf

  (
    g498_n_spl_,
    g498_n
  );


  buf

  (
    g515_p_spl_,
    g515_p
  );


  buf

  (
    g498_p_spl_,
    g498_p
  );


  buf

  (
    g515_n_spl_,
    g515_n
  );


  buf

  (
    g516_n_spl_,
    g516_n
  );


  buf

  (
    g516_p_spl_,
    g516_p
  );


  buf

  (
    g497_p_spl_,
    g497_p
  );


  buf

  (
    g518_n_spl_,
    g518_n
  );


  buf

  (
    g519_p_spl_,
    g519_p
  );


  buf

  (
    ffc_6_p_spl_,
    ffc_6_p
  );


  buf

  (
    ffc_6_n_spl_,
    ffc_6_n
  );


  buf

  (
    ffc_7_p_spl_,
    ffc_7_p
  );


  buf

  (
    ffc_7_p_spl_0,
    ffc_7_p_spl_
  );


  buf

  (
    ffc_7_n_spl_,
    ffc_7_n
  );


  buf

  (
    ffc_7_n_spl_0,
    ffc_7_n_spl_
  );


  buf

  (
    g527_n_spl_,
    g527_n
  );


  buf

  (
    g528_n_spl_,
    g528_n
  );


  buf

  (
    g527_p_spl_,
    g527_p
  );


  buf

  (
    g528_p_spl_,
    g528_p
  );


  buf

  (
    g529_n_spl_,
    g529_n
  );


  buf

  (
    g529_p_spl_,
    g529_p
  );


  buf

  (
    g526_n_spl_,
    g526_n
  );


  buf

  (
    g531_p_spl_,
    g531_p
  );


  buf

  (
    g526_p_spl_,
    g526_p
  );


  buf

  (
    g531_n_spl_,
    g531_n
  );


  buf

  (
    g532_n_spl_,
    g532_n
  );


  buf

  (
    g532_p_spl_,
    g532_p
  );


  buf

  (
    g525_n_spl_,
    g525_n
  );


  buf

  (
    g534_p_spl_,
    g534_p
  );


  buf

  (
    g525_p_spl_,
    g525_p
  );


  buf

  (
    g534_n_spl_,
    g534_n
  );


  buf

  (
    g535_n_spl_,
    g535_n
  );


  buf

  (
    g535_p_spl_,
    g535_p
  );


  buf

  (
    g524_n_spl_,
    g524_n
  );


  buf

  (
    g537_p_spl_,
    g537_p
  );


  buf

  (
    g524_p_spl_,
    g524_p
  );


  buf

  (
    g537_n_spl_,
    g537_n
  );


  buf

  (
    g538_n_spl_,
    g538_n
  );


  buf

  (
    g538_p_spl_,
    g538_p
  );


  buf

  (
    g523_n_spl_,
    g523_n
  );


  buf

  (
    g540_p_spl_,
    g540_p
  );


  buf

  (
    g523_p_spl_,
    g523_p
  );


  buf

  (
    g540_n_spl_,
    g540_n
  );


  buf

  (
    g541_n_spl_,
    g541_n
  );


  buf

  (
    g541_p_spl_,
    g541_p
  );


  buf

  (
    g522_p_spl_,
    g522_p
  );


  buf

  (
    g543_n_spl_,
    g543_n
  );


  buf

  (
    g544_p_spl_,
    g544_p
  );


  buf

  (
    g550_n_spl_,
    g550_n
  );


  buf

  (
    g551_n_spl_,
    g551_n
  );


  buf

  (
    g550_p_spl_,
    g550_p
  );


  buf

  (
    g551_p_spl_,
    g551_p
  );


  buf

  (
    g552_n_spl_,
    g552_n
  );


  buf

  (
    g552_p_spl_,
    g552_p
  );


  buf

  (
    g549_n_spl_,
    g549_n
  );


  buf

  (
    g554_p_spl_,
    g554_p
  );


  buf

  (
    g549_p_spl_,
    g549_p
  );


  buf

  (
    g554_n_spl_,
    g554_n
  );


  buf

  (
    g555_n_spl_,
    g555_n
  );


  buf

  (
    g555_p_spl_,
    g555_p
  );


  buf

  (
    g548_n_spl_,
    g548_n
  );


  buf

  (
    g557_p_spl_,
    g557_p
  );


  buf

  (
    g548_p_spl_,
    g548_p
  );


  buf

  (
    g557_n_spl_,
    g557_n
  );


  buf

  (
    g558_n_spl_,
    g558_n
  );


  buf

  (
    g558_p_spl_,
    g558_p
  );


  buf

  (
    g547_p_spl_,
    g547_p
  );


  buf

  (
    g560_n_spl_,
    g560_n
  );


  buf

  (
    g561_p_spl_,
    g561_p
  );


  buf

  (
    g564_n_spl_,
    g564_n
  );


  buf

  (
    g565_n_spl_,
    g565_n
  );


  buf

  (
    g564_p_spl_,
    g564_p
  );


  buf

  (
    g565_p_spl_,
    g565_p
  );


  buf

  (
    g566_n_spl_,
    g566_n
  );


  buf

  (
    g570_n_spl_,
    g570_n
  );


  buf

  (
    ffc_25_p_spl_,
    ffc_25_p
  );


  buf

  (
    ffc_25_p_spl_0,
    ffc_25_p_spl_
  );


  buf

  (
    ffc_25_p_spl_00,
    ffc_25_p_spl_0
  );


  buf

  (
    ffc_25_p_spl_000,
    ffc_25_p_spl_00
  );


  buf

  (
    ffc_25_p_spl_001,
    ffc_25_p_spl_00
  );


  buf

  (
    ffc_25_p_spl_01,
    ffc_25_p_spl_0
  );


  buf

  (
    ffc_25_p_spl_010,
    ffc_25_p_spl_01
  );


  buf

  (
    ffc_25_p_spl_011,
    ffc_25_p_spl_01
  );


  buf

  (
    ffc_25_p_spl_1,
    ffc_25_p_spl_
  );


  buf

  (
    ffc_25_p_spl_10,
    ffc_25_p_spl_1
  );


  buf

  (
    ffc_25_p_spl_11,
    ffc_25_p_spl_1
  );


  buf

  (
    ffc_80_p_spl_,
    ffc_80_p
  );


  buf

  (
    ffc_25_n_spl_,
    ffc_25_n
  );


  buf

  (
    ffc_25_n_spl_0,
    ffc_25_n_spl_
  );


  buf

  (
    ffc_25_n_spl_00,
    ffc_25_n_spl_0
  );


  buf

  (
    ffc_25_n_spl_000,
    ffc_25_n_spl_00
  );


  buf

  (
    ffc_25_n_spl_001,
    ffc_25_n_spl_00
  );


  buf

  (
    ffc_25_n_spl_01,
    ffc_25_n_spl_0
  );


  buf

  (
    ffc_25_n_spl_010,
    ffc_25_n_spl_01
  );


  buf

  (
    ffc_25_n_spl_011,
    ffc_25_n_spl_01
  );


  buf

  (
    ffc_25_n_spl_1,
    ffc_25_n_spl_
  );


  buf

  (
    ffc_25_n_spl_10,
    ffc_25_n_spl_1
  );


  buf

  (
    ffc_25_n_spl_11,
    ffc_25_n_spl_1
  );


  buf

  (
    ffc_80_n_spl_,
    ffc_80_n
  );


  buf

  (
    ffc_272_p_spl_,
    ffc_272_p
  );


  buf

  (
    g575_n_spl_,
    g575_n
  );


  buf

  (
    g576_p_spl_,
    g576_p
  );


  buf

  (
    g575_p_spl_,
    g575_p
  );


  buf

  (
    g576_n_spl_,
    g576_n
  );


  buf

  (
    g577_n_spl_,
    g577_n
  );


  buf

  (
    g577_p_spl_,
    g577_p
  );


  buf

  (
    g579_p_spl_,
    g579_p
  );


  buf

  (
    g574_p_spl_,
    g574_p
  );


  buf

  (
    ffc_29_n_spl_,
    ffc_29_n
  );


  buf

  (
    ffc_29_n_spl_0,
    ffc_29_n_spl_
  );


  buf

  (
    ffc_29_n_spl_00,
    ffc_29_n_spl_0
  );


  buf

  (
    ffc_29_n_spl_000,
    ffc_29_n_spl_00
  );


  buf

  (
    ffc_29_n_spl_01,
    ffc_29_n_spl_0
  );


  buf

  (
    ffc_29_n_spl_1,
    ffc_29_n_spl_
  );


  buf

  (
    ffc_29_n_spl_10,
    ffc_29_n_spl_1
  );


  buf

  (
    ffc_29_n_spl_11,
    ffc_29_n_spl_1
  );


  buf

  (
    g580_p_spl_,
    g580_p
  );


  buf

  (
    ffc_79_p_spl_,
    ffc_79_p
  );


  buf

  (
    ffc_79_n_spl_,
    ffc_79_n
  );


  buf

  (
    ffc_270_n_spl_,
    ffc_270_n
  );


  buf

  (
    ffc_275_n_spl_,
    ffc_275_n
  );


  buf

  (
    ffc_270_p_spl_,
    ffc_270_p
  );


  buf

  (
    ffc_275_p_spl_,
    ffc_275_p
  );


  buf

  (
    g584_n_spl_,
    g584_n
  );


  buf

  (
    g584_p_spl_,
    g584_p
  );


  buf

  (
    g583_n_spl_,
    g583_n
  );


  buf

  (
    g586_p_spl_,
    g586_p
  );


  buf

  (
    g583_p_spl_,
    g583_p
  );


  buf

  (
    g586_n_spl_,
    g586_n
  );


  buf

  (
    g587_n_spl_,
    g587_n
  );


  buf

  (
    g587_p_spl_,
    g587_p
  );


  buf

  (
    g582_n_spl_,
    g582_n
  );


  buf

  (
    g589_p_spl_,
    g589_p
  );


  buf

  (
    g581_n_spl_,
    g581_n
  );


  buf

  (
    g592_p_spl_,
    g592_p
  );


  buf

  (
    g593_p_spl_,
    g593_p
  );


  buf

  (
    ffc_29_p_spl_,
    ffc_29_p
  );


  buf

  (
    ffc_29_p_spl_0,
    ffc_29_p_spl_
  );


  buf

  (
    ffc_29_p_spl_00,
    ffc_29_p_spl_0
  );


  buf

  (
    ffc_29_p_spl_01,
    ffc_29_p_spl_0
  );


  buf

  (
    ffc_29_p_spl_1,
    ffc_29_p_spl_
  );


  buf

  (
    ffc_29_p_spl_10,
    ffc_29_p_spl_1
  );


  buf

  (
    ffc_29_p_spl_11,
    ffc_29_p_spl_1
  );


  buf

  (
    ffc_64_p_spl_,
    ffc_64_p
  );


  buf

  (
    ffc_64_n_spl_,
    ffc_64_n
  );


  buf

  (
    ffc_268_n_spl_,
    ffc_268_n
  );


  buf

  (
    ffc_276_n_spl_,
    ffc_276_n
  );


  buf

  (
    ffc_268_p_spl_,
    ffc_268_p
  );


  buf

  (
    ffc_276_p_spl_,
    ffc_276_p
  );


  buf

  (
    g598_n_spl_,
    g598_n
  );


  buf

  (
    g598_p_spl_,
    g598_p
  );


  buf

  (
    g597_n_spl_,
    g597_n
  );


  buf

  (
    g600_p_spl_,
    g600_p
  );


  buf

  (
    g597_p_spl_,
    g597_p
  );


  buf

  (
    g600_n_spl_,
    g600_n
  );


  buf

  (
    g601_n_spl_,
    g601_n
  );


  buf

  (
    g601_p_spl_,
    g601_p
  );


  buf

  (
    g596_n_spl_,
    g596_n
  );


  buf

  (
    g603_p_spl_,
    g603_p
  );


  buf

  (
    g596_p_spl_,
    g596_p
  );


  buf

  (
    g603_n_spl_,
    g603_n
  );


  buf

  (
    g604_n_spl_,
    g604_n
  );


  buf

  (
    g604_p_spl_,
    g604_p
  );


  buf

  (
    g595_n_spl_,
    g595_n
  );


  buf

  (
    g606_p_spl_,
    g606_p
  );


  buf

  (
    g607_n_spl_,
    g607_n
  );


  buf

  (
    g594_n_spl_,
    g594_n
  );


  buf

  (
    g609_p_spl_,
    g609_p
  );


  buf

  (
    ffc_65_p_spl_,
    ffc_65_p
  );


  buf

  (
    ffc_65_n_spl_,
    ffc_65_n
  );


  buf

  (
    ffc_269_n_spl_,
    ffc_269_n
  );


  buf

  (
    ffc_277_n_spl_,
    ffc_277_n
  );


  buf

  (
    ffc_269_p_spl_,
    ffc_269_p
  );


  buf

  (
    ffc_277_p_spl_,
    ffc_277_p
  );


  buf

  (
    g615_n_spl_,
    g615_n
  );


  buf

  (
    g615_p_spl_,
    g615_p
  );


  buf

  (
    g614_n_spl_,
    g614_n
  );


  buf

  (
    g617_p_spl_,
    g617_p
  );


  buf

  (
    g614_p_spl_,
    g614_p
  );


  buf

  (
    g617_n_spl_,
    g617_n
  );


  buf

  (
    g618_n_spl_,
    g618_n
  );


  buf

  (
    g618_p_spl_,
    g618_p
  );


  buf

  (
    g613_n_spl_,
    g613_n
  );


  buf

  (
    g620_p_spl_,
    g620_p
  );


  buf

  (
    g613_p_spl_,
    g613_p
  );


  buf

  (
    g620_n_spl_,
    g620_n
  );


  buf

  (
    g621_n_spl_,
    g621_n
  );


  buf

  (
    g621_p_spl_,
    g621_p
  );


  buf

  (
    g612_n_spl_,
    g612_n
  );


  buf

  (
    g623_p_spl_,
    g623_p
  );


  buf

  (
    g612_p_spl_,
    g612_p
  );


  buf

  (
    g623_n_spl_,
    g623_n
  );


  buf

  (
    g624_n_spl_,
    g624_n
  );


  buf

  (
    g624_p_spl_,
    g624_p
  );


  buf

  (
    g611_n_spl_,
    g611_n
  );


  buf

  (
    g626_p_spl_,
    g626_p
  );


  buf

  (
    ffc_135_p_spl_,
    ffc_135_p
  );


  buf

  (
    ffc_135_p_spl_0,
    ffc_135_p_spl_
  );


  buf

  (
    ffc_135_p_spl_00,
    ffc_135_p_spl_0
  );


  buf

  (
    ffc_135_p_spl_1,
    ffc_135_p_spl_
  );


  buf

  (
    ffc_287_p_spl_,
    ffc_287_p
  );


  buf

  (
    ffc_287_p_spl_0,
    ffc_287_p_spl_
  );


  buf

  (
    ffc_287_p_spl_00,
    ffc_287_p_spl_0
  );


  buf

  (
    ffc_287_p_spl_000,
    ffc_287_p_spl_00
  );


  buf

  (
    ffc_287_p_spl_001,
    ffc_287_p_spl_00
  );


  buf

  (
    ffc_287_p_spl_01,
    ffc_287_p_spl_0
  );


  buf

  (
    ffc_287_p_spl_010,
    ffc_287_p_spl_01
  );


  buf

  (
    ffc_287_p_spl_011,
    ffc_287_p_spl_01
  );


  buf

  (
    ffc_287_p_spl_1,
    ffc_287_p_spl_
  );


  buf

  (
    ffc_287_p_spl_10,
    ffc_287_p_spl_1
  );


  buf

  (
    ffc_287_p_spl_100,
    ffc_287_p_spl_10
  );


  buf

  (
    ffc_287_p_spl_101,
    ffc_287_p_spl_10
  );


  buf

  (
    ffc_287_p_spl_11,
    ffc_287_p_spl_1
  );


  buf

  (
    ffc_287_p_spl_110,
    ffc_287_p_spl_11
  );


  buf

  (
    ffc_287_p_spl_111,
    ffc_287_p_spl_11
  );


  buf

  (
    ffc_135_n_spl_,
    ffc_135_n
  );


  buf

  (
    ffc_135_n_spl_0,
    ffc_135_n_spl_
  );


  buf

  (
    ffc_135_n_spl_00,
    ffc_135_n_spl_0
  );


  buf

  (
    ffc_135_n_spl_1,
    ffc_135_n_spl_
  );


  buf

  (
    ffc_287_n_spl_,
    ffc_287_n
  );


  buf

  (
    ffc_287_n_spl_0,
    ffc_287_n_spl_
  );


  buf

  (
    ffc_287_n_spl_00,
    ffc_287_n_spl_0
  );


  buf

  (
    ffc_287_n_spl_000,
    ffc_287_n_spl_00
  );


  buf

  (
    ffc_287_n_spl_001,
    ffc_287_n_spl_00
  );


  buf

  (
    ffc_287_n_spl_01,
    ffc_287_n_spl_0
  );


  buf

  (
    ffc_287_n_spl_010,
    ffc_287_n_spl_01
  );


  buf

  (
    ffc_287_n_spl_011,
    ffc_287_n_spl_01
  );


  buf

  (
    ffc_287_n_spl_1,
    ffc_287_n_spl_
  );


  buf

  (
    ffc_287_n_spl_10,
    ffc_287_n_spl_1
  );


  buf

  (
    ffc_287_n_spl_100,
    ffc_287_n_spl_10
  );


  buf

  (
    ffc_287_n_spl_101,
    ffc_287_n_spl_10
  );


  buf

  (
    ffc_287_n_spl_11,
    ffc_287_n_spl_1
  );


  buf

  (
    ffc_287_n_spl_110,
    ffc_287_n_spl_11
  );


  buf

  (
    ffc_287_n_spl_111,
    ffc_287_n_spl_11
  );


  buf

  (
    g610_n_spl_,
    g610_n
  );


  buf

  (
    g629_p_spl_,
    g629_p
  );


  buf

  (
    ffc_285_n_spl_,
    ffc_285_n
  );


  buf

  (
    ffc_286_n_spl_,
    ffc_286_n
  );


  buf

  (
    ffc_285_p_spl_,
    ffc_285_p
  );


  buf

  (
    ffc_286_p_spl_,
    ffc_286_p
  );


  buf

  (
    g632_n_spl_,
    g632_n
  );


  buf

  (
    g632_p_spl_,
    g632_p
  );


  buf

  (
    g634_p_spl_,
    g634_p
  );


  buf

  (
    g630_p_spl_,
    g630_p
  );


  buf

  (
    g631_p_spl_,
    g631_p
  );


  buf

  (
    ffc_66_p_spl_,
    ffc_66_p
  );


  buf

  (
    ffc_66_n_spl_,
    ffc_66_n
  );


  buf

  (
    ffc_261_n_spl_,
    ffc_261_n
  );


  buf

  (
    ffc_284_p_spl_,
    ffc_284_p
  );


  buf

  (
    ffc_261_p_spl_,
    ffc_261_p
  );


  buf

  (
    ffc_284_n_spl_,
    ffc_284_n
  );


  buf

  (
    g642_n_spl_,
    g642_n
  );


  buf

  (
    g642_p_spl_,
    g642_p
  );


  buf

  (
    g641_n_spl_,
    g641_n
  );


  buf

  (
    g644_p_spl_,
    g644_p
  );


  buf

  (
    g641_p_spl_,
    g641_p
  );


  buf

  (
    g644_n_spl_,
    g644_n
  );


  buf

  (
    g645_n_spl_,
    g645_n
  );


  buf

  (
    g645_p_spl_,
    g645_p
  );


  buf

  (
    g640_n_spl_,
    g640_n
  );


  buf

  (
    g647_p_spl_,
    g647_p
  );


  buf

  (
    g640_p_spl_,
    g640_p
  );


  buf

  (
    g647_n_spl_,
    g647_n
  );


  buf

  (
    g648_n_spl_,
    g648_n
  );


  buf

  (
    g648_p_spl_,
    g648_p
  );


  buf

  (
    g639_n_spl_,
    g639_n
  );


  buf

  (
    g650_p_spl_,
    g650_p
  );


  buf

  (
    g639_p_spl_,
    g639_p
  );


  buf

  (
    g650_n_spl_,
    g650_n
  );


  buf

  (
    g651_n_spl_,
    g651_n
  );


  buf

  (
    g651_p_spl_,
    g651_p
  );


  buf

  (
    g638_n_spl_,
    g638_n
  );


  buf

  (
    g653_p_spl_,
    g653_p
  );


  buf

  (
    g638_p_spl_,
    g638_p
  );


  buf

  (
    g653_n_spl_,
    g653_n
  );


  buf

  (
    g654_n_spl_,
    g654_n
  );


  buf

  (
    g654_p_spl_,
    g654_p
  );


  buf

  (
    g637_n_spl_,
    g637_n
  );


  buf

  (
    g656_p_spl_,
    g656_p
  );


  buf

  (
    ffc_15_p_spl_,
    ffc_15_p
  );


  buf

  (
    ffc_15_p_spl_0,
    ffc_15_p_spl_
  );


  buf

  (
    ffc_15_p_spl_00,
    ffc_15_p_spl_0
  );


  buf

  (
    ffc_15_p_spl_000,
    ffc_15_p_spl_00
  );


  buf

  (
    ffc_15_p_spl_001,
    ffc_15_p_spl_00
  );


  buf

  (
    ffc_15_p_spl_01,
    ffc_15_p_spl_0
  );


  buf

  (
    ffc_15_p_spl_010,
    ffc_15_p_spl_01
  );


  buf

  (
    ffc_15_p_spl_011,
    ffc_15_p_spl_01
  );


  buf

  (
    ffc_15_p_spl_1,
    ffc_15_p_spl_
  );


  buf

  (
    ffc_15_p_spl_10,
    ffc_15_p_spl_1
  );


  buf

  (
    ffc_15_p_spl_100,
    ffc_15_p_spl_10
  );


  buf

  (
    ffc_15_p_spl_101,
    ffc_15_p_spl_10
  );


  buf

  (
    ffc_15_p_spl_11,
    ffc_15_p_spl_1
  );


  buf

  (
    ffc_15_p_spl_110,
    ffc_15_p_spl_11
  );


  buf

  (
    ffc_15_p_spl_111,
    ffc_15_p_spl_11
  );


  buf

  (
    ffc_15_n_spl_,
    ffc_15_n
  );


  buf

  (
    ffc_15_n_spl_0,
    ffc_15_n_spl_
  );


  buf

  (
    ffc_15_n_spl_00,
    ffc_15_n_spl_0
  );


  buf

  (
    ffc_15_n_spl_000,
    ffc_15_n_spl_00
  );


  buf

  (
    ffc_15_n_spl_001,
    ffc_15_n_spl_00
  );


  buf

  (
    ffc_15_n_spl_01,
    ffc_15_n_spl_0
  );


  buf

  (
    ffc_15_n_spl_010,
    ffc_15_n_spl_01
  );


  buf

  (
    ffc_15_n_spl_011,
    ffc_15_n_spl_01
  );


  buf

  (
    ffc_15_n_spl_1,
    ffc_15_n_spl_
  );


  buf

  (
    ffc_15_n_spl_10,
    ffc_15_n_spl_1
  );


  buf

  (
    ffc_15_n_spl_100,
    ffc_15_n_spl_10
  );


  buf

  (
    ffc_15_n_spl_101,
    ffc_15_n_spl_10
  );


  buf

  (
    ffc_15_n_spl_11,
    ffc_15_n_spl_1
  );


  buf

  (
    g636_n_spl_,
    g636_n
  );


  buf

  (
    g659_p_spl_,
    g659_p
  );


  buf

  (
    g635_p_spl_,
    g635_p
  );


  buf

  (
    ffc_133_p_spl_,
    ffc_133_p
  );


  buf

  (
    ffc_133_p_spl_0,
    ffc_133_p_spl_
  );


  buf

  (
    ffc_133_p_spl_00,
    ffc_133_p_spl_0
  );


  buf

  (
    ffc_133_p_spl_1,
    ffc_133_p_spl_
  );


  buf

  (
    ffc_133_n_spl_,
    ffc_133_n
  );


  buf

  (
    ffc_133_n_spl_0,
    ffc_133_n_spl_
  );


  buf

  (
    ffc_133_n_spl_00,
    ffc_133_n_spl_0
  );


  buf

  (
    ffc_133_n_spl_1,
    ffc_133_n_spl_
  );


  buf

  (
    ffc_310_p_spl_,
    ffc_310_p
  );


  buf

  (
    ffc_310_n_spl_,
    ffc_310_n
  );


  buf

  (
    g663_n_spl_,
    g663_n
  );


  buf

  (
    g664_p_spl_,
    g664_p
  );


  buf

  (
    g663_p_spl_,
    g663_p
  );


  buf

  (
    g664_n_spl_,
    g664_n
  );


  buf

  (
    g665_n_spl_,
    g665_n
  );


  buf

  (
    g665_p_spl_,
    g665_p
  );


  buf

  (
    g662_n_spl_,
    g662_n
  );


  buf

  (
    g667_p_spl_,
    g667_p
  );


  buf

  (
    g662_p_spl_,
    g662_p
  );


  buf

  (
    g667_n_spl_,
    g667_n
  );


  buf

  (
    g668_n_spl_,
    g668_n
  );


  buf

  (
    g668_p_spl_,
    g668_p
  );


  buf

  (
    g670_p_spl_,
    g670_p
  );


  buf

  (
    g660_p_spl_,
    g660_p
  );


  buf

  (
    ffc_207_p_spl_,
    ffc_207_p
  );


  buf

  (
    ffc_207_p_spl_0,
    ffc_207_p_spl_
  );


  buf

  (
    ffc_207_p_spl_00,
    ffc_207_p_spl_0
  );


  buf

  (
    ffc_207_p_spl_1,
    ffc_207_p_spl_
  );


  buf

  (
    ffc_325_p_spl_,
    ffc_325_p
  );


  buf

  (
    ffc_325_p_spl_0,
    ffc_325_p_spl_
  );


  buf

  (
    ffc_207_n_spl_,
    ffc_207_n
  );


  buf

  (
    ffc_207_n_spl_0,
    ffc_207_n_spl_
  );


  buf

  (
    ffc_207_n_spl_00,
    ffc_207_n_spl_0
  );


  buf

  (
    ffc_207_n_spl_1,
    ffc_207_n_spl_
  );


  buf

  (
    ffc_325_n_spl_,
    ffc_325_n
  );


  buf

  (
    ffc_325_n_spl_0,
    ffc_325_n_spl_
  );


  buf

  (
    ffc_341_p_spl_,
    ffc_341_p
  );


  buf

  (
    ffc_341_n_spl_,
    ffc_341_n
  );


  buf

  (
    g661_p_spl_,
    g661_p
  );


  buf

  (
    ffc_67_p_spl_,
    ffc_67_p
  );


  buf

  (
    ffc_67_n_spl_,
    ffc_67_n
  );


  buf

  (
    ffc_68_p_spl_,
    ffc_68_p
  );


  buf

  (
    ffc_68_p_spl_0,
    ffc_68_p_spl_
  );


  buf

  (
    ffc_214_p_spl_,
    ffc_214_p
  );


  buf

  (
    ffc_214_p_spl_0,
    ffc_214_p_spl_
  );


  buf

  (
    ffc_214_p_spl_00,
    ffc_214_p_spl_0
  );


  buf

  (
    ffc_214_p_spl_000,
    ffc_214_p_spl_00
  );


  buf

  (
    ffc_214_p_spl_01,
    ffc_214_p_spl_0
  );


  buf

  (
    ffc_214_p_spl_1,
    ffc_214_p_spl_
  );


  buf

  (
    ffc_214_p_spl_10,
    ffc_214_p_spl_1
  );


  buf

  (
    ffc_214_p_spl_11,
    ffc_214_p_spl_1
  );


  buf

  (
    ffc_68_n_spl_,
    ffc_68_n
  );


  buf

  (
    ffc_68_n_spl_0,
    ffc_68_n_spl_
  );


  buf

  (
    ffc_214_n_spl_,
    ffc_214_n
  );


  buf

  (
    ffc_214_n_spl_0,
    ffc_214_n_spl_
  );


  buf

  (
    ffc_214_n_spl_00,
    ffc_214_n_spl_0
  );


  buf

  (
    ffc_214_n_spl_000,
    ffc_214_n_spl_00
  );


  buf

  (
    ffc_214_n_spl_01,
    ffc_214_n_spl_0
  );


  buf

  (
    ffc_214_n_spl_1,
    ffc_214_n_spl_
  );


  buf

  (
    ffc_214_n_spl_10,
    ffc_214_n_spl_1
  );


  buf

  (
    ffc_214_n_spl_11,
    ffc_214_n_spl_1
  );


  buf

  (
    ffc_267_n_spl_,
    ffc_267_n
  );


  buf

  (
    ffc_278_n_spl_,
    ffc_278_n
  );


  buf

  (
    ffc_267_p_spl_,
    ffc_267_p
  );


  buf

  (
    ffc_278_p_spl_,
    ffc_278_p
  );


  buf

  (
    g681_n_spl_,
    g681_n
  );


  buf

  (
    g681_p_spl_,
    g681_p
  );


  buf

  (
    g680_n_spl_,
    g680_n
  );


  buf

  (
    g683_p_spl_,
    g683_p
  );


  buf

  (
    g680_p_spl_,
    g680_p
  );


  buf

  (
    g683_n_spl_,
    g683_n
  );


  buf

  (
    g684_n_spl_,
    g684_n
  );


  buf

  (
    g684_p_spl_,
    g684_p
  );


  buf

  (
    g679_n_spl_,
    g679_n
  );


  buf

  (
    g686_p_spl_,
    g686_p
  );


  buf

  (
    g679_p_spl_,
    g679_p
  );


  buf

  (
    g686_n_spl_,
    g686_n
  );


  buf

  (
    g687_n_spl_,
    g687_n
  );


  buf

  (
    g687_p_spl_,
    g687_p
  );


  buf

  (
    g678_n_spl_,
    g678_n
  );


  buf

  (
    g689_p_spl_,
    g689_p
  );


  buf

  (
    g678_p_spl_,
    g678_p
  );


  buf

  (
    g689_n_spl_,
    g689_n
  );


  buf

  (
    g690_n_spl_,
    g690_n
  );


  buf

  (
    g690_p_spl_,
    g690_p
  );


  buf

  (
    g677_n_spl_,
    g677_n
  );


  buf

  (
    g692_p_spl_,
    g692_p
  );


  buf

  (
    g677_p_spl_,
    g677_p
  );


  buf

  (
    g692_n_spl_,
    g692_n
  );


  buf

  (
    g693_n_spl_,
    g693_n
  );


  buf

  (
    g693_p_spl_,
    g693_p
  );


  buf

  (
    g676_n_spl_,
    g676_n
  );


  buf

  (
    g695_p_spl_,
    g695_p
  );


  buf

  (
    g676_p_spl_,
    g676_p
  );


  buf

  (
    g695_n_spl_,
    g695_n
  );


  buf

  (
    g696_n_spl_,
    g696_n
  );


  buf

  (
    g696_p_spl_,
    g696_p
  );


  buf

  (
    g675_n_spl_,
    g675_n
  );


  buf

  (
    g698_p_spl_,
    g698_p
  );


  buf

  (
    g673_p_spl_,
    g673_p
  );


  buf

  (
    g672_p_spl_,
    g672_p
  );


  buf

  (
    ffc_17_p_spl_,
    ffc_17_p
  );


  buf

  (
    ffc_17_p_spl_0,
    ffc_17_p_spl_
  );


  buf

  (
    ffc_17_p_spl_00,
    ffc_17_p_spl_0
  );


  buf

  (
    ffc_17_p_spl_000,
    ffc_17_p_spl_00
  );


  buf

  (
    ffc_17_p_spl_001,
    ffc_17_p_spl_00
  );


  buf

  (
    ffc_17_p_spl_01,
    ffc_17_p_spl_0
  );


  buf

  (
    ffc_17_p_spl_010,
    ffc_17_p_spl_01
  );


  buf

  (
    ffc_17_p_spl_011,
    ffc_17_p_spl_01
  );


  buf

  (
    ffc_17_p_spl_1,
    ffc_17_p_spl_
  );


  buf

  (
    ffc_17_p_spl_10,
    ffc_17_p_spl_1
  );


  buf

  (
    ffc_17_p_spl_100,
    ffc_17_p_spl_10
  );


  buf

  (
    ffc_17_p_spl_11,
    ffc_17_p_spl_1
  );


  buf

  (
    ffc_17_n_spl_,
    ffc_17_n
  );


  buf

  (
    ffc_17_n_spl_0,
    ffc_17_n_spl_
  );


  buf

  (
    ffc_17_n_spl_00,
    ffc_17_n_spl_0
  );


  buf

  (
    ffc_17_n_spl_000,
    ffc_17_n_spl_00
  );


  buf

  (
    ffc_17_n_spl_001,
    ffc_17_n_spl_00
  );


  buf

  (
    ffc_17_n_spl_01,
    ffc_17_n_spl_0
  );


  buf

  (
    ffc_17_n_spl_010,
    ffc_17_n_spl_01
  );


  buf

  (
    ffc_17_n_spl_1,
    ffc_17_n_spl_
  );


  buf

  (
    ffc_17_n_spl_10,
    ffc_17_n_spl_1
  );


  buf

  (
    ffc_17_n_spl_11,
    ffc_17_n_spl_1
  );


  buf

  (
    ffc_9_p_spl_,
    ffc_9_p
  );


  buf

  (
    ffc_9_p_spl_0,
    ffc_9_p_spl_
  );


  buf

  (
    ffc_9_p_spl_00,
    ffc_9_p_spl_0
  );


  buf

  (
    ffc_9_p_spl_000,
    ffc_9_p_spl_00
  );


  buf

  (
    ffc_9_p_spl_001,
    ffc_9_p_spl_00
  );


  buf

  (
    ffc_9_p_spl_01,
    ffc_9_p_spl_0
  );


  buf

  (
    ffc_9_p_spl_010,
    ffc_9_p_spl_01
  );


  buf

  (
    ffc_9_p_spl_011,
    ffc_9_p_spl_01
  );


  buf

  (
    ffc_9_p_spl_1,
    ffc_9_p_spl_
  );


  buf

  (
    ffc_9_p_spl_10,
    ffc_9_p_spl_1
  );


  buf

  (
    ffc_9_p_spl_100,
    ffc_9_p_spl_10
  );


  buf

  (
    ffc_9_p_spl_101,
    ffc_9_p_spl_10
  );


  buf

  (
    ffc_9_p_spl_11,
    ffc_9_p_spl_1
  );


  buf

  (
    ffc_9_p_spl_110,
    ffc_9_p_spl_11
  );


  buf

  (
    ffc_9_p_spl_111,
    ffc_9_p_spl_11
  );


  buf

  (
    ffc_9_n_spl_,
    ffc_9_n
  );


  buf

  (
    ffc_9_n_spl_0,
    ffc_9_n_spl_
  );


  buf

  (
    ffc_9_n_spl_00,
    ffc_9_n_spl_0
  );


  buf

  (
    ffc_9_n_spl_000,
    ffc_9_n_spl_00
  );


  buf

  (
    ffc_9_n_spl_001,
    ffc_9_n_spl_00
  );


  buf

  (
    ffc_9_n_spl_01,
    ffc_9_n_spl_0
  );


  buf

  (
    ffc_9_n_spl_010,
    ffc_9_n_spl_01
  );


  buf

  (
    ffc_9_n_spl_011,
    ffc_9_n_spl_01
  );


  buf

  (
    ffc_9_n_spl_1,
    ffc_9_n_spl_
  );


  buf

  (
    ffc_9_n_spl_10,
    ffc_9_n_spl_1
  );


  buf

  (
    ffc_9_n_spl_100,
    ffc_9_n_spl_10
  );


  buf

  (
    ffc_9_n_spl_101,
    ffc_9_n_spl_10
  );


  buf

  (
    ffc_9_n_spl_11,
    ffc_9_n_spl_1
  );


  buf

  (
    ffc_9_n_spl_110,
    ffc_9_n_spl_11
  );


  buf

  (
    ffc_9_n_spl_111,
    ffc_9_n_spl_11
  );


  buf

  (
    ffc_264_n_spl_,
    ffc_264_n
  );


  buf

  (
    ffc_281_p_spl_,
    ffc_281_p
  );


  buf

  (
    ffc_264_p_spl_,
    ffc_264_p
  );


  buf

  (
    ffc_281_n_spl_,
    ffc_281_n
  );


  buf

  (
    g706_n_spl_,
    g706_n
  );


  buf

  (
    g706_p_spl_,
    g706_p
  );


  buf

  (
    g705_n_spl_,
    g705_n
  );


  buf

  (
    g708_p_spl_,
    g708_p
  );


  buf

  (
    g705_p_spl_,
    g705_p
  );


  buf

  (
    g708_n_spl_,
    g708_n
  );


  buf

  (
    ffc_75_p_spl_,
    ffc_75_p
  );


  buf

  (
    ffc_75_p_spl_0,
    ffc_75_p_spl_
  );


  buf

  (
    ffc_75_p_spl_1,
    ffc_75_p_spl_
  );


  buf

  (
    ffc_160_p_spl_,
    ffc_160_p
  );


  buf

  (
    ffc_160_p_spl_0,
    ffc_160_p_spl_
  );


  buf

  (
    ffc_160_p_spl_1,
    ffc_160_p_spl_
  );


  buf

  (
    ffc_75_n_spl_,
    ffc_75_n
  );


  buf

  (
    ffc_75_n_spl_0,
    ffc_75_n_spl_
  );


  buf

  (
    ffc_160_n_spl_,
    ffc_160_n
  );


  buf

  (
    ffc_160_n_spl_0,
    ffc_160_n_spl_
  );


  buf

  (
    ffc_160_n_spl_1,
    ffc_160_n_spl_
  );


  buf

  (
    g709_n_spl_,
    g709_n
  );


  buf

  (
    g709_p_spl_,
    g709_p
  );


  buf

  (
    g710_n_spl_,
    g710_n
  );


  buf

  (
    g712_p_spl_,
    g712_p
  );


  buf

  (
    g710_p_spl_,
    g710_p
  );


  buf

  (
    g712_n_spl_,
    g712_n
  );


  buf

  (
    g713_n_spl_,
    g713_n
  );


  buf

  (
    g713_p_spl_,
    g713_p
  );


  buf

  (
    ffc_76_p_spl_,
    ffc_76_p
  );


  buf

  (
    ffc_76_p_spl_0,
    ffc_76_p_spl_
  );


  buf

  (
    ffc_76_n_spl_,
    ffc_76_n
  );


  buf

  (
    ffc_76_n_spl_0,
    ffc_76_n_spl_
  );


  buf

  (
    ffc_77_p_spl_,
    ffc_77_p
  );


  buf

  (
    ffc_77_p_spl_0,
    ffc_77_p_spl_
  );


  buf

  (
    ffc_77_p_spl_1,
    ffc_77_p_spl_
  );


  buf

  (
    ffc_77_n_spl_,
    ffc_77_n
  );


  buf

  (
    ffc_77_n_spl_0,
    ffc_77_n_spl_
  );


  buf

  (
    g716_n_spl_,
    g716_n
  );


  buf

  (
    g717_n_spl_,
    g717_n
  );


  buf

  (
    g716_p_spl_,
    g716_p
  );


  buf

  (
    g717_p_spl_,
    g717_p
  );


  buf

  (
    g718_n_spl_,
    g718_n
  );


  buf

  (
    g718_p_spl_,
    g718_p
  );


  buf

  (
    g715_n_spl_,
    g715_n
  );


  buf

  (
    g720_p_spl_,
    g720_p
  );


  buf

  (
    g715_p_spl_,
    g715_p
  );


  buf

  (
    g720_n_spl_,
    g720_n
  );


  buf

  (
    g721_n_spl_,
    g721_n
  );


  buf

  (
    g721_p_spl_,
    g721_p
  );


  buf

  (
    g714_n_spl_,
    g714_n
  );


  buf

  (
    g723_p_spl_,
    g723_p
  );


  buf

  (
    g714_p_spl_,
    g714_p
  );


  buf

  (
    g723_n_spl_,
    g723_n
  );


  buf

  (
    ffc_174_p_spl_,
    ffc_174_p
  );


  buf

  (
    ffc_174_p_spl_0,
    ffc_174_p_spl_
  );


  buf

  (
    ffc_174_p_spl_00,
    ffc_174_p_spl_0
  );


  buf

  (
    ffc_174_p_spl_01,
    ffc_174_p_spl_0
  );


  buf

  (
    ffc_174_p_spl_1,
    ffc_174_p_spl_
  );


  buf

  (
    ffc_174_p_spl_10,
    ffc_174_p_spl_1
  );


  buf

  (
    ffc_174_n_spl_,
    ffc_174_n
  );


  buf

  (
    ffc_174_n_spl_0,
    ffc_174_n_spl_
  );


  buf

  (
    ffc_174_n_spl_00,
    ffc_174_n_spl_0
  );


  buf

  (
    ffc_174_n_spl_01,
    ffc_174_n_spl_0
  );


  buf

  (
    ffc_174_n_spl_1,
    ffc_174_n_spl_
  );


  buf

  (
    ffc_174_n_spl_10,
    ffc_174_n_spl_1
  );


  buf

  (
    g724_n_spl_,
    g724_n
  );


  buf

  (
    g724_p_spl_,
    g724_p
  );


  buf

  (
    g725_n_spl_,
    g725_n
  );


  buf

  (
    g727_p_spl_,
    g727_p
  );


  buf

  (
    g725_p_spl_,
    g725_p
  );


  buf

  (
    g727_n_spl_,
    g727_n
  );


  buf

  (
    g728_n_spl_,
    g728_n
  );


  buf

  (
    g728_p_spl_,
    g728_p
  );


  buf

  (
    g731_n_spl_,
    g731_n
  );


  buf

  (
    g732_n_spl_,
    g732_n
  );


  buf

  (
    g731_p_spl_,
    g731_p
  );


  buf

  (
    g732_p_spl_,
    g732_p
  );


  buf

  (
    g733_n_spl_,
    g733_n
  );


  buf

  (
    g733_p_spl_,
    g733_p
  );


  buf

  (
    g730_n_spl_,
    g730_n
  );


  buf

  (
    g735_p_spl_,
    g735_p
  );


  buf

  (
    g730_p_spl_,
    g730_p
  );


  buf

  (
    g735_n_spl_,
    g735_n
  );


  buf

  (
    g736_n_spl_,
    g736_n
  );


  buf

  (
    g736_p_spl_,
    g736_p
  );


  buf

  (
    g729_n_spl_,
    g729_n
  );


  buf

  (
    g738_p_spl_,
    g738_p
  );


  buf

  (
    g729_p_spl_,
    g729_p
  );


  buf

  (
    g738_n_spl_,
    g738_n
  );


  buf

  (
    ffc_263_n_spl_,
    ffc_263_n
  );


  buf

  (
    ffc_282_p_spl_,
    ffc_282_p
  );


  buf

  (
    ffc_263_p_spl_,
    ffc_263_p
  );


  buf

  (
    ffc_282_n_spl_,
    ffc_282_n
  );


  buf

  (
    g741_n_spl_,
    g741_n
  );


  buf

  (
    g741_p_spl_,
    g741_p
  );


  buf

  (
    g740_n_spl_,
    g740_n
  );


  buf

  (
    g743_p_spl_,
    g743_p
  );


  buf

  (
    g740_p_spl_,
    g740_p
  );


  buf

  (
    g743_n_spl_,
    g743_n
  );


  buf

  (
    ffc_72_p_spl_,
    ffc_72_p
  );


  buf

  (
    ffc_72_p_spl_0,
    ffc_72_p_spl_
  );


  buf

  (
    ffc_72_p_spl_1,
    ffc_72_p_spl_
  );


  buf

  (
    ffc_72_n_spl_,
    ffc_72_n
  );


  buf

  (
    ffc_72_n_spl_0,
    ffc_72_n_spl_
  );


  buf

  (
    g744_n_spl_,
    g744_n
  );


  buf

  (
    g744_p_spl_,
    g744_p
  );


  buf

  (
    g745_n_spl_,
    g745_n
  );


  buf

  (
    g747_p_spl_,
    g747_p
  );


  buf

  (
    g745_p_spl_,
    g745_p
  );


  buf

  (
    g747_n_spl_,
    g747_n
  );


  buf

  (
    g748_n_spl_,
    g748_n
  );


  buf

  (
    g748_p_spl_,
    g748_p
  );


  buf

  (
    ffc_73_p_spl_,
    ffc_73_p
  );


  buf

  (
    ffc_73_p_spl_0,
    ffc_73_p_spl_
  );


  buf

  (
    ffc_73_n_spl_,
    ffc_73_n
  );


  buf

  (
    ffc_73_n_spl_0,
    ffc_73_n_spl_
  );


  buf

  (
    ffc_74_p_spl_,
    ffc_74_p
  );


  buf

  (
    ffc_74_p_spl_0,
    ffc_74_p_spl_
  );


  buf

  (
    ffc_74_p_spl_1,
    ffc_74_p_spl_
  );


  buf

  (
    ffc_74_n_spl_,
    ffc_74_n
  );


  buf

  (
    ffc_74_n_spl_0,
    ffc_74_n_spl_
  );


  buf

  (
    ffc_265_n_spl_,
    ffc_265_n
  );


  buf

  (
    ffc_280_n_spl_,
    ffc_280_n
  );


  buf

  (
    ffc_265_p_spl_,
    ffc_265_p
  );


  buf

  (
    ffc_280_p_spl_,
    ffc_280_p
  );


  buf

  (
    g753_n_spl_,
    g753_n
  );


  buf

  (
    g753_p_spl_,
    g753_p
  );


  buf

  (
    g752_n_spl_,
    g752_n
  );


  buf

  (
    g755_p_spl_,
    g755_p
  );


  buf

  (
    g752_p_spl_,
    g752_p
  );


  buf

  (
    g755_n_spl_,
    g755_n
  );


  buf

  (
    g756_n_spl_,
    g756_n
  );


  buf

  (
    g756_p_spl_,
    g756_p
  );


  buf

  (
    g751_n_spl_,
    g751_n
  );


  buf

  (
    g758_p_spl_,
    g758_p
  );


  buf

  (
    g751_p_spl_,
    g751_p
  );


  buf

  (
    g758_n_spl_,
    g758_n
  );


  buf

  (
    g759_n_spl_,
    g759_n
  );


  buf

  (
    g759_p_spl_,
    g759_p
  );


  buf

  (
    g750_n_spl_,
    g750_n
  );


  buf

  (
    g761_p_spl_,
    g761_p
  );


  buf

  (
    g750_p_spl_,
    g750_p
  );


  buf

  (
    g761_n_spl_,
    g761_n
  );


  buf

  (
    g762_n_spl_,
    g762_n
  );


  buf

  (
    g762_p_spl_,
    g762_p
  );


  buf

  (
    g749_n_spl_,
    g749_n
  );


  buf

  (
    g764_p_spl_,
    g764_p
  );


  buf

  (
    g749_p_spl_,
    g749_p
  );


  buf

  (
    g764_n_spl_,
    g764_n
  );


  buf

  (
    g765_n_spl_,
    g765_n
  );


  buf

  (
    g765_p_spl_,
    g765_p
  );


  buf

  (
    g766_n_spl_,
    g766_n
  );


  buf

  (
    g768_p_spl_,
    g768_p
  );


  buf

  (
    g766_p_spl_,
    g766_p
  );


  buf

  (
    g768_n_spl_,
    g768_n
  );


  buf

  (
    g769_n_spl_,
    g769_n
  );


  buf

  (
    g769_p_spl_,
    g769_p
  );


  buf

  (
    g774_n_spl_,
    g774_n
  );


  buf

  (
    g776_p_spl_,
    g776_p
  );


  buf

  (
    g774_p_spl_,
    g774_p
  );


  buf

  (
    g776_n_spl_,
    g776_n
  );


  buf

  (
    g777_n_spl_,
    g777_n
  );


  buf

  (
    g777_p_spl_,
    g777_p
  );


  buf

  (
    g773_n_spl_,
    g773_n
  );


  buf

  (
    g779_p_spl_,
    g779_p
  );


  buf

  (
    g773_p_spl_,
    g773_p
  );


  buf

  (
    g779_n_spl_,
    g779_n
  );


  buf

  (
    g780_n_spl_,
    g780_n
  );


  buf

  (
    g780_p_spl_,
    g780_p
  );


  buf

  (
    g772_n_spl_,
    g772_n
  );


  buf

  (
    g782_p_spl_,
    g782_p
  );


  buf

  (
    g772_p_spl_,
    g772_p
  );


  buf

  (
    g782_n_spl_,
    g782_n
  );


  buf

  (
    g783_n_spl_,
    g783_n
  );


  buf

  (
    g783_p_spl_,
    g783_p
  );


  buf

  (
    g771_n_spl_,
    g771_n
  );


  buf

  (
    g785_p_spl_,
    g785_p
  );


  buf

  (
    g771_p_spl_,
    g771_p
  );


  buf

  (
    g785_n_spl_,
    g785_n
  );


  buf

  (
    g786_n_spl_,
    g786_n
  );


  buf

  (
    g786_p_spl_,
    g786_p
  );


  buf

  (
    g770_n_spl_,
    g770_n
  );


  buf

  (
    g788_p_spl_,
    g788_p
  );


  buf

  (
    g770_p_spl_,
    g770_p
  );


  buf

  (
    g788_n_spl_,
    g788_n
  );


  buf

  (
    ffc_262_n_spl_,
    ffc_262_n
  );


  buf

  (
    ffc_283_p_spl_,
    ffc_283_p
  );


  buf

  (
    ffc_262_p_spl_,
    ffc_262_p
  );


  buf

  (
    ffc_283_n_spl_,
    ffc_283_n
  );


  buf

  (
    g791_n_spl_,
    g791_n
  );


  buf

  (
    g791_p_spl_,
    g791_p
  );


  buf

  (
    g790_n_spl_,
    g790_n
  );


  buf

  (
    g793_p_spl_,
    g793_p
  );


  buf

  (
    g790_p_spl_,
    g790_p
  );


  buf

  (
    g793_n_spl_,
    g793_n
  );


  buf

  (
    ffc_69_p_spl_,
    ffc_69_p
  );


  buf

  (
    ffc_69_p_spl_0,
    ffc_69_p_spl_
  );


  buf

  (
    ffc_69_n_spl_,
    ffc_69_n
  );


  buf

  (
    ffc_69_n_spl_0,
    ffc_69_n_spl_
  );


  buf

  (
    g794_n_spl_,
    g794_n
  );


  buf

  (
    g794_p_spl_,
    g794_p
  );


  buf

  (
    g795_n_spl_,
    g795_n
  );


  buf

  (
    g797_p_spl_,
    g797_p
  );


  buf

  (
    g795_p_spl_,
    g795_p
  );


  buf

  (
    g797_n_spl_,
    g797_n
  );


  buf

  (
    g798_n_spl_,
    g798_n
  );


  buf

  (
    g798_p_spl_,
    g798_p
  );


  buf

  (
    ffc_70_p_spl_,
    ffc_70_p
  );


  buf

  (
    ffc_70_n_spl_,
    ffc_70_n
  );


  buf

  (
    ffc_70_n_spl_0,
    ffc_70_n_spl_
  );


  buf

  (
    ffc_71_p_spl_,
    ffc_71_p
  );


  buf

  (
    ffc_71_p_spl_0,
    ffc_71_p_spl_
  );


  buf

  (
    ffc_71_p_spl_1,
    ffc_71_p_spl_
  );


  buf

  (
    ffc_71_n_spl_,
    ffc_71_n
  );


  buf

  (
    ffc_71_n_spl_0,
    ffc_71_n_spl_
  );


  buf

  (
    ffc_266_n_spl_,
    ffc_266_n
  );


  buf

  (
    ffc_279_n_spl_,
    ffc_279_n
  );


  buf

  (
    ffc_266_p_spl_,
    ffc_266_p
  );


  buf

  (
    ffc_279_p_spl_,
    ffc_279_p
  );


  buf

  (
    g803_n_spl_,
    g803_n
  );


  buf

  (
    g803_p_spl_,
    g803_p
  );


  buf

  (
    g802_n_spl_,
    g802_n
  );


  buf

  (
    g805_p_spl_,
    g805_p
  );


  buf

  (
    g802_p_spl_,
    g802_p
  );


  buf

  (
    g805_n_spl_,
    g805_n
  );


  buf

  (
    g806_n_spl_,
    g806_n
  );


  buf

  (
    g806_p_spl_,
    g806_p
  );


  buf

  (
    g801_n_spl_,
    g801_n
  );


  buf

  (
    g808_p_spl_,
    g808_p
  );


  buf

  (
    g801_p_spl_,
    g801_p
  );


  buf

  (
    g808_n_spl_,
    g808_n
  );


  buf

  (
    g809_n_spl_,
    g809_n
  );


  buf

  (
    g809_p_spl_,
    g809_p
  );


  buf

  (
    g800_n_spl_,
    g800_n
  );


  buf

  (
    g811_p_spl_,
    g811_p
  );


  buf

  (
    g800_p_spl_,
    g800_p
  );


  buf

  (
    g811_n_spl_,
    g811_n
  );


  buf

  (
    g812_n_spl_,
    g812_n
  );


  buf

  (
    g812_p_spl_,
    g812_p
  );


  buf

  (
    g799_n_spl_,
    g799_n
  );


  buf

  (
    g814_p_spl_,
    g814_p
  );


  buf

  (
    g799_p_spl_,
    g799_p
  );


  buf

  (
    g814_n_spl_,
    g814_n
  );


  buf

  (
    g815_n_spl_,
    g815_n
  );


  buf

  (
    g815_p_spl_,
    g815_p
  );


  buf

  (
    g816_n_spl_,
    g816_n
  );


  buf

  (
    g818_p_spl_,
    g818_p
  );


  buf

  (
    g816_p_spl_,
    g816_p
  );


  buf

  (
    g818_n_spl_,
    g818_n
  );


  buf

  (
    g819_n_spl_,
    g819_n
  );


  buf

  (
    g819_p_spl_,
    g819_p
  );


  buf

  (
    g824_n_spl_,
    g824_n
  );


  buf

  (
    g826_p_spl_,
    g826_p
  );


  buf

  (
    g824_p_spl_,
    g824_p
  );


  buf

  (
    g826_n_spl_,
    g826_n
  );


  buf

  (
    g827_n_spl_,
    g827_n
  );


  buf

  (
    g827_p_spl_,
    g827_p
  );


  buf

  (
    g823_n_spl_,
    g823_n
  );


  buf

  (
    g829_p_spl_,
    g829_p
  );


  buf

  (
    g823_p_spl_,
    g823_p
  );


  buf

  (
    g829_n_spl_,
    g829_n
  );


  buf

  (
    g830_n_spl_,
    g830_n
  );


  buf

  (
    g830_p_spl_,
    g830_p
  );


  buf

  (
    g822_n_spl_,
    g822_n
  );


  buf

  (
    g832_p_spl_,
    g832_p
  );


  buf

  (
    g822_p_spl_,
    g822_p
  );


  buf

  (
    g832_n_spl_,
    g832_n
  );


  buf

  (
    g833_n_spl_,
    g833_n
  );


  buf

  (
    g833_p_spl_,
    g833_p
  );


  buf

  (
    g821_n_spl_,
    g821_n
  );


  buf

  (
    g835_p_spl_,
    g835_p
  );


  buf

  (
    g821_p_spl_,
    g821_p
  );


  buf

  (
    g835_n_spl_,
    g835_n
  );


  buf

  (
    g836_n_spl_,
    g836_n
  );


  buf

  (
    g836_p_spl_,
    g836_p
  );


  buf

  (
    g820_n_spl_,
    g820_n
  );


  buf

  (
    g838_p_spl_,
    g838_p
  );


  buf

  (
    g820_p_spl_,
    g820_p
  );


  buf

  (
    g838_n_spl_,
    g838_n
  );


  buf

  (
    g674_n_spl_,
    g674_n
  );


  buf

  (
    g701_p_spl_,
    g701_p
  );


  buf

  (
    g671_p_spl_,
    g671_p
  );


  buf

  (
    ffc_118_p_spl_,
    ffc_118_p
  );


  buf

  (
    ffc_118_p_spl_0,
    ffc_118_p_spl_
  );


  buf

  (
    ffc_118_p_spl_00,
    ffc_118_p_spl_0
  );


  buf

  (
    ffc_118_p_spl_01,
    ffc_118_p_spl_0
  );


  buf

  (
    ffc_118_p_spl_1,
    ffc_118_p_spl_
  );


  buf

  (
    ffc_118_n_spl_,
    ffc_118_n
  );


  buf

  (
    ffc_118_n_spl_0,
    ffc_118_n_spl_
  );


  buf

  (
    ffc_118_n_spl_00,
    ffc_118_n_spl_0
  );


  buf

  (
    ffc_118_n_spl_1,
    ffc_118_n_spl_
  );


  buf

  (
    ffc_296_p_spl_,
    ffc_296_p
  );


  buf

  (
    ffc_296_n_spl_,
    ffc_296_n
  );


  buf

  (
    g844_n_spl_,
    g844_n
  );


  buf

  (
    g845_p_spl_,
    g845_p
  );


  buf

  (
    g844_p_spl_,
    g844_p
  );


  buf

  (
    g845_n_spl_,
    g845_n
  );


  buf

  (
    g846_n_spl_,
    g846_n
  );


  buf

  (
    g846_p_spl_,
    g846_p
  );


  buf

  (
    g843_n_spl_,
    g843_n
  );


  buf

  (
    g848_p_spl_,
    g848_p
  );


  buf

  (
    g843_p_spl_,
    g843_p
  );


  buf

  (
    g848_n_spl_,
    g848_n
  );


  buf

  (
    g849_n_spl_,
    g849_n
  );


  buf

  (
    g849_p_spl_,
    g849_p
  );


  buf

  (
    g842_n_spl_,
    g842_n
  );


  buf

  (
    g851_p_spl_,
    g851_p
  );


  buf

  (
    g842_p_spl_,
    g842_p
  );


  buf

  (
    g851_n_spl_,
    g851_n
  );


  buf

  (
    g852_n_spl_,
    g852_n
  );


  buf

  (
    g852_p_spl_,
    g852_p
  );


  buf

  (
    g841_n_spl_,
    g841_n
  );


  buf

  (
    g854_p_spl_,
    g854_p
  );


  buf

  (
    g841_p_spl_,
    g841_p
  );


  buf

  (
    g854_n_spl_,
    g854_n
  );


  buf

  (
    g855_n_spl_,
    g855_n
  );


  buf

  (
    g855_p_spl_,
    g855_p
  );


  buf

  (
    g702_p_spl_,
    g702_p
  );


  buf

  (
    ffc_339_n_spl_,
    ffc_339_n
  );


  buf

  (
    ffc_355_p_spl_,
    ffc_355_p
  );


  buf

  (
    ffc_339_p_spl_,
    ffc_339_p
  );


  buf

  (
    ffc_355_n_spl_,
    ffc_355_n
  );


  buf

  (
    g859_n_spl_,
    g859_n
  );


  buf

  (
    g859_p_spl_,
    g859_p
  );


  buf

  (
    g858_n_spl_,
    g858_n
  );


  buf

  (
    g861_p_spl_,
    g861_p
  );


  buf

  (
    g858_p_spl_,
    g858_p
  );


  buf

  (
    g861_n_spl_,
    g861_n
  );


  buf

  (
    g862_n_spl_,
    g862_n
  );


  buf

  (
    g862_p_spl_,
    g862_p
  );


  buf

  (
    g857_p_spl_,
    g857_p
  );


  buf

  (
    g703_p_spl_,
    g703_p
  );


  buf

  (
    g864_p_spl_,
    g864_p
  );


  buf

  (
    g704_p_spl_,
    g704_p
  );


  buf

  (
    g840_p_spl_,
    g840_p
  );


  buf

  (
    g872_n_spl_,
    g872_n
  );


  buf

  (
    g874_p_spl_,
    g874_p
  );


  buf

  (
    g872_p_spl_,
    g872_p
  );


  buf

  (
    g874_n_spl_,
    g874_n
  );


  buf

  (
    g875_n_spl_,
    g875_n
  );


  buf

  (
    g875_p_spl_,
    g875_p
  );


  buf

  (
    g871_n_spl_,
    g871_n
  );


  buf

  (
    g877_p_spl_,
    g877_p
  );


  buf

  (
    g871_p_spl_,
    g871_p
  );


  buf

  (
    g877_n_spl_,
    g877_n
  );


  buf

  (
    g878_n_spl_,
    g878_n
  );


  buf

  (
    g878_p_spl_,
    g878_p
  );


  buf

  (
    g870_n_spl_,
    g870_n
  );


  buf

  (
    g880_p_spl_,
    g880_p
  );


  buf

  (
    g870_p_spl_,
    g870_p
  );


  buf

  (
    g880_n_spl_,
    g880_n
  );


  buf

  (
    g881_n_spl_,
    g881_n
  );


  buf

  (
    g881_p_spl_,
    g881_p
  );


  buf

  (
    g869_n_spl_,
    g869_n
  );


  buf

  (
    g883_p_spl_,
    g883_p
  );


  buf

  (
    g869_p_spl_,
    g869_p
  );


  buf

  (
    g883_n_spl_,
    g883_n
  );


  buf

  (
    g884_n_spl_,
    g884_n
  );


  buf

  (
    g884_p_spl_,
    g884_p
  );


  buf

  (
    g868_n_spl_,
    g868_n
  );


  buf

  (
    g886_p_spl_,
    g886_p
  );


  buf

  (
    ffc_10_p_spl_,
    ffc_10_p
  );


  buf

  (
    ffc_10_p_spl_0,
    ffc_10_p_spl_
  );


  buf

  (
    ffc_10_p_spl_00,
    ffc_10_p_spl_0
  );


  buf

  (
    ffc_10_p_spl_000,
    ffc_10_p_spl_00
  );


  buf

  (
    ffc_10_p_spl_001,
    ffc_10_p_spl_00
  );


  buf

  (
    ffc_10_p_spl_01,
    ffc_10_p_spl_0
  );


  buf

  (
    ffc_10_p_spl_010,
    ffc_10_p_spl_01
  );


  buf

  (
    ffc_10_p_spl_011,
    ffc_10_p_spl_01
  );


  buf

  (
    ffc_10_p_spl_1,
    ffc_10_p_spl_
  );


  buf

  (
    ffc_10_p_spl_10,
    ffc_10_p_spl_1
  );


  buf

  (
    ffc_10_p_spl_100,
    ffc_10_p_spl_10
  );


  buf

  (
    ffc_10_p_spl_101,
    ffc_10_p_spl_10
  );


  buf

  (
    ffc_10_p_spl_11,
    ffc_10_p_spl_1
  );


  buf

  (
    ffc_10_p_spl_110,
    ffc_10_p_spl_11
  );


  buf

  (
    ffc_10_n_spl_,
    ffc_10_n
  );


  buf

  (
    ffc_10_n_spl_0,
    ffc_10_n_spl_
  );


  buf

  (
    ffc_10_n_spl_00,
    ffc_10_n_spl_0
  );


  buf

  (
    ffc_10_n_spl_000,
    ffc_10_n_spl_00
  );


  buf

  (
    ffc_10_n_spl_001,
    ffc_10_n_spl_00
  );


  buf

  (
    ffc_10_n_spl_01,
    ffc_10_n_spl_0
  );


  buf

  (
    ffc_10_n_spl_010,
    ffc_10_n_spl_01
  );


  buf

  (
    ffc_10_n_spl_011,
    ffc_10_n_spl_01
  );


  buf

  (
    ffc_10_n_spl_1,
    ffc_10_n_spl_
  );


  buf

  (
    ffc_10_n_spl_10,
    ffc_10_n_spl_1
  );


  buf

  (
    ffc_10_n_spl_100,
    ffc_10_n_spl_10
  );


  buf

  (
    ffc_10_n_spl_101,
    ffc_10_n_spl_10
  );


  buf

  (
    ffc_10_n_spl_11,
    ffc_10_n_spl_1
  );


  buf

  (
    ffc_10_n_spl_110,
    ffc_10_n_spl_11
  );


  buf

  (
    ffc_10_n_spl_111,
    ffc_10_n_spl_11
  );


  buf

  (
    g866_p_spl_,
    g866_p
  );


  buf

  (
    ffc_195_p_spl_,
    ffc_195_p
  );


  buf

  (
    ffc_195_p_spl_0,
    ffc_195_p_spl_
  );


  buf

  (
    ffc_195_p_spl_00,
    ffc_195_p_spl_0
  );


  buf

  (
    ffc_195_p_spl_1,
    ffc_195_p_spl_
  );


  buf

  (
    ffc_195_n_spl_,
    ffc_195_n
  );


  buf

  (
    ffc_195_n_spl_0,
    ffc_195_n_spl_
  );


  buf

  (
    ffc_195_n_spl_1,
    ffc_195_n_spl_
  );


  buf

  (
    ffc_326_n_spl_,
    ffc_326_n
  );


  buf

  (
    ffc_343_p_spl_,
    ffc_343_p
  );


  buf

  (
    ffc_326_p_spl_,
    ffc_326_p
  );


  buf

  (
    ffc_343_n_spl_,
    ffc_343_n
  );


  buf

  (
    g894_n_spl_,
    g894_n
  );


  buf

  (
    g894_p_spl_,
    g894_p
  );


  buf

  (
    g893_n_spl_,
    g893_n
  );


  buf

  (
    g896_p_spl_,
    g896_p
  );


  buf

  (
    g893_p_spl_,
    g893_p
  );


  buf

  (
    g896_n_spl_,
    g896_n
  );


  buf

  (
    g897_n_spl_,
    g897_n
  );


  buf

  (
    g897_p_spl_,
    g897_p
  );


  buf

  (
    g892_n_spl_,
    g892_n
  );


  buf

  (
    g899_p_spl_,
    g899_p
  );


  buf

  (
    g892_p_spl_,
    g892_p
  );


  buf

  (
    g899_n_spl_,
    g899_n
  );


  buf

  (
    g900_n_spl_,
    g900_n
  );


  buf

  (
    g900_p_spl_,
    g900_p
  );


  buf

  (
    g891_n_spl_,
    g891_n
  );


  buf

  (
    g902_p_spl_,
    g902_p
  );


  buf

  (
    g891_p_spl_,
    g891_p
  );


  buf

  (
    g902_n_spl_,
    g902_n
  );


  buf

  (
    g903_n_spl_,
    g903_n
  );


  buf

  (
    g903_p_spl_,
    g903_p
  );


  buf

  (
    g905_p_spl_,
    g905_p
  );


  buf

  (
    g890_p_spl_,
    g890_p
  );


  buf

  (
    ffc_19_p_spl_,
    ffc_19_p
  );


  buf

  (
    ffc_19_p_spl_0,
    ffc_19_p_spl_
  );


  buf

  (
    ffc_19_p_spl_00,
    ffc_19_p_spl_0
  );


  buf

  (
    ffc_19_p_spl_000,
    ffc_19_p_spl_00
  );


  buf

  (
    ffc_19_p_spl_001,
    ffc_19_p_spl_00
  );


  buf

  (
    ffc_19_p_spl_01,
    ffc_19_p_spl_0
  );


  buf

  (
    ffc_19_p_spl_1,
    ffc_19_p_spl_
  );


  buf

  (
    ffc_19_p_spl_10,
    ffc_19_p_spl_1
  );


  buf

  (
    ffc_19_p_spl_11,
    ffc_19_p_spl_1
  );


  buf

  (
    ffc_19_n_spl_,
    ffc_19_n
  );


  buf

  (
    ffc_19_n_spl_0,
    ffc_19_n_spl_
  );


  buf

  (
    ffc_19_n_spl_00,
    ffc_19_n_spl_0
  );


  buf

  (
    ffc_19_n_spl_01,
    ffc_19_n_spl_0
  );


  buf

  (
    ffc_19_n_spl_1,
    ffc_19_n_spl_
  );


  buf

  (
    ffc_19_n_spl_10,
    ffc_19_n_spl_1
  );


  buf

  (
    ffc_19_n_spl_11,
    ffc_19_n_spl_1
  );


  buf

  (
    g839_n_spl_,
    g839_n
  );


  buf

  (
    g789_n_spl_,
    g789_n
  );


  buf

  (
    g739_n_spl_,
    g739_n
  );


  buf

  (
    g925_n_spl_,
    g925_n
  );


  buf

  (
    g927_p_spl_,
    g927_p
  );


  buf

  (
    g925_p_spl_,
    g925_p
  );


  buf

  (
    g927_n_spl_,
    g927_n
  );


  buf

  (
    g928_p_spl_,
    g928_p
  );


  buf

  (
    g924_n_spl_,
    g924_n
  );


  buf

  (
    g930_p_spl_,
    g930_p
  );


  buf

  (
    g924_p_spl_,
    g924_p
  );


  buf

  (
    g930_n_spl_,
    g930_n
  );


  buf

  (
    g931_p_spl_,
    g931_p
  );


  buf

  (
    g937_n_spl_,
    g937_n
  );


  buf

  (
    g939_p_spl_,
    g939_p
  );


  buf

  (
    g937_p_spl_,
    g937_p
  );


  buf

  (
    g939_n_spl_,
    g939_n
  );


  buf

  (
    g940_p_spl_,
    g940_p
  );


  buf

  (
    g936_n_spl_,
    g936_n
  );


  buf

  (
    g942_p_spl_,
    g942_p
  );


  buf

  (
    g936_p_spl_,
    g936_p
  );


  buf

  (
    g942_n_spl_,
    g942_n
  );


  buf

  (
    g943_p_spl_,
    g943_p
  );


  buf

  (
    g949_n_spl_,
    g949_n
  );


  buf

  (
    g951_p_spl_,
    g951_p
  );


  buf

  (
    g949_p_spl_,
    g949_p
  );


  buf

  (
    g951_n_spl_,
    g951_n
  );


  buf

  (
    g952_p_spl_,
    g952_p
  );


  buf

  (
    g948_n_spl_,
    g948_n
  );


  buf

  (
    g954_p_spl_,
    g954_p
  );


  buf

  (
    g948_p_spl_,
    g948_p
  );


  buf

  (
    g954_n_spl_,
    g954_n
  );


  buf

  (
    g955_p_spl_,
    g955_p
  );


  buf

  (
    g867_n_spl_,
    g867_n
  );


  buf

  (
    g889_p_spl_,
    g889_p
  );


  buf

  (
    g865_p_spl_,
    g865_p
  );


  buf

  (
    ffc_119_p_spl_,
    ffc_119_p
  );


  buf

  (
    ffc_119_p_spl_0,
    ffc_119_p_spl_
  );


  buf

  (
    ffc_119_p_spl_00,
    ffc_119_p_spl_0
  );


  buf

  (
    ffc_119_p_spl_01,
    ffc_119_p_spl_0
  );


  buf

  (
    ffc_119_p_spl_1,
    ffc_119_p_spl_
  );


  buf

  (
    ffc_119_n_spl_,
    ffc_119_n
  );


  buf

  (
    ffc_119_n_spl_0,
    ffc_119_n_spl_
  );


  buf

  (
    ffc_119_n_spl_00,
    ffc_119_n_spl_0
  );


  buf

  (
    ffc_119_n_spl_1,
    ffc_119_n_spl_
  );


  buf

  (
    ffc_298_p_spl_,
    ffc_298_p
  );


  buf

  (
    ffc_298_n_spl_,
    ffc_298_n
  );


  buf

  (
    g965_n_spl_,
    g965_n
  );


  buf

  (
    g966_p_spl_,
    g966_p
  );


  buf

  (
    g965_p_spl_,
    g965_p
  );


  buf

  (
    g966_n_spl_,
    g966_n
  );


  buf

  (
    g967_n_spl_,
    g967_n
  );


  buf

  (
    g967_p_spl_,
    g967_p
  );


  buf

  (
    g964_n_spl_,
    g964_n
  );


  buf

  (
    g969_p_spl_,
    g969_p
  );


  buf

  (
    g964_p_spl_,
    g964_p
  );


  buf

  (
    g969_n_spl_,
    g969_n
  );


  buf

  (
    g970_n_spl_,
    g970_n
  );


  buf

  (
    g970_p_spl_,
    g970_p
  );


  buf

  (
    g963_n_spl_,
    g963_n
  );


  buf

  (
    g972_p_spl_,
    g972_p
  );


  buf

  (
    g963_p_spl_,
    g963_p
  );


  buf

  (
    g972_n_spl_,
    g972_n
  );


  buf

  (
    g973_n_spl_,
    g973_n
  );


  buf

  (
    g973_p_spl_,
    g973_p
  );


  buf

  (
    g962_n_spl_,
    g962_n
  );


  buf

  (
    g975_p_spl_,
    g975_p
  );


  buf

  (
    g962_p_spl_,
    g962_p
  );


  buf

  (
    g975_n_spl_,
    g975_n
  );


  buf

  (
    g976_n_spl_,
    g976_n
  );


  buf

  (
    g976_p_spl_,
    g976_p
  );


  buf

  (
    g961_n_spl_,
    g961_n
  );


  buf

  (
    g978_p_spl_,
    g978_p
  );


  buf

  (
    g961_p_spl_,
    g961_p
  );


  buf

  (
    g978_n_spl_,
    g978_n
  );


  buf

  (
    g979_n_spl_,
    g979_n
  );


  buf

  (
    g979_p_spl_,
    g979_p
  );


  buf

  (
    g960_n_spl_,
    g960_n
  );


  buf

  (
    g981_p_spl_,
    g981_p
  );


  buf

  (
    g960_p_spl_,
    g960_p
  );


  buf

  (
    g981_n_spl_,
    g981_n
  );


  buf

  (
    g982_n_spl_,
    g982_n
  );


  buf

  (
    g982_p_spl_,
    g982_p
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G2_p_spl_0,
    G2_p_spl_
  );


  buf

  (
    G2_p_spl_00,
    G2_p_spl_0
  );


  buf

  (
    G2_p_spl_01,
    G2_p_spl_0
  );


  buf

  (
    G2_p_spl_1,
    G2_p_spl_
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    G17_p_spl_0,
    G17_p_spl_
  );


  buf

  (
    G17_p_spl_00,
    G17_p_spl_0
  );


  buf

  (
    G17_p_spl_000,
    G17_p_spl_00
  );


  buf

  (
    G17_p_spl_001,
    G17_p_spl_00
  );


  buf

  (
    G17_p_spl_01,
    G17_p_spl_0
  );


  buf

  (
    G17_p_spl_010,
    G17_p_spl_01
  );


  buf

  (
    G17_p_spl_011,
    G17_p_spl_01
  );


  buf

  (
    G17_p_spl_1,
    G17_p_spl_
  );


  buf

  (
    G17_p_spl_10,
    G17_p_spl_1
  );


  buf

  (
    G17_p_spl_100,
    G17_p_spl_10
  );


  buf

  (
    G17_p_spl_101,
    G17_p_spl_10
  );


  buf

  (
    G17_p_spl_11,
    G17_p_spl_1
  );


  buf

  (
    G17_p_spl_110,
    G17_p_spl_11
  );


  buf

  (
    G17_p_spl_111,
    G17_p_spl_11
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G2_n_spl_0,
    G2_n_spl_
  );


  buf

  (
    G2_n_spl_1,
    G2_n_spl_
  );


  buf

  (
    G17_n_spl_,
    G17_n
  );


  buf

  (
    G17_n_spl_0,
    G17_n_spl_
  );


  buf

  (
    G17_n_spl_00,
    G17_n_spl_0
  );


  buf

  (
    G17_n_spl_000,
    G17_n_spl_00
  );


  buf

  (
    G17_n_spl_001,
    G17_n_spl_00
  );


  buf

  (
    G17_n_spl_01,
    G17_n_spl_0
  );


  buf

  (
    G17_n_spl_010,
    G17_n_spl_01
  );


  buf

  (
    G17_n_spl_011,
    G17_n_spl_01
  );


  buf

  (
    G17_n_spl_1,
    G17_n_spl_
  );


  buf

  (
    G17_n_spl_10,
    G17_n_spl_1
  );


  buf

  (
    G17_n_spl_100,
    G17_n_spl_10
  );


  buf

  (
    G17_n_spl_101,
    G17_n_spl_10
  );


  buf

  (
    G17_n_spl_11,
    G17_n_spl_1
  );


  buf

  (
    G17_n_spl_110,
    G17_n_spl_11
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G1_p_spl_0,
    G1_p_spl_
  );


  buf

  (
    G18_p_spl_,
    G18_p
  );


  buf

  (
    G18_p_spl_0,
    G18_p_spl_
  );


  buf

  (
    G18_p_spl_00,
    G18_p_spl_0
  );


  buf

  (
    G18_p_spl_000,
    G18_p_spl_00
  );


  buf

  (
    G18_p_spl_001,
    G18_p_spl_00
  );


  buf

  (
    G18_p_spl_01,
    G18_p_spl_0
  );


  buf

  (
    G18_p_spl_010,
    G18_p_spl_01
  );


  buf

  (
    G18_p_spl_011,
    G18_p_spl_01
  );


  buf

  (
    G18_p_spl_1,
    G18_p_spl_
  );


  buf

  (
    G18_p_spl_10,
    G18_p_spl_1
  );


  buf

  (
    G18_p_spl_100,
    G18_p_spl_10
  );


  buf

  (
    G18_p_spl_101,
    G18_p_spl_10
  );


  buf

  (
    G18_p_spl_11,
    G18_p_spl_1
  );


  buf

  (
    G18_p_spl_110,
    G18_p_spl_11
  );


  buf

  (
    G18_p_spl_111,
    G18_p_spl_11
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    G18_n_spl_,
    G18_n
  );


  buf

  (
    G18_n_spl_0,
    G18_n_spl_
  );


  buf

  (
    G18_n_spl_00,
    G18_n_spl_0
  );


  buf

  (
    G18_n_spl_000,
    G18_n_spl_00
  );


  buf

  (
    G18_n_spl_001,
    G18_n_spl_00
  );


  buf

  (
    G18_n_spl_01,
    G18_n_spl_0
  );


  buf

  (
    G18_n_spl_010,
    G18_n_spl_01
  );


  buf

  (
    G18_n_spl_011,
    G18_n_spl_01
  );


  buf

  (
    G18_n_spl_1,
    G18_n_spl_
  );


  buf

  (
    G18_n_spl_10,
    G18_n_spl_1
  );


  buf

  (
    G18_n_spl_100,
    G18_n_spl_10
  );


  buf

  (
    G18_n_spl_101,
    G18_n_spl_10
  );


  buf

  (
    G18_n_spl_11,
    G18_n_spl_1
  );


  buf

  (
    G18_n_spl_110,
    G18_n_spl_11
  );


  buf

  (
    G18_n_spl_111,
    G18_n_spl_11
  );


  buf

  (
    g984_p_spl_,
    g984_p
  );


  buf

  (
    g907_p_spl_,
    g907_p
  );


  buf

  (
    ffc_11_p_spl_,
    ffc_11_p
  );


  buf

  (
    ffc_11_p_spl_0,
    ffc_11_p_spl_
  );


  buf

  (
    ffc_11_p_spl_00,
    ffc_11_p_spl_0
  );


  buf

  (
    ffc_11_p_spl_000,
    ffc_11_p_spl_00
  );


  buf

  (
    ffc_11_p_spl_001,
    ffc_11_p_spl_00
  );


  buf

  (
    ffc_11_p_spl_01,
    ffc_11_p_spl_0
  );


  buf

  (
    ffc_11_p_spl_010,
    ffc_11_p_spl_01
  );


  buf

  (
    ffc_11_p_spl_011,
    ffc_11_p_spl_01
  );


  buf

  (
    ffc_11_p_spl_1,
    ffc_11_p_spl_
  );


  buf

  (
    ffc_11_p_spl_10,
    ffc_11_p_spl_1
  );


  buf

  (
    ffc_11_p_spl_100,
    ffc_11_p_spl_10
  );


  buf

  (
    ffc_11_p_spl_101,
    ffc_11_p_spl_10
  );


  buf

  (
    ffc_11_p_spl_11,
    ffc_11_p_spl_1
  );


  buf

  (
    ffc_11_n_spl_,
    ffc_11_n
  );


  buf

  (
    ffc_11_n_spl_0,
    ffc_11_n_spl_
  );


  buf

  (
    ffc_11_n_spl_00,
    ffc_11_n_spl_0
  );


  buf

  (
    ffc_11_n_spl_000,
    ffc_11_n_spl_00
  );


  buf

  (
    ffc_11_n_spl_001,
    ffc_11_n_spl_00
  );


  buf

  (
    ffc_11_n_spl_01,
    ffc_11_n_spl_0
  );


  buf

  (
    ffc_11_n_spl_010,
    ffc_11_n_spl_01
  );


  buf

  (
    ffc_11_n_spl_011,
    ffc_11_n_spl_01
  );


  buf

  (
    ffc_11_n_spl_1,
    ffc_11_n_spl_
  );


  buf

  (
    ffc_11_n_spl_10,
    ffc_11_n_spl_1
  );


  buf

  (
    ffc_11_n_spl_100,
    ffc_11_n_spl_10
  );


  buf

  (
    ffc_11_n_spl_101,
    ffc_11_n_spl_10
  );


  buf

  (
    ffc_11_n_spl_11,
    ffc_11_n_spl_1
  );


  buf

  (
    g985_p_spl_,
    g985_p
  );


  buf

  (
    g986_p_spl_,
    g986_p
  );


  buf

  (
    g906_p_spl_,
    g906_p
  );


  buf

  (
    ffc_180_p_spl_,
    ffc_180_p
  );


  buf

  (
    ffc_180_p_spl_0,
    ffc_180_p_spl_
  );


  buf

  (
    ffc_180_p_spl_00,
    ffc_180_p_spl_0
  );


  buf

  (
    ffc_180_p_spl_1,
    ffc_180_p_spl_
  );


  buf

  (
    ffc_180_n_spl_,
    ffc_180_n
  );


  buf

  (
    ffc_180_n_spl_0,
    ffc_180_n_spl_
  );


  buf

  (
    ffc_180_n_spl_1,
    ffc_180_n_spl_
  );


  buf

  (
    ffc_327_n_spl_,
    ffc_327_n
  );


  buf

  (
    ffc_344_p_spl_,
    ffc_344_p
  );


  buf

  (
    ffc_327_p_spl_,
    ffc_327_p
  );


  buf

  (
    ffc_344_n_spl_,
    ffc_344_n
  );


  buf

  (
    g995_n_spl_,
    g995_n
  );


  buf

  (
    g995_p_spl_,
    g995_p
  );


  buf

  (
    g994_n_spl_,
    g994_n
  );


  buf

  (
    g997_p_spl_,
    g997_p
  );


  buf

  (
    g994_p_spl_,
    g994_p
  );


  buf

  (
    g997_n_spl_,
    g997_n
  );


  buf

  (
    g998_n_spl_,
    g998_n
  );


  buf

  (
    g998_p_spl_,
    g998_p
  );


  buf

  (
    g993_n_spl_,
    g993_n
  );


  buf

  (
    g1000_p_spl_,
    g1000_p
  );


  buf

  (
    g993_p_spl_,
    g993_p
  );


  buf

  (
    g1000_n_spl_,
    g1000_n
  );


  buf

  (
    g1001_n_spl_,
    g1001_n
  );


  buf

  (
    g1001_p_spl_,
    g1001_p
  );


  buf

  (
    g992_n_spl_,
    g992_n
  );


  buf

  (
    g1003_p_spl_,
    g1003_p
  );


  buf

  (
    g992_p_spl_,
    g992_p
  );


  buf

  (
    g1003_n_spl_,
    g1003_n
  );


  buf

  (
    g1004_n_spl_,
    g1004_n
  );


  buf

  (
    g1004_p_spl_,
    g1004_p
  );


  buf

  (
    g991_n_spl_,
    g991_n
  );


  buf

  (
    g1006_p_spl_,
    g1006_p
  );


  buf

  (
    g991_p_spl_,
    g991_p
  );


  buf

  (
    g1006_n_spl_,
    g1006_n
  );


  buf

  (
    g1007_n_spl_,
    g1007_n
  );


  buf

  (
    g1007_p_spl_,
    g1007_p
  );


  buf

  (
    g990_n_spl_,
    g990_n
  );


  buf

  (
    g1009_p_spl_,
    g1009_p
  );


  buf

  (
    g990_p_spl_,
    g990_p
  );


  buf

  (
    g1009_n_spl_,
    g1009_n
  );


  buf

  (
    g1010_n_spl_,
    g1010_n
  );


  buf

  (
    g1010_p_spl_,
    g1010_p
  );


  buf

  (
    g959_p_spl_,
    g959_p
  );


  buf

  (
    g958_n_spl_,
    g958_n
  );


  buf

  (
    G19_p_spl_,
    G19_p
  );


  buf

  (
    G19_p_spl_0,
    G19_p_spl_
  );


  buf

  (
    G19_p_spl_00,
    G19_p_spl_0
  );


  buf

  (
    G19_p_spl_000,
    G19_p_spl_00
  );


  buf

  (
    G19_p_spl_001,
    G19_p_spl_00
  );


  buf

  (
    G19_p_spl_01,
    G19_p_spl_0
  );


  buf

  (
    G19_p_spl_010,
    G19_p_spl_01
  );


  buf

  (
    G19_p_spl_011,
    G19_p_spl_01
  );


  buf

  (
    G19_p_spl_1,
    G19_p_spl_
  );


  buf

  (
    G19_p_spl_10,
    G19_p_spl_1
  );


  buf

  (
    G19_p_spl_100,
    G19_p_spl_10
  );


  buf

  (
    G19_p_spl_101,
    G19_p_spl_10
  );


  buf

  (
    G19_p_spl_11,
    G19_p_spl_1
  );


  buf

  (
    G19_p_spl_110,
    G19_p_spl_11
  );


  buf

  (
    G19_p_spl_111,
    G19_p_spl_11
  );


  buf

  (
    G19_n_spl_,
    G19_n
  );


  buf

  (
    G19_n_spl_0,
    G19_n_spl_
  );


  buf

  (
    G19_n_spl_00,
    G19_n_spl_0
  );


  buf

  (
    G19_n_spl_000,
    G19_n_spl_00
  );


  buf

  (
    G19_n_spl_001,
    G19_n_spl_00
  );


  buf

  (
    G19_n_spl_01,
    G19_n_spl_0
  );


  buf

  (
    G19_n_spl_010,
    G19_n_spl_01
  );


  buf

  (
    G19_n_spl_011,
    G19_n_spl_01
  );


  buf

  (
    G19_n_spl_1,
    G19_n_spl_
  );


  buf

  (
    G19_n_spl_10,
    G19_n_spl_1
  );


  buf

  (
    G19_n_spl_100,
    G19_n_spl_10
  );


  buf

  (
    G19_n_spl_101,
    G19_n_spl_10
  );


  buf

  (
    G19_n_spl_11,
    G19_n_spl_1
  );


  buf

  (
    G19_n_spl_110,
    G19_n_spl_11
  );


  buf

  (
    G19_n_spl_111,
    G19_n_spl_11
  );


  buf

  (
    ffc_290_n_spl_,
    ffc_290_n
  );


  buf

  (
    ffc_290_p_spl_,
    ffc_290_p
  );


  buf

  (
    ffc_130_p_spl_,
    ffc_130_p
  );


  buf

  (
    ffc_130_p_spl_0,
    ffc_130_p_spl_
  );


  buf

  (
    ffc_130_p_spl_00,
    ffc_130_p_spl_0
  );


  buf

  (
    ffc_130_p_spl_1,
    ffc_130_p_spl_
  );


  buf

  (
    ffc_206_p_spl_,
    ffc_206_p
  );


  buf

  (
    ffc_130_n_spl_,
    ffc_130_n
  );


  buf

  (
    ffc_130_n_spl_0,
    ffc_130_n_spl_
  );


  buf

  (
    ffc_206_n_spl_,
    ffc_206_n
  );


  buf

  (
    ffc_292_p_spl_,
    ffc_292_p
  );


  buf

  (
    ffc_292_n_spl_,
    ffc_292_n
  );


  buf

  (
    g1018_n_spl_,
    g1018_n
  );


  buf

  (
    g1019_p_spl_,
    g1019_p
  );


  buf

  (
    g1018_p_spl_,
    g1018_p
  );


  buf

  (
    g1019_n_spl_,
    g1019_n
  );


  buf

  (
    g1020_n_spl_,
    g1020_n
  );


  buf

  (
    g1020_p_spl_,
    g1020_p
  );


  buf

  (
    g1017_n_spl_,
    g1017_n
  );


  buf

  (
    g1022_p_spl_,
    g1022_p
  );


  buf

  (
    g1017_p_spl_,
    g1017_p
  );


  buf

  (
    g1022_n_spl_,
    g1022_n
  );


  buf

  (
    ffc_129_p_spl_,
    ffc_129_p
  );


  buf

  (
    ffc_129_p_spl_0,
    ffc_129_p_spl_
  );


  buf

  (
    ffc_129_p_spl_1,
    ffc_129_p_spl_
  );


  buf

  (
    ffc_224_p_spl_,
    ffc_224_p
  );


  buf

  (
    ffc_224_p_spl_0,
    ffc_224_p_spl_
  );


  buf

  (
    ffc_224_p_spl_00,
    ffc_224_p_spl_0
  );


  buf

  (
    ffc_224_p_spl_1,
    ffc_224_p_spl_
  );


  buf

  (
    ffc_129_n_spl_,
    ffc_129_n
  );


  buf

  (
    ffc_129_n_spl_0,
    ffc_129_n_spl_
  );


  buf

  (
    ffc_224_n_spl_,
    ffc_224_n
  );


  buf

  (
    ffc_224_n_spl_0,
    ffc_224_n_spl_
  );


  buf

  (
    ffc_224_n_spl_00,
    ffc_224_n_spl_0
  );


  buf

  (
    ffc_224_n_spl_1,
    ffc_224_n_spl_
  );


  buf

  (
    g1023_n_spl_,
    g1023_n
  );


  buf

  (
    g1023_p_spl_,
    g1023_p
  );


  buf

  (
    g1024_n_spl_,
    g1024_n
  );


  buf

  (
    g1026_p_spl_,
    g1026_p
  );


  buf

  (
    g1024_p_spl_,
    g1024_p
  );


  buf

  (
    g1026_n_spl_,
    g1026_n
  );


  buf

  (
    g1027_n_spl_,
    g1027_n
  );


  buf

  (
    g1027_p_spl_,
    g1027_p
  );


  buf

  (
    ffc_131_p_spl_,
    ffc_131_p
  );


  buf

  (
    ffc_131_p_spl_0,
    ffc_131_p_spl_
  );


  buf

  (
    ffc_131_p_spl_1,
    ffc_131_p_spl_
  );


  buf

  (
    ffc_131_n_spl_,
    ffc_131_n
  );


  buf

  (
    ffc_131_n_spl_0,
    ffc_131_n_spl_
  );


  buf

  (
    g1030_n_spl_,
    g1030_n
  );


  buf

  (
    g1031_n_spl_,
    g1031_n
  );


  buf

  (
    g1030_p_spl_,
    g1030_p
  );


  buf

  (
    g1031_p_spl_,
    g1031_p
  );


  buf

  (
    g1032_n_spl_,
    g1032_n
  );


  buf

  (
    g1032_p_spl_,
    g1032_p
  );


  buf

  (
    g1029_n_spl_,
    g1029_n
  );


  buf

  (
    g1034_p_spl_,
    g1034_p
  );


  buf

  (
    g1029_p_spl_,
    g1029_p
  );


  buf

  (
    g1034_n_spl_,
    g1034_n
  );


  buf

  (
    g1035_n_spl_,
    g1035_n
  );


  buf

  (
    g1035_p_spl_,
    g1035_p
  );


  buf

  (
    g1028_n_spl_,
    g1028_n
  );


  buf

  (
    g1037_p_spl_,
    g1037_p
  );


  buf

  (
    g1028_p_spl_,
    g1028_p
  );


  buf

  (
    g1037_n_spl_,
    g1037_n
  );


  buf

  (
    g1038_n_spl_,
    g1038_n
  );


  buf

  (
    g1038_p_spl_,
    g1038_p
  );


  buf

  (
    g1039_n_spl_,
    g1039_n
  );


  buf

  (
    g1041_p_spl_,
    g1041_p
  );


  buf

  (
    g1039_p_spl_,
    g1039_p
  );


  buf

  (
    g1041_n_spl_,
    g1041_n
  );


  buf

  (
    g1042_n_spl_,
    g1042_n
  );


  buf

  (
    g1042_p_spl_,
    g1042_p
  );


  buf

  (
    g1045_n_spl_,
    g1045_n
  );


  buf

  (
    g1046_n_spl_,
    g1046_n
  );


  buf

  (
    g1045_p_spl_,
    g1045_p
  );


  buf

  (
    g1046_p_spl_,
    g1046_p
  );


  buf

  (
    g1047_n_spl_,
    g1047_n
  );


  buf

  (
    g1047_p_spl_,
    g1047_p
  );


  buf

  (
    g1044_n_spl_,
    g1044_n
  );


  buf

  (
    g1049_p_spl_,
    g1049_p
  );


  buf

  (
    g1044_p_spl_,
    g1044_p
  );


  buf

  (
    g1049_n_spl_,
    g1049_n
  );


  buf

  (
    g1050_n_spl_,
    g1050_n
  );


  buf

  (
    g1050_p_spl_,
    g1050_p
  );


  buf

  (
    g1043_n_spl_,
    g1043_n
  );


  buf

  (
    g1052_p_spl_,
    g1052_p
  );


  buf

  (
    g1043_p_spl_,
    g1043_p
  );


  buf

  (
    g1052_n_spl_,
    g1052_n
  );


  buf

  (
    ffc_288_n_spl_,
    ffc_288_n
  );


  buf

  (
    ffc_288_p_spl_,
    ffc_288_p
  );


  buf

  (
    ffc_127_p_spl_,
    ffc_127_p
  );


  buf

  (
    ffc_127_p_spl_0,
    ffc_127_p_spl_
  );


  buf

  (
    ffc_127_p_spl_00,
    ffc_127_p_spl_0
  );


  buf

  (
    ffc_127_p_spl_1,
    ffc_127_p_spl_
  );


  buf

  (
    ffc_127_n_spl_,
    ffc_127_n
  );


  buf

  (
    ffc_127_n_spl_0,
    ffc_127_n_spl_
  );


  buf

  (
    ffc_294_p_spl_,
    ffc_294_p
  );


  buf

  (
    ffc_294_n_spl_,
    ffc_294_n
  );


  buf

  (
    g1055_n_spl_,
    g1055_n
  );


  buf

  (
    g1056_p_spl_,
    g1056_p
  );


  buf

  (
    g1055_p_spl_,
    g1055_p
  );


  buf

  (
    g1056_n_spl_,
    g1056_n
  );


  buf

  (
    g1057_n_spl_,
    g1057_n
  );


  buf

  (
    g1057_p_spl_,
    g1057_p
  );


  buf

  (
    g1054_n_spl_,
    g1054_n
  );


  buf

  (
    g1059_p_spl_,
    g1059_p
  );


  buf

  (
    g1054_p_spl_,
    g1054_p
  );


  buf

  (
    g1059_n_spl_,
    g1059_n
  );


  buf

  (
    ffc_126_p_spl_,
    ffc_126_p
  );


  buf

  (
    ffc_126_p_spl_0,
    ffc_126_p_spl_
  );


  buf

  (
    ffc_126_p_spl_1,
    ffc_126_p_spl_
  );


  buf

  (
    ffc_126_n_spl_,
    ffc_126_n
  );


  buf

  (
    ffc_126_n_spl_0,
    ffc_126_n_spl_
  );


  buf

  (
    g1060_n_spl_,
    g1060_n
  );


  buf

  (
    g1060_p_spl_,
    g1060_p
  );


  buf

  (
    g1061_n_spl_,
    g1061_n
  );


  buf

  (
    g1063_p_spl_,
    g1063_p
  );


  buf

  (
    g1061_p_spl_,
    g1061_p
  );


  buf

  (
    g1063_n_spl_,
    g1063_n
  );


  buf

  (
    g1064_n_spl_,
    g1064_n
  );


  buf

  (
    g1064_p_spl_,
    g1064_p
  );


  buf

  (
    ffc_128_p_spl_,
    ffc_128_p
  );


  buf

  (
    ffc_128_p_spl_0,
    ffc_128_p_spl_
  );


  buf

  (
    ffc_128_p_spl_1,
    ffc_128_p_spl_
  );


  buf

  (
    ffc_128_n_spl_,
    ffc_128_n
  );


  buf

  (
    ffc_128_n_spl_0,
    ffc_128_n_spl_
  );


  buf

  (
    g1069_n_spl_,
    g1069_n
  );


  buf

  (
    g1070_p_spl_,
    g1070_p
  );


  buf

  (
    g1069_p_spl_,
    g1069_p
  );


  buf

  (
    g1070_n_spl_,
    g1070_n
  );


  buf

  (
    g1071_n_spl_,
    g1071_n
  );


  buf

  (
    g1071_p_spl_,
    g1071_p
  );


  buf

  (
    g1068_n_spl_,
    g1068_n
  );


  buf

  (
    g1073_p_spl_,
    g1073_p
  );


  buf

  (
    g1068_p_spl_,
    g1068_p
  );


  buf

  (
    g1073_n_spl_,
    g1073_n
  );


  buf

  (
    g1074_n_spl_,
    g1074_n
  );


  buf

  (
    g1074_p_spl_,
    g1074_p
  );


  buf

  (
    g1067_n_spl_,
    g1067_n
  );


  buf

  (
    g1076_p_spl_,
    g1076_p
  );


  buf

  (
    g1067_p_spl_,
    g1067_p
  );


  buf

  (
    g1076_n_spl_,
    g1076_n
  );


  buf

  (
    g1077_n_spl_,
    g1077_n
  );


  buf

  (
    g1077_p_spl_,
    g1077_p
  );


  buf

  (
    g1066_n_spl_,
    g1066_n
  );


  buf

  (
    g1079_p_spl_,
    g1079_p
  );


  buf

  (
    g1066_p_spl_,
    g1066_p
  );


  buf

  (
    g1079_n_spl_,
    g1079_n
  );


  buf

  (
    g1080_n_spl_,
    g1080_n
  );


  buf

  (
    g1080_p_spl_,
    g1080_p
  );


  buf

  (
    g1065_n_spl_,
    g1065_n
  );


  buf

  (
    g1082_p_spl_,
    g1082_p
  );


  buf

  (
    g1065_p_spl_,
    g1065_p
  );


  buf

  (
    g1082_n_spl_,
    g1082_n
  );


  buf

  (
    g1083_n_spl_,
    g1083_n
  );


  buf

  (
    g1083_p_spl_,
    g1083_p
  );


  buf

  (
    g1084_n_spl_,
    g1084_n
  );


  buf

  (
    g1086_p_spl_,
    g1086_p
  );


  buf

  (
    g1084_p_spl_,
    g1084_p
  );


  buf

  (
    g1086_n_spl_,
    g1086_n
  );


  buf

  (
    g1087_n_spl_,
    g1087_n
  );


  buf

  (
    g1087_p_spl_,
    g1087_p
  );


  buf

  (
    g1092_n_spl_,
    g1092_n
  );


  buf

  (
    g1094_p_spl_,
    g1094_p
  );


  buf

  (
    g1092_p_spl_,
    g1092_p
  );


  buf

  (
    g1094_n_spl_,
    g1094_n
  );


  buf

  (
    g1095_n_spl_,
    g1095_n
  );


  buf

  (
    g1095_p_spl_,
    g1095_p
  );


  buf

  (
    g1091_n_spl_,
    g1091_n
  );


  buf

  (
    g1097_p_spl_,
    g1097_p
  );


  buf

  (
    g1091_p_spl_,
    g1091_p
  );


  buf

  (
    g1097_n_spl_,
    g1097_n
  );


  buf

  (
    g1098_n_spl_,
    g1098_n
  );


  buf

  (
    g1098_p_spl_,
    g1098_p
  );


  buf

  (
    g1090_n_spl_,
    g1090_n
  );


  buf

  (
    g1100_p_spl_,
    g1100_p
  );


  buf

  (
    g1090_p_spl_,
    g1090_p
  );


  buf

  (
    g1100_n_spl_,
    g1100_n
  );


  buf

  (
    g1101_n_spl_,
    g1101_n
  );


  buf

  (
    g1101_p_spl_,
    g1101_p
  );


  buf

  (
    g1089_n_spl_,
    g1089_n
  );


  buf

  (
    g1103_p_spl_,
    g1103_p
  );


  buf

  (
    g1089_p_spl_,
    g1089_p
  );


  buf

  (
    g1103_n_spl_,
    g1103_n
  );


  buf

  (
    g1104_n_spl_,
    g1104_n
  );


  buf

  (
    g1104_p_spl_,
    g1104_p
  );


  buf

  (
    g1088_n_spl_,
    g1088_n
  );


  buf

  (
    g1106_p_spl_,
    g1106_p
  );


  buf

  (
    g1088_p_spl_,
    g1088_p
  );


  buf

  (
    g1106_n_spl_,
    g1106_n
  );


  buf

  (
    ffc_123_p_spl_,
    ffc_123_p
  );


  buf

  (
    ffc_123_p_spl_0,
    ffc_123_p_spl_
  );


  buf

  (
    ffc_123_p_spl_00,
    ffc_123_p_spl_0
  );


  buf

  (
    ffc_123_p_spl_1,
    ffc_123_p_spl_
  );


  buf

  (
    ffc_123_n_spl_,
    ffc_123_n
  );


  buf

  (
    ffc_123_n_spl_0,
    ffc_123_n_spl_
  );


  buf

  (
    ffc_123_n_spl_1,
    ffc_123_n_spl_
  );


  buf

  (
    ffc_306_p_spl_,
    ffc_306_p
  );


  buf

  (
    ffc_306_n_spl_,
    ffc_306_n
  );


  buf

  (
    g1108_n_spl_,
    g1108_n
  );


  buf

  (
    g1109_p_spl_,
    g1109_p
  );


  buf

  (
    g1108_p_spl_,
    g1108_p
  );


  buf

  (
    g1109_n_spl_,
    g1109_n
  );


  buf

  (
    g1110_n_spl_,
    g1110_n
  );


  buf

  (
    g1110_p_spl_,
    g1110_p
  );


  buf

  (
    ffc_124_p_spl_,
    ffc_124_p
  );


  buf

  (
    ffc_124_p_spl_0,
    ffc_124_p_spl_
  );


  buf

  (
    ffc_124_p_spl_00,
    ffc_124_p_spl_0
  );


  buf

  (
    ffc_124_p_spl_1,
    ffc_124_p_spl_
  );


  buf

  (
    ffc_124_n_spl_,
    ffc_124_n
  );


  buf

  (
    ffc_124_n_spl_0,
    ffc_124_n_spl_
  );


  buf

  (
    ffc_308_p_spl_,
    ffc_308_p
  );


  buf

  (
    ffc_308_n_spl_,
    ffc_308_n
  );


  buf

  (
    g1112_n_spl_,
    g1112_n
  );


  buf

  (
    g1113_p_spl_,
    g1113_p
  );


  buf

  (
    g1112_p_spl_,
    g1112_p
  );


  buf

  (
    g1113_n_spl_,
    g1113_n
  );


  buf

  (
    g1114_n_spl_,
    g1114_n
  );


  buf

  (
    g1114_p_spl_,
    g1114_p
  );


  buf

  (
    g1111_n_spl_,
    g1111_n
  );


  buf

  (
    g1116_p_spl_,
    g1116_p
  );


  buf

  (
    g1111_p_spl_,
    g1111_p
  );


  buf

  (
    g1116_n_spl_,
    g1116_n
  );


  buf

  (
    g1117_n_spl_,
    g1117_n
  );


  buf

  (
    g1117_p_spl_,
    g1117_p
  );


  buf

  (
    g1118_n_spl_,
    g1118_n
  );


  buf

  (
    g1120_p_spl_,
    g1120_p
  );


  buf

  (
    g1118_p_spl_,
    g1118_p
  );


  buf

  (
    g1120_n_spl_,
    g1120_n
  );


  buf

  (
    g1121_n_spl_,
    g1121_n
  );


  buf

  (
    g1121_p_spl_,
    g1121_p
  );


  buf

  (
    ffc_125_p_spl_,
    ffc_125_p
  );


  buf

  (
    ffc_125_p_spl_0,
    ffc_125_p_spl_
  );


  buf

  (
    ffc_125_p_spl_1,
    ffc_125_p_spl_
  );


  buf

  (
    ffc_125_n_spl_,
    ffc_125_n
  );


  buf

  (
    ffc_125_n_spl_0,
    ffc_125_n_spl_
  );


  buf

  (
    g1126_n_spl_,
    g1126_n
  );


  buf

  (
    g1127_p_spl_,
    g1127_p
  );


  buf

  (
    g1126_p_spl_,
    g1126_p
  );


  buf

  (
    g1127_n_spl_,
    g1127_n
  );


  buf

  (
    g1128_n_spl_,
    g1128_n
  );


  buf

  (
    g1128_p_spl_,
    g1128_p
  );


  buf

  (
    g1125_n_spl_,
    g1125_n
  );


  buf

  (
    g1130_p_spl_,
    g1130_p
  );


  buf

  (
    g1125_p_spl_,
    g1125_p
  );


  buf

  (
    g1130_n_spl_,
    g1130_n
  );


  buf

  (
    g1131_n_spl_,
    g1131_n
  );


  buf

  (
    g1131_p_spl_,
    g1131_p
  );


  buf

  (
    g1124_n_spl_,
    g1124_n
  );


  buf

  (
    g1133_p_spl_,
    g1133_p
  );


  buf

  (
    g1124_p_spl_,
    g1124_p
  );


  buf

  (
    g1133_n_spl_,
    g1133_n
  );


  buf

  (
    g1134_n_spl_,
    g1134_n
  );


  buf

  (
    g1134_p_spl_,
    g1134_p
  );


  buf

  (
    g1123_n_spl_,
    g1123_n
  );


  buf

  (
    g1136_p_spl_,
    g1136_p
  );


  buf

  (
    g1123_p_spl_,
    g1123_p
  );


  buf

  (
    g1136_n_spl_,
    g1136_n
  );


  buf

  (
    g1137_n_spl_,
    g1137_n
  );


  buf

  (
    g1137_p_spl_,
    g1137_p
  );


  buf

  (
    g1122_n_spl_,
    g1122_n
  );


  buf

  (
    g1139_p_spl_,
    g1139_p
  );


  buf

  (
    g1122_p_spl_,
    g1122_p
  );


  buf

  (
    g1139_n_spl_,
    g1139_n
  );


  buf

  (
    g1140_n_spl_,
    g1140_n
  );


  buf

  (
    g1140_p_spl_,
    g1140_p
  );


  buf

  (
    g1141_n_spl_,
    g1141_n
  );


  buf

  (
    g1143_p_spl_,
    g1143_p
  );


  buf

  (
    g1141_p_spl_,
    g1141_p
  );


  buf

  (
    g1143_n_spl_,
    g1143_n
  );


  buf

  (
    g1144_n_spl_,
    g1144_n
  );


  buf

  (
    g1144_p_spl_,
    g1144_p
  );


  buf

  (
    g1149_n_spl_,
    g1149_n
  );


  buf

  (
    g1151_p_spl_,
    g1151_p
  );


  buf

  (
    g1149_p_spl_,
    g1149_p
  );


  buf

  (
    g1151_n_spl_,
    g1151_n
  );


  buf

  (
    g1152_n_spl_,
    g1152_n
  );


  buf

  (
    g1152_p_spl_,
    g1152_p
  );


  buf

  (
    g1148_n_spl_,
    g1148_n
  );


  buf

  (
    g1154_p_spl_,
    g1154_p
  );


  buf

  (
    g1148_p_spl_,
    g1148_p
  );


  buf

  (
    g1154_n_spl_,
    g1154_n
  );


  buf

  (
    g1155_n_spl_,
    g1155_n
  );


  buf

  (
    g1155_p_spl_,
    g1155_p
  );


  buf

  (
    g1147_n_spl_,
    g1147_n
  );


  buf

  (
    g1157_p_spl_,
    g1157_p
  );


  buf

  (
    g1147_p_spl_,
    g1147_p
  );


  buf

  (
    g1157_n_spl_,
    g1157_n
  );


  buf

  (
    g1158_n_spl_,
    g1158_n
  );


  buf

  (
    g1158_p_spl_,
    g1158_p
  );


  buf

  (
    g1146_n_spl_,
    g1146_n
  );


  buf

  (
    g1160_p_spl_,
    g1160_p
  );


  buf

  (
    g1146_p_spl_,
    g1146_p
  );


  buf

  (
    g1160_n_spl_,
    g1160_n
  );


  buf

  (
    g1161_n_spl_,
    g1161_n
  );


  buf

  (
    g1161_p_spl_,
    g1161_p
  );


  buf

  (
    g1145_n_spl_,
    g1145_n
  );


  buf

  (
    g1163_p_spl_,
    g1163_p
  );


  buf

  (
    g1145_p_spl_,
    g1145_p
  );


  buf

  (
    g1163_n_spl_,
    g1163_n
  );


  buf

  (
    ffc_120_p_spl_,
    ffc_120_p
  );


  buf

  (
    ffc_120_p_spl_0,
    ffc_120_p_spl_
  );


  buf

  (
    ffc_120_p_spl_00,
    ffc_120_p_spl_0
  );


  buf

  (
    ffc_120_p_spl_01,
    ffc_120_p_spl_0
  );


  buf

  (
    ffc_120_p_spl_1,
    ffc_120_p_spl_
  );


  buf

  (
    ffc_120_n_spl_,
    ffc_120_n
  );


  buf

  (
    ffc_120_n_spl_0,
    ffc_120_n_spl_
  );


  buf

  (
    ffc_120_n_spl_00,
    ffc_120_n_spl_0
  );


  buf

  (
    ffc_120_n_spl_1,
    ffc_120_n_spl_
  );


  buf

  (
    ffc_300_p_spl_,
    ffc_300_p
  );


  buf

  (
    ffc_300_n_spl_,
    ffc_300_n
  );


  buf

  (
    g1165_n_spl_,
    g1165_n
  );


  buf

  (
    g1166_p_spl_,
    g1166_p
  );


  buf

  (
    g1165_p_spl_,
    g1165_p
  );


  buf

  (
    g1166_n_spl_,
    g1166_n
  );


  buf

  (
    g1167_n_spl_,
    g1167_n
  );


  buf

  (
    g1167_p_spl_,
    g1167_p
  );


  buf

  (
    ffc_121_p_spl_,
    ffc_121_p
  );


  buf

  (
    ffc_121_p_spl_0,
    ffc_121_p_spl_
  );


  buf

  (
    ffc_121_p_spl_00,
    ffc_121_p_spl_0
  );


  buf

  (
    ffc_121_p_spl_01,
    ffc_121_p_spl_0
  );


  buf

  (
    ffc_121_p_spl_1,
    ffc_121_p_spl_
  );


  buf

  (
    ffc_121_n_spl_,
    ffc_121_n
  );


  buf

  (
    ffc_121_n_spl_0,
    ffc_121_n_spl_
  );


  buf

  (
    ffc_121_n_spl_1,
    ffc_121_n_spl_
  );


  buf

  (
    ffc_302_p_spl_,
    ffc_302_p
  );


  buf

  (
    ffc_302_n_spl_,
    ffc_302_n
  );


  buf

  (
    g1169_n_spl_,
    g1169_n
  );


  buf

  (
    g1170_p_spl_,
    g1170_p
  );


  buf

  (
    g1169_p_spl_,
    g1169_p
  );


  buf

  (
    g1170_n_spl_,
    g1170_n
  );


  buf

  (
    g1171_n_spl_,
    g1171_n
  );


  buf

  (
    g1171_p_spl_,
    g1171_p
  );


  buf

  (
    g1168_n_spl_,
    g1168_n
  );


  buf

  (
    g1173_p_spl_,
    g1173_p
  );


  buf

  (
    g1168_p_spl_,
    g1168_p
  );


  buf

  (
    g1173_n_spl_,
    g1173_n
  );


  buf

  (
    g1174_n_spl_,
    g1174_n
  );


  buf

  (
    g1174_p_spl_,
    g1174_p
  );


  buf

  (
    g1175_n_spl_,
    g1175_n
  );


  buf

  (
    g1177_p_spl_,
    g1177_p
  );


  buf

  (
    g1175_p_spl_,
    g1175_p
  );


  buf

  (
    g1177_n_spl_,
    g1177_n
  );


  buf

  (
    g1178_n_spl_,
    g1178_n
  );


  buf

  (
    g1178_p_spl_,
    g1178_p
  );


  buf

  (
    ffc_122_p_spl_,
    ffc_122_p
  );


  buf

  (
    ffc_122_p_spl_0,
    ffc_122_p_spl_
  );


  buf

  (
    ffc_122_p_spl_00,
    ffc_122_p_spl_0
  );


  buf

  (
    ffc_122_p_spl_1,
    ffc_122_p_spl_
  );


  buf

  (
    ffc_122_n_spl_,
    ffc_122_n
  );


  buf

  (
    ffc_122_n_spl_0,
    ffc_122_n_spl_
  );


  buf

  (
    ffc_122_n_spl_1,
    ffc_122_n_spl_
  );


  buf

  (
    ffc_304_p_spl_,
    ffc_304_p
  );


  buf

  (
    ffc_304_n_spl_,
    ffc_304_n
  );


  buf

  (
    g1182_n_spl_,
    g1182_n
  );


  buf

  (
    g1183_p_spl_,
    g1183_p
  );


  buf

  (
    g1182_p_spl_,
    g1182_p
  );


  buf

  (
    g1183_n_spl_,
    g1183_n
  );


  buf

  (
    g1184_n_spl_,
    g1184_n
  );


  buf

  (
    g1184_p_spl_,
    g1184_p
  );


  buf

  (
    g1181_n_spl_,
    g1181_n
  );


  buf

  (
    g1186_p_spl_,
    g1186_p
  );


  buf

  (
    g1181_p_spl_,
    g1181_p
  );


  buf

  (
    g1186_n_spl_,
    g1186_n
  );


  buf

  (
    g1187_n_spl_,
    g1187_n
  );


  buf

  (
    g1187_p_spl_,
    g1187_p
  );


  buf

  (
    g1180_n_spl_,
    g1180_n
  );


  buf

  (
    g1189_p_spl_,
    g1189_p
  );


  buf

  (
    g1180_p_spl_,
    g1180_p
  );


  buf

  (
    g1189_n_spl_,
    g1189_n
  );


  buf

  (
    g1190_n_spl_,
    g1190_n
  );


  buf

  (
    g1190_p_spl_,
    g1190_p
  );


  buf

  (
    g1179_n_spl_,
    g1179_n
  );


  buf

  (
    g1192_p_spl_,
    g1192_p
  );


  buf

  (
    g1179_p_spl_,
    g1179_p
  );


  buf

  (
    g1192_n_spl_,
    g1192_n
  );


  buf

  (
    g1193_n_spl_,
    g1193_n
  );


  buf

  (
    g1193_p_spl_,
    g1193_p
  );


  buf

  (
    g1194_n_spl_,
    g1194_n
  );


  buf

  (
    g1196_p_spl_,
    g1196_p
  );


  buf

  (
    g1194_p_spl_,
    g1194_p
  );


  buf

  (
    g1196_n_spl_,
    g1196_n
  );


  buf

  (
    g1197_n_spl_,
    g1197_n
  );


  buf

  (
    g1197_p_spl_,
    g1197_p
  );


  buf

  (
    g1202_n_spl_,
    g1202_n
  );


  buf

  (
    g1204_p_spl_,
    g1204_p
  );


  buf

  (
    g1202_p_spl_,
    g1202_p
  );


  buf

  (
    g1204_n_spl_,
    g1204_n
  );


  buf

  (
    g1205_n_spl_,
    g1205_n
  );


  buf

  (
    g1205_p_spl_,
    g1205_p
  );


  buf

  (
    g1201_n_spl_,
    g1201_n
  );


  buf

  (
    g1207_p_spl_,
    g1207_p
  );


  buf

  (
    g1201_p_spl_,
    g1201_p
  );


  buf

  (
    g1207_n_spl_,
    g1207_n
  );


  buf

  (
    g1208_n_spl_,
    g1208_n
  );


  buf

  (
    g1208_p_spl_,
    g1208_p
  );


  buf

  (
    g1200_n_spl_,
    g1200_n
  );


  buf

  (
    g1210_p_spl_,
    g1210_p
  );


  buf

  (
    g1200_p_spl_,
    g1200_p
  );


  buf

  (
    g1210_n_spl_,
    g1210_n
  );


  buf

  (
    g1211_n_spl_,
    g1211_n
  );


  buf

  (
    g1211_p_spl_,
    g1211_p
  );


  buf

  (
    g1199_n_spl_,
    g1199_n
  );


  buf

  (
    g1213_p_spl_,
    g1213_p
  );


  buf

  (
    g1199_p_spl_,
    g1199_p
  );


  buf

  (
    g1213_n_spl_,
    g1213_n
  );


  buf

  (
    g1214_n_spl_,
    g1214_n
  );


  buf

  (
    g1214_p_spl_,
    g1214_p
  );


  buf

  (
    g1198_n_spl_,
    g1198_n
  );


  buf

  (
    g1216_p_spl_,
    g1216_p
  );


  buf

  (
    g1198_p_spl_,
    g1198_p
  );


  buf

  (
    g1216_n_spl_,
    g1216_n
  );


  buf

  (
    g1217_n_spl_,
    g1217_n
  );


  buf

  (
    g1217_p_spl_,
    g1217_p
  );


  buf

  (
    g1218_n_spl_,
    g1218_n
  );


  buf

  (
    g1220_p_spl_,
    g1220_p
  );


  buf

  (
    g1218_p_spl_,
    g1218_p
  );


  buf

  (
    g1220_n_spl_,
    g1220_n
  );


  buf

  (
    g1221_n_spl_,
    g1221_n
  );


  buf

  (
    g1221_p_spl_,
    g1221_p
  );


  buf

  (
    g1226_n_spl_,
    g1226_n
  );


  buf

  (
    g1228_p_spl_,
    g1228_p
  );


  buf

  (
    g1226_p_spl_,
    g1226_p
  );


  buf

  (
    g1228_n_spl_,
    g1228_n
  );


  buf

  (
    g1229_n_spl_,
    g1229_n
  );


  buf

  (
    g1229_p_spl_,
    g1229_p
  );


  buf

  (
    g1225_n_spl_,
    g1225_n
  );


  buf

  (
    g1231_p_spl_,
    g1231_p
  );


  buf

  (
    g1225_p_spl_,
    g1225_p
  );


  buf

  (
    g1231_n_spl_,
    g1231_n
  );


  buf

  (
    g1232_n_spl_,
    g1232_n
  );


  buf

  (
    g1232_p_spl_,
    g1232_p
  );


  buf

  (
    g1224_n_spl_,
    g1224_n
  );


  buf

  (
    g1234_p_spl_,
    g1234_p
  );


  buf

  (
    g1224_p_spl_,
    g1224_p
  );


  buf

  (
    g1234_n_spl_,
    g1234_n
  );


  buf

  (
    g1235_n_spl_,
    g1235_n
  );


  buf

  (
    g1235_p_spl_,
    g1235_p
  );


  buf

  (
    g1223_n_spl_,
    g1223_n
  );


  buf

  (
    g1237_p_spl_,
    g1237_p
  );


  buf

  (
    g1223_p_spl_,
    g1223_p
  );


  buf

  (
    g1237_n_spl_,
    g1237_n
  );


  buf

  (
    g1238_n_spl_,
    g1238_n
  );


  buf

  (
    g1238_p_spl_,
    g1238_p
  );


  buf

  (
    g1222_n_spl_,
    g1222_n
  );


  buf

  (
    g1240_p_spl_,
    g1240_p
  );


  buf

  (
    g1222_p_spl_,
    g1222_p
  );


  buf

  (
    g1240_n_spl_,
    g1240_n
  );


  buf

  (
    g1012_p_spl_,
    g1012_p
  );


  buf

  (
    g988_p_spl_,
    g988_p
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G3_p_spl_0,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_00,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_01,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_1,
    G3_p_spl_
  );


  buf

  (
    G3_n_spl_,
    G3_n
  );


  buf

  (
    G3_n_spl_0,
    G3_n_spl_
  );


  buf

  (
    G3_n_spl_1,
    G3_n_spl_
  );


  buf

  (
    g1243_p_spl_,
    g1243_p
  );


  buf

  (
    g1244_p_spl_,
    g1244_p
  );


  buf

  (
    g1243_n_spl_,
    g1243_n
  );


  buf

  (
    g1244_n_spl_,
    g1244_n
  );


  buf

  (
    g1245_n_spl_,
    g1245_n
  );


  buf

  (
    g1245_n_spl_0,
    g1245_n_spl_
  );


  buf

  (
    g1245_p_spl_,
    g1245_p
  );


  buf

  (
    g1245_p_spl_0,
    g1245_p_spl_
  );


  buf

  (
    g989_n_spl_,
    g989_n
  );


  buf

  (
    g1247_n_spl_,
    g1247_n
  );


  buf

  (
    g989_p_spl_,
    g989_p
  );


  buf

  (
    g989_p_spl_0,
    g989_p_spl_
  );


  buf

  (
    g1247_p_spl_,
    g1247_p
  );


  buf

  (
    g1248_n_spl_,
    g1248_n
  );


  buf

  (
    g1248_p_spl_,
    g1248_p
  );


  buf

  (
    g987_p_spl_,
    g987_p
  );


  buf

  (
    g1257_n_spl_,
    g1257_n
  );


  buf

  (
    g1259_p_spl_,
    g1259_p
  );


  buf

  (
    g1257_p_spl_,
    g1257_p
  );


  buf

  (
    g1259_n_spl_,
    g1259_n
  );


  buf

  (
    g1260_n_spl_,
    g1260_n
  );


  buf

  (
    g1260_p_spl_,
    g1260_p
  );


  buf

  (
    g1256_n_spl_,
    g1256_n
  );


  buf

  (
    g1262_p_spl_,
    g1262_p
  );


  buf

  (
    g1256_p_spl_,
    g1256_p
  );


  buf

  (
    g1262_n_spl_,
    g1262_n
  );


  buf

  (
    g1263_n_spl_,
    g1263_n
  );


  buf

  (
    g1263_p_spl_,
    g1263_p
  );


  buf

  (
    g1255_n_spl_,
    g1255_n
  );


  buf

  (
    g1265_p_spl_,
    g1265_p
  );


  buf

  (
    g1255_p_spl_,
    g1255_p
  );


  buf

  (
    g1265_n_spl_,
    g1265_n
  );


  buf

  (
    g1266_n_spl_,
    g1266_n
  );


  buf

  (
    g1266_p_spl_,
    g1266_p
  );


  buf

  (
    g1254_n_spl_,
    g1254_n
  );


  buf

  (
    g1268_p_spl_,
    g1268_p
  );


  buf

  (
    g1254_p_spl_,
    g1254_p
  );


  buf

  (
    g1268_n_spl_,
    g1268_n
  );


  buf

  (
    g1269_n_spl_,
    g1269_n
  );


  buf

  (
    g1269_p_spl_,
    g1269_p
  );


  buf

  (
    g1253_n_spl_,
    g1253_n
  );


  buf

  (
    g1271_p_spl_,
    g1271_p
  );


  buf

  (
    g1253_p_spl_,
    g1253_p
  );


  buf

  (
    g1271_n_spl_,
    g1271_n
  );


  buf

  (
    g1272_n_spl_,
    g1272_n
  );


  buf

  (
    g1272_p_spl_,
    g1272_p
  );


  buf

  (
    g1252_n_spl_,
    g1252_n
  );


  buf

  (
    g1274_p_spl_,
    g1274_p
  );


  buf

  (
    g1252_p_spl_,
    g1252_p
  );


  buf

  (
    g1274_n_spl_,
    g1274_n
  );


  buf

  (
    g1275_n_spl_,
    g1275_n
  );


  buf

  (
    g1275_p_spl_,
    g1275_p
  );


  buf

  (
    ffc_336_n_spl_,
    ffc_336_n
  );


  buf

  (
    ffc_353_p_spl_,
    ffc_353_p
  );


  buf

  (
    ffc_336_p_spl_,
    ffc_336_p
  );


  buf

  (
    ffc_353_n_spl_,
    ffc_353_n
  );


  buf

  (
    g1279_n_spl_,
    g1279_n
  );


  buf

  (
    g1279_p_spl_,
    g1279_p
  );


  buf

  (
    ffc_337_n_spl_,
    ffc_337_n
  );


  buf

  (
    ffc_354_p_spl_,
    ffc_354_p
  );


  buf

  (
    ffc_337_p_spl_,
    ffc_337_p
  );


  buf

  (
    ffc_354_n_spl_,
    ffc_354_n
  );


  buf

  (
    g1281_n_spl_,
    g1281_n
  );


  buf

  (
    g1281_p_spl_,
    g1281_p
  );


  buf

  (
    g1280_n_spl_,
    g1280_n
  );


  buf

  (
    g1283_p_spl_,
    g1283_p
  );


  buf

  (
    g1280_p_spl_,
    g1280_p
  );


  buf

  (
    g1283_n_spl_,
    g1283_n
  );


  buf

  (
    ffc_190_p_spl_,
    ffc_190_p
  );


  buf

  (
    ffc_190_p_spl_0,
    ffc_190_p_spl_
  );


  buf

  (
    ffc_190_p_spl_1,
    ffc_190_p_spl_
  );


  buf

  (
    ffc_190_n_spl_,
    ffc_190_n
  );


  buf

  (
    ffc_190_n_spl_0,
    ffc_190_n_spl_
  );


  buf

  (
    g1284_n_spl_,
    g1284_n
  );


  buf

  (
    g1284_p_spl_,
    g1284_p
  );


  buf

  (
    g1285_n_spl_,
    g1285_n
  );


  buf

  (
    g1287_p_spl_,
    g1287_p
  );


  buf

  (
    g1285_p_spl_,
    g1285_p
  );


  buf

  (
    g1287_n_spl_,
    g1287_n
  );


  buf

  (
    g1288_n_spl_,
    g1288_n
  );


  buf

  (
    g1288_p_spl_,
    g1288_p
  );


  buf

  (
    ffc_191_p_spl_,
    ffc_191_p
  );


  buf

  (
    ffc_191_p_spl_0,
    ffc_191_p_spl_
  );


  buf

  (
    ffc_191_n_spl_,
    ffc_191_n
  );


  buf

  (
    ffc_191_n_spl_0,
    ffc_191_n_spl_
  );


  buf

  (
    ffc_192_p_spl_,
    ffc_192_p
  );


  buf

  (
    ffc_192_p_spl_0,
    ffc_192_p_spl_
  );


  buf

  (
    ffc_192_p_spl_1,
    ffc_192_p_spl_
  );


  buf

  (
    ffc_192_n_spl_,
    ffc_192_n
  );


  buf

  (
    ffc_192_n_spl_0,
    ffc_192_n_spl_
  );


  buf

  (
    ffc_338_n_spl_,
    ffc_338_n
  );


  buf

  (
    ffc_340_n_spl_,
    ffc_340_n
  );


  buf

  (
    ffc_338_p_spl_,
    ffc_338_p
  );


  buf

  (
    ffc_340_p_spl_,
    ffc_340_p
  );


  buf

  (
    g1293_n_spl_,
    g1293_n
  );


  buf

  (
    g1293_p_spl_,
    g1293_p
  );


  buf

  (
    g1292_n_spl_,
    g1292_n
  );


  buf

  (
    g1295_p_spl_,
    g1295_p
  );


  buf

  (
    g1292_p_spl_,
    g1292_p
  );


  buf

  (
    g1295_n_spl_,
    g1295_n
  );


  buf

  (
    g1296_n_spl_,
    g1296_n
  );


  buf

  (
    g1296_p_spl_,
    g1296_p
  );


  buf

  (
    g1291_n_spl_,
    g1291_n
  );


  buf

  (
    g1298_p_spl_,
    g1298_p
  );


  buf

  (
    g1291_p_spl_,
    g1291_p
  );


  buf

  (
    g1298_n_spl_,
    g1298_n
  );


  buf

  (
    g1299_n_spl_,
    g1299_n
  );


  buf

  (
    g1299_p_spl_,
    g1299_p
  );


  buf

  (
    g1290_n_spl_,
    g1290_n
  );


  buf

  (
    g1301_p_spl_,
    g1301_p
  );


  buf

  (
    g1290_p_spl_,
    g1290_p
  );


  buf

  (
    g1301_n_spl_,
    g1301_n
  );


  buf

  (
    g1302_n_spl_,
    g1302_n
  );


  buf

  (
    g1302_p_spl_,
    g1302_p
  );


  buf

  (
    g1289_n_spl_,
    g1289_n
  );


  buf

  (
    g1304_p_spl_,
    g1304_p
  );


  buf

  (
    g1289_p_spl_,
    g1289_p
  );


  buf

  (
    g1304_n_spl_,
    g1304_n
  );


  buf

  (
    g1305_n_spl_,
    g1305_n
  );


  buf

  (
    g1305_p_spl_,
    g1305_p
  );


  buf

  (
    g1306_n_spl_,
    g1306_n
  );


  buf

  (
    g1308_p_spl_,
    g1308_p
  );


  buf

  (
    g1306_p_spl_,
    g1306_p
  );


  buf

  (
    g1308_n_spl_,
    g1308_n
  );


  buf

  (
    g1309_n_spl_,
    g1309_n
  );


  buf

  (
    g1309_p_spl_,
    g1309_p
  );


  buf

  (
    ffc_193_p_spl_,
    ffc_193_p
  );


  buf

  (
    ffc_193_p_spl_0,
    ffc_193_p_spl_
  );


  buf

  (
    ffc_193_n_spl_,
    ffc_193_n
  );


  buf

  (
    ffc_193_n_spl_0,
    ffc_193_n_spl_
  );


  buf

  (
    g1314_n_spl_,
    g1314_n
  );


  buf

  (
    g1315_n_spl_,
    g1315_n
  );


  buf

  (
    g1314_p_spl_,
    g1314_p
  );


  buf

  (
    g1315_p_spl_,
    g1315_p
  );


  buf

  (
    g1316_n_spl_,
    g1316_n
  );


  buf

  (
    g1316_p_spl_,
    g1316_p
  );


  buf

  (
    g1313_n_spl_,
    g1313_n
  );


  buf

  (
    g1318_p_spl_,
    g1318_p
  );


  buf

  (
    g1313_p_spl_,
    g1313_p
  );


  buf

  (
    g1318_n_spl_,
    g1318_n
  );


  buf

  (
    g1319_n_spl_,
    g1319_n
  );


  buf

  (
    g1319_p_spl_,
    g1319_p
  );


  buf

  (
    g1312_n_spl_,
    g1312_n
  );


  buf

  (
    g1321_p_spl_,
    g1321_p
  );


  buf

  (
    g1312_p_spl_,
    g1312_p
  );


  buf

  (
    g1321_n_spl_,
    g1321_n
  );


  buf

  (
    g1322_n_spl_,
    g1322_n
  );


  buf

  (
    g1322_p_spl_,
    g1322_p
  );


  buf

  (
    g1311_n_spl_,
    g1311_n
  );


  buf

  (
    g1324_p_spl_,
    g1324_p
  );


  buf

  (
    g1311_p_spl_,
    g1311_p
  );


  buf

  (
    g1324_n_spl_,
    g1324_n
  );


  buf

  (
    g1325_n_spl_,
    g1325_n
  );


  buf

  (
    g1325_p_spl_,
    g1325_p
  );


  buf

  (
    g1310_n_spl_,
    g1310_n
  );


  buf

  (
    g1327_p_spl_,
    g1327_p
  );


  buf

  (
    g1310_p_spl_,
    g1310_p
  );


  buf

  (
    g1327_n_spl_,
    g1327_n
  );


  buf

  (
    ffc_333_n_spl_,
    ffc_333_n
  );


  buf

  (
    ffc_350_p_spl_,
    ffc_350_p
  );


  buf

  (
    ffc_333_p_spl_,
    ffc_333_p
  );


  buf

  (
    ffc_350_n_spl_,
    ffc_350_n
  );


  buf

  (
    g1329_n_spl_,
    g1329_n
  );


  buf

  (
    g1329_p_spl_,
    g1329_p
  );


  buf

  (
    ffc_334_n_spl_,
    ffc_334_n
  );


  buf

  (
    ffc_351_p_spl_,
    ffc_351_p
  );


  buf

  (
    ffc_334_p_spl_,
    ffc_334_p
  );


  buf

  (
    ffc_351_n_spl_,
    ffc_351_n
  );


  buf

  (
    g1331_n_spl_,
    g1331_n
  );


  buf

  (
    g1331_p_spl_,
    g1331_p
  );


  buf

  (
    g1330_n_spl_,
    g1330_n
  );


  buf

  (
    g1333_p_spl_,
    g1333_p
  );


  buf

  (
    g1330_p_spl_,
    g1330_p
  );


  buf

  (
    g1333_n_spl_,
    g1333_n
  );


  buf

  (
    ffc_187_p_spl_,
    ffc_187_p
  );


  buf

  (
    ffc_187_p_spl_0,
    ffc_187_p_spl_
  );


  buf

  (
    ffc_187_p_spl_00,
    ffc_187_p_spl_0
  );


  buf

  (
    ffc_187_p_spl_1,
    ffc_187_p_spl_
  );


  buf

  (
    ffc_187_n_spl_,
    ffc_187_n
  );


  buf

  (
    ffc_187_n_spl_0,
    ffc_187_n_spl_
  );


  buf

  (
    ffc_187_n_spl_1,
    ffc_187_n_spl_
  );


  buf

  (
    g1334_n_spl_,
    g1334_n
  );


  buf

  (
    g1334_p_spl_,
    g1334_p
  );


  buf

  (
    g1335_n_spl_,
    g1335_n
  );


  buf

  (
    g1337_p_spl_,
    g1337_p
  );


  buf

  (
    g1335_p_spl_,
    g1335_p
  );


  buf

  (
    g1337_n_spl_,
    g1337_n
  );


  buf

  (
    g1338_n_spl_,
    g1338_n
  );


  buf

  (
    g1338_p_spl_,
    g1338_p
  );


  buf

  (
    ffc_188_p_spl_,
    ffc_188_p
  );


  buf

  (
    ffc_188_p_spl_0,
    ffc_188_p_spl_
  );


  buf

  (
    ffc_188_p_spl_1,
    ffc_188_p_spl_
  );


  buf

  (
    ffc_188_n_spl_,
    ffc_188_n
  );


  buf

  (
    ffc_188_n_spl_0,
    ffc_188_n_spl_
  );


  buf

  (
    ffc_188_n_spl_1,
    ffc_188_n_spl_
  );


  buf

  (
    ffc_335_n_spl_,
    ffc_335_n
  );


  buf

  (
    ffc_352_p_spl_,
    ffc_352_p
  );


  buf

  (
    ffc_335_p_spl_,
    ffc_335_p
  );


  buf

  (
    ffc_352_n_spl_,
    ffc_352_n
  );


  buf

  (
    g1342_n_spl_,
    g1342_n
  );


  buf

  (
    g1342_p_spl_,
    g1342_p
  );


  buf

  (
    g1341_n_spl_,
    g1341_n
  );


  buf

  (
    g1344_p_spl_,
    g1344_p
  );


  buf

  (
    g1341_p_spl_,
    g1341_p
  );


  buf

  (
    g1344_n_spl_,
    g1344_n
  );


  buf

  (
    g1345_n_spl_,
    g1345_n
  );


  buf

  (
    g1345_p_spl_,
    g1345_p
  );


  buf

  (
    g1340_n_spl_,
    g1340_n
  );


  buf

  (
    g1347_p_spl_,
    g1347_p
  );


  buf

  (
    g1340_p_spl_,
    g1340_p
  );


  buf

  (
    g1347_n_spl_,
    g1347_n
  );


  buf

  (
    g1348_n_spl_,
    g1348_n
  );


  buf

  (
    g1348_p_spl_,
    g1348_p
  );


  buf

  (
    g1339_n_spl_,
    g1339_n
  );


  buf

  (
    g1350_p_spl_,
    g1350_p
  );


  buf

  (
    g1339_p_spl_,
    g1339_p
  );


  buf

  (
    g1350_n_spl_,
    g1350_n
  );


  buf

  (
    g1351_n_spl_,
    g1351_n
  );


  buf

  (
    g1351_p_spl_,
    g1351_p
  );


  buf

  (
    g1352_n_spl_,
    g1352_n
  );


  buf

  (
    g1354_p_spl_,
    g1354_p
  );


  buf

  (
    g1352_p_spl_,
    g1352_p
  );


  buf

  (
    g1354_n_spl_,
    g1354_n
  );


  buf

  (
    g1355_n_spl_,
    g1355_n
  );


  buf

  (
    g1355_p_spl_,
    g1355_p
  );


  buf

  (
    ffc_189_p_spl_,
    ffc_189_p
  );


  buf

  (
    ffc_189_p_spl_0,
    ffc_189_p_spl_
  );


  buf

  (
    ffc_189_p_spl_1,
    ffc_189_p_spl_
  );


  buf

  (
    ffc_189_n_spl_,
    ffc_189_n
  );


  buf

  (
    ffc_189_n_spl_0,
    ffc_189_n_spl_
  );


  buf

  (
    g1360_n_spl_,
    g1360_n
  );


  buf

  (
    g1362_p_spl_,
    g1362_p
  );


  buf

  (
    g1360_p_spl_,
    g1360_p
  );


  buf

  (
    g1362_n_spl_,
    g1362_n
  );


  buf

  (
    g1363_n_spl_,
    g1363_n
  );


  buf

  (
    g1363_p_spl_,
    g1363_p
  );


  buf

  (
    g1359_n_spl_,
    g1359_n
  );


  buf

  (
    g1365_p_spl_,
    g1365_p
  );


  buf

  (
    g1359_p_spl_,
    g1359_p
  );


  buf

  (
    g1365_n_spl_,
    g1365_n
  );


  buf

  (
    g1366_n_spl_,
    g1366_n
  );


  buf

  (
    g1366_p_spl_,
    g1366_p
  );


  buf

  (
    g1358_n_spl_,
    g1358_n
  );


  buf

  (
    g1368_p_spl_,
    g1368_p
  );


  buf

  (
    g1358_p_spl_,
    g1358_p
  );


  buf

  (
    g1368_n_spl_,
    g1368_n
  );


  buf

  (
    g1369_n_spl_,
    g1369_n
  );


  buf

  (
    g1369_p_spl_,
    g1369_p
  );


  buf

  (
    g1357_n_spl_,
    g1357_n
  );


  buf

  (
    g1371_p_spl_,
    g1371_p
  );


  buf

  (
    g1357_p_spl_,
    g1357_p
  );


  buf

  (
    g1371_n_spl_,
    g1371_n
  );


  buf

  (
    g1372_n_spl_,
    g1372_n
  );


  buf

  (
    g1372_p_spl_,
    g1372_p
  );


  buf

  (
    g1356_n_spl_,
    g1356_n
  );


  buf

  (
    g1374_p_spl_,
    g1374_p
  );


  buf

  (
    g1356_p_spl_,
    g1356_p
  );


  buf

  (
    g1374_n_spl_,
    g1374_n
  );


  buf

  (
    g1375_n_spl_,
    g1375_n
  );


  buf

  (
    g1375_p_spl_,
    g1375_p
  );


  buf

  (
    g1376_n_spl_,
    g1376_n
  );


  buf

  (
    g1378_p_spl_,
    g1378_p
  );


  buf

  (
    g1376_p_spl_,
    g1376_p
  );


  buf

  (
    g1378_n_spl_,
    g1378_n
  );


  buf

  (
    g1379_n_spl_,
    g1379_n
  );


  buf

  (
    g1379_p_spl_,
    g1379_p
  );


  buf

  (
    g1384_n_spl_,
    g1384_n
  );


  buf

  (
    g1386_p_spl_,
    g1386_p
  );


  buf

  (
    g1384_p_spl_,
    g1384_p
  );


  buf

  (
    g1386_n_spl_,
    g1386_n
  );


  buf

  (
    g1387_n_spl_,
    g1387_n
  );


  buf

  (
    g1387_p_spl_,
    g1387_p
  );


  buf

  (
    g1383_n_spl_,
    g1383_n
  );


  buf

  (
    g1389_p_spl_,
    g1389_p
  );


  buf

  (
    g1383_p_spl_,
    g1383_p
  );


  buf

  (
    g1389_n_spl_,
    g1389_n
  );


  buf

  (
    g1390_n_spl_,
    g1390_n
  );


  buf

  (
    g1390_p_spl_,
    g1390_p
  );


  buf

  (
    g1382_n_spl_,
    g1382_n
  );


  buf

  (
    g1392_p_spl_,
    g1392_p
  );


  buf

  (
    g1382_p_spl_,
    g1382_p
  );


  buf

  (
    g1392_n_spl_,
    g1392_n
  );


  buf

  (
    g1393_n_spl_,
    g1393_n
  );


  buf

  (
    g1393_p_spl_,
    g1393_p
  );


  buf

  (
    g1381_n_spl_,
    g1381_n
  );


  buf

  (
    g1395_p_spl_,
    g1395_p
  );


  buf

  (
    g1381_p_spl_,
    g1381_p
  );


  buf

  (
    g1395_n_spl_,
    g1395_n
  );


  buf

  (
    g1396_n_spl_,
    g1396_n
  );


  buf

  (
    g1396_p_spl_,
    g1396_p
  );


  buf

  (
    g1380_n_spl_,
    g1380_n
  );


  buf

  (
    g1398_p_spl_,
    g1398_p
  );


  buf

  (
    g1380_p_spl_,
    g1380_p
  );


  buf

  (
    g1398_n_spl_,
    g1398_n
  );


  buf

  (
    g1250_p_spl_,
    g1250_p
  );


  buf

  (
    g1016_p_spl_,
    g1016_p
  );


  buf

  (
    ffc_21_n_spl_,
    ffc_21_n
  );


  buf

  (
    ffc_21_n_spl_0,
    ffc_21_n_spl_
  );


  buf

  (
    ffc_21_n_spl_00,
    ffc_21_n_spl_0
  );


  buf

  (
    ffc_21_n_spl_1,
    ffc_21_n_spl_
  );


  buf

  (
    ffc_12_n_spl_,
    ffc_12_n
  );


  buf

  (
    ffc_12_n_spl_0,
    ffc_12_n_spl_
  );


  buf

  (
    ffc_12_n_spl_00,
    ffc_12_n_spl_0
  );


  buf

  (
    ffc_12_n_spl_000,
    ffc_12_n_spl_00
  );


  buf

  (
    ffc_12_n_spl_001,
    ffc_12_n_spl_00
  );


  buf

  (
    ffc_12_n_spl_01,
    ffc_12_n_spl_0
  );


  buf

  (
    ffc_12_n_spl_010,
    ffc_12_n_spl_01
  );


  buf

  (
    ffc_12_n_spl_1,
    ffc_12_n_spl_
  );


  buf

  (
    ffc_12_n_spl_10,
    ffc_12_n_spl_1
  );


  buf

  (
    ffc_12_n_spl_11,
    ffc_12_n_spl_1
  );


  buf

  (
    G20_n_spl_,
    G20_n
  );


  buf

  (
    G20_n_spl_0,
    G20_n_spl_
  );


  buf

  (
    G20_n_spl_00,
    G20_n_spl_0
  );


  buf

  (
    G20_n_spl_000,
    G20_n_spl_00
  );


  buf

  (
    G20_n_spl_001,
    G20_n_spl_00
  );


  buf

  (
    G20_n_spl_01,
    G20_n_spl_0
  );


  buf

  (
    G20_n_spl_010,
    G20_n_spl_01
  );


  buf

  (
    G20_n_spl_011,
    G20_n_spl_01
  );


  buf

  (
    G20_n_spl_1,
    G20_n_spl_
  );


  buf

  (
    G20_n_spl_10,
    G20_n_spl_1
  );


  buf

  (
    G20_n_spl_100,
    G20_n_spl_10
  );


  buf

  (
    G20_n_spl_101,
    G20_n_spl_10
  );


  buf

  (
    G20_n_spl_11,
    G20_n_spl_1
  );


  buf

  (
    G20_n_spl_110,
    G20_n_spl_11
  );


  buf

  (
    g946_n_spl_,
    g946_n
  );


  buf

  (
    g1404_n_spl_,
    g1404_n
  );


  buf

  (
    g1406_p_spl_,
    g1406_p
  );


  buf

  (
    g934_n_spl_,
    g934_n
  );


  buf

  (
    g1409_n_spl_,
    g1409_n
  );


  buf

  (
    g1411_p_spl_,
    g1411_p
  );


  buf

  (
    g922_n_spl_,
    g922_n
  );


  buf

  (
    g1414_n_spl_,
    g1414_n
  );


  buf

  (
    g1416_p_spl_,
    g1416_p
  );


  buf

  (
    g919_n_spl_,
    g919_n
  );


  buf

  (
    g1419_n_spl_,
    g1419_n
  );


  buf

  (
    g1421_p_spl_,
    g1421_p
  );


  buf

  (
    g915_n_spl_,
    g915_n
  );


  buf

  (
    g1424_n_spl_,
    g1424_n
  );


  buf

  (
    g1426_p_spl_,
    g1426_p
  );


  buf

  (
    g911_n_spl_,
    g911_n
  );


  buf

  (
    g1429_n_spl_,
    g1429_n
  );


  buf

  (
    g1431_p_spl_,
    g1431_p
  );


  buf

  (
    g1013_n_spl_,
    g1013_n
  );


  buf

  (
    g1015_p_spl_,
    g1015_p
  );


  buf

  (
    ffc_21_p_spl_,
    ffc_21_p
  );


  buf

  (
    ffc_21_p_spl_0,
    ffc_21_p_spl_
  );


  buf

  (
    ffc_21_p_spl_00,
    ffc_21_p_spl_0
  );


  buf

  (
    ffc_21_p_spl_1,
    ffc_21_p_spl_
  );


  buf

  (
    g1241_n_spl_,
    g1241_n
  );


  buf

  (
    g1164_n_spl_,
    g1164_n
  );


  buf

  (
    g1107_n_spl_,
    g1107_n
  );


  buf

  (
    g1053_n_spl_,
    g1053_n
  );


  buf

  (
    g1459_n_spl_,
    g1459_n
  );


  buf

  (
    g1461_p_spl_,
    g1461_p
  );


  buf

  (
    g1459_p_spl_,
    g1459_p
  );


  buf

  (
    g1461_n_spl_,
    g1461_n
  );


  buf

  (
    g1462_n_spl_,
    g1462_n
  );


  buf

  (
    g1462_p_spl_,
    g1462_p
  );


  buf

  (
    g1458_n_spl_,
    g1458_n
  );


  buf

  (
    g1464_p_spl_,
    g1464_p
  );


  buf

  (
    g1458_p_spl_,
    g1458_p
  );


  buf

  (
    g1464_n_spl_,
    g1464_n
  );


  buf

  (
    g1465_n_spl_,
    g1465_n
  );


  buf

  (
    g1465_p_spl_,
    g1465_p
  );


  buf

  (
    g1457_n_spl_,
    g1457_n
  );


  buf

  (
    g1467_p_spl_,
    g1467_p
  );


  buf

  (
    g1457_p_spl_,
    g1457_p
  );


  buf

  (
    g1467_n_spl_,
    g1467_n
  );


  buf

  (
    g1468_n_spl_,
    g1468_n
  );


  buf

  (
    g1468_p_spl_,
    g1468_p
  );


  buf

  (
    g1456_n_spl_,
    g1456_n
  );


  buf

  (
    g1470_p_spl_,
    g1470_p
  );


  buf

  (
    g1456_p_spl_,
    g1456_p
  );


  buf

  (
    g1470_n_spl_,
    g1470_n
  );


  buf

  (
    g1471_n_spl_,
    g1471_n
  );


  buf

  (
    g1471_p_spl_,
    g1471_p
  );


  buf

  (
    g1455_n_spl_,
    g1455_n
  );


  buf

  (
    g1473_p_spl_,
    g1473_p
  );


  buf

  (
    g1454_n_spl_,
    g1454_n
  );


  buf

  (
    g1476_p_spl_,
    g1476_p
  );


  buf

  (
    g1480_n_spl_,
    g1480_n
  );


  buf

  (
    g1482_p_spl_,
    g1482_p
  );


  buf

  (
    g1480_p_spl_,
    g1480_p
  );


  buf

  (
    g1482_n_spl_,
    g1482_n
  );


  buf

  (
    g1483_n_spl_,
    g1483_n
  );


  buf

  (
    g1479_n_spl_,
    g1479_n
  );


  buf

  (
    g1485_p_spl_,
    g1485_p
  );


  buf

  (
    g1479_p_spl_,
    g1479_p
  );


  buf

  (
    g1485_n_spl_,
    g1485_n
  );


  buf

  (
    g1486_n_spl_,
    g1486_n
  );


  buf

  (
    g1492_n_spl_,
    g1492_n
  );


  buf

  (
    g1494_p_spl_,
    g1494_p
  );


  buf

  (
    g1492_p_spl_,
    g1492_p
  );


  buf

  (
    g1494_n_spl_,
    g1494_n
  );


  buf

  (
    g1495_n_spl_,
    g1495_n
  );


  buf

  (
    g1491_n_spl_,
    g1491_n
  );


  buf

  (
    g1497_p_spl_,
    g1497_p
  );


  buf

  (
    g1491_p_spl_,
    g1491_p
  );


  buf

  (
    g1497_n_spl_,
    g1497_n
  );


  buf

  (
    g1498_n_spl_,
    g1498_n
  );


  buf

  (
    g1504_n_spl_,
    g1504_n
  );


  buf

  (
    g1506_p_spl_,
    g1506_p
  );


  buf

  (
    g1504_p_spl_,
    g1504_p
  );


  buf

  (
    g1506_n_spl_,
    g1506_n
  );


  buf

  (
    g1507_n_spl_,
    g1507_n
  );


  buf

  (
    g1503_n_spl_,
    g1503_n
  );


  buf

  (
    g1509_p_spl_,
    g1509_p
  );


  buf

  (
    g1503_p_spl_,
    g1503_p
  );


  buf

  (
    g1509_n_spl_,
    g1509_n
  );


  buf

  (
    g1510_n_spl_,
    g1510_n
  );


  buf

  (
    g1278_n_spl_,
    g1278_n
  );


  buf

  (
    ffc_12_p_spl_,
    ffc_12_p
  );


  buf

  (
    ffc_12_p_spl_0,
    ffc_12_p_spl_
  );


  buf

  (
    ffc_12_p_spl_00,
    ffc_12_p_spl_0
  );


  buf

  (
    ffc_12_p_spl_000,
    ffc_12_p_spl_00
  );


  buf

  (
    ffc_12_p_spl_001,
    ffc_12_p_spl_00
  );


  buf

  (
    ffc_12_p_spl_01,
    ffc_12_p_spl_0
  );


  buf

  (
    ffc_12_p_spl_1,
    ffc_12_p_spl_
  );


  buf

  (
    ffc_12_p_spl_10,
    ffc_12_p_spl_1
  );


  buf

  (
    ffc_12_p_spl_11,
    ffc_12_p_spl_1
  );


  buf

  (
    g1399_n_spl_,
    g1399_n
  );


  buf

  (
    g1328_n_spl_,
    g1328_n
  );


  buf

  (
    g1526_n_spl_,
    g1526_n
  );


  buf

  (
    g1527_n_spl_,
    g1527_n
  );


  buf

  (
    g1526_p_spl_,
    g1526_p
  );


  buf

  (
    g1527_p_spl_,
    g1527_p
  );


  buf

  (
    g1528_p_spl_,
    g1528_p
  );


  buf

  (
    g1525_n_spl_,
    g1525_n
  );


  buf

  (
    g1530_p_spl_,
    g1530_p
  );


  buf

  (
    g1525_p_spl_,
    g1525_p
  );


  buf

  (
    g1530_n_spl_,
    g1530_n
  );


  buf

  (
    g1531_p_spl_,
    g1531_p
  );


  buf

  (
    g1537_n_spl_,
    g1537_n
  );


  buf

  (
    g1539_p_spl_,
    g1539_p
  );


  buf

  (
    g1537_p_spl_,
    g1537_p
  );


  buf

  (
    g1539_n_spl_,
    g1539_n
  );


  buf

  (
    g1540_p_spl_,
    g1540_p
  );


  buf

  (
    g1536_n_spl_,
    g1536_n
  );


  buf

  (
    g1542_p_spl_,
    g1542_p
  );


  buf

  (
    g1536_p_spl_,
    g1536_p
  );


  buf

  (
    g1542_n_spl_,
    g1542_n
  );


  buf

  (
    g1543_p_spl_,
    g1543_p
  );


  buf

  (
    g1242_p_spl_,
    g1242_p
  );


  buf

  (
    ffc_181_p_spl_,
    ffc_181_p
  );


  buf

  (
    ffc_181_p_spl_0,
    ffc_181_p_spl_
  );


  buf

  (
    ffc_181_p_spl_00,
    ffc_181_p_spl_0
  );


  buf

  (
    ffc_181_p_spl_1,
    ffc_181_p_spl_
  );


  buf

  (
    ffc_181_n_spl_,
    ffc_181_n
  );


  buf

  (
    ffc_181_n_spl_0,
    ffc_181_n_spl_
  );


  buf

  (
    ffc_181_n_spl_1,
    ffc_181_n_spl_
  );


  buf

  (
    ffc_328_n_spl_,
    ffc_328_n
  );


  buf

  (
    ffc_345_p_spl_,
    ffc_345_p
  );


  buf

  (
    ffc_328_p_spl_,
    ffc_328_p
  );


  buf

  (
    ffc_345_n_spl_,
    ffc_345_n
  );


  buf

  (
    g1554_n_spl_,
    g1554_n
  );


  buf

  (
    g1554_p_spl_,
    g1554_p
  );


  buf

  (
    g1553_n_spl_,
    g1553_n
  );


  buf

  (
    g1556_p_spl_,
    g1556_p
  );


  buf

  (
    g1553_p_spl_,
    g1553_p
  );


  buf

  (
    g1556_n_spl_,
    g1556_n
  );


  buf

  (
    g1557_n_spl_,
    g1557_n
  );


  buf

  (
    g1557_p_spl_,
    g1557_p
  );


  buf

  (
    g1552_n_spl_,
    g1552_n
  );


  buf

  (
    g1559_p_spl_,
    g1559_p
  );


  buf

  (
    g1552_p_spl_,
    g1552_p
  );


  buf

  (
    g1559_n_spl_,
    g1559_n
  );


  buf

  (
    g1560_n_spl_,
    g1560_n
  );


  buf

  (
    g1560_p_spl_,
    g1560_p
  );


  buf

  (
    g1551_n_spl_,
    g1551_n
  );


  buf

  (
    g1562_p_spl_,
    g1562_p
  );


  buf

  (
    g1551_p_spl_,
    g1551_p
  );


  buf

  (
    g1562_n_spl_,
    g1562_n
  );


  buf

  (
    g1563_n_spl_,
    g1563_n
  );


  buf

  (
    g1563_p_spl_,
    g1563_p
  );


  buf

  (
    g1550_n_spl_,
    g1550_n
  );


  buf

  (
    g1565_p_spl_,
    g1565_p
  );


  buf

  (
    g1550_p_spl_,
    g1550_p
  );


  buf

  (
    g1565_n_spl_,
    g1565_n
  );


  buf

  (
    g1566_n_spl_,
    g1566_n
  );


  buf

  (
    g1566_p_spl_,
    g1566_p
  );


  buf

  (
    g1549_n_spl_,
    g1549_n
  );


  buf

  (
    g1568_p_spl_,
    g1568_p
  );


  buf

  (
    g1549_p_spl_,
    g1549_p
  );


  buf

  (
    g1568_n_spl_,
    g1568_n
  );


  buf

  (
    g1569_n_spl_,
    g1569_n
  );


  buf

  (
    g1569_p_spl_,
    g1569_p
  );


  buf

  (
    g1548_n_spl_,
    g1548_n
  );


  buf

  (
    g1571_p_spl_,
    g1571_p
  );


  buf

  (
    g1548_p_spl_,
    g1548_p
  );


  buf

  (
    g1571_n_spl_,
    g1571_n
  );


  buf

  (
    g1572_n_spl_,
    g1572_n
  );


  buf

  (
    g1572_p_spl_,
    g1572_p
  );


  buf

  (
    g1547_n_spl_,
    g1547_n
  );


  buf

  (
    g1574_p_spl_,
    g1574_p
  );


  buf

  (
    g1400_p_spl_,
    g1400_p
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_00,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_01,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    G4_n_spl_0,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_1,
    G4_n_spl_
  );


  buf

  (
    g1580_p_spl_,
    g1580_p
  );


  buf

  (
    g1581_p_spl_,
    g1581_p
  );


  buf

  (
    g1580_n_spl_,
    g1580_n
  );


  buf

  (
    g1581_n_spl_,
    g1581_n
  );


  buf

  (
    g1582_n_spl_,
    g1582_n
  );


  buf

  (
    g1582_n_spl_0,
    g1582_n_spl_
  );


  buf

  (
    g1582_p_spl_,
    g1582_p
  );


  buf

  (
    g1582_p_spl_0,
    g1582_p_spl_
  );


  buf

  (
    g1584_n_spl_,
    g1584_n
  );


  buf

  (
    g1584_p_spl_,
    g1584_p
  );


  buf

  (
    g1585_n_spl_,
    g1585_n
  );


  buf

  (
    g1585_p_spl_,
    g1585_p
  );


  buf

  (
    g1579_n_spl_,
    g1579_n
  );


  buf

  (
    g1587_p_spl_,
    g1587_p
  );


  buf

  (
    g1579_p_spl_,
    g1579_p
  );


  buf

  (
    g1587_n_spl_,
    g1587_n
  );


  buf

  (
    g1588_n_spl_,
    g1588_n
  );


  buf

  (
    g1588_p_spl_,
    g1588_p
  );


  buf

  (
    g1578_n_spl_,
    g1578_n
  );


  buf

  (
    g1590_p_spl_,
    g1590_p
  );


  buf

  (
    g1603_n_spl_,
    g1603_n
  );


  buf

  (
    g1605_p_spl_,
    g1605_p
  );


  buf

  (
    g1603_p_spl_,
    g1603_p
  );


  buf

  (
    g1605_n_spl_,
    g1605_n
  );


  buf

  (
    g1606_n_spl_,
    g1606_n
  );


  buf

  (
    g1606_p_spl_,
    g1606_p
  );


  buf

  (
    g1602_n_spl_,
    g1602_n
  );


  buf

  (
    g1608_p_spl_,
    g1608_p
  );


  buf

  (
    g1602_p_spl_,
    g1602_p
  );


  buf

  (
    g1608_n_spl_,
    g1608_n
  );


  buf

  (
    g1609_n_spl_,
    g1609_n
  );


  buf

  (
    g1609_p_spl_,
    g1609_p
  );


  buf

  (
    g1601_n_spl_,
    g1601_n
  );


  buf

  (
    g1611_p_spl_,
    g1611_p
  );


  buf

  (
    g1601_p_spl_,
    g1601_p
  );


  buf

  (
    g1611_n_spl_,
    g1611_n
  );


  buf

  (
    g1612_n_spl_,
    g1612_n
  );


  buf

  (
    g1616_n_spl_,
    g1616_n
  );


  buf

  (
    g1618_n_spl_,
    g1618_n
  );


  buf

  (
    g1620_p_spl_,
    g1620_p
  );


  buf

  (
    g1618_p_spl_,
    g1618_p
  );


  buf

  (
    g1620_n_spl_,
    g1620_n
  );


  buf

  (
    g1621_n_spl_,
    g1621_n
  );


  buf

  (
    g1625_n_spl_,
    g1625_n
  );


  buf

  (
    g1477_p_spl_,
    g1477_p
  );


  buf

  (
    g1401_n_spl_,
    g1401_n
  );


  buf

  (
    g1515_p_spl_,
    g1515_p
  );


  buf

  (
    g1402_n_spl_,
    g1402_n
  );


  buf

  (
    g1577_p_spl_,
    g1577_p
  );


  buf

  (
    g1403_n_spl_,
    g1403_n
  );


  buf

  (
    g1593_p_spl_,
    g1593_p
  );


  buf

  (
    g1438_n_spl_,
    g1438_n
  );


  buf

  (
    g1442_n_spl_,
    g1442_n
  );


  buf

  (
    g1446_n_spl_,
    g1446_n
  );


  buf

  (
    g1450_n_spl_,
    g1450_n
  );


  buf

  (
    g1453_n_spl_,
    g1453_n
  );


  buf

  (
    g1489_n_spl_,
    g1489_n
  );


  buf

  (
    g1501_n_spl_,
    g1501_n
  );


  buf

  (
    g1513_n_spl_,
    g1513_n
  );


  buf

  (
    g1630_p_spl_,
    g1630_p
  );


  buf

  (
    ffc_182_p_spl_,
    ffc_182_p
  );


  buf

  (
    ffc_182_p_spl_0,
    ffc_182_p_spl_
  );


  buf

  (
    ffc_182_p_spl_00,
    ffc_182_p_spl_0
  );


  buf

  (
    ffc_182_p_spl_1,
    ffc_182_p_spl_
  );


  buf

  (
    ffc_182_n_spl_,
    ffc_182_n
  );


  buf

  (
    ffc_182_n_spl_0,
    ffc_182_n_spl_
  );


  buf

  (
    ffc_182_n_spl_1,
    ffc_182_n_spl_
  );


  buf

  (
    ffc_329_n_spl_,
    ffc_329_n
  );


  buf

  (
    ffc_346_p_spl_,
    ffc_346_p
  );


  buf

  (
    ffc_329_p_spl_,
    ffc_329_p
  );


  buf

  (
    ffc_346_n_spl_,
    ffc_346_n
  );


  buf

  (
    g1661_n_spl_,
    g1661_n
  );


  buf

  (
    g1661_p_spl_,
    g1661_p
  );


  buf

  (
    g1660_n_spl_,
    g1660_n
  );


  buf

  (
    g1663_p_spl_,
    g1663_p
  );


  buf

  (
    g1660_p_spl_,
    g1660_p
  );


  buf

  (
    g1663_n_spl_,
    g1663_n
  );


  buf

  (
    g1664_n_spl_,
    g1664_n
  );


  buf

  (
    g1664_p_spl_,
    g1664_p
  );


  buf

  (
    g1659_n_spl_,
    g1659_n
  );


  buf

  (
    g1666_p_spl_,
    g1666_p
  );


  buf

  (
    g1659_p_spl_,
    g1659_p
  );


  buf

  (
    g1666_n_spl_,
    g1666_n
  );


  buf

  (
    g1667_n_spl_,
    g1667_n
  );


  buf

  (
    g1667_p_spl_,
    g1667_p
  );


  buf

  (
    g1658_n_spl_,
    g1658_n
  );


  buf

  (
    g1669_p_spl_,
    g1669_p
  );


  buf

  (
    g1658_p_spl_,
    g1658_p
  );


  buf

  (
    g1669_n_spl_,
    g1669_n
  );


  buf

  (
    g1670_n_spl_,
    g1670_n
  );


  buf

  (
    g1670_p_spl_,
    g1670_p
  );


  buf

  (
    g1657_n_spl_,
    g1657_n
  );


  buf

  (
    g1672_p_spl_,
    g1672_p
  );


  buf

  (
    g1657_p_spl_,
    g1657_p
  );


  buf

  (
    g1672_n_spl_,
    g1672_n
  );


  buf

  (
    g1673_n_spl_,
    g1673_n
  );


  buf

  (
    g1673_p_spl_,
    g1673_p
  );


  buf

  (
    g1656_n_spl_,
    g1656_n
  );


  buf

  (
    g1675_p_spl_,
    g1675_p
  );


  buf

  (
    g1656_p_spl_,
    g1656_p
  );


  buf

  (
    g1675_n_spl_,
    g1675_n
  );


  buf

  (
    g1676_n_spl_,
    g1676_n
  );


  buf

  (
    g1676_p_spl_,
    g1676_p
  );


  buf

  (
    g1655_n_spl_,
    g1655_n
  );


  buf

  (
    g1678_p_spl_,
    g1678_p
  );


  buf

  (
    g1655_p_spl_,
    g1655_p
  );


  buf

  (
    g1678_n_spl_,
    g1678_n
  );


  buf

  (
    g1679_n_spl_,
    g1679_n
  );


  buf

  (
    g1679_p_spl_,
    g1679_p
  );


  buf

  (
    g1654_n_spl_,
    g1654_n
  );


  buf

  (
    g1681_p_spl_,
    g1681_p
  );


  buf

  (
    g1654_p_spl_,
    g1654_p
  );


  buf

  (
    g1681_n_spl_,
    g1681_n
  );


  buf

  (
    g1682_n_spl_,
    g1682_n
  );


  buf

  (
    g1685_n_spl_,
    g1685_n
  );


  buf

  (
    g1546_n_spl_,
    g1546_n
  );


  buf

  (
    g1688_n_spl_,
    g1688_n
  );


  buf

  (
    g1690_p_spl_,
    g1690_p
  );


  buf

  (
    g1534_n_spl_,
    g1534_n
  );


  buf

  (
    g1693_n_spl_,
    g1693_n
  );


  buf

  (
    g1695_p_spl_,
    g1695_p
  );


  buf

  (
    g1698_n_spl_,
    g1698_n
  );


  buf

  (
    g1699_n_spl_,
    g1699_n
  );


  buf

  (
    g1523_n_spl_,
    g1523_n
  );


  buf

  (
    g1702_n_spl_,
    g1702_n
  );


  buf

  (
    g1704_p_spl_,
    g1704_p
  );


  buf

  (
    ffc_183_p_spl_,
    ffc_183_p
  );


  buf

  (
    ffc_183_p_spl_0,
    ffc_183_p_spl_
  );


  buf

  (
    ffc_183_p_spl_00,
    ffc_183_p_spl_0
  );


  buf

  (
    ffc_183_p_spl_1,
    ffc_183_p_spl_
  );


  buf

  (
    ffc_183_n_spl_,
    ffc_183_n
  );


  buf

  (
    ffc_183_n_spl_0,
    ffc_183_n_spl_
  );


  buf

  (
    ffc_183_n_spl_1,
    ffc_183_n_spl_
  );


  buf

  (
    ffc_330_n_spl_,
    ffc_330_n
  );


  buf

  (
    ffc_347_p_spl_,
    ffc_347_p
  );


  buf

  (
    ffc_330_p_spl_,
    ffc_330_p
  );


  buf

  (
    ffc_347_n_spl_,
    ffc_347_n
  );


  buf

  (
    g1714_n_spl_,
    g1714_n
  );


  buf

  (
    g1714_p_spl_,
    g1714_p
  );


  buf

  (
    g1713_n_spl_,
    g1713_n
  );


  buf

  (
    g1716_p_spl_,
    g1716_p
  );


  buf

  (
    g1713_p_spl_,
    g1713_p
  );


  buf

  (
    g1716_n_spl_,
    g1716_n
  );


  buf

  (
    g1717_n_spl_,
    g1717_n
  );


  buf

  (
    g1717_p_spl_,
    g1717_p
  );


  buf

  (
    g1712_n_spl_,
    g1712_n
  );


  buf

  (
    g1719_p_spl_,
    g1719_p
  );


  buf

  (
    g1712_p_spl_,
    g1712_p
  );


  buf

  (
    g1719_n_spl_,
    g1719_n
  );


  buf

  (
    g1720_n_spl_,
    g1720_n
  );


  buf

  (
    g1720_p_spl_,
    g1720_p
  );


  buf

  (
    g1711_n_spl_,
    g1711_n
  );


  buf

  (
    g1722_p_spl_,
    g1722_p
  );


  buf

  (
    g1711_p_spl_,
    g1711_p
  );


  buf

  (
    g1722_n_spl_,
    g1722_n
  );


  buf

  (
    g1723_n_spl_,
    g1723_n
  );


  buf

  (
    g1723_p_spl_,
    g1723_p
  );


  buf

  (
    g1710_n_spl_,
    g1710_n
  );


  buf

  (
    g1725_p_spl_,
    g1725_p
  );


  buf

  (
    g1710_p_spl_,
    g1710_p
  );


  buf

  (
    g1725_n_spl_,
    g1725_n
  );


  buf

  (
    g1726_n_spl_,
    g1726_n
  );


  buf

  (
    g1726_p_spl_,
    g1726_p
  );


  buf

  (
    g1709_n_spl_,
    g1709_n
  );


  buf

  (
    g1728_p_spl_,
    g1728_p
  );


  buf

  (
    g1709_p_spl_,
    g1709_p
  );


  buf

  (
    g1728_n_spl_,
    g1728_n
  );


  buf

  (
    g1729_n_spl_,
    g1729_n
  );


  buf

  (
    g1729_p_spl_,
    g1729_p
  );


  buf

  (
    g1708_n_spl_,
    g1708_n
  );


  buf

  (
    g1731_p_spl_,
    g1731_p
  );


  buf

  (
    g1708_p_spl_,
    g1708_p
  );


  buf

  (
    g1731_n_spl_,
    g1731_n
  );


  buf

  (
    g1732_n_spl_,
    g1732_n
  );


  buf

  (
    g1732_p_spl_,
    g1732_p
  );


  buf

  (
    g1707_n_spl_,
    g1707_n
  );


  buf

  (
    g1734_p_spl_,
    g1734_p
  );


  buf

  (
    g1707_p_spl_,
    g1707_p
  );


  buf

  (
    g1734_n_spl_,
    g1734_n
  );


  buf

  (
    g1735_p_spl_,
    g1735_p
  );


  buf

  (
    g1739_p_spl_,
    g1739_p
  );


  buf

  (
    ffc_184_p_spl_,
    ffc_184_p
  );


  buf

  (
    ffc_184_p_spl_0,
    ffc_184_p_spl_
  );


  buf

  (
    ffc_184_p_spl_00,
    ffc_184_p_spl_0
  );


  buf

  (
    ffc_184_p_spl_1,
    ffc_184_p_spl_
  );


  buf

  (
    ffc_184_n_spl_,
    ffc_184_n
  );


  buf

  (
    ffc_184_n_spl_0,
    ffc_184_n_spl_
  );


  buf

  (
    ffc_184_n_spl_1,
    ffc_184_n_spl_
  );


  buf

  (
    ffc_331_n_spl_,
    ffc_331_n
  );


  buf

  (
    ffc_348_p_spl_,
    ffc_348_p
  );


  buf

  (
    ffc_331_p_spl_,
    ffc_331_p
  );


  buf

  (
    ffc_348_n_spl_,
    ffc_348_n
  );


  buf

  (
    g1749_n_spl_,
    g1749_n
  );


  buf

  (
    g1749_p_spl_,
    g1749_p
  );


  buf

  (
    g1748_n_spl_,
    g1748_n
  );


  buf

  (
    g1751_p_spl_,
    g1751_p
  );


  buf

  (
    g1748_p_spl_,
    g1748_p
  );


  buf

  (
    g1751_n_spl_,
    g1751_n
  );


  buf

  (
    g1752_n_spl_,
    g1752_n
  );


  buf

  (
    g1752_p_spl_,
    g1752_p
  );


  buf

  (
    g1747_n_spl_,
    g1747_n
  );


  buf

  (
    g1754_p_spl_,
    g1754_p
  );


  buf

  (
    g1747_p_spl_,
    g1747_p
  );


  buf

  (
    g1754_n_spl_,
    g1754_n
  );


  buf

  (
    g1755_n_spl_,
    g1755_n
  );


  buf

  (
    g1755_p_spl_,
    g1755_p
  );


  buf

  (
    g1746_n_spl_,
    g1746_n
  );


  buf

  (
    g1757_p_spl_,
    g1757_p
  );


  buf

  (
    g1746_p_spl_,
    g1746_p
  );


  buf

  (
    g1757_n_spl_,
    g1757_n
  );


  buf

  (
    g1758_n_spl_,
    g1758_n
  );


  buf

  (
    g1758_p_spl_,
    g1758_p
  );


  buf

  (
    g1745_n_spl_,
    g1745_n
  );


  buf

  (
    g1760_p_spl_,
    g1760_p
  );


  buf

  (
    g1745_p_spl_,
    g1745_p
  );


  buf

  (
    g1760_n_spl_,
    g1760_n
  );


  buf

  (
    g1761_n_spl_,
    g1761_n
  );


  buf

  (
    g1761_p_spl_,
    g1761_p
  );


  buf

  (
    g1744_n_spl_,
    g1744_n
  );


  buf

  (
    g1763_p_spl_,
    g1763_p
  );


  buf

  (
    g1744_p_spl_,
    g1744_p
  );


  buf

  (
    g1763_n_spl_,
    g1763_n
  );


  buf

  (
    g1764_n_spl_,
    g1764_n
  );


  buf

  (
    g1764_p_spl_,
    g1764_p
  );


  buf

  (
    g1743_n_spl_,
    g1743_n
  );


  buf

  (
    g1766_p_spl_,
    g1766_p
  );


  buf

  (
    g1743_p_spl_,
    g1743_p
  );


  buf

  (
    g1766_n_spl_,
    g1766_n
  );


  buf

  (
    g1767_n_spl_,
    g1767_n
  );


  buf

  (
    g1767_p_spl_,
    g1767_p
  );


  buf

  (
    g1742_n_spl_,
    g1742_n
  );


  buf

  (
    g1769_p_spl_,
    g1769_p
  );


  buf

  (
    g1742_p_spl_,
    g1742_p
  );


  buf

  (
    g1769_n_spl_,
    g1769_n
  );


  buf

  (
    g1770_p_spl_,
    g1770_p
  );


  buf

  (
    g1741_n_spl_,
    g1741_n
  );


  buf

  (
    g1772_p_spl_,
    g1772_p
  );


  buf

  (
    g1740_n_spl_,
    g1740_n
  );


  buf

  (
    g1775_p_spl_,
    g1775_p
  );


  buf

  (
    ffc_185_p_spl_,
    ffc_185_p
  );


  buf

  (
    ffc_185_p_spl_0,
    ffc_185_p_spl_
  );


  buf

  (
    ffc_185_p_spl_00,
    ffc_185_p_spl_0
  );


  buf

  (
    ffc_185_p_spl_1,
    ffc_185_p_spl_
  );


  buf

  (
    ffc_185_n_spl_,
    ffc_185_n
  );


  buf

  (
    ffc_185_n_spl_0,
    ffc_185_n_spl_
  );


  buf

  (
    ffc_185_n_spl_1,
    ffc_185_n_spl_
  );


  buf

  (
    ffc_332_n_spl_,
    ffc_332_n
  );


  buf

  (
    ffc_349_p_spl_,
    ffc_349_p
  );


  buf

  (
    ffc_332_p_spl_,
    ffc_332_p
  );


  buf

  (
    ffc_349_n_spl_,
    ffc_349_n
  );


  buf

  (
    g1787_n_spl_,
    g1787_n
  );


  buf

  (
    g1787_p_spl_,
    g1787_p
  );


  buf

  (
    g1786_n_spl_,
    g1786_n
  );


  buf

  (
    g1789_p_spl_,
    g1789_p
  );


  buf

  (
    g1786_p_spl_,
    g1786_p
  );


  buf

  (
    g1789_n_spl_,
    g1789_n
  );


  buf

  (
    g1790_n_spl_,
    g1790_n
  );


  buf

  (
    g1790_p_spl_,
    g1790_p
  );


  buf

  (
    g1785_n_spl_,
    g1785_n
  );


  buf

  (
    g1792_p_spl_,
    g1792_p
  );


  buf

  (
    g1785_p_spl_,
    g1785_p
  );


  buf

  (
    g1792_n_spl_,
    g1792_n
  );


  buf

  (
    g1793_n_spl_,
    g1793_n
  );


  buf

  (
    g1793_p_spl_,
    g1793_p
  );


  buf

  (
    g1784_n_spl_,
    g1784_n
  );


  buf

  (
    g1795_p_spl_,
    g1795_p
  );


  buf

  (
    g1784_p_spl_,
    g1784_p
  );


  buf

  (
    g1795_n_spl_,
    g1795_n
  );


  buf

  (
    g1796_n_spl_,
    g1796_n
  );


  buf

  (
    g1796_p_spl_,
    g1796_p
  );


  buf

  (
    g1783_n_spl_,
    g1783_n
  );


  buf

  (
    g1798_p_spl_,
    g1798_p
  );


  buf

  (
    g1783_p_spl_,
    g1783_p
  );


  buf

  (
    g1798_n_spl_,
    g1798_n
  );


  buf

  (
    g1799_n_spl_,
    g1799_n
  );


  buf

  (
    g1799_p_spl_,
    g1799_p
  );


  buf

  (
    g1782_n_spl_,
    g1782_n
  );


  buf

  (
    g1801_p_spl_,
    g1801_p
  );


  buf

  (
    g1782_p_spl_,
    g1782_p
  );


  buf

  (
    g1801_n_spl_,
    g1801_n
  );


  buf

  (
    g1802_n_spl_,
    g1802_n
  );


  buf

  (
    g1802_p_spl_,
    g1802_p
  );


  buf

  (
    g1781_n_spl_,
    g1781_n
  );


  buf

  (
    g1804_p_spl_,
    g1804_p
  );


  buf

  (
    g1781_p_spl_,
    g1781_p
  );


  buf

  (
    g1804_n_spl_,
    g1804_n
  );


  buf

  (
    g1805_n_spl_,
    g1805_n
  );


  buf

  (
    g1805_p_spl_,
    g1805_p
  );


  buf

  (
    g1780_n_spl_,
    g1780_n
  );


  buf

  (
    g1807_p_spl_,
    g1807_p
  );


  buf

  (
    g1780_p_spl_,
    g1780_p
  );


  buf

  (
    g1807_n_spl_,
    g1807_n
  );


  buf

  (
    g1808_p_spl_,
    g1808_p
  );


  buf

  (
    g1779_n_spl_,
    g1779_n
  );


  buf

  (
    g1810_p_spl_,
    g1810_p
  );


  buf

  (
    g1778_n_spl_,
    g1778_n
  );


  buf

  (
    g1813_p_spl_,
    g1813_p
  );


  buf

  (
    ffc_186_p_spl_,
    ffc_186_p
  );


  buf

  (
    ffc_186_p_spl_0,
    ffc_186_p_spl_
  );


  buf

  (
    ffc_186_p_spl_00,
    ffc_186_p_spl_0
  );


  buf

  (
    ffc_186_p_spl_1,
    ffc_186_p_spl_
  );


  buf

  (
    ffc_186_n_spl_,
    ffc_186_n
  );


  buf

  (
    ffc_186_n_spl_0,
    ffc_186_n_spl_
  );


  buf

  (
    ffc_186_n_spl_1,
    ffc_186_n_spl_
  );


  buf

  (
    g1824_n_spl_,
    g1824_n
  );


  buf

  (
    g1826_p_spl_,
    g1826_p
  );


  buf

  (
    g1824_p_spl_,
    g1824_p
  );


  buf

  (
    g1826_n_spl_,
    g1826_n
  );


  buf

  (
    g1827_n_spl_,
    g1827_n
  );


  buf

  (
    g1827_p_spl_,
    g1827_p
  );


  buf

  (
    g1823_n_spl_,
    g1823_n
  );


  buf

  (
    g1829_p_spl_,
    g1829_p
  );


  buf

  (
    g1823_p_spl_,
    g1823_p
  );


  buf

  (
    g1829_n_spl_,
    g1829_n
  );


  buf

  (
    g1830_n_spl_,
    g1830_n
  );


  buf

  (
    g1830_p_spl_,
    g1830_p
  );


  buf

  (
    g1822_n_spl_,
    g1822_n
  );


  buf

  (
    g1832_p_spl_,
    g1832_p
  );


  buf

  (
    g1822_p_spl_,
    g1822_p
  );


  buf

  (
    g1832_n_spl_,
    g1832_n
  );


  buf

  (
    g1833_n_spl_,
    g1833_n
  );


  buf

  (
    g1833_p_spl_,
    g1833_p
  );


  buf

  (
    g1821_n_spl_,
    g1821_n
  );


  buf

  (
    g1835_p_spl_,
    g1835_p
  );


  buf

  (
    g1821_p_spl_,
    g1821_p
  );


  buf

  (
    g1835_n_spl_,
    g1835_n
  );


  buf

  (
    g1836_n_spl_,
    g1836_n
  );


  buf

  (
    g1836_p_spl_,
    g1836_p
  );


  buf

  (
    g1820_n_spl_,
    g1820_n
  );


  buf

  (
    g1838_p_spl_,
    g1838_p
  );


  buf

  (
    g1820_p_spl_,
    g1820_p
  );


  buf

  (
    g1838_n_spl_,
    g1838_n
  );


  buf

  (
    g1839_n_spl_,
    g1839_n
  );


  buf

  (
    g1839_p_spl_,
    g1839_p
  );


  buf

  (
    g1819_n_spl_,
    g1819_n
  );


  buf

  (
    g1841_p_spl_,
    g1841_p
  );


  buf

  (
    g1819_p_spl_,
    g1819_p
  );


  buf

  (
    g1841_n_spl_,
    g1841_n
  );


  buf

  (
    g1842_n_spl_,
    g1842_n
  );


  buf

  (
    g1842_p_spl_,
    g1842_p
  );


  buf

  (
    g1818_n_spl_,
    g1818_n
  );


  buf

  (
    g1844_p_spl_,
    g1844_p
  );


  buf

  (
    g1818_p_spl_,
    g1818_p
  );


  buf

  (
    g1844_n_spl_,
    g1844_n
  );


  buf

  (
    g1845_p_spl_,
    g1845_p
  );


  buf

  (
    g1817_n_spl_,
    g1817_n
  );


  buf

  (
    g1847_p_spl_,
    g1847_p
  );


  buf

  (
    g1816_n_spl_,
    g1816_n
  );


  buf

  (
    g1850_p_spl_,
    g1850_p
  );


  buf

  (
    g1859_n_spl_,
    g1859_n
  );


  buf

  (
    g1861_p_spl_,
    g1861_p
  );


  buf

  (
    g1859_p_spl_,
    g1859_p
  );


  buf

  (
    g1861_n_spl_,
    g1861_n
  );


  buf

  (
    g1862_n_spl_,
    g1862_n
  );


  buf

  (
    g1862_p_spl_,
    g1862_p
  );


  buf

  (
    g1858_n_spl_,
    g1858_n
  );


  buf

  (
    g1864_p_spl_,
    g1864_p
  );


  buf

  (
    g1858_p_spl_,
    g1858_p
  );


  buf

  (
    g1864_n_spl_,
    g1864_n
  );


  buf

  (
    g1865_n_spl_,
    g1865_n
  );


  buf

  (
    g1865_p_spl_,
    g1865_p
  );


  buf

  (
    g1857_n_spl_,
    g1857_n
  );


  buf

  (
    g1867_p_spl_,
    g1867_p
  );


  buf

  (
    g1857_p_spl_,
    g1857_p
  );


  buf

  (
    g1867_n_spl_,
    g1867_n
  );


  buf

  (
    g1868_n_spl_,
    g1868_n
  );


  buf

  (
    g1868_p_spl_,
    g1868_p
  );


  buf

  (
    g1856_n_spl_,
    g1856_n
  );


  buf

  (
    g1870_p_spl_,
    g1870_p
  );


  buf

  (
    g1856_p_spl_,
    g1856_p
  );


  buf

  (
    g1870_n_spl_,
    g1870_n
  );


  buf

  (
    g1871_n_spl_,
    g1871_n
  );


  buf

  (
    g1871_p_spl_,
    g1871_p
  );


  buf

  (
    g1855_n_spl_,
    g1855_n
  );


  buf

  (
    g1873_p_spl_,
    g1873_p
  );


  buf

  (
    g1855_p_spl_,
    g1855_p
  );


  buf

  (
    g1873_n_spl_,
    g1873_n
  );


  buf

  (
    g1874_p_spl_,
    g1874_p
  );


  buf

  (
    g1854_n_spl_,
    g1854_n
  );


  buf

  (
    g1876_p_spl_,
    g1876_p
  );


  buf

  (
    g1853_n_spl_,
    g1853_n
  );


  buf

  (
    g1879_p_spl_,
    g1879_p
  );


  buf

  (
    g1886_n_spl_,
    g1886_n
  );


  buf

  (
    g1888_p_spl_,
    g1888_p
  );


  buf

  (
    g1886_p_spl_,
    g1886_p
  );


  buf

  (
    g1888_n_spl_,
    g1888_n
  );


  buf

  (
    g1889_n_spl_,
    g1889_n
  );


  buf

  (
    g1889_p_spl_,
    g1889_p
  );


  buf

  (
    g1885_n_spl_,
    g1885_n
  );


  buf

  (
    g1891_p_spl_,
    g1891_p
  );


  buf

  (
    g1885_p_spl_,
    g1885_p
  );


  buf

  (
    g1891_n_spl_,
    g1891_n
  );


  buf

  (
    g1892_n_spl_,
    g1892_n
  );


  buf

  (
    g1892_p_spl_,
    g1892_p
  );


  buf

  (
    g1884_n_spl_,
    g1884_n
  );


  buf

  (
    g1894_p_spl_,
    g1894_p
  );


  buf

  (
    g1884_p_spl_,
    g1884_p
  );


  buf

  (
    g1894_n_spl_,
    g1894_n
  );


  buf

  (
    g1895_p_spl_,
    g1895_p
  );


  buf

  (
    g1883_n_spl_,
    g1883_n
  );


  buf

  (
    g1897_p_spl_,
    g1897_p
  );


  buf

  (
    g1882_n_spl_,
    g1882_n
  );


  buf

  (
    g1900_p_spl_,
    g1900_p
  );


  buf

  (
    g1905_n_spl_,
    g1905_n
  );


  buf

  (
    g1907_p_spl_,
    g1907_p
  );


  buf

  (
    g1905_p_spl_,
    g1905_p
  );


  buf

  (
    g1907_n_spl_,
    g1907_n
  );


  buf

  (
    g1908_p_spl_,
    g1908_p
  );


  buf

  (
    g1904_n_spl_,
    g1904_n
  );


  buf

  (
    g1910_p_spl_,
    g1910_p
  );


  buf

  (
    g1903_n_spl_,
    g1903_n
  );


  buf

  (
    g1913_p_spl_,
    g1913_p
  );


  buf

  (
    g1519_n_spl_,
    g1519_n
  );


  buf

  (
    g1916_n_spl_,
    g1916_n
  );


  buf

  (
    g1918_p_spl_,
    g1918_p
  );


  buf

  (
    g1921_p_spl_,
    g1921_p
  );


  buf

  (
    g1923_n_spl_,
    g1923_n
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G5_p_spl_0,
    G5_p_spl_
  );


  buf

  (
    G5_p_spl_00,
    G5_p_spl_0
  );


  buf

  (
    G5_p_spl_01,
    G5_p_spl_0
  );


  buf

  (
    G5_p_spl_1,
    G5_p_spl_
  );


  buf

  (
    G5_n_spl_,
    G5_n
  );


  buf

  (
    G5_n_spl_0,
    G5_n_spl_
  );


  buf

  (
    G5_n_spl_1,
    G5_n_spl_
  );


  buf

  (
    g1926_p_spl_,
    g1926_p
  );


  buf

  (
    g1927_p_spl_,
    g1927_p
  );


  buf

  (
    g1926_n_spl_,
    g1926_n
  );


  buf

  (
    g1927_n_spl_,
    g1927_n
  );


  buf

  (
    g1928_n_spl_,
    g1928_n
  );


  buf

  (
    g1928_n_spl_0,
    g1928_n_spl_
  );


  buf

  (
    g1928_p_spl_,
    g1928_p
  );


  buf

  (
    g1928_p_spl_0,
    g1928_p_spl_
  );


  buf

  (
    g1930_n_spl_,
    g1930_n
  );


  buf

  (
    g1930_p_spl_,
    g1930_p
  );


  buf

  (
    g1931_n_spl_,
    g1931_n
  );


  buf

  (
    g1931_p_spl_,
    g1931_p
  );


  buf

  (
    g1932_n_spl_,
    g1932_n
  );


  buf

  (
    g1934_p_spl_,
    g1934_p
  );


  buf

  (
    g1932_p_spl_,
    g1932_p
  );


  buf

  (
    g1934_n_spl_,
    g1934_n
  );


  buf

  (
    g1935_n_spl_,
    g1935_n
  );


  buf

  (
    g1935_p_spl_,
    g1935_p
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G6_p_spl_0,
    G6_p_spl_
  );


  buf

  (
    G6_p_spl_00,
    G6_p_spl_0
  );


  buf

  (
    G6_p_spl_01,
    G6_p_spl_0
  );


  buf

  (
    G6_p_spl_1,
    G6_p_spl_
  );


  buf

  (
    G6_n_spl_,
    G6_n
  );


  buf

  (
    G6_n_spl_0,
    G6_n_spl_
  );


  buf

  (
    G6_n_spl_1,
    G6_n_spl_
  );


  buf

  (
    g1938_p_spl_,
    g1938_p
  );


  buf

  (
    g1939_p_spl_,
    g1939_p
  );


  buf

  (
    g1938_n_spl_,
    g1938_n
  );


  buf

  (
    g1939_n_spl_,
    g1939_n
  );


  buf

  (
    g1940_n_spl_,
    g1940_n
  );


  buf

  (
    g1940_n_spl_0,
    g1940_n_spl_
  );


  buf

  (
    g1940_p_spl_,
    g1940_p
  );


  buf

  (
    g1940_p_spl_0,
    g1940_p_spl_
  );


  buf

  (
    g1942_n_spl_,
    g1942_n
  );


  buf

  (
    g1942_p_spl_,
    g1942_p
  );


  buf

  (
    g1943_n_spl_,
    g1943_n
  );


  buf

  (
    g1943_p_spl_,
    g1943_p
  );


  buf

  (
    g1937_n_spl_,
    g1937_n
  );


  buf

  (
    g1945_p_spl_,
    g1945_p
  );


  buf

  (
    g1937_p_spl_,
    g1937_p
  );


  buf

  (
    g1945_n_spl_,
    g1945_n
  );


  buf

  (
    g1946_n_spl_,
    g1946_n
  );


  buf

  (
    g1946_p_spl_,
    g1946_p
  );


  buf

  (
    g1936_n_spl_,
    g1936_n
  );


  buf

  (
    g1948_p_spl_,
    g1948_p
  );


  buf

  (
    g1936_p_spl_,
    g1936_p
  );


  buf

  (
    g1948_n_spl_,
    g1948_n
  );


  buf

  (
    G20_p_spl_,
    G20_p
  );


  buf

  (
    G20_p_spl_0,
    G20_p_spl_
  );


  buf

  (
    G20_p_spl_00,
    G20_p_spl_0
  );


  buf

  (
    G20_p_spl_000,
    G20_p_spl_00
  );


  buf

  (
    G20_p_spl_001,
    G20_p_spl_00
  );


  buf

  (
    G20_p_spl_01,
    G20_p_spl_0
  );


  buf

  (
    G20_p_spl_010,
    G20_p_spl_01
  );


  buf

  (
    G20_p_spl_011,
    G20_p_spl_01
  );


  buf

  (
    G20_p_spl_1,
    G20_p_spl_
  );


  buf

  (
    G20_p_spl_10,
    G20_p_spl_1
  );


  buf

  (
    G20_p_spl_100,
    G20_p_spl_10
  );


  buf

  (
    G20_p_spl_101,
    G20_p_spl_10
  );


  buf

  (
    G20_p_spl_11,
    G20_p_spl_1
  );


  buf

  (
    G20_p_spl_110,
    G20_p_spl_11
  );


  buf

  (
    g1949_n_spl_,
    g1949_n
  );


  buf

  (
    g1949_p_spl_,
    g1949_p
  );


  buf

  (
    g1950_n_spl_,
    g1950_n
  );


  buf

  (
    g1952_p_spl_,
    g1952_p
  );


  buf

  (
    g1950_p_spl_,
    g1950_p
  );


  buf

  (
    g1952_n_spl_,
    g1952_n
  );


  buf

  (
    g1953_n_spl_,
    g1953_n
  );


  buf

  (
    g1953_p_spl_,
    g1953_p
  );


  buf

  (
    G7_p_spl_,
    G7_p
  );


  buf

  (
    G7_p_spl_0,
    G7_p_spl_
  );


  buf

  (
    G7_p_spl_00,
    G7_p_spl_0
  );


  buf

  (
    G7_p_spl_01,
    G7_p_spl_0
  );


  buf

  (
    G7_p_spl_1,
    G7_p_spl_
  );


  buf

  (
    G7_n_spl_,
    G7_n
  );


  buf

  (
    G7_n_spl_0,
    G7_n_spl_
  );


  buf

  (
    G7_n_spl_1,
    G7_n_spl_
  );


  buf

  (
    g1958_p_spl_,
    g1958_p
  );


  buf

  (
    g1959_p_spl_,
    g1959_p
  );


  buf

  (
    g1958_n_spl_,
    g1958_n
  );


  buf

  (
    g1959_n_spl_,
    g1959_n
  );


  buf

  (
    g1960_n_spl_,
    g1960_n
  );


  buf

  (
    g1960_n_spl_0,
    g1960_n_spl_
  );


  buf

  (
    g1960_p_spl_,
    g1960_p
  );


  buf

  (
    g1960_p_spl_0,
    g1960_p_spl_
  );


  buf

  (
    g1962_n_spl_,
    g1962_n
  );


  buf

  (
    g1962_p_spl_,
    g1962_p
  );


  buf

  (
    g1963_n_spl_,
    g1963_n
  );


  buf

  (
    g1963_p_spl_,
    g1963_p
  );


  buf

  (
    g1957_n_spl_,
    g1957_n
  );


  buf

  (
    g1965_p_spl_,
    g1965_p
  );


  buf

  (
    g1957_p_spl_,
    g1957_p
  );


  buf

  (
    g1965_n_spl_,
    g1965_n
  );


  buf

  (
    g1966_n_spl_,
    g1966_n
  );


  buf

  (
    g1966_p_spl_,
    g1966_p
  );


  buf

  (
    g1956_n_spl_,
    g1956_n
  );


  buf

  (
    g1968_p_spl_,
    g1968_p
  );


  buf

  (
    g1956_p_spl_,
    g1956_p
  );


  buf

  (
    g1968_n_spl_,
    g1968_n
  );


  buf

  (
    g1969_n_spl_,
    g1969_n
  );


  buf

  (
    g1969_p_spl_,
    g1969_p
  );


  buf

  (
    g1955_n_spl_,
    g1955_n
  );


  buf

  (
    g1971_p_spl_,
    g1971_p
  );


  buf

  (
    g1955_p_spl_,
    g1955_p
  );


  buf

  (
    g1971_n_spl_,
    g1971_n
  );


  buf

  (
    g1972_n_spl_,
    g1972_n
  );


  buf

  (
    g1972_p_spl_,
    g1972_p
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_00,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_01,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_1,
    G8_p_spl_
  );


  buf

  (
    G8_n_spl_,
    G8_n
  );


  buf

  (
    G8_n_spl_0,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_1,
    G8_n_spl_
  );


  buf

  (
    g1980_p_spl_,
    g1980_p
  );


  buf

  (
    g1981_p_spl_,
    g1981_p
  );


  buf

  (
    g1980_n_spl_,
    g1980_n
  );


  buf

  (
    g1981_n_spl_,
    g1981_n
  );


  buf

  (
    g1982_n_spl_,
    g1982_n
  );


  buf

  (
    g1982_n_spl_0,
    g1982_n_spl_
  );


  buf

  (
    g1982_p_spl_,
    g1982_p
  );


  buf

  (
    g1982_p_spl_0,
    g1982_p_spl_
  );


  buf

  (
    g1984_n_spl_,
    g1984_n
  );


  buf

  (
    g1984_p_spl_,
    g1984_p
  );


  buf

  (
    g1985_n_spl_,
    g1985_n
  );


  buf

  (
    g1985_p_spl_,
    g1985_p
  );


  buf

  (
    g1979_n_spl_,
    g1979_n
  );


  buf

  (
    g1987_p_spl_,
    g1987_p
  );


  buf

  (
    g1979_p_spl_,
    g1979_p
  );


  buf

  (
    g1987_n_spl_,
    g1987_n
  );


  buf

  (
    g1988_n_spl_,
    g1988_n
  );


  buf

  (
    g1988_p_spl_,
    g1988_p
  );


  buf

  (
    g1978_n_spl_,
    g1978_n
  );


  buf

  (
    g1990_p_spl_,
    g1990_p
  );


  buf

  (
    g1978_p_spl_,
    g1978_p
  );


  buf

  (
    g1990_n_spl_,
    g1990_n
  );


  buf

  (
    g1991_n_spl_,
    g1991_n
  );


  buf

  (
    g1991_p_spl_,
    g1991_p
  );


  buf

  (
    g1977_n_spl_,
    g1977_n
  );


  buf

  (
    g1993_p_spl_,
    g1993_p
  );


  buf

  (
    g1977_p_spl_,
    g1977_p
  );


  buf

  (
    g1993_n_spl_,
    g1993_n
  );


  buf

  (
    g1994_n_spl_,
    g1994_n
  );


  buf

  (
    g1994_p_spl_,
    g1994_p
  );


  buf

  (
    G9_p_spl_,
    G9_p
  );


  buf

  (
    G9_p_spl_0,
    G9_p_spl_
  );


  buf

  (
    G9_p_spl_00,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_01,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_1,
    G9_p_spl_
  );


  buf

  (
    G9_n_spl_,
    G9_n
  );


  buf

  (
    G9_n_spl_0,
    G9_n_spl_
  );


  buf

  (
    G9_n_spl_1,
    G9_n_spl_
  );


  buf

  (
    g2002_p_spl_,
    g2002_p
  );


  buf

  (
    g2003_p_spl_,
    g2003_p
  );


  buf

  (
    g2002_n_spl_,
    g2002_n
  );


  buf

  (
    g2003_n_spl_,
    g2003_n
  );


  buf

  (
    g2004_n_spl_,
    g2004_n
  );


  buf

  (
    g2004_n_spl_0,
    g2004_n_spl_
  );


  buf

  (
    g2004_p_spl_,
    g2004_p
  );


  buf

  (
    g2004_p_spl_0,
    g2004_p_spl_
  );


  buf

  (
    g2006_n_spl_,
    g2006_n
  );


  buf

  (
    g2006_p_spl_,
    g2006_p
  );


  buf

  (
    g2007_n_spl_,
    g2007_n
  );


  buf

  (
    g2007_p_spl_,
    g2007_p
  );


  buf

  (
    g2001_n_spl_,
    g2001_n
  );


  buf

  (
    g2009_p_spl_,
    g2009_p
  );


  buf

  (
    g2001_p_spl_,
    g2001_p
  );


  buf

  (
    g2009_n_spl_,
    g2009_n
  );


  buf

  (
    g2010_n_spl_,
    g2010_n
  );


  buf

  (
    g2010_p_spl_,
    g2010_p
  );


  buf

  (
    g2000_n_spl_,
    g2000_n
  );


  buf

  (
    g2012_p_spl_,
    g2012_p
  );


  buf

  (
    g2000_p_spl_,
    g2000_p
  );


  buf

  (
    g2012_n_spl_,
    g2012_n
  );


  buf

  (
    g2013_n_spl_,
    g2013_n
  );


  buf

  (
    g2013_p_spl_,
    g2013_p
  );


  buf

  (
    g1999_n_spl_,
    g1999_n
  );


  buf

  (
    g2015_p_spl_,
    g2015_p
  );


  buf

  (
    g1999_p_spl_,
    g1999_p
  );


  buf

  (
    g2015_n_spl_,
    g2015_n
  );


  buf

  (
    g2016_n_spl_,
    g2016_n
  );


  buf

  (
    g2016_p_spl_,
    g2016_p
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


  buf

  (
    G10_p_spl_0,
    G10_p_spl_
  );


  buf

  (
    G10_p_spl_00,
    G10_p_spl_0
  );


  buf

  (
    G10_p_spl_01,
    G10_p_spl_0
  );


  buf

  (
    G10_p_spl_1,
    G10_p_spl_
  );


  buf

  (
    G10_n_spl_,
    G10_n
  );


  buf

  (
    G10_n_spl_0,
    G10_n_spl_
  );


  buf

  (
    G10_n_spl_1,
    G10_n_spl_
  );


  buf

  (
    g2024_p_spl_,
    g2024_p
  );


  buf

  (
    g2025_p_spl_,
    g2025_p
  );


  buf

  (
    g2024_n_spl_,
    g2024_n
  );


  buf

  (
    g2025_n_spl_,
    g2025_n
  );


  buf

  (
    g2026_n_spl_,
    g2026_n
  );


  buf

  (
    g2026_n_spl_0,
    g2026_n_spl_
  );


  buf

  (
    g2026_p_spl_,
    g2026_p
  );


  buf

  (
    g2026_p_spl_0,
    g2026_p_spl_
  );


  buf

  (
    g2028_n_spl_,
    g2028_n
  );


  buf

  (
    g2028_p_spl_,
    g2028_p
  );


  buf

  (
    g2029_n_spl_,
    g2029_n
  );


  buf

  (
    g2029_p_spl_,
    g2029_p
  );


  buf

  (
    g2023_n_spl_,
    g2023_n
  );


  buf

  (
    g2031_p_spl_,
    g2031_p
  );


  buf

  (
    g2023_p_spl_,
    g2023_p
  );


  buf

  (
    g2031_n_spl_,
    g2031_n
  );


  buf

  (
    g2032_n_spl_,
    g2032_n
  );


  buf

  (
    g2032_p_spl_,
    g2032_p
  );


  buf

  (
    g2022_n_spl_,
    g2022_n
  );


  buf

  (
    g2034_p_spl_,
    g2034_p
  );


  buf

  (
    g2022_p_spl_,
    g2022_p
  );


  buf

  (
    g2034_n_spl_,
    g2034_n
  );


  buf

  (
    g2035_n_spl_,
    g2035_n
  );


  buf

  (
    g2035_p_spl_,
    g2035_p
  );


  buf

  (
    g2021_n_spl_,
    g2021_n
  );


  buf

  (
    g2037_p_spl_,
    g2037_p
  );


  buf

  (
    g2021_p_spl_,
    g2021_p
  );


  buf

  (
    g2037_n_spl_,
    g2037_n
  );


  buf

  (
    g2038_n_spl_,
    g2038_n
  );


  buf

  (
    g2038_p_spl_,
    g2038_p
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    G11_p_spl_0,
    G11_p_spl_
  );


  buf

  (
    G11_p_spl_00,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_01,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_1,
    G11_p_spl_
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    G11_n_spl_0,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_1,
    G11_n_spl_
  );


  buf

  (
    g2046_p_spl_,
    g2046_p
  );


  buf

  (
    g2047_p_spl_,
    g2047_p
  );


  buf

  (
    g2046_n_spl_,
    g2046_n
  );


  buf

  (
    g2047_n_spl_,
    g2047_n
  );


  buf

  (
    g2048_n_spl_,
    g2048_n
  );


  buf

  (
    g2048_n_spl_0,
    g2048_n_spl_
  );


  buf

  (
    g2048_p_spl_,
    g2048_p
  );


  buf

  (
    g2048_p_spl_0,
    g2048_p_spl_
  );


  buf

  (
    g2050_n_spl_,
    g2050_n
  );


  buf

  (
    g2050_p_spl_,
    g2050_p
  );


  buf

  (
    g2051_n_spl_,
    g2051_n
  );


  buf

  (
    g2051_p_spl_,
    g2051_p
  );


  buf

  (
    g2045_n_spl_,
    g2045_n
  );


  buf

  (
    g2053_p_spl_,
    g2053_p
  );


  buf

  (
    g2045_p_spl_,
    g2045_p
  );


  buf

  (
    g2053_n_spl_,
    g2053_n
  );


  buf

  (
    g2054_n_spl_,
    g2054_n
  );


  buf

  (
    g2054_p_spl_,
    g2054_p
  );


  buf

  (
    g2044_n_spl_,
    g2044_n
  );


  buf

  (
    g2056_p_spl_,
    g2056_p
  );


  buf

  (
    g2044_p_spl_,
    g2044_p
  );


  buf

  (
    g2056_n_spl_,
    g2056_n
  );


  buf

  (
    g2057_n_spl_,
    g2057_n
  );


  buf

  (
    g2057_p_spl_,
    g2057_p
  );


  buf

  (
    g2043_n_spl_,
    g2043_n
  );


  buf

  (
    g2059_p_spl_,
    g2059_p
  );


  buf

  (
    g2043_p_spl_,
    g2043_p
  );


  buf

  (
    g2059_n_spl_,
    g2059_n
  );


  buf

  (
    g2060_n_spl_,
    g2060_n
  );


  buf

  (
    g2060_p_spl_,
    g2060_p
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_00,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_01,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_1,
    G12_p_spl_
  );


  buf

  (
    G12_n_spl_,
    G12_n
  );


  buf

  (
    G12_n_spl_0,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_1,
    G12_n_spl_
  );


  buf

  (
    g2068_p_spl_,
    g2068_p
  );


  buf

  (
    g2069_p_spl_,
    g2069_p
  );


  buf

  (
    g2068_n_spl_,
    g2068_n
  );


  buf

  (
    g2069_n_spl_,
    g2069_n
  );


  buf

  (
    g2070_n_spl_,
    g2070_n
  );


  buf

  (
    g2070_n_spl_0,
    g2070_n_spl_
  );


  buf

  (
    g2070_p_spl_,
    g2070_p
  );


  buf

  (
    g2070_p_spl_0,
    g2070_p_spl_
  );


  buf

  (
    g2072_n_spl_,
    g2072_n
  );


  buf

  (
    g2072_p_spl_,
    g2072_p
  );


  buf

  (
    g2073_n_spl_,
    g2073_n
  );


  buf

  (
    g2073_p_spl_,
    g2073_p
  );


  buf

  (
    g2067_n_spl_,
    g2067_n
  );


  buf

  (
    g2075_p_spl_,
    g2075_p
  );


  buf

  (
    g2067_p_spl_,
    g2067_p
  );


  buf

  (
    g2075_n_spl_,
    g2075_n
  );


  buf

  (
    g2076_n_spl_,
    g2076_n
  );


  buf

  (
    g2076_p_spl_,
    g2076_p
  );


  buf

  (
    g2066_n_spl_,
    g2066_n
  );


  buf

  (
    g2078_p_spl_,
    g2078_p
  );


  buf

  (
    g2066_p_spl_,
    g2066_p
  );


  buf

  (
    g2078_n_spl_,
    g2078_n
  );


  buf

  (
    g2079_n_spl_,
    g2079_n
  );


  buf

  (
    g2079_p_spl_,
    g2079_p
  );


  buf

  (
    g2065_n_spl_,
    g2065_n
  );


  buf

  (
    g2081_p_spl_,
    g2081_p
  );


  buf

  (
    g2065_p_spl_,
    g2065_p
  );


  buf

  (
    g2081_n_spl_,
    g2081_n
  );


  buf

  (
    g2082_n_spl_,
    g2082_n
  );


  buf

  (
    g2082_p_spl_,
    g2082_p
  );


  buf

  (
    G13_p_spl_,
    G13_p
  );


  buf

  (
    G13_p_spl_0,
    G13_p_spl_
  );


  buf

  (
    G13_p_spl_00,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_01,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_1,
    G13_p_spl_
  );


  buf

  (
    G13_n_spl_,
    G13_n
  );


  buf

  (
    G13_n_spl_0,
    G13_n_spl_
  );


  buf

  (
    G13_n_spl_1,
    G13_n_spl_
  );


  buf

  (
    g2090_p_spl_,
    g2090_p
  );


  buf

  (
    g2091_p_spl_,
    g2091_p
  );


  buf

  (
    g2090_n_spl_,
    g2090_n
  );


  buf

  (
    g2091_n_spl_,
    g2091_n
  );


  buf

  (
    g2092_n_spl_,
    g2092_n
  );


  buf

  (
    g2092_n_spl_0,
    g2092_n_spl_
  );


  buf

  (
    g2092_p_spl_,
    g2092_p
  );


  buf

  (
    g2092_p_spl_0,
    g2092_p_spl_
  );


  buf

  (
    g2094_n_spl_,
    g2094_n
  );


  buf

  (
    g2094_p_spl_,
    g2094_p
  );


  buf

  (
    g2095_n_spl_,
    g2095_n
  );


  buf

  (
    g2095_p_spl_,
    g2095_p
  );


  buf

  (
    g2089_n_spl_,
    g2089_n
  );


  buf

  (
    g2097_p_spl_,
    g2097_p
  );


  buf

  (
    g2089_p_spl_,
    g2089_p
  );


  buf

  (
    g2097_n_spl_,
    g2097_n
  );


  buf

  (
    g2098_n_spl_,
    g2098_n
  );


  buf

  (
    g2098_p_spl_,
    g2098_p
  );


  buf

  (
    g2088_n_spl_,
    g2088_n
  );


  buf

  (
    g2100_p_spl_,
    g2100_p
  );


  buf

  (
    g2088_p_spl_,
    g2088_p
  );


  buf

  (
    g2100_n_spl_,
    g2100_n
  );


  buf

  (
    g2101_n_spl_,
    g2101_n
  );


  buf

  (
    g2101_p_spl_,
    g2101_p
  );


  buf

  (
    g2087_n_spl_,
    g2087_n
  );


  buf

  (
    g2103_p_spl_,
    g2103_p
  );


  buf

  (
    g2087_p_spl_,
    g2087_p
  );


  buf

  (
    g2103_n_spl_,
    g2103_n
  );


  buf

  (
    g2104_n_spl_,
    g2104_n
  );


  buf

  (
    g2104_p_spl_,
    g2104_p
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G14_p_spl_0,
    G14_p_spl_
  );


  buf

  (
    G14_p_spl_00,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_01,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_1,
    G14_p_spl_
  );


  buf

  (
    G14_n_spl_,
    G14_n
  );


  buf

  (
    G14_n_spl_0,
    G14_n_spl_
  );


  buf

  (
    G14_n_spl_1,
    G14_n_spl_
  );


  buf

  (
    g2112_p_spl_,
    g2112_p
  );


  buf

  (
    g2113_p_spl_,
    g2113_p
  );


  buf

  (
    g2112_n_spl_,
    g2112_n
  );


  buf

  (
    g2113_n_spl_,
    g2113_n
  );


  buf

  (
    g2114_n_spl_,
    g2114_n
  );


  buf

  (
    g2114_n_spl_0,
    g2114_n_spl_
  );


  buf

  (
    g2114_p_spl_,
    g2114_p
  );


  buf

  (
    g2114_p_spl_0,
    g2114_p_spl_
  );


  buf

  (
    g2116_n_spl_,
    g2116_n
  );


  buf

  (
    g2116_p_spl_,
    g2116_p
  );


  buf

  (
    g2117_n_spl_,
    g2117_n
  );


  buf

  (
    g2117_p_spl_,
    g2117_p
  );


  buf

  (
    g2111_n_spl_,
    g2111_n
  );


  buf

  (
    g2119_p_spl_,
    g2119_p
  );


  buf

  (
    g2111_p_spl_,
    g2111_p
  );


  buf

  (
    g2119_n_spl_,
    g2119_n
  );


  buf

  (
    g2120_n_spl_,
    g2120_n
  );


  buf

  (
    g2120_p_spl_,
    g2120_p
  );


  buf

  (
    g2110_n_spl_,
    g2110_n
  );


  buf

  (
    g2122_p_spl_,
    g2122_p
  );


  buf

  (
    g2110_p_spl_,
    g2110_p
  );


  buf

  (
    g2122_n_spl_,
    g2122_n
  );


  buf

  (
    g2123_n_spl_,
    g2123_n
  );


  buf

  (
    g2123_p_spl_,
    g2123_p
  );


  buf

  (
    g2109_n_spl_,
    g2109_n
  );


  buf

  (
    g2125_p_spl_,
    g2125_p
  );


  buf

  (
    g2109_p_spl_,
    g2109_p
  );


  buf

  (
    g2125_n_spl_,
    g2125_n
  );


  buf

  (
    g2126_n_spl_,
    g2126_n
  );


  buf

  (
    g2126_p_spl_,
    g2126_p
  );


  buf

  (
    G15_p_spl_,
    G15_p
  );


  buf

  (
    G15_p_spl_0,
    G15_p_spl_
  );


  buf

  (
    G15_p_spl_00,
    G15_p_spl_0
  );


  buf

  (
    G15_p_spl_1,
    G15_p_spl_
  );


  buf

  (
    G15_n_spl_,
    G15_n
  );


  buf

  (
    G15_n_spl_0,
    G15_n_spl_
  );


  buf

  (
    G15_n_spl_1,
    G15_n_spl_
  );


  buf

  (
    g2134_p_spl_,
    g2134_p
  );


  buf

  (
    g2135_p_spl_,
    g2135_p
  );


  buf

  (
    g2134_n_spl_,
    g2134_n
  );


  buf

  (
    g2135_n_spl_,
    g2135_n
  );


  buf

  (
    g2136_n_spl_,
    g2136_n
  );


  buf

  (
    g2136_n_spl_0,
    g2136_n_spl_
  );


  buf

  (
    g2136_p_spl_,
    g2136_p
  );


  buf

  (
    g2136_p_spl_0,
    g2136_p_spl_
  );


  buf

  (
    g2138_n_spl_,
    g2138_n
  );


  buf

  (
    g2138_p_spl_,
    g2138_p
  );


  buf

  (
    g2139_n_spl_,
    g2139_n
  );


  buf

  (
    g2139_p_spl_,
    g2139_p
  );


  buf

  (
    g2133_n_spl_,
    g2133_n
  );


  buf

  (
    g2141_p_spl_,
    g2141_p
  );


  buf

  (
    g2133_p_spl_,
    g2133_p
  );


  buf

  (
    g2141_n_spl_,
    g2141_n
  );


  buf

  (
    g2142_n_spl_,
    g2142_n
  );


  buf

  (
    g2142_p_spl_,
    g2142_p
  );


  buf

  (
    g2132_n_spl_,
    g2132_n
  );


  buf

  (
    g2144_p_spl_,
    g2144_p
  );


  buf

  (
    g2132_p_spl_,
    g2132_p
  );


  buf

  (
    g2144_n_spl_,
    g2144_n
  );


  buf

  (
    g2145_n_spl_,
    g2145_n
  );


  buf

  (
    g2145_p_spl_,
    g2145_p
  );


  buf

  (
    g2131_n_spl_,
    g2131_n
  );


  buf

  (
    g2147_p_spl_,
    g2147_p
  );


  buf

  (
    g2131_p_spl_,
    g2131_p
  );


  buf

  (
    g2147_n_spl_,
    g2147_n
  );


  buf

  (
    g2148_n_spl_,
    g2148_n
  );


  buf

  (
    g2148_p_spl_,
    g2148_p
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    G16_p_spl_0,
    G16_p_spl_
  );


  buf

  (
    G16_p_spl_00,
    G16_p_spl_0
  );


  buf

  (
    G16_p_spl_1,
    G16_p_spl_
  );


  buf

  (
    G16_n_spl_,
    G16_n
  );


  buf

  (
    G16_n_spl_0,
    G16_n_spl_
  );


  buf

  (
    g2156_p_spl_,
    g2156_p
  );


  buf

  (
    g2157_p_spl_,
    g2157_p
  );


  buf

  (
    g2156_n_spl_,
    g2156_n
  );


  buf

  (
    g2157_n_spl_,
    g2157_n
  );


  buf

  (
    g2158_n_spl_,
    g2158_n
  );


  buf

  (
    g2158_p_spl_,
    g2158_p
  );


  buf

  (
    g2160_n_spl_,
    g2160_n
  );


  buf

  (
    g2160_p_spl_,
    g2160_p
  );


  buf

  (
    g2161_n_spl_,
    g2161_n
  );


  buf

  (
    g2161_p_spl_,
    g2161_p
  );


  buf

  (
    g2155_n_spl_,
    g2155_n
  );


  buf

  (
    g2163_p_spl_,
    g2163_p
  );


  buf

  (
    g2155_p_spl_,
    g2155_p
  );


  buf

  (
    g2163_n_spl_,
    g2163_n
  );


  buf

  (
    g2164_n_spl_,
    g2164_n
  );


  buf

  (
    g2164_p_spl_,
    g2164_p
  );


  buf

  (
    g2154_n_spl_,
    g2154_n
  );


  buf

  (
    g2166_p_spl_,
    g2166_p
  );


  buf

  (
    g2154_p_spl_,
    g2154_p
  );


  buf

  (
    g2166_n_spl_,
    g2166_n
  );


  buf

  (
    g2167_n_spl_,
    g2167_n
  );


  buf

  (
    g2167_p_spl_,
    g2167_p
  );


  buf

  (
    g2153_n_spl_,
    g2153_n
  );


  buf

  (
    g2169_p_spl_,
    g2169_p
  );


  buf

  (
    g2153_p_spl_,
    g2153_p
  );


  buf

  (
    g2169_n_spl_,
    g2169_n
  );


  buf

  (
    g2170_n_spl_,
    g2170_n
  );


  buf

  (
    g2170_p_spl_,
    g2170_p
  );


  buf

  (
    g2177_p_spl_,
    g2177_p
  );


  buf

  (
    g2177_n_spl_,
    g2177_n
  );


  buf

  (
    g2178_p_spl_,
    g2178_p
  );


  buf

  (
    g2179_n_spl_,
    g2179_n
  );


  buf

  (
    g2178_n_spl_,
    g2178_n
  );


  buf

  (
    g2179_p_spl_,
    g2179_p
  );


  buf

  (
    g2180_n_spl_,
    g2180_n
  );


  buf

  (
    g2180_p_spl_,
    g2180_p
  );


  buf

  (
    g2176_n_spl_,
    g2176_n
  );


  buf

  (
    g2182_p_spl_,
    g2182_p
  );


  buf

  (
    g2176_p_spl_,
    g2176_p
  );


  buf

  (
    g2182_n_spl_,
    g2182_n
  );


  buf

  (
    g2183_n_spl_,
    g2183_n
  );


  buf

  (
    g2183_p_spl_,
    g2183_p
  );


  buf

  (
    g2175_n_spl_,
    g2175_n
  );


  buf

  (
    g2185_p_spl_,
    g2185_p
  );


  buf

  (
    g2175_p_spl_,
    g2175_p
  );


  buf

  (
    g2185_n_spl_,
    g2185_n
  );


  buf

  (
    g2186_n_spl_,
    g2186_n
  );


  buf

  (
    g2186_p_spl_,
    g2186_p
  );


  buf

  (
    g2192_n_spl_,
    g2192_n
  );


  buf

  (
    g2193_n_spl_,
    g2193_n
  );


  buf

  (
    g2192_p_spl_,
    g2192_p
  );


  buf

  (
    g2193_p_spl_,
    g2193_p
  );


  buf

  (
    g2194_n_spl_,
    g2194_n
  );


  buf

  (
    g2191_n_spl_,
    g2191_n
  );


  buf

  (
    g2196_p_spl_,
    g2196_p
  );


  buf

  (
    g2191_p_spl_,
    g2191_p
  );


  buf

  (
    g2196_n_spl_,
    g2196_n
  );


  buf

  (
    g2197_n_spl_,
    g2197_n
  );


  buf

  (
    g2201_n_spl_,
    g2201_n
  );


  buf

  (
    g2203_p_spl_,
    g2203_p
  );


  buf

  (
    g2201_p_spl_,
    g2201_p
  );


  buf

  (
    g2203_n_spl_,
    g2203_n
  );


  buf

  (
    g2204_n_spl_,
    g2204_n
  );


  buf

  (
    g2204_p_spl_,
    g2204_p
  );


  buf

  (
    g2205_n_spl_,
    g2205_n
  );


  buf

  (
    g2207_p_spl_,
    g2207_p
  );


  buf

  (
    g2208_n_spl_,
    g2208_n
  );


  buf

  (
    G21_p_spl_,
    G21_p
  );


  buf

  (
    G21_p_spl_0,
    G21_p_spl_
  );


  buf

  (
    G21_p_spl_00,
    G21_p_spl_0
  );


  buf

  (
    G21_p_spl_000,
    G21_p_spl_00
  );


  buf

  (
    G21_p_spl_001,
    G21_p_spl_00
  );


  buf

  (
    G21_p_spl_01,
    G21_p_spl_0
  );


  buf

  (
    G21_p_spl_010,
    G21_p_spl_01
  );


  buf

  (
    G21_p_spl_011,
    G21_p_spl_01
  );


  buf

  (
    G21_p_spl_1,
    G21_p_spl_
  );


  buf

  (
    G21_p_spl_10,
    G21_p_spl_1
  );


  buf

  (
    G21_p_spl_100,
    G21_p_spl_10
  );


  buf

  (
    G21_p_spl_101,
    G21_p_spl_10
  );


  buf

  (
    G21_p_spl_11,
    G21_p_spl_1
  );


  buf

  (
    g1631_p_spl_,
    g1631_p
  );


  buf

  (
    g2228_n_spl_,
    g2228_n
  );


  buf

  (
    g2230_p_spl_,
    g2230_p
  );


  buf

  (
    g1975_n_spl_,
    g1975_n
  );


  buf

  (
    g1997_n_spl_,
    g1997_n
  );


  buf

  (
    g2019_n_spl_,
    g2019_n
  );


  buf

  (
    g2041_n_spl_,
    g2041_n
  );


  buf

  (
    g2063_n_spl_,
    g2063_n
  );


  buf

  (
    g2085_n_spl_,
    g2085_n
  );


  buf

  (
    g2107_n_spl_,
    g2107_n
  );


  buf

  (
    g2129_n_spl_,
    g2129_n
  );


  buf

  (
    g2151_n_spl_,
    g2151_n
  );


  buf

  (
    g2173_n_spl_,
    g2173_n
  );


  buf

  (
    g2189_n_spl_,
    g2189_n
  );


  buf

  (
    g2200_n_spl_,
    g2200_n
  );


  buf

  (
    g2212_n_spl_,
    g2212_n
  );


endmodule
