// Benchmark "mymod" written by ABC on Sun Oct 29 23:44:41 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41,
    G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
    G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
    G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
    G1354, G1355  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
    G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
    G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
    G1354, G1355;
  reg n621_lo, n630_lo, n633_lo, n642_lo, n645_lo, n654_lo, n657_lo,
    n666_lo, n669_lo, n678_lo, n681_lo, n690_lo, n693_lo, n702_lo, n705_lo,
    n714_lo, n717_lo, n726_lo, n729_lo, n738_lo, n741_lo, n750_lo, n753_lo,
    n762_lo, n765_lo, n774_lo, n777_lo, n786_lo, n789_lo, n798_lo, n801_lo,
    n810_lo, n813_lo, n822_lo, n825_lo, n834_lo, n837_lo, n846_lo, n849_lo,
    n858_lo, n861_lo, n870_lo, n873_lo, n882_lo, n885_lo, n894_lo, n897_lo,
    n906_lo, n909_lo, n918_lo, n921_lo, n930_lo, n933_lo, n942_lo, n945_lo,
    n954_lo, n957_lo, n966_lo, n969_lo, n978_lo, n981_lo, n990_lo, n993_lo,
    n1002_lo, n1005_lo, n1017_lo, n1029_lo, n1041_lo, n1053_lo, n1065_lo,
    n1077_lo, n1089_lo, n1101_lo, n602_o2, n639_o2, n678_o2, n658_o2,
    n783_o2, n802_o2, n726_o2, n763_o2, n1644_o2, n1645_o2, n1646_o2,
    n1647_o2, n1648_o2, n1649_o2, n1650_o2, n1651_o2, n1652_o2, n1653_o2,
    n1654_o2, n1655_o2, n1656_o2, n1657_o2, n1658_o2, n1659_o2, n1660_o2,
    n1661_o2, n1662_o2, n1663_o2, n1664_o2, n1665_o2, n1666_o2, n1667_o2,
    n1668_o2, n1669_o2, n1670_o2, n1671_o2, n1672_o2, n1673_o2, n1674_o2,
    n1675_o2, n685_o2, n680_o2, n822_o2, n843_o2, n842_o2, n681_o2,
    n684_o2, n686_o2, n823_o2, n683_o2, n688_o2, n803_o2, n862_o2, n764_o2,
    n863_o2, n886_o2, lo002_buf_o2, lo006_buf_o2, lo010_buf_o2,
    lo014_buf_o2, lo018_buf_o2, lo022_buf_o2, lo026_buf_o2, lo030_buf_o2,
    lo034_buf_o2, lo038_buf_o2, lo042_buf_o2, lo046_buf_o2, lo050_buf_o2,
    lo054_buf_o2, lo058_buf_o2, lo062_buf_o2, lo066_buf_o2, lo070_buf_o2,
    lo074_buf_o2, lo078_buf_o2, lo082_buf_o2, lo086_buf_o2, lo090_buf_o2,
    lo094_buf_o2, lo098_buf_o2, lo102_buf_o2, lo106_buf_o2, lo110_buf_o2,
    lo114_buf_o2, lo118_buf_o2, lo122_buf_o2, lo126_buf_o2, n600_o2,
    n601_o2, n637_o2, n638_o2, n676_o2, n677_o2, n656_o2, n657_o2, n781_o2,
    n782_o2, n800_o2, n801_o2, n724_o2, n725_o2, n761_o2, n762_o2,
    lo129_buf_o2, lo133_buf_o2, lo137_buf_o2, lo141_buf_o2, lo145_buf_o2,
    lo149_buf_o2, lo153_buf_o2, lo157_buf_o2, lo161_buf_o2, n571_o2,
    n708_o2, n608_o2, n665_o2, n705_o2, n645_o2, n745_o2, n742_o2, n568_o2,
    n717_o2, n605_o2, n662_o2, n714_o2, n642_o2, n754_o2, n751_o2, n584_o2,
    n770_o2, n789_o2, n581_o2, n695_o2, n732_o2, n593_o2, n590_o2, n630_o2,
    n767_o2, n786_o2, n627_o2, n692_o2, n729_o2, n621_o2, n618_o2;
  wire new_new_n510__, new_new_n512__, new_new_n514__, new_new_n516__,
    new_new_n518__, new_new_n520__, new_new_n522__, new_new_n524__,
    new_new_n526__, new_new_n528__, new_new_n530__, new_new_n532__,
    new_new_n534__, new_new_n536__, new_new_n538__, new_new_n540__,
    new_new_n542__, new_new_n544__, new_new_n546__, new_new_n548__,
    new_new_n550__, new_new_n552__, new_new_n554__, new_new_n556__,
    new_new_n558__, new_new_n560__, new_new_n562__, new_new_n564__,
    new_new_n566__, new_new_n568__, new_new_n570__, new_new_n572__,
    new_new_n574__, new_new_n576__, new_new_n578__, new_new_n580__,
    new_new_n582__, new_new_n584__, new_new_n586__, new_new_n588__,
    new_new_n590__, new_new_n592__, new_new_n593__, new_new_n594__,
    new_new_n595__, new_new_n596__, new_new_n597__, new_new_n598__,
    new_new_n599__, new_new_n600__, new_new_n601__, new_new_n602__,
    new_new_n603__, new_new_n604__, new_new_n605__, new_new_n606__,
    new_new_n607__, new_new_n608__, new_new_n609__, new_new_n610__,
    new_new_n611__, new_new_n612__, new_new_n613__, new_new_n614__,
    new_new_n615__, new_new_n616__, new_new_n617__, new_new_n618__,
    new_new_n619__, new_new_n620__, new_new_n621__, new_new_n622__,
    new_new_n623__, new_new_n624__, new_new_n625__, new_new_n626__,
    new_new_n627__, new_new_n628__, new_new_n629__, new_new_n630__,
    new_new_n631__, new_new_n632__, new_new_n633__, new_new_n634__,
    new_new_n635__, new_new_n636__, new_new_n637__, new_new_n638__,
    new_new_n639__, new_new_n640__, new_new_n641__, new_new_n642__,
    new_new_n643__, new_new_n644__, new_new_n645__, new_new_n646__,
    new_new_n647__, new_new_n648__, new_new_n649__, new_new_n650__,
    new_new_n651__, new_new_n652__, new_new_n653__, new_new_n654__,
    new_new_n655__, new_new_n656__, new_new_n657__, new_new_n658__,
    new_new_n659__, new_new_n660__, new_new_n661__, new_new_n662__,
    new_new_n663__, new_new_n664__, new_new_n665__, new_new_n666__,
    new_new_n667__, new_new_n668__, new_new_n669__, new_new_n670__,
    new_new_n671__, new_new_n672__, new_new_n673__, new_new_n674__,
    new_new_n675__, new_new_n676__, new_new_n677__, new_new_n678__,
    new_new_n679__, new_new_n680__, new_new_n681__, new_new_n682__,
    new_new_n683__, new_new_n684__, new_new_n685__, new_new_n686__,
    new_new_n687__, new_new_n688__, new_new_n689__, new_new_n690__,
    new_new_n691__, new_new_n692__, new_new_n693__, new_new_n694__,
    new_new_n695__, new_new_n696__, new_new_n697__, new_new_n698__,
    new_new_n699__, new_new_n700__, new_new_n701__, new_new_n702__,
    new_new_n703__, new_new_n704__, new_new_n705__, new_new_n706__,
    new_new_n707__, new_new_n708__, new_new_n709__, new_new_n710__,
    new_new_n711__, new_new_n712__, new_new_n713__, new_new_n714__,
    new_new_n715__, new_new_n716__, new_new_n717__, new_new_n718__,
    new_new_n719__, new_new_n720__, new_new_n722__, new_new_n724__,
    new_new_n726__, new_new_n728__, new_new_n730__, new_new_n732__,
    new_new_n734__, new_new_n736__, new_new_n738__, new_new_n739__,
    new_new_n740__, new_new_n741__, new_new_n742__, new_new_n743__,
    new_new_n744__, new_new_n745__, new_new_n746__, new_new_n747__,
    new_new_n748__, new_new_n749__, new_new_n750__, new_new_n751__,
    new_new_n752__, new_new_n753__, new_new_n754__, new_new_n756__,
    new_new_n758__, new_new_n760__, new_new_n762__, new_new_n764__,
    new_new_n766__, new_new_n768__, new_new_n770__, new_new_n772__,
    new_new_n774__, new_new_n776__, new_new_n778__, new_new_n780__,
    new_new_n782__, new_new_n784__, new_new_n786__, new_new_n788__,
    new_new_n790__, new_new_n792__, new_new_n794__, new_new_n796__,
    new_new_n798__, new_new_n800__, new_new_n802__, new_new_n804__,
    new_new_n806__, new_new_n808__, new_new_n810__, new_new_n812__,
    new_new_n814__, new_new_n816__, new_new_n818__, new_new_n819__,
    new_new_n820__, new_new_n821__, new_new_n822__, new_new_n823__,
    new_new_n824__, new_new_n825__, new_new_n826__, new_new_n827__,
    new_new_n828__, new_new_n829__, new_new_n830__, new_new_n831__,
    new_new_n832__, new_new_n833__, new_new_n834__, new_new_n835__,
    new_new_n836__, new_new_n837__, new_new_n838__, new_new_n839__,
    new_new_n840__, new_new_n841__, new_new_n842__, new_new_n843__,
    new_new_n844__, new_new_n845__, new_new_n846__, new_new_n847__,
    new_new_n848__, new_new_n849__, new_new_n850__, new_new_n852__,
    new_new_n854__, new_new_n856__, new_new_n858__, new_new_n860__,
    new_new_n862__, new_new_n864__, new_new_n866__, new_new_n868__,
    new_new_n870__, new_new_n872__, new_new_n874__, new_new_n876__,
    new_new_n878__, new_new_n880__, new_new_n882__, new_new_n884__,
    new_new_n886__, new_new_n888__, new_new_n890__, new_new_n892__,
    new_new_n894__, new_new_n896__, new_new_n898__, new_new_n900__,
    new_new_n902__, new_new_n904__, new_new_n906__, new_new_n908__,
    new_new_n910__, new_new_n912__, new_new_n914__, new_new_n915__,
    new_new_n916__, new_new_n917__, new_new_n918__, new_new_n919__,
    new_new_n920__, new_new_n921__, new_new_n922__, new_new_n923__,
    new_new_n924__, new_new_n925__, new_new_n926__, new_new_n927__,
    new_new_n928__, new_new_n929__, new_new_n930__, new_new_n931__,
    new_new_n932__, new_new_n933__, new_new_n934__, new_new_n935__,
    new_new_n936__, new_new_n937__, new_new_n938__, new_new_n939__,
    new_new_n940__, new_new_n941__, new_new_n942__, new_new_n943__,
    new_new_n944__, new_new_n945__, new_new_n946__, new_new_n947__,
    new_new_n948__, new_new_n949__, new_new_n950__, new_new_n951__,
    new_new_n952__, new_new_n953__, new_new_n954__, new_new_n955__,
    new_new_n956__, new_new_n957__, new_new_n958__, new_new_n959__,
    new_new_n960__, new_new_n961__, new_new_n962__, new_new_n963__,
    new_new_n964__, new_new_n965__, new_new_n966__, new_new_n967__,
    new_new_n968__, new_new_n969__, new_new_n970__, new_new_n971__,
    new_new_n972__, new_new_n973__, new_new_n974__, new_new_n975__,
    new_new_n976__, new_new_n977__, new_new_n978__, new_new_n979__,
    new_new_n980__, new_new_n981__, new_new_n982__, new_new_n983__,
    new_new_n984__, new_new_n985__, new_new_n986__, new_new_n987__,
    new_new_n988__, new_new_n989__, new_new_n990__, new_new_n991__,
    new_new_n992__, new_new_n993__, new_new_n994__, new_new_n995__,
    new_new_n996__, new_new_n997__, new_new_n998__, new_new_n999__,
    new_new_n1000__, new_new_n1001__, new_new_n1002__, new_new_n1003__,
    new_new_n1004__, new_new_n1005__, new_new_n1006__, new_new_n1007__,
    new_new_n1008__, new_new_n1009__, new_new_n1010__, new_new_n1011__,
    new_new_n1012__, new_new_n1013__, new_new_n1014__, new_new_n1015__,
    new_new_n1016__, new_new_n1017__, new_new_n1018__, new_new_n1019__,
    new_new_n1020__, new_new_n1021__, new_new_n1022__, new_new_n1023__,
    new_new_n1024__, new_new_n1025__, new_new_n1026__, new_new_n1027__,
    new_new_n1028__, new_new_n1029__, new_new_n1030__, new_new_n1031__,
    new_new_n1032__, new_new_n1033__, new_new_n1034__, new_new_n1035__,
    new_new_n1036__, new_new_n1037__, new_new_n1038__, new_new_n1039__,
    new_new_n1040__, new_new_n1041__, new_new_n1042__, new_new_n1043__,
    new_new_n1044__, new_new_n1045__, new_new_n1046__, new_new_n1047__,
    new_new_n1048__, new_new_n1049__, new_new_n1050__, new_new_n1051__,
    new_new_n1052__, new_new_n1053__, new_new_n1054__, new_new_n1055__,
    new_new_n1056__, new_new_n1057__, new_new_n1058__, new_new_n1059__,
    new_new_n1060__, new_new_n1061__, new_new_n1062__, new_new_n1063__,
    new_new_n1064__, new_new_n1065__, new_new_n1066__, new_new_n1067__,
    new_new_n1068__, new_new_n1069__, new_new_n1070__, new_new_n1071__,
    new_new_n1072__, new_new_n1073__, new_new_n1074__, new_new_n1075__,
    new_new_n1076__, new_new_n1077__, new_new_n1078__, new_new_n1079__,
    new_new_n1080__, new_new_n1081__, new_new_n1082__, new_new_n1083__,
    new_new_n1084__, new_new_n1085__, new_new_n1086__, new_new_n1087__,
    new_new_n1088__, new_new_n1089__, new_new_n1090__, new_new_n1091__,
    new_new_n1092__, new_new_n1093__, new_new_n1094__, new_new_n1095__,
    new_new_n1096__, new_new_n1097__, new_new_n1098__, new_new_n1099__,
    new_new_n1100__, new_new_n1101__, new_new_n1102__, new_new_n1103__,
    new_new_n1104__, new_new_n1105__, new_new_n1106__, new_new_n1107__,
    new_new_n1108__, new_new_n1109__, new_new_n1110__, new_new_n1111__,
    new_new_n1112__, new_new_n1113__, new_new_n1114__, new_new_n1115__,
    new_new_n1116__, new_new_n1117__, new_new_n1118__, new_new_n1119__,
    new_new_n1120__, new_new_n1121__, new_new_n1122__, new_new_n1123__,
    new_new_n1124__, new_new_n1125__, new_new_n1126__, new_new_n1127__,
    new_new_n1128__, new_new_n1129__, new_new_n1130__, new_new_n1131__,
    new_new_n1132__, new_new_n1133__, new_new_n1134__, new_new_n1135__,
    new_new_n1136__, new_new_n1137__, new_new_n1138__, new_new_n1139__,
    new_new_n1140__, new_new_n1141__, new_new_n1142__, new_new_n1143__,
    new_new_n1144__, new_new_n1145__, new_new_n1146__, new_new_n1147__,
    new_new_n1148__, new_new_n1149__, new_new_n1150__, new_new_n1151__,
    new_new_n1152__, new_new_n1153__, new_new_n1154__, new_new_n1155__,
    new_new_n1156__, new_new_n1157__, new_new_n1158__, new_new_n1159__,
    new_new_n1160__, new_new_n1161__, new_new_n1162__, new_new_n1163__,
    new_new_n1164__, new_new_n1165__, new_new_n1166__, new_new_n1167__,
    new_new_n1168__, new_new_n1169__, new_new_n1170__, new_new_n1171__,
    new_new_n1172__, new_new_n1173__, new_new_n1174__, new_new_n1175__,
    new_new_n1176__, new_new_n1177__, new_new_n1178__, new_new_n1179__,
    new_new_n1180__, new_new_n1181__, new_new_n1182__, new_new_n1183__,
    new_new_n1184__, new_new_n1185__, new_new_n1186__, new_new_n1187__,
    new_new_n1188__, new_new_n1189__, new_new_n1190__, new_new_n1191__,
    new_new_n1192__, new_new_n1193__, new_new_n1194__, new_new_n1195__,
    new_new_n1196__, new_new_n1197__, new_new_n1198__, new_new_n1199__,
    new_new_n1200__, new_new_n1201__, new_new_n1202__, new_new_n1203__,
    new_new_n1204__, new_new_n1205__, new_new_n1206__, new_new_n1207__,
    new_new_n1208__, new_new_n1209__, new_new_n1210__, new_new_n1211__,
    new_new_n1212__, new_new_n1213__, new_new_n1214__, new_new_n1215__,
    new_new_n1216__, new_new_n1217__, new_new_n1218__, new_new_n1219__,
    new_new_n1220__, new_new_n1221__, new_new_n1222__, new_new_n1223__,
    new_new_n1224__, new_new_n1225__, new_new_n1226__, new_new_n1227__,
    new_new_n1228__, new_new_n1229__, new_new_n1230__, new_new_n1231__,
    new_new_n1232__, new_new_n1233__, new_new_n1234__, new_new_n1235__,
    new_new_n1236__, new_new_n1237__, new_new_n1238__, new_new_n1239__,
    new_new_n1240__, new_new_n1241__, new_new_n1242__, new_new_n1243__,
    new_new_n1244__, new_new_n1245__, new_new_n1246__, new_new_n1247__,
    new_new_n1248__, new_new_n1249__, new_new_n1250__, new_new_n1251__,
    new_new_n1252__, new_new_n1253__, new_new_n1254__, new_new_n1255__,
    new_new_n1256__, new_new_n1257__, new_new_n1258__, new_new_n1259__,
    new_new_n1260__, new_new_n1261__, new_new_n1262__, new_new_n1263__,
    new_new_n1264__, new_new_n1265__, new_new_n1266__, new_new_n1267__,
    new_new_n1268__, new_new_n1269__, new_new_n1270__, new_new_n1271__,
    new_new_n1272__, new_new_n1273__, new_new_n1274__, new_new_n1275__,
    new_new_n1276__, new_new_n1277__, new_new_n1278__, new_new_n1279__,
    new_new_n1280__, new_new_n1281__, new_new_n1282__, new_new_n1283__,
    new_new_n1284__, new_new_n1285__, new_new_n1286__, new_new_n1287__,
    new_new_n1288__, new_new_n1289__, new_new_n1290__, new_new_n1291__,
    new_new_n1292__, new_new_n1293__, new_new_n1294__, new_new_n1295__,
    new_new_n1296__, new_new_n1297__, new_new_n1298__, new_new_n1299__,
    new_new_n1300__, new_new_n1301__, new_new_n1302__, new_new_n1303__,
    new_new_n1304__, new_new_n1305__, new_new_n1306__, new_new_n1307__,
    new_new_n1308__, new_new_n1309__, new_new_n1310__, new_new_n1311__,
    new_new_n1312__, new_new_n1313__, new_new_n1314__, new_new_n1315__,
    new_new_n1316__, new_new_n1317__, new_new_n1318__, new_new_n1319__,
    new_new_n1320__, new_new_n1321__, new_new_n1322__, new_new_n1323__,
    new_new_n1324__, new_new_n1325__, new_new_n1326__, new_new_n1327__,
    new_new_n1328__, new_new_n1329__, new_new_n1330__, new_new_n1331__,
    new_new_n1332__, new_new_n1333__, new_new_n1334__, new_new_n1335__,
    new_new_n1336__, new_new_n1337__, new_new_n1338__, new_new_n1339__,
    new_new_n1340__, new_new_n1341__, new_new_n1342__, new_new_n1343__,
    new_new_n1344__, new_new_n1345__, new_new_n1346__, new_new_n1347__,
    new_new_n1348__, new_new_n1349__, new_new_n1350__, new_new_n1351__,
    new_new_n1352__, new_new_n1353__, new_new_n1354__, new_new_n1355__,
    new_new_n1356__, new_new_n1357__, new_new_n1358__, new_new_n1359__,
    new_new_n1360__, new_new_n1361__, new_new_n1362__, new_new_n1363__,
    new_new_n1364__, new_new_n1365__, new_new_n1366__, new_new_n1367__,
    new_new_n1368__, new_new_n1369__, new_new_n1370__, new_new_n1371__,
    new_new_n1372__, new_new_n1373__, new_new_n1374__, new_new_n1375__,
    new_new_n1376__, new_new_n1377__, new_new_n1378__, new_new_n1379__,
    new_new_n1380__, new_new_n1381__, new_new_n1382__, new_new_n1383__,
    new_new_n1384__, new_new_n1385__, new_new_n1386__, new_new_n1387__,
    new_new_n1388__, new_new_n1389__, new_new_n1390__, new_new_n1391__,
    new_new_n1392__, new_new_n1393__, new_new_n1394__, new_new_n1395__,
    new_new_n1396__, new_new_n1397__, new_new_n1398__, new_new_n1399__,
    new_new_n1400__, new_new_n1401__, new_new_n1402__, new_new_n1403__,
    new_new_n1404__, new_new_n1405__, new_new_n1406__, new_new_n1407__,
    new_new_n1408__, new_new_n1409__, new_new_n1410__, new_new_n1411__,
    new_new_n1412__, new_new_n1413__, new_new_n1414__, new_new_n1415__,
    new_new_n1416__, new_new_n1417__, new_new_n1418__, new_new_n1419__,
    new_new_n1420__, new_new_n1421__, new_new_n1422__, new_new_n1423__,
    new_new_n1424__, new_new_n1425__, new_new_n1426__, new_new_n1427__,
    new_new_n1428__, new_new_n1429__, new_new_n1430__, new_new_n1431__,
    new_new_n1432__, new_new_n1433__, new_new_n1434__, new_new_n1435__,
    new_new_n1436__, new_new_n1437__, new_new_n1438__, new_new_n1439__,
    new_new_n1440__, new_new_n1441__, new_new_n1442__, new_new_n1443__,
    new_new_n1444__, new_new_n1445__, new_new_n1446__, new_new_n1447__,
    new_new_n1448__, new_new_n1449__, new_new_n1450__, new_new_n1451__,
    new_new_n1452__, new_new_n1453__, new_new_n1454__, new_new_n1455__,
    new_new_n1456__, new_new_n1457__, new_new_n1458__, new_new_n1459__,
    new_new_n1460__, new_new_n1461__, new_new_n1462__, new_new_n1463__,
    new_new_n1464__, new_new_n1465__, new_new_n1466__, new_new_n1467__,
    new_new_n1468__, new_new_n1469__, new_new_n1470__, new_new_n1471__,
    new_new_n1472__, new_new_n1473__, new_new_n1474__, new_new_n1475__,
    new_new_n1476__, new_new_n1477__, new_new_n1478__, new_new_n1479__,
    new_new_n1480__, new_new_n1481__, new_new_n1482__, new_new_n1483__,
    new_new_n1484__, new_new_n1485__, new_new_n1486__, new_new_n1487__,
    new_new_n1488__, new_new_n1489__, new_new_n1490__, new_new_n1491__,
    new_new_n1492__, new_new_n1493__, new_new_n1494__, new_new_n1495__,
    new_new_n1496__, new_new_n1497__, new_new_n1498__, new_new_n1499__,
    new_new_n1500__, new_new_n1501__, new_new_n1502__, new_new_n1503__,
    new_new_n1504__, new_new_n1505__, new_new_n1506__, new_new_n1507__,
    new_new_n1508__, new_new_n1509__, new_new_n1510__, new_new_n1511__,
    new_new_n1512__, new_new_n1513__, new_new_n1514__, new_new_n1515__,
    new_new_n1516__, new_new_n1517__, new_new_n1518__, new_new_n1519__,
    new_new_n1520__, new_new_n1521__, new_new_n1522__, new_new_n1523__,
    new_new_n1524__, new_new_n1525__, new_new_n1526__, new_new_n1527__,
    new_new_n1528__, new_new_n1529__, new_new_n1530__, new_new_n1531__,
    new_new_n1532__, new_new_n1533__, new_new_n1534__, new_new_n1535__,
    new_new_n1786__, new_new_n1787__, new_new_n1788__, new_new_n1789__,
    new_new_n1790__, new_new_n1791__, new_new_n1792__, new_new_n1793__,
    new_new_n1794__, new_new_n1795__, new_new_n1796__, new_new_n1797__,
    new_new_n1798__, new_new_n1799__, new_new_n1800__, new_new_n1801__,
    new_new_n1802__, new_new_n1803__, new_new_n1804__, new_new_n1805__,
    new_new_n1806__, new_new_n1807__, new_new_n1808__, new_new_n1809__,
    new_new_n1810__, new_new_n1811__, new_new_n1812__, new_new_n1813__,
    new_new_n1814__, new_new_n1815__, new_new_n1816__, new_new_n1817__,
    new_new_n1818__, new_new_n1819__, new_new_n1820__, new_new_n1821__,
    new_new_n1822__, new_new_n1823__, new_new_n1824__, new_new_n1825__,
    new_new_n1826__, new_new_n1827__, new_new_n1828__, new_new_n1829__,
    new_new_n1830__, new_new_n1831__, new_new_n1832__, new_new_n1833__,
    new_new_n1834__, new_new_n1835__, new_new_n1836__, new_new_n1837__,
    new_new_n1838__, new_new_n1839__, new_new_n1840__, new_new_n1841__,
    new_new_n1842__, new_new_n1843__, new_new_n1844__, new_new_n1845__,
    new_new_n1846__, new_new_n1847__, new_new_n1848__, new_new_n1849__,
    new_new_n1850__, new_new_n1851__, new_new_n1852__, new_new_n1853__,
    new_new_n1854__, new_new_n1855__, new_new_n1856__, new_new_n1857__,
    new_new_n1858__, new_new_n1859__, new_new_n1860__, new_new_n1861__,
    new_new_n1862__, new_new_n1863__, new_new_n1864__, new_new_n1865__,
    new_new_n1866__, new_new_n1867__, new_new_n1868__, new_new_n1869__,
    new_new_n1870__, new_new_n1871__, new_new_n1872__, new_new_n1873__,
    new_new_n1874__, new_new_n1875__, new_new_n1876__, new_new_n1877__,
    new_new_n1878__, new_new_n1879__, new_new_n1880__, new_new_n1881__,
    new_new_n1882__, new_new_n1883__, new_new_n1884__, new_new_n1885__,
    new_new_n1886__, new_new_n1887__, new_new_n1888__, new_new_n1889__,
    new_new_n1890__, new_new_n1891__, new_new_n1892__, new_new_n1893__,
    new_new_n1894__, new_new_n1895__, new_new_n1896__, new_new_n1897__,
    new_new_n1898__, new_new_n1899__, new_new_n1900__, new_new_n1901__,
    new_new_n1902__, new_new_n1903__, new_new_n1904__, new_new_n1905__,
    new_new_n1906__, new_new_n1907__, new_new_n1908__, new_new_n1909__,
    new_new_n1910__, new_new_n1911__, new_new_n1912__, new_new_n1913__,
    new_new_n1914__, new_new_n1915__, new_new_n1916__, new_new_n1917__,
    new_new_n1918__, new_new_n1919__, new_new_n1920__, new_new_n1921__,
    new_new_n1922__, new_new_n1923__, new_new_n1924__, new_new_n1925__,
    new_new_n1926__, new_new_n1927__, new_new_n1928__, new_new_n1929__,
    new_new_n1930__, new_new_n1931__, new_new_n1932__, new_new_n1933__,
    new_new_n1934__, new_new_n1935__, new_new_n1936__, new_new_n1937__,
    new_new_n1938__, new_new_n1939__, new_new_n1940__, new_new_n1941__,
    new_new_n1942__, new_new_n1943__, new_new_n1944__, new_new_n1945__,
    new_new_n1946__, new_new_n1947__, new_new_n1948__, new_new_n1949__,
    new_new_n1950__, new_new_n1951__, new_new_n1952__, new_new_n1953__,
    new_new_n1954__, new_new_n1955__, new_new_n1956__, new_new_n1957__,
    new_new_n1958__, new_new_n1959__, new_new_n1960__, new_new_n1961__,
    new_new_n1962__, new_new_n1963__, new_new_n1964__, new_new_n1965__,
    new_new_n1966__, new_new_n1967__, new_new_n1968__, new_new_n1969__,
    new_new_n1970__, new_new_n1971__, new_new_n1972__, new_new_n1973__,
    new_new_n1974__, new_new_n1975__, new_new_n1976__, new_new_n1977__,
    new_new_n1978__, new_new_n1979__, new_new_n1980__, new_new_n1981__,
    new_new_n1982__, new_new_n1983__, new_new_n1984__, new_new_n1985__,
    new_new_n1986__, new_new_n1987__, new_new_n1988__, new_new_n1989__,
    new_new_n1990__, new_new_n1991__, new_new_n1992__, new_new_n1993__,
    new_new_n1994__, new_new_n1995__, new_new_n1996__, new_new_n1997__,
    new_new_n1998__, new_new_n1999__, new_new_n2000__, new_new_n2001__,
    new_new_n2002__, new_new_n2003__, new_new_n2004__, new_new_n2005__,
    new_new_n2006__, new_new_n2007__, new_new_n2008__, new_new_n2009__,
    new_new_n2010__, new_new_n2011__, new_new_n2012__, new_new_n2013__,
    new_new_n2014__, new_new_n2015__, new_new_n2016__, new_new_n2017__,
    new_new_n2018__, new_new_n2019__, new_new_n2020__, new_new_n2021__,
    new_new_n2022__, new_new_n2023__, new_new_n2024__, new_new_n2025__,
    new_new_n2026__, new_new_n2027__, new_new_n2028__, new_new_n2029__,
    new_new_n2030__, new_new_n2031__, new_new_n2032__, new_new_n2033__,
    new_new_n2034__, new_new_n2035__, new_new_n2036__, new_new_n2037__,
    new_new_n2038__, new_new_n2039__, new_new_n2040__, new_new_n2041__,
    new_new_n2042__, new_new_n2043__, new_new_n2044__, new_new_n2045__,
    new_new_n2046__, new_new_n2047__, new_new_n2048__, new_new_n2049__,
    new_new_n2050__, new_new_n2051__, new_new_n2052__, new_new_n2053__,
    new_new_n2054__, new_new_n2055__, new_new_n2056__, new_new_n2057__,
    new_new_n2058__, new_new_n2059__, new_new_n2060__, new_new_n2061__,
    new_new_n2062__, new_new_n2063__, new_new_n2064__, new_new_n2065__,
    new_new_n2066__, new_new_n2067__, new_new_n2068__, new_new_n2069__,
    new_new_n2070__, new_new_n2071__, new_new_n2072__, new_new_n2073__,
    new_new_n2074__, new_new_n2075__, new_new_n2076__, new_new_n2077__,
    new_new_n2078__, new_new_n2079__, new_new_n2080__, new_new_n2081__,
    new_new_n2082__, new_new_n2083__, new_new_n2084__, new_new_n2085__,
    new_new_n2086__, new_new_n2087__, new_new_n2088__, new_new_n2089__,
    new_new_n2090__, new_new_n2091__, new_new_n2092__, new_new_n2093__,
    new_new_n2094__, new_new_n2095__, new_new_n2096__, new_new_n2097__,
    new_new_n2098__, new_new_n2099__, new_new_n2100__, new_new_n2101__,
    new_new_n2102__, new_new_n2103__, new_new_n2104__, new_new_n2105__,
    new_new_n2106__, new_new_n2107__, new_new_n2108__, new_new_n2109__,
    new_new_n2110__, new_new_n2111__, new_new_n2112__, new_new_n2113__,
    new_new_n2114__, new_new_n2115__, new_new_n2116__, new_new_n2117__,
    new_new_n2118__, new_new_n2119__, new_new_n2120__, new_new_n2121__,
    new_new_n2122__, new_new_n2123__, new_new_n2124__, new_new_n2125__,
    new_new_n2126__, new_new_n2127__, new_new_n2128__, new_new_n2129__,
    new_new_n2130__, new_new_n2131__, new_new_n2132__, new_new_n2133__,
    new_new_n2134__, new_new_n2135__, new_new_n2136__, new_new_n2137__,
    new_new_n2138__, new_new_n2139__, n3365, n3368, n3371, n3374, n3377,
    n3380, n3383, n3386, n3389, n3392, n3395, n3398, n3401, n3404, n3407,
    n3410, n3413, n3416, n3419, n3422, n3425, n3428, n3431, n3434, n3437,
    n3440, n3443, n3446, n3449, n3452, n3455, n3458, n3461, n3464, n3467,
    n3470, n3473, n3476, n3479, n3482, n3485, n3488, n3491, n3494, n3497,
    n3500, n3503, n3506, n3509, n3512, n3515, n3518, n3521, n3524, n3527,
    n3530, n3533, n3536, n3539, n3542, n3545, n3548, n3551, n3554, n3557,
    n3560, n3563, n3566, n3569, n3572, n3575, n3578, n3581, n3584, n3587,
    n3590, n3593, n3596, n3599, n3602, n3605, n3608, n3611, n3614, n3617,
    n3620, n3623, n3626, n3629, n3632, n3635, n3638, n3641, n3644, n3647,
    n3650, n3653, n3656, n3659, n3662, n3665, n3668, n3671, n3674, n3677,
    n3680, n3683, n3686, n3689, n3692, n3695, n3698, n3701, n3704, n3707,
    n3710, n3713, n3716, n3719, n3722, n3725, n3728, n3731, n3734, n3737,
    n3740, n3743, n3746, n3749, n3752, n3755, n3758, n3761, n3764, n3767,
    n3770, n3773, n3776, n3779, n3782, n3785, n3788, n3791, n3794, n3797,
    n3800, n3803, n3806, n3809, n3812, n3815, n3818, n3821, n3824, n3827,
    n3830, n3833, n3836, n3839, n3842, n3845, n3848, n3851, n3854, n3857,
    n3860, n3863, n3866, n3869, n3872, n3875, n3878, n3881, n3884, n3887,
    n3890, n3893, n3896, n3899, n3902, n3905, n3908, n3911, n3914, n3917,
    n3920, n3923, n3926, n3929, n3932, n3935, n3938, n3941, n3944, n3947,
    n3950, n3953, n3956, n3959, n3962, n3965, n3968, n3971, n3974, n3977,
    n3980, n3983, n3986, n3989, n3992, n3995, n3998, n4001, n4004, n4007,
    n4010, n4013, n4016;
  buf1  g0000(.din(G1), .dout(new_new_n510__));
  buf1  g0001(.din(G2), .dout(new_new_n512__));
  buf1  g0002(.din(G3), .dout(new_new_n514__));
  buf1  g0003(.din(G4), .dout(new_new_n516__));
  buf1  g0004(.din(G5), .dout(new_new_n518__));
  buf1  g0005(.din(G6), .dout(new_new_n520__));
  buf1  g0006(.din(G7), .dout(new_new_n522__));
  buf1  g0007(.din(G8), .dout(new_new_n524__));
  buf1  g0008(.din(G9), .dout(new_new_n526__));
  buf1  g0009(.din(G10), .dout(new_new_n528__));
  buf1  g0010(.din(G11), .dout(new_new_n530__));
  buf1  g0011(.din(G12), .dout(new_new_n532__));
  buf1  g0012(.din(G13), .dout(new_new_n534__));
  buf1  g0013(.din(G14), .dout(new_new_n536__));
  buf1  g0014(.din(G15), .dout(new_new_n538__));
  buf1  g0015(.din(G16), .dout(new_new_n540__));
  buf1  g0016(.din(G17), .dout(new_new_n542__));
  buf1  g0017(.din(G18), .dout(new_new_n544__));
  buf1  g0018(.din(G19), .dout(new_new_n546__));
  buf1  g0019(.din(G20), .dout(new_new_n548__));
  buf1  g0020(.din(G21), .dout(new_new_n550__));
  buf1  g0021(.din(G22), .dout(new_new_n552__));
  buf1  g0022(.din(G23), .dout(new_new_n554__));
  buf1  g0023(.din(G24), .dout(new_new_n556__));
  buf1  g0024(.din(G25), .dout(new_new_n558__));
  buf1  g0025(.din(G26), .dout(new_new_n560__));
  buf1  g0026(.din(G27), .dout(new_new_n562__));
  buf1  g0027(.din(G28), .dout(new_new_n564__));
  buf1  g0028(.din(G29), .dout(new_new_n566__));
  buf1  g0029(.din(G30), .dout(new_new_n568__));
  buf1  g0030(.din(G31), .dout(new_new_n570__));
  buf1  g0031(.din(G32), .dout(new_new_n572__));
  buf1  g0032(.din(G33), .dout(new_new_n574__));
  buf1  g0033(.din(G34), .dout(new_new_n576__));
  buf1  g0034(.din(G35), .dout(new_new_n578__));
  buf1  g0035(.din(G36), .dout(new_new_n580__));
  buf1  g0036(.din(G37), .dout(new_new_n582__));
  buf1  g0037(.din(G38), .dout(new_new_n584__));
  buf1  g0038(.din(G39), .dout(new_new_n586__));
  buf1  g0039(.din(G40), .dout(new_new_n588__));
  buf1  g0040(.din(G41), .dout(new_new_n590__));
  buf1  g0041(.din(n621_lo), .dout(new_new_n592__));
  not1  g0042(.din(n621_lo), .dout(new_new_n593__));
  buf1  g0043(.din(n630_lo), .dout(new_new_n594__));
  not1  g0044(.din(n630_lo), .dout(new_new_n595__));
  buf1  g0045(.din(n633_lo), .dout(new_new_n596__));
  not1  g0046(.din(n633_lo), .dout(new_new_n597__));
  buf1  g0047(.din(n642_lo), .dout(new_new_n598__));
  not1  g0048(.din(n642_lo), .dout(new_new_n599__));
  buf1  g0049(.din(n645_lo), .dout(new_new_n600__));
  not1  g0050(.din(n645_lo), .dout(new_new_n601__));
  buf1  g0051(.din(n654_lo), .dout(new_new_n602__));
  not1  g0052(.din(n654_lo), .dout(new_new_n603__));
  buf1  g0053(.din(n657_lo), .dout(new_new_n604__));
  not1  g0054(.din(n657_lo), .dout(new_new_n605__));
  buf1  g0055(.din(n666_lo), .dout(new_new_n606__));
  not1  g0056(.din(n666_lo), .dout(new_new_n607__));
  buf1  g0057(.din(n669_lo), .dout(new_new_n608__));
  not1  g0058(.din(n669_lo), .dout(new_new_n609__));
  buf1  g0059(.din(n678_lo), .dout(new_new_n610__));
  not1  g0060(.din(n678_lo), .dout(new_new_n611__));
  buf1  g0061(.din(n681_lo), .dout(new_new_n612__));
  not1  g0062(.din(n681_lo), .dout(new_new_n613__));
  buf1  g0063(.din(n690_lo), .dout(new_new_n614__));
  not1  g0064(.din(n690_lo), .dout(new_new_n615__));
  buf1  g0065(.din(n693_lo), .dout(new_new_n616__));
  not1  g0066(.din(n693_lo), .dout(new_new_n617__));
  buf1  g0067(.din(n702_lo), .dout(new_new_n618__));
  not1  g0068(.din(n702_lo), .dout(new_new_n619__));
  buf1  g0069(.din(n705_lo), .dout(new_new_n620__));
  not1  g0070(.din(n705_lo), .dout(new_new_n621__));
  buf1  g0071(.din(n714_lo), .dout(new_new_n622__));
  not1  g0072(.din(n714_lo), .dout(new_new_n623__));
  buf1  g0073(.din(n717_lo), .dout(new_new_n624__));
  not1  g0074(.din(n717_lo), .dout(new_new_n625__));
  buf1  g0075(.din(n726_lo), .dout(new_new_n626__));
  not1  g0076(.din(n726_lo), .dout(new_new_n627__));
  buf1  g0077(.din(n729_lo), .dout(new_new_n628__));
  not1  g0078(.din(n729_lo), .dout(new_new_n629__));
  buf1  g0079(.din(n738_lo), .dout(new_new_n630__));
  not1  g0080(.din(n738_lo), .dout(new_new_n631__));
  buf1  g0081(.din(n741_lo), .dout(new_new_n632__));
  not1  g0082(.din(n741_lo), .dout(new_new_n633__));
  buf1  g0083(.din(n750_lo), .dout(new_new_n634__));
  not1  g0084(.din(n750_lo), .dout(new_new_n635__));
  buf1  g0085(.din(n753_lo), .dout(new_new_n636__));
  not1  g0086(.din(n753_lo), .dout(new_new_n637__));
  buf1  g0087(.din(n762_lo), .dout(new_new_n638__));
  not1  g0088(.din(n762_lo), .dout(new_new_n639__));
  buf1  g0089(.din(n765_lo), .dout(new_new_n640__));
  not1  g0090(.din(n765_lo), .dout(new_new_n641__));
  buf1  g0091(.din(n774_lo), .dout(new_new_n642__));
  not1  g0092(.din(n774_lo), .dout(new_new_n643__));
  buf1  g0093(.din(n777_lo), .dout(new_new_n644__));
  not1  g0094(.din(n777_lo), .dout(new_new_n645__));
  buf1  g0095(.din(n786_lo), .dout(new_new_n646__));
  not1  g0096(.din(n786_lo), .dout(new_new_n647__));
  buf1  g0097(.din(n789_lo), .dout(new_new_n648__));
  not1  g0098(.din(n789_lo), .dout(new_new_n649__));
  buf1  g0099(.din(n798_lo), .dout(new_new_n650__));
  not1  g0100(.din(n798_lo), .dout(new_new_n651__));
  buf1  g0101(.din(n801_lo), .dout(new_new_n652__));
  not1  g0102(.din(n801_lo), .dout(new_new_n653__));
  buf1  g0103(.din(n810_lo), .dout(new_new_n654__));
  not1  g0104(.din(n810_lo), .dout(new_new_n655__));
  buf1  g0105(.din(n813_lo), .dout(new_new_n656__));
  not1  g0106(.din(n813_lo), .dout(new_new_n657__));
  buf1  g0107(.din(n822_lo), .dout(new_new_n658__));
  not1  g0108(.din(n822_lo), .dout(new_new_n659__));
  buf1  g0109(.din(n825_lo), .dout(new_new_n660__));
  not1  g0110(.din(n825_lo), .dout(new_new_n661__));
  buf1  g0111(.din(n834_lo), .dout(new_new_n662__));
  not1  g0112(.din(n834_lo), .dout(new_new_n663__));
  buf1  g0113(.din(n837_lo), .dout(new_new_n664__));
  not1  g0114(.din(n837_lo), .dout(new_new_n665__));
  buf1  g0115(.din(n846_lo), .dout(new_new_n666__));
  not1  g0116(.din(n846_lo), .dout(new_new_n667__));
  buf1  g0117(.din(n849_lo), .dout(new_new_n668__));
  not1  g0118(.din(n849_lo), .dout(new_new_n669__));
  buf1  g0119(.din(n858_lo), .dout(new_new_n670__));
  not1  g0120(.din(n858_lo), .dout(new_new_n671__));
  buf1  g0121(.din(n861_lo), .dout(new_new_n672__));
  not1  g0122(.din(n861_lo), .dout(new_new_n673__));
  buf1  g0123(.din(n870_lo), .dout(new_new_n674__));
  not1  g0124(.din(n870_lo), .dout(new_new_n675__));
  buf1  g0125(.din(n873_lo), .dout(new_new_n676__));
  not1  g0126(.din(n873_lo), .dout(new_new_n677__));
  buf1  g0127(.din(n882_lo), .dout(new_new_n678__));
  not1  g0128(.din(n882_lo), .dout(new_new_n679__));
  buf1  g0129(.din(n885_lo), .dout(new_new_n680__));
  not1  g0130(.din(n885_lo), .dout(new_new_n681__));
  buf1  g0131(.din(n894_lo), .dout(new_new_n682__));
  not1  g0132(.din(n894_lo), .dout(new_new_n683__));
  buf1  g0133(.din(n897_lo), .dout(new_new_n684__));
  not1  g0134(.din(n897_lo), .dout(new_new_n685__));
  buf1  g0135(.din(n906_lo), .dout(new_new_n686__));
  not1  g0136(.din(n906_lo), .dout(new_new_n687__));
  buf1  g0137(.din(n909_lo), .dout(new_new_n688__));
  not1  g0138(.din(n909_lo), .dout(new_new_n689__));
  buf1  g0139(.din(n918_lo), .dout(new_new_n690__));
  not1  g0140(.din(n918_lo), .dout(new_new_n691__));
  buf1  g0141(.din(n921_lo), .dout(new_new_n692__));
  not1  g0142(.din(n921_lo), .dout(new_new_n693__));
  buf1  g0143(.din(n930_lo), .dout(new_new_n694__));
  not1  g0144(.din(n930_lo), .dout(new_new_n695__));
  buf1  g0145(.din(n933_lo), .dout(new_new_n696__));
  not1  g0146(.din(n933_lo), .dout(new_new_n697__));
  buf1  g0147(.din(n942_lo), .dout(new_new_n698__));
  not1  g0148(.din(n942_lo), .dout(new_new_n699__));
  buf1  g0149(.din(n945_lo), .dout(new_new_n700__));
  not1  g0150(.din(n945_lo), .dout(new_new_n701__));
  buf1  g0151(.din(n954_lo), .dout(new_new_n702__));
  not1  g0152(.din(n954_lo), .dout(new_new_n703__));
  buf1  g0153(.din(n957_lo), .dout(new_new_n704__));
  not1  g0154(.din(n957_lo), .dout(new_new_n705__));
  buf1  g0155(.din(n966_lo), .dout(new_new_n706__));
  not1  g0156(.din(n966_lo), .dout(new_new_n707__));
  buf1  g0157(.din(n969_lo), .dout(new_new_n708__));
  not1  g0158(.din(n969_lo), .dout(new_new_n709__));
  buf1  g0159(.din(n978_lo), .dout(new_new_n710__));
  not1  g0160(.din(n978_lo), .dout(new_new_n711__));
  buf1  g0161(.din(n981_lo), .dout(new_new_n712__));
  not1  g0162(.din(n981_lo), .dout(new_new_n713__));
  buf1  g0163(.din(n990_lo), .dout(new_new_n714__));
  not1  g0164(.din(n990_lo), .dout(new_new_n715__));
  buf1  g0165(.din(n993_lo), .dout(new_new_n716__));
  not1  g0166(.din(n993_lo), .dout(new_new_n717__));
  buf1  g0167(.din(n1002_lo), .dout(new_new_n718__));
  not1  g0168(.din(n1002_lo), .dout(new_new_n719__));
  buf1  g0169(.din(n1005_lo), .dout(new_new_n720__));
  buf1  g0170(.din(n1017_lo), .dout(new_new_n722__));
  buf1  g0171(.din(n1029_lo), .dout(new_new_n724__));
  buf1  g0172(.din(n1041_lo), .dout(new_new_n726__));
  buf1  g0173(.din(n1053_lo), .dout(new_new_n728__));
  buf1  g0174(.din(n1065_lo), .dout(new_new_n730__));
  buf1  g0175(.din(n1077_lo), .dout(new_new_n732__));
  buf1  g0176(.din(n1089_lo), .dout(new_new_n734__));
  buf1  g0177(.din(n1101_lo), .dout(new_new_n736__));
  buf1  g0178(.din(n602_o2), .dout(new_new_n738__));
  not1  g0179(.din(n602_o2), .dout(new_new_n739__));
  buf1  g0180(.din(n639_o2), .dout(new_new_n740__));
  not1  g0181(.din(n639_o2), .dout(new_new_n741__));
  buf1  g0182(.din(n678_o2), .dout(new_new_n742__));
  not1  g0183(.din(n678_o2), .dout(new_new_n743__));
  buf1  g0184(.din(n658_o2), .dout(new_new_n744__));
  not1  g0185(.din(n658_o2), .dout(new_new_n745__));
  buf1  g0186(.din(n783_o2), .dout(new_new_n746__));
  not1  g0187(.din(n783_o2), .dout(new_new_n747__));
  buf1  g0188(.din(n802_o2), .dout(new_new_n748__));
  not1  g0189(.din(n802_o2), .dout(new_new_n749__));
  buf1  g0190(.din(n726_o2), .dout(new_new_n750__));
  not1  g0191(.din(n726_o2), .dout(new_new_n751__));
  buf1  g0192(.din(n763_o2), .dout(new_new_n752__));
  not1  g0193(.din(n763_o2), .dout(new_new_n753__));
  buf1  g0194(.din(n1644_o2), .dout(new_new_n754__));
  buf1  g0195(.din(n1645_o2), .dout(new_new_n756__));
  buf1  g0196(.din(n1646_o2), .dout(new_new_n758__));
  buf1  g0197(.din(n1647_o2), .dout(new_new_n760__));
  buf1  g0198(.din(n1648_o2), .dout(new_new_n762__));
  buf1  g0199(.din(n1649_o2), .dout(new_new_n764__));
  buf1  g0200(.din(n1650_o2), .dout(new_new_n766__));
  buf1  g0201(.din(n1651_o2), .dout(new_new_n768__));
  buf1  g0202(.din(n1652_o2), .dout(new_new_n770__));
  buf1  g0203(.din(n1653_o2), .dout(new_new_n772__));
  buf1  g0204(.din(n1654_o2), .dout(new_new_n774__));
  buf1  g0205(.din(n1655_o2), .dout(new_new_n776__));
  buf1  g0206(.din(n1656_o2), .dout(new_new_n778__));
  buf1  g0207(.din(n1657_o2), .dout(new_new_n780__));
  buf1  g0208(.din(n1658_o2), .dout(new_new_n782__));
  buf1  g0209(.din(n1659_o2), .dout(new_new_n784__));
  buf1  g0210(.din(n1660_o2), .dout(new_new_n786__));
  buf1  g0211(.din(n1661_o2), .dout(new_new_n788__));
  buf1  g0212(.din(n1662_o2), .dout(new_new_n790__));
  buf1  g0213(.din(n1663_o2), .dout(new_new_n792__));
  buf1  g0214(.din(n1664_o2), .dout(new_new_n794__));
  buf1  g0215(.din(n1665_o2), .dout(new_new_n796__));
  buf1  g0216(.din(n1666_o2), .dout(new_new_n798__));
  buf1  g0217(.din(n1667_o2), .dout(new_new_n800__));
  buf1  g0218(.din(n1668_o2), .dout(new_new_n802__));
  buf1  g0219(.din(n1669_o2), .dout(new_new_n804__));
  buf1  g0220(.din(n1670_o2), .dout(new_new_n806__));
  buf1  g0221(.din(n1671_o2), .dout(new_new_n808__));
  buf1  g0222(.din(n1672_o2), .dout(new_new_n810__));
  buf1  g0223(.din(n1673_o2), .dout(new_new_n812__));
  buf1  g0224(.din(n1674_o2), .dout(new_new_n814__));
  buf1  g0225(.din(n1675_o2), .dout(new_new_n816__));
  buf1  g0226(.din(n685_o2), .dout(new_new_n818__));
  not1  g0227(.din(n685_o2), .dout(new_new_n819__));
  buf1  g0228(.din(n680_o2), .dout(new_new_n820__));
  not1  g0229(.din(n680_o2), .dout(new_new_n821__));
  buf1  g0230(.din(n822_o2), .dout(new_new_n822__));
  not1  g0231(.din(n822_o2), .dout(new_new_n823__));
  buf1  g0232(.din(n843_o2), .dout(new_new_n824__));
  not1  g0233(.din(n843_o2), .dout(new_new_n825__));
  buf1  g0234(.din(n842_o2), .dout(new_new_n826__));
  not1  g0235(.din(n842_o2), .dout(new_new_n827__));
  buf1  g0236(.din(n681_o2), .dout(new_new_n828__));
  not1  g0237(.din(n681_o2), .dout(new_new_n829__));
  buf1  g0238(.din(n684_o2), .dout(new_new_n830__));
  not1  g0239(.din(n684_o2), .dout(new_new_n831__));
  buf1  g0240(.din(n686_o2), .dout(new_new_n832__));
  not1  g0241(.din(n686_o2), .dout(new_new_n833__));
  buf1  g0242(.din(n823_o2), .dout(new_new_n834__));
  not1  g0243(.din(n823_o2), .dout(new_new_n835__));
  buf1  g0244(.din(n683_o2), .dout(new_new_n836__));
  not1  g0245(.din(n683_o2), .dout(new_new_n837__));
  buf1  g0246(.din(n688_o2), .dout(new_new_n838__));
  not1  g0247(.din(n688_o2), .dout(new_new_n839__));
  buf1  g0248(.din(n803_o2), .dout(new_new_n840__));
  not1  g0249(.din(n803_o2), .dout(new_new_n841__));
  buf1  g0250(.din(n862_o2), .dout(new_new_n842__));
  not1  g0251(.din(n862_o2), .dout(new_new_n843__));
  buf1  g0252(.din(n764_o2), .dout(new_new_n844__));
  not1  g0253(.din(n764_o2), .dout(new_new_n845__));
  buf1  g0254(.din(n863_o2), .dout(new_new_n846__));
  not1  g0255(.din(n863_o2), .dout(new_new_n847__));
  buf1  g0256(.din(n886_o2), .dout(new_new_n848__));
  not1  g0257(.din(n886_o2), .dout(new_new_n849__));
  buf1  g0258(.din(lo002_buf_o2), .dout(new_new_n850__));
  buf1  g0259(.din(lo006_buf_o2), .dout(new_new_n852__));
  buf1  g0260(.din(lo010_buf_o2), .dout(new_new_n854__));
  buf1  g0261(.din(lo014_buf_o2), .dout(new_new_n856__));
  buf1  g0262(.din(lo018_buf_o2), .dout(new_new_n858__));
  buf1  g0263(.din(lo022_buf_o2), .dout(new_new_n860__));
  buf1  g0264(.din(lo026_buf_o2), .dout(new_new_n862__));
  buf1  g0265(.din(lo030_buf_o2), .dout(new_new_n864__));
  buf1  g0266(.din(lo034_buf_o2), .dout(new_new_n866__));
  buf1  g0267(.din(lo038_buf_o2), .dout(new_new_n868__));
  buf1  g0268(.din(lo042_buf_o2), .dout(new_new_n870__));
  buf1  g0269(.din(lo046_buf_o2), .dout(new_new_n872__));
  buf1  g0270(.din(lo050_buf_o2), .dout(new_new_n874__));
  buf1  g0271(.din(lo054_buf_o2), .dout(new_new_n876__));
  buf1  g0272(.din(lo058_buf_o2), .dout(new_new_n878__));
  buf1  g0273(.din(lo062_buf_o2), .dout(new_new_n880__));
  buf1  g0274(.din(lo066_buf_o2), .dout(new_new_n882__));
  buf1  g0275(.din(lo070_buf_o2), .dout(new_new_n884__));
  buf1  g0276(.din(lo074_buf_o2), .dout(new_new_n886__));
  buf1  g0277(.din(lo078_buf_o2), .dout(new_new_n888__));
  buf1  g0278(.din(lo082_buf_o2), .dout(new_new_n890__));
  buf1  g0279(.din(lo086_buf_o2), .dout(new_new_n892__));
  buf1  g0280(.din(lo090_buf_o2), .dout(new_new_n894__));
  buf1  g0281(.din(lo094_buf_o2), .dout(new_new_n896__));
  buf1  g0282(.din(lo098_buf_o2), .dout(new_new_n898__));
  buf1  g0283(.din(lo102_buf_o2), .dout(new_new_n900__));
  buf1  g0284(.din(lo106_buf_o2), .dout(new_new_n902__));
  buf1  g0285(.din(lo110_buf_o2), .dout(new_new_n904__));
  buf1  g0286(.din(lo114_buf_o2), .dout(new_new_n906__));
  buf1  g0287(.din(lo118_buf_o2), .dout(new_new_n908__));
  buf1  g0288(.din(lo122_buf_o2), .dout(new_new_n910__));
  buf1  g0289(.din(lo126_buf_o2), .dout(new_new_n912__));
  buf1  g0290(.din(n600_o2), .dout(new_new_n914__));
  not1  g0291(.din(n600_o2), .dout(new_new_n915__));
  buf1  g0292(.din(n601_o2), .dout(new_new_n916__));
  not1  g0293(.din(n601_o2), .dout(new_new_n917__));
  buf1  g0294(.din(n637_o2), .dout(new_new_n918__));
  not1  g0295(.din(n637_o2), .dout(new_new_n919__));
  buf1  g0296(.din(n638_o2), .dout(new_new_n920__));
  not1  g0297(.din(n638_o2), .dout(new_new_n921__));
  buf1  g0298(.din(n676_o2), .dout(new_new_n922__));
  not1  g0299(.din(n676_o2), .dout(new_new_n923__));
  buf1  g0300(.din(n677_o2), .dout(new_new_n924__));
  not1  g0301(.din(n677_o2), .dout(new_new_n925__));
  buf1  g0302(.din(n656_o2), .dout(new_new_n926__));
  not1  g0303(.din(n656_o2), .dout(new_new_n927__));
  buf1  g0304(.din(n657_o2), .dout(new_new_n928__));
  not1  g0305(.din(n657_o2), .dout(new_new_n929__));
  buf1  g0306(.din(n781_o2), .dout(new_new_n930__));
  not1  g0307(.din(n781_o2), .dout(new_new_n931__));
  buf1  g0308(.din(n782_o2), .dout(new_new_n932__));
  not1  g0309(.din(n782_o2), .dout(new_new_n933__));
  buf1  g0310(.din(n800_o2), .dout(new_new_n934__));
  not1  g0311(.din(n800_o2), .dout(new_new_n935__));
  buf1  g0312(.din(n801_o2), .dout(new_new_n936__));
  not1  g0313(.din(n801_o2), .dout(new_new_n937__));
  buf1  g0314(.din(n724_o2), .dout(new_new_n938__));
  not1  g0315(.din(n724_o2), .dout(new_new_n939__));
  buf1  g0316(.din(n725_o2), .dout(new_new_n940__));
  not1  g0317(.din(n725_o2), .dout(new_new_n941__));
  buf1  g0318(.din(n761_o2), .dout(new_new_n942__));
  not1  g0319(.din(n761_o2), .dout(new_new_n943__));
  buf1  g0320(.din(n762_o2), .dout(new_new_n944__));
  not1  g0321(.din(n762_o2), .dout(new_new_n945__));
  buf1  g0322(.din(lo129_buf_o2), .dout(new_new_n946__));
  not1  g0323(.din(lo129_buf_o2), .dout(new_new_n947__));
  buf1  g0324(.din(lo133_buf_o2), .dout(new_new_n948__));
  not1  g0325(.din(lo133_buf_o2), .dout(new_new_n949__));
  buf1  g0326(.din(lo137_buf_o2), .dout(new_new_n950__));
  not1  g0327(.din(lo137_buf_o2), .dout(new_new_n951__));
  buf1  g0328(.din(lo141_buf_o2), .dout(new_new_n952__));
  not1  g0329(.din(lo141_buf_o2), .dout(new_new_n953__));
  buf1  g0330(.din(lo145_buf_o2), .dout(new_new_n954__));
  not1  g0331(.din(lo145_buf_o2), .dout(new_new_n955__));
  buf1  g0332(.din(lo149_buf_o2), .dout(new_new_n956__));
  not1  g0333(.din(lo149_buf_o2), .dout(new_new_n957__));
  buf1  g0334(.din(lo153_buf_o2), .dout(new_new_n958__));
  not1  g0335(.din(lo153_buf_o2), .dout(new_new_n959__));
  buf1  g0336(.din(lo157_buf_o2), .dout(new_new_n960__));
  not1  g0337(.din(lo157_buf_o2), .dout(new_new_n961__));
  buf1  g0338(.din(lo161_buf_o2), .dout(new_new_n962__));
  not1  g0339(.din(lo161_buf_o2), .dout(new_new_n963__));
  buf1  g0340(.din(n571_o2), .dout(new_new_n964__));
  not1  g0341(.din(n571_o2), .dout(new_new_n965__));
  buf1  g0342(.din(n708_o2), .dout(new_new_n966__));
  not1  g0343(.din(n708_o2), .dout(new_new_n967__));
  buf1  g0344(.din(n608_o2), .dout(new_new_n968__));
  not1  g0345(.din(n608_o2), .dout(new_new_n969__));
  buf1  g0346(.din(n665_o2), .dout(new_new_n970__));
  not1  g0347(.din(n665_o2), .dout(new_new_n971__));
  buf1  g0348(.din(n705_o2), .dout(new_new_n972__));
  not1  g0349(.din(n705_o2), .dout(new_new_n973__));
  buf1  g0350(.din(n645_o2), .dout(new_new_n974__));
  not1  g0351(.din(n645_o2), .dout(new_new_n975__));
  buf1  g0352(.din(n745_o2), .dout(new_new_n976__));
  not1  g0353(.din(n745_o2), .dout(new_new_n977__));
  buf1  g0354(.din(n742_o2), .dout(new_new_n978__));
  not1  g0355(.din(n742_o2), .dout(new_new_n979__));
  buf1  g0356(.din(n568_o2), .dout(new_new_n980__));
  not1  g0357(.din(n568_o2), .dout(new_new_n981__));
  buf1  g0358(.din(n717_o2), .dout(new_new_n982__));
  not1  g0359(.din(n717_o2), .dout(new_new_n983__));
  buf1  g0360(.din(n605_o2), .dout(new_new_n984__));
  not1  g0361(.din(n605_o2), .dout(new_new_n985__));
  buf1  g0362(.din(n662_o2), .dout(new_new_n986__));
  not1  g0363(.din(n662_o2), .dout(new_new_n987__));
  buf1  g0364(.din(n714_o2), .dout(new_new_n988__));
  not1  g0365(.din(n714_o2), .dout(new_new_n989__));
  buf1  g0366(.din(n642_o2), .dout(new_new_n990__));
  not1  g0367(.din(n642_o2), .dout(new_new_n991__));
  buf1  g0368(.din(n754_o2), .dout(new_new_n992__));
  not1  g0369(.din(n754_o2), .dout(new_new_n993__));
  buf1  g0370(.din(n751_o2), .dout(new_new_n994__));
  not1  g0371(.din(n751_o2), .dout(new_new_n995__));
  buf1  g0372(.din(n584_o2), .dout(new_new_n996__));
  not1  g0373(.din(n584_o2), .dout(new_new_n997__));
  buf1  g0374(.din(n770_o2), .dout(new_new_n998__));
  not1  g0375(.din(n770_o2), .dout(new_new_n999__));
  buf1  g0376(.din(n789_o2), .dout(new_new_n1000__));
  not1  g0377(.din(n789_o2), .dout(new_new_n1001__));
  buf1  g0378(.din(n581_o2), .dout(new_new_n1002__));
  not1  g0379(.din(n581_o2), .dout(new_new_n1003__));
  buf1  g0380(.din(n695_o2), .dout(new_new_n1004__));
  not1  g0381(.din(n695_o2), .dout(new_new_n1005__));
  buf1  g0382(.din(n732_o2), .dout(new_new_n1006__));
  not1  g0383(.din(n732_o2), .dout(new_new_n1007__));
  buf1  g0384(.din(n593_o2), .dout(new_new_n1008__));
  not1  g0385(.din(n593_o2), .dout(new_new_n1009__));
  buf1  g0386(.din(n590_o2), .dout(new_new_n1010__));
  not1  g0387(.din(n590_o2), .dout(new_new_n1011__));
  buf1  g0388(.din(n630_o2), .dout(new_new_n1012__));
  not1  g0389(.din(n630_o2), .dout(new_new_n1013__));
  buf1  g0390(.din(n767_o2), .dout(new_new_n1014__));
  not1  g0391(.din(n767_o2), .dout(new_new_n1015__));
  buf1  g0392(.din(n786_o2), .dout(new_new_n1016__));
  not1  g0393(.din(n786_o2), .dout(new_new_n1017__));
  buf1  g0394(.din(n627_o2), .dout(new_new_n1018__));
  not1  g0395(.din(n627_o2), .dout(new_new_n1019__));
  buf1  g0396(.din(n692_o2), .dout(new_new_n1020__));
  not1  g0397(.din(n692_o2), .dout(new_new_n1021__));
  buf1  g0398(.din(n729_o2), .dout(new_new_n1022__));
  not1  g0399(.din(n729_o2), .dout(new_new_n1023__));
  buf1  g0400(.din(n621_o2), .dout(new_new_n1024__));
  not1  g0401(.din(n621_o2), .dout(new_new_n1025__));
  buf1  g0402(.din(n618_o2), .dout(new_new_n1026__));
  not1  g0403(.din(n618_o2), .dout(new_new_n1027__));
  and1  g0404(.dina(new_new_n839__), .dinb(new_new_n837__), .dout(new_new_n1028__));
  or1   g0405(.dina(new_new_n838__), .dinb(new_new_n836__), .dout(new_new_n1029__));
  and1  g0406(.dina(new_new_n844__), .dinb(new_new_n840__), .dout(new_new_n1030__));
  or1   g0407(.dina(new_new_n845__), .dinb(new_new_n841__), .dout(new_new_n1031__));
  and1  g0408(.dina(new_new_n1030__), .dinb(new_new_n1787__), .dout(new_new_n1032__));
  or1   g0409(.dina(new_new_n1031__), .dinb(new_new_n1790__), .dout(new_new_n1033__));
  and1  g0410(.dina(new_new_n1793__), .dinb(new_new_n1796__), .dout(new_new_n1034__));
  or1   g0411(.dina(new_new_n1799__), .dinb(new_new_n1802__), .dout(new_new_n1035__));
  or1   g0412(.dina(new_new_n1034__), .dinb(new_new_n595__), .dout(new_new_n1036__));
  or1   g0413(.dina(new_new_n1035__), .dinb(new_new_n594__), .dout(new_new_n1037__));
  and1  g0414(.dina(new_new_n1037__), .dinb(new_new_n1036__), .dout(new_new_n1038__));
  and1  g0415(.dina(new_new_n1793__), .dinb(new_new_n1806__), .dout(new_new_n1039__));
  or1   g0416(.dina(new_new_n1799__), .dinb(new_new_n1810__), .dout(new_new_n1040__));
  or1   g0417(.dina(new_new_n1039__), .dinb(new_new_n599__), .dout(new_new_n1041__));
  or1   g0418(.dina(new_new_n1040__), .dinb(new_new_n598__), .dout(new_new_n1042__));
  and1  g0419(.dina(new_new_n1042__), .dinb(new_new_n1041__), .dout(new_new_n1043__));
  and1  g0420(.dina(new_new_n1794__), .dinb(new_new_n1814__), .dout(new_new_n1044__));
  or1   g0421(.dina(new_new_n1800__), .dinb(new_new_n1819__), .dout(new_new_n1045__));
  or1   g0422(.dina(new_new_n1044__), .dinb(new_new_n603__), .dout(new_new_n1046__));
  or1   g0423(.dina(new_new_n1045__), .dinb(new_new_n602__), .dout(new_new_n1047__));
  and1  g0424(.dina(new_new_n1047__), .dinb(new_new_n1046__), .dout(new_new_n1048__));
  and1  g0425(.dina(new_new_n1794__), .dinb(new_new_n1823__), .dout(new_new_n1049__));
  or1   g0426(.dina(new_new_n1800__), .dinb(new_new_n1826__), .dout(new_new_n1050__));
  or1   g0427(.dina(new_new_n1049__), .dinb(new_new_n607__), .dout(new_new_n1051__));
  or1   g0428(.dina(new_new_n1050__), .dinb(new_new_n606__), .dout(new_new_n1052__));
  and1  g0429(.dina(new_new_n1052__), .dinb(new_new_n1051__), .dout(new_new_n1053__));
  and1  g0430(.dina(new_new_n835__), .dinb(new_new_n822__), .dout(new_new_n1054__));
  or1   g0431(.dina(new_new_n834__), .dinb(new_new_n823__), .dout(new_new_n1055__));
  and1  g0432(.dina(new_new_n1054__), .dinb(new_new_n1787__), .dout(new_new_n1056__));
  or1   g0433(.dina(new_new_n1055__), .dinb(new_new_n1790__), .dout(new_new_n1057__));
  and1  g0434(.dina(new_new_n1829__), .dinb(new_new_n1796__), .dout(new_new_n1058__));
  or1   g0435(.dina(new_new_n1832__), .dinb(new_new_n1802__), .dout(new_new_n1059__));
  or1   g0436(.dina(new_new_n1058__), .dinb(new_new_n611__), .dout(new_new_n1060__));
  or1   g0437(.dina(new_new_n1059__), .dinb(new_new_n610__), .dout(new_new_n1061__));
  and1  g0438(.dina(new_new_n1061__), .dinb(new_new_n1060__), .dout(new_new_n1062__));
  and1  g0439(.dina(new_new_n1829__), .dinb(new_new_n1806__), .dout(new_new_n1063__));
  or1   g0440(.dina(new_new_n1832__), .dinb(new_new_n1810__), .dout(new_new_n1064__));
  or1   g0441(.dina(new_new_n1063__), .dinb(new_new_n615__), .dout(new_new_n1065__));
  or1   g0442(.dina(new_new_n1064__), .dinb(new_new_n614__), .dout(new_new_n1066__));
  and1  g0443(.dina(new_new_n1066__), .dinb(new_new_n1065__), .dout(new_new_n1067__));
  and1  g0444(.dina(new_new_n1830__), .dinb(new_new_n1814__), .dout(new_new_n1068__));
  or1   g0445(.dina(new_new_n1833__), .dinb(new_new_n1819__), .dout(new_new_n1069__));
  or1   g0446(.dina(new_new_n1068__), .dinb(new_new_n619__), .dout(new_new_n1070__));
  or1   g0447(.dina(new_new_n1069__), .dinb(new_new_n618__), .dout(new_new_n1071__));
  and1  g0448(.dina(new_new_n1071__), .dinb(new_new_n1070__), .dout(new_new_n1072__));
  and1  g0449(.dina(new_new_n1830__), .dinb(new_new_n1823__), .dout(new_new_n1073__));
  or1   g0450(.dina(new_new_n1833__), .dinb(new_new_n1826__), .dout(new_new_n1074__));
  or1   g0451(.dina(new_new_n1073__), .dinb(new_new_n623__), .dout(new_new_n1075__));
  or1   g0452(.dina(new_new_n1074__), .dinb(new_new_n622__), .dout(new_new_n1076__));
  and1  g0453(.dina(new_new_n1076__), .dinb(new_new_n1075__), .dout(new_new_n1077__));
  and1  g0454(.dina(new_new_n826__), .dinb(new_new_n825__), .dout(new_new_n1078__));
  or1   g0455(.dina(new_new_n827__), .dinb(new_new_n824__), .dout(new_new_n1079__));
  and1  g0456(.dina(new_new_n1078__), .dinb(new_new_n1788__), .dout(new_new_n1080__));
  or1   g0457(.dina(new_new_n1079__), .dinb(new_new_n1791__), .dout(new_new_n1081__));
  and1  g0458(.dina(new_new_n1835__), .dinb(new_new_n1797__), .dout(new_new_n1082__));
  or1   g0459(.dina(new_new_n1838__), .dinb(new_new_n1803__), .dout(new_new_n1083__));
  or1   g0460(.dina(new_new_n1082__), .dinb(new_new_n627__), .dout(new_new_n1084__));
  or1   g0461(.dina(new_new_n1083__), .dinb(new_new_n626__), .dout(new_new_n1085__));
  and1  g0462(.dina(new_new_n1085__), .dinb(new_new_n1084__), .dout(new_new_n1086__));
  and1  g0463(.dina(new_new_n1835__), .dinb(new_new_n1805__), .dout(new_new_n1087__));
  or1   g0464(.dina(new_new_n1838__), .dinb(new_new_n1809__), .dout(new_new_n1088__));
  or1   g0465(.dina(new_new_n1087__), .dinb(new_new_n631__), .dout(new_new_n1089__));
  or1   g0466(.dina(new_new_n1088__), .dinb(new_new_n630__), .dout(new_new_n1090__));
  and1  g0467(.dina(new_new_n1090__), .dinb(new_new_n1089__), .dout(new_new_n1091__));
  and1  g0468(.dina(new_new_n1836__), .dinb(new_new_n1815__), .dout(new_new_n1092__));
  or1   g0469(.dina(new_new_n1839__), .dinb(new_new_n1820__), .dout(new_new_n1093__));
  or1   g0470(.dina(new_new_n1092__), .dinb(new_new_n635__), .dout(new_new_n1094__));
  or1   g0471(.dina(new_new_n1093__), .dinb(new_new_n634__), .dout(new_new_n1095__));
  and1  g0472(.dina(new_new_n1095__), .dinb(new_new_n1094__), .dout(new_new_n1096__));
  and1  g0473(.dina(new_new_n1836__), .dinb(new_new_n1824__), .dout(new_new_n1097__));
  or1   g0474(.dina(new_new_n1839__), .dinb(new_new_n1827__), .dout(new_new_n1098__));
  or1   g0475(.dina(new_new_n1097__), .dinb(new_new_n639__), .dout(new_new_n1099__));
  or1   g0476(.dina(new_new_n1098__), .dinb(new_new_n638__), .dout(new_new_n1100__));
  and1  g0477(.dina(new_new_n1100__), .dinb(new_new_n1099__), .dout(new_new_n1101__));
  and1  g0478(.dina(new_new_n846__), .dinb(new_new_n842__), .dout(new_new_n1102__));
  or1   g0479(.dina(new_new_n847__), .dinb(new_new_n843__), .dout(new_new_n1103__));
  and1  g0480(.dina(new_new_n1102__), .dinb(new_new_n1788__), .dout(new_new_n1104__));
  or1   g0481(.dina(new_new_n1103__), .dinb(new_new_n1791__), .dout(new_new_n1105__));
  and1  g0482(.dina(new_new_n1841__), .dinb(new_new_n1797__), .dout(new_new_n1106__));
  or1   g0483(.dina(new_new_n1844__), .dinb(new_new_n1803__), .dout(new_new_n1107__));
  or1   g0484(.dina(new_new_n1106__), .dinb(new_new_n643__), .dout(new_new_n1108__));
  or1   g0485(.dina(new_new_n1107__), .dinb(new_new_n642__), .dout(new_new_n1109__));
  and1  g0486(.dina(new_new_n1109__), .dinb(new_new_n1108__), .dout(new_new_n1110__));
  and1  g0487(.dina(new_new_n1841__), .dinb(new_new_n1807__), .dout(new_new_n1111__));
  or1   g0488(.dina(new_new_n1844__), .dinb(new_new_n1811__), .dout(new_new_n1112__));
  or1   g0489(.dina(new_new_n1111__), .dinb(new_new_n647__), .dout(new_new_n1113__));
  or1   g0490(.dina(new_new_n1112__), .dinb(new_new_n646__), .dout(new_new_n1114__));
  and1  g0491(.dina(new_new_n1114__), .dinb(new_new_n1113__), .dout(new_new_n1115__));
  and1  g0492(.dina(new_new_n1842__), .dinb(new_new_n1815__), .dout(new_new_n1116__));
  or1   g0493(.dina(new_new_n1845__), .dinb(new_new_n1820__), .dout(new_new_n1117__));
  or1   g0494(.dina(new_new_n1116__), .dinb(new_new_n651__), .dout(new_new_n1118__));
  or1   g0495(.dina(new_new_n1117__), .dinb(new_new_n650__), .dout(new_new_n1119__));
  and1  g0496(.dina(new_new_n1119__), .dinb(new_new_n1118__), .dout(new_new_n1120__));
  and1  g0497(.dina(new_new_n1842__), .dinb(new_new_n1824__), .dout(new_new_n1121__));
  or1   g0498(.dina(new_new_n1845__), .dinb(new_new_n1827__), .dout(new_new_n1122__));
  or1   g0499(.dina(new_new_n1121__), .dinb(new_new_n655__), .dout(new_new_n1123__));
  or1   g0500(.dina(new_new_n1122__), .dinb(new_new_n654__), .dout(new_new_n1124__));
  and1  g0501(.dina(new_new_n1124__), .dinb(new_new_n1123__), .dout(new_new_n1125__));
  and1  g0502(.dina(new_new_n1847__), .dinb(new_new_n832__), .dout(new_new_n1126__));
  or1   g0503(.dina(new_new_n1850__), .dinb(new_new_n833__), .dout(new_new_n1127__));
  and1  g0504(.dina(new_new_n1126__), .dinb(new_new_n1816__), .dout(new_new_n1128__));
  or1   g0505(.dina(new_new_n1127__), .dinb(new_new_n1821__), .dout(new_new_n1129__));
  and1  g0506(.dina(new_new_n1853__), .dinb(new_new_n1856__), .dout(new_new_n1130__));
  or1   g0507(.dina(new_new_n1859__), .dinb(new_new_n1862__), .dout(new_new_n1131__));
  or1   g0508(.dina(new_new_n1130__), .dinb(new_new_n659__), .dout(new_new_n1132__));
  or1   g0509(.dina(new_new_n1131__), .dinb(new_new_n658__), .dout(new_new_n1133__));
  and1  g0510(.dina(new_new_n1133__), .dinb(new_new_n1132__), .dout(new_new_n1134__));
  and1  g0511(.dina(new_new_n1853__), .dinb(new_new_n1865__), .dout(new_new_n1135__));
  or1   g0512(.dina(new_new_n1859__), .dinb(new_new_n1868__), .dout(new_new_n1136__));
  or1   g0513(.dina(new_new_n1135__), .dinb(new_new_n663__), .dout(new_new_n1137__));
  or1   g0514(.dina(new_new_n1136__), .dinb(new_new_n662__), .dout(new_new_n1138__));
  and1  g0515(.dina(new_new_n1138__), .dinb(new_new_n1137__), .dout(new_new_n1139__));
  and1  g0516(.dina(new_new_n1854__), .dinb(new_new_n1871__), .dout(new_new_n1140__));
  or1   g0517(.dina(new_new_n1860__), .dinb(new_new_n1874__), .dout(new_new_n1141__));
  or1   g0518(.dina(new_new_n1140__), .dinb(new_new_n667__), .dout(new_new_n1142__));
  or1   g0519(.dina(new_new_n1141__), .dinb(new_new_n666__), .dout(new_new_n1143__));
  and1  g0520(.dina(new_new_n1143__), .dinb(new_new_n1142__), .dout(new_new_n1144__));
  and1  g0521(.dina(new_new_n1854__), .dinb(new_new_n1877__), .dout(new_new_n1145__));
  or1   g0522(.dina(new_new_n1860__), .dinb(new_new_n1880__), .dout(new_new_n1146__));
  or1   g0523(.dina(new_new_n1145__), .dinb(new_new_n671__), .dout(new_new_n1147__));
  or1   g0524(.dina(new_new_n1146__), .dinb(new_new_n670__), .dout(new_new_n1148__));
  and1  g0525(.dina(new_new_n1148__), .dinb(new_new_n1147__), .dout(new_new_n1149__));
  and1  g0526(.dina(new_new_n820__), .dinb(new_new_n818__), .dout(new_new_n1150__));
  or1   g0527(.dina(new_new_n821__), .dinb(new_new_n819__), .dout(new_new_n1151__));
  and1  g0528(.dina(new_new_n1150__), .dinb(new_new_n1847__), .dout(new_new_n1152__));
  or1   g0529(.dina(new_new_n1151__), .dinb(new_new_n1850__), .dout(new_new_n1153__));
  and1  g0530(.dina(new_new_n1883__), .dinb(new_new_n1856__), .dout(new_new_n1154__));
  or1   g0531(.dina(new_new_n1886__), .dinb(new_new_n1862__), .dout(new_new_n1155__));
  or1   g0532(.dina(new_new_n1154__), .dinb(new_new_n675__), .dout(new_new_n1156__));
  or1   g0533(.dina(new_new_n1155__), .dinb(new_new_n674__), .dout(new_new_n1157__));
  and1  g0534(.dina(new_new_n1157__), .dinb(new_new_n1156__), .dout(new_new_n1158__));
  and1  g0535(.dina(new_new_n1883__), .dinb(new_new_n1865__), .dout(new_new_n1159__));
  or1   g0536(.dina(new_new_n1886__), .dinb(new_new_n1868__), .dout(new_new_n1160__));
  or1   g0537(.dina(new_new_n1159__), .dinb(new_new_n679__), .dout(new_new_n1161__));
  or1   g0538(.dina(new_new_n1160__), .dinb(new_new_n678__), .dout(new_new_n1162__));
  and1  g0539(.dina(new_new_n1162__), .dinb(new_new_n1161__), .dout(new_new_n1163__));
  and1  g0540(.dina(new_new_n1884__), .dinb(new_new_n1871__), .dout(new_new_n1164__));
  or1   g0541(.dina(new_new_n1887__), .dinb(new_new_n1874__), .dout(new_new_n1165__));
  or1   g0542(.dina(new_new_n1164__), .dinb(new_new_n683__), .dout(new_new_n1166__));
  or1   g0543(.dina(new_new_n1165__), .dinb(new_new_n682__), .dout(new_new_n1167__));
  and1  g0544(.dina(new_new_n1167__), .dinb(new_new_n1166__), .dout(new_new_n1168__));
  and1  g0545(.dina(new_new_n1884__), .dinb(new_new_n1877__), .dout(new_new_n1169__));
  or1   g0546(.dina(new_new_n1887__), .dinb(new_new_n1880__), .dout(new_new_n1170__));
  or1   g0547(.dina(new_new_n1169__), .dinb(new_new_n687__), .dout(new_new_n1171__));
  or1   g0548(.dina(new_new_n1170__), .dinb(new_new_n686__), .dout(new_new_n1172__));
  and1  g0549(.dina(new_new_n1172__), .dinb(new_new_n1171__), .dout(new_new_n1173__));
  and1  g0550(.dina(new_new_n830__), .dinb(new_new_n1816__), .dout(new_new_n1174__));
  or1   g0551(.dina(new_new_n831__), .dinb(new_new_n1821__), .dout(new_new_n1175__));
  and1  g0552(.dina(new_new_n1174__), .dinb(new_new_n1848__), .dout(new_new_n1176__));
  or1   g0553(.dina(new_new_n1175__), .dinb(new_new_n1851__), .dout(new_new_n1177__));
  and1  g0554(.dina(new_new_n1889__), .dinb(new_new_n1857__), .dout(new_new_n1178__));
  or1   g0555(.dina(new_new_n1892__), .dinb(new_new_n1863__), .dout(new_new_n1179__));
  or1   g0556(.dina(new_new_n1178__), .dinb(new_new_n691__), .dout(new_new_n1180__));
  or1   g0557(.dina(new_new_n1179__), .dinb(new_new_n690__), .dout(new_new_n1181__));
  and1  g0558(.dina(new_new_n1181__), .dinb(new_new_n1180__), .dout(new_new_n1182__));
  and1  g0559(.dina(new_new_n1889__), .dinb(new_new_n1866__), .dout(new_new_n1183__));
  or1   g0560(.dina(new_new_n1892__), .dinb(new_new_n1869__), .dout(new_new_n1184__));
  or1   g0561(.dina(new_new_n1183__), .dinb(new_new_n695__), .dout(new_new_n1185__));
  or1   g0562(.dina(new_new_n1184__), .dinb(new_new_n694__), .dout(new_new_n1186__));
  and1  g0563(.dina(new_new_n1186__), .dinb(new_new_n1185__), .dout(new_new_n1187__));
  and1  g0564(.dina(new_new_n1890__), .dinb(new_new_n1872__), .dout(new_new_n1188__));
  or1   g0565(.dina(new_new_n1893__), .dinb(new_new_n1875__), .dout(new_new_n1189__));
  or1   g0566(.dina(new_new_n1188__), .dinb(new_new_n699__), .dout(new_new_n1190__));
  or1   g0567(.dina(new_new_n1189__), .dinb(new_new_n698__), .dout(new_new_n1191__));
  and1  g0568(.dina(new_new_n1191__), .dinb(new_new_n1190__), .dout(new_new_n1192__));
  and1  g0569(.dina(new_new_n1890__), .dinb(new_new_n1878__), .dout(new_new_n1193__));
  or1   g0570(.dina(new_new_n1893__), .dinb(new_new_n1881__), .dout(new_new_n1194__));
  or1   g0571(.dina(new_new_n1193__), .dinb(new_new_n703__), .dout(new_new_n1195__));
  or1   g0572(.dina(new_new_n1194__), .dinb(new_new_n702__), .dout(new_new_n1196__));
  and1  g0573(.dina(new_new_n1196__), .dinb(new_new_n1195__), .dout(new_new_n1197__));
  and1  g0574(.dina(new_new_n828__), .dinb(new_new_n1807__), .dout(new_new_n1198__));
  or1   g0575(.dina(new_new_n829__), .dinb(new_new_n1811__), .dout(new_new_n1199__));
  and1  g0576(.dina(new_new_n1198__), .dinb(new_new_n1848__), .dout(new_new_n1200__));
  or1   g0577(.dina(new_new_n1199__), .dinb(new_new_n1851__), .dout(new_new_n1201__));
  and1  g0578(.dina(new_new_n1895__), .dinb(new_new_n1857__), .dout(new_new_n1202__));
  or1   g0579(.dina(new_new_n1898__), .dinb(new_new_n1863__), .dout(new_new_n1203__));
  or1   g0580(.dina(new_new_n1202__), .dinb(new_new_n707__), .dout(new_new_n1204__));
  or1   g0581(.dina(new_new_n1203__), .dinb(new_new_n706__), .dout(new_new_n1205__));
  and1  g0582(.dina(new_new_n1205__), .dinb(new_new_n1204__), .dout(new_new_n1206__));
  and1  g0583(.dina(new_new_n1895__), .dinb(new_new_n1866__), .dout(new_new_n1207__));
  or1   g0584(.dina(new_new_n1898__), .dinb(new_new_n1869__), .dout(new_new_n1208__));
  or1   g0585(.dina(new_new_n1207__), .dinb(new_new_n711__), .dout(new_new_n1209__));
  or1   g0586(.dina(new_new_n1208__), .dinb(new_new_n710__), .dout(new_new_n1210__));
  and1  g0587(.dina(new_new_n1210__), .dinb(new_new_n1209__), .dout(new_new_n1211__));
  and1  g0588(.dina(new_new_n1896__), .dinb(new_new_n1872__), .dout(new_new_n1212__));
  or1   g0589(.dina(new_new_n1899__), .dinb(new_new_n1875__), .dout(new_new_n1213__));
  or1   g0590(.dina(new_new_n1212__), .dinb(new_new_n715__), .dout(new_new_n1214__));
  or1   g0591(.dina(new_new_n1213__), .dinb(new_new_n714__), .dout(new_new_n1215__));
  and1  g0592(.dina(new_new_n1215__), .dinb(new_new_n1214__), .dout(new_new_n1216__));
  and1  g0593(.dina(new_new_n1896__), .dinb(new_new_n1878__), .dout(new_new_n1217__));
  or1   g0594(.dina(new_new_n1899__), .dinb(new_new_n1881__), .dout(new_new_n1218__));
  or1   g0595(.dina(new_new_n1217__), .dinb(new_new_n719__), .dout(new_new_n1219__));
  or1   g0596(.dina(new_new_n1218__), .dinb(new_new_n718__), .dout(new_new_n1220__));
  and1  g0597(.dina(new_new_n1220__), .dinb(new_new_n1219__), .dout(new_new_n1221__));
  and1  g0598(.dina(new_new_n917__), .dinb(new_new_n915__), .dout(new_new_n1222__));
  or1   g0599(.dina(new_new_n916__), .dinb(new_new_n914__), .dout(new_new_n1223__));
  and1  g0600(.dina(new_new_n921__), .dinb(new_new_n919__), .dout(new_new_n1224__));
  or1   g0601(.dina(new_new_n920__), .dinb(new_new_n918__), .dout(new_new_n1225__));
  and1  g0602(.dina(new_new_n925__), .dinb(new_new_n923__), .dout(new_new_n1226__));
  or1   g0603(.dina(new_new_n924__), .dinb(new_new_n922__), .dout(new_new_n1227__));
  and1  g0604(.dina(new_new_n929__), .dinb(new_new_n927__), .dout(new_new_n1228__));
  or1   g0605(.dina(new_new_n928__), .dinb(new_new_n926__), .dout(new_new_n1229__));
  and1  g0606(.dina(new_new_n933__), .dinb(new_new_n931__), .dout(new_new_n1230__));
  or1   g0607(.dina(new_new_n932__), .dinb(new_new_n930__), .dout(new_new_n1231__));
  and1  g0608(.dina(new_new_n937__), .dinb(new_new_n935__), .dout(new_new_n1232__));
  or1   g0609(.dina(new_new_n936__), .dinb(new_new_n934__), .dout(new_new_n1233__));
  and1  g0610(.dina(new_new_n941__), .dinb(new_new_n939__), .dout(new_new_n1234__));
  or1   g0611(.dina(new_new_n940__), .dinb(new_new_n938__), .dout(new_new_n1235__));
  and1  g0612(.dina(new_new_n945__), .dinb(new_new_n943__), .dout(new_new_n1236__));
  or1   g0613(.dina(new_new_n944__), .dinb(new_new_n942__), .dout(new_new_n1237__));
  or1   g0614(.dina(new_new_n1901__), .dinb(new_new_n1222__), .dout(new_new_n1238__));
  or1   g0615(.dina(new_new_n1228__), .dinb(new_new_n1903__), .dout(new_new_n1239__));
  or1   g0616(.dina(new_new_n1905__), .dinb(new_new_n1907__), .dout(new_new_n1240__));
  and1  g0617(.dina(new_new_n1905__), .dinb(new_new_n1907__), .dout(new_new_n1241__));
  or1   g0618(.dina(new_new_n1909__), .dinb(new_new_n1911__), .dout(new_new_n1242__));
  or1   g0619(.dina(new_new_n1913__), .dinb(new_new_n1915__), .dout(new_new_n1243__));
  or1   g0620(.dina(new_new_n1916__), .dinb(new_new_n1918__), .dout(new_new_n1244__));
  or1   g0621(.dina(new_new_n1920__), .dinb(new_new_n1918__), .dout(new_new_n1245__));
  or1   g0622(.dina(new_new_n1921__), .dinb(new_new_n1224__), .dout(new_new_n1246__));
  or1   g0623(.dina(new_new_n1922__), .dinb(new_new_n1920__), .dout(new_new_n1247__));
  and1  g0624(.dina(new_new_n1913__), .dinb(new_new_n1915__), .dout(new_new_n1248__));
  or1   g0625(.dina(new_new_n1924__), .dinb(new_new_n1926__), .dout(new_new_n1249__));
  or1   g0626(.dina(new_new_n1921__), .dinb(new_new_n1226__), .dout(new_new_n1250__));
  and1  g0627(.dina(new_new_n1250__), .dinb(new_new_n1927__), .dout(new_new_n1251__));
  or1   g0628(.dina(new_new_n1251__), .dinb(new_new_n1901__), .dout(new_new_n1252__));
  and1  g0629(.dina(new_new_n1928__), .dinb(new_new_n1929__), .dout(new_new_n1253__));
  or1   g0630(.dina(new_new_n1253__), .dinb(new_new_n1903__), .dout(new_new_n1254__));
  and1  g0631(.dina(new_new_n1914__), .dinb(new_new_n1911__), .dout(new_new_n1255__));
  and1  g0632(.dina(new_new_n1926__), .dinb(new_new_n1906__), .dout(new_new_n1256__));
  and1  g0633(.dina(new_new_n1904__), .dinb(new_new_n1924__), .dout(new_new_n1257__));
  and1  g0634(.dina(new_new_n1909__), .dinb(new_new_n1912__), .dout(new_new_n1258__));
  and1  g0635(.dina(new_new_n1930__), .dinb(new_new_n1931__), .dout(new_new_n1259__));
  or1   g0636(.dina(new_new_n1259__), .dinb(new_new_n1932__), .dout(new_new_n1260__));
  and1  g0637(.dina(new_new_n1933__), .dinb(new_new_n1241__), .dout(new_new_n1261__));
  or1   g0638(.dina(new_new_n1261__), .dinb(new_new_n1248__), .dout(new_new_n1262__));
  and1  g0639(.dina(new_new_n1262__), .dinb(new_new_n1260__), .dout(new_new_n1263__));
  and1  g0640(.dina(new_new_n1934__), .dinb(new_new_n1935__), .dout(new_new_n1264__));
  or1   g0641(.dina(new_new_n1936__), .dinb(new_new_n1937__), .dout(new_new_n1265__));
  and1  g0642(.dina(new_new_n1936__), .dinb(new_new_n1937__), .dout(new_new_n1266__));
  or1   g0643(.dina(new_new_n1934__), .dinb(new_new_n1935__), .dout(new_new_n1267__));
  and1  g0644(.dina(new_new_n1267__), .dinb(new_new_n1265__), .dout(new_new_n1268__));
  or1   g0645(.dina(new_new_n1266__), .dinb(new_new_n1264__), .dout(new_new_n1269__));
  and1  g0646(.dina(new_new_n1940__), .dinb(new_new_n946__), .dout(new_new_n1270__));
  or1   g0647(.dina(new_new_n1947__), .dinb(new_new_n947__), .dout(new_new_n1271__));
  and1  g0648(.dina(new_new_n1270__), .dinb(new_new_n1269__), .dout(new_new_n1272__));
  and1  g0649(.dina(new_new_n1271__), .dinb(new_new_n1268__), .dout(new_new_n1273__));
  or1   g0650(.dina(new_new_n1273__), .dinb(new_new_n1272__), .dout(new_new_n1274__));
  and1  g0651(.dina(new_new_n1952__), .dinb(new_new_n1953__), .dout(new_new_n1275__));
  or1   g0652(.dina(new_new_n1954__), .dinb(new_new_n1955__), .dout(new_new_n1276__));
  and1  g0653(.dina(new_new_n1954__), .dinb(new_new_n1955__), .dout(new_new_n1277__));
  or1   g0654(.dina(new_new_n1952__), .dinb(new_new_n1953__), .dout(new_new_n1278__));
  and1  g0655(.dina(new_new_n1278__), .dinb(new_new_n1276__), .dout(new_new_n1279__));
  or1   g0656(.dina(new_new_n1277__), .dinb(new_new_n1275__), .dout(new_new_n1280__));
  and1  g0657(.dina(new_new_n1956__), .dinb(new_new_n1957__), .dout(new_new_n1281__));
  or1   g0658(.dina(new_new_n1958__), .dinb(new_new_n1959__), .dout(new_new_n1282__));
  and1  g0659(.dina(new_new_n1958__), .dinb(new_new_n1959__), .dout(new_new_n1283__));
  or1   g0660(.dina(new_new_n1956__), .dinb(new_new_n1957__), .dout(new_new_n1284__));
  and1  g0661(.dina(new_new_n1284__), .dinb(new_new_n1282__), .dout(new_new_n1285__));
  or1   g0662(.dina(new_new_n1283__), .dinb(new_new_n1281__), .dout(new_new_n1286__));
  and1  g0663(.dina(new_new_n1960__), .dinb(new_new_n1961__), .dout(new_new_n1287__));
  and1  g0664(.dina(new_new_n1962__), .dinb(new_new_n1963__), .dout(new_new_n1288__));
  or1   g0665(.dina(new_new_n1288__), .dinb(new_new_n1287__), .dout(new_new_n1289__));
  and1  g0666(.dina(new_new_n1964__), .dinb(new_new_n1965__), .dout(new_new_n1290__));
  or1   g0667(.dina(new_new_n1964__), .dinb(new_new_n1965__), .dout(new_new_n1291__));
  and1  g0668(.dina(new_new_n1966__), .dinb(new_new_n1967__), .dout(new_new_n1292__));
  or1   g0669(.dina(new_new_n1968__), .dinb(new_new_n1969__), .dout(new_new_n1293__));
  and1  g0670(.dina(new_new_n1968__), .dinb(new_new_n1969__), .dout(new_new_n1294__));
  or1   g0671(.dina(new_new_n1966__), .dinb(new_new_n1967__), .dout(new_new_n1295__));
  and1  g0672(.dina(new_new_n1295__), .dinb(new_new_n1293__), .dout(new_new_n1296__));
  or1   g0673(.dina(new_new_n1294__), .dinb(new_new_n1292__), .dout(new_new_n1297__));
  and1  g0674(.dina(new_new_n1940__), .dinb(new_new_n948__), .dout(new_new_n1298__));
  or1   g0675(.dina(new_new_n1947__), .dinb(new_new_n949__), .dout(new_new_n1299__));
  and1  g0676(.dina(new_new_n1298__), .dinb(new_new_n1297__), .dout(new_new_n1300__));
  and1  g0677(.dina(new_new_n1299__), .dinb(new_new_n1296__), .dout(new_new_n1301__));
  or1   g0678(.dina(new_new_n1301__), .dinb(new_new_n1300__), .dout(new_new_n1302__));
  and1  g0679(.dina(new_new_n1970__), .dinb(new_new_n1971__), .dout(new_new_n1303__));
  or1   g0680(.dina(new_new_n1972__), .dinb(new_new_n1973__), .dout(new_new_n1304__));
  and1  g0681(.dina(new_new_n1972__), .dinb(new_new_n1973__), .dout(new_new_n1305__));
  or1   g0682(.dina(new_new_n1970__), .dinb(new_new_n1971__), .dout(new_new_n1306__));
  and1  g0683(.dina(new_new_n1306__), .dinb(new_new_n1304__), .dout(new_new_n1307__));
  or1   g0684(.dina(new_new_n1305__), .dinb(new_new_n1303__), .dout(new_new_n1308__));
  and1  g0685(.dina(new_new_n1974__), .dinb(new_new_n1975__), .dout(new_new_n1309__));
  or1   g0686(.dina(new_new_n1976__), .dinb(new_new_n1977__), .dout(new_new_n1310__));
  and1  g0687(.dina(new_new_n1976__), .dinb(new_new_n1977__), .dout(new_new_n1311__));
  or1   g0688(.dina(new_new_n1974__), .dinb(new_new_n1975__), .dout(new_new_n1312__));
  and1  g0689(.dina(new_new_n1312__), .dinb(new_new_n1310__), .dout(new_new_n1313__));
  or1   g0690(.dina(new_new_n1311__), .dinb(new_new_n1309__), .dout(new_new_n1314__));
  and1  g0691(.dina(new_new_n1978__), .dinb(new_new_n1979__), .dout(new_new_n1315__));
  and1  g0692(.dina(new_new_n1980__), .dinb(new_new_n1981__), .dout(new_new_n1316__));
  or1   g0693(.dina(new_new_n1316__), .dinb(new_new_n1315__), .dout(new_new_n1317__));
  and1  g0694(.dina(new_new_n1982__), .dinb(new_new_n1983__), .dout(new_new_n1318__));
  or1   g0695(.dina(new_new_n1982__), .dinb(new_new_n1983__), .dout(new_new_n1319__));
  and1  g0696(.dina(new_new_n1984__), .dinb(new_new_n1985__), .dout(new_new_n1320__));
  or1   g0697(.dina(new_new_n1986__), .dinb(new_new_n1987__), .dout(new_new_n1321__));
  and1  g0698(.dina(new_new_n1986__), .dinb(new_new_n1987__), .dout(new_new_n1322__));
  or1   g0699(.dina(new_new_n1984__), .dinb(new_new_n1985__), .dout(new_new_n1323__));
  and1  g0700(.dina(new_new_n1323__), .dinb(new_new_n1321__), .dout(new_new_n1324__));
  or1   g0701(.dina(new_new_n1322__), .dinb(new_new_n1320__), .dout(new_new_n1325__));
  and1  g0702(.dina(new_new_n1941__), .dinb(new_new_n950__), .dout(new_new_n1326__));
  or1   g0703(.dina(new_new_n1948__), .dinb(new_new_n951__), .dout(new_new_n1327__));
  and1  g0704(.dina(new_new_n1326__), .dinb(new_new_n1325__), .dout(new_new_n1328__));
  and1  g0705(.dina(new_new_n1327__), .dinb(new_new_n1324__), .dout(new_new_n1329__));
  or1   g0706(.dina(new_new_n1329__), .dinb(new_new_n1328__), .dout(new_new_n1330__));
  and1  g0707(.dina(new_new_n1978__), .dinb(new_new_n1961__), .dout(new_new_n1331__));
  and1  g0708(.dina(new_new_n1980__), .dinb(new_new_n1963__), .dout(new_new_n1332__));
  or1   g0709(.dina(new_new_n1332__), .dinb(new_new_n1331__), .dout(new_new_n1333__));
  and1  g0710(.dina(new_new_n1988__), .dinb(new_new_n1989__), .dout(new_new_n1334__));
  or1   g0711(.dina(new_new_n1988__), .dinb(new_new_n1989__), .dout(new_new_n1335__));
  and1  g0712(.dina(new_new_n1990__), .dinb(new_new_n1991__), .dout(new_new_n1336__));
  or1   g0713(.dina(new_new_n1992__), .dinb(new_new_n1993__), .dout(new_new_n1337__));
  and1  g0714(.dina(new_new_n1992__), .dinb(new_new_n1993__), .dout(new_new_n1338__));
  or1   g0715(.dina(new_new_n1990__), .dinb(new_new_n1991__), .dout(new_new_n1339__));
  and1  g0716(.dina(new_new_n1339__), .dinb(new_new_n1337__), .dout(new_new_n1340__));
  or1   g0717(.dina(new_new_n1338__), .dinb(new_new_n1336__), .dout(new_new_n1341__));
  and1  g0718(.dina(new_new_n1941__), .dinb(new_new_n952__), .dout(new_new_n1342__));
  or1   g0719(.dina(new_new_n1948__), .dinb(new_new_n953__), .dout(new_new_n1343__));
  and1  g0720(.dina(new_new_n1342__), .dinb(new_new_n1341__), .dout(new_new_n1344__));
  and1  g0721(.dina(new_new_n1343__), .dinb(new_new_n1340__), .dout(new_new_n1345__));
  or1   g0722(.dina(new_new_n1345__), .dinb(new_new_n1344__), .dout(new_new_n1346__));
  and1  g0723(.dina(new_new_n1981__), .dinb(new_new_n1962__), .dout(new_new_n1347__));
  and1  g0724(.dina(new_new_n1979__), .dinb(new_new_n1960__), .dout(new_new_n1348__));
  or1   g0725(.dina(new_new_n1348__), .dinb(new_new_n1347__), .dout(new_new_n1349__));
  and1  g0726(.dina(new_new_n1994__), .dinb(new_new_n1995__), .dout(new_new_n1350__));
  or1   g0727(.dina(new_new_n1994__), .dinb(new_new_n1995__), .dout(new_new_n1351__));
  and1  g0728(.dina(new_new_n1996__), .dinb(new_new_n1997__), .dout(new_new_n1352__));
  or1   g0729(.dina(new_new_n1998__), .dinb(new_new_n1999__), .dout(new_new_n1353__));
  and1  g0730(.dina(new_new_n1998__), .dinb(new_new_n1999__), .dout(new_new_n1354__));
  or1   g0731(.dina(new_new_n1996__), .dinb(new_new_n1997__), .dout(new_new_n1355__));
  and1  g0732(.dina(new_new_n1355__), .dinb(new_new_n1353__), .dout(new_new_n1356__));
  or1   g0733(.dina(new_new_n1354__), .dinb(new_new_n1352__), .dout(new_new_n1357__));
  and1  g0734(.dina(new_new_n1943__), .dinb(new_new_n954__), .dout(new_new_n1358__));
  or1   g0735(.dina(new_new_n1950__), .dinb(new_new_n955__), .dout(new_new_n1359__));
  and1  g0736(.dina(new_new_n1358__), .dinb(new_new_n1357__), .dout(new_new_n1360__));
  and1  g0737(.dina(new_new_n1359__), .dinb(new_new_n1356__), .dout(new_new_n1361__));
  or1   g0738(.dina(new_new_n1361__), .dinb(new_new_n1360__), .dout(new_new_n1362__));
  and1  g0739(.dina(new_new_n2000__), .dinb(new_new_n2001__), .dout(new_new_n1363__));
  or1   g0740(.dina(new_new_n2002__), .dinb(new_new_n2003__), .dout(new_new_n1364__));
  and1  g0741(.dina(new_new_n2002__), .dinb(new_new_n2003__), .dout(new_new_n1365__));
  or1   g0742(.dina(new_new_n2000__), .dinb(new_new_n2001__), .dout(new_new_n1366__));
  and1  g0743(.dina(new_new_n1366__), .dinb(new_new_n1364__), .dout(new_new_n1367__));
  or1   g0744(.dina(new_new_n1365__), .dinb(new_new_n1363__), .dout(new_new_n1368__));
  and1  g0745(.dina(new_new_n2004__), .dinb(new_new_n2005__), .dout(new_new_n1369__));
  or1   g0746(.dina(new_new_n2006__), .dinb(new_new_n2007__), .dout(new_new_n1370__));
  and1  g0747(.dina(new_new_n2006__), .dinb(new_new_n2007__), .dout(new_new_n1371__));
  or1   g0748(.dina(new_new_n2004__), .dinb(new_new_n2005__), .dout(new_new_n1372__));
  and1  g0749(.dina(new_new_n1372__), .dinb(new_new_n1370__), .dout(new_new_n1373__));
  or1   g0750(.dina(new_new_n1371__), .dinb(new_new_n1369__), .dout(new_new_n1374__));
  and1  g0751(.dina(new_new_n2008__), .dinb(new_new_n2009__), .dout(new_new_n1375__));
  and1  g0752(.dina(new_new_n2010__), .dinb(new_new_n2011__), .dout(new_new_n1376__));
  or1   g0753(.dina(new_new_n1376__), .dinb(new_new_n1375__), .dout(new_new_n1377__));
  and1  g0754(.dina(new_new_n2012__), .dinb(new_new_n2013__), .dout(new_new_n1378__));
  or1   g0755(.dina(new_new_n2012__), .dinb(new_new_n2013__), .dout(new_new_n1379__));
  and1  g0756(.dina(new_new_n2014__), .dinb(new_new_n2015__), .dout(new_new_n1380__));
  or1   g0757(.dina(new_new_n2016__), .dinb(new_new_n2017__), .dout(new_new_n1381__));
  and1  g0758(.dina(new_new_n2016__), .dinb(new_new_n2017__), .dout(new_new_n1382__));
  or1   g0759(.dina(new_new_n2014__), .dinb(new_new_n2015__), .dout(new_new_n1383__));
  and1  g0760(.dina(new_new_n1383__), .dinb(new_new_n1381__), .dout(new_new_n1384__));
  or1   g0761(.dina(new_new_n1382__), .dinb(new_new_n1380__), .dout(new_new_n1385__));
  and1  g0762(.dina(new_new_n1943__), .dinb(new_new_n956__), .dout(new_new_n1386__));
  or1   g0763(.dina(new_new_n1950__), .dinb(new_new_n957__), .dout(new_new_n1387__));
  and1  g0764(.dina(new_new_n1386__), .dinb(new_new_n1385__), .dout(new_new_n1388__));
  and1  g0765(.dina(new_new_n1387__), .dinb(new_new_n1384__), .dout(new_new_n1389__));
  or1   g0766(.dina(new_new_n1389__), .dinb(new_new_n1388__), .dout(new_new_n1390__));
  and1  g0767(.dina(new_new_n2018__), .dinb(new_new_n2019__), .dout(new_new_n1391__));
  or1   g0768(.dina(new_new_n2020__), .dinb(new_new_n2021__), .dout(new_new_n1392__));
  and1  g0769(.dina(new_new_n2020__), .dinb(new_new_n2021__), .dout(new_new_n1393__));
  or1   g0770(.dina(new_new_n2018__), .dinb(new_new_n2019__), .dout(new_new_n1394__));
  and1  g0771(.dina(new_new_n1394__), .dinb(new_new_n1392__), .dout(new_new_n1395__));
  or1   g0772(.dina(new_new_n1393__), .dinb(new_new_n1391__), .dout(new_new_n1396__));
  and1  g0773(.dina(new_new_n2022__), .dinb(new_new_n2023__), .dout(new_new_n1397__));
  or1   g0774(.dina(new_new_n2024__), .dinb(new_new_n2025__), .dout(new_new_n1398__));
  and1  g0775(.dina(new_new_n2024__), .dinb(new_new_n2025__), .dout(new_new_n1399__));
  or1   g0776(.dina(new_new_n2022__), .dinb(new_new_n2023__), .dout(new_new_n1400__));
  and1  g0777(.dina(new_new_n1400__), .dinb(new_new_n1398__), .dout(new_new_n1401__));
  or1   g0778(.dina(new_new_n1399__), .dinb(new_new_n1397__), .dout(new_new_n1402__));
  and1  g0779(.dina(new_new_n2026__), .dinb(new_new_n2027__), .dout(new_new_n1403__));
  and1  g0780(.dina(new_new_n2028__), .dinb(new_new_n2029__), .dout(new_new_n1404__));
  or1   g0781(.dina(new_new_n1404__), .dinb(new_new_n1403__), .dout(new_new_n1405__));
  and1  g0782(.dina(new_new_n2030__), .dinb(new_new_n2031__), .dout(new_new_n1406__));
  or1   g0783(.dina(new_new_n2030__), .dinb(new_new_n2031__), .dout(new_new_n1407__));
  and1  g0784(.dina(new_new_n2032__), .dinb(new_new_n2033__), .dout(new_new_n1408__));
  or1   g0785(.dina(new_new_n2034__), .dinb(new_new_n2035__), .dout(new_new_n1409__));
  and1  g0786(.dina(new_new_n2034__), .dinb(new_new_n2035__), .dout(new_new_n1410__));
  or1   g0787(.dina(new_new_n2032__), .dinb(new_new_n2033__), .dout(new_new_n1411__));
  and1  g0788(.dina(new_new_n1411__), .dinb(new_new_n1409__), .dout(new_new_n1412__));
  or1   g0789(.dina(new_new_n1410__), .dinb(new_new_n1408__), .dout(new_new_n1413__));
  and1  g0790(.dina(new_new_n1944__), .dinb(new_new_n958__), .dout(new_new_n1414__));
  or1   g0791(.dina(new_new_n1951__), .dinb(new_new_n959__), .dout(new_new_n1415__));
  and1  g0792(.dina(new_new_n1414__), .dinb(new_new_n1413__), .dout(new_new_n1416__));
  and1  g0793(.dina(new_new_n1415__), .dinb(new_new_n1412__), .dout(new_new_n1417__));
  or1   g0794(.dina(new_new_n1417__), .dinb(new_new_n1416__), .dout(new_new_n1418__));
  and1  g0795(.dina(new_new_n2029__), .dinb(new_new_n2009__), .dout(new_new_n1419__));
  and1  g0796(.dina(new_new_n2027__), .dinb(new_new_n2011__), .dout(new_new_n1420__));
  or1   g0797(.dina(new_new_n1420__), .dinb(new_new_n1419__), .dout(new_new_n1421__));
  and1  g0798(.dina(new_new_n2036__), .dinb(new_new_n2037__), .dout(new_new_n1422__));
  or1   g0799(.dina(new_new_n2036__), .dinb(new_new_n2037__), .dout(new_new_n1423__));
  and1  g0800(.dina(new_new_n2038__), .dinb(new_new_n2039__), .dout(new_new_n1424__));
  or1   g0801(.dina(new_new_n2040__), .dinb(new_new_n2041__), .dout(new_new_n1425__));
  and1  g0802(.dina(new_new_n2040__), .dinb(new_new_n2041__), .dout(new_new_n1426__));
  or1   g0803(.dina(new_new_n2038__), .dinb(new_new_n2039__), .dout(new_new_n1427__));
  and1  g0804(.dina(new_new_n1427__), .dinb(new_new_n1425__), .dout(new_new_n1428__));
  or1   g0805(.dina(new_new_n1426__), .dinb(new_new_n1424__), .dout(new_new_n1429__));
  and1  g0806(.dina(new_new_n1944__), .dinb(new_new_n960__), .dout(new_new_n1430__));
  or1   g0807(.dina(new_new_n1951__), .dinb(new_new_n961__), .dout(new_new_n1431__));
  and1  g0808(.dina(new_new_n1430__), .dinb(new_new_n1429__), .dout(new_new_n1432__));
  and1  g0809(.dina(new_new_n1431__), .dinb(new_new_n1428__), .dout(new_new_n1433__));
  or1   g0810(.dina(new_new_n1433__), .dinb(new_new_n1432__), .dout(new_new_n1434__));
  and1  g0811(.dina(new_new_n2026__), .dinb(new_new_n2010__), .dout(new_new_n1435__));
  and1  g0812(.dina(new_new_n2028__), .dinb(new_new_n2008__), .dout(new_new_n1436__));
  or1   g0813(.dina(new_new_n1436__), .dinb(new_new_n1435__), .dout(new_new_n1437__));
  and1  g0814(.dina(new_new_n2042__), .dinb(new_new_n2043__), .dout(new_new_n1438__));
  or1   g0815(.dina(new_new_n2042__), .dinb(new_new_n2043__), .dout(new_new_n1439__));
  or1   g0816(.dina(new_new_n2045__), .dinb(new_new_n2047__), .dout(new_new_n1440__));
  or1   g0817(.dina(new_new_n2048__), .dinb(new_new_n2049__), .dout(new_new_n1441__));
  and1  g0818(.dina(new_new_n1441__), .dinb(new_new_n1440__), .dout(new_new_n1442__));
  or1   g0819(.dina(new_new_n2051__), .dinb(new_new_n2047__), .dout(new_new_n1443__));
  or1   g0820(.dina(new_new_n2052__), .dinb(new_new_n2049__), .dout(new_new_n1444__));
  and1  g0821(.dina(new_new_n1444__), .dinb(new_new_n1443__), .dout(new_new_n1445__));
  or1   g0822(.dina(new_new_n2054__), .dinb(new_new_n2051__), .dout(new_new_n1446__));
  or1   g0823(.dina(new_new_n2055__), .dinb(new_new_n2052__), .dout(new_new_n1447__));
  and1  g0824(.dina(new_new_n1447__), .dinb(new_new_n1446__), .dout(new_new_n1448__));
  or1   g0825(.dina(new_new_n2057__), .dinb(new_new_n2059__), .dout(new_new_n1449__));
  or1   g0826(.dina(new_new_n2060__), .dinb(new_new_n2061__), .dout(new_new_n1450__));
  and1  g0827(.dina(new_new_n1450__), .dinb(new_new_n1449__), .dout(new_new_n1451__));
  and1  g0828(.dina(new_new_n2062__), .dinb(new_new_n2059__), .dout(new_new_n1452__));
  and1  g0829(.dina(new_new_n2064__), .dinb(new_new_n2061__), .dout(new_new_n1453__));
  or1   g0830(.dina(new_new_n1453__), .dinb(new_new_n1452__), .dout(new_new_n1454__));
  or1   g0831(.dina(new_new_n2066__), .dinb(new_new_n2064__), .dout(new_new_n1455__));
  or1   g0832(.dina(new_new_n2067__), .dinb(new_new_n2062__), .dout(new_new_n1456__));
  and1  g0833(.dina(new_new_n1456__), .dinb(new_new_n1455__), .dout(new_new_n1457__));
  or1   g0834(.dina(new_new_n2054__), .dinb(new_new_n2045__), .dout(new_new_n1458__));
  or1   g0835(.dina(new_new_n2055__), .dinb(new_new_n2048__), .dout(new_new_n1459__));
  and1  g0836(.dina(new_new_n1459__), .dinb(new_new_n1458__), .dout(new_new_n1460__));
  and1  g0837(.dina(new_new_n2067__), .dinb(new_new_n2057__), .dout(new_new_n1461__));
  and1  g0838(.dina(new_new_n2066__), .dinb(new_new_n2060__), .dout(new_new_n1462__));
  or1   g0839(.dina(new_new_n1462__), .dinb(new_new_n1461__), .dout(new_new_n1463__));
  and1  g0840(.dina(new_new_n2068__), .dinb(new_new_n2070__), .dout(new_new_n1464__));
  and1  g0841(.dina(new_new_n2072__), .dinb(new_new_n2073__), .dout(new_new_n1465__));
  or1   g0842(.dina(new_new_n1465__), .dinb(new_new_n1464__), .dout(new_new_n1466__));
  or1   g0843(.dina(new_new_n2075__), .dinb(new_new_n2070__), .dout(new_new_n1467__));
  or1   g0844(.dina(new_new_n2076__), .dinb(new_new_n2073__), .dout(new_new_n1468__));
  and1  g0845(.dina(new_new_n1468__), .dinb(new_new_n1467__), .dout(new_new_n1469__));
  and1  g0846(.dina(new_new_n2077__), .dinb(new_new_n2075__), .dout(new_new_n1470__));
  and1  g0847(.dina(new_new_n2079__), .dinb(new_new_n2076__), .dout(new_new_n1471__));
  or1   g0848(.dina(new_new_n1471__), .dinb(new_new_n1470__), .dout(new_new_n1472__));
  and1  g0849(.dina(new_new_n2080__), .dinb(new_new_n2082__), .dout(new_new_n1473__));
  and1  g0850(.dina(new_new_n2084__), .dinb(new_new_n2085__), .dout(new_new_n1474__));
  or1   g0851(.dina(new_new_n1474__), .dinb(new_new_n1473__), .dout(new_new_n1475__));
  and1  g0852(.dina(new_new_n2086__), .dinb(new_new_n2082__), .dout(new_new_n1476__));
  and1  g0853(.dina(new_new_n2088__), .dinb(new_new_n2085__), .dout(new_new_n1477__));
  or1   g0854(.dina(new_new_n1477__), .dinb(new_new_n1476__), .dout(new_new_n1478__));
  and1  g0855(.dina(new_new_n2089__), .dinb(new_new_n2088__), .dout(new_new_n1479__));
  and1  g0856(.dina(new_new_n2091__), .dinb(new_new_n2086__), .dout(new_new_n1480__));
  or1   g0857(.dina(new_new_n1480__), .dinb(new_new_n1479__), .dout(new_new_n1481__));
  or1   g0858(.dina(new_new_n2079__), .dinb(new_new_n2072__), .dout(new_new_n1482__));
  or1   g0859(.dina(new_new_n2077__), .dinb(new_new_n2068__), .dout(new_new_n1483__));
  and1  g0860(.dina(new_new_n1483__), .dinb(new_new_n1482__), .dout(new_new_n1484__));
  and1  g0861(.dina(new_new_n2089__), .dinb(new_new_n2084__), .dout(new_new_n1485__));
  and1  g0862(.dina(new_new_n2091__), .dinb(new_new_n2080__), .dout(new_new_n1486__));
  or1   g0863(.dina(new_new_n1486__), .dinb(new_new_n1485__), .dout(new_new_n1487__));
  or1   g0864(.dina(new_new_n2093__), .dinb(new_new_n2095__), .dout(new_new_n1488__));
  or1   g0865(.dina(new_new_n2096__), .dinb(new_new_n2097__), .dout(new_new_n1489__));
  and1  g0866(.dina(new_new_n1489__), .dinb(new_new_n1488__), .dout(new_new_n1490__));
  or1   g0867(.dina(new_new_n2099__), .dinb(new_new_n2095__), .dout(new_new_n1491__));
  or1   g0868(.dina(new_new_n2100__), .dinb(new_new_n2097__), .dout(new_new_n1492__));
  and1  g0869(.dina(new_new_n1492__), .dinb(new_new_n1491__), .dout(new_new_n1493__));
  or1   g0870(.dina(new_new_n2102__), .dinb(new_new_n2093__), .dout(new_new_n1494__));
  or1   g0871(.dina(new_new_n2103__), .dinb(new_new_n2096__), .dout(new_new_n1495__));
  and1  g0872(.dina(new_new_n1495__), .dinb(new_new_n1494__), .dout(new_new_n1496__));
  and1  g0873(.dina(new_new_n2104__), .dinb(new_new_n2106__), .dout(new_new_n1497__));
  and1  g0874(.dina(new_new_n2108__), .dinb(new_new_n2109__), .dout(new_new_n1498__));
  or1   g0875(.dina(new_new_n1498__), .dinb(new_new_n1497__), .dout(new_new_n1499__));
  or1   g0876(.dina(new_new_n2111__), .dinb(new_new_n2106__), .dout(new_new_n1500__));
  or1   g0877(.dina(new_new_n2112__), .dinb(new_new_n2109__), .dout(new_new_n1501__));
  and1  g0878(.dina(new_new_n1501__), .dinb(new_new_n1500__), .dout(new_new_n1502__));
  or1   g0879(.dina(new_new_n2114__), .dinb(new_new_n2108__), .dout(new_new_n1503__));
  or1   g0880(.dina(new_new_n2115__), .dinb(new_new_n2104__), .dout(new_new_n1504__));
  and1  g0881(.dina(new_new_n1504__), .dinb(new_new_n1503__), .dout(new_new_n1505__));
  or1   g0882(.dina(new_new_n2102__), .dinb(new_new_n2099__), .dout(new_new_n1506__));
  or1   g0883(.dina(new_new_n2103__), .dinb(new_new_n2100__), .dout(new_new_n1507__));
  and1  g0884(.dina(new_new_n1507__), .dinb(new_new_n1506__), .dout(new_new_n1508__));
  and1  g0885(.dina(new_new_n2115__), .dinb(new_new_n2111__), .dout(new_new_n1509__));
  and1  g0886(.dina(new_new_n2114__), .dinb(new_new_n2112__), .dout(new_new_n1510__));
  or1   g0887(.dina(new_new_n1510__), .dinb(new_new_n1509__), .dout(new_new_n1511__));
  or1   g0888(.dina(new_new_n2117__), .dinb(new_new_n2119__), .dout(new_new_n1512__));
  or1   g0889(.dina(new_new_n2120__), .dinb(new_new_n2121__), .dout(new_new_n1513__));
  and1  g0890(.dina(new_new_n1513__), .dinb(new_new_n1512__), .dout(new_new_n1514__));
  and1  g0891(.dina(new_new_n2122__), .dinb(new_new_n2119__), .dout(new_new_n1515__));
  and1  g0892(.dina(new_new_n2124__), .dinb(new_new_n2121__), .dout(new_new_n1516__));
  or1   g0893(.dina(new_new_n1516__), .dinb(new_new_n1515__), .dout(new_new_n1517__));
  and1  g0894(.dina(new_new_n2125__), .dinb(new_new_n2117__), .dout(new_new_n1518__));
  and1  g0895(.dina(new_new_n2127__), .dinb(new_new_n2120__), .dout(new_new_n1519__));
  or1   g0896(.dina(new_new_n1519__), .dinb(new_new_n1518__), .dout(new_new_n1520__));
  and1  g0897(.dina(new_new_n2128__), .dinb(new_new_n2130__), .dout(new_new_n1521__));
  and1  g0898(.dina(new_new_n2132__), .dinb(new_new_n2133__), .dout(new_new_n1522__));
  or1   g0899(.dina(new_new_n1522__), .dinb(new_new_n1521__), .dout(new_new_n1523__));
  and1  g0900(.dina(new_new_n2134__), .dinb(new_new_n2130__), .dout(new_new_n1524__));
  and1  g0901(.dina(new_new_n2136__), .dinb(new_new_n2133__), .dout(new_new_n1525__));
  or1   g0902(.dina(new_new_n1525__), .dinb(new_new_n1524__), .dout(new_new_n1526__));
  and1  g0903(.dina(new_new_n2137__), .dinb(new_new_n2132__), .dout(new_new_n1527__));
  and1  g0904(.dina(new_new_n2139__), .dinb(new_new_n2128__), .dout(new_new_n1528__));
  or1   g0905(.dina(new_new_n1528__), .dinb(new_new_n1527__), .dout(new_new_n1529__));
  or1   g0906(.dina(new_new_n2127__), .dinb(new_new_n2124__), .dout(new_new_n1530__));
  or1   g0907(.dina(new_new_n2125__), .dinb(new_new_n2122__), .dout(new_new_n1531__));
  and1  g0908(.dina(new_new_n1531__), .dinb(new_new_n1530__), .dout(new_new_n1532__));
  and1  g0909(.dina(new_new_n2137__), .dinb(new_new_n2136__), .dout(new_new_n1533__));
  and1  g0910(.dina(new_new_n2139__), .dinb(new_new_n2134__), .dout(new_new_n1534__));
  or1   g0911(.dina(new_new_n1534__), .dinb(new_new_n1533__), .dout(new_new_n1535__));
  buf1  g0912(.din(new_new_n1038__), .dout(G1324));
  buf1  g0913(.din(new_new_n1043__), .dout(G1325));
  buf1  g0914(.din(new_new_n1048__), .dout(G1326));
  buf1  g0915(.din(new_new_n1053__), .dout(G1327));
  buf1  g0916(.din(new_new_n1062__), .dout(G1328));
  buf1  g0917(.din(new_new_n1067__), .dout(G1329));
  buf1  g0918(.din(new_new_n1072__), .dout(G1330));
  buf1  g0919(.din(new_new_n1077__), .dout(G1331));
  buf1  g0920(.din(new_new_n1086__), .dout(G1332));
  buf1  g0921(.din(new_new_n1091__), .dout(G1333));
  buf1  g0922(.din(new_new_n1096__), .dout(G1334));
  buf1  g0923(.din(new_new_n1101__), .dout(G1335));
  buf1  g0924(.din(new_new_n1110__), .dout(G1336));
  buf1  g0925(.din(new_new_n1115__), .dout(G1337));
  buf1  g0926(.din(new_new_n1120__), .dout(G1338));
  buf1  g0927(.din(new_new_n1125__), .dout(G1339));
  buf1  g0928(.din(new_new_n1134__), .dout(G1340));
  buf1  g0929(.din(new_new_n1139__), .dout(G1341));
  buf1  g0930(.din(new_new_n1144__), .dout(G1342));
  buf1  g0931(.din(new_new_n1149__), .dout(G1343));
  buf1  g0932(.din(new_new_n1158__), .dout(G1344));
  buf1  g0933(.din(new_new_n1163__), .dout(G1345));
  buf1  g0934(.din(new_new_n1168__), .dout(G1346));
  buf1  g0935(.din(new_new_n1173__), .dout(G1347));
  buf1  g0936(.din(new_new_n1182__), .dout(G1348));
  buf1  g0937(.din(new_new_n1187__), .dout(G1349));
  buf1  g0938(.din(new_new_n1192__), .dout(G1350));
  buf1  g0939(.din(new_new_n1197__), .dout(G1351));
  buf1  g0940(.din(new_new_n1206__), .dout(G1352));
  buf1  g0941(.din(new_new_n1211__), .dout(G1353));
  buf1  g0942(.din(new_new_n1216__), .dout(G1354));
  buf1  g0943(.din(new_new_n1221__), .dout(G1355));
  buf1  g0944(.din(new_new_n510__), .dout(n3365));
  buf1  g0945(.din(new_new_n754__), .dout(n3368));
  buf1  g0946(.din(new_new_n512__), .dout(n3371));
  buf1  g0947(.din(new_new_n756__), .dout(n3374));
  buf1  g0948(.din(new_new_n514__), .dout(n3377));
  buf1  g0949(.din(new_new_n758__), .dout(n3380));
  buf1  g0950(.din(new_new_n516__), .dout(n3383));
  buf1  g0951(.din(new_new_n760__), .dout(n3386));
  buf1  g0952(.din(new_new_n518__), .dout(n3389));
  buf1  g0953(.din(new_new_n762__), .dout(n3392));
  buf1  g0954(.din(new_new_n520__), .dout(n3395));
  buf1  g0955(.din(new_new_n764__), .dout(n3398));
  buf1  g0956(.din(new_new_n522__), .dout(n3401));
  buf1  g0957(.din(new_new_n766__), .dout(n3404));
  buf1  g0958(.din(new_new_n524__), .dout(n3407));
  buf1  g0959(.din(new_new_n768__), .dout(n3410));
  buf1  g0960(.din(new_new_n526__), .dout(n3413));
  buf1  g0961(.din(new_new_n770__), .dout(n3416));
  buf1  g0962(.din(new_new_n528__), .dout(n3419));
  buf1  g0963(.din(new_new_n772__), .dout(n3422));
  buf1  g0964(.din(new_new_n530__), .dout(n3425));
  buf1  g0965(.din(new_new_n774__), .dout(n3428));
  buf1  g0966(.din(new_new_n532__), .dout(n3431));
  buf1  g0967(.din(new_new_n776__), .dout(n3434));
  buf1  g0968(.din(new_new_n534__), .dout(n3437));
  buf1  g0969(.din(new_new_n778__), .dout(n3440));
  buf1  g0970(.din(new_new_n536__), .dout(n3443));
  buf1  g0971(.din(new_new_n780__), .dout(n3446));
  buf1  g0972(.din(new_new_n538__), .dout(n3449));
  buf1  g0973(.din(new_new_n782__), .dout(n3452));
  buf1  g0974(.din(new_new_n540__), .dout(n3455));
  buf1  g0975(.din(new_new_n784__), .dout(n3458));
  buf1  g0976(.din(new_new_n542__), .dout(n3461));
  buf1  g0977(.din(new_new_n786__), .dout(n3464));
  buf1  g0978(.din(new_new_n544__), .dout(n3467));
  buf1  g0979(.din(new_new_n788__), .dout(n3470));
  buf1  g0980(.din(new_new_n546__), .dout(n3473));
  buf1  g0981(.din(new_new_n790__), .dout(n3476));
  buf1  g0982(.din(new_new_n548__), .dout(n3479));
  buf1  g0983(.din(new_new_n792__), .dout(n3482));
  buf1  g0984(.din(new_new_n550__), .dout(n3485));
  buf1  g0985(.din(new_new_n794__), .dout(n3488));
  buf1  g0986(.din(new_new_n552__), .dout(n3491));
  buf1  g0987(.din(new_new_n796__), .dout(n3494));
  buf1  g0988(.din(new_new_n554__), .dout(n3497));
  buf1  g0989(.din(new_new_n798__), .dout(n3500));
  buf1  g0990(.din(new_new_n556__), .dout(n3503));
  buf1  g0991(.din(new_new_n800__), .dout(n3506));
  buf1  g0992(.din(new_new_n558__), .dout(n3509));
  buf1  g0993(.din(new_new_n802__), .dout(n3512));
  buf1  g0994(.din(new_new_n560__), .dout(n3515));
  buf1  g0995(.din(new_new_n804__), .dout(n3518));
  buf1  g0996(.din(new_new_n562__), .dout(n3521));
  buf1  g0997(.din(new_new_n806__), .dout(n3524));
  buf1  g0998(.din(new_new_n564__), .dout(n3527));
  buf1  g0999(.din(new_new_n808__), .dout(n3530));
  buf1  g1000(.din(new_new_n566__), .dout(n3533));
  buf1  g1001(.din(new_new_n810__), .dout(n3536));
  buf1  g1002(.din(new_new_n568__), .dout(n3539));
  buf1  g1003(.din(new_new_n812__), .dout(n3542));
  buf1  g1004(.din(new_new_n570__), .dout(n3545));
  buf1  g1005(.din(new_new_n814__), .dout(n3548));
  buf1  g1006(.din(new_new_n572__), .dout(n3551));
  buf1  g1007(.din(new_new_n816__), .dout(n3554));
  buf1  g1008(.din(new_new_n574__), .dout(n3557));
  buf1  g1009(.din(new_new_n576__), .dout(n3560));
  buf1  g1010(.din(new_new_n578__), .dout(n3563));
  buf1  g1011(.din(new_new_n580__), .dout(n3566));
  buf1  g1012(.din(new_new_n582__), .dout(n3569));
  buf1  g1013(.din(new_new_n584__), .dout(n3572));
  buf1  g1014(.din(new_new_n586__), .dout(n3575));
  buf1  g1015(.din(new_new_n588__), .dout(n3578));
  buf1  g1016(.din(new_new_n590__), .dout(n3581));
  buf1  g1017(.din(new_new_n1917__), .dout(n3584));
  buf1  g1018(.din(new_new_n1900__), .dout(n3587));
  buf1  g1019(.din(new_new_n1902__), .dout(n3590));
  buf1  g1020(.din(new_new_n1919__), .dout(n3593));
  buf1  g1021(.din(new_new_n1910__), .dout(n3596));
  buf1  g1022(.din(new_new_n1925__), .dout(n3599));
  buf1  g1023(.din(new_new_n1923__), .dout(n3602));
  buf1  g1024(.din(new_new_n1908__), .dout(n3605));
  buf1  g1025(.din(new_new_n850__), .dout(n3608));
  buf1  g1026(.din(new_new_n852__), .dout(n3611));
  buf1  g1027(.din(new_new_n854__), .dout(n3614));
  buf1  g1028(.din(new_new_n856__), .dout(n3617));
  buf1  g1029(.din(new_new_n858__), .dout(n3620));
  buf1  g1030(.din(new_new_n860__), .dout(n3623));
  buf1  g1031(.din(new_new_n862__), .dout(n3626));
  buf1  g1032(.din(new_new_n864__), .dout(n3629));
  buf1  g1033(.din(new_new_n866__), .dout(n3632));
  buf1  g1034(.din(new_new_n868__), .dout(n3635));
  buf1  g1035(.din(new_new_n870__), .dout(n3638));
  buf1  g1036(.din(new_new_n872__), .dout(n3641));
  buf1  g1037(.din(new_new_n874__), .dout(n3644));
  buf1  g1038(.din(new_new_n876__), .dout(n3647));
  buf1  g1039(.din(new_new_n878__), .dout(n3650));
  buf1  g1040(.din(new_new_n880__), .dout(n3653));
  buf1  g1041(.din(new_new_n882__), .dout(n3656));
  buf1  g1042(.din(new_new_n884__), .dout(n3659));
  buf1  g1043(.din(new_new_n886__), .dout(n3662));
  buf1  g1044(.din(new_new_n888__), .dout(n3665));
  buf1  g1045(.din(new_new_n890__), .dout(n3668));
  buf1  g1046(.din(new_new_n892__), .dout(n3671));
  buf1  g1047(.din(new_new_n894__), .dout(n3674));
  buf1  g1048(.din(new_new_n896__), .dout(n3677));
  buf1  g1049(.din(new_new_n898__), .dout(n3680));
  buf1  g1050(.din(new_new_n900__), .dout(n3683));
  buf1  g1051(.din(new_new_n902__), .dout(n3686));
  buf1  g1052(.din(new_new_n904__), .dout(n3689));
  buf1  g1053(.din(new_new_n906__), .dout(n3692));
  buf1  g1054(.din(new_new_n908__), .dout(n3695));
  buf1  g1055(.din(new_new_n910__), .dout(n3698));
  buf1  g1056(.din(new_new_n912__), .dout(n3701));
  not1  g1057(.din(new_new_n1922__), .dout(n3704));
  not1  g1058(.din(new_new_n1916__), .dout(n3707));
  not1  g1059(.din(new_new_n1931__), .dout(n3710));
  buf1  g1060(.din(new_new_n1930__), .dout(n3713));
  not1  g1061(.din(new_new_n1933__), .dout(n3716));
  not1  g1062(.din(new_new_n1927__), .dout(n3719));
  not1  g1063(.din(new_new_n1929__), .dout(n3722));
  not1  g1064(.din(new_new_n1928__), .dout(n3725));
  buf1  g1065(.din(new_new_n1932__), .dout(n3728));
  not1  g1066(.din(new_new_n1252__), .dout(n3731));
  not1  g1067(.din(new_new_n1254__), .dout(n3734));
  buf1  g1068(.din(new_new_n1255__), .dout(n3737));
  buf1  g1069(.din(new_new_n1256__), .dout(n3740));
  buf1  g1070(.din(new_new_n1257__), .dout(n3743));
  buf1  g1071(.din(new_new_n1258__), .dout(n3746));
  buf1  g1072(.din(new_new_n1263__), .dout(n3749));
  buf1  g1073(.din(new_new_n2046__), .dout(n3752));
  buf1  g1074(.din(new_new_n2050__), .dout(n3755));
  buf1  g1075(.din(new_new_n2058__), .dout(n3758));
  buf1  g1076(.din(new_new_n2063__), .dout(n3761));
  buf1  g1077(.din(new_new_n2044__), .dout(n3764));
  buf1  g1078(.din(new_new_n2053__), .dout(n3767));
  buf1  g1079(.din(new_new_n2056__), .dout(n3770));
  buf1  g1080(.din(new_new_n2065__), .dout(n3773));
  buf1  g1081(.din(new_new_n2069__), .dout(n3776));
  buf1  g1082(.din(new_new_n2074__), .dout(n3779));
  buf1  g1083(.din(new_new_n2081__), .dout(n3782));
  buf1  g1084(.din(new_new_n2087__), .dout(n3785));
  buf1  g1085(.din(new_new_n2071__), .dout(n3788));
  buf1  g1086(.din(new_new_n2078__), .dout(n3791));
  buf1  g1087(.din(new_new_n2083__), .dout(n3794));
  buf1  g1088(.din(new_new_n2090__), .dout(n3797));
  buf1  g1089(.din(new_new_n2094__), .dout(n3800));
  buf1  g1090(.din(new_new_n2092__), .dout(n3803));
  buf1  g1091(.din(new_new_n2105__), .dout(n3806));
  buf1  g1092(.din(new_new_n2107__), .dout(n3809));
  buf1  g1093(.din(new_new_n2098__), .dout(n3812));
  buf1  g1094(.din(new_new_n2101__), .dout(n3815));
  buf1  g1095(.din(new_new_n2110__), .dout(n3818));
  buf1  g1096(.din(new_new_n2113__), .dout(n3821));
  buf1  g1097(.din(new_new_n2118__), .dout(n3824));
  buf1  g1098(.din(new_new_n2116__), .dout(n3827));
  buf1  g1099(.din(new_new_n2129__), .dout(n3830));
  buf1  g1100(.din(new_new_n2131__), .dout(n3833));
  buf1  g1101(.din(new_new_n2123__), .dout(n3836));
  buf1  g1102(.din(new_new_n2126__), .dout(n3839));
  buf1  g1103(.din(new_new_n2135__), .dout(n3842));
  buf1  g1104(.din(new_new_n2138__), .dout(n3845));
  buf1  g1105(.din(new_new_n1290__), .dout(n3848));
  not1  g1106(.din(new_new_n1291__), .dout(n3851));
  buf1  g1107(.din(new_new_n1318__), .dout(n3854));
  not1  g1108(.din(new_new_n1319__), .dout(n3857));
  buf1  g1109(.din(new_new_n1334__), .dout(n3860));
  not1  g1110(.din(new_new_n1335__), .dout(n3863));
  buf1  g1111(.din(new_new_n1350__), .dout(n3866));
  not1  g1112(.din(new_new_n1351__), .dout(n3869));
  buf1  g1113(.din(new_new_n1378__), .dout(n3872));
  not1  g1114(.din(new_new_n1379__), .dout(n3875));
  buf1  g1115(.din(new_new_n1406__), .dout(n3878));
  not1  g1116(.din(new_new_n1407__), .dout(n3881));
  buf1  g1117(.din(new_new_n1422__), .dout(n3884));
  not1  g1118(.din(new_new_n1423__), .dout(n3887));
  buf1  g1119(.din(new_new_n1438__), .dout(n3890));
  not1  g1120(.din(new_new_n1439__), .dout(n3893));
  buf1  g1121(.din(new_new_n720__), .dout(n3896));
  buf1  g1122(.din(new_new_n722__), .dout(n3899));
  buf1  g1123(.din(new_new_n724__), .dout(n3902));
  buf1  g1124(.din(new_new_n726__), .dout(n3905));
  buf1  g1125(.din(new_new_n728__), .dout(n3908));
  buf1  g1126(.din(new_new_n730__), .dout(n3911));
  buf1  g1127(.din(new_new_n732__), .dout(n3914));
  buf1  g1128(.din(new_new_n734__), .dout(n3917));
  buf1  g1129(.din(new_new_n736__), .dout(n3920));
  buf1  g1130(.din(new_new_n1442__), .dout(n3923));
  buf1  g1131(.din(new_new_n1445__), .dout(n3926));
  buf1  g1132(.din(new_new_n1448__), .dout(n3929));
  buf1  g1133(.din(new_new_n1451__), .dout(n3932));
  buf1  g1134(.din(new_new_n1454__), .dout(n3935));
  buf1  g1135(.din(new_new_n1457__), .dout(n3938));
  buf1  g1136(.din(new_new_n1460__), .dout(n3941));
  buf1  g1137(.din(new_new_n1463__), .dout(n3944));
  buf1  g1138(.din(new_new_n1466__), .dout(n3947));
  buf1  g1139(.din(new_new_n1469__), .dout(n3950));
  buf1  g1140(.din(new_new_n1472__), .dout(n3953));
  buf1  g1141(.din(new_new_n1475__), .dout(n3956));
  buf1  g1142(.din(new_new_n1478__), .dout(n3959));
  buf1  g1143(.din(new_new_n1481__), .dout(n3962));
  buf1  g1144(.din(new_new_n1484__), .dout(n3965));
  buf1  g1145(.din(new_new_n1487__), .dout(n3968));
  buf1  g1146(.din(new_new_n1490__), .dout(n3971));
  buf1  g1147(.din(new_new_n1493__), .dout(n3974));
  buf1  g1148(.din(new_new_n1496__), .dout(n3977));
  buf1  g1149(.din(new_new_n1499__), .dout(n3980));
  buf1  g1150(.din(new_new_n1502__), .dout(n3983));
  buf1  g1151(.din(new_new_n1505__), .dout(n3986));
  buf1  g1152(.din(new_new_n1508__), .dout(n3989));
  buf1  g1153(.din(new_new_n1511__), .dout(n3992));
  buf1  g1154(.din(new_new_n1514__), .dout(n3995));
  buf1  g1155(.din(new_new_n1517__), .dout(n3998));
  buf1  g1156(.din(new_new_n1520__), .dout(n4001));
  buf1  g1157(.din(new_new_n1523__), .dout(n4004));
  buf1  g1158(.din(new_new_n1526__), .dout(n4007));
  buf1  g1159(.din(new_new_n1529__), .dout(n4010));
  buf1  g1160(.din(new_new_n1532__), .dout(n4013));
  buf1  g1161(.din(new_new_n1535__), .dout(n4016));
  buf1  g1162(.din(new_new_n1029__), .dout(new_new_n1786__));
  buf1  g1163(.din(new_new_n1786__), .dout(new_new_n1787__));
  buf1  g1164(.din(new_new_n1786__), .dout(new_new_n1788__));
  buf1  g1165(.din(new_new_n1028__), .dout(new_new_n1789__));
  buf1  g1166(.din(new_new_n1789__), .dout(new_new_n1790__));
  buf1  g1167(.din(new_new_n1789__), .dout(new_new_n1791__));
  buf1  g1168(.din(new_new_n1032__), .dout(new_new_n1792__));
  buf1  g1169(.din(new_new_n1792__), .dout(new_new_n1793__));
  buf1  g1170(.din(new_new_n1792__), .dout(new_new_n1794__));
  buf1  g1171(.din(new_new_n738__), .dout(new_new_n1795__));
  buf1  g1172(.din(new_new_n1795__), .dout(new_new_n1796__));
  buf1  g1173(.din(new_new_n1795__), .dout(new_new_n1797__));
  buf1  g1174(.din(new_new_n1033__), .dout(new_new_n1798__));
  buf1  g1175(.din(new_new_n1798__), .dout(new_new_n1799__));
  buf1  g1176(.din(new_new_n1798__), .dout(new_new_n1800__));
  buf1  g1177(.din(new_new_n739__), .dout(new_new_n1801__));
  buf1  g1178(.din(new_new_n1801__), .dout(new_new_n1802__));
  buf1  g1179(.din(new_new_n1801__), .dout(new_new_n1803__));
  buf1  g1180(.din(new_new_n740__), .dout(new_new_n1804__));
  buf1  g1181(.din(new_new_n1804__), .dout(new_new_n1805__));
  buf1  g1182(.din(new_new_n1805__), .dout(new_new_n1806__));
  buf1  g1183(.din(new_new_n1804__), .dout(new_new_n1807__));
  buf1  g1184(.din(new_new_n741__), .dout(new_new_n1808__));
  buf1  g1185(.din(new_new_n1808__), .dout(new_new_n1809__));
  buf1  g1186(.din(new_new_n1809__), .dout(new_new_n1810__));
  buf1  g1187(.din(new_new_n1808__), .dout(new_new_n1811__));
  buf1  g1188(.din(new_new_n742__), .dout(new_new_n1812__));
  buf1  g1189(.din(new_new_n1812__), .dout(new_new_n1813__));
  buf1  g1190(.din(new_new_n1813__), .dout(new_new_n1814__));
  buf1  g1191(.din(new_new_n1813__), .dout(new_new_n1815__));
  buf1  g1192(.din(new_new_n1812__), .dout(new_new_n1816__));
  buf1  g1193(.din(new_new_n743__), .dout(new_new_n1817__));
  buf1  g1194(.din(new_new_n1817__), .dout(new_new_n1818__));
  buf1  g1195(.din(new_new_n1818__), .dout(new_new_n1819__));
  buf1  g1196(.din(new_new_n1818__), .dout(new_new_n1820__));
  buf1  g1197(.din(new_new_n1817__), .dout(new_new_n1821__));
  buf1  g1198(.din(new_new_n744__), .dout(new_new_n1822__));
  buf1  g1199(.din(new_new_n1822__), .dout(new_new_n1823__));
  buf1  g1200(.din(new_new_n1822__), .dout(new_new_n1824__));
  buf1  g1201(.din(new_new_n745__), .dout(new_new_n1825__));
  buf1  g1202(.din(new_new_n1825__), .dout(new_new_n1826__));
  buf1  g1203(.din(new_new_n1825__), .dout(new_new_n1827__));
  buf1  g1204(.din(new_new_n1056__), .dout(new_new_n1828__));
  buf1  g1205(.din(new_new_n1828__), .dout(new_new_n1829__));
  buf1  g1206(.din(new_new_n1828__), .dout(new_new_n1830__));
  buf1  g1207(.din(new_new_n1057__), .dout(new_new_n1831__));
  buf1  g1208(.din(new_new_n1831__), .dout(new_new_n1832__));
  buf1  g1209(.din(new_new_n1831__), .dout(new_new_n1833__));
  buf1  g1210(.din(new_new_n1080__), .dout(new_new_n1834__));
  buf1  g1211(.din(new_new_n1834__), .dout(new_new_n1835__));
  buf1  g1212(.din(new_new_n1834__), .dout(new_new_n1836__));
  buf1  g1213(.din(new_new_n1081__), .dout(new_new_n1837__));
  buf1  g1214(.din(new_new_n1837__), .dout(new_new_n1838__));
  buf1  g1215(.din(new_new_n1837__), .dout(new_new_n1839__));
  buf1  g1216(.din(new_new_n1104__), .dout(new_new_n1840__));
  buf1  g1217(.din(new_new_n1840__), .dout(new_new_n1841__));
  buf1  g1218(.din(new_new_n1840__), .dout(new_new_n1842__));
  buf1  g1219(.din(new_new_n1105__), .dout(new_new_n1843__));
  buf1  g1220(.din(new_new_n1843__), .dout(new_new_n1844__));
  buf1  g1221(.din(new_new_n1843__), .dout(new_new_n1845__));
  buf1  g1222(.din(new_new_n848__), .dout(new_new_n1846__));
  buf1  g1223(.din(new_new_n1846__), .dout(new_new_n1847__));
  buf1  g1224(.din(new_new_n1846__), .dout(new_new_n1848__));
  buf1  g1225(.din(new_new_n849__), .dout(new_new_n1849__));
  buf1  g1226(.din(new_new_n1849__), .dout(new_new_n1850__));
  buf1  g1227(.din(new_new_n1849__), .dout(new_new_n1851__));
  buf1  g1228(.din(new_new_n1128__), .dout(new_new_n1852__));
  buf1  g1229(.din(new_new_n1852__), .dout(new_new_n1853__));
  buf1  g1230(.din(new_new_n1852__), .dout(new_new_n1854__));
  buf1  g1231(.din(new_new_n746__), .dout(new_new_n1855__));
  buf1  g1232(.din(new_new_n1855__), .dout(new_new_n1856__));
  buf1  g1233(.din(new_new_n1855__), .dout(new_new_n1857__));
  buf1  g1234(.din(new_new_n1129__), .dout(new_new_n1858__));
  buf1  g1235(.din(new_new_n1858__), .dout(new_new_n1859__));
  buf1  g1236(.din(new_new_n1858__), .dout(new_new_n1860__));
  buf1  g1237(.din(new_new_n747__), .dout(new_new_n1861__));
  buf1  g1238(.din(new_new_n1861__), .dout(new_new_n1862__));
  buf1  g1239(.din(new_new_n1861__), .dout(new_new_n1863__));
  buf1  g1240(.din(new_new_n748__), .dout(new_new_n1864__));
  buf1  g1241(.din(new_new_n1864__), .dout(new_new_n1865__));
  buf1  g1242(.din(new_new_n1864__), .dout(new_new_n1866__));
  buf1  g1243(.din(new_new_n749__), .dout(new_new_n1867__));
  buf1  g1244(.din(new_new_n1867__), .dout(new_new_n1868__));
  buf1  g1245(.din(new_new_n1867__), .dout(new_new_n1869__));
  buf1  g1246(.din(new_new_n750__), .dout(new_new_n1870__));
  buf1  g1247(.din(new_new_n1870__), .dout(new_new_n1871__));
  buf1  g1248(.din(new_new_n1870__), .dout(new_new_n1872__));
  buf1  g1249(.din(new_new_n751__), .dout(new_new_n1873__));
  buf1  g1250(.din(new_new_n1873__), .dout(new_new_n1874__));
  buf1  g1251(.din(new_new_n1873__), .dout(new_new_n1875__));
  buf1  g1252(.din(new_new_n752__), .dout(new_new_n1876__));
  buf1  g1253(.din(new_new_n1876__), .dout(new_new_n1877__));
  buf1  g1254(.din(new_new_n1876__), .dout(new_new_n1878__));
  buf1  g1255(.din(new_new_n753__), .dout(new_new_n1879__));
  buf1  g1256(.din(new_new_n1879__), .dout(new_new_n1880__));
  buf1  g1257(.din(new_new_n1879__), .dout(new_new_n1881__));
  buf1  g1258(.din(new_new_n1152__), .dout(new_new_n1882__));
  buf1  g1259(.din(new_new_n1882__), .dout(new_new_n1883__));
  buf1  g1260(.din(new_new_n1882__), .dout(new_new_n1884__));
  buf1  g1261(.din(new_new_n1153__), .dout(new_new_n1885__));
  buf1  g1262(.din(new_new_n1885__), .dout(new_new_n1886__));
  buf1  g1263(.din(new_new_n1885__), .dout(new_new_n1887__));
  buf1  g1264(.din(new_new_n1176__), .dout(new_new_n1888__));
  buf1  g1265(.din(new_new_n1888__), .dout(new_new_n1889__));
  buf1  g1266(.din(new_new_n1888__), .dout(new_new_n1890__));
  buf1  g1267(.din(new_new_n1177__), .dout(new_new_n1891__));
  buf1  g1268(.din(new_new_n1891__), .dout(new_new_n1892__));
  buf1  g1269(.din(new_new_n1891__), .dout(new_new_n1893__));
  buf1  g1270(.din(new_new_n1200__), .dout(new_new_n1894__));
  buf1  g1271(.din(new_new_n1894__), .dout(new_new_n1895__));
  buf1  g1272(.din(new_new_n1894__), .dout(new_new_n1896__));
  buf1  g1273(.din(new_new_n1201__), .dout(new_new_n1897__));
  buf1  g1274(.din(new_new_n1897__), .dout(new_new_n1898__));
  buf1  g1275(.din(new_new_n1897__), .dout(new_new_n1899__));
  buf1  g1276(.din(new_new_n1225__), .dout(new_new_n1900__));
  buf1  g1277(.din(new_new_n1900__), .dout(new_new_n1901__));
  buf1  g1278(.din(new_new_n1227__), .dout(new_new_n1902__));
  buf1  g1279(.din(new_new_n1902__), .dout(new_new_n1903__));
  buf1  g1280(.din(new_new_n1236__), .dout(new_new_n1904__));
  buf1  g1281(.din(new_new_n1904__), .dout(new_new_n1905__));
  buf1  g1282(.din(new_new_n1230__), .dout(new_new_n1906__));
  buf1  g1283(.din(new_new_n1906__), .dout(new_new_n1907__));
  buf1  g1284(.din(new_new_n1237__), .dout(new_new_n1908__));
  buf1  g1285(.din(new_new_n1908__), .dout(new_new_n1909__));
  buf1  g1286(.din(new_new_n1231__), .dout(new_new_n1910__));
  buf1  g1287(.din(new_new_n1910__), .dout(new_new_n1911__));
  buf1  g1288(.din(new_new_n1234__), .dout(new_new_n1912__));
  buf1  g1289(.din(new_new_n1912__), .dout(new_new_n1913__));
  buf1  g1290(.din(new_new_n1232__), .dout(new_new_n1914__));
  buf1  g1291(.din(new_new_n1914__), .dout(new_new_n1915__));
  buf1  g1292(.din(new_new_n1239__), .dout(new_new_n1916__));
  buf1  g1293(.din(new_new_n1223__), .dout(new_new_n1917__));
  buf1  g1294(.din(new_new_n1917__), .dout(new_new_n1918__));
  buf1  g1295(.din(new_new_n1229__), .dout(new_new_n1919__));
  buf1  g1296(.din(new_new_n1919__), .dout(new_new_n1920__));
  buf1  g1297(.din(new_new_n1245__), .dout(new_new_n1921__));
  buf1  g1298(.din(new_new_n1238__), .dout(new_new_n1922__));
  buf1  g1299(.din(new_new_n1235__), .dout(new_new_n1923__));
  buf1  g1300(.din(new_new_n1923__), .dout(new_new_n1924__));
  buf1  g1301(.din(new_new_n1233__), .dout(new_new_n1925__));
  buf1  g1302(.din(new_new_n1925__), .dout(new_new_n1926__));
  buf1  g1303(.din(new_new_n1244__), .dout(new_new_n1927__));
  buf1  g1304(.din(new_new_n1247__), .dout(new_new_n1928__));
  buf1  g1305(.din(new_new_n1246__), .dout(new_new_n1929__));
  buf1  g1306(.din(new_new_n1242__), .dout(new_new_n1930__));
  buf1  g1307(.din(new_new_n1240__), .dout(new_new_n1931__));
  buf1  g1308(.din(new_new_n1249__), .dout(new_new_n1932__));
  buf1  g1309(.din(new_new_n1243__), .dout(new_new_n1933__));
  buf1  g1310(.din(new_new_n981__), .dout(new_new_n1934__));
  buf1  g1311(.din(new_new_n964__), .dout(new_new_n1935__));
  buf1  g1312(.din(new_new_n980__), .dout(new_new_n1936__));
  buf1  g1313(.din(new_new_n965__), .dout(new_new_n1937__));
  buf1  g1314(.din(new_new_n962__), .dout(new_new_n1938__));
  buf1  g1315(.din(new_new_n1938__), .dout(new_new_n1939__));
  buf1  g1316(.din(new_new_n1939__), .dout(new_new_n1940__));
  buf1  g1317(.din(new_new_n1939__), .dout(new_new_n1941__));
  buf1  g1318(.din(new_new_n1938__), .dout(new_new_n1942__));
  buf1  g1319(.din(new_new_n1942__), .dout(new_new_n1943__));
  buf1  g1320(.din(new_new_n1942__), .dout(new_new_n1944__));
  buf1  g1321(.din(new_new_n963__), .dout(new_new_n1945__));
  buf1  g1322(.din(new_new_n1945__), .dout(new_new_n1946__));
  buf1  g1323(.din(new_new_n1946__), .dout(new_new_n1947__));
  buf1  g1324(.din(new_new_n1946__), .dout(new_new_n1948__));
  buf1  g1325(.din(new_new_n1945__), .dout(new_new_n1949__));
  buf1  g1326(.din(new_new_n1949__), .dout(new_new_n1950__));
  buf1  g1327(.din(new_new_n1949__), .dout(new_new_n1951__));
  buf1  g1328(.din(new_new_n1003__), .dout(new_new_n1952__));
  buf1  g1329(.din(new_new_n996__), .dout(new_new_n1953__));
  buf1  g1330(.din(new_new_n1002__), .dout(new_new_n1954__));
  buf1  g1331(.din(new_new_n997__), .dout(new_new_n1955__));
  buf1  g1332(.din(new_new_n1011__), .dout(new_new_n1956__));
  buf1  g1333(.din(new_new_n1008__), .dout(new_new_n1957__));
  buf1  g1334(.din(new_new_n1010__), .dout(new_new_n1958__));
  buf1  g1335(.din(new_new_n1009__), .dout(new_new_n1959__));
  buf1  g1336(.din(new_new_n1286__), .dout(new_new_n1960__));
  buf1  g1337(.din(new_new_n1279__), .dout(new_new_n1961__));
  buf1  g1338(.din(new_new_n1285__), .dout(new_new_n1962__));
  buf1  g1339(.din(new_new_n1280__), .dout(new_new_n1963__));
  buf1  g1340(.din(new_new_n1289__), .dout(new_new_n1964__));
  buf1  g1341(.din(new_new_n1274__), .dout(new_new_n1965__));
  buf1  g1342(.din(new_new_n985__), .dout(new_new_n1966__));
  buf1  g1343(.din(new_new_n968__), .dout(new_new_n1967__));
  buf1  g1344(.din(new_new_n984__), .dout(new_new_n1968__));
  buf1  g1345(.din(new_new_n969__), .dout(new_new_n1969__));
  buf1  g1346(.din(new_new_n1027__), .dout(new_new_n1970__));
  buf1  g1347(.din(new_new_n1024__), .dout(new_new_n1971__));
  buf1  g1348(.din(new_new_n1026__), .dout(new_new_n1972__));
  buf1  g1349(.din(new_new_n1025__), .dout(new_new_n1973__));
  buf1  g1350(.din(new_new_n1019__), .dout(new_new_n1974__));
  buf1  g1351(.din(new_new_n1012__), .dout(new_new_n1975__));
  buf1  g1352(.din(new_new_n1018__), .dout(new_new_n1976__));
  buf1  g1353(.din(new_new_n1013__), .dout(new_new_n1977__));
  buf1  g1354(.din(new_new_n1314__), .dout(new_new_n1978__));
  buf1  g1355(.din(new_new_n1307__), .dout(new_new_n1979__));
  buf1  g1356(.din(new_new_n1313__), .dout(new_new_n1980__));
  buf1  g1357(.din(new_new_n1308__), .dout(new_new_n1981__));
  buf1  g1358(.din(new_new_n1317__), .dout(new_new_n1982__));
  buf1  g1359(.din(new_new_n1302__), .dout(new_new_n1983__));
  buf1  g1360(.din(new_new_n987__), .dout(new_new_n1984__));
  buf1  g1361(.din(new_new_n970__), .dout(new_new_n1985__));
  buf1  g1362(.din(new_new_n986__), .dout(new_new_n1986__));
  buf1  g1363(.din(new_new_n971__), .dout(new_new_n1987__));
  buf1  g1364(.din(new_new_n1333__), .dout(new_new_n1988__));
  buf1  g1365(.din(new_new_n1330__), .dout(new_new_n1989__));
  buf1  g1366(.din(new_new_n991__), .dout(new_new_n1990__));
  buf1  g1367(.din(new_new_n974__), .dout(new_new_n1991__));
  buf1  g1368(.din(new_new_n990__), .dout(new_new_n1992__));
  buf1  g1369(.din(new_new_n975__), .dout(new_new_n1993__));
  buf1  g1370(.din(new_new_n1349__), .dout(new_new_n1994__));
  buf1  g1371(.din(new_new_n1346__), .dout(new_new_n1995__));
  buf1  g1372(.din(new_new_n1015__), .dout(new_new_n1996__));
  buf1  g1373(.din(new_new_n998__), .dout(new_new_n1997__));
  buf1  g1374(.din(new_new_n1014__), .dout(new_new_n1998__));
  buf1  g1375(.din(new_new_n999__), .dout(new_new_n1999__));
  buf1  g1376(.din(new_new_n973__), .dout(new_new_n2000__));
  buf1  g1377(.din(new_new_n966__), .dout(new_new_n2001__));
  buf1  g1378(.din(new_new_n972__), .dout(new_new_n2002__));
  buf1  g1379(.din(new_new_n967__), .dout(new_new_n2003__));
  buf1  g1380(.din(new_new_n979__), .dout(new_new_n2004__));
  buf1  g1381(.din(new_new_n976__), .dout(new_new_n2005__));
  buf1  g1382(.din(new_new_n978__), .dout(new_new_n2006__));
  buf1  g1383(.din(new_new_n977__), .dout(new_new_n2007__));
  buf1  g1384(.din(new_new_n1374__), .dout(new_new_n2008__));
  buf1  g1385(.din(new_new_n1367__), .dout(new_new_n2009__));
  buf1  g1386(.din(new_new_n1373__), .dout(new_new_n2010__));
  buf1  g1387(.din(new_new_n1368__), .dout(new_new_n2011__));
  buf1  g1388(.din(new_new_n1377__), .dout(new_new_n2012__));
  buf1  g1389(.din(new_new_n1362__), .dout(new_new_n2013__));
  buf1  g1390(.din(new_new_n1017__), .dout(new_new_n2014__));
  buf1  g1391(.din(new_new_n1000__), .dout(new_new_n2015__));
  buf1  g1392(.din(new_new_n1016__), .dout(new_new_n2016__));
  buf1  g1393(.din(new_new_n1001__), .dout(new_new_n2017__));
  buf1  g1394(.din(new_new_n989__), .dout(new_new_n2018__));
  buf1  g1395(.din(new_new_n982__), .dout(new_new_n2019__));
  buf1  g1396(.din(new_new_n988__), .dout(new_new_n2020__));
  buf1  g1397(.din(new_new_n983__), .dout(new_new_n2021__));
  buf1  g1398(.din(new_new_n995__), .dout(new_new_n2022__));
  buf1  g1399(.din(new_new_n992__), .dout(new_new_n2023__));
  buf1  g1400(.din(new_new_n994__), .dout(new_new_n2024__));
  buf1  g1401(.din(new_new_n993__), .dout(new_new_n2025__));
  buf1  g1402(.din(new_new_n1402__), .dout(new_new_n2026__));
  buf1  g1403(.din(new_new_n1395__), .dout(new_new_n2027__));
  buf1  g1404(.din(new_new_n1401__), .dout(new_new_n2028__));
  buf1  g1405(.din(new_new_n1396__), .dout(new_new_n2029__));
  buf1  g1406(.din(new_new_n1405__), .dout(new_new_n2030__));
  buf1  g1407(.din(new_new_n1390__), .dout(new_new_n2031__));
  buf1  g1408(.din(new_new_n1021__), .dout(new_new_n2032__));
  buf1  g1409(.din(new_new_n1004__), .dout(new_new_n2033__));
  buf1  g1410(.din(new_new_n1020__), .dout(new_new_n2034__));
  buf1  g1411(.din(new_new_n1005__), .dout(new_new_n2035__));
  buf1  g1412(.din(new_new_n1421__), .dout(new_new_n2036__));
  buf1  g1413(.din(new_new_n1418__), .dout(new_new_n2037__));
  buf1  g1414(.din(new_new_n1023__), .dout(new_new_n2038__));
  buf1  g1415(.din(new_new_n1006__), .dout(new_new_n2039__));
  buf1  g1416(.din(new_new_n1022__), .dout(new_new_n2040__));
  buf1  g1417(.din(new_new_n1007__), .dout(new_new_n2041__));
  buf1  g1418(.din(new_new_n1437__), .dout(new_new_n2042__));
  buf1  g1419(.din(new_new_n1434__), .dout(new_new_n2043__));
  buf1  g1420(.din(new_new_n608__), .dout(new_new_n2044__));
  buf1  g1421(.din(new_new_n2044__), .dout(new_new_n2045__));
  buf1  g1422(.din(new_new_n592__), .dout(new_new_n2046__));
  buf1  g1423(.din(new_new_n2046__), .dout(new_new_n2047__));
  buf1  g1424(.din(new_new_n609__), .dout(new_new_n2048__));
  buf1  g1425(.din(new_new_n593__), .dout(new_new_n2049__));
  buf1  g1426(.din(new_new_n596__), .dout(new_new_n2050__));
  buf1  g1427(.din(new_new_n2050__), .dout(new_new_n2051__));
  buf1  g1428(.din(new_new_n597__), .dout(new_new_n2052__));
  buf1  g1429(.din(new_new_n612__), .dout(new_new_n2053__));
  buf1  g1430(.din(new_new_n2053__), .dout(new_new_n2054__));
  buf1  g1431(.din(new_new_n613__), .dout(new_new_n2055__));
  buf1  g1432(.din(new_new_n616__), .dout(new_new_n2056__));
  buf1  g1433(.din(new_new_n2056__), .dout(new_new_n2057__));
  buf1  g1434(.din(new_new_n600__), .dout(new_new_n2058__));
  buf1  g1435(.din(new_new_n2058__), .dout(new_new_n2059__));
  buf1  g1436(.din(new_new_n617__), .dout(new_new_n2060__));
  buf1  g1437(.din(new_new_n601__), .dout(new_new_n2061__));
  buf1  g1438(.din(new_new_n605__), .dout(new_new_n2062__));
  buf1  g1439(.din(new_new_n604__), .dout(new_new_n2063__));
  buf1  g1440(.din(new_new_n2063__), .dout(new_new_n2064__));
  buf1  g1441(.din(new_new_n620__), .dout(new_new_n2065__));
  buf1  g1442(.din(new_new_n2065__), .dout(new_new_n2066__));
  buf1  g1443(.din(new_new_n621__), .dout(new_new_n2067__));
  buf1  g1444(.din(new_new_n641__), .dout(new_new_n2068__));
  buf1  g1445(.din(new_new_n624__), .dout(new_new_n2069__));
  buf1  g1446(.din(new_new_n2069__), .dout(new_new_n2070__));
  buf1  g1447(.din(new_new_n640__), .dout(new_new_n2071__));
  buf1  g1448(.din(new_new_n2071__), .dout(new_new_n2072__));
  buf1  g1449(.din(new_new_n625__), .dout(new_new_n2073__));
  buf1  g1450(.din(new_new_n628__), .dout(new_new_n2074__));
  buf1  g1451(.din(new_new_n2074__), .dout(new_new_n2075__));
  buf1  g1452(.din(new_new_n629__), .dout(new_new_n2076__));
  buf1  g1453(.din(new_new_n645__), .dout(new_new_n2077__));
  buf1  g1454(.din(new_new_n644__), .dout(new_new_n2078__));
  buf1  g1455(.din(new_new_n2078__), .dout(new_new_n2079__));
  buf1  g1456(.din(new_new_n649__), .dout(new_new_n2080__));
  buf1  g1457(.din(new_new_n632__), .dout(new_new_n2081__));
  buf1  g1458(.din(new_new_n2081__), .dout(new_new_n2082__));
  buf1  g1459(.din(new_new_n648__), .dout(new_new_n2083__));
  buf1  g1460(.din(new_new_n2083__), .dout(new_new_n2084__));
  buf1  g1461(.din(new_new_n633__), .dout(new_new_n2085__));
  buf1  g1462(.din(new_new_n637__), .dout(new_new_n2086__));
  buf1  g1463(.din(new_new_n636__), .dout(new_new_n2087__));
  buf1  g1464(.din(new_new_n2087__), .dout(new_new_n2088__));
  buf1  g1465(.din(new_new_n653__), .dout(new_new_n2089__));
  buf1  g1466(.din(new_new_n652__), .dout(new_new_n2090__));
  buf1  g1467(.din(new_new_n2090__), .dout(new_new_n2091__));
  buf1  g1468(.din(new_new_n660__), .dout(new_new_n2092__));
  buf1  g1469(.din(new_new_n2092__), .dout(new_new_n2093__));
  buf1  g1470(.din(new_new_n656__), .dout(new_new_n2094__));
  buf1  g1471(.din(new_new_n2094__), .dout(new_new_n2095__));
  buf1  g1472(.din(new_new_n661__), .dout(new_new_n2096__));
  buf1  g1473(.din(new_new_n657__), .dout(new_new_n2097__));
  buf1  g1474(.din(new_new_n672__), .dout(new_new_n2098__));
  buf1  g1475(.din(new_new_n2098__), .dout(new_new_n2099__));
  buf1  g1476(.din(new_new_n673__), .dout(new_new_n2100__));
  buf1  g1477(.din(new_new_n676__), .dout(new_new_n2101__));
  buf1  g1478(.din(new_new_n2101__), .dout(new_new_n2102__));
  buf1  g1479(.din(new_new_n677__), .dout(new_new_n2103__));
  buf1  g1480(.din(new_new_n669__), .dout(new_new_n2104__));
  buf1  g1481(.din(new_new_n664__), .dout(new_new_n2105__));
  buf1  g1482(.din(new_new_n2105__), .dout(new_new_n2106__));
  buf1  g1483(.din(new_new_n668__), .dout(new_new_n2107__));
  buf1  g1484(.din(new_new_n2107__), .dout(new_new_n2108__));
  buf1  g1485(.din(new_new_n665__), .dout(new_new_n2109__));
  buf1  g1486(.din(new_new_n680__), .dout(new_new_n2110__));
  buf1  g1487(.din(new_new_n2110__), .dout(new_new_n2111__));
  buf1  g1488(.din(new_new_n681__), .dout(new_new_n2112__));
  buf1  g1489(.din(new_new_n684__), .dout(new_new_n2113__));
  buf1  g1490(.din(new_new_n2113__), .dout(new_new_n2114__));
  buf1  g1491(.din(new_new_n685__), .dout(new_new_n2115__));
  buf1  g1492(.din(new_new_n692__), .dout(new_new_n2116__));
  buf1  g1493(.din(new_new_n2116__), .dout(new_new_n2117__));
  buf1  g1494(.din(new_new_n688__), .dout(new_new_n2118__));
  buf1  g1495(.din(new_new_n2118__), .dout(new_new_n2119__));
  buf1  g1496(.din(new_new_n693__), .dout(new_new_n2120__));
  buf1  g1497(.din(new_new_n689__), .dout(new_new_n2121__));
  buf1  g1498(.din(new_new_n705__), .dout(new_new_n2122__));
  buf1  g1499(.din(new_new_n704__), .dout(new_new_n2123__));
  buf1  g1500(.din(new_new_n2123__), .dout(new_new_n2124__));
  buf1  g1501(.din(new_new_n709__), .dout(new_new_n2125__));
  buf1  g1502(.din(new_new_n708__), .dout(new_new_n2126__));
  buf1  g1503(.din(new_new_n2126__), .dout(new_new_n2127__));
  buf1  g1504(.din(new_new_n701__), .dout(new_new_n2128__));
  buf1  g1505(.din(new_new_n696__), .dout(new_new_n2129__));
  buf1  g1506(.din(new_new_n2129__), .dout(new_new_n2130__));
  buf1  g1507(.din(new_new_n700__), .dout(new_new_n2131__));
  buf1  g1508(.din(new_new_n2131__), .dout(new_new_n2132__));
  buf1  g1509(.din(new_new_n697__), .dout(new_new_n2133__));
  buf1  g1510(.din(new_new_n713__), .dout(new_new_n2134__));
  buf1  g1511(.din(new_new_n712__), .dout(new_new_n2135__));
  buf1  g1512(.din(new_new_n2135__), .dout(new_new_n2136__));
  buf1  g1513(.din(new_new_n717__), .dout(new_new_n2137__));
  buf1  g1514(.din(new_new_n716__), .dout(new_new_n2138__));
  buf1  g1515(.din(new_new_n2138__), .dout(new_new_n2139__));
  always @ (posedge clock) begin
    n621_lo <= n3365;
    n630_lo <= n3368;
    n633_lo <= n3371;
    n642_lo <= n3374;
    n645_lo <= n3377;
    n654_lo <= n3380;
    n657_lo <= n3383;
    n666_lo <= n3386;
    n669_lo <= n3389;
    n678_lo <= n3392;
    n681_lo <= n3395;
    n690_lo <= n3398;
    n693_lo <= n3401;
    n702_lo <= n3404;
    n705_lo <= n3407;
    n714_lo <= n3410;
    n717_lo <= n3413;
    n726_lo <= n3416;
    n729_lo <= n3419;
    n738_lo <= n3422;
    n741_lo <= n3425;
    n750_lo <= n3428;
    n753_lo <= n3431;
    n762_lo <= n3434;
    n765_lo <= n3437;
    n774_lo <= n3440;
    n777_lo <= n3443;
    n786_lo <= n3446;
    n789_lo <= n3449;
    n798_lo <= n3452;
    n801_lo <= n3455;
    n810_lo <= n3458;
    n813_lo <= n3461;
    n822_lo <= n3464;
    n825_lo <= n3467;
    n834_lo <= n3470;
    n837_lo <= n3473;
    n846_lo <= n3476;
    n849_lo <= n3479;
    n858_lo <= n3482;
    n861_lo <= n3485;
    n870_lo <= n3488;
    n873_lo <= n3491;
    n882_lo <= n3494;
    n885_lo <= n3497;
    n894_lo <= n3500;
    n897_lo <= n3503;
    n906_lo <= n3506;
    n909_lo <= n3509;
    n918_lo <= n3512;
    n921_lo <= n3515;
    n930_lo <= n3518;
    n933_lo <= n3521;
    n942_lo <= n3524;
    n945_lo <= n3527;
    n954_lo <= n3530;
    n957_lo <= n3533;
    n966_lo <= n3536;
    n969_lo <= n3539;
    n978_lo <= n3542;
    n981_lo <= n3545;
    n990_lo <= n3548;
    n993_lo <= n3551;
    n1002_lo <= n3554;
    n1005_lo <= n3557;
    n1017_lo <= n3560;
    n1029_lo <= n3563;
    n1041_lo <= n3566;
    n1053_lo <= n3569;
    n1065_lo <= n3572;
    n1077_lo <= n3575;
    n1089_lo <= n3578;
    n1101_lo <= n3581;
    n602_o2 <= n3584;
    n639_o2 <= n3587;
    n678_o2 <= n3590;
    n658_o2 <= n3593;
    n783_o2 <= n3596;
    n802_o2 <= n3599;
    n726_o2 <= n3602;
    n763_o2 <= n3605;
    n1644_o2 <= n3608;
    n1645_o2 <= n3611;
    n1646_o2 <= n3614;
    n1647_o2 <= n3617;
    n1648_o2 <= n3620;
    n1649_o2 <= n3623;
    n1650_o2 <= n3626;
    n1651_o2 <= n3629;
    n1652_o2 <= n3632;
    n1653_o2 <= n3635;
    n1654_o2 <= n3638;
    n1655_o2 <= n3641;
    n1656_o2 <= n3644;
    n1657_o2 <= n3647;
    n1658_o2 <= n3650;
    n1659_o2 <= n3653;
    n1660_o2 <= n3656;
    n1661_o2 <= n3659;
    n1662_o2 <= n3662;
    n1663_o2 <= n3665;
    n1664_o2 <= n3668;
    n1665_o2 <= n3671;
    n1666_o2 <= n3674;
    n1667_o2 <= n3677;
    n1668_o2 <= n3680;
    n1669_o2 <= n3683;
    n1670_o2 <= n3686;
    n1671_o2 <= n3689;
    n1672_o2 <= n3692;
    n1673_o2 <= n3695;
    n1674_o2 <= n3698;
    n1675_o2 <= n3701;
    n685_o2 <= n3704;
    n680_o2 <= n3707;
    n822_o2 <= n3710;
    n843_o2 <= n3713;
    n842_o2 <= n3716;
    n681_o2 <= n3719;
    n684_o2 <= n3722;
    n686_o2 <= n3725;
    n823_o2 <= n3728;
    n683_o2 <= n3731;
    n688_o2 <= n3734;
    n803_o2 <= n3737;
    n862_o2 <= n3740;
    n764_o2 <= n3743;
    n863_o2 <= n3746;
    n886_o2 <= n3749;
    lo002_buf_o2 <= n3752;
    lo006_buf_o2 <= n3755;
    lo010_buf_o2 <= n3758;
    lo014_buf_o2 <= n3761;
    lo018_buf_o2 <= n3764;
    lo022_buf_o2 <= n3767;
    lo026_buf_o2 <= n3770;
    lo030_buf_o2 <= n3773;
    lo034_buf_o2 <= n3776;
    lo038_buf_o2 <= n3779;
    lo042_buf_o2 <= n3782;
    lo046_buf_o2 <= n3785;
    lo050_buf_o2 <= n3788;
    lo054_buf_o2 <= n3791;
    lo058_buf_o2 <= n3794;
    lo062_buf_o2 <= n3797;
    lo066_buf_o2 <= n3800;
    lo070_buf_o2 <= n3803;
    lo074_buf_o2 <= n3806;
    lo078_buf_o2 <= n3809;
    lo082_buf_o2 <= n3812;
    lo086_buf_o2 <= n3815;
    lo090_buf_o2 <= n3818;
    lo094_buf_o2 <= n3821;
    lo098_buf_o2 <= n3824;
    lo102_buf_o2 <= n3827;
    lo106_buf_o2 <= n3830;
    lo110_buf_o2 <= n3833;
    lo114_buf_o2 <= n3836;
    lo118_buf_o2 <= n3839;
    lo122_buf_o2 <= n3842;
    lo126_buf_o2 <= n3845;
    n600_o2 <= n3848;
    n601_o2 <= n3851;
    n637_o2 <= n3854;
    n638_o2 <= n3857;
    n676_o2 <= n3860;
    n677_o2 <= n3863;
    n656_o2 <= n3866;
    n657_o2 <= n3869;
    n781_o2 <= n3872;
    n782_o2 <= n3875;
    n800_o2 <= n3878;
    n801_o2 <= n3881;
    n724_o2 <= n3884;
    n725_o2 <= n3887;
    n761_o2 <= n3890;
    n762_o2 <= n3893;
    lo129_buf_o2 <= n3896;
    lo133_buf_o2 <= n3899;
    lo137_buf_o2 <= n3902;
    lo141_buf_o2 <= n3905;
    lo145_buf_o2 <= n3908;
    lo149_buf_o2 <= n3911;
    lo153_buf_o2 <= n3914;
    lo157_buf_o2 <= n3917;
    lo161_buf_o2 <= n3920;
    n571_o2 <= n3923;
    n708_o2 <= n3926;
    n608_o2 <= n3929;
    n665_o2 <= n3932;
    n705_o2 <= n3935;
    n645_o2 <= n3938;
    n745_o2 <= n3941;
    n742_o2 <= n3944;
    n568_o2 <= n3947;
    n717_o2 <= n3950;
    n605_o2 <= n3953;
    n662_o2 <= n3956;
    n714_o2 <= n3959;
    n642_o2 <= n3962;
    n754_o2 <= n3965;
    n751_o2 <= n3968;
    n584_o2 <= n3971;
    n770_o2 <= n3974;
    n789_o2 <= n3977;
    n581_o2 <= n3980;
    n695_o2 <= n3983;
    n732_o2 <= n3986;
    n593_o2 <= n3989;
    n590_o2 <= n3992;
    n630_o2 <= n3995;
    n767_o2 <= n3998;
    n786_o2 <= n4001;
    n627_o2 <= n4004;
    n692_o2 <= n4007;
    n729_o2 <= n4010;
    n621_o2 <= n4013;
    n618_o2 <= n4016;
  end
  initial begin
    n621_lo <= 1'b0;
    n630_lo <= 1'b0;
    n633_lo <= 1'b0;
    n642_lo <= 1'b0;
    n645_lo <= 1'b0;
    n654_lo <= 1'b0;
    n657_lo <= 1'b0;
    n666_lo <= 1'b0;
    n669_lo <= 1'b0;
    n678_lo <= 1'b0;
    n681_lo <= 1'b0;
    n690_lo <= 1'b0;
    n693_lo <= 1'b0;
    n702_lo <= 1'b0;
    n705_lo <= 1'b0;
    n714_lo <= 1'b0;
    n717_lo <= 1'b0;
    n726_lo <= 1'b0;
    n729_lo <= 1'b0;
    n738_lo <= 1'b0;
    n741_lo <= 1'b0;
    n750_lo <= 1'b0;
    n753_lo <= 1'b0;
    n762_lo <= 1'b0;
    n765_lo <= 1'b0;
    n774_lo <= 1'b0;
    n777_lo <= 1'b0;
    n786_lo <= 1'b0;
    n789_lo <= 1'b0;
    n798_lo <= 1'b0;
    n801_lo <= 1'b0;
    n810_lo <= 1'b0;
    n813_lo <= 1'b0;
    n822_lo <= 1'b0;
    n825_lo <= 1'b0;
    n834_lo <= 1'b0;
    n837_lo <= 1'b0;
    n846_lo <= 1'b0;
    n849_lo <= 1'b0;
    n858_lo <= 1'b0;
    n861_lo <= 1'b0;
    n870_lo <= 1'b0;
    n873_lo <= 1'b0;
    n882_lo <= 1'b0;
    n885_lo <= 1'b0;
    n894_lo <= 1'b0;
    n897_lo <= 1'b0;
    n906_lo <= 1'b0;
    n909_lo <= 1'b0;
    n918_lo <= 1'b0;
    n921_lo <= 1'b0;
    n930_lo <= 1'b0;
    n933_lo <= 1'b0;
    n942_lo <= 1'b0;
    n945_lo <= 1'b0;
    n954_lo <= 1'b0;
    n957_lo <= 1'b0;
    n966_lo <= 1'b0;
    n969_lo <= 1'b0;
    n978_lo <= 1'b0;
    n981_lo <= 1'b0;
    n990_lo <= 1'b0;
    n993_lo <= 1'b0;
    n1002_lo <= 1'b0;
    n1005_lo <= 1'b0;
    n1017_lo <= 1'b0;
    n1029_lo <= 1'b0;
    n1041_lo <= 1'b0;
    n1053_lo <= 1'b0;
    n1065_lo <= 1'b0;
    n1077_lo <= 1'b0;
    n1089_lo <= 1'b0;
    n1101_lo <= 1'b0;
    n602_o2 <= 1'b0;
    n639_o2 <= 1'b0;
    n678_o2 <= 1'b0;
    n658_o2 <= 1'b0;
    n783_o2 <= 1'b0;
    n802_o2 <= 1'b0;
    n726_o2 <= 1'b0;
    n763_o2 <= 1'b0;
    n1644_o2 <= 1'b0;
    n1645_o2 <= 1'b0;
    n1646_o2 <= 1'b0;
    n1647_o2 <= 1'b0;
    n1648_o2 <= 1'b0;
    n1649_o2 <= 1'b0;
    n1650_o2 <= 1'b0;
    n1651_o2 <= 1'b0;
    n1652_o2 <= 1'b0;
    n1653_o2 <= 1'b0;
    n1654_o2 <= 1'b0;
    n1655_o2 <= 1'b0;
    n1656_o2 <= 1'b0;
    n1657_o2 <= 1'b0;
    n1658_o2 <= 1'b0;
    n1659_o2 <= 1'b0;
    n1660_o2 <= 1'b0;
    n1661_o2 <= 1'b0;
    n1662_o2 <= 1'b0;
    n1663_o2 <= 1'b0;
    n1664_o2 <= 1'b0;
    n1665_o2 <= 1'b0;
    n1666_o2 <= 1'b0;
    n1667_o2 <= 1'b0;
    n1668_o2 <= 1'b0;
    n1669_o2 <= 1'b0;
    n1670_o2 <= 1'b0;
    n1671_o2 <= 1'b0;
    n1672_o2 <= 1'b0;
    n1673_o2 <= 1'b0;
    n1674_o2 <= 1'b0;
    n1675_o2 <= 1'b0;
    n685_o2 <= 1'b0;
    n680_o2 <= 1'b0;
    n822_o2 <= 1'b0;
    n843_o2 <= 1'b0;
    n842_o2 <= 1'b0;
    n681_o2 <= 1'b0;
    n684_o2 <= 1'b0;
    n686_o2 <= 1'b0;
    n823_o2 <= 1'b0;
    n683_o2 <= 1'b0;
    n688_o2 <= 1'b0;
    n803_o2 <= 1'b0;
    n862_o2 <= 1'b0;
    n764_o2 <= 1'b0;
    n863_o2 <= 1'b0;
    n886_o2 <= 1'b0;
    lo002_buf_o2 <= 1'b0;
    lo006_buf_o2 <= 1'b0;
    lo010_buf_o2 <= 1'b0;
    lo014_buf_o2 <= 1'b0;
    lo018_buf_o2 <= 1'b0;
    lo022_buf_o2 <= 1'b0;
    lo026_buf_o2 <= 1'b0;
    lo030_buf_o2 <= 1'b0;
    lo034_buf_o2 <= 1'b0;
    lo038_buf_o2 <= 1'b0;
    lo042_buf_o2 <= 1'b0;
    lo046_buf_o2 <= 1'b0;
    lo050_buf_o2 <= 1'b0;
    lo054_buf_o2 <= 1'b0;
    lo058_buf_o2 <= 1'b0;
    lo062_buf_o2 <= 1'b0;
    lo066_buf_o2 <= 1'b0;
    lo070_buf_o2 <= 1'b0;
    lo074_buf_o2 <= 1'b0;
    lo078_buf_o2 <= 1'b0;
    lo082_buf_o2 <= 1'b0;
    lo086_buf_o2 <= 1'b0;
    lo090_buf_o2 <= 1'b0;
    lo094_buf_o2 <= 1'b0;
    lo098_buf_o2 <= 1'b0;
    lo102_buf_o2 <= 1'b0;
    lo106_buf_o2 <= 1'b0;
    lo110_buf_o2 <= 1'b0;
    lo114_buf_o2 <= 1'b0;
    lo118_buf_o2 <= 1'b0;
    lo122_buf_o2 <= 1'b0;
    lo126_buf_o2 <= 1'b0;
    n600_o2 <= 1'b0;
    n601_o2 <= 1'b0;
    n637_o2 <= 1'b0;
    n638_o2 <= 1'b0;
    n676_o2 <= 1'b0;
    n677_o2 <= 1'b0;
    n656_o2 <= 1'b0;
    n657_o2 <= 1'b0;
    n781_o2 <= 1'b0;
    n782_o2 <= 1'b0;
    n800_o2 <= 1'b0;
    n801_o2 <= 1'b0;
    n724_o2 <= 1'b0;
    n725_o2 <= 1'b0;
    n761_o2 <= 1'b0;
    n762_o2 <= 1'b0;
    lo129_buf_o2 <= 1'b0;
    lo133_buf_o2 <= 1'b0;
    lo137_buf_o2 <= 1'b0;
    lo141_buf_o2 <= 1'b0;
    lo145_buf_o2 <= 1'b0;
    lo149_buf_o2 <= 1'b0;
    lo153_buf_o2 <= 1'b0;
    lo157_buf_o2 <= 1'b0;
    lo161_buf_o2 <= 1'b0;
    n571_o2 <= 1'b0;
    n708_o2 <= 1'b0;
    n608_o2 <= 1'b0;
    n665_o2 <= 1'b0;
    n705_o2 <= 1'b0;
    n645_o2 <= 1'b0;
    n745_o2 <= 1'b0;
    n742_o2 <= 1'b0;
    n568_o2 <= 1'b0;
    n717_o2 <= 1'b0;
    n605_o2 <= 1'b0;
    n662_o2 <= 1'b0;
    n714_o2 <= 1'b0;
    n642_o2 <= 1'b0;
    n754_o2 <= 1'b0;
    n751_o2 <= 1'b0;
    n584_o2 <= 1'b0;
    n770_o2 <= 1'b0;
    n789_o2 <= 1'b0;
    n581_o2 <= 1'b0;
    n695_o2 <= 1'b0;
    n732_o2 <= 1'b0;
    n593_o2 <= 1'b0;
    n590_o2 <= 1'b0;
    n630_o2 <= 1'b0;
    n767_o2 <= 1'b0;
    n786_o2 <= 1'b0;
    n627_o2 <= 1'b0;
    n692_o2 <= 1'b0;
    n729_o2 <= 1'b0;
    n621_o2 <= 1'b0;
    n618_o2 <= 1'b0;
  end
endmodule


