
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  G42,
  G43,
  G44,
  G45,
  G46,
  G47,
  G48,
  G49,
  G50,
  G51,
  G52,
  G53,
  G54,
  G55,
  G56,
  G57,
  G58,
  G59,
  G60,
  n492_lo,
  n495_lo,
  n498_lo,
  n501_lo,
  n516_lo,
  n528_lo,
  n540_lo,
  n543_lo,
  n546_lo,
  n549_lo,
  n552_lo,
  n564_lo,
  n600_lo,
  n603_lo,
  n606_lo,
  n609_lo,
  n615_lo,
  n618_lo,
  n621_lo,
  n627_lo,
  n630_lo,
  n633_lo,
  n639_lo,
  n642_lo,
  n645_lo,
  n648_lo,
  n660_lo,
  n672_lo,
  n675_lo,
  n678_lo,
  n681_lo,
  n684_lo,
  n687_lo,
  n690_lo,
  n693_lo,
  n696_lo,
  n699_lo,
  n702_lo,
  n705_lo,
  n708_lo,
  n711_lo,
  n714_lo,
  n717_lo,
  n720_lo,
  n723_lo,
  n726_lo,
  n729_lo,
  n732_lo,
  n735_lo,
  n738_lo,
  n741_lo,
  n744_lo,
  n747_lo,
  n750_lo,
  n753_lo,
  n756_lo,
  n759_lo,
  n762_lo,
  n765_lo,
  n768_lo,
  n771_lo,
  n774_lo,
  n777_lo,
  n780_lo,
  n783_lo,
  n786_lo,
  n792_lo,
  n795_lo,
  n798_lo,
  n807_lo,
  n816_lo,
  n819_lo,
  n828_lo,
  n831_lo,
  n843_lo,
  n846_lo,
  n849_lo,
  n852_lo,
  n855_lo,
  n858_lo,
  n861_lo,
  n864_lo,
  n867_lo,
  n870_lo,
  n879_lo,
  n882_lo,
  n891_lo,
  n903_lo,
  n915_lo,
  n918_lo,
  n951_lo,
  n954_lo,
  n957_lo,
  n960_lo,
  n963_lo,
  n966_lo,
  n969_lo,
  n972_lo,
  n975_lo,
  n978_lo,
  n981_lo,
  n984_lo,
  n987_lo,
  n990_lo,
  n993_lo,
  n996_lo,
  n999_lo,
  n1002_lo,
  n1008_lo,
  n1011_lo,
  n1014_lo,
  n1020_lo,
  n1023_lo,
  n1032_lo,
  n1035_lo,
  n1044_lo,
  n1047_lo,
  n1050_lo,
  n1053_lo,
  n1056_lo,
  n1059_lo,
  n1062_lo,
  n1065_lo,
  n1068_lo,
  n1071_lo,
  n1074_lo,
  n1077_lo,
  n1080_lo,
  n1083_lo,
  n1086_lo,
  n1089_lo,
  n1092_lo,
  n1095_lo,
  n1098_lo,
  n1101_lo,
  n1104_lo,
  n1107_lo,
  n1110_lo,
  n1113_lo,
  n1116_lo,
  n1119_lo,
  n1122_lo,
  n1125_lo,
  n1128_lo,
  n1131_lo,
  n1134_lo,
  n1137_lo,
  n1143_lo,
  n1146_lo,
  n1149_lo,
  n1152_lo,
  n1155_lo,
  n1164_lo,
  n1167_lo,
  n1170_lo,
  n1173_lo,
  n1176_lo,
  n1188_lo,
  n563_inv,
  n1429_o2,
  n1427_o2,
  n1471_o2,
  n1476_o2,
  n1499_o2,
  n1500_o2,
  n1501_o2,
  n1516_o2,
  n1517_o2,
  n1562_o2,
  n1563_o2,
  n1564_o2,
  n1582_o2,
  n1583_o2,
  n1618_o2,
  n1622_o2,
  n1502_o2,
  n1503_o2,
  n1504_o2,
  n1505_o2,
  n1506_o2,
  n1512_o2,
  n1513_o2,
  n1514_o2,
  n1515_o2,
  n1644_o2,
  n1647_o2,
  n1527_o2,
  n650_inv,
  n653_inv,
  n656_inv,
  n1567_o2,
  n955_o2,
  n1568_o2,
  n1037_o2,
  n960_o2,
  n1587_o2,
  n1040_o2,
  n1039_o2,
  n1589_o2,
  n1624_o2,
  n1643_o2,
  n1038_o2,
  n1645_o2,
  n1029_o2,
  n701_inv,
  n1662_o2,
  n1663_o2,
  n710_inv,
  n813_o2,
  lo114_buf_o2,
  n1031_o2,
  lo186_buf_o2,
  n1042_o2,
  n728_inv,
  n917_o2,
  n734_inv,
  n1649_o2,
  n1650_o2,
  n1651_o2,
  n1652_o2,
  n1653_o2,
  lo138_buf_o2,
  n1664_o2,
  n1665_o2,
  n1666_o2,
  n1667_o2,
  n944_o2,
  n770_inv,
  n1672_o2,
  n776_inv,
  n1679_o2,
  n782_inv,
  n785_inv,
  lo110_buf_o2,
  lo134_buf_o2,
  n1030_o2,
  lo182_buf_o2,
  n830_o2,
  n1021_o2,
  n806_inv,
  n809_inv,
  n946_o2,
  lo038_buf_o2,
  lo238_buf_o2,
  n1010_o2,
  n1006_o2,
  n907_o2,
  n902_o2,
  lo154_buf_o2,
  n836_inv,
  n839_inv,
  lo122_buf_o2,
  n845_inv,
  n904_o2,
  lo106_buf_o2,
  n980_o2,
  n1023_o2,
  lo178_buf_o2,
  n981_o2,
  n837_o2,
  n1013_o2,
  n840_o2,
  n849_o2,
  n852_o2,
  n864_o2,
  n867_o2,
  n1044_o2,
  n876_o2,
  n893_inv,
  n879_o2,
  n925_o2,
  n902_inv,
  lo146_buf_o2,
  n1026_o2,
  n1032_o2,
  lo118_buf_o2,
  n917_inv,
  lo190_buf_o2,
  n1036_o2,
  n926_inv,
  n929_inv,
  lo002_buf_o2,
  lo014_buf_o2,
  lo030_buf_o2,
  lo034_buf_o2,
  lo042_buf_o2,
  lo113_buf_o2,
  lo185_buf_o2,
  n939_o2,
  n941_o2,
  lo142_buf_o2,
  lo230_buf_o2,
  lo006_buf_o2,
  lo018_buf_o2,
  lo022_buf_o2,
  lo066_buf_o2,
  n977_inv,
  n826_o2,
  n892_o2,
  lo152_buf_o2,
  n896_o2,
  n905_o2,
  n995_inv,
  lo037_buf_o2,
  lo237_buf_o2,
  lo062_buf_o2,
  n1007_inv,
  n1010_inv,
  n891_o2,
  G855,
  G856,
  G857,
  G858,
  G859,
  G860,
  G861,
  G862,
  G863,
  G864,
  G865,
  G866,
  G867,
  G868,
  G869,
  G870,
  G871,
  G872,
  G873,
  G874,
  G875,
  G876,
  G877,
  G878,
  G879,
  G880,
  n1654_li007_li007,
  n1657_li008_li008,
  n1660_li009_li009,
  n1663_li010_li010,
  n1678_li015_li015,
  n1690_li019_li019,
  n1702_li023_li023,
  n1705_li024_li024,
  n1708_li025_li025,
  n1711_li026_li026,
  n1714_li027_li027,
  n1726_li031_li031,
  n1762_li043_li043,
  n1765_li044_li044,
  n1768_li045_li045,
  n1771_li046_li046,
  n1777_li048_li048,
  n1780_li049_li049,
  n1783_li050_li050,
  n1789_li052_li052,
  n1792_li053_li053,
  n1795_li054_li054,
  n1801_li056_li056,
  n1804_li057_li057,
  n1807_li058_li058,
  n1810_li059_li059,
  n1822_li063_li063,
  n1834_li067_li067,
  n1837_li068_li068,
  n1840_li069_li069,
  n1843_li070_li070,
  n1846_li071_li071,
  n1849_li072_li072,
  n1852_li073_li073,
  n1855_li074_li074,
  n1858_li075_li075,
  n1861_li076_li076,
  n1864_li077_li077,
  n1867_li078_li078,
  n1870_li079_li079,
  n1873_li080_li080,
  n1876_li081_li081,
  n1879_li082_li082,
  n1882_li083_li083,
  n1885_li084_li084,
  n1888_li085_li085,
  n1891_li086_li086,
  n1894_li087_li087,
  n1897_li088_li088,
  n1900_li089_li089,
  n1903_li090_li090,
  n1906_li091_li091,
  n1909_li092_li092,
  n1912_li093_li093,
  n1915_li094_li094,
  n1918_li095_li095,
  n1921_li096_li096,
  n1924_li097_li097,
  n1927_li098_li098,
  n1930_li099_li099,
  n1933_li100_li100,
  n1936_li101_li101,
  n1939_li102_li102,
  n1942_li103_li103,
  n1945_li104_li104,
  n1948_li105_li105,
  n1954_li107_li107,
  n1957_li108_li108,
  n1960_li109_li109,
  n1969_li112_li112,
  n1978_li115_li115,
  n1981_li116_li116,
  n1990_li119_li119,
  n1993_li120_li120,
  n2005_li124_li124,
  n2008_li125_li125,
  n2011_li126_li126,
  n2014_li127_li127,
  n2017_li128_li128,
  n2020_li129_li129,
  n2023_li130_li130,
  n2026_li131_li131,
  n2029_li132_li132,
  n2032_li133_li133,
  n2041_li136_li136,
  n2044_li137_li137,
  n2053_li140_li140,
  n2065_li144_li144,
  n2077_li148_li148,
  n2080_li149_li149,
  n2113_li160_li160,
  n2116_li161_li161,
  n2119_li162_li162,
  n2122_li163_li163,
  n2125_li164_li164,
  n2128_li165_li165,
  n2131_li166_li166,
  n2134_li167_li167,
  n2137_li168_li168,
  n2140_li169_li169,
  n2143_li170_li170,
  n2146_li171_li171,
  n2149_li172_li172,
  n2152_li173_li173,
  n2155_li174_li174,
  n2158_li175_li175,
  n2161_li176_li176,
  n2164_li177_li177,
  n2170_li179_li179,
  n2173_li180_li180,
  n2176_li181_li181,
  n2182_li183_li183,
  n2185_li184_li184,
  n2194_li187_li187,
  n2197_li188_li188,
  n2206_li191_li191,
  n2209_li192_li192,
  n2212_li193_li193,
  n2215_li194_li194,
  n2218_li195_li195,
  n2221_li196_li196,
  n2224_li197_li197,
  n2227_li198_li198,
  n2230_li199_li199,
  n2233_li200_li200,
  n2236_li201_li201,
  n2239_li202_li202,
  n2242_li203_li203,
  n2245_li204_li204,
  n2248_li205_li205,
  n2251_li206_li206,
  n2254_li207_li207,
  n2257_li208_li208,
  n2260_li209_li209,
  n2263_li210_li210,
  n2266_li211_li211,
  n2269_li212_li212,
  n2272_li213_li213,
  n2275_li214_li214,
  n2278_li215_li215,
  n2281_li216_li216,
  n2284_li217_li217,
  n2287_li218_li218,
  n2290_li219_li219,
  n2293_li220_li220,
  n2296_li221_li221,
  n2299_li222_li222,
  n2305_li224_li224,
  n2308_li225_li225,
  n2311_li226_li226,
  n2314_li227_li227,
  n2317_li228_li228,
  n2326_li231_li231,
  n2329_li232_li232,
  n2332_li233_li233,
  n2335_li234_li234,
  n2338_li235_li235,
  n2350_li239_li239,
  n1428_i2,
  n1429_i2,
  n1427_i2,
  n1471_i2,
  n1476_i2,
  n1499_i2,
  n1500_i2,
  n1501_i2,
  n1516_i2,
  n1517_i2,
  n1562_i2,
  n1563_i2,
  n1564_i2,
  n1582_i2,
  n1583_i2,
  n1618_i2,
  n1622_i2,
  n1502_i2,
  n1503_i2,
  n1504_i2,
  n1505_i2,
  n1506_i2,
  n1512_i2,
  n1513_i2,
  n1514_i2,
  n1515_i2,
  n1644_i2,
  n1647_i2,
  n1527_i2,
  n1526_i2,
  n1528_i2,
  n1529_i2,
  n1567_i2,
  n955_i2,
  n1568_i2,
  n1037_i2,
  n960_i2,
  n1587_i2,
  n1040_i2,
  n1039_i2,
  n1589_i2,
  n1624_i2,
  n1643_i2,
  n1038_i2,
  n1645_i2,
  n1029_i2,
  n1648_i2,
  n1662_i2,
  n1663_i2,
  n1668_i2,
  n813_i2,
  lo114_buf_i2,
  n1031_i2,
  lo186_buf_i2,
  n1042_i2,
  n911_i2,
  n917_i2,
  n942_i2,
  n1649_i2,
  n1650_i2,
  n1651_i2,
  n1652_i2,
  n1653_i2,
  lo138_buf_i2,
  n1664_i2,
  n1665_i2,
  n1666_i2,
  n1667_i2,
  n944_i2,
  n945_i2,
  n1672_i2,
  n1676_i2,
  n1679_i2,
  n1680_i2,
  n1681_i2,
  lo110_buf_i2,
  lo134_buf_i2,
  n1030_i2,
  lo182_buf_i2,
  n830_i2,
  n1021_i2,
  n943_i2,
  n936_i2,
  n946_i2,
  lo038_buf_i2,
  lo238_buf_i2,
  n1010_i2,
  n1006_i2,
  n907_i2,
  n902_i2,
  lo154_buf_i2,
  n938_i2,
  n947_i2,
  lo122_buf_i2,
  n899_i2,
  n904_i2,
  lo106_buf_i2,
  n980_i2,
  n1023_i2,
  lo178_buf_i2,
  n981_i2,
  n837_i2,
  n1013_i2,
  n840_i2,
  n849_i2,
  n852_i2,
  n864_i2,
  n867_i2,
  n1044_i2,
  n876_i2,
  n937_i2,
  n879_i2,
  n925_i2,
  n954_i2,
  lo146_buf_i2,
  n1026_i2,
  n1032_i2,
  lo118_buf_i2,
  n957_i2,
  lo190_buf_i2,
  n1036_i2,
  n949_i2,
  n910_i2,
  lo002_buf_i2,
  lo014_buf_i2,
  lo030_buf_i2,
  lo034_buf_i2,
  lo042_buf_i2,
  lo113_buf_i2,
  lo185_buf_i2,
  n939_i2,
  n941_i2,
  lo142_buf_i2,
  lo230_buf_i2,
  lo006_buf_i2,
  lo018_buf_i2,
  lo022_buf_i2,
  lo066_buf_i2,
  n913_i2,
  n826_i2,
  n892_i2,
  lo152_buf_i2,
  n896_i2,
  n905_i2,
  n821_i2,
  lo037_buf_i2,
  lo237_buf_i2,
  lo062_buf_i2,
  n827_i2,
  n809_i2,
  n891_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input G42;input G43;input G44;input G45;input G46;input G47;input G48;input G49;input G50;input G51;input G52;input G53;input G54;input G55;input G56;input G57;input G58;input G59;input G60;input n492_lo;input n495_lo;input n498_lo;input n501_lo;input n516_lo;input n528_lo;input n540_lo;input n543_lo;input n546_lo;input n549_lo;input n552_lo;input n564_lo;input n600_lo;input n603_lo;input n606_lo;input n609_lo;input n615_lo;input n618_lo;input n621_lo;input n627_lo;input n630_lo;input n633_lo;input n639_lo;input n642_lo;input n645_lo;input n648_lo;input n660_lo;input n672_lo;input n675_lo;input n678_lo;input n681_lo;input n684_lo;input n687_lo;input n690_lo;input n693_lo;input n696_lo;input n699_lo;input n702_lo;input n705_lo;input n708_lo;input n711_lo;input n714_lo;input n717_lo;input n720_lo;input n723_lo;input n726_lo;input n729_lo;input n732_lo;input n735_lo;input n738_lo;input n741_lo;input n744_lo;input n747_lo;input n750_lo;input n753_lo;input n756_lo;input n759_lo;input n762_lo;input n765_lo;input n768_lo;input n771_lo;input n774_lo;input n777_lo;input n780_lo;input n783_lo;input n786_lo;input n792_lo;input n795_lo;input n798_lo;input n807_lo;input n816_lo;input n819_lo;input n828_lo;input n831_lo;input n843_lo;input n846_lo;input n849_lo;input n852_lo;input n855_lo;input n858_lo;input n861_lo;input n864_lo;input n867_lo;input n870_lo;input n879_lo;input n882_lo;input n891_lo;input n903_lo;input n915_lo;input n918_lo;input n951_lo;input n954_lo;input n957_lo;input n960_lo;input n963_lo;input n966_lo;input n969_lo;input n972_lo;input n975_lo;input n978_lo;input n981_lo;input n984_lo;input n987_lo;input n990_lo;input n993_lo;input n996_lo;input n999_lo;input n1002_lo;input n1008_lo;input n1011_lo;input n1014_lo;input n1020_lo;input n1023_lo;input n1032_lo;input n1035_lo;input n1044_lo;input n1047_lo;input n1050_lo;input n1053_lo;input n1056_lo;input n1059_lo;input n1062_lo;input n1065_lo;input n1068_lo;input n1071_lo;input n1074_lo;input n1077_lo;input n1080_lo;input n1083_lo;input n1086_lo;input n1089_lo;input n1092_lo;input n1095_lo;input n1098_lo;input n1101_lo;input n1104_lo;input n1107_lo;input n1110_lo;input n1113_lo;input n1116_lo;input n1119_lo;input n1122_lo;input n1125_lo;input n1128_lo;input n1131_lo;input n1134_lo;input n1137_lo;input n1143_lo;input n1146_lo;input n1149_lo;input n1152_lo;input n1155_lo;input n1164_lo;input n1167_lo;input n1170_lo;input n1173_lo;input n1176_lo;input n1188_lo;input n563_inv;input n1429_o2;input n1427_o2;input n1471_o2;input n1476_o2;input n1499_o2;input n1500_o2;input n1501_o2;input n1516_o2;input n1517_o2;input n1562_o2;input n1563_o2;input n1564_o2;input n1582_o2;input n1583_o2;input n1618_o2;input n1622_o2;input n1502_o2;input n1503_o2;input n1504_o2;input n1505_o2;input n1506_o2;input n1512_o2;input n1513_o2;input n1514_o2;input n1515_o2;input n1644_o2;input n1647_o2;input n1527_o2;input n650_inv;input n653_inv;input n656_inv;input n1567_o2;input n955_o2;input n1568_o2;input n1037_o2;input n960_o2;input n1587_o2;input n1040_o2;input n1039_o2;input n1589_o2;input n1624_o2;input n1643_o2;input n1038_o2;input n1645_o2;input n1029_o2;input n701_inv;input n1662_o2;input n1663_o2;input n710_inv;input n813_o2;input lo114_buf_o2;input n1031_o2;input lo186_buf_o2;input n1042_o2;input n728_inv;input n917_o2;input n734_inv;input n1649_o2;input n1650_o2;input n1651_o2;input n1652_o2;input n1653_o2;input lo138_buf_o2;input n1664_o2;input n1665_o2;input n1666_o2;input n1667_o2;input n944_o2;input n770_inv;input n1672_o2;input n776_inv;input n1679_o2;input n782_inv;input n785_inv;input lo110_buf_o2;input lo134_buf_o2;input n1030_o2;input lo182_buf_o2;input n830_o2;input n1021_o2;input n806_inv;input n809_inv;input n946_o2;input lo038_buf_o2;input lo238_buf_o2;input n1010_o2;input n1006_o2;input n907_o2;input n902_o2;input lo154_buf_o2;input n836_inv;input n839_inv;input lo122_buf_o2;input n845_inv;input n904_o2;input lo106_buf_o2;input n980_o2;input n1023_o2;input lo178_buf_o2;input n981_o2;input n837_o2;input n1013_o2;input n840_o2;input n849_o2;input n852_o2;input n864_o2;input n867_o2;input n1044_o2;input n876_o2;input n893_inv;input n879_o2;input n925_o2;input n902_inv;input lo146_buf_o2;input n1026_o2;input n1032_o2;input lo118_buf_o2;input n917_inv;input lo190_buf_o2;input n1036_o2;input n926_inv;input n929_inv;input lo002_buf_o2;input lo014_buf_o2;input lo030_buf_o2;input lo034_buf_o2;input lo042_buf_o2;input lo113_buf_o2;input lo185_buf_o2;input n939_o2;input n941_o2;input lo142_buf_o2;input lo230_buf_o2;input lo006_buf_o2;input lo018_buf_o2;input lo022_buf_o2;input lo066_buf_o2;input n977_inv;input n826_o2;input n892_o2;input lo152_buf_o2;input n896_o2;input n905_o2;input n995_inv;input lo037_buf_o2;input lo237_buf_o2;input lo062_buf_o2;input n1007_inv;input n1010_inv;input n891_o2;
  output G855;output G856;output G857;output G858;output G859;output G860;output G861;output G862;output G863;output G864;output G865;output G866;output G867;output G868;output G869;output G870;output G871;output G872;output G873;output G874;output G875;output G876;output G877;output G878;output G879;output G880;output n1654_li007_li007;output n1657_li008_li008;output n1660_li009_li009;output n1663_li010_li010;output n1678_li015_li015;output n1690_li019_li019;output n1702_li023_li023;output n1705_li024_li024;output n1708_li025_li025;output n1711_li026_li026;output n1714_li027_li027;output n1726_li031_li031;output n1762_li043_li043;output n1765_li044_li044;output n1768_li045_li045;output n1771_li046_li046;output n1777_li048_li048;output n1780_li049_li049;output n1783_li050_li050;output n1789_li052_li052;output n1792_li053_li053;output n1795_li054_li054;output n1801_li056_li056;output n1804_li057_li057;output n1807_li058_li058;output n1810_li059_li059;output n1822_li063_li063;output n1834_li067_li067;output n1837_li068_li068;output n1840_li069_li069;output n1843_li070_li070;output n1846_li071_li071;output n1849_li072_li072;output n1852_li073_li073;output n1855_li074_li074;output n1858_li075_li075;output n1861_li076_li076;output n1864_li077_li077;output n1867_li078_li078;output n1870_li079_li079;output n1873_li080_li080;output n1876_li081_li081;output n1879_li082_li082;output n1882_li083_li083;output n1885_li084_li084;output n1888_li085_li085;output n1891_li086_li086;output n1894_li087_li087;output n1897_li088_li088;output n1900_li089_li089;output n1903_li090_li090;output n1906_li091_li091;output n1909_li092_li092;output n1912_li093_li093;output n1915_li094_li094;output n1918_li095_li095;output n1921_li096_li096;output n1924_li097_li097;output n1927_li098_li098;output n1930_li099_li099;output n1933_li100_li100;output n1936_li101_li101;output n1939_li102_li102;output n1942_li103_li103;output n1945_li104_li104;output n1948_li105_li105;output n1954_li107_li107;output n1957_li108_li108;output n1960_li109_li109;output n1969_li112_li112;output n1978_li115_li115;output n1981_li116_li116;output n1990_li119_li119;output n1993_li120_li120;output n2005_li124_li124;output n2008_li125_li125;output n2011_li126_li126;output n2014_li127_li127;output n2017_li128_li128;output n2020_li129_li129;output n2023_li130_li130;output n2026_li131_li131;output n2029_li132_li132;output n2032_li133_li133;output n2041_li136_li136;output n2044_li137_li137;output n2053_li140_li140;output n2065_li144_li144;output n2077_li148_li148;output n2080_li149_li149;output n2113_li160_li160;output n2116_li161_li161;output n2119_li162_li162;output n2122_li163_li163;output n2125_li164_li164;output n2128_li165_li165;output n2131_li166_li166;output n2134_li167_li167;output n2137_li168_li168;output n2140_li169_li169;output n2143_li170_li170;output n2146_li171_li171;output n2149_li172_li172;output n2152_li173_li173;output n2155_li174_li174;output n2158_li175_li175;output n2161_li176_li176;output n2164_li177_li177;output n2170_li179_li179;output n2173_li180_li180;output n2176_li181_li181;output n2182_li183_li183;output n2185_li184_li184;output n2194_li187_li187;output n2197_li188_li188;output n2206_li191_li191;output n2209_li192_li192;output n2212_li193_li193;output n2215_li194_li194;output n2218_li195_li195;output n2221_li196_li196;output n2224_li197_li197;output n2227_li198_li198;output n2230_li199_li199;output n2233_li200_li200;output n2236_li201_li201;output n2239_li202_li202;output n2242_li203_li203;output n2245_li204_li204;output n2248_li205_li205;output n2251_li206_li206;output n2254_li207_li207;output n2257_li208_li208;output n2260_li209_li209;output n2263_li210_li210;output n2266_li211_li211;output n2269_li212_li212;output n2272_li213_li213;output n2275_li214_li214;output n2278_li215_li215;output n2281_li216_li216;output n2284_li217_li217;output n2287_li218_li218;output n2290_li219_li219;output n2293_li220_li220;output n2296_li221_li221;output n2299_li222_li222;output n2305_li224_li224;output n2308_li225_li225;output n2311_li226_li226;output n2314_li227_li227;output n2317_li228_li228;output n2326_li231_li231;output n2329_li232_li232;output n2332_li233_li233;output n2335_li234_li234;output n2338_li235_li235;output n2350_li239_li239;output n1428_i2;output n1429_i2;output n1427_i2;output n1471_i2;output n1476_i2;output n1499_i2;output n1500_i2;output n1501_i2;output n1516_i2;output n1517_i2;output n1562_i2;output n1563_i2;output n1564_i2;output n1582_i2;output n1583_i2;output n1618_i2;output n1622_i2;output n1502_i2;output n1503_i2;output n1504_i2;output n1505_i2;output n1506_i2;output n1512_i2;output n1513_i2;output n1514_i2;output n1515_i2;output n1644_i2;output n1647_i2;output n1527_i2;output n1526_i2;output n1528_i2;output n1529_i2;output n1567_i2;output n955_i2;output n1568_i2;output n1037_i2;output n960_i2;output n1587_i2;output n1040_i2;output n1039_i2;output n1589_i2;output n1624_i2;output n1643_i2;output n1038_i2;output n1645_i2;output n1029_i2;output n1648_i2;output n1662_i2;output n1663_i2;output n1668_i2;output n813_i2;output lo114_buf_i2;output n1031_i2;output lo186_buf_i2;output n1042_i2;output n911_i2;output n917_i2;output n942_i2;output n1649_i2;output n1650_i2;output n1651_i2;output n1652_i2;output n1653_i2;output lo138_buf_i2;output n1664_i2;output n1665_i2;output n1666_i2;output n1667_i2;output n944_i2;output n945_i2;output n1672_i2;output n1676_i2;output n1679_i2;output n1680_i2;output n1681_i2;output lo110_buf_i2;output lo134_buf_i2;output n1030_i2;output lo182_buf_i2;output n830_i2;output n1021_i2;output n943_i2;output n936_i2;output n946_i2;output lo038_buf_i2;output lo238_buf_i2;output n1010_i2;output n1006_i2;output n907_i2;output n902_i2;output lo154_buf_i2;output n938_i2;output n947_i2;output lo122_buf_i2;output n899_i2;output n904_i2;output lo106_buf_i2;output n980_i2;output n1023_i2;output lo178_buf_i2;output n981_i2;output n837_i2;output n1013_i2;output n840_i2;output n849_i2;output n852_i2;output n864_i2;output n867_i2;output n1044_i2;output n876_i2;output n937_i2;output n879_i2;output n925_i2;output n954_i2;output lo146_buf_i2;output n1026_i2;output n1032_i2;output lo118_buf_i2;output n957_i2;output lo190_buf_i2;output n1036_i2;output n949_i2;output n910_i2;output lo002_buf_i2;output lo014_buf_i2;output lo030_buf_i2;output lo034_buf_i2;output lo042_buf_i2;output lo113_buf_i2;output lo185_buf_i2;output n939_i2;output n941_i2;output lo142_buf_i2;output lo230_buf_i2;output lo006_buf_i2;output lo018_buf_i2;output lo022_buf_i2;output lo066_buf_i2;output n913_i2;output n826_i2;output n892_i2;output lo152_buf_i2;output n896_i2;output n905_i2;output n821_i2;output lo037_buf_i2;output lo237_buf_i2;output lo062_buf_i2;output n827_i2;output n809_i2;output n891_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire G51_p;
  wire G51_n;
  wire G52_p;
  wire G52_n;
  wire G53_p;
  wire G53_n;
  wire G54_p;
  wire G54_n;
  wire G55_p;
  wire G55_n;
  wire G56_p;
  wire G56_n;
  wire G57_p;
  wire G57_n;
  wire G58_p;
  wire G58_n;
  wire G59_p;
  wire G59_n;
  wire G60_p;
  wire G60_n;
  wire n492_lo_p;
  wire n492_lo_n;
  wire n495_lo_p;
  wire n495_lo_n;
  wire n498_lo_p;
  wire n498_lo_n;
  wire n501_lo_p;
  wire n501_lo_n;
  wire n516_lo_p;
  wire n516_lo_n;
  wire n528_lo_p;
  wire n528_lo_n;
  wire n540_lo_p;
  wire n540_lo_n;
  wire n543_lo_p;
  wire n543_lo_n;
  wire n546_lo_p;
  wire n546_lo_n;
  wire n549_lo_p;
  wire n549_lo_n;
  wire n552_lo_p;
  wire n552_lo_n;
  wire n564_lo_p;
  wire n564_lo_n;
  wire n600_lo_p;
  wire n600_lo_n;
  wire n603_lo_p;
  wire n603_lo_n;
  wire n606_lo_p;
  wire n606_lo_n;
  wire n609_lo_p;
  wire n609_lo_n;
  wire n615_lo_p;
  wire n615_lo_n;
  wire n618_lo_p;
  wire n618_lo_n;
  wire n621_lo_p;
  wire n621_lo_n;
  wire n627_lo_p;
  wire n627_lo_n;
  wire n630_lo_p;
  wire n630_lo_n;
  wire n633_lo_p;
  wire n633_lo_n;
  wire n639_lo_p;
  wire n639_lo_n;
  wire n642_lo_p;
  wire n642_lo_n;
  wire n645_lo_p;
  wire n645_lo_n;
  wire n648_lo_p;
  wire n648_lo_n;
  wire n660_lo_p;
  wire n660_lo_n;
  wire n672_lo_p;
  wire n672_lo_n;
  wire n675_lo_p;
  wire n675_lo_n;
  wire n678_lo_p;
  wire n678_lo_n;
  wire n681_lo_p;
  wire n681_lo_n;
  wire n684_lo_p;
  wire n684_lo_n;
  wire n687_lo_p;
  wire n687_lo_n;
  wire n690_lo_p;
  wire n690_lo_n;
  wire n693_lo_p;
  wire n693_lo_n;
  wire n696_lo_p;
  wire n696_lo_n;
  wire n699_lo_p;
  wire n699_lo_n;
  wire n702_lo_p;
  wire n702_lo_n;
  wire n705_lo_p;
  wire n705_lo_n;
  wire n708_lo_p;
  wire n708_lo_n;
  wire n711_lo_p;
  wire n711_lo_n;
  wire n714_lo_p;
  wire n714_lo_n;
  wire n717_lo_p;
  wire n717_lo_n;
  wire n720_lo_p;
  wire n720_lo_n;
  wire n723_lo_p;
  wire n723_lo_n;
  wire n726_lo_p;
  wire n726_lo_n;
  wire n729_lo_p;
  wire n729_lo_n;
  wire n732_lo_p;
  wire n732_lo_n;
  wire n735_lo_p;
  wire n735_lo_n;
  wire n738_lo_p;
  wire n738_lo_n;
  wire n741_lo_p;
  wire n741_lo_n;
  wire n744_lo_p;
  wire n744_lo_n;
  wire n747_lo_p;
  wire n747_lo_n;
  wire n750_lo_p;
  wire n750_lo_n;
  wire n753_lo_p;
  wire n753_lo_n;
  wire n756_lo_p;
  wire n756_lo_n;
  wire n759_lo_p;
  wire n759_lo_n;
  wire n762_lo_p;
  wire n762_lo_n;
  wire n765_lo_p;
  wire n765_lo_n;
  wire n768_lo_p;
  wire n768_lo_n;
  wire n771_lo_p;
  wire n771_lo_n;
  wire n774_lo_p;
  wire n774_lo_n;
  wire n777_lo_p;
  wire n777_lo_n;
  wire n780_lo_p;
  wire n780_lo_n;
  wire n783_lo_p;
  wire n783_lo_n;
  wire n786_lo_p;
  wire n786_lo_n;
  wire n792_lo_p;
  wire n792_lo_n;
  wire n795_lo_p;
  wire n795_lo_n;
  wire n798_lo_p;
  wire n798_lo_n;
  wire n807_lo_p;
  wire n807_lo_n;
  wire n816_lo_p;
  wire n816_lo_n;
  wire n819_lo_p;
  wire n819_lo_n;
  wire n828_lo_p;
  wire n828_lo_n;
  wire n831_lo_p;
  wire n831_lo_n;
  wire n843_lo_p;
  wire n843_lo_n;
  wire n846_lo_p;
  wire n846_lo_n;
  wire n849_lo_p;
  wire n849_lo_n;
  wire n852_lo_p;
  wire n852_lo_n;
  wire n855_lo_p;
  wire n855_lo_n;
  wire n858_lo_p;
  wire n858_lo_n;
  wire n861_lo_p;
  wire n861_lo_n;
  wire n864_lo_p;
  wire n864_lo_n;
  wire n867_lo_p;
  wire n867_lo_n;
  wire n870_lo_p;
  wire n870_lo_n;
  wire n879_lo_p;
  wire n879_lo_n;
  wire n882_lo_p;
  wire n882_lo_n;
  wire n891_lo_p;
  wire n891_lo_n;
  wire n903_lo_p;
  wire n903_lo_n;
  wire n915_lo_p;
  wire n915_lo_n;
  wire n918_lo_p;
  wire n918_lo_n;
  wire n951_lo_p;
  wire n951_lo_n;
  wire n954_lo_p;
  wire n954_lo_n;
  wire n957_lo_p;
  wire n957_lo_n;
  wire n960_lo_p;
  wire n960_lo_n;
  wire n963_lo_p;
  wire n963_lo_n;
  wire n966_lo_p;
  wire n966_lo_n;
  wire n969_lo_p;
  wire n969_lo_n;
  wire n972_lo_p;
  wire n972_lo_n;
  wire n975_lo_p;
  wire n975_lo_n;
  wire n978_lo_p;
  wire n978_lo_n;
  wire n981_lo_p;
  wire n981_lo_n;
  wire n984_lo_p;
  wire n984_lo_n;
  wire n987_lo_p;
  wire n987_lo_n;
  wire n990_lo_p;
  wire n990_lo_n;
  wire n993_lo_p;
  wire n993_lo_n;
  wire n996_lo_p;
  wire n996_lo_n;
  wire n999_lo_p;
  wire n999_lo_n;
  wire n1002_lo_p;
  wire n1002_lo_n;
  wire n1008_lo_p;
  wire n1008_lo_n;
  wire n1011_lo_p;
  wire n1011_lo_n;
  wire n1014_lo_p;
  wire n1014_lo_n;
  wire n1020_lo_p;
  wire n1020_lo_n;
  wire n1023_lo_p;
  wire n1023_lo_n;
  wire n1032_lo_p;
  wire n1032_lo_n;
  wire n1035_lo_p;
  wire n1035_lo_n;
  wire n1044_lo_p;
  wire n1044_lo_n;
  wire n1047_lo_p;
  wire n1047_lo_n;
  wire n1050_lo_p;
  wire n1050_lo_n;
  wire n1053_lo_p;
  wire n1053_lo_n;
  wire n1056_lo_p;
  wire n1056_lo_n;
  wire n1059_lo_p;
  wire n1059_lo_n;
  wire n1062_lo_p;
  wire n1062_lo_n;
  wire n1065_lo_p;
  wire n1065_lo_n;
  wire n1068_lo_p;
  wire n1068_lo_n;
  wire n1071_lo_p;
  wire n1071_lo_n;
  wire n1074_lo_p;
  wire n1074_lo_n;
  wire n1077_lo_p;
  wire n1077_lo_n;
  wire n1080_lo_p;
  wire n1080_lo_n;
  wire n1083_lo_p;
  wire n1083_lo_n;
  wire n1086_lo_p;
  wire n1086_lo_n;
  wire n1089_lo_p;
  wire n1089_lo_n;
  wire n1092_lo_p;
  wire n1092_lo_n;
  wire n1095_lo_p;
  wire n1095_lo_n;
  wire n1098_lo_p;
  wire n1098_lo_n;
  wire n1101_lo_p;
  wire n1101_lo_n;
  wire n1104_lo_p;
  wire n1104_lo_n;
  wire n1107_lo_p;
  wire n1107_lo_n;
  wire n1110_lo_p;
  wire n1110_lo_n;
  wire n1113_lo_p;
  wire n1113_lo_n;
  wire n1116_lo_p;
  wire n1116_lo_n;
  wire n1119_lo_p;
  wire n1119_lo_n;
  wire n1122_lo_p;
  wire n1122_lo_n;
  wire n1125_lo_p;
  wire n1125_lo_n;
  wire n1128_lo_p;
  wire n1128_lo_n;
  wire n1131_lo_p;
  wire n1131_lo_n;
  wire n1134_lo_p;
  wire n1134_lo_n;
  wire n1137_lo_p;
  wire n1137_lo_n;
  wire n1143_lo_p;
  wire n1143_lo_n;
  wire n1146_lo_p;
  wire n1146_lo_n;
  wire n1149_lo_p;
  wire n1149_lo_n;
  wire n1152_lo_p;
  wire n1152_lo_n;
  wire n1155_lo_p;
  wire n1155_lo_n;
  wire n1164_lo_p;
  wire n1164_lo_n;
  wire n1167_lo_p;
  wire n1167_lo_n;
  wire n1170_lo_p;
  wire n1170_lo_n;
  wire n1173_lo_p;
  wire n1173_lo_n;
  wire n1176_lo_p;
  wire n1176_lo_n;
  wire n1188_lo_p;
  wire n1188_lo_n;
  wire n563_inv_p;
  wire n563_inv_n;
  wire n1429_o2_p;
  wire n1429_o2_n;
  wire n1427_o2_p;
  wire n1427_o2_n;
  wire n1471_o2_p;
  wire n1471_o2_n;
  wire n1476_o2_p;
  wire n1476_o2_n;
  wire n1499_o2_p;
  wire n1499_o2_n;
  wire n1500_o2_p;
  wire n1500_o2_n;
  wire n1501_o2_p;
  wire n1501_o2_n;
  wire n1516_o2_p;
  wire n1516_o2_n;
  wire n1517_o2_p;
  wire n1517_o2_n;
  wire n1562_o2_p;
  wire n1562_o2_n;
  wire n1563_o2_p;
  wire n1563_o2_n;
  wire n1564_o2_p;
  wire n1564_o2_n;
  wire n1582_o2_p;
  wire n1582_o2_n;
  wire n1583_o2_p;
  wire n1583_o2_n;
  wire n1618_o2_p;
  wire n1618_o2_n;
  wire n1622_o2_p;
  wire n1622_o2_n;
  wire n1502_o2_p;
  wire n1502_o2_n;
  wire n1503_o2_p;
  wire n1503_o2_n;
  wire n1504_o2_p;
  wire n1504_o2_n;
  wire n1505_o2_p;
  wire n1505_o2_n;
  wire n1506_o2_p;
  wire n1506_o2_n;
  wire n1512_o2_p;
  wire n1512_o2_n;
  wire n1513_o2_p;
  wire n1513_o2_n;
  wire n1514_o2_p;
  wire n1514_o2_n;
  wire n1515_o2_p;
  wire n1515_o2_n;
  wire n1644_o2_p;
  wire n1644_o2_n;
  wire n1647_o2_p;
  wire n1647_o2_n;
  wire n1527_o2_p;
  wire n1527_o2_n;
  wire n650_inv_p;
  wire n650_inv_n;
  wire n653_inv_p;
  wire n653_inv_n;
  wire n656_inv_p;
  wire n656_inv_n;
  wire n1567_o2_p;
  wire n1567_o2_n;
  wire n955_o2_p;
  wire n955_o2_n;
  wire n1568_o2_p;
  wire n1568_o2_n;
  wire n1037_o2_p;
  wire n1037_o2_n;
  wire n960_o2_p;
  wire n960_o2_n;
  wire n1587_o2_p;
  wire n1587_o2_n;
  wire n1040_o2_p;
  wire n1040_o2_n;
  wire n1039_o2_p;
  wire n1039_o2_n;
  wire n1589_o2_p;
  wire n1589_o2_n;
  wire n1624_o2_p;
  wire n1624_o2_n;
  wire n1643_o2_p;
  wire n1643_o2_n;
  wire n1038_o2_p;
  wire n1038_o2_n;
  wire n1645_o2_p;
  wire n1645_o2_n;
  wire n1029_o2_p;
  wire n1029_o2_n;
  wire n701_inv_p;
  wire n701_inv_n;
  wire n1662_o2_p;
  wire n1662_o2_n;
  wire n1663_o2_p;
  wire n1663_o2_n;
  wire n710_inv_p;
  wire n710_inv_n;
  wire n813_o2_p;
  wire n813_o2_n;
  wire lo114_buf_o2_p;
  wire lo114_buf_o2_n;
  wire n1031_o2_p;
  wire n1031_o2_n;
  wire lo186_buf_o2_p;
  wire lo186_buf_o2_n;
  wire n1042_o2_p;
  wire n1042_o2_n;
  wire n728_inv_p;
  wire n728_inv_n;
  wire n917_o2_p;
  wire n917_o2_n;
  wire n734_inv_p;
  wire n734_inv_n;
  wire n1649_o2_p;
  wire n1649_o2_n;
  wire n1650_o2_p;
  wire n1650_o2_n;
  wire n1651_o2_p;
  wire n1651_o2_n;
  wire n1652_o2_p;
  wire n1652_o2_n;
  wire n1653_o2_p;
  wire n1653_o2_n;
  wire lo138_buf_o2_p;
  wire lo138_buf_o2_n;
  wire n1664_o2_p;
  wire n1664_o2_n;
  wire n1665_o2_p;
  wire n1665_o2_n;
  wire n1666_o2_p;
  wire n1666_o2_n;
  wire n1667_o2_p;
  wire n1667_o2_n;
  wire n944_o2_p;
  wire n944_o2_n;
  wire n770_inv_p;
  wire n770_inv_n;
  wire n1672_o2_p;
  wire n1672_o2_n;
  wire n776_inv_p;
  wire n776_inv_n;
  wire n1679_o2_p;
  wire n1679_o2_n;
  wire n782_inv_p;
  wire n782_inv_n;
  wire n785_inv_p;
  wire n785_inv_n;
  wire lo110_buf_o2_p;
  wire lo110_buf_o2_n;
  wire lo134_buf_o2_p;
  wire lo134_buf_o2_n;
  wire n1030_o2_p;
  wire n1030_o2_n;
  wire lo182_buf_o2_p;
  wire lo182_buf_o2_n;
  wire n830_o2_p;
  wire n830_o2_n;
  wire n1021_o2_p;
  wire n1021_o2_n;
  wire n806_inv_p;
  wire n806_inv_n;
  wire n809_inv_p;
  wire n809_inv_n;
  wire n946_o2_p;
  wire n946_o2_n;
  wire lo038_buf_o2_p;
  wire lo038_buf_o2_n;
  wire lo238_buf_o2_p;
  wire lo238_buf_o2_n;
  wire n1010_o2_p;
  wire n1010_o2_n;
  wire n1006_o2_p;
  wire n1006_o2_n;
  wire n907_o2_p;
  wire n907_o2_n;
  wire n902_o2_p;
  wire n902_o2_n;
  wire lo154_buf_o2_p;
  wire lo154_buf_o2_n;
  wire n836_inv_p;
  wire n836_inv_n;
  wire n839_inv_p;
  wire n839_inv_n;
  wire lo122_buf_o2_p;
  wire lo122_buf_o2_n;
  wire n845_inv_p;
  wire n845_inv_n;
  wire n904_o2_p;
  wire n904_o2_n;
  wire lo106_buf_o2_p;
  wire lo106_buf_o2_n;
  wire n980_o2_p;
  wire n980_o2_n;
  wire n1023_o2_p;
  wire n1023_o2_n;
  wire lo178_buf_o2_p;
  wire lo178_buf_o2_n;
  wire n981_o2_p;
  wire n981_o2_n;
  wire n837_o2_p;
  wire n837_o2_n;
  wire n1013_o2_p;
  wire n1013_o2_n;
  wire n840_o2_p;
  wire n840_o2_n;
  wire n849_o2_p;
  wire n849_o2_n;
  wire n852_o2_p;
  wire n852_o2_n;
  wire n864_o2_p;
  wire n864_o2_n;
  wire n867_o2_p;
  wire n867_o2_n;
  wire n1044_o2_p;
  wire n1044_o2_n;
  wire n876_o2_p;
  wire n876_o2_n;
  wire n893_inv_p;
  wire n893_inv_n;
  wire n879_o2_p;
  wire n879_o2_n;
  wire n925_o2_p;
  wire n925_o2_n;
  wire n902_inv_p;
  wire n902_inv_n;
  wire lo146_buf_o2_p;
  wire lo146_buf_o2_n;
  wire n1026_o2_p;
  wire n1026_o2_n;
  wire n1032_o2_p;
  wire n1032_o2_n;
  wire lo118_buf_o2_p;
  wire lo118_buf_o2_n;
  wire n917_inv_p;
  wire n917_inv_n;
  wire lo190_buf_o2_p;
  wire lo190_buf_o2_n;
  wire n1036_o2_p;
  wire n1036_o2_n;
  wire n926_inv_p;
  wire n926_inv_n;
  wire n929_inv_p;
  wire n929_inv_n;
  wire lo002_buf_o2_p;
  wire lo002_buf_o2_n;
  wire lo014_buf_o2_p;
  wire lo014_buf_o2_n;
  wire lo030_buf_o2_p;
  wire lo030_buf_o2_n;
  wire lo034_buf_o2_p;
  wire lo034_buf_o2_n;
  wire lo042_buf_o2_p;
  wire lo042_buf_o2_n;
  wire lo113_buf_o2_p;
  wire lo113_buf_o2_n;
  wire lo185_buf_o2_p;
  wire lo185_buf_o2_n;
  wire n939_o2_p;
  wire n939_o2_n;
  wire n941_o2_p;
  wire n941_o2_n;
  wire lo142_buf_o2_p;
  wire lo142_buf_o2_n;
  wire lo230_buf_o2_p;
  wire lo230_buf_o2_n;
  wire lo006_buf_o2_p;
  wire lo006_buf_o2_n;
  wire lo018_buf_o2_p;
  wire lo018_buf_o2_n;
  wire lo022_buf_o2_p;
  wire lo022_buf_o2_n;
  wire lo066_buf_o2_p;
  wire lo066_buf_o2_n;
  wire n977_inv_p;
  wire n977_inv_n;
  wire n826_o2_p;
  wire n826_o2_n;
  wire n892_o2_p;
  wire n892_o2_n;
  wire lo152_buf_o2_p;
  wire lo152_buf_o2_n;
  wire n896_o2_p;
  wire n896_o2_n;
  wire n905_o2_p;
  wire n905_o2_n;
  wire n995_inv_p;
  wire n995_inv_n;
  wire lo037_buf_o2_p;
  wire lo037_buf_o2_n;
  wire lo237_buf_o2_p;
  wire lo237_buf_o2_n;
  wire lo062_buf_o2_p;
  wire lo062_buf_o2_n;
  wire n1007_inv_p;
  wire n1007_inv_n;
  wire n1010_inv_p;
  wire n1010_inv_n;
  wire n891_o2_p;
  wire n891_o2_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire n540_lo_n_spl_;
  wire n660_lo_n_spl_;
  wire g370_n_spl_;
  wire n552_lo_n_spl_;
  wire n552_lo_n_spl_0;
  wire n552_lo_p_spl_;
  wire g375_n_spl_;
  wire g377_n_spl_;
  wire n600_lo_n_spl_;
  wire g379_n_spl_;
  wire g383_n_spl_;
  wire g373_n_spl_;
  wire n830_o2_n_spl_;
  wire n837_o2_n_spl_;
  wire n840_o2_n_spl_;
  wire n837_o2_p_spl_;
  wire n840_o2_p_spl_;
  wire n852_lo_p_spl_;
  wire n852_lo_p_spl_0;
  wire n852_lo_p_spl_1;
  wire g392_p_spl_;
  wire n852_lo_n_spl_;
  wire n852_lo_n_spl_0;
  wire n852_lo_n_spl_1;
  wire g392_n_spl_;
  wire n849_o2_n_spl_;
  wire n852_o2_n_spl_;
  wire n849_o2_p_spl_;
  wire n852_o2_p_spl_;
  wire n864_lo_p_spl_;
  wire g398_p_spl_;
  wire n864_lo_n_spl_;
  wire g398_n_spl_;
  wire n864_o2_n_spl_;
  wire n867_o2_n_spl_;
  wire n864_o2_p_spl_;
  wire n867_o2_p_spl_;
  wire g407_p_spl_;
  wire g407_n_spl_;
  wire n876_o2_n_spl_;
  wire n879_o2_n_spl_;
  wire n876_o2_p_spl_;
  wire n879_o2_p_spl_;
  wire n1056_lo_p_spl_;
  wire g413_p_spl_;
  wire n1056_lo_n_spl_;
  wire g413_n_spl_;
  wire n1104_lo_n_spl_;
  wire n1104_lo_n_spl_0;
  wire n1104_lo_n_spl_00;
  wire n1104_lo_n_spl_01;
  wire n1104_lo_n_spl_1;
  wire n1104_lo_n_spl_10;
  wire n1104_lo_n_spl_11;
  wire n1080_lo_n_spl_;
  wire n1080_lo_n_spl_0;
  wire n1080_lo_n_spl_00;
  wire n1080_lo_n_spl_000;
  wire n1080_lo_n_spl_001;
  wire n1080_lo_n_spl_01;
  wire n1080_lo_n_spl_010;
  wire n1080_lo_n_spl_1;
  wire n1080_lo_n_spl_10;
  wire n1080_lo_n_spl_11;
  wire n1092_lo_n_spl_;
  wire n1092_lo_n_spl_0;
  wire n1092_lo_n_spl_00;
  wire n1092_lo_n_spl_01;
  wire n1092_lo_n_spl_1;
  wire n1092_lo_n_spl_10;
  wire n1092_lo_n_spl_11;
  wire n1116_lo_n_spl_;
  wire n1116_lo_n_spl_0;
  wire n1116_lo_n_spl_00;
  wire n1116_lo_n_spl_01;
  wire n1116_lo_n_spl_1;
  wire n1116_lo_n_spl_10;
  wire n1116_lo_n_spl_11;
  wire n925_o2_n_spl_;
  wire n925_o2_n_spl_0;
  wire n925_o2_n_spl_00;
  wire n925_o2_n_spl_01;
  wire n925_o2_n_spl_1;
  wire n925_o2_n_spl_10;
  wire n925_o2_n_spl_11;
  wire n1068_lo_n_spl_;
  wire n1068_lo_n_spl_0;
  wire n1068_lo_n_spl_00;
  wire n1068_lo_n_spl_01;
  wire n1068_lo_n_spl_1;
  wire n1068_lo_n_spl_10;
  wire n1128_lo_n_spl_;
  wire n1582_o2_n_spl_;
  wire g450_n_spl_;
  wire n960_lo_p_spl_;
  wire n1013_o2_p_spl_;
  wire n960_lo_n_spl_;
  wire n960_lo_n_spl_0;
  wire n1013_o2_n_spl_;
  wire n1013_o2_n_spl_0;
  wire n972_lo_n_spl_;
  wire n1021_o2_n_spl_;
  wire n1023_o2_n_spl_;
  wire n1023_o2_n_spl_0;
  wire n1044_o2_n_spl_;
  wire n1023_o2_p_spl_;
  wire n1044_o2_p_spl_;
  wire g483_n_spl_;
  wire g483_p_spl_;
  wire g482_p_spl_;
  wire g485_n_spl_;
  wire g481_n_spl_;
  wire g481_n_spl_0;
  wire n1038_o2_n_spl_;
  wire g488_n_spl_;
  wire g503_n_spl_;
  wire g518_n_spl_;
  wire n1030_o2_n_spl_;
  wire g533_n_spl_;
  wire lo178_buf_o2_n_spl_;
  wire n993_lo_n_spl_;
  wire n993_lo_n_spl_0;
  wire g549_p_spl_;
  wire g549_p_spl_0;
  wire g548_n_spl_;
  wire g550_n_spl_;
  wire n777_lo_n_spl_;
  wire n981_lo_n_spl_;
  wire n981_lo_n_spl_0;
  wire g558_p_spl_;
  wire g558_p_spl_0;
  wire g551_p_spl_;
  wire g552_p_spl_;
  wire g553_n_spl_;
  wire lo185_buf_o2_n_spl_;
  wire g565_p_spl_;
  wire g565_p_spl_0;
  wire g563_n_spl_;
  wire g564_n_spl_;
  wire g559_n_spl_;
  wire n765_lo_p_spl_;
  wire n765_lo_p_spl_0;
  wire n1589_o2_p_spl_;
  wire n1010_o2_p_spl_;
  wire lo134_buf_o2_p_spl_;
  wire n1006_o2_p_spl_;
  wire g566_p_spl_;
  wire g567_p_spl_;
  wire lo238_buf_o2_p_spl_;
  wire n1007_inv_p_spl_;
  wire n1007_inv_p_spl_0;
  wire n1007_inv_p_spl_1;
  wire lo062_buf_o2_p_spl_;
  wire n1010_inv_p_spl_;
  wire n1014_lo_n_spl_;
  wire g582_p_spl_;
  wire g582_p_spl_0;
  wire g578_n_spl_;
  wire g583_n_spl_;
  wire n892_o2_p_spl_;
  wire lo037_buf_o2_p_spl_;
  wire g591_p_spl_;
  wire n1065_lo_p_spl_;
  wire lo110_buf_o2_p_spl_;
  wire n969_lo_p_spl_;
  wire n969_lo_p_spl_0;
  wire g577_n_spl_;
  wire n1125_lo_p_spl_;
  wire n753_lo_p_spl_;
  wire n753_lo_p_spl_0;
  wire n1512_o2_p_spl_;
  wire n777_lo_p_spl_;
  wire lo106_buf_o2_p_spl_;
  wire lo114_buf_o2_p_spl_;
  wire n1643_o2_p_spl_;
  wire n957_lo_p_spl_;
  wire n981_lo_p_spl_;
  wire n993_lo_p_spl_;
  wire g560_p_spl_;
  wire g562_p_spl_;
  wire g568_n_spl_;
  wire lo182_buf_o2_p_spl_;
  wire lo178_buf_o2_p_spl_;
  wire n1645_o2_p_spl_;
  wire lo186_buf_o2_p_spl_;
  wire g571_n_spl_;
  wire n798_lo_p_spl_;
  wire n845_inv_p_spl_;
  wire n845_inv_p_spl_0;
  wire n882_lo_p_spl_;
  wire n870_lo_p_spl_;
  wire n1650_o2_p_spl_;
  wire n786_lo_p_spl_;
  wire n1002_lo_p_spl_;
  wire g644_n_spl_;
  wire g585_n_spl_;
  wire g587_n_spl_;
  wire g592_n_spl_;
  wire g593_p_spl_;
  wire g634_p_spl_;
  wire n831_lo_p_spl_;
  wire g599_n_spl_;
  wire g599_n_spl_0;
  wire lo152_buf_o2_p_spl_;
  wire g589_n_spl_;
  wire g589_n_spl_0;
  wire g601_p_spl_;
  wire g601_p_spl_0;
  wire n819_lo_p_spl_;
  wire n903_lo_p_spl_;
  wire n1035_lo_p_spl_;
  wire g657_n_spl_;
  wire G2_p_spl_;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_1;
  wire g663_n_spl_;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire G11_p_spl_;
  wire g662_n_spl_;
  wire G6_p_spl_;
  wire G17_p_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  buf

  (
    G42_p,
    G42
  );


  not

  (
    G42_n,
    G42
  );


  buf

  (
    G43_p,
    G43
  );


  not

  (
    G43_n,
    G43
  );


  buf

  (
    G44_p,
    G44
  );


  not

  (
    G44_n,
    G44
  );


  buf

  (
    G45_p,
    G45
  );


  not

  (
    G45_n,
    G45
  );


  buf

  (
    G46_p,
    G46
  );


  not

  (
    G46_n,
    G46
  );


  buf

  (
    G47_p,
    G47
  );


  not

  (
    G47_n,
    G47
  );


  buf

  (
    G48_p,
    G48
  );


  not

  (
    G48_n,
    G48
  );


  buf

  (
    G49_p,
    G49
  );


  not

  (
    G49_n,
    G49
  );


  buf

  (
    G50_p,
    G50
  );


  not

  (
    G50_n,
    G50
  );


  buf

  (
    G51_p,
    G51
  );


  not

  (
    G51_n,
    G51
  );


  buf

  (
    G52_p,
    G52
  );


  not

  (
    G52_n,
    G52
  );


  buf

  (
    G53_p,
    G53
  );


  not

  (
    G53_n,
    G53
  );


  buf

  (
    G54_p,
    G54
  );


  not

  (
    G54_n,
    G54
  );


  buf

  (
    G55_p,
    G55
  );


  not

  (
    G55_n,
    G55
  );


  buf

  (
    G56_p,
    G56
  );


  not

  (
    G56_n,
    G56
  );


  buf

  (
    G57_p,
    G57
  );


  not

  (
    G57_n,
    G57
  );


  buf

  (
    G58_p,
    G58
  );


  not

  (
    G58_n,
    G58
  );


  buf

  (
    G59_p,
    G59
  );


  not

  (
    G59_n,
    G59
  );


  buf

  (
    G60_p,
    G60
  );


  not

  (
    G60_n,
    G60
  );


  buf

  (
    n492_lo_p,
    n492_lo
  );


  not

  (
    n492_lo_n,
    n492_lo
  );


  buf

  (
    n495_lo_p,
    n495_lo
  );


  not

  (
    n495_lo_n,
    n495_lo
  );


  buf

  (
    n498_lo_p,
    n498_lo
  );


  not

  (
    n498_lo_n,
    n498_lo
  );


  buf

  (
    n501_lo_p,
    n501_lo
  );


  not

  (
    n501_lo_n,
    n501_lo
  );


  buf

  (
    n516_lo_p,
    n516_lo
  );


  not

  (
    n516_lo_n,
    n516_lo
  );


  buf

  (
    n528_lo_p,
    n528_lo
  );


  not

  (
    n528_lo_n,
    n528_lo
  );


  buf

  (
    n540_lo_p,
    n540_lo
  );


  not

  (
    n540_lo_n,
    n540_lo
  );


  buf

  (
    n543_lo_p,
    n543_lo
  );


  not

  (
    n543_lo_n,
    n543_lo
  );


  buf

  (
    n546_lo_p,
    n546_lo
  );


  not

  (
    n546_lo_n,
    n546_lo
  );


  buf

  (
    n549_lo_p,
    n549_lo
  );


  not

  (
    n549_lo_n,
    n549_lo
  );


  buf

  (
    n552_lo_p,
    n552_lo
  );


  not

  (
    n552_lo_n,
    n552_lo
  );


  buf

  (
    n564_lo_p,
    n564_lo
  );


  not

  (
    n564_lo_n,
    n564_lo
  );


  buf

  (
    n600_lo_p,
    n600_lo
  );


  not

  (
    n600_lo_n,
    n600_lo
  );


  buf

  (
    n603_lo_p,
    n603_lo
  );


  not

  (
    n603_lo_n,
    n603_lo
  );


  buf

  (
    n606_lo_p,
    n606_lo
  );


  not

  (
    n606_lo_n,
    n606_lo
  );


  buf

  (
    n609_lo_p,
    n609_lo
  );


  not

  (
    n609_lo_n,
    n609_lo
  );


  buf

  (
    n615_lo_p,
    n615_lo
  );


  not

  (
    n615_lo_n,
    n615_lo
  );


  buf

  (
    n618_lo_p,
    n618_lo
  );


  not

  (
    n618_lo_n,
    n618_lo
  );


  buf

  (
    n621_lo_p,
    n621_lo
  );


  not

  (
    n621_lo_n,
    n621_lo
  );


  buf

  (
    n627_lo_p,
    n627_lo
  );


  not

  (
    n627_lo_n,
    n627_lo
  );


  buf

  (
    n630_lo_p,
    n630_lo
  );


  not

  (
    n630_lo_n,
    n630_lo
  );


  buf

  (
    n633_lo_p,
    n633_lo
  );


  not

  (
    n633_lo_n,
    n633_lo
  );


  buf

  (
    n639_lo_p,
    n639_lo
  );


  not

  (
    n639_lo_n,
    n639_lo
  );


  buf

  (
    n642_lo_p,
    n642_lo
  );


  not

  (
    n642_lo_n,
    n642_lo
  );


  buf

  (
    n645_lo_p,
    n645_lo
  );


  not

  (
    n645_lo_n,
    n645_lo
  );


  buf

  (
    n648_lo_p,
    n648_lo
  );


  not

  (
    n648_lo_n,
    n648_lo
  );


  buf

  (
    n660_lo_p,
    n660_lo
  );


  not

  (
    n660_lo_n,
    n660_lo
  );


  buf

  (
    n672_lo_p,
    n672_lo
  );


  not

  (
    n672_lo_n,
    n672_lo
  );


  buf

  (
    n675_lo_p,
    n675_lo
  );


  not

  (
    n675_lo_n,
    n675_lo
  );


  buf

  (
    n678_lo_p,
    n678_lo
  );


  not

  (
    n678_lo_n,
    n678_lo
  );


  buf

  (
    n681_lo_p,
    n681_lo
  );


  not

  (
    n681_lo_n,
    n681_lo
  );


  buf

  (
    n684_lo_p,
    n684_lo
  );


  not

  (
    n684_lo_n,
    n684_lo
  );


  buf

  (
    n687_lo_p,
    n687_lo
  );


  not

  (
    n687_lo_n,
    n687_lo
  );


  buf

  (
    n690_lo_p,
    n690_lo
  );


  not

  (
    n690_lo_n,
    n690_lo
  );


  buf

  (
    n693_lo_p,
    n693_lo
  );


  not

  (
    n693_lo_n,
    n693_lo
  );


  buf

  (
    n696_lo_p,
    n696_lo
  );


  not

  (
    n696_lo_n,
    n696_lo
  );


  buf

  (
    n699_lo_p,
    n699_lo
  );


  not

  (
    n699_lo_n,
    n699_lo
  );


  buf

  (
    n702_lo_p,
    n702_lo
  );


  not

  (
    n702_lo_n,
    n702_lo
  );


  buf

  (
    n705_lo_p,
    n705_lo
  );


  not

  (
    n705_lo_n,
    n705_lo
  );


  buf

  (
    n708_lo_p,
    n708_lo
  );


  not

  (
    n708_lo_n,
    n708_lo
  );


  buf

  (
    n711_lo_p,
    n711_lo
  );


  not

  (
    n711_lo_n,
    n711_lo
  );


  buf

  (
    n714_lo_p,
    n714_lo
  );


  not

  (
    n714_lo_n,
    n714_lo
  );


  buf

  (
    n717_lo_p,
    n717_lo
  );


  not

  (
    n717_lo_n,
    n717_lo
  );


  buf

  (
    n720_lo_p,
    n720_lo
  );


  not

  (
    n720_lo_n,
    n720_lo
  );


  buf

  (
    n723_lo_p,
    n723_lo
  );


  not

  (
    n723_lo_n,
    n723_lo
  );


  buf

  (
    n726_lo_p,
    n726_lo
  );


  not

  (
    n726_lo_n,
    n726_lo
  );


  buf

  (
    n729_lo_p,
    n729_lo
  );


  not

  (
    n729_lo_n,
    n729_lo
  );


  buf

  (
    n732_lo_p,
    n732_lo
  );


  not

  (
    n732_lo_n,
    n732_lo
  );


  buf

  (
    n735_lo_p,
    n735_lo
  );


  not

  (
    n735_lo_n,
    n735_lo
  );


  buf

  (
    n738_lo_p,
    n738_lo
  );


  not

  (
    n738_lo_n,
    n738_lo
  );


  buf

  (
    n741_lo_p,
    n741_lo
  );


  not

  (
    n741_lo_n,
    n741_lo
  );


  buf

  (
    n744_lo_p,
    n744_lo
  );


  not

  (
    n744_lo_n,
    n744_lo
  );


  buf

  (
    n747_lo_p,
    n747_lo
  );


  not

  (
    n747_lo_n,
    n747_lo
  );


  buf

  (
    n750_lo_p,
    n750_lo
  );


  not

  (
    n750_lo_n,
    n750_lo
  );


  buf

  (
    n753_lo_p,
    n753_lo
  );


  not

  (
    n753_lo_n,
    n753_lo
  );


  buf

  (
    n756_lo_p,
    n756_lo
  );


  not

  (
    n756_lo_n,
    n756_lo
  );


  buf

  (
    n759_lo_p,
    n759_lo
  );


  not

  (
    n759_lo_n,
    n759_lo
  );


  buf

  (
    n762_lo_p,
    n762_lo
  );


  not

  (
    n762_lo_n,
    n762_lo
  );


  buf

  (
    n765_lo_p,
    n765_lo
  );


  not

  (
    n765_lo_n,
    n765_lo
  );


  buf

  (
    n768_lo_p,
    n768_lo
  );


  not

  (
    n768_lo_n,
    n768_lo
  );


  buf

  (
    n771_lo_p,
    n771_lo
  );


  not

  (
    n771_lo_n,
    n771_lo
  );


  buf

  (
    n774_lo_p,
    n774_lo
  );


  not

  (
    n774_lo_n,
    n774_lo
  );


  buf

  (
    n777_lo_p,
    n777_lo
  );


  not

  (
    n777_lo_n,
    n777_lo
  );


  buf

  (
    n780_lo_p,
    n780_lo
  );


  not

  (
    n780_lo_n,
    n780_lo
  );


  buf

  (
    n783_lo_p,
    n783_lo
  );


  not

  (
    n783_lo_n,
    n783_lo
  );


  buf

  (
    n786_lo_p,
    n786_lo
  );


  not

  (
    n786_lo_n,
    n786_lo
  );


  buf

  (
    n792_lo_p,
    n792_lo
  );


  not

  (
    n792_lo_n,
    n792_lo
  );


  buf

  (
    n795_lo_p,
    n795_lo
  );


  not

  (
    n795_lo_n,
    n795_lo
  );


  buf

  (
    n798_lo_p,
    n798_lo
  );


  not

  (
    n798_lo_n,
    n798_lo
  );


  buf

  (
    n807_lo_p,
    n807_lo
  );


  not

  (
    n807_lo_n,
    n807_lo
  );


  buf

  (
    n816_lo_p,
    n816_lo
  );


  not

  (
    n816_lo_n,
    n816_lo
  );


  buf

  (
    n819_lo_p,
    n819_lo
  );


  not

  (
    n819_lo_n,
    n819_lo
  );


  buf

  (
    n828_lo_p,
    n828_lo
  );


  not

  (
    n828_lo_n,
    n828_lo
  );


  buf

  (
    n831_lo_p,
    n831_lo
  );


  not

  (
    n831_lo_n,
    n831_lo
  );


  buf

  (
    n843_lo_p,
    n843_lo
  );


  not

  (
    n843_lo_n,
    n843_lo
  );


  buf

  (
    n846_lo_p,
    n846_lo
  );


  not

  (
    n846_lo_n,
    n846_lo
  );


  buf

  (
    n849_lo_p,
    n849_lo
  );


  not

  (
    n849_lo_n,
    n849_lo
  );


  buf

  (
    n852_lo_p,
    n852_lo
  );


  not

  (
    n852_lo_n,
    n852_lo
  );


  buf

  (
    n855_lo_p,
    n855_lo
  );


  not

  (
    n855_lo_n,
    n855_lo
  );


  buf

  (
    n858_lo_p,
    n858_lo
  );


  not

  (
    n858_lo_n,
    n858_lo
  );


  buf

  (
    n861_lo_p,
    n861_lo
  );


  not

  (
    n861_lo_n,
    n861_lo
  );


  buf

  (
    n864_lo_p,
    n864_lo
  );


  not

  (
    n864_lo_n,
    n864_lo
  );


  buf

  (
    n867_lo_p,
    n867_lo
  );


  not

  (
    n867_lo_n,
    n867_lo
  );


  buf

  (
    n870_lo_p,
    n870_lo
  );


  not

  (
    n870_lo_n,
    n870_lo
  );


  buf

  (
    n879_lo_p,
    n879_lo
  );


  not

  (
    n879_lo_n,
    n879_lo
  );


  buf

  (
    n882_lo_p,
    n882_lo
  );


  not

  (
    n882_lo_n,
    n882_lo
  );


  buf

  (
    n891_lo_p,
    n891_lo
  );


  not

  (
    n891_lo_n,
    n891_lo
  );


  buf

  (
    n903_lo_p,
    n903_lo
  );


  not

  (
    n903_lo_n,
    n903_lo
  );


  buf

  (
    n915_lo_p,
    n915_lo
  );


  not

  (
    n915_lo_n,
    n915_lo
  );


  buf

  (
    n918_lo_p,
    n918_lo
  );


  not

  (
    n918_lo_n,
    n918_lo
  );


  buf

  (
    n951_lo_p,
    n951_lo
  );


  not

  (
    n951_lo_n,
    n951_lo
  );


  buf

  (
    n954_lo_p,
    n954_lo
  );


  not

  (
    n954_lo_n,
    n954_lo
  );


  buf

  (
    n957_lo_p,
    n957_lo
  );


  not

  (
    n957_lo_n,
    n957_lo
  );


  buf

  (
    n960_lo_p,
    n960_lo
  );


  not

  (
    n960_lo_n,
    n960_lo
  );


  buf

  (
    n963_lo_p,
    n963_lo
  );


  not

  (
    n963_lo_n,
    n963_lo
  );


  buf

  (
    n966_lo_p,
    n966_lo
  );


  not

  (
    n966_lo_n,
    n966_lo
  );


  buf

  (
    n969_lo_p,
    n969_lo
  );


  not

  (
    n969_lo_n,
    n969_lo
  );


  buf

  (
    n972_lo_p,
    n972_lo
  );


  not

  (
    n972_lo_n,
    n972_lo
  );


  buf

  (
    n975_lo_p,
    n975_lo
  );


  not

  (
    n975_lo_n,
    n975_lo
  );


  buf

  (
    n978_lo_p,
    n978_lo
  );


  not

  (
    n978_lo_n,
    n978_lo
  );


  buf

  (
    n981_lo_p,
    n981_lo
  );


  not

  (
    n981_lo_n,
    n981_lo
  );


  buf

  (
    n984_lo_p,
    n984_lo
  );


  not

  (
    n984_lo_n,
    n984_lo
  );


  buf

  (
    n987_lo_p,
    n987_lo
  );


  not

  (
    n987_lo_n,
    n987_lo
  );


  buf

  (
    n990_lo_p,
    n990_lo
  );


  not

  (
    n990_lo_n,
    n990_lo
  );


  buf

  (
    n993_lo_p,
    n993_lo
  );


  not

  (
    n993_lo_n,
    n993_lo
  );


  buf

  (
    n996_lo_p,
    n996_lo
  );


  not

  (
    n996_lo_n,
    n996_lo
  );


  buf

  (
    n999_lo_p,
    n999_lo
  );


  not

  (
    n999_lo_n,
    n999_lo
  );


  buf

  (
    n1002_lo_p,
    n1002_lo
  );


  not

  (
    n1002_lo_n,
    n1002_lo
  );


  buf

  (
    n1008_lo_p,
    n1008_lo
  );


  not

  (
    n1008_lo_n,
    n1008_lo
  );


  buf

  (
    n1011_lo_p,
    n1011_lo
  );


  not

  (
    n1011_lo_n,
    n1011_lo
  );


  buf

  (
    n1014_lo_p,
    n1014_lo
  );


  not

  (
    n1014_lo_n,
    n1014_lo
  );


  buf

  (
    n1020_lo_p,
    n1020_lo
  );


  not

  (
    n1020_lo_n,
    n1020_lo
  );


  buf

  (
    n1023_lo_p,
    n1023_lo
  );


  not

  (
    n1023_lo_n,
    n1023_lo
  );


  buf

  (
    n1032_lo_p,
    n1032_lo
  );


  not

  (
    n1032_lo_n,
    n1032_lo
  );


  buf

  (
    n1035_lo_p,
    n1035_lo
  );


  not

  (
    n1035_lo_n,
    n1035_lo
  );


  buf

  (
    n1044_lo_p,
    n1044_lo
  );


  not

  (
    n1044_lo_n,
    n1044_lo
  );


  buf

  (
    n1047_lo_p,
    n1047_lo
  );


  not

  (
    n1047_lo_n,
    n1047_lo
  );


  buf

  (
    n1050_lo_p,
    n1050_lo
  );


  not

  (
    n1050_lo_n,
    n1050_lo
  );


  buf

  (
    n1053_lo_p,
    n1053_lo
  );


  not

  (
    n1053_lo_n,
    n1053_lo
  );


  buf

  (
    n1056_lo_p,
    n1056_lo
  );


  not

  (
    n1056_lo_n,
    n1056_lo
  );


  buf

  (
    n1059_lo_p,
    n1059_lo
  );


  not

  (
    n1059_lo_n,
    n1059_lo
  );


  buf

  (
    n1062_lo_p,
    n1062_lo
  );


  not

  (
    n1062_lo_n,
    n1062_lo
  );


  buf

  (
    n1065_lo_p,
    n1065_lo
  );


  not

  (
    n1065_lo_n,
    n1065_lo
  );


  buf

  (
    n1068_lo_p,
    n1068_lo
  );


  not

  (
    n1068_lo_n,
    n1068_lo
  );


  buf

  (
    n1071_lo_p,
    n1071_lo
  );


  not

  (
    n1071_lo_n,
    n1071_lo
  );


  buf

  (
    n1074_lo_p,
    n1074_lo
  );


  not

  (
    n1074_lo_n,
    n1074_lo
  );


  buf

  (
    n1077_lo_p,
    n1077_lo
  );


  not

  (
    n1077_lo_n,
    n1077_lo
  );


  buf

  (
    n1080_lo_p,
    n1080_lo
  );


  not

  (
    n1080_lo_n,
    n1080_lo
  );


  buf

  (
    n1083_lo_p,
    n1083_lo
  );


  not

  (
    n1083_lo_n,
    n1083_lo
  );


  buf

  (
    n1086_lo_p,
    n1086_lo
  );


  not

  (
    n1086_lo_n,
    n1086_lo
  );


  buf

  (
    n1089_lo_p,
    n1089_lo
  );


  not

  (
    n1089_lo_n,
    n1089_lo
  );


  buf

  (
    n1092_lo_p,
    n1092_lo
  );


  not

  (
    n1092_lo_n,
    n1092_lo
  );


  buf

  (
    n1095_lo_p,
    n1095_lo
  );


  not

  (
    n1095_lo_n,
    n1095_lo
  );


  buf

  (
    n1098_lo_p,
    n1098_lo
  );


  not

  (
    n1098_lo_n,
    n1098_lo
  );


  buf

  (
    n1101_lo_p,
    n1101_lo
  );


  not

  (
    n1101_lo_n,
    n1101_lo
  );


  buf

  (
    n1104_lo_p,
    n1104_lo
  );


  not

  (
    n1104_lo_n,
    n1104_lo
  );


  buf

  (
    n1107_lo_p,
    n1107_lo
  );


  not

  (
    n1107_lo_n,
    n1107_lo
  );


  buf

  (
    n1110_lo_p,
    n1110_lo
  );


  not

  (
    n1110_lo_n,
    n1110_lo
  );


  buf

  (
    n1113_lo_p,
    n1113_lo
  );


  not

  (
    n1113_lo_n,
    n1113_lo
  );


  buf

  (
    n1116_lo_p,
    n1116_lo
  );


  not

  (
    n1116_lo_n,
    n1116_lo
  );


  buf

  (
    n1119_lo_p,
    n1119_lo
  );


  not

  (
    n1119_lo_n,
    n1119_lo
  );


  buf

  (
    n1122_lo_p,
    n1122_lo
  );


  not

  (
    n1122_lo_n,
    n1122_lo
  );


  buf

  (
    n1125_lo_p,
    n1125_lo
  );


  not

  (
    n1125_lo_n,
    n1125_lo
  );


  buf

  (
    n1128_lo_p,
    n1128_lo
  );


  not

  (
    n1128_lo_n,
    n1128_lo
  );


  buf

  (
    n1131_lo_p,
    n1131_lo
  );


  not

  (
    n1131_lo_n,
    n1131_lo
  );


  buf

  (
    n1134_lo_p,
    n1134_lo
  );


  not

  (
    n1134_lo_n,
    n1134_lo
  );


  buf

  (
    n1137_lo_p,
    n1137_lo
  );


  not

  (
    n1137_lo_n,
    n1137_lo
  );


  buf

  (
    n1143_lo_p,
    n1143_lo
  );


  not

  (
    n1143_lo_n,
    n1143_lo
  );


  buf

  (
    n1146_lo_p,
    n1146_lo
  );


  not

  (
    n1146_lo_n,
    n1146_lo
  );


  buf

  (
    n1149_lo_p,
    n1149_lo
  );


  not

  (
    n1149_lo_n,
    n1149_lo
  );


  buf

  (
    n1152_lo_p,
    n1152_lo
  );


  not

  (
    n1152_lo_n,
    n1152_lo
  );


  buf

  (
    n1155_lo_p,
    n1155_lo
  );


  not

  (
    n1155_lo_n,
    n1155_lo
  );


  buf

  (
    n1164_lo_p,
    n1164_lo
  );


  not

  (
    n1164_lo_n,
    n1164_lo
  );


  buf

  (
    n1167_lo_p,
    n1167_lo
  );


  not

  (
    n1167_lo_n,
    n1167_lo
  );


  buf

  (
    n1170_lo_p,
    n1170_lo
  );


  not

  (
    n1170_lo_n,
    n1170_lo
  );


  buf

  (
    n1173_lo_p,
    n1173_lo
  );


  not

  (
    n1173_lo_n,
    n1173_lo
  );


  buf

  (
    n1176_lo_p,
    n1176_lo
  );


  not

  (
    n1176_lo_n,
    n1176_lo
  );


  buf

  (
    n1188_lo_p,
    n1188_lo
  );


  not

  (
    n1188_lo_n,
    n1188_lo
  );


  buf

  (
    n563_inv_p,
    n563_inv
  );


  not

  (
    n563_inv_n,
    n563_inv
  );


  buf

  (
    n1429_o2_p,
    n1429_o2
  );


  not

  (
    n1429_o2_n,
    n1429_o2
  );


  buf

  (
    n1427_o2_p,
    n1427_o2
  );


  not

  (
    n1427_o2_n,
    n1427_o2
  );


  buf

  (
    n1471_o2_p,
    n1471_o2
  );


  not

  (
    n1471_o2_n,
    n1471_o2
  );


  buf

  (
    n1476_o2_p,
    n1476_o2
  );


  not

  (
    n1476_o2_n,
    n1476_o2
  );


  buf

  (
    n1499_o2_p,
    n1499_o2
  );


  not

  (
    n1499_o2_n,
    n1499_o2
  );


  buf

  (
    n1500_o2_p,
    n1500_o2
  );


  not

  (
    n1500_o2_n,
    n1500_o2
  );


  buf

  (
    n1501_o2_p,
    n1501_o2
  );


  not

  (
    n1501_o2_n,
    n1501_o2
  );


  buf

  (
    n1516_o2_p,
    n1516_o2
  );


  not

  (
    n1516_o2_n,
    n1516_o2
  );


  buf

  (
    n1517_o2_p,
    n1517_o2
  );


  not

  (
    n1517_o2_n,
    n1517_o2
  );


  buf

  (
    n1562_o2_p,
    n1562_o2
  );


  not

  (
    n1562_o2_n,
    n1562_o2
  );


  buf

  (
    n1563_o2_p,
    n1563_o2
  );


  not

  (
    n1563_o2_n,
    n1563_o2
  );


  buf

  (
    n1564_o2_p,
    n1564_o2
  );


  not

  (
    n1564_o2_n,
    n1564_o2
  );


  buf

  (
    n1582_o2_p,
    n1582_o2
  );


  not

  (
    n1582_o2_n,
    n1582_o2
  );


  buf

  (
    n1583_o2_p,
    n1583_o2
  );


  not

  (
    n1583_o2_n,
    n1583_o2
  );


  buf

  (
    n1618_o2_p,
    n1618_o2
  );


  not

  (
    n1618_o2_n,
    n1618_o2
  );


  buf

  (
    n1622_o2_p,
    n1622_o2
  );


  not

  (
    n1622_o2_n,
    n1622_o2
  );


  buf

  (
    n1502_o2_p,
    n1502_o2
  );


  not

  (
    n1502_o2_n,
    n1502_o2
  );


  buf

  (
    n1503_o2_p,
    n1503_o2
  );


  not

  (
    n1503_o2_n,
    n1503_o2
  );


  buf

  (
    n1504_o2_p,
    n1504_o2
  );


  not

  (
    n1504_o2_n,
    n1504_o2
  );


  buf

  (
    n1505_o2_p,
    n1505_o2
  );


  not

  (
    n1505_o2_n,
    n1505_o2
  );


  buf

  (
    n1506_o2_p,
    n1506_o2
  );


  not

  (
    n1506_o2_n,
    n1506_o2
  );


  buf

  (
    n1512_o2_p,
    n1512_o2
  );


  not

  (
    n1512_o2_n,
    n1512_o2
  );


  buf

  (
    n1513_o2_p,
    n1513_o2
  );


  not

  (
    n1513_o2_n,
    n1513_o2
  );


  buf

  (
    n1514_o2_p,
    n1514_o2
  );


  not

  (
    n1514_o2_n,
    n1514_o2
  );


  buf

  (
    n1515_o2_p,
    n1515_o2
  );


  not

  (
    n1515_o2_n,
    n1515_o2
  );


  buf

  (
    n1644_o2_p,
    n1644_o2
  );


  not

  (
    n1644_o2_n,
    n1644_o2
  );


  buf

  (
    n1647_o2_p,
    n1647_o2
  );


  not

  (
    n1647_o2_n,
    n1647_o2
  );


  buf

  (
    n1527_o2_p,
    n1527_o2
  );


  not

  (
    n1527_o2_n,
    n1527_o2
  );


  buf

  (
    n650_inv_p,
    n650_inv
  );


  not

  (
    n650_inv_n,
    n650_inv
  );


  buf

  (
    n653_inv_p,
    n653_inv
  );


  not

  (
    n653_inv_n,
    n653_inv
  );


  buf

  (
    n656_inv_p,
    n656_inv
  );


  not

  (
    n656_inv_n,
    n656_inv
  );


  buf

  (
    n1567_o2_p,
    n1567_o2
  );


  not

  (
    n1567_o2_n,
    n1567_o2
  );


  buf

  (
    n955_o2_p,
    n955_o2
  );


  not

  (
    n955_o2_n,
    n955_o2
  );


  buf

  (
    n1568_o2_p,
    n1568_o2
  );


  not

  (
    n1568_o2_n,
    n1568_o2
  );


  buf

  (
    n1037_o2_p,
    n1037_o2
  );


  not

  (
    n1037_o2_n,
    n1037_o2
  );


  buf

  (
    n960_o2_p,
    n960_o2
  );


  not

  (
    n960_o2_n,
    n960_o2
  );


  buf

  (
    n1587_o2_p,
    n1587_o2
  );


  not

  (
    n1587_o2_n,
    n1587_o2
  );


  buf

  (
    n1040_o2_p,
    n1040_o2
  );


  not

  (
    n1040_o2_n,
    n1040_o2
  );


  buf

  (
    n1039_o2_p,
    n1039_o2
  );


  not

  (
    n1039_o2_n,
    n1039_o2
  );


  buf

  (
    n1589_o2_p,
    n1589_o2
  );


  not

  (
    n1589_o2_n,
    n1589_o2
  );


  buf

  (
    n1624_o2_p,
    n1624_o2
  );


  not

  (
    n1624_o2_n,
    n1624_o2
  );


  buf

  (
    n1643_o2_p,
    n1643_o2
  );


  not

  (
    n1643_o2_n,
    n1643_o2
  );


  buf

  (
    n1038_o2_p,
    n1038_o2
  );


  not

  (
    n1038_o2_n,
    n1038_o2
  );


  buf

  (
    n1645_o2_p,
    n1645_o2
  );


  not

  (
    n1645_o2_n,
    n1645_o2
  );


  buf

  (
    n1029_o2_p,
    n1029_o2
  );


  not

  (
    n1029_o2_n,
    n1029_o2
  );


  buf

  (
    n701_inv_p,
    n701_inv
  );


  not

  (
    n701_inv_n,
    n701_inv
  );


  buf

  (
    n1662_o2_p,
    n1662_o2
  );


  not

  (
    n1662_o2_n,
    n1662_o2
  );


  buf

  (
    n1663_o2_p,
    n1663_o2
  );


  not

  (
    n1663_o2_n,
    n1663_o2
  );


  buf

  (
    n710_inv_p,
    n710_inv
  );


  not

  (
    n710_inv_n,
    n710_inv
  );


  buf

  (
    n813_o2_p,
    n813_o2
  );


  not

  (
    n813_o2_n,
    n813_o2
  );


  buf

  (
    lo114_buf_o2_p,
    lo114_buf_o2
  );


  not

  (
    lo114_buf_o2_n,
    lo114_buf_o2
  );


  buf

  (
    n1031_o2_p,
    n1031_o2
  );


  not

  (
    n1031_o2_n,
    n1031_o2
  );


  buf

  (
    lo186_buf_o2_p,
    lo186_buf_o2
  );


  not

  (
    lo186_buf_o2_n,
    lo186_buf_o2
  );


  buf

  (
    n1042_o2_p,
    n1042_o2
  );


  not

  (
    n1042_o2_n,
    n1042_o2
  );


  buf

  (
    n728_inv_p,
    n728_inv
  );


  not

  (
    n728_inv_n,
    n728_inv
  );


  buf

  (
    n917_o2_p,
    n917_o2
  );


  not

  (
    n917_o2_n,
    n917_o2
  );


  buf

  (
    n734_inv_p,
    n734_inv
  );


  not

  (
    n734_inv_n,
    n734_inv
  );


  buf

  (
    n1649_o2_p,
    n1649_o2
  );


  not

  (
    n1649_o2_n,
    n1649_o2
  );


  buf

  (
    n1650_o2_p,
    n1650_o2
  );


  not

  (
    n1650_o2_n,
    n1650_o2
  );


  buf

  (
    n1651_o2_p,
    n1651_o2
  );


  not

  (
    n1651_o2_n,
    n1651_o2
  );


  buf

  (
    n1652_o2_p,
    n1652_o2
  );


  not

  (
    n1652_o2_n,
    n1652_o2
  );


  buf

  (
    n1653_o2_p,
    n1653_o2
  );


  not

  (
    n1653_o2_n,
    n1653_o2
  );


  buf

  (
    lo138_buf_o2_p,
    lo138_buf_o2
  );


  not

  (
    lo138_buf_o2_n,
    lo138_buf_o2
  );


  buf

  (
    n1664_o2_p,
    n1664_o2
  );


  not

  (
    n1664_o2_n,
    n1664_o2
  );


  buf

  (
    n1665_o2_p,
    n1665_o2
  );


  not

  (
    n1665_o2_n,
    n1665_o2
  );


  buf

  (
    n1666_o2_p,
    n1666_o2
  );


  not

  (
    n1666_o2_n,
    n1666_o2
  );


  buf

  (
    n1667_o2_p,
    n1667_o2
  );


  not

  (
    n1667_o2_n,
    n1667_o2
  );


  buf

  (
    n944_o2_p,
    n944_o2
  );


  not

  (
    n944_o2_n,
    n944_o2
  );


  buf

  (
    n770_inv_p,
    n770_inv
  );


  not

  (
    n770_inv_n,
    n770_inv
  );


  buf

  (
    n1672_o2_p,
    n1672_o2
  );


  not

  (
    n1672_o2_n,
    n1672_o2
  );


  buf

  (
    n776_inv_p,
    n776_inv
  );


  not

  (
    n776_inv_n,
    n776_inv
  );


  buf

  (
    n1679_o2_p,
    n1679_o2
  );


  not

  (
    n1679_o2_n,
    n1679_o2
  );


  buf

  (
    n782_inv_p,
    n782_inv
  );


  not

  (
    n782_inv_n,
    n782_inv
  );


  buf

  (
    n785_inv_p,
    n785_inv
  );


  not

  (
    n785_inv_n,
    n785_inv
  );


  buf

  (
    lo110_buf_o2_p,
    lo110_buf_o2
  );


  not

  (
    lo110_buf_o2_n,
    lo110_buf_o2
  );


  buf

  (
    lo134_buf_o2_p,
    lo134_buf_o2
  );


  not

  (
    lo134_buf_o2_n,
    lo134_buf_o2
  );


  buf

  (
    n1030_o2_p,
    n1030_o2
  );


  not

  (
    n1030_o2_n,
    n1030_o2
  );


  buf

  (
    lo182_buf_o2_p,
    lo182_buf_o2
  );


  not

  (
    lo182_buf_o2_n,
    lo182_buf_o2
  );


  buf

  (
    n830_o2_p,
    n830_o2
  );


  not

  (
    n830_o2_n,
    n830_o2
  );


  buf

  (
    n1021_o2_p,
    n1021_o2
  );


  not

  (
    n1021_o2_n,
    n1021_o2
  );


  buf

  (
    n806_inv_p,
    n806_inv
  );


  not

  (
    n806_inv_n,
    n806_inv
  );


  buf

  (
    n809_inv_p,
    n809_inv
  );


  not

  (
    n809_inv_n,
    n809_inv
  );


  buf

  (
    n946_o2_p,
    n946_o2
  );


  not

  (
    n946_o2_n,
    n946_o2
  );


  buf

  (
    lo038_buf_o2_p,
    lo038_buf_o2
  );


  not

  (
    lo038_buf_o2_n,
    lo038_buf_o2
  );


  buf

  (
    lo238_buf_o2_p,
    lo238_buf_o2
  );


  not

  (
    lo238_buf_o2_n,
    lo238_buf_o2
  );


  buf

  (
    n1010_o2_p,
    n1010_o2
  );


  not

  (
    n1010_o2_n,
    n1010_o2
  );


  buf

  (
    n1006_o2_p,
    n1006_o2
  );


  not

  (
    n1006_o2_n,
    n1006_o2
  );


  buf

  (
    n907_o2_p,
    n907_o2
  );


  not

  (
    n907_o2_n,
    n907_o2
  );


  buf

  (
    n902_o2_p,
    n902_o2
  );


  not

  (
    n902_o2_n,
    n902_o2
  );


  buf

  (
    lo154_buf_o2_p,
    lo154_buf_o2
  );


  not

  (
    lo154_buf_o2_n,
    lo154_buf_o2
  );


  buf

  (
    n836_inv_p,
    n836_inv
  );


  not

  (
    n836_inv_n,
    n836_inv
  );


  buf

  (
    n839_inv_p,
    n839_inv
  );


  not

  (
    n839_inv_n,
    n839_inv
  );


  buf

  (
    lo122_buf_o2_p,
    lo122_buf_o2
  );


  not

  (
    lo122_buf_o2_n,
    lo122_buf_o2
  );


  buf

  (
    n845_inv_p,
    n845_inv
  );


  not

  (
    n845_inv_n,
    n845_inv
  );


  buf

  (
    n904_o2_p,
    n904_o2
  );


  not

  (
    n904_o2_n,
    n904_o2
  );


  buf

  (
    lo106_buf_o2_p,
    lo106_buf_o2
  );


  not

  (
    lo106_buf_o2_n,
    lo106_buf_o2
  );


  buf

  (
    n980_o2_p,
    n980_o2
  );


  not

  (
    n980_o2_n,
    n980_o2
  );


  buf

  (
    n1023_o2_p,
    n1023_o2
  );


  not

  (
    n1023_o2_n,
    n1023_o2
  );


  buf

  (
    lo178_buf_o2_p,
    lo178_buf_o2
  );


  not

  (
    lo178_buf_o2_n,
    lo178_buf_o2
  );


  buf

  (
    n981_o2_p,
    n981_o2
  );


  not

  (
    n981_o2_n,
    n981_o2
  );


  buf

  (
    n837_o2_p,
    n837_o2
  );


  not

  (
    n837_o2_n,
    n837_o2
  );


  buf

  (
    n1013_o2_p,
    n1013_o2
  );


  not

  (
    n1013_o2_n,
    n1013_o2
  );


  buf

  (
    n840_o2_p,
    n840_o2
  );


  not

  (
    n840_o2_n,
    n840_o2
  );


  buf

  (
    n849_o2_p,
    n849_o2
  );


  not

  (
    n849_o2_n,
    n849_o2
  );


  buf

  (
    n852_o2_p,
    n852_o2
  );


  not

  (
    n852_o2_n,
    n852_o2
  );


  buf

  (
    n864_o2_p,
    n864_o2
  );


  not

  (
    n864_o2_n,
    n864_o2
  );


  buf

  (
    n867_o2_p,
    n867_o2
  );


  not

  (
    n867_o2_n,
    n867_o2
  );


  buf

  (
    n1044_o2_p,
    n1044_o2
  );


  not

  (
    n1044_o2_n,
    n1044_o2
  );


  buf

  (
    n876_o2_p,
    n876_o2
  );


  not

  (
    n876_o2_n,
    n876_o2
  );


  buf

  (
    n893_inv_p,
    n893_inv
  );


  not

  (
    n893_inv_n,
    n893_inv
  );


  buf

  (
    n879_o2_p,
    n879_o2
  );


  not

  (
    n879_o2_n,
    n879_o2
  );


  buf

  (
    n925_o2_p,
    n925_o2
  );


  not

  (
    n925_o2_n,
    n925_o2
  );


  buf

  (
    n902_inv_p,
    n902_inv
  );


  not

  (
    n902_inv_n,
    n902_inv
  );


  buf

  (
    lo146_buf_o2_p,
    lo146_buf_o2
  );


  not

  (
    lo146_buf_o2_n,
    lo146_buf_o2
  );


  buf

  (
    n1026_o2_p,
    n1026_o2
  );


  not

  (
    n1026_o2_n,
    n1026_o2
  );


  buf

  (
    n1032_o2_p,
    n1032_o2
  );


  not

  (
    n1032_o2_n,
    n1032_o2
  );


  buf

  (
    lo118_buf_o2_p,
    lo118_buf_o2
  );


  not

  (
    lo118_buf_o2_n,
    lo118_buf_o2
  );


  buf

  (
    n917_inv_p,
    n917_inv
  );


  not

  (
    n917_inv_n,
    n917_inv
  );


  buf

  (
    lo190_buf_o2_p,
    lo190_buf_o2
  );


  not

  (
    lo190_buf_o2_n,
    lo190_buf_o2
  );


  buf

  (
    n1036_o2_p,
    n1036_o2
  );


  not

  (
    n1036_o2_n,
    n1036_o2
  );


  buf

  (
    n926_inv_p,
    n926_inv
  );


  not

  (
    n926_inv_n,
    n926_inv
  );


  buf

  (
    n929_inv_p,
    n929_inv
  );


  not

  (
    n929_inv_n,
    n929_inv
  );


  buf

  (
    lo002_buf_o2_p,
    lo002_buf_o2
  );


  not

  (
    lo002_buf_o2_n,
    lo002_buf_o2
  );


  buf

  (
    lo014_buf_o2_p,
    lo014_buf_o2
  );


  not

  (
    lo014_buf_o2_n,
    lo014_buf_o2
  );


  buf

  (
    lo030_buf_o2_p,
    lo030_buf_o2
  );


  not

  (
    lo030_buf_o2_n,
    lo030_buf_o2
  );


  buf

  (
    lo034_buf_o2_p,
    lo034_buf_o2
  );


  not

  (
    lo034_buf_o2_n,
    lo034_buf_o2
  );


  buf

  (
    lo042_buf_o2_p,
    lo042_buf_o2
  );


  not

  (
    lo042_buf_o2_n,
    lo042_buf_o2
  );


  buf

  (
    lo113_buf_o2_p,
    lo113_buf_o2
  );


  not

  (
    lo113_buf_o2_n,
    lo113_buf_o2
  );


  buf

  (
    lo185_buf_o2_p,
    lo185_buf_o2
  );


  not

  (
    lo185_buf_o2_n,
    lo185_buf_o2
  );


  buf

  (
    n939_o2_p,
    n939_o2
  );


  not

  (
    n939_o2_n,
    n939_o2
  );


  buf

  (
    n941_o2_p,
    n941_o2
  );


  not

  (
    n941_o2_n,
    n941_o2
  );


  buf

  (
    lo142_buf_o2_p,
    lo142_buf_o2
  );


  not

  (
    lo142_buf_o2_n,
    lo142_buf_o2
  );


  buf

  (
    lo230_buf_o2_p,
    lo230_buf_o2
  );


  not

  (
    lo230_buf_o2_n,
    lo230_buf_o2
  );


  buf

  (
    lo006_buf_o2_p,
    lo006_buf_o2
  );


  not

  (
    lo006_buf_o2_n,
    lo006_buf_o2
  );


  buf

  (
    lo018_buf_o2_p,
    lo018_buf_o2
  );


  not

  (
    lo018_buf_o2_n,
    lo018_buf_o2
  );


  buf

  (
    lo022_buf_o2_p,
    lo022_buf_o2
  );


  not

  (
    lo022_buf_o2_n,
    lo022_buf_o2
  );


  buf

  (
    lo066_buf_o2_p,
    lo066_buf_o2
  );


  not

  (
    lo066_buf_o2_n,
    lo066_buf_o2
  );


  buf

  (
    n977_inv_p,
    n977_inv
  );


  not

  (
    n977_inv_n,
    n977_inv
  );


  buf

  (
    n826_o2_p,
    n826_o2
  );


  not

  (
    n826_o2_n,
    n826_o2
  );


  buf

  (
    n892_o2_p,
    n892_o2
  );


  not

  (
    n892_o2_n,
    n892_o2
  );


  buf

  (
    lo152_buf_o2_p,
    lo152_buf_o2
  );


  not

  (
    lo152_buf_o2_n,
    lo152_buf_o2
  );


  buf

  (
    n896_o2_p,
    n896_o2
  );


  not

  (
    n896_o2_n,
    n896_o2
  );


  buf

  (
    n905_o2_p,
    n905_o2
  );


  not

  (
    n905_o2_n,
    n905_o2
  );


  buf

  (
    n995_inv_p,
    n995_inv
  );


  not

  (
    n995_inv_n,
    n995_inv
  );


  buf

  (
    lo037_buf_o2_p,
    lo037_buf_o2
  );


  not

  (
    lo037_buf_o2_n,
    lo037_buf_o2
  );


  buf

  (
    lo237_buf_o2_p,
    lo237_buf_o2
  );


  not

  (
    lo237_buf_o2_n,
    lo237_buf_o2
  );


  buf

  (
    lo062_buf_o2_p,
    lo062_buf_o2
  );


  not

  (
    lo062_buf_o2_n,
    lo062_buf_o2
  );


  buf

  (
    n1007_inv_p,
    n1007_inv
  );


  not

  (
    n1007_inv_n,
    n1007_inv
  );


  buf

  (
    n1010_inv_p,
    n1010_inv
  );


  not

  (
    n1010_inv_n,
    n1010_inv
  );


  buf

  (
    n891_o2_p,
    n891_o2
  );


  not

  (
    n891_o2_n,
    n891_o2
  );


  and

  (
    g370_p,
    n540_lo_p,
    n564_lo_p
  );


  or

  (
    g370_n,
    n540_lo_n_spl_,
    n564_lo_n
  );


  or

  (
    g371_n,
    n660_lo_n_spl_,
    g370_n_spl_
  );


  or

  (
    g372_n,
    n552_lo_n_spl_0,
    n1429_o2_n
  );


  and

  (
    g373_p,
    n552_lo_p_spl_,
    g370_p
  );


  or

  (
    g373_n,
    n552_lo_n_spl_0,
    g370_n_spl_
  );


  or

  (
    g374_n,
    n684_lo_n,
    n696_lo_n
  );


  or

  (
    g375_n,
    n516_lo_n,
    n813_o2_n
  );


  or

  (
    g376_n,
    n492_lo_n,
    g375_n_spl_
  );


  or

  (
    g377_n,
    n528_lo_n,
    g375_n_spl_
  );


  or

  (
    g378_n,
    g373_p,
    g377_n_spl_
  );


  or

  (
    g379_n,
    n600_lo_n_spl_,
    n672_lo_n
  );


  or

  (
    g380_n,
    n660_lo_n_spl_,
    g379_n_spl_
  );


  or

  (
    g381_n,
    n552_lo_n_spl_,
    g379_n_spl_
  );


  and

  (
    g382_p,
    n552_lo_p_spl_,
    n1427_o2_p
  );


  or

  (
    g383_n,
    n708_lo_p,
    n720_lo_p
  );


  and

  (
    g384_p,
    n744_lo_p,
    g383_n_spl_
  );


  or

  (
    g385_n,
    g373_n_spl_,
    g377_n_spl_
  );


  or

  (
    g386_n,
    n540_lo_n_spl_,
    n830_o2_n_spl_
  );


  or

  (
    g387_n,
    n600_lo_n_spl_,
    n648_lo_n
  );


  or

  (
    g388_n,
    n830_o2_n_spl_,
    g387_n
  );


  and

  (
    g389_p,
    n732_lo_p,
    g383_n_spl_
  );


  and

  (
    g390_p,
    n837_o2_n_spl_,
    n840_o2_n_spl_
  );


  or

  (
    g390_n,
    n837_o2_p_spl_,
    n840_o2_p_spl_
  );


  and

  (
    g391_p,
    n837_o2_p_spl_,
    n840_o2_p_spl_
  );


  or

  (
    g391_n,
    n837_o2_n_spl_,
    n840_o2_n_spl_
  );


  and

  (
    g392_p,
    g390_n,
    g391_n
  );


  or

  (
    g392_n,
    g390_p,
    g391_p
  );


  and

  (
    g393_p,
    n852_lo_p_spl_0,
    g392_p_spl_
  );


  or

  (
    g393_n,
    n852_lo_n_spl_0,
    g392_n_spl_
  );


  and

  (
    g394_p,
    n852_lo_n_spl_0,
    g392_n_spl_
  );


  or

  (
    g394_n,
    n852_lo_p_spl_0,
    g392_p_spl_
  );


  and

  (
    g395_p,
    g393_n,
    g394_n
  );


  or

  (
    g395_n,
    g393_p,
    g394_p
  );


  and

  (
    g396_p,
    n849_o2_n_spl_,
    n852_o2_n_spl_
  );


  or

  (
    g396_n,
    n849_o2_p_spl_,
    n852_o2_p_spl_
  );


  and

  (
    g397_p,
    n849_o2_p_spl_,
    n852_o2_p_spl_
  );


  or

  (
    g397_n,
    n849_o2_n_spl_,
    n852_o2_n_spl_
  );


  and

  (
    g398_p,
    g396_n,
    g397_n
  );


  or

  (
    g398_n,
    g396_p,
    g397_p
  );


  and

  (
    g399_p,
    n864_lo_p_spl_,
    g398_p_spl_
  );


  or

  (
    g399_n,
    n864_lo_n_spl_,
    g398_n_spl_
  );


  and

  (
    g400_p,
    n864_lo_n_spl_,
    g398_n_spl_
  );


  or

  (
    g400_n,
    n864_lo_p_spl_,
    g398_p_spl_
  );


  and

  (
    g401_p,
    g399_n,
    g400_n
  );


  or

  (
    g401_n,
    g399_p,
    g400_p
  );


  and

  (
    g402_p,
    g395_n,
    g401_n
  );


  and

  (
    g403_p,
    g395_p,
    g401_p
  );


  or

  (
    g404_n,
    g402_p,
    g403_p
  );


  and

  (
    g405_p,
    n864_o2_n_spl_,
    n867_o2_n_spl_
  );


  or

  (
    g405_n,
    n864_o2_p_spl_,
    n867_o2_p_spl_
  );


  and

  (
    g406_p,
    n864_o2_p_spl_,
    n867_o2_p_spl_
  );


  or

  (
    g406_n,
    n864_o2_n_spl_,
    n867_o2_n_spl_
  );


  and

  (
    g407_p,
    g405_n,
    g406_n
  );


  or

  (
    g407_n,
    g405_p,
    g406_p
  );


  and

  (
    g408_p,
    n852_lo_p_spl_1,
    g407_p_spl_
  );


  or

  (
    g408_n,
    n852_lo_n_spl_1,
    g407_n_spl_
  );


  and

  (
    g409_p,
    n852_lo_n_spl_1,
    g407_n_spl_
  );


  or

  (
    g409_n,
    n852_lo_p_spl_1,
    g407_p_spl_
  );


  and

  (
    g410_p,
    g408_n,
    g409_n
  );


  or

  (
    g410_n,
    g408_p,
    g409_p
  );


  and

  (
    g411_p,
    n876_o2_n_spl_,
    n879_o2_n_spl_
  );


  or

  (
    g411_n,
    n876_o2_p_spl_,
    n879_o2_p_spl_
  );


  and

  (
    g412_p,
    n876_o2_p_spl_,
    n879_o2_p_spl_
  );


  or

  (
    g412_n,
    n876_o2_n_spl_,
    n879_o2_n_spl_
  );


  and

  (
    g413_p,
    g411_n,
    g412_n
  );


  or

  (
    g413_n,
    g411_p,
    g412_p
  );


  and

  (
    g414_p,
    n1056_lo_p_spl_,
    g413_p_spl_
  );


  or

  (
    g414_n,
    n1056_lo_n_spl_,
    g413_n_spl_
  );


  and

  (
    g415_p,
    n1056_lo_n_spl_,
    g413_n_spl_
  );


  or

  (
    g415_n,
    n1056_lo_p_spl_,
    g413_p_spl_
  );


  and

  (
    g416_p,
    g414_n,
    g415_n
  );


  or

  (
    g416_n,
    g414_p,
    g415_p
  );


  and

  (
    g417_p,
    g410_n,
    g416_n
  );


  and

  (
    g418_p,
    g410_p,
    g416_p
  );


  or

  (
    g419_n,
    g417_p,
    g418_p
  );


  and

  (
    g420_p,
    n1104_lo_n_spl_00,
    n1499_o2_p
  );


  or

  (
    g421_n,
    n1476_o2_n,
    g420_p
  );


  or

  (
    g422_n,
    n1080_lo_n_spl_000,
    n1164_lo_n
  );


  and

  (
    g423_p,
    g421_n,
    g422_n
  );


  or

  (
    g424_n,
    n1080_lo_n_spl_000,
    n1500_o2_p
  );


  and

  (
    g425_p,
    n1092_lo_n_spl_00,
    n1499_o2_n
  );


  and

  (
    g426_p,
    g424_n,
    g425_p
  );


  or

  (
    g427_n,
    g423_p,
    g426_p
  );


  or

  (
    g428_n,
    n1116_lo_n_spl_00,
    n1471_o2_n
  );


  or

  (
    g429_n,
    n1044_lo_n,
    n925_o2_n_spl_00
  );


  or

  (
    g430_n,
    n828_lo_n,
    n1068_lo_n_spl_00
  );


  or

  (
    g431_n,
    n1128_lo_n_spl_,
    n1176_lo_n
  );


  and

  (
    g432_p,
    g430_n,
    g431_n
  );


  and

  (
    g433_p,
    g429_n,
    g432_p
  );


  and

  (
    g434_p,
    g428_n,
    g433_p
  );


  and

  (
    g435_p,
    g427_n,
    g434_p
  );


  or

  (
    g436_n,
    n1080_lo_n_spl_001,
    n1647_o2_n
  );


  and

  (
    g437_p,
    n1104_lo_n_spl_00,
    n955_o2_p
  );


  or

  (
    g438_n,
    n1644_o2_n,
    g437_p
  );


  and

  (
    g439_p,
    g436_n,
    g438_n
  );


  or

  (
    g440_n,
    n1080_lo_n_spl_001,
    n960_o2_p
  );


  and

  (
    g441_p,
    n1092_lo_n_spl_00,
    n955_o2_n
  );


  and

  (
    g442_p,
    g440_n,
    g441_p
  );


  or

  (
    g443_n,
    g439_p,
    g442_p
  );


  or

  (
    g444_n,
    n1116_lo_n_spl_00,
    n1622_o2_n
  );


  or

  (
    g445_n,
    n792_lo_n,
    n1068_lo_n_spl_00
  );


  or

  (
    g446_n,
    n1008_lo_n,
    n925_o2_n_spl_00
  );


  and

  (
    g447_p,
    g445_n,
    g446_n
  );


  and

  (
    g448_p,
    g444_n,
    g447_p
  );


  and

  (
    g449_p,
    g443_n,
    g448_p
  );


  and

  (
    g450_p,
    n1582_o2_n_spl_,
    n1618_o2_p
  );


  or

  (
    g450_n,
    n1582_o2_p,
    n1618_o2_n
  );


  or

  (
    g451_n,
    n1583_o2_n,
    g450_p
  );


  or

  (
    g452_n,
    n1583_o2_p,
    g450_n_spl_
  );


  and

  (
    g453_p,
    g451_n,
    g452_n
  );


  or

  (
    g454_n,
    n1080_lo_n_spl_010,
    g453_p
  );


  or

  (
    g455_n,
    n1092_lo_n_spl_01,
    g450_n_spl_
  );


  or

  (
    g456_n,
    n1104_lo_n_spl_01,
    n1582_o2_n_spl_
  );


  or

  (
    g457_n,
    n1116_lo_n_spl_01,
    n1563_o2_n
  );


  or

  (
    g458_n,
    n1020_lo_n,
    n925_o2_n_spl_01
  );


  and

  (
    g459_p,
    n980_o2_n,
    n981_o2_n
  );


  and

  (
    g460_p,
    g458_n,
    g459_p
  );


  and

  (
    g461_p,
    g457_n,
    g460_p
  );


  and

  (
    g462_p,
    g456_n,
    g461_p
  );


  and

  (
    g463_p,
    g455_n,
    g462_p
  );


  and

  (
    g464_p,
    g454_n,
    g463_p
  );


  and

  (
    g465_p,
    n1104_lo_n_spl_01,
    n1562_o2_p
  );


  or

  (
    g466_n,
    n1516_o2_n,
    g465_p
  );


  or

  (
    g467_n,
    n1080_lo_n_spl_010,
    n1517_o2_n
  );


  and

  (
    g468_p,
    g466_n,
    g467_n
  );


  or

  (
    g469_n,
    n1080_lo_n_spl_01,
    n1564_o2_p
  );


  and

  (
    g470_p,
    n1092_lo_n_spl_01,
    n1562_o2_n
  );


  and

  (
    g471_p,
    g469_n,
    g470_p
  );


  or

  (
    g472_n,
    g468_p,
    g471_p
  );


  or

  (
    g473_n,
    n1116_lo_n_spl_01,
    n1501_o2_n
  );


  or

  (
    g474_n,
    n1032_lo_n,
    n925_o2_n_spl_01
  );


  or

  (
    g475_n,
    n816_lo_n,
    n1068_lo_n_spl_01
  );


  or

  (
    g476_n,
    n1128_lo_n_spl_,
    n1152_lo_n
  );


  and

  (
    g477_p,
    g475_n,
    g476_n
  );


  and

  (
    g478_p,
    g474_n,
    g477_p
  );


  and

  (
    g479_p,
    g473_n,
    g478_p
  );


  and

  (
    g480_p,
    g472_n,
    g479_p
  );


  and

  (
    g481_p,
    n960_lo_p_spl_,
    n1013_o2_p_spl_
  );


  or

  (
    g481_n,
    n960_lo_n_spl_0,
    n1013_o2_n_spl_0
  );


  and

  (
    g482_p,
    n960_lo_n_spl_0,
    n1013_o2_n_spl_0
  );


  or

  (
    g482_n,
    n960_lo_p_spl_,
    n1013_o2_p_spl_
  );


  and

  (
    g483_p,
    n972_lo_n_spl_,
    n1021_o2_n_spl_
  );


  or

  (
    g483_n,
    n972_lo_p,
    n1021_o2_p
  );


  and

  (
    g484_p,
    n1023_o2_n_spl_0,
    n1044_o2_n_spl_
  );


  or

  (
    g484_n,
    n1023_o2_p_spl_,
    n1044_o2_p_spl_
  );


  and

  (
    g485_p,
    g483_n_spl_,
    g484_n
  );


  or

  (
    g485_n,
    g483_p_spl_,
    g484_p
  );


  or

  (
    g486_n,
    g482_p_spl_,
    g485_n_spl_
  );


  and

  (
    g487_p,
    g481_n_spl_0,
    g486_n
  );


  and

  (
    g488_p,
    n1040_o2_p,
    n1038_o2_n_spl_
  );


  or

  (
    g488_n,
    n1040_o2_n,
    n1038_o2_p
  );


  or

  (
    g489_n,
    n1039_o2_n,
    g488_p
  );


  or

  (
    g490_n,
    n1039_o2_p,
    g488_n_spl_
  );


  and

  (
    g491_p,
    g489_n,
    g490_n
  );


  or

  (
    g492_n,
    n1080_lo_n_spl_10,
    g491_p
  );


  or

  (
    g493_n,
    n1092_lo_n_spl_10,
    g488_n_spl_
  );


  or

  (
    g494_n,
    n1104_lo_n_spl_10,
    n1038_o2_n_spl_
  );


  or

  (
    g495_n,
    n1116_lo_n_spl_10,
    n1037_o2_n
  );


  or

  (
    g496_n,
    n996_lo_n,
    n925_o2_n_spl_10
  );


  or

  (
    g497_n,
    n780_lo_n,
    n1068_lo_n_spl_01
  );


  and

  (
    g498_p,
    g496_n,
    g497_n
  );


  and

  (
    g499_p,
    g495_n,
    g498_p
  );


  and

  (
    g500_p,
    g494_n,
    g499_p
  );


  and

  (
    g501_p,
    g493_n,
    g500_p
  );


  and

  (
    g502_p,
    g492_n,
    g501_p
  );


  and

  (
    g503_p,
    g481_n_spl_0,
    g482_n
  );


  or

  (
    g503_n,
    g481_p,
    g482_p_spl_
  );


  and

  (
    g504_p,
    g485_p,
    g503_p
  );


  and

  (
    g505_p,
    g485_n_spl_,
    g503_n_spl_
  );


  or

  (
    g506_n,
    n1080_lo_n_spl_10,
    g505_p
  );


  or

  (
    g507_n,
    g504_p,
    g506_n
  );


  or

  (
    g508_n,
    n1092_lo_n_spl_10,
    g503_n_spl_
  );


  or

  (
    g509_n,
    n1104_lo_n_spl_10,
    g481_n_spl_
  );


  or

  (
    g510_n,
    n1116_lo_n_spl_10,
    n1013_o2_n_spl_
  );


  or

  (
    g511_n,
    n1068_lo_n_spl_10,
    n1188_lo_n
  );


  or

  (
    g512_n,
    n960_lo_n_spl_,
    n925_o2_n_spl_10
  );


  and

  (
    g513_p,
    g511_n,
    g512_n
  );


  and

  (
    g514_p,
    g510_n,
    g513_p
  );


  and

  (
    g515_p,
    g509_n,
    g514_p
  );


  and

  (
    g516_p,
    g508_n,
    g515_p
  );


  and

  (
    g517_p,
    g507_n,
    g516_p
  );


  and

  (
    g518_p,
    n1023_o2_n_spl_0,
    g483_n_spl_
  );


  or

  (
    g518_n,
    n1023_o2_p_spl_,
    g483_p_spl_
  );


  and

  (
    g519_p,
    n1044_o2_p_spl_,
    g518_p
  );


  and

  (
    g520_p,
    n1044_o2_n_spl_,
    g518_n_spl_
  );


  or

  (
    g521_n,
    n1080_lo_n_spl_11,
    g520_p
  );


  or

  (
    g522_n,
    g519_p,
    g521_n
  );


  or

  (
    g523_n,
    n1092_lo_n_spl_11,
    g518_n_spl_
  );


  or

  (
    g524_n,
    n1104_lo_n_spl_11,
    n1023_o2_n_spl_
  );


  or

  (
    g525_n,
    n1116_lo_n_spl_11,
    n1021_o2_n_spl_
  );


  or

  (
    g526_n,
    n756_lo_n,
    n1068_lo_n_spl_10
  );


  or

  (
    g527_n,
    n972_lo_n_spl_,
    n925_o2_n_spl_11
  );


  and

  (
    g528_p,
    g526_n,
    g527_n
  );


  and

  (
    g529_p,
    g525_n,
    g528_p
  );


  and

  (
    g530_p,
    g524_n,
    g529_p
  );


  and

  (
    g531_p,
    g523_n,
    g530_p
  );


  and

  (
    g532_p,
    g522_n,
    g531_p
  );


  and

  (
    g533_p,
    n1031_o2_p,
    n1030_o2_n_spl_
  );


  or

  (
    g533_n,
    n1031_o2_n,
    n1030_o2_p
  );


  and

  (
    g534_p,
    n1042_o2_n,
    g533_n_spl_
  );


  and

  (
    g535_p,
    n1042_o2_p,
    g533_p
  );


  or

  (
    g536_n,
    n1080_lo_n_spl_11,
    g535_p
  );


  or

  (
    g537_n,
    g534_p,
    g536_n
  );


  or

  (
    g538_n,
    n1092_lo_n_spl_11,
    g533_n_spl_
  );


  or

  (
    g539_n,
    n1104_lo_n_spl_11,
    n1030_o2_n_spl_
  );


  or

  (
    g540_n,
    n1116_lo_n_spl_11,
    n1029_o2_n
  );


  or

  (
    g541_n,
    n768_lo_n,
    n1068_lo_n_spl_1
  );


  or

  (
    g542_n,
    n984_lo_n,
    n925_o2_n_spl_11
  );


  and

  (
    g543_p,
    g541_n,
    g542_n
  );


  and

  (
    g544_p,
    g540_n,
    g543_p
  );


  and

  (
    g545_p,
    g539_n,
    g544_p
  );


  and

  (
    g546_p,
    g538_n,
    g545_p
  );


  and

  (
    g547_p,
    g537_n,
    g546_p
  );


  or

  (
    g548_n,
    lo178_buf_o2_n_spl_,
    n902_inv_n
  );


  and

  (
    g549_p,
    n1032_o2_n,
    n1036_o2_n
  );


  or

  (
    g550_n,
    n917_inv_n,
    n926_inv_n
  );


  and

  (
    g551_p,
    n993_lo_n_spl_0,
    g549_p_spl_0
  );


  and

  (
    g552_p,
    g548_n_spl_,
    g550_n_spl_
  );


  or

  (
    g553_n,
    n993_lo_n_spl_0,
    g549_p_spl_0
  );


  or

  (
    g554_n,
    n777_lo_n_spl_,
    n1589_o2_n
  );


  or

  (
    g555_n,
    n1624_o2_n,
    n1010_o2_n
  );


  and

  (
    g556_p,
    n1006_o2_n,
    n1026_o2_n
  );


  and

  (
    g557_p,
    g555_n,
    g556_p
  );


  and

  (
    g558_p,
    g554_n,
    g557_p
  );


  or

  (
    g559_n,
    n501_lo_n,
    n1502_o2_n
  );


  and

  (
    g560_p,
    n981_lo_n_spl_0,
    g558_p_spl_0
  );


  or

  (
    g561_n,
    g551_p_spl_,
    g552_p_spl_
  );


  and

  (
    g562_p,
    g553_n_spl_,
    g561_n
  );


  or

  (
    g563_n,
    lo190_buf_o2_n,
    n929_inv_n
  );


  or

  (
    g564_n,
    lo230_buf_o2_n,
    n977_inv_n
  );


  and

  (
    g565_p,
    n939_o2_n,
    n941_o2_n
  );


  and

  (
    g566_p,
    lo185_buf_o2_n_spl_,
    g565_p_spl_0
  );


  and

  (
    g567_p,
    g563_n_spl_,
    g564_n_spl_
  );


  or

  (
    g568_n,
    n981_lo_n_spl_0,
    g558_p_spl_0
  );


  or

  (
    g569_n,
    n1512_o2_n,
    n1567_o2_n
  );


  or

  (
    g570_n,
    n609_lo_n,
    g569_n
  );


  or

  (
    g571_n,
    g559_n_spl_,
    g570_n
  );


  and

  (
    g572_p,
    n765_lo_p_spl_0,
    n1589_o2_p_spl_
  );


  and

  (
    g573_p,
    n1662_o2_p,
    n1010_o2_p_spl_
  );


  and

  (
    g574_p,
    n1505_o2_p,
    lo134_buf_o2_p_spl_
  );


  or

  (
    g575_n,
    n1006_o2_p_spl_,
    g574_p
  );


  or

  (
    g576_n,
    g573_p,
    g575_n
  );


  or

  (
    g577_n,
    g572_p,
    g576_n
  );


  or

  (
    g578_n,
    lo185_buf_o2_n_spl_,
    g565_p_spl_0
  );


  or

  (
    g579_n,
    n845_inv_n,
    lo113_buf_o2_n
  );


  or

  (
    g580_n,
    n907_o2_p,
    lo142_buf_o2_n
  );


  and

  (
    g581_p,
    n904_o2_n,
    g580_n
  );


  and

  (
    g582_p,
    g579_n,
    g581_p
  );


  or

  (
    g583_n,
    g566_p_spl_,
    g567_p_spl_
  );


  or

  (
    g584_n,
    n1672_o2_p,
    lo038_buf_o2_n
  );


  or

  (
    g585_n,
    n782_inv_n,
    g584_n
  );


  or

  (
    g586_n,
    n1650_o2_n,
    lo238_buf_o2_p_spl_
  );


  or

  (
    g587_n,
    n902_o2_n,
    g586_n
  );


  and

  (
    g588_p,
    n905_o2_p,
    n1007_inv_p_spl_0
  );


  or

  (
    g589_n,
    lo002_buf_o2_n,
    g588_p
  );


  and

  (
    g590_p,
    lo062_buf_o2_p_spl_,
    n1010_inv_p_spl_
  );


  and

  (
    g591_p,
    n1007_inv_p_spl_0,
    g590_p
  );


  or

  (
    g592_n,
    n1014_lo_n_spl_,
    g582_p_spl_0
  );


  and

  (
    g593_p,
    g578_n_spl_,
    g583_n_spl_
  );


  and

  (
    g594_p,
    n892_o2_p_spl_,
    n891_o2_p
  );


  and

  (
    g595_p,
    n1007_inv_p_spl_1,
    g594_p
  );


  or

  (
    g596_n,
    n995_inv_n,
    lo062_buf_o2_n
  );


  and

  (
    g597_p,
    n826_o2_p,
    n896_o2_p
  );


  and

  (
    g598_p,
    g596_n,
    g597_p
  );


  or

  (
    g599_n,
    g595_p,
    g598_p
  );


  and

  (
    g600_p,
    lo037_buf_o2_p_spl_,
    lo237_buf_o2_n
  );


  and

  (
    g601_p,
    g591_p_spl_,
    g600_p
  );


  and

  (
    g602_p,
    n1065_lo_p_spl_,
    lo110_buf_o2_p_spl_
  );


  and

  (
    g603_p,
    n969_lo_p_spl_0,
    g577_n_spl_
  );


  and

  (
    g604_p,
    n1125_lo_p_spl_,
    n1137_lo_p
  );


  or

  (
    g605_n,
    n753_lo_p_spl_0,
    n765_lo_p_spl_0
  );


  or

  (
    g606_n,
    n753_lo_n,
    n765_lo_n
  );


  and

  (
    g607_p,
    g605_n,
    g606_n
  );


  and

  (
    g608_p,
    n753_lo_p_spl_0,
    n1589_o2_p_spl_
  );


  and

  (
    g609_p,
    n1512_o2_p_spl_,
    lo134_buf_o2_p_spl_
  );


  or

  (
    g610_n,
    n1006_o2_p_spl_,
    g609_p
  );


  and

  (
    g611_p,
    lo138_buf_o2_p,
    n1010_o2_p_spl_
  );


  or

  (
    g612_n,
    g610_n,
    g611_p
  );


  or

  (
    g613_n,
    g608_p,
    g612_n
  );


  or

  (
    g614_n,
    n777_lo_p_spl_,
    lo106_buf_o2_p_spl_
  );


  or

  (
    g615_n,
    n777_lo_n_spl_,
    lo106_buf_o2_n
  );


  and

  (
    g616_p,
    g614_n,
    g615_n
  );


  or

  (
    g617_n,
    lo114_buf_o2_p_spl_,
    lo110_buf_o2_p_spl_
  );


  or

  (
    g618_n,
    lo114_buf_o2_n,
    lo110_buf_o2_n
  );


  and

  (
    g619_p,
    g617_n,
    g618_n
  );


  or

  (
    g620_n,
    n1587_o2_p,
    n1643_o2_p_spl_
  );


  or

  (
    g621_n,
    n1587_o2_n,
    n1643_o2_n
  );


  and

  (
    g622_p,
    g620_n,
    g621_n
  );


  or

  (
    g623_n,
    n957_lo_p_spl_,
    n969_lo_p_spl_0
  );


  or

  (
    g624_n,
    n957_lo_n,
    n969_lo_n
  );


  and

  (
    g625_p,
    g623_n,
    g624_n
  );


  or

  (
    g626_n,
    n981_lo_p_spl_,
    n993_lo_p_spl_
  );


  or

  (
    g627_n,
    n981_lo_n_spl_,
    n993_lo_n_spl_
  );


  and

  (
    g628_p,
    g626_n,
    g627_n
  );


  or

  (
    g629_n,
    g560_p_spl_,
    g562_p_spl_
  );


  and

  (
    g630_p,
    g568_n_spl_,
    g629_n
  );


  or

  (
    g631_n,
    lo182_buf_o2_p_spl_,
    lo178_buf_o2_p_spl_
  );


  or

  (
    g632_n,
    lo182_buf_o2_n,
    lo178_buf_o2_n_spl_
  );


  and

  (
    g633_p,
    g631_n,
    g632_n
  );


  and

  (
    g634_p,
    n1014_lo_n_spl_,
    g582_p_spl_0
  );


  or

  (
    g635_n,
    n1645_o2_p_spl_,
    lo186_buf_o2_p_spl_
  );


  or

  (
    g636_n,
    n1645_o2_n,
    lo186_buf_o2_n
  );


  and

  (
    g637_p,
    g635_n,
    g636_n
  );


  or

  (
    g638_n,
    n621_lo_n,
    n633_lo_n
  );


  or

  (
    g639_n,
    n650_inv_n,
    g638_n
  );


  or

  (
    g640_n,
    g571_n_spl_,
    g639_n
  );


  and

  (
    g641_p,
    n798_lo_p_spl_,
    n845_inv_p_spl_0
  );


  and

  (
    g642_p,
    n882_lo_p_spl_,
    n907_o2_n
  );


  or

  (
    g643_n,
    n904_o2_p,
    g642_p
  );


  or

  (
    g644_n,
    g641_p,
    g643_n
  );


  and

  (
    g645_p,
    n870_lo_p_spl_,
    n1650_o2_p_spl_
  );


  and

  (
    g646_p,
    n786_lo_p_spl_,
    n845_inv_p_spl_0
  );


  or

  (
    g647_n,
    n1002_lo_p_spl_,
    g644_n_spl_
  );


  or

  (
    g648_n,
    lo154_buf_o2_n,
    g585_n_spl_
  );


  or

  (
    g649_n,
    n870_lo_n,
    n918_lo_n
  );


  and

  (
    g650_p,
    g587_n_spl_,
    g649_n
  );


  and

  (
    g651_p,
    g648_n,
    g650_p
  );


  and

  (
    g652_p,
    g592_n_spl_,
    g593_p_spl_
  );


  or

  (
    g653_n,
    g634_p_spl_,
    g652_p
  );


  and

  (
    g654_p,
    n831_lo_p_spl_,
    g599_n_spl_0
  );


  and

  (
    g655_p,
    lo152_buf_o2_p_spl_,
    g589_n_spl_0
  );


  or

  (
    g656_n,
    g601_p_spl_0,
    g655_p
  );


  or

  (
    g657_n,
    g654_p,
    g656_n
  );


  and

  (
    g658_p,
    n819_lo_p_spl_,
    g599_n_spl_0
  );


  and

  (
    g659_p,
    n903_lo_p_spl_,
    g589_n_spl_0
  );


  or

  (
    g660_n,
    g601_p_spl_0,
    g659_p
  );


  or

  (
    g661_n,
    n1035_lo_p_spl_,
    g657_n_spl_
  );


  or

  (
    g662_n,
    G1_n,
    G9_n
  );


  or

  (
    g663_n,
    G11_n,
    G40_n
  );


  and

  (
    g664_p,
    G2_p_spl_,
    G4_p_spl_0
  );


  and

  (
    g665_p,
    G4_p_spl_0,
    g663_n_spl_
  );


  and

  (
    g666_p,
    G8_p_spl_0,
    G11_p_spl_
  );


  or

  (
    g667_n,
    G5_n,
    g662_n_spl_
  );


  and

  (
    g668_p,
    G6_p_spl_,
    G17_p_spl_
  );


  and

  (
    g669_p,
    G4_p_spl_1,
    G8_n
  );


  and

  (
    g670_p,
    G4_n,
    G8_p_spl_0
  );


  or

  (
    g671_n,
    g669_p,
    g670_p
  );


  buf

  (
    G855,
    g371_n
  );


  buf

  (
    G856,
    g372_n
  );


  buf

  (
    G857,
    g373_n_spl_
  );


  buf

  (
    G858,
    g374_n
  );


  buf

  (
    G859,
    g376_n
  );


  not

  (
    G860,
    g378_n
  );


  not

  (
    G861,
    g380_n
  );


  not

  (
    G862,
    g381_n
  );


  buf

  (
    G863,
    g382_p
  );


  not

  (
    G864,
    g384_p
  );


  not

  (
    G865,
    g385_n
  );


  buf

  (
    G866,
    n563_inv_n
  );


  buf

  (
    G867,
    g386_n
  );


  buf

  (
    G868,
    g388_n
  );


  not

  (
    G869,
    g389_p
  );


  buf

  (
    G870,
    g404_n
  );


  buf

  (
    G871,
    g419_n
  );


  buf

  (
    G872,
    g435_p
  );


  buf

  (
    G873,
    g449_p
  );


  buf

  (
    G874,
    g464_p
  );


  buf

  (
    G875,
    g480_p
  );


  buf

  (
    G876,
    g487_p
  );


  buf

  (
    G877,
    g502_p
  );


  buf

  (
    G878,
    g517_p
  );


  buf

  (
    G879,
    g532_p
  );


  buf

  (
    G880,
    g547_p
  );


  buf

  (
    n1654_li007_li007,
    n1512_o2_p_spl_
  );


  buf

  (
    n1657_li008_li008,
    G3_p
  );


  buf

  (
    n1660_li009_li009,
    n495_lo_p
  );


  buf

  (
    n1663_li010_li010,
    n498_lo_p
  );


  buf

  (
    n1678_li015_li015,
    n1503_o2_p
  );


  buf

  (
    n1690_li019_li019,
    n1513_o2_p
  );


  buf

  (
    n1702_li023_li023,
    n1514_o2_p
  );


  buf

  (
    n1705_li024_li024,
    G7_p
  );


  buf

  (
    n1708_li025_li025,
    n543_lo_p
  );


  buf

  (
    n1711_li026_li026,
    n546_lo_p
  );


  buf

  (
    n1714_li027_li027,
    n549_lo_p
  );


  buf

  (
    n1726_li031_li031,
    n1504_o2_p
  );


  buf

  (
    n1762_li043_li043,
    n1506_o2_p
  );


  buf

  (
    n1765_li044_li044,
    G12_p
  );


  buf

  (
    n1768_li045_li045,
    n603_lo_p
  );


  buf

  (
    n1771_li046_li046,
    n606_lo_p
  );


  buf

  (
    n1777_li048_li048,
    G13_p
  );


  buf

  (
    n1780_li049_li049,
    n615_lo_p
  );


  buf

  (
    n1783_li050_li050,
    n618_lo_p
  );


  buf

  (
    n1789_li052_li052,
    G14_p
  );


  buf

  (
    n1792_li053_li053,
    n627_lo_p
  );


  buf

  (
    n1795_li054_li054,
    n630_lo_p
  );


  buf

  (
    n1801_li056_li056,
    G15_p
  );


  buf

  (
    n1804_li057_li057,
    n639_lo_p
  );


  buf

  (
    n1807_li058_li058,
    n642_lo_p
  );


  buf

  (
    n1810_li059_li059,
    n645_lo_p
  );


  buf

  (
    n1822_li063_li063,
    n1527_o2_p
  );


  buf

  (
    n1834_li067_li067,
    n1515_o2_p
  );


  buf

  (
    n1837_li068_li068,
    G18_p
  );


  buf

  (
    n1840_li069_li069,
    n675_lo_p
  );


  buf

  (
    n1843_li070_li070,
    n678_lo_p
  );


  buf

  (
    n1846_li071_li071,
    n681_lo_p
  );


  buf

  (
    n1849_li072_li072,
    G19_p
  );


  buf

  (
    n1852_li073_li073,
    n687_lo_p
  );


  buf

  (
    n1855_li074_li074,
    n690_lo_p
  );


  buf

  (
    n1858_li075_li075,
    n693_lo_p
  );


  buf

  (
    n1861_li076_li076,
    G20_p
  );


  buf

  (
    n1864_li077_li077,
    n699_lo_p
  );


  buf

  (
    n1867_li078_li078,
    n702_lo_p
  );


  buf

  (
    n1870_li079_li079,
    n705_lo_p
  );


  buf

  (
    n1873_li080_li080,
    G21_p
  );


  buf

  (
    n1876_li081_li081,
    n711_lo_p
  );


  buf

  (
    n1879_li082_li082,
    n714_lo_p
  );


  buf

  (
    n1882_li083_li083,
    n717_lo_p
  );


  buf

  (
    n1885_li084_li084,
    G22_p
  );


  buf

  (
    n1888_li085_li085,
    n723_lo_p
  );


  buf

  (
    n1891_li086_li086,
    n726_lo_p
  );


  buf

  (
    n1894_li087_li087,
    n729_lo_p
  );


  buf

  (
    n1897_li088_li088,
    G23_p
  );


  buf

  (
    n1900_li089_li089,
    n735_lo_p
  );


  buf

  (
    n1903_li090_li090,
    n738_lo_p
  );


  buf

  (
    n1906_li091_li091,
    n741_lo_p
  );


  buf

  (
    n1909_li092_li092,
    G24_p
  );


  buf

  (
    n1912_li093_li093,
    n747_lo_p
  );


  buf

  (
    n1915_li094_li094,
    n750_lo_p
  );


  buf

  (
    n1918_li095_li095,
    n753_lo_p_spl_
  );


  buf

  (
    n1921_li096_li096,
    G25_p
  );


  buf

  (
    n1924_li097_li097,
    n759_lo_p
  );


  buf

  (
    n1927_li098_li098,
    n762_lo_p
  );


  buf

  (
    n1930_li099_li099,
    n765_lo_p_spl_
  );


  buf

  (
    n1933_li100_li100,
    G26_p
  );


  buf

  (
    n1936_li101_li101,
    n771_lo_p
  );


  buf

  (
    n1939_li102_li102,
    n774_lo_p
  );


  buf

  (
    n1942_li103_li103,
    n777_lo_p_spl_
  );


  buf

  (
    n1945_li104_li104,
    G27_p
  );


  buf

  (
    n1948_li105_li105,
    n783_lo_p
  );


  buf

  (
    n1954_li107_li107,
    lo106_buf_o2_p_spl_
  );


  buf

  (
    n1957_li108_li108,
    G28_p
  );


  buf

  (
    n1960_li109_li109,
    n795_lo_p
  );


  buf

  (
    n1969_li112_li112,
    G29_p
  );


  buf

  (
    n1978_li115_li115,
    lo114_buf_o2_p_spl_
  );


  buf

  (
    n1981_li116_li116,
    G30_p
  );


  buf

  (
    n1990_li119_li119,
    n1643_o2_p_spl_
  );


  buf

  (
    n1993_li120_li120,
    G31_p
  );


  buf

  (
    n2005_li124_li124,
    G32_p
  );


  buf

  (
    n2008_li125_li125,
    n843_lo_p
  );


  buf

  (
    n2011_li126_li126,
    n846_lo_p
  );


  buf

  (
    n2014_li127_li127,
    n849_lo_p
  );


  buf

  (
    n2017_li128_li128,
    G33_p
  );


  buf

  (
    n2020_li129_li129,
    n855_lo_p
  );


  buf

  (
    n2023_li130_li130,
    n858_lo_p
  );


  buf

  (
    n2026_li131_li131,
    n861_lo_p
  );


  buf

  (
    n2029_li132_li132,
    G34_p
  );


  buf

  (
    n2032_li133_li133,
    n867_lo_p
  );


  buf

  (
    n2041_li136_li136,
    G35_p
  );


  buf

  (
    n2044_li137_li137,
    n879_lo_p
  );


  buf

  (
    n2053_li140_li140,
    G36_p
  );


  buf

  (
    n2065_li144_li144,
    G37_p
  );


  buf

  (
    n2077_li148_li148,
    G38_p
  );


  buf

  (
    n2080_li149_li149,
    n915_lo_p
  );


  buf

  (
    n2113_li160_li160,
    G41_p
  );


  buf

  (
    n2116_li161_li161,
    n951_lo_p
  );


  buf

  (
    n2119_li162_li162,
    n954_lo_p
  );


  buf

  (
    n2122_li163_li163,
    n957_lo_p_spl_
  );


  buf

  (
    n2125_li164_li164,
    G42_p
  );


  buf

  (
    n2128_li165_li165,
    n963_lo_p
  );


  buf

  (
    n2131_li166_li166,
    n966_lo_p
  );


  buf

  (
    n2134_li167_li167,
    n969_lo_p_spl_
  );


  buf

  (
    n2137_li168_li168,
    G43_p
  );


  buf

  (
    n2140_li169_li169,
    n975_lo_p
  );


  buf

  (
    n2143_li170_li170,
    n978_lo_p
  );


  buf

  (
    n2146_li171_li171,
    n981_lo_p_spl_
  );


  buf

  (
    n2149_li172_li172,
    G44_p
  );


  buf

  (
    n2152_li173_li173,
    n987_lo_p
  );


  buf

  (
    n2155_li174_li174,
    n990_lo_p
  );


  buf

  (
    n2158_li175_li175,
    n993_lo_p_spl_
  );


  buf

  (
    n2161_li176_li176,
    G45_p
  );


  buf

  (
    n2164_li177_li177,
    n999_lo_p
  );


  buf

  (
    n2170_li179_li179,
    lo178_buf_o2_p_spl_
  );


  buf

  (
    n2173_li180_li180,
    G46_p
  );


  buf

  (
    n2176_li181_li181,
    n1011_lo_p
  );


  buf

  (
    n2182_li183_li183,
    lo182_buf_o2_p_spl_
  );


  buf

  (
    n2185_li184_li184,
    G47_p
  );


  buf

  (
    n2194_li187_li187,
    lo186_buf_o2_p_spl_
  );


  buf

  (
    n2197_li188_li188,
    G48_p
  );


  buf

  (
    n2206_li191_li191,
    n1645_o2_p_spl_
  );


  buf

  (
    n2209_li192_li192,
    G49_p
  );


  buf

  (
    n2212_li193_li193,
    n1047_lo_p
  );


  buf

  (
    n2215_li194_li194,
    n1050_lo_p
  );


  buf

  (
    n2218_li195_li195,
    n1053_lo_p
  );


  buf

  (
    n2221_li196_li196,
    G50_p
  );


  buf

  (
    n2224_li197_li197,
    n1059_lo_p
  );


  buf

  (
    n2227_li198_li198,
    n1062_lo_p
  );


  buf

  (
    n2230_li199_li199,
    n1065_lo_p_spl_
  );


  buf

  (
    n2233_li200_li200,
    G51_p
  );


  buf

  (
    n2236_li201_li201,
    n1071_lo_p
  );


  buf

  (
    n2239_li202_li202,
    n1074_lo_p
  );


  buf

  (
    n2242_li203_li203,
    n1077_lo_p
  );


  buf

  (
    n2245_li204_li204,
    G52_p
  );


  buf

  (
    n2248_li205_li205,
    n1083_lo_p
  );


  buf

  (
    n2251_li206_li206,
    n1086_lo_p
  );


  buf

  (
    n2254_li207_li207,
    n1089_lo_p
  );


  buf

  (
    n2257_li208_li208,
    G53_p
  );


  buf

  (
    n2260_li209_li209,
    n1095_lo_p
  );


  buf

  (
    n2263_li210_li210,
    n1098_lo_p
  );


  buf

  (
    n2266_li211_li211,
    n1101_lo_p
  );


  buf

  (
    n2269_li212_li212,
    G54_p
  );


  buf

  (
    n2272_li213_li213,
    n1107_lo_p
  );


  buf

  (
    n2275_li214_li214,
    n1110_lo_p
  );


  buf

  (
    n2278_li215_li215,
    n1113_lo_p
  );


  buf

  (
    n2281_li216_li216,
    G55_p
  );


  buf

  (
    n2284_li217_li217,
    n1119_lo_p
  );


  buf

  (
    n2287_li218_li218,
    n1122_lo_p
  );


  buf

  (
    n2290_li219_li219,
    n1125_lo_p_spl_
  );


  buf

  (
    n2293_li220_li220,
    G56_p
  );


  buf

  (
    n2296_li221_li221,
    n1131_lo_p
  );


  buf

  (
    n2299_li222_li222,
    n1134_lo_p
  );


  buf

  (
    n2305_li224_li224,
    G57_p
  );


  buf

  (
    n2308_li225_li225,
    n1143_lo_p
  );


  buf

  (
    n2311_li226_li226,
    n1146_lo_p
  );


  buf

  (
    n2314_li227_li227,
    n1149_lo_p
  );


  buf

  (
    n2317_li228_li228,
    G58_p
  );


  buf

  (
    n2326_li231_li231,
    n1663_o2_p
  );


  buf

  (
    n2329_li232_li232,
    G59_p
  );


  buf

  (
    n2332_li233_li233,
    n1167_lo_p
  );


  buf

  (
    n2335_li234_li234,
    n1170_lo_p
  );


  buf

  (
    n2338_li235_li235,
    n1173_lo_p
  );


  buf

  (
    n2350_li239_li239,
    n1568_o2_p
  );


  buf

  (
    n1428_i2,
    n653_inv_p
  );


  buf

  (
    n1429_i2,
    n656_inv_p
  );


  buf

  (
    n1427_i2,
    n650_inv_p
  );


  buf

  (
    n1471_i2,
    n701_inv_p
  );


  buf

  (
    n1476_i2,
    n710_inv_p
  );


  buf

  (
    n1499_i2,
    n728_inv_p
  );


  buf

  (
    n1500_i2,
    n917_o2_p
  );


  buf

  (
    n1501_i2,
    n734_inv_p
  );


  buf

  (
    n1516_i2,
    n944_o2_p
  );


  buf

  (
    n1517_i2,
    n770_inv_p
  );


  buf

  (
    n1562_i2,
    n806_inv_p
  );


  buf

  (
    n1563_i2,
    n809_inv_p
  );


  buf

  (
    n1564_i2,
    n946_o2_p
  );


  buf

  (
    n1582_i2,
    n836_inv_p
  );


  buf

  (
    n1583_i2,
    n839_inv_p
  );


  buf

  (
    n1618_i2,
    n893_inv_p
  );


  buf

  (
    n1622_i2,
    n902_inv_p
  );


  buf

  (
    n1502_i2,
    n1649_o2_p
  );


  buf

  (
    n1503_i2,
    n1650_o2_p_spl_
  );


  buf

  (
    n1504_i2,
    n1651_o2_p
  );


  buf

  (
    n1505_i2,
    n1652_o2_p
  );


  buf

  (
    n1506_i2,
    n1653_o2_p
  );


  buf

  (
    n1512_i2,
    n1664_o2_p
  );


  buf

  (
    n1513_i2,
    n1665_o2_p
  );


  buf

  (
    n1514_i2,
    n1666_o2_p
  );


  buf

  (
    n1515_i2,
    n1667_o2_p
  );


  buf

  (
    n1644_i2,
    n917_inv_p
  );


  buf

  (
    n1647_i2,
    n926_inv_p
  );


  buf

  (
    n1527_i2,
    n1679_o2_p
  );


  buf

  (
    n1526_i2,
    n776_inv_p
  );


  buf

  (
    n1528_i2,
    n782_inv_p
  );


  buf

  (
    n1529_i2,
    n785_inv_p
  );


  buf

  (
    n1567_i2,
    lo038_buf_o2_p
  );


  not

  (
    n955_i2,
    g548_n_spl_
  );


  buf

  (
    n1568_i2,
    lo238_buf_o2_p_spl_
  );


  not

  (
    n1037_i2,
    g549_p_spl_
  );


  not

  (
    n960_i2,
    g550_n_spl_
  );


  buf

  (
    n1587_i2,
    lo122_buf_o2_p
  );


  not

  (
    n1040_i2,
    g551_p_spl_
  );


  not

  (
    n1039_i2,
    g552_p_spl_
  );


  buf

  (
    n1589_i2,
    n845_inv_p_spl_
  );


  buf

  (
    n1624_i2,
    lo146_buf_o2_p
  );


  buf

  (
    n1643_i2,
    lo118_buf_o2_p
  );


  not

  (
    n1038_i2,
    g553_n_spl_
  );


  buf

  (
    n1645_i2,
    lo190_buf_o2_p
  );


  not

  (
    n1029_i2,
    g558_p_spl_
  );


  buf

  (
    n1648_i2,
    n929_inv_p
  );


  buf

  (
    n1662_i2,
    lo142_buf_o2_p
  );


  buf

  (
    n1663_i2,
    lo230_buf_o2_p
  );


  buf

  (
    n1668_i2,
    n977_inv_p
  );


  not

  (
    n813_i2,
    g559_n_spl_
  );


  buf

  (
    lo114_buf_i2,
    lo113_buf_o2_p
  );


  not

  (
    n1031_i2,
    g560_p_spl_
  );


  buf

  (
    lo186_buf_i2,
    lo185_buf_o2_p
  );


  not

  (
    n1042_i2,
    g562_p_spl_
  );


  not

  (
    n911_i2,
    g563_n_spl_
  );


  not

  (
    n917_i2,
    g564_n_spl_
  );


  not

  (
    n942_i2,
    g565_p_spl_
  );


  buf

  (
    n1649_i2,
    lo002_buf_o2_p
  );


  buf

  (
    n1650_i2,
    lo014_buf_o2_p
  );


  buf

  (
    n1651_i2,
    lo030_buf_o2_p
  );


  buf

  (
    n1652_i2,
    lo034_buf_o2_p
  );


  buf

  (
    n1653_i2,
    lo042_buf_o2_p
  );


  buf

  (
    lo138_buf_i2,
    n882_lo_p_spl_
  );


  buf

  (
    n1664_i2,
    lo006_buf_o2_p
  );


  buf

  (
    n1665_i2,
    lo018_buf_o2_p
  );


  buf

  (
    n1666_i2,
    lo022_buf_o2_p
  );


  buf

  (
    n1667_i2,
    lo066_buf_o2_p
  );


  not

  (
    n944_i2,
    g566_p_spl_
  );


  not

  (
    n945_i2,
    g567_p_spl_
  );


  buf

  (
    n1672_i2,
    n892_o2_p_spl_
  );


  buf

  (
    n1676_i2,
    n995_inv_p
  );


  buf

  (
    n1679_i2,
    lo062_buf_o2_p_spl_
  );


  buf

  (
    n1680_i2,
    n1007_inv_p_spl_1
  );


  buf

  (
    n1681_i2,
    n1010_inv_p_spl_
  );


  buf

  (
    lo110_buf_i2,
    n798_lo_p_spl_
  );


  buf

  (
    lo134_buf_i2,
    n870_lo_p_spl_
  );


  not

  (
    n1030_i2,
    g568_n_spl_
  );


  buf

  (
    lo182_buf_i2,
    n1014_lo_p
  );


  not

  (
    n830_i2,
    g571_n_spl_
  );


  buf

  (
    n1021_i2,
    g577_n_spl_
  );


  not

  (
    n943_i2,
    g578_n_spl_
  );


  not

  (
    n936_i2,
    g582_p_spl_
  );


  not

  (
    n946_i2,
    g583_n_spl_
  );


  buf

  (
    lo038_buf_i2,
    lo037_buf_o2_p_spl_
  );


  buf

  (
    lo238_buf_i2,
    lo237_buf_o2_p
  );


  not

  (
    n1010_i2,
    g585_n_spl_
  );


  not

  (
    n1006_i2,
    g587_n_spl_
  );


  not

  (
    n907_i2,
    g589_n_spl_
  );


  buf

  (
    n902_i2,
    g591_p_spl_
  );


  buf

  (
    lo154_buf_i2,
    lo152_buf_o2_p_spl_
  );


  not

  (
    n938_i2,
    g592_n_spl_
  );


  not

  (
    n947_i2,
    g593_p_spl_
  );


  buf

  (
    lo122_buf_i2,
    n831_lo_p_spl_
  );


  buf

  (
    n899_i2,
    g599_n_spl_
  );


  buf

  (
    n904_i2,
    g601_p_spl_
  );


  buf

  (
    lo106_buf_i2,
    n786_lo_p_spl_
  );


  buf

  (
    n980_i2,
    g602_p
  );


  buf

  (
    n1023_i2,
    g603_p
  );


  buf

  (
    lo178_buf_i2,
    n1002_lo_p_spl_
  );


  buf

  (
    n981_i2,
    g604_p
  );


  buf

  (
    n837_i2,
    g607_p
  );


  buf

  (
    n1013_i2,
    g613_n
  );


  buf

  (
    n840_i2,
    g616_p
  );


  buf

  (
    n849_i2,
    g619_p
  );


  buf

  (
    n852_i2,
    g622_p
  );


  buf

  (
    n864_i2,
    g625_p
  );


  buf

  (
    n867_i2,
    g628_p
  );


  not

  (
    n1044_i2,
    g630_p
  );


  buf

  (
    n876_i2,
    g633_p
  );


  not

  (
    n937_i2,
    g634_p_spl_
  );


  buf

  (
    n879_i2,
    g637_p
  );


  not

  (
    n925_i2,
    g640_n
  );


  buf

  (
    n954_i2,
    g644_n_spl_
  );


  buf

  (
    lo146_buf_i2,
    n903_lo_p_spl_
  );


  buf

  (
    n1026_i2,
    g645_p
  );


  buf

  (
    n1032_i2,
    g646_p
  );


  buf

  (
    lo118_buf_i2,
    n819_lo_p_spl_
  );


  buf

  (
    n957_i2,
    g647_n
  );


  buf

  (
    lo190_buf_i2,
    n1035_lo_p_spl_
  );


  not

  (
    n1036_i2,
    g651_p
  );


  not

  (
    n949_i2,
    g653_n
  );


  buf

  (
    n910_i2,
    g657_n_spl_
  );


  buf

  (
    lo002_buf_i2,
    G1_p
  );


  buf

  (
    lo014_buf_i2,
    G4_p_spl_1
  );


  buf

  (
    lo030_buf_i2,
    G8_p_spl_
  );


  buf

  (
    lo034_buf_i2,
    G9_p
  );


  buf

  (
    lo042_buf_i2,
    G11_p_spl_
  );


  buf

  (
    lo113_buf_i2,
    n807_lo_p
  );


  buf

  (
    lo185_buf_i2,
    n1023_lo_p
  );


  buf

  (
    n939_i2,
    g658_p
  );


  buf

  (
    n941_i2,
    g660_n
  );


  buf

  (
    lo142_buf_i2,
    n891_lo_p
  );


  buf

  (
    lo230_buf_i2,
    n1155_lo_p
  );


  buf

  (
    lo006_buf_i2,
    G2_p_spl_
  );


  buf

  (
    lo018_buf_i2,
    G5_p
  );


  buf

  (
    lo022_buf_i2,
    G6_p_spl_
  );


  buf

  (
    lo066_buf_i2,
    G17_p_spl_
  );


  buf

  (
    n913_i2,
    g661_n
  );


  not

  (
    n826_i2,
    g662_n_spl_
  );


  not

  (
    n892_i2,
    g663_n_spl_
  );


  buf

  (
    lo152_buf_i2,
    G39_p
  );


  buf

  (
    n896_i2,
    g664_p
  );


  buf

  (
    n905_i2,
    g665_p
  );


  buf

  (
    n821_i2,
    g666_p
  );


  buf

  (
    lo037_buf_i2,
    G10_p
  );


  buf

  (
    lo237_buf_i2,
    G60_p
  );


  buf

  (
    lo062_buf_i2,
    G16_p
  );


  not

  (
    n827_i2,
    g667_n
  );


  buf

  (
    n809_i2,
    g668_p
  );


  buf

  (
    n891_i2,
    g671_n
  );


  buf

  (
    n540_lo_n_spl_,
    n540_lo_n
  );


  buf

  (
    n660_lo_n_spl_,
    n660_lo_n
  );


  buf

  (
    g370_n_spl_,
    g370_n
  );


  buf

  (
    n552_lo_n_spl_,
    n552_lo_n
  );


  buf

  (
    n552_lo_n_spl_0,
    n552_lo_n_spl_
  );


  buf

  (
    n552_lo_p_spl_,
    n552_lo_p
  );


  buf

  (
    g375_n_spl_,
    g375_n
  );


  buf

  (
    g377_n_spl_,
    g377_n
  );


  buf

  (
    n600_lo_n_spl_,
    n600_lo_n
  );


  buf

  (
    g379_n_spl_,
    g379_n
  );


  buf

  (
    g383_n_spl_,
    g383_n
  );


  buf

  (
    g373_n_spl_,
    g373_n
  );


  buf

  (
    n830_o2_n_spl_,
    n830_o2_n
  );


  buf

  (
    n837_o2_n_spl_,
    n837_o2_n
  );


  buf

  (
    n840_o2_n_spl_,
    n840_o2_n
  );


  buf

  (
    n837_o2_p_spl_,
    n837_o2_p
  );


  buf

  (
    n840_o2_p_spl_,
    n840_o2_p
  );


  buf

  (
    n852_lo_p_spl_,
    n852_lo_p
  );


  buf

  (
    n852_lo_p_spl_0,
    n852_lo_p_spl_
  );


  buf

  (
    n852_lo_p_spl_1,
    n852_lo_p_spl_
  );


  buf

  (
    g392_p_spl_,
    g392_p
  );


  buf

  (
    n852_lo_n_spl_,
    n852_lo_n
  );


  buf

  (
    n852_lo_n_spl_0,
    n852_lo_n_spl_
  );


  buf

  (
    n852_lo_n_spl_1,
    n852_lo_n_spl_
  );


  buf

  (
    g392_n_spl_,
    g392_n
  );


  buf

  (
    n849_o2_n_spl_,
    n849_o2_n
  );


  buf

  (
    n852_o2_n_spl_,
    n852_o2_n
  );


  buf

  (
    n849_o2_p_spl_,
    n849_o2_p
  );


  buf

  (
    n852_o2_p_spl_,
    n852_o2_p
  );


  buf

  (
    n864_lo_p_spl_,
    n864_lo_p
  );


  buf

  (
    g398_p_spl_,
    g398_p
  );


  buf

  (
    n864_lo_n_spl_,
    n864_lo_n
  );


  buf

  (
    g398_n_spl_,
    g398_n
  );


  buf

  (
    n864_o2_n_spl_,
    n864_o2_n
  );


  buf

  (
    n867_o2_n_spl_,
    n867_o2_n
  );


  buf

  (
    n864_o2_p_spl_,
    n864_o2_p
  );


  buf

  (
    n867_o2_p_spl_,
    n867_o2_p
  );


  buf

  (
    g407_p_spl_,
    g407_p
  );


  buf

  (
    g407_n_spl_,
    g407_n
  );


  buf

  (
    n876_o2_n_spl_,
    n876_o2_n
  );


  buf

  (
    n879_o2_n_spl_,
    n879_o2_n
  );


  buf

  (
    n876_o2_p_spl_,
    n876_o2_p
  );


  buf

  (
    n879_o2_p_spl_,
    n879_o2_p
  );


  buf

  (
    n1056_lo_p_spl_,
    n1056_lo_p
  );


  buf

  (
    g413_p_spl_,
    g413_p
  );


  buf

  (
    n1056_lo_n_spl_,
    n1056_lo_n
  );


  buf

  (
    g413_n_spl_,
    g413_n
  );


  buf

  (
    n1104_lo_n_spl_,
    n1104_lo_n
  );


  buf

  (
    n1104_lo_n_spl_0,
    n1104_lo_n_spl_
  );


  buf

  (
    n1104_lo_n_spl_00,
    n1104_lo_n_spl_0
  );


  buf

  (
    n1104_lo_n_spl_01,
    n1104_lo_n_spl_0
  );


  buf

  (
    n1104_lo_n_spl_1,
    n1104_lo_n_spl_
  );


  buf

  (
    n1104_lo_n_spl_10,
    n1104_lo_n_spl_1
  );


  buf

  (
    n1104_lo_n_spl_11,
    n1104_lo_n_spl_1
  );


  buf

  (
    n1080_lo_n_spl_,
    n1080_lo_n
  );


  buf

  (
    n1080_lo_n_spl_0,
    n1080_lo_n_spl_
  );


  buf

  (
    n1080_lo_n_spl_00,
    n1080_lo_n_spl_0
  );


  buf

  (
    n1080_lo_n_spl_000,
    n1080_lo_n_spl_00
  );


  buf

  (
    n1080_lo_n_spl_001,
    n1080_lo_n_spl_00
  );


  buf

  (
    n1080_lo_n_spl_01,
    n1080_lo_n_spl_0
  );


  buf

  (
    n1080_lo_n_spl_010,
    n1080_lo_n_spl_01
  );


  buf

  (
    n1080_lo_n_spl_1,
    n1080_lo_n_spl_
  );


  buf

  (
    n1080_lo_n_spl_10,
    n1080_lo_n_spl_1
  );


  buf

  (
    n1080_lo_n_spl_11,
    n1080_lo_n_spl_1
  );


  buf

  (
    n1092_lo_n_spl_,
    n1092_lo_n
  );


  buf

  (
    n1092_lo_n_spl_0,
    n1092_lo_n_spl_
  );


  buf

  (
    n1092_lo_n_spl_00,
    n1092_lo_n_spl_0
  );


  buf

  (
    n1092_lo_n_spl_01,
    n1092_lo_n_spl_0
  );


  buf

  (
    n1092_lo_n_spl_1,
    n1092_lo_n_spl_
  );


  buf

  (
    n1092_lo_n_spl_10,
    n1092_lo_n_spl_1
  );


  buf

  (
    n1092_lo_n_spl_11,
    n1092_lo_n_spl_1
  );


  buf

  (
    n1116_lo_n_spl_,
    n1116_lo_n
  );


  buf

  (
    n1116_lo_n_spl_0,
    n1116_lo_n_spl_
  );


  buf

  (
    n1116_lo_n_spl_00,
    n1116_lo_n_spl_0
  );


  buf

  (
    n1116_lo_n_spl_01,
    n1116_lo_n_spl_0
  );


  buf

  (
    n1116_lo_n_spl_1,
    n1116_lo_n_spl_
  );


  buf

  (
    n1116_lo_n_spl_10,
    n1116_lo_n_spl_1
  );


  buf

  (
    n1116_lo_n_spl_11,
    n1116_lo_n_spl_1
  );


  buf

  (
    n925_o2_n_spl_,
    n925_o2_n
  );


  buf

  (
    n925_o2_n_spl_0,
    n925_o2_n_spl_
  );


  buf

  (
    n925_o2_n_spl_00,
    n925_o2_n_spl_0
  );


  buf

  (
    n925_o2_n_spl_01,
    n925_o2_n_spl_0
  );


  buf

  (
    n925_o2_n_spl_1,
    n925_o2_n_spl_
  );


  buf

  (
    n925_o2_n_spl_10,
    n925_o2_n_spl_1
  );


  buf

  (
    n925_o2_n_spl_11,
    n925_o2_n_spl_1
  );


  buf

  (
    n1068_lo_n_spl_,
    n1068_lo_n
  );


  buf

  (
    n1068_lo_n_spl_0,
    n1068_lo_n_spl_
  );


  buf

  (
    n1068_lo_n_spl_00,
    n1068_lo_n_spl_0
  );


  buf

  (
    n1068_lo_n_spl_01,
    n1068_lo_n_spl_0
  );


  buf

  (
    n1068_lo_n_spl_1,
    n1068_lo_n_spl_
  );


  buf

  (
    n1068_lo_n_spl_10,
    n1068_lo_n_spl_1
  );


  buf

  (
    n1128_lo_n_spl_,
    n1128_lo_n
  );


  buf

  (
    n1582_o2_n_spl_,
    n1582_o2_n
  );


  buf

  (
    g450_n_spl_,
    g450_n
  );


  buf

  (
    n960_lo_p_spl_,
    n960_lo_p
  );


  buf

  (
    n1013_o2_p_spl_,
    n1013_o2_p
  );


  buf

  (
    n960_lo_n_spl_,
    n960_lo_n
  );


  buf

  (
    n960_lo_n_spl_0,
    n960_lo_n_spl_
  );


  buf

  (
    n1013_o2_n_spl_,
    n1013_o2_n
  );


  buf

  (
    n1013_o2_n_spl_0,
    n1013_o2_n_spl_
  );


  buf

  (
    n972_lo_n_spl_,
    n972_lo_n
  );


  buf

  (
    n1021_o2_n_spl_,
    n1021_o2_n
  );


  buf

  (
    n1023_o2_n_spl_,
    n1023_o2_n
  );


  buf

  (
    n1023_o2_n_spl_0,
    n1023_o2_n_spl_
  );


  buf

  (
    n1044_o2_n_spl_,
    n1044_o2_n
  );


  buf

  (
    n1023_o2_p_spl_,
    n1023_o2_p
  );


  buf

  (
    n1044_o2_p_spl_,
    n1044_o2_p
  );


  buf

  (
    g483_n_spl_,
    g483_n
  );


  buf

  (
    g483_p_spl_,
    g483_p
  );


  buf

  (
    g482_p_spl_,
    g482_p
  );


  buf

  (
    g485_n_spl_,
    g485_n
  );


  buf

  (
    g481_n_spl_,
    g481_n
  );


  buf

  (
    g481_n_spl_0,
    g481_n_spl_
  );


  buf

  (
    n1038_o2_n_spl_,
    n1038_o2_n
  );


  buf

  (
    g488_n_spl_,
    g488_n
  );


  buf

  (
    g503_n_spl_,
    g503_n
  );


  buf

  (
    g518_n_spl_,
    g518_n
  );


  buf

  (
    n1030_o2_n_spl_,
    n1030_o2_n
  );


  buf

  (
    g533_n_spl_,
    g533_n
  );


  buf

  (
    lo178_buf_o2_n_spl_,
    lo178_buf_o2_n
  );


  buf

  (
    n993_lo_n_spl_,
    n993_lo_n
  );


  buf

  (
    n993_lo_n_spl_0,
    n993_lo_n_spl_
  );


  buf

  (
    g549_p_spl_,
    g549_p
  );


  buf

  (
    g549_p_spl_0,
    g549_p_spl_
  );


  buf

  (
    g548_n_spl_,
    g548_n
  );


  buf

  (
    g550_n_spl_,
    g550_n
  );


  buf

  (
    n777_lo_n_spl_,
    n777_lo_n
  );


  buf

  (
    n981_lo_n_spl_,
    n981_lo_n
  );


  buf

  (
    n981_lo_n_spl_0,
    n981_lo_n_spl_
  );


  buf

  (
    g558_p_spl_,
    g558_p
  );


  buf

  (
    g558_p_spl_0,
    g558_p_spl_
  );


  buf

  (
    g551_p_spl_,
    g551_p
  );


  buf

  (
    g552_p_spl_,
    g552_p
  );


  buf

  (
    g553_n_spl_,
    g553_n
  );


  buf

  (
    lo185_buf_o2_n_spl_,
    lo185_buf_o2_n
  );


  buf

  (
    g565_p_spl_,
    g565_p
  );


  buf

  (
    g565_p_spl_0,
    g565_p_spl_
  );


  buf

  (
    g563_n_spl_,
    g563_n
  );


  buf

  (
    g564_n_spl_,
    g564_n
  );


  buf

  (
    g559_n_spl_,
    g559_n
  );


  buf

  (
    n765_lo_p_spl_,
    n765_lo_p
  );


  buf

  (
    n765_lo_p_spl_0,
    n765_lo_p_spl_
  );


  buf

  (
    n1589_o2_p_spl_,
    n1589_o2_p
  );


  buf

  (
    n1010_o2_p_spl_,
    n1010_o2_p
  );


  buf

  (
    lo134_buf_o2_p_spl_,
    lo134_buf_o2_p
  );


  buf

  (
    n1006_o2_p_spl_,
    n1006_o2_p
  );


  buf

  (
    g566_p_spl_,
    g566_p
  );


  buf

  (
    g567_p_spl_,
    g567_p
  );


  buf

  (
    lo238_buf_o2_p_spl_,
    lo238_buf_o2_p
  );


  buf

  (
    n1007_inv_p_spl_,
    n1007_inv_p
  );


  buf

  (
    n1007_inv_p_spl_0,
    n1007_inv_p_spl_
  );


  buf

  (
    n1007_inv_p_spl_1,
    n1007_inv_p_spl_
  );


  buf

  (
    lo062_buf_o2_p_spl_,
    lo062_buf_o2_p
  );


  buf

  (
    n1010_inv_p_spl_,
    n1010_inv_p
  );


  buf

  (
    n1014_lo_n_spl_,
    n1014_lo_n
  );


  buf

  (
    g582_p_spl_,
    g582_p
  );


  buf

  (
    g582_p_spl_0,
    g582_p_spl_
  );


  buf

  (
    g578_n_spl_,
    g578_n
  );


  buf

  (
    g583_n_spl_,
    g583_n
  );


  buf

  (
    n892_o2_p_spl_,
    n892_o2_p
  );


  buf

  (
    lo037_buf_o2_p_spl_,
    lo037_buf_o2_p
  );


  buf

  (
    g591_p_spl_,
    g591_p
  );


  buf

  (
    n1065_lo_p_spl_,
    n1065_lo_p
  );


  buf

  (
    lo110_buf_o2_p_spl_,
    lo110_buf_o2_p
  );


  buf

  (
    n969_lo_p_spl_,
    n969_lo_p
  );


  buf

  (
    n969_lo_p_spl_0,
    n969_lo_p_spl_
  );


  buf

  (
    g577_n_spl_,
    g577_n
  );


  buf

  (
    n1125_lo_p_spl_,
    n1125_lo_p
  );


  buf

  (
    n753_lo_p_spl_,
    n753_lo_p
  );


  buf

  (
    n753_lo_p_spl_0,
    n753_lo_p_spl_
  );


  buf

  (
    n1512_o2_p_spl_,
    n1512_o2_p
  );


  buf

  (
    n777_lo_p_spl_,
    n777_lo_p
  );


  buf

  (
    lo106_buf_o2_p_spl_,
    lo106_buf_o2_p
  );


  buf

  (
    lo114_buf_o2_p_spl_,
    lo114_buf_o2_p
  );


  buf

  (
    n1643_o2_p_spl_,
    n1643_o2_p
  );


  buf

  (
    n957_lo_p_spl_,
    n957_lo_p
  );


  buf

  (
    n981_lo_p_spl_,
    n981_lo_p
  );


  buf

  (
    n993_lo_p_spl_,
    n993_lo_p
  );


  buf

  (
    g560_p_spl_,
    g560_p
  );


  buf

  (
    g562_p_spl_,
    g562_p
  );


  buf

  (
    g568_n_spl_,
    g568_n
  );


  buf

  (
    lo182_buf_o2_p_spl_,
    lo182_buf_o2_p
  );


  buf

  (
    lo178_buf_o2_p_spl_,
    lo178_buf_o2_p
  );


  buf

  (
    n1645_o2_p_spl_,
    n1645_o2_p
  );


  buf

  (
    lo186_buf_o2_p_spl_,
    lo186_buf_o2_p
  );


  buf

  (
    g571_n_spl_,
    g571_n
  );


  buf

  (
    n798_lo_p_spl_,
    n798_lo_p
  );


  buf

  (
    n845_inv_p_spl_,
    n845_inv_p
  );


  buf

  (
    n845_inv_p_spl_0,
    n845_inv_p_spl_
  );


  buf

  (
    n882_lo_p_spl_,
    n882_lo_p
  );


  buf

  (
    n870_lo_p_spl_,
    n870_lo_p
  );


  buf

  (
    n1650_o2_p_spl_,
    n1650_o2_p
  );


  buf

  (
    n786_lo_p_spl_,
    n786_lo_p
  );


  buf

  (
    n1002_lo_p_spl_,
    n1002_lo_p
  );


  buf

  (
    g644_n_spl_,
    g644_n
  );


  buf

  (
    g585_n_spl_,
    g585_n
  );


  buf

  (
    g587_n_spl_,
    g587_n
  );


  buf

  (
    g592_n_spl_,
    g592_n
  );


  buf

  (
    g593_p_spl_,
    g593_p
  );


  buf

  (
    g634_p_spl_,
    g634_p
  );


  buf

  (
    n831_lo_p_spl_,
    n831_lo_p
  );


  buf

  (
    g599_n_spl_,
    g599_n
  );


  buf

  (
    g599_n_spl_0,
    g599_n_spl_
  );


  buf

  (
    lo152_buf_o2_p_spl_,
    lo152_buf_o2_p
  );


  buf

  (
    g589_n_spl_,
    g589_n
  );


  buf

  (
    g589_n_spl_0,
    g589_n_spl_
  );


  buf

  (
    g601_p_spl_,
    g601_p
  );


  buf

  (
    g601_p_spl_0,
    g601_p_spl_
  );


  buf

  (
    n819_lo_p_spl_,
    n819_lo_p
  );


  buf

  (
    n903_lo_p_spl_,
    n903_lo_p
  );


  buf

  (
    n1035_lo_p_spl_,
    n1035_lo_p
  );


  buf

  (
    g657_n_spl_,
    g657_n
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    g663_n_spl_,
    g663_n
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    g662_n_spl_,
    g662_n
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


endmodule
