
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  G42,
  G43,
  G44,
  G45,
  G46,
  G47,
  G48,
  G49,
  G50,
  G51,
  G52,
  G53,
  G54,
  G55,
  G56,
  G57,
  G58,
  G59,
  G60,
  G61,
  G62,
  G63,
  G64,
  G65,
  G66,
  G67,
  G68,
  G69,
  G70,
  G71,
  G72,
  G73,
  G74,
  G75,
  G76,
  G77,
  G78,
  G79,
  G80,
  G81,
  G82,
  G83,
  G84,
  G85,
  G86,
  G87,
  G88,
  G89,
  G90,
  G91,
  G92,
  G93,
  G94,
  G95,
  G96,
  G97,
  G98,
  G99,
  G100,
  G101,
  G102,
  G103,
  G104,
  G105,
  G106,
  G107,
  G108,
  G109,
  G110,
  G111,
  G112,
  G113,
  G114,
  G115,
  G116,
  G117,
  G118,
  G119,
  G120,
  G121,
  G122,
  G123,
  G124,
  G125,
  G126,
  G127,
  G128,
  G129,
  G130,
  G131,
  G132,
  G133,
  G134,
  G135,
  G136,
  G137,
  G138,
  G139,
  G140,
  G141,
  G142,
  G143,
  G144,
  G145,
  G146,
  G147,
  G148,
  G149,
  G150,
  G151,
  G152,
  G153,
  G154,
  G155,
  G156,
  G157,
  G158,
  G159,
  G160,
  G161,
  G162,
  G163,
  G164,
  G165,
  G166,
  G167,
  G168,
  G169,
  G170,
  G171,
  G172,
  G173,
  G174,
  G175,
  G176,
  G177,
  G178,
  G5193,
  G5194,
  G5195,
  G5196,
  G5197,
  G5198,
  G5199,
  G5200,
  G5201,
  G5202,
  G5203,
  G5204,
  G5205,
  G5206,
  G5207,
  G5208,
  G5209,
  G5210,
  G5211,
  G5212,
  G5213,
  G5214,
  G5215,
  G5216,
  G5217,
  G5218,
  G5219,
  G5220,
  G5221,
  G5222,
  G5223,
  G5224,
  G5225,
  G5226,
  G5227,
  G5228,
  G5229,
  G5230,
  G5231,
  G5232,
  G5233,
  G5234,
  G5235,
  G5236,
  G5237,
  G5238,
  G5239,
  G5240,
  G5241,
  G5242,
  G5243,
  G5244,
  G5245,
  G5246,
  G5247,
  G5248,
  G5249,
  G5250,
  G5251,
  G5252,
  G5253,
  G5254,
  G5255,
  G5256,
  G5257,
  G5258,
  G5259,
  G5260,
  G5261,
  G5262,
  G5263,
  G5264,
  G5265,
  G5266,
  G5267,
  G5268,
  G5269,
  G5270,
  G5271,
  G5272,
  G5273,
  G5274,
  G5275,
  G5276,
  G5277,
  G5278,
  G5279,
  G5280,
  G5281,
  G5282,
  G5283,
  G5284,
  G5285,
  G5286,
  G5287,
  G5288,
  G5289,
  G5290,
  G5291,
  G5292,
  G5293,
  G5294,
  G5295,
  G5296,
  G5297,
  G5298,
  G5299,
  G5300,
  G5301,
  G5302,
  G5303,
  G5304,
  G5305,
  G5306,
  G5307,
  G5308,
  G5309,
  G5310,
  G5311,
  G5312,
  G5313,
  G5314,
  G5315
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input G42;input G43;input G44;input G45;input G46;input G47;input G48;input G49;input G50;input G51;input G52;input G53;input G54;input G55;input G56;input G57;input G58;input G59;input G60;input G61;input G62;input G63;input G64;input G65;input G66;input G67;input G68;input G69;input G70;input G71;input G72;input G73;input G74;input G75;input G76;input G77;input G78;input G79;input G80;input G81;input G82;input G83;input G84;input G85;input G86;input G87;input G88;input G89;input G90;input G91;input G92;input G93;input G94;input G95;input G96;input G97;input G98;input G99;input G100;input G101;input G102;input G103;input G104;input G105;input G106;input G107;input G108;input G109;input G110;input G111;input G112;input G113;input G114;input G115;input G116;input G117;input G118;input G119;input G120;input G121;input G122;input G123;input G124;input G125;input G126;input G127;input G128;input G129;input G130;input G131;input G132;input G133;input G134;input G135;input G136;input G137;input G138;input G139;input G140;input G141;input G142;input G143;input G144;input G145;input G146;input G147;input G148;input G149;input G150;input G151;input G152;input G153;input G154;input G155;input G156;input G157;input G158;input G159;input G160;input G161;input G162;input G163;input G164;input G165;input G166;input G167;input G168;input G169;input G170;input G171;input G172;input G173;input G174;input G175;input G176;input G177;input G178;
  output G5193;output G5194;output G5195;output G5196;output G5197;output G5198;output G5199;output G5200;output G5201;output G5202;output G5203;output G5204;output G5205;output G5206;output G5207;output G5208;output G5209;output G5210;output G5211;output G5212;output G5213;output G5214;output G5215;output G5216;output G5217;output G5218;output G5219;output G5220;output G5221;output G5222;output G5223;output G5224;output G5225;output G5226;output G5227;output G5228;output G5229;output G5230;output G5231;output G5232;output G5233;output G5234;output G5235;output G5236;output G5237;output G5238;output G5239;output G5240;output G5241;output G5242;output G5243;output G5244;output G5245;output G5246;output G5247;output G5248;output G5249;output G5250;output G5251;output G5252;output G5253;output G5254;output G5255;output G5256;output G5257;output G5258;output G5259;output G5260;output G5261;output G5262;output G5263;output G5264;output G5265;output G5266;output G5267;output G5268;output G5269;output G5270;output G5271;output G5272;output G5273;output G5274;output G5275;output G5276;output G5277;output G5278;output G5279;output G5280;output G5281;output G5282;output G5283;output G5284;output G5285;output G5286;output G5287;output G5288;output G5289;output G5290;output G5291;output G5292;output G5293;output G5294;output G5295;output G5296;output G5297;output G5298;output G5299;output G5300;output G5301;output G5302;output G5303;output G5304;output G5305;output G5306;output G5307;output G5308;output G5309;output G5310;output G5311;output G5312;output G5313;output G5314;output G5315;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire G51_p;
  wire G51_n;
  wire G52_p;
  wire G52_n;
  wire G53_p;
  wire G53_n;
  wire G54_p;
  wire G54_n;
  wire G55_p;
  wire G55_n;
  wire G56_p;
  wire G56_n;
  wire G57_p;
  wire G57_n;
  wire G58_p;
  wire G58_n;
  wire G59_p;
  wire G59_n;
  wire G60_p;
  wire G60_n;
  wire G61_p;
  wire G61_n;
  wire G62_p;
  wire G62_n;
  wire G63_p;
  wire G63_n;
  wire G64_p;
  wire G64_n;
  wire G65_p;
  wire G65_n;
  wire G66_p;
  wire G66_n;
  wire G67_p;
  wire G67_n;
  wire G68_p;
  wire G68_n;
  wire G69_p;
  wire G69_n;
  wire G70_p;
  wire G70_n;
  wire G71_p;
  wire G71_n;
  wire G72_p;
  wire G72_n;
  wire G73_p;
  wire G73_n;
  wire G74_p;
  wire G74_n;
  wire G75_p;
  wire G75_n;
  wire G76_p;
  wire G76_n;
  wire G77_p;
  wire G77_n;
  wire G78_p;
  wire G78_n;
  wire G79_p;
  wire G79_n;
  wire G80_p;
  wire G80_n;
  wire G81_p;
  wire G81_n;
  wire G82_p;
  wire G82_n;
  wire G83_p;
  wire G83_n;
  wire G84_p;
  wire G84_n;
  wire G85_p;
  wire G85_n;
  wire G86_p;
  wire G86_n;
  wire G87_p;
  wire G87_n;
  wire G88_p;
  wire G88_n;
  wire G89_p;
  wire G89_n;
  wire G90_p;
  wire G90_n;
  wire G91_p;
  wire G91_n;
  wire G92_p;
  wire G92_n;
  wire G93_p;
  wire G93_n;
  wire G94_p;
  wire G94_n;
  wire G95_p;
  wire G95_n;
  wire G96_p;
  wire G96_n;
  wire G97_p;
  wire G97_n;
  wire G98_p;
  wire G98_n;
  wire G99_p;
  wire G99_n;
  wire G100_p;
  wire G100_n;
  wire G101_p;
  wire G101_n;
  wire G102_p;
  wire G102_n;
  wire G103_p;
  wire G103_n;
  wire G104_p;
  wire G104_n;
  wire G105_p;
  wire G105_n;
  wire G106_p;
  wire G106_n;
  wire G107_p;
  wire G107_n;
  wire G108_p;
  wire G108_n;
  wire G109_p;
  wire G109_n;
  wire G110_p;
  wire G110_n;
  wire G111_p;
  wire G111_n;
  wire G112_p;
  wire G112_n;
  wire G113_p;
  wire G113_n;
  wire G114_p;
  wire G114_n;
  wire G115_p;
  wire G115_n;
  wire G116_p;
  wire G116_n;
  wire G117_p;
  wire G117_n;
  wire G118_p;
  wire G118_n;
  wire G119_p;
  wire G119_n;
  wire G120_p;
  wire G120_n;
  wire G121_p;
  wire G121_n;
  wire G122_p;
  wire G122_n;
  wire G123_p;
  wire G123_n;
  wire G124_p;
  wire G124_n;
  wire G125_p;
  wire G125_n;
  wire G126_p;
  wire G126_n;
  wire G127_p;
  wire G127_n;
  wire G128_p;
  wire G128_n;
  wire G129_p;
  wire G129_n;
  wire G130_p;
  wire G130_n;
  wire G131_p;
  wire G131_n;
  wire G132_p;
  wire G132_n;
  wire G133_p;
  wire G133_n;
  wire G134_p;
  wire G134_n;
  wire G135_p;
  wire G135_n;
  wire G136_p;
  wire G136_n;
  wire G137_p;
  wire G137_n;
  wire G138_p;
  wire G138_n;
  wire G139_p;
  wire G139_n;
  wire G140_p;
  wire G140_n;
  wire G141_p;
  wire G141_n;
  wire G142_p;
  wire G142_n;
  wire G143_p;
  wire G143_n;
  wire G144_p;
  wire G144_n;
  wire G145_p;
  wire G145_n;
  wire G146_p;
  wire G146_n;
  wire G147_p;
  wire G147_n;
  wire G148_p;
  wire G148_n;
  wire G149_p;
  wire G149_n;
  wire G150_p;
  wire G150_n;
  wire G151_p;
  wire G151_n;
  wire G152_p;
  wire G152_n;
  wire G153_p;
  wire G153_n;
  wire G154_p;
  wire G154_n;
  wire G155_p;
  wire G155_n;
  wire G156_p;
  wire G156_n;
  wire G157_p;
  wire G157_n;
  wire G158_p;
  wire G158_n;
  wire G159_p;
  wire G159_n;
  wire G160_p;
  wire G160_n;
  wire G161_p;
  wire G161_n;
  wire G162_p;
  wire G162_n;
  wire G163_p;
  wire G163_n;
  wire G164_p;
  wire G164_n;
  wire G165_p;
  wire G165_n;
  wire G166_p;
  wire G166_n;
  wire G167_p;
  wire G167_n;
  wire G168_p;
  wire G168_n;
  wire G169_p;
  wire G169_n;
  wire G170_p;
  wire G170_n;
  wire G171_p;
  wire G171_n;
  wire G172_p;
  wire G172_n;
  wire G173_p;
  wire G173_n;
  wire G174_p;
  wire G174_n;
  wire G175_p;
  wire G175_n;
  wire G176_p;
  wire G176_n;
  wire G177_p;
  wire G177_n;
  wire G178_p;
  wire G178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire g693_p;
  wire g693_n;
  wire g694_p;
  wire g694_n;
  wire g695_p;
  wire g695_n;
  wire g696_p;
  wire g696_n;
  wire g697_p;
  wire g697_n;
  wire g698_p;
  wire g698_n;
  wire g699_p;
  wire g699_n;
  wire g700_p;
  wire g700_n;
  wire g701_p;
  wire g701_n;
  wire g702_p;
  wire g702_n;
  wire g703_p;
  wire g703_n;
  wire g704_p;
  wire g704_n;
  wire g705_p;
  wire g705_n;
  wire g706_p;
  wire g706_n;
  wire g707_p;
  wire g707_n;
  wire g708_p;
  wire g708_n;
  wire g709_p;
  wire g709_n;
  wire g710_p;
  wire g710_n;
  wire g711_p;
  wire g711_n;
  wire g712_p;
  wire g712_n;
  wire g713_p;
  wire g713_n;
  wire g714_p;
  wire g714_n;
  wire g715_p;
  wire g715_n;
  wire g716_p;
  wire g716_n;
  wire g717_p;
  wire g717_n;
  wire g718_p;
  wire g718_n;
  wire g719_p;
  wire g719_n;
  wire g720_p;
  wire g720_n;
  wire g721_p;
  wire g721_n;
  wire g722_p;
  wire g722_n;
  wire g723_p;
  wire g723_n;
  wire g724_p;
  wire g724_n;
  wire g725_p;
  wire g725_n;
  wire g726_p;
  wire g726_n;
  wire g727_p;
  wire g727_n;
  wire g728_p;
  wire g728_n;
  wire g729_p;
  wire g729_n;
  wire g730_p;
  wire g730_n;
  wire g731_p;
  wire g731_n;
  wire g732_p;
  wire g732_n;
  wire g733_p;
  wire g733_n;
  wire g734_p;
  wire g734_n;
  wire g735_p;
  wire g735_n;
  wire g736_p;
  wire g736_n;
  wire g737_p;
  wire g737_n;
  wire g738_p;
  wire g738_n;
  wire g739_p;
  wire g739_n;
  wire g740_p;
  wire g740_n;
  wire g741_p;
  wire g741_n;
  wire g742_p;
  wire g742_n;
  wire g743_p;
  wire g743_n;
  wire g744_p;
  wire g744_n;
  wire g745_p;
  wire g745_n;
  wire g746_p;
  wire g746_n;
  wire g747_p;
  wire g747_n;
  wire g748_p;
  wire g748_n;
  wire g749_p;
  wire g749_n;
  wire g750_p;
  wire g750_n;
  wire g751_p;
  wire g751_n;
  wire g752_p;
  wire g752_n;
  wire g753_p;
  wire g753_n;
  wire g754_p;
  wire g754_n;
  wire g755_p;
  wire g755_n;
  wire g756_p;
  wire g756_n;
  wire g757_p;
  wire g757_n;
  wire g758_p;
  wire g758_n;
  wire g759_p;
  wire g759_n;
  wire g760_p;
  wire g760_n;
  wire g761_p;
  wire g761_n;
  wire g762_p;
  wire g762_n;
  wire g763_p;
  wire g763_n;
  wire g764_p;
  wire g764_n;
  wire g765_p;
  wire g765_n;
  wire g766_p;
  wire g766_n;
  wire g767_p;
  wire g767_n;
  wire g768_p;
  wire g768_n;
  wire g769_p;
  wire g769_n;
  wire g770_p;
  wire g770_n;
  wire g771_p;
  wire g771_n;
  wire g772_p;
  wire g772_n;
  wire g773_p;
  wire g773_n;
  wire g774_p;
  wire g774_n;
  wire g775_p;
  wire g775_n;
  wire g776_p;
  wire g776_n;
  wire g777_p;
  wire g777_n;
  wire g778_p;
  wire g778_n;
  wire g779_p;
  wire g779_n;
  wire g780_p;
  wire g780_n;
  wire g781_p;
  wire g781_n;
  wire g782_p;
  wire g782_n;
  wire g783_p;
  wire g783_n;
  wire g784_p;
  wire g784_n;
  wire g785_p;
  wire g785_n;
  wire g786_p;
  wire g786_n;
  wire g787_p;
  wire g787_n;
  wire g788_p;
  wire g788_n;
  wire g789_p;
  wire g789_n;
  wire g790_p;
  wire g790_n;
  wire g791_p;
  wire g791_n;
  wire g792_p;
  wire g792_n;
  wire g793_p;
  wire g793_n;
  wire g794_p;
  wire g794_n;
  wire g795_p;
  wire g795_n;
  wire g796_p;
  wire g796_n;
  wire g797_p;
  wire g797_n;
  wire g798_p;
  wire g798_n;
  wire g799_p;
  wire g799_n;
  wire g800_p;
  wire g800_n;
  wire g801_p;
  wire g801_n;
  wire g802_p;
  wire g802_n;
  wire g803_p;
  wire g803_n;
  wire g804_p;
  wire g804_n;
  wire g805_p;
  wire g805_n;
  wire g806_p;
  wire g806_n;
  wire g807_p;
  wire g807_n;
  wire g808_p;
  wire g808_n;
  wire g809_p;
  wire g809_n;
  wire g810_p;
  wire g810_n;
  wire g811_p;
  wire g811_n;
  wire g812_p;
  wire g812_n;
  wire g813_p;
  wire g813_n;
  wire g814_p;
  wire g814_n;
  wire g815_p;
  wire g815_n;
  wire g816_p;
  wire g816_n;
  wire g817_p;
  wire g817_n;
  wire g818_p;
  wire g818_n;
  wire g819_p;
  wire g819_n;
  wire g820_p;
  wire g820_n;
  wire g821_p;
  wire g821_n;
  wire g822_p;
  wire g822_n;
  wire g823_p;
  wire g823_n;
  wire g824_p;
  wire g824_n;
  wire g825_p;
  wire g825_n;
  wire g826_p;
  wire g826_n;
  wire g827_p;
  wire g827_n;
  wire g828_p;
  wire g828_n;
  wire g829_p;
  wire g829_n;
  wire g830_p;
  wire g830_n;
  wire g831_p;
  wire g831_n;
  wire g832_p;
  wire g832_n;
  wire g833_p;
  wire g833_n;
  wire g834_p;
  wire g834_n;
  wire g835_p;
  wire g835_n;
  wire g836_p;
  wire g836_n;
  wire g837_p;
  wire g837_n;
  wire g838_p;
  wire g838_n;
  wire g839_p;
  wire g839_n;
  wire g840_p;
  wire g840_n;
  wire g841_p;
  wire g841_n;
  wire g842_p;
  wire g842_n;
  wire g843_p;
  wire g843_n;
  wire g844_p;
  wire g844_n;
  wire g845_p;
  wire g845_n;
  wire g846_p;
  wire g846_n;
  wire g847_p;
  wire g847_n;
  wire g848_p;
  wire g848_n;
  wire g849_p;
  wire g849_n;
  wire g850_p;
  wire g850_n;
  wire g851_p;
  wire g851_n;
  wire g852_p;
  wire g852_n;
  wire g853_p;
  wire g853_n;
  wire g854_p;
  wire g854_n;
  wire g855_p;
  wire g855_n;
  wire g856_p;
  wire g856_n;
  wire g857_p;
  wire g857_n;
  wire g858_p;
  wire g858_n;
  wire g859_p;
  wire g859_n;
  wire g860_p;
  wire g860_n;
  wire g861_p;
  wire g861_n;
  wire g862_p;
  wire g862_n;
  wire g863_p;
  wire g863_n;
  wire g864_p;
  wire g864_n;
  wire g865_p;
  wire g865_n;
  wire g866_p;
  wire g866_n;
  wire g867_p;
  wire g867_n;
  wire g868_p;
  wire g868_n;
  wire g869_p;
  wire g869_n;
  wire g870_p;
  wire g870_n;
  wire g871_p;
  wire g871_n;
  wire g872_p;
  wire g872_n;
  wire g873_p;
  wire g873_n;
  wire g874_p;
  wire g874_n;
  wire g875_p;
  wire g875_n;
  wire g876_p;
  wire g876_n;
  wire g877_p;
  wire g877_n;
  wire g878_p;
  wire g878_n;
  wire g879_p;
  wire g879_n;
  wire g880_p;
  wire g880_n;
  wire g881_p;
  wire g881_n;
  wire g882_p;
  wire g882_n;
  wire g883_p;
  wire g883_n;
  wire g884_p;
  wire g884_n;
  wire g885_p;
  wire g885_n;
  wire g886_p;
  wire g886_n;
  wire g887_p;
  wire g887_n;
  wire g888_p;
  wire g888_n;
  wire g889_p;
  wire g889_n;
  wire g890_p;
  wire g890_n;
  wire g891_p;
  wire g891_n;
  wire g892_p;
  wire g892_n;
  wire g893_p;
  wire g893_n;
  wire g894_p;
  wire g894_n;
  wire g895_p;
  wire g895_n;
  wire g896_p;
  wire g896_n;
  wire g897_p;
  wire g897_n;
  wire g898_p;
  wire g898_n;
  wire g899_p;
  wire g899_n;
  wire g900_p;
  wire g900_n;
  wire g901_p;
  wire g901_n;
  wire g902_p;
  wire g902_n;
  wire g903_p;
  wire g903_n;
  wire g904_p;
  wire g904_n;
  wire g905_p;
  wire g905_n;
  wire g906_p;
  wire g906_n;
  wire g907_p;
  wire g907_n;
  wire g908_p;
  wire g908_n;
  wire g909_p;
  wire g909_n;
  wire g910_p;
  wire g910_n;
  wire g911_p;
  wire g911_n;
  wire g912_p;
  wire g912_n;
  wire g913_p;
  wire g913_n;
  wire g914_p;
  wire g914_n;
  wire g915_p;
  wire g915_n;
  wire g916_p;
  wire g916_n;
  wire g917_p;
  wire g917_n;
  wire g918_p;
  wire g918_n;
  wire g919_p;
  wire g919_n;
  wire g920_p;
  wire g920_n;
  wire g921_p;
  wire g921_n;
  wire g922_p;
  wire g922_n;
  wire g923_p;
  wire g923_n;
  wire g924_p;
  wire g924_n;
  wire g925_p;
  wire g925_n;
  wire g926_p;
  wire g926_n;
  wire g927_p;
  wire g927_n;
  wire g928_p;
  wire g928_n;
  wire g929_p;
  wire g929_n;
  wire g930_p;
  wire g930_n;
  wire g931_p;
  wire g931_n;
  wire g932_p;
  wire g932_n;
  wire g933_p;
  wire g933_n;
  wire g934_p;
  wire g934_n;
  wire g935_p;
  wire g935_n;
  wire g936_p;
  wire g936_n;
  wire g937_p;
  wire g937_n;
  wire g938_p;
  wire g938_n;
  wire g939_p;
  wire g939_n;
  wire g940_p;
  wire g940_n;
  wire g941_p;
  wire g941_n;
  wire g942_p;
  wire g942_n;
  wire g943_p;
  wire g943_n;
  wire g944_p;
  wire g944_n;
  wire g945_p;
  wire g945_n;
  wire g946_p;
  wire g946_n;
  wire g947_p;
  wire g947_n;
  wire g948_p;
  wire g948_n;
  wire g949_p;
  wire g949_n;
  wire g950_p;
  wire g950_n;
  wire g951_p;
  wire g951_n;
  wire g952_p;
  wire g952_n;
  wire g953_p;
  wire g953_n;
  wire g954_p;
  wire g954_n;
  wire g955_p;
  wire g955_n;
  wire g956_p;
  wire g956_n;
  wire g957_p;
  wire g957_n;
  wire g958_p;
  wire g958_n;
  wire g959_p;
  wire g959_n;
  wire g960_p;
  wire g960_n;
  wire g961_p;
  wire g961_n;
  wire g962_p;
  wire g962_n;
  wire g963_p;
  wire g963_n;
  wire g964_p;
  wire g964_n;
  wire g965_p;
  wire g965_n;
  wire g966_p;
  wire g966_n;
  wire g967_p;
  wire g967_n;
  wire g968_p;
  wire g968_n;
  wire g969_p;
  wire g969_n;
  wire g970_p;
  wire g970_n;
  wire g971_p;
  wire g971_n;
  wire g972_p;
  wire g972_n;
  wire g973_p;
  wire g973_n;
  wire g974_p;
  wire g974_n;
  wire g975_p;
  wire g975_n;
  wire g976_p;
  wire g976_n;
  wire g977_p;
  wire g977_n;
  wire g978_p;
  wire g978_n;
  wire g979_p;
  wire g979_n;
  wire g980_p;
  wire g980_n;
  wire g981_p;
  wire g981_n;
  wire g982_p;
  wire g982_n;
  wire g983_p;
  wire g983_n;
  wire g984_p;
  wire g984_n;
  wire g985_p;
  wire g985_n;
  wire g986_p;
  wire g986_n;
  wire g987_p;
  wire g987_n;
  wire g988_p;
  wire g988_n;
  wire g989_p;
  wire g989_n;
  wire g990_p;
  wire g990_n;
  wire g991_p;
  wire g991_n;
  wire g992_p;
  wire g992_n;
  wire g993_p;
  wire g993_n;
  wire g994_p;
  wire g994_n;
  wire g995_p;
  wire g995_n;
  wire g996_p;
  wire g996_n;
  wire g997_p;
  wire g997_n;
  wire g998_p;
  wire g998_n;
  wire g999_p;
  wire g999_n;
  wire g1000_p;
  wire g1000_n;
  wire g1001_p;
  wire g1001_n;
  wire g1002_p;
  wire g1002_n;
  wire g1003_p;
  wire g1003_n;
  wire g1004_p;
  wire g1004_n;
  wire g1005_p;
  wire g1005_n;
  wire g1006_p;
  wire g1006_n;
  wire g1007_p;
  wire g1007_n;
  wire g1008_p;
  wire g1008_n;
  wire g1009_p;
  wire g1009_n;
  wire g1010_p;
  wire g1010_n;
  wire g1011_p;
  wire g1011_n;
  wire g1012_p;
  wire g1012_n;
  wire g1013_p;
  wire g1013_n;
  wire g1014_p;
  wire g1014_n;
  wire g1015_p;
  wire g1015_n;
  wire g1016_p;
  wire g1016_n;
  wire g1017_p;
  wire g1017_n;
  wire g1018_p;
  wire g1018_n;
  wire g1019_p;
  wire g1019_n;
  wire g1020_p;
  wire g1020_n;
  wire g1021_p;
  wire g1021_n;
  wire g1022_p;
  wire g1022_n;
  wire g1023_p;
  wire g1023_n;
  wire g1024_p;
  wire g1024_n;
  wire g1025_p;
  wire g1025_n;
  wire g1026_p;
  wire g1026_n;
  wire g1027_p;
  wire g1027_n;
  wire g1028_p;
  wire g1028_n;
  wire g1029_p;
  wire g1029_n;
  wire g1030_p;
  wire g1030_n;
  wire g1031_p;
  wire g1031_n;
  wire g1032_p;
  wire g1032_n;
  wire g1033_p;
  wire g1033_n;
  wire g1034_p;
  wire g1034_n;
  wire g1035_p;
  wire g1035_n;
  wire g1036_p;
  wire g1036_n;
  wire g1037_p;
  wire g1037_n;
  wire g1038_p;
  wire g1038_n;
  wire g1039_p;
  wire g1039_n;
  wire g1040_p;
  wire g1040_n;
  wire g1041_p;
  wire g1041_n;
  wire g1042_p;
  wire g1042_n;
  wire g1043_p;
  wire g1043_n;
  wire g1044_p;
  wire g1044_n;
  wire g1045_p;
  wire g1045_n;
  wire g1046_p;
  wire g1046_n;
  wire g1047_p;
  wire g1047_n;
  wire g1048_p;
  wire g1048_n;
  wire g1049_p;
  wire g1049_n;
  wire g1050_p;
  wire g1050_n;
  wire g1051_p;
  wire g1051_n;
  wire g1052_p;
  wire g1052_n;
  wire g1053_p;
  wire g1053_n;
  wire g1054_p;
  wire g1054_n;
  wire g1055_p;
  wire g1055_n;
  wire g1056_p;
  wire g1056_n;
  wire g1057_p;
  wire g1057_n;
  wire g1058_p;
  wire g1058_n;
  wire g1059_p;
  wire g1059_n;
  wire g1060_p;
  wire g1060_n;
  wire g1061_p;
  wire g1061_n;
  wire g1062_p;
  wire g1062_n;
  wire g1063_p;
  wire g1063_n;
  wire g1064_p;
  wire g1064_n;
  wire g1065_p;
  wire g1065_n;
  wire g1066_p;
  wire g1066_n;
  wire g1067_p;
  wire g1067_n;
  wire g1068_p;
  wire g1068_n;
  wire g1069_p;
  wire g1069_n;
  wire g1070_p;
  wire g1070_n;
  wire g1071_p;
  wire g1071_n;
  wire g1072_p;
  wire g1072_n;
  wire g1073_p;
  wire g1073_n;
  wire g1074_p;
  wire g1074_n;
  wire g1075_p;
  wire g1075_n;
  wire g1076_p;
  wire g1076_n;
  wire g1077_p;
  wire g1077_n;
  wire g1078_p;
  wire g1078_n;
  wire g1079_p;
  wire g1079_n;
  wire g1080_p;
  wire g1080_n;
  wire g1081_p;
  wire g1081_n;
  wire g1082_p;
  wire g1082_n;
  wire g1083_p;
  wire g1083_n;
  wire g1084_p;
  wire g1084_n;
  wire g1085_p;
  wire g1085_n;
  wire g1086_p;
  wire g1086_n;
  wire g1087_p;
  wire g1087_n;
  wire g1088_p;
  wire g1088_n;
  wire g1089_p;
  wire g1089_n;
  wire g1090_p;
  wire g1090_n;
  wire g1091_p;
  wire g1091_n;
  wire g1092_p;
  wire g1092_n;
  wire g1093_p;
  wire g1093_n;
  wire g1094_p;
  wire g1094_n;
  wire g1095_p;
  wire g1095_n;
  wire g1096_p;
  wire g1096_n;
  wire g1097_p;
  wire g1097_n;
  wire g1098_p;
  wire g1098_n;
  wire g1099_p;
  wire g1099_n;
  wire g1100_p;
  wire g1100_n;
  wire g1101_p;
  wire g1101_n;
  wire g1102_p;
  wire g1102_n;
  wire g1103_p;
  wire g1103_n;
  wire g1104_p;
  wire g1104_n;
  wire g1105_p;
  wire g1105_n;
  wire g1106_p;
  wire g1106_n;
  wire g1107_p;
  wire g1107_n;
  wire g1108_p;
  wire g1108_n;
  wire g1109_p;
  wire g1109_n;
  wire g1110_p;
  wire g1110_n;
  wire g1111_p;
  wire g1111_n;
  wire g1112_p;
  wire g1112_n;
  wire g1113_p;
  wire g1113_n;
  wire g1114_p;
  wire g1114_n;
  wire g1115_p;
  wire g1115_n;
  wire g1116_p;
  wire g1116_n;
  wire g1117_p;
  wire g1117_n;
  wire g1118_p;
  wire g1118_n;
  wire g1119_p;
  wire g1119_n;
  wire g1120_p;
  wire g1120_n;
  wire g1121_p;
  wire g1121_n;
  wire g1122_p;
  wire g1122_n;
  wire g1123_p;
  wire g1123_n;
  wire g1124_p;
  wire g1124_n;
  wire g1125_p;
  wire g1125_n;
  wire g1126_p;
  wire g1126_n;
  wire g1127_p;
  wire g1127_n;
  wire g1128_p;
  wire g1128_n;
  wire g1129_p;
  wire g1129_n;
  wire g1130_p;
  wire g1130_n;
  wire g1131_p;
  wire g1131_n;
  wire g1132_p;
  wire g1132_n;
  wire g1133_p;
  wire g1133_n;
  wire g1134_p;
  wire g1134_n;
  wire g1135_p;
  wire g1135_n;
  wire g1136_p;
  wire g1136_n;
  wire g1137_p;
  wire g1137_n;
  wire g1138_p;
  wire g1138_n;
  wire g1139_p;
  wire g1139_n;
  wire g1140_p;
  wire g1140_n;
  wire g1141_p;
  wire g1141_n;
  wire g1142_p;
  wire g1142_n;
  wire g1143_p;
  wire g1143_n;
  wire g1144_p;
  wire g1144_n;
  wire g1145_p;
  wire g1145_n;
  wire g1146_p;
  wire g1146_n;
  wire g1147_p;
  wire g1147_n;
  wire g1148_p;
  wire g1148_n;
  wire g1149_p;
  wire g1149_n;
  wire g1150_p;
  wire g1150_n;
  wire g1151_p;
  wire g1151_n;
  wire g1152_p;
  wire g1152_n;
  wire g1153_p;
  wire g1153_n;
  wire g1154_p;
  wire g1154_n;
  wire g1155_p;
  wire g1155_n;
  wire g1156_p;
  wire g1156_n;
  wire g1157_p;
  wire g1157_n;
  wire g1158_p;
  wire g1158_n;
  wire g1159_p;
  wire g1159_n;
  wire g1160_p;
  wire g1160_n;
  wire g1161_p;
  wire g1161_n;
  wire g1162_p;
  wire g1162_n;
  wire g1163_p;
  wire g1163_n;
  wire g1164_p;
  wire g1164_n;
  wire g1165_p;
  wire g1165_n;
  wire g1166_p;
  wire g1166_n;
  wire g1167_p;
  wire g1167_n;
  wire g1168_p;
  wire g1168_n;
  wire g1169_p;
  wire g1169_n;
  wire g1170_p;
  wire g1170_n;
  wire g1171_p;
  wire g1171_n;
  wire g1172_p;
  wire g1172_n;
  wire g1173_p;
  wire g1173_n;
  wire g1174_p;
  wire g1174_n;
  wire g1175_p;
  wire g1175_n;
  wire g1176_p;
  wire g1176_n;
  wire g1177_p;
  wire g1177_n;
  wire g1178_p;
  wire g1178_n;
  wire g1179_p;
  wire g1179_n;
  wire g1180_p;
  wire g1180_n;
  wire g1181_p;
  wire g1181_n;
  wire g1182_p;
  wire g1182_n;
  wire g1183_p;
  wire g1183_n;
  wire g1184_p;
  wire g1184_n;
  wire g1185_p;
  wire g1185_n;
  wire g1186_p;
  wire g1186_n;
  wire g1187_p;
  wire g1187_n;
  wire g1188_p;
  wire g1188_n;
  wire g1189_p;
  wire g1189_n;
  wire g1190_p;
  wire g1190_n;
  wire g1191_p;
  wire g1191_n;
  wire g1192_p;
  wire g1192_n;
  wire g1193_p;
  wire g1193_n;
  wire g1194_p;
  wire g1194_n;
  wire g1195_p;
  wire g1195_n;
  wire g1196_p;
  wire g1196_n;
  wire g1197_p;
  wire g1197_n;
  wire g1198_p;
  wire g1198_n;
  wire g1199_p;
  wire g1199_n;
  wire g1200_p;
  wire g1200_n;
  wire g1201_p;
  wire g1201_n;
  wire g1202_p;
  wire g1202_n;
  wire g1203_p;
  wire g1203_n;
  wire g1204_p;
  wire g1204_n;
  wire g1205_p;
  wire g1205_n;
  wire g1206_p;
  wire g1206_n;
  wire g1207_p;
  wire g1207_n;
  wire g1208_p;
  wire g1208_n;
  wire g1209_p;
  wire g1209_n;
  wire g1210_p;
  wire g1210_n;
  wire g1211_p;
  wire g1211_n;
  wire g1212_p;
  wire g1212_n;
  wire g1213_p;
  wire g1213_n;
  wire g1214_p;
  wire g1214_n;
  wire g1215_p;
  wire g1215_n;
  wire g1216_p;
  wire g1216_n;
  wire g1217_p;
  wire g1217_n;
  wire g1218_p;
  wire g1218_n;
  wire g1219_p;
  wire g1219_n;
  wire g1220_p;
  wire g1220_n;
  wire g1221_p;
  wire g1221_n;
  wire g1222_p;
  wire g1222_n;
  wire g1223_p;
  wire g1223_n;
  wire g1224_p;
  wire g1224_n;
  wire g1225_p;
  wire g1225_n;
  wire g1226_p;
  wire g1226_n;
  wire g1227_p;
  wire g1227_n;
  wire g1228_p;
  wire g1228_n;
  wire g1229_p;
  wire g1229_n;
  wire g1230_p;
  wire g1230_n;
  wire g1231_p;
  wire g1231_n;
  wire g1232_p;
  wire g1232_n;
  wire g1233_p;
  wire g1233_n;
  wire g1234_p;
  wire g1234_n;
  wire g1235_p;
  wire g1235_n;
  wire g1236_p;
  wire g1236_n;
  wire g1237_p;
  wire g1237_n;
  wire g1238_p;
  wire g1238_n;
  wire g1239_p;
  wire g1239_n;
  wire g1240_p;
  wire g1240_n;
  wire g1241_p;
  wire g1241_n;
  wire g1242_p;
  wire g1242_n;
  wire g1243_p;
  wire g1243_n;
  wire g1244_p;
  wire g1244_n;
  wire g1245_p;
  wire g1245_n;
  wire g1246_p;
  wire g1246_n;
  wire g1247_p;
  wire g1247_n;
  wire g1248_p;
  wire g1248_n;
  wire g1249_p;
  wire g1249_n;
  wire g1250_p;
  wire g1250_n;
  wire g1251_p;
  wire g1251_n;
  wire g1252_p;
  wire g1252_n;
  wire g1253_p;
  wire g1253_n;
  wire g1254_p;
  wire g1254_n;
  wire g1255_p;
  wire g1255_n;
  wire g1256_p;
  wire g1256_n;
  wire g1257_p;
  wire g1257_n;
  wire g1258_p;
  wire g1258_n;
  wire g1259_p;
  wire g1259_n;
  wire g1260_p;
  wire g1260_n;
  wire g1261_p;
  wire g1261_n;
  wire g1262_p;
  wire g1262_n;
  wire g1263_p;
  wire g1263_n;
  wire g1264_p;
  wire g1264_n;
  wire g1265_p;
  wire g1265_n;
  wire g1266_p;
  wire g1266_n;
  wire g1267_p;
  wire g1267_n;
  wire g1268_p;
  wire g1268_n;
  wire g1269_p;
  wire g1269_n;
  wire g1270_p;
  wire g1270_n;
  wire g1271_p;
  wire g1271_n;
  wire g1272_p;
  wire g1272_n;
  wire g1273_p;
  wire g1273_n;
  wire g1274_p;
  wire g1274_n;
  wire g1275_p;
  wire g1275_n;
  wire g1276_p;
  wire g1276_n;
  wire g1277_p;
  wire g1277_n;
  wire g1278_p;
  wire g1278_n;
  wire g1279_p;
  wire g1279_n;
  wire g1280_p;
  wire g1280_n;
  wire g1281_p;
  wire g1281_n;
  wire g1282_p;
  wire g1282_n;
  wire g1283_p;
  wire g1283_n;
  wire g1284_p;
  wire g1284_n;
  wire g1285_p;
  wire g1285_n;
  wire g1286_p;
  wire g1286_n;
  wire g1287_p;
  wire g1287_n;
  wire g1288_p;
  wire g1288_n;
  wire g1289_p;
  wire g1289_n;
  wire g1290_p;
  wire g1290_n;
  wire g1291_p;
  wire g1291_n;
  wire g1292_p;
  wire g1292_n;
  wire g1293_p;
  wire g1293_n;
  wire g1294_p;
  wire g1294_n;
  wire g1295_p;
  wire g1295_n;
  wire g1296_p;
  wire g1296_n;
  wire g1297_p;
  wire g1297_n;
  wire g1298_p;
  wire g1298_n;
  wire g1299_p;
  wire g1299_n;
  wire g1300_p;
  wire g1300_n;
  wire g1301_p;
  wire g1301_n;
  wire g1302_p;
  wire g1302_n;
  wire g1303_p;
  wire g1303_n;
  wire g1304_p;
  wire g1304_n;
  wire g1305_p;
  wire g1305_n;
  wire g1306_p;
  wire g1306_n;
  wire g1307_p;
  wire g1307_n;
  wire g1308_p;
  wire g1308_n;
  wire g1309_p;
  wire g1309_n;
  wire g1310_p;
  wire g1310_n;
  wire g1311_p;
  wire g1311_n;
  wire g1312_p;
  wire g1312_n;
  wire g1313_p;
  wire g1313_n;
  wire g1314_p;
  wire g1314_n;
  wire g1315_p;
  wire g1315_n;
  wire g1316_p;
  wire g1316_n;
  wire g1317_p;
  wire g1317_n;
  wire g1318_p;
  wire g1318_n;
  wire g1319_p;
  wire g1319_n;
  wire g1320_p;
  wire g1320_n;
  wire g1321_p;
  wire g1321_n;
  wire g1322_p;
  wire g1322_n;
  wire g1323_p;
  wire g1323_n;
  wire g1324_p;
  wire g1324_n;
  wire g1325_p;
  wire g1325_n;
  wire g1326_p;
  wire g1326_n;
  wire g1327_p;
  wire g1327_n;
  wire g1328_p;
  wire g1328_n;
  wire g1329_p;
  wire g1329_n;
  wire g1330_p;
  wire g1330_n;
  wire g1331_p;
  wire g1331_n;
  wire g1332_p;
  wire g1332_n;
  wire g1333_p;
  wire g1333_n;
  wire g1334_p;
  wire g1334_n;
  wire g1335_p;
  wire g1335_n;
  wire g1336_p;
  wire g1336_n;
  wire g1337_p;
  wire g1337_n;
  wire g1338_p;
  wire g1338_n;
  wire g1339_p;
  wire g1339_n;
  wire g1340_p;
  wire g1340_n;
  wire g1341_p;
  wire g1341_n;
  wire g1342_p;
  wire g1342_n;
  wire g1343_p;
  wire g1343_n;
  wire g1344_p;
  wire g1344_n;
  wire g1345_p;
  wire g1345_n;
  wire g1346_p;
  wire g1346_n;
  wire g1347_p;
  wire g1347_n;
  wire g1348_p;
  wire g1348_n;
  wire g1349_p;
  wire g1349_n;
  wire g1350_p;
  wire g1350_n;
  wire g1351_p;
  wire g1351_n;
  wire g1352_p;
  wire g1352_n;
  wire g1353_p;
  wire g1353_n;
  wire g1354_p;
  wire g1354_n;
  wire g1355_p;
  wire g1355_n;
  wire g1356_p;
  wire g1356_n;
  wire g1357_p;
  wire g1357_n;
  wire g1358_p;
  wire g1358_n;
  wire g1359_p;
  wire g1359_n;
  wire g1360_p;
  wire g1360_n;
  wire g1361_p;
  wire g1361_n;
  wire g1362_p;
  wire g1362_n;
  wire g1363_p;
  wire g1363_n;
  wire g1364_p;
  wire g1364_n;
  wire g1365_p;
  wire g1365_n;
  wire g1366_p;
  wire g1366_n;
  wire g1367_p;
  wire g1367_n;
  wire g1368_p;
  wire g1368_n;
  wire g1369_p;
  wire g1369_n;
  wire g1370_p;
  wire g1370_n;
  wire g1371_p;
  wire g1371_n;
  wire g1372_p;
  wire g1372_n;
  wire g1373_p;
  wire g1373_n;
  wire g1374_p;
  wire g1374_n;
  wire g1375_p;
  wire g1375_n;
  wire g1376_p;
  wire g1376_n;
  wire g1377_p;
  wire g1377_n;
  wire g1378_p;
  wire g1378_n;
  wire g1379_p;
  wire g1379_n;
  wire g1380_p;
  wire g1380_n;
  wire g1381_p;
  wire g1381_n;
  wire g1382_p;
  wire g1382_n;
  wire g1383_p;
  wire g1383_n;
  wire g1384_p;
  wire g1384_n;
  wire g1385_p;
  wire g1385_n;
  wire g1386_p;
  wire g1386_n;
  wire g1387_p;
  wire g1387_n;
  wire g1388_p;
  wire g1388_n;
  wire g1389_p;
  wire g1389_n;
  wire g1390_p;
  wire g1390_n;
  wire g1391_p;
  wire g1391_n;
  wire g1392_p;
  wire g1392_n;
  wire g1393_p;
  wire g1393_n;
  wire g1394_p;
  wire g1394_n;
  wire g1395_p;
  wire g1395_n;
  wire g1396_p;
  wire g1396_n;
  wire g1397_p;
  wire g1397_n;
  wire g1398_p;
  wire g1398_n;
  wire g1399_p;
  wire g1399_n;
  wire g1400_p;
  wire g1400_n;
  wire g1401_p;
  wire g1401_n;
  wire g1402_p;
  wire g1402_n;
  wire g1403_p;
  wire g1403_n;
  wire g1404_p;
  wire g1404_n;
  wire g1405_p;
  wire g1405_n;
  wire g1406_p;
  wire g1406_n;
  wire g1407_p;
  wire g1407_n;
  wire g1408_p;
  wire g1408_n;
  wire g1409_p;
  wire g1409_n;
  wire g1410_p;
  wire g1410_n;
  wire g1411_p;
  wire g1411_n;
  wire g1412_p;
  wire g1412_n;
  wire g1413_p;
  wire g1413_n;
  wire g1414_p;
  wire g1414_n;
  wire g1415_p;
  wire g1415_n;
  wire g1416_p;
  wire g1416_n;
  wire g1417_p;
  wire g1417_n;
  wire g1418_p;
  wire g1418_n;
  wire g1419_p;
  wire g1419_n;
  wire g1420_p;
  wire g1420_n;
  wire g1421_p;
  wire g1421_n;
  wire g1422_p;
  wire g1422_n;
  wire g1423_p;
  wire g1423_n;
  wire g1424_p;
  wire g1424_n;
  wire g1425_p;
  wire g1425_n;
  wire g1426_p;
  wire g1426_n;
  wire g1427_p;
  wire g1427_n;
  wire g1428_p;
  wire g1428_n;
  wire g1429_p;
  wire g1429_n;
  wire g1430_p;
  wire g1430_n;
  wire g1431_p;
  wire g1431_n;
  wire g1432_p;
  wire g1432_n;
  wire g1433_p;
  wire g1433_n;
  wire g1434_p;
  wire g1434_n;
  wire g1435_p;
  wire g1435_n;
  wire g1436_p;
  wire g1436_n;
  wire g1437_p;
  wire g1437_n;
  wire g1438_p;
  wire g1438_n;
  wire g1439_p;
  wire g1439_n;
  wire g1440_p;
  wire g1440_n;
  wire g1441_p;
  wire g1441_n;
  wire g1442_p;
  wire g1442_n;
  wire g1443_p;
  wire g1443_n;
  wire g1444_p;
  wire g1444_n;
  wire g1445_p;
  wire g1445_n;
  wire g1446_p;
  wire g1446_n;
  wire g1447_p;
  wire g1447_n;
  wire g1448_p;
  wire g1448_n;
  wire g1449_p;
  wire g1449_n;
  wire g1450_p;
  wire g1450_n;
  wire g1451_p;
  wire g1451_n;
  wire g1452_p;
  wire g1452_n;
  wire g1453_p;
  wire g1453_n;
  wire g1454_p;
  wire g1454_n;
  wire g1455_p;
  wire g1455_n;
  wire g1456_p;
  wire g1456_n;
  wire g1457_p;
  wire g1457_n;
  wire g1458_p;
  wire g1458_n;
  wire g1459_p;
  wire g1459_n;
  wire g1460_p;
  wire g1460_n;
  wire g1461_p;
  wire g1461_n;
  wire g1462_p;
  wire g1462_n;
  wire g1463_p;
  wire g1463_n;
  wire g1464_p;
  wire g1464_n;
  wire g1465_p;
  wire g1465_n;
  wire g1466_p;
  wire g1466_n;
  wire g1467_p;
  wire g1467_n;
  wire g1468_p;
  wire g1468_n;
  wire g1469_p;
  wire g1469_n;
  wire g1470_p;
  wire g1470_n;
  wire g1471_p;
  wire g1471_n;
  wire g1472_p;
  wire g1472_n;
  wire g1473_p;
  wire g1473_n;
  wire g1474_p;
  wire g1474_n;
  wire g1475_p;
  wire g1475_n;
  wire g1476_p;
  wire g1476_n;
  wire g1477_p;
  wire g1477_n;
  wire g1478_p;
  wire g1478_n;
  wire g1479_p;
  wire g1479_n;
  wire g1480_p;
  wire g1480_n;
  wire g1481_p;
  wire g1481_n;
  wire g1482_p;
  wire g1482_n;
  wire g1483_p;
  wire g1483_n;
  wire g1484_p;
  wire g1484_n;
  wire g1485_p;
  wire g1485_n;
  wire g1486_p;
  wire g1486_n;
  wire g1487_p;
  wire g1487_n;
  wire g1488_p;
  wire g1488_n;
  wire g1489_p;
  wire g1489_n;
  wire g1490_p;
  wire g1490_n;
  wire g1491_p;
  wire g1491_n;
  wire g1492_p;
  wire g1492_n;
  wire g1493_p;
  wire g1493_n;
  wire g1494_p;
  wire g1494_n;
  wire g1495_p;
  wire g1495_n;
  wire g1496_p;
  wire g1496_n;
  wire g1497_p;
  wire g1497_n;
  wire g1498_p;
  wire g1498_n;
  wire g1499_p;
  wire g1499_n;
  wire g1500_p;
  wire g1500_n;
  wire g1501_p;
  wire g1501_n;
  wire g1502_p;
  wire g1502_n;
  wire g1503_p;
  wire g1503_n;
  wire g1504_p;
  wire g1504_n;
  wire g1505_p;
  wire g1505_n;
  wire g1506_p;
  wire g1506_n;
  wire g1507_p;
  wire g1507_n;
  wire g1508_p;
  wire g1508_n;
  wire g1509_p;
  wire g1509_n;
  wire g1510_p;
  wire g1510_n;
  wire g1511_p;
  wire g1511_n;
  wire g1512_p;
  wire g1512_n;
  wire g1513_p;
  wire g1513_n;
  wire g1514_p;
  wire g1514_n;
  wire g1515_p;
  wire g1515_n;
  wire g1516_p;
  wire g1516_n;
  wire g1517_p;
  wire g1517_n;
  wire g1518_p;
  wire g1518_n;
  wire g1519_p;
  wire g1519_n;
  wire g1520_p;
  wire g1520_n;
  wire g1521_p;
  wire g1521_n;
  wire g1522_p;
  wire g1522_n;
  wire g1523_p;
  wire g1523_n;
  wire g1524_p;
  wire g1524_n;
  wire g1525_p;
  wire g1525_n;
  wire g1526_p;
  wire g1526_n;
  wire g1527_p;
  wire g1527_n;
  wire g1528_p;
  wire g1528_n;
  wire g1529_p;
  wire g1529_n;
  wire g1530_p;
  wire g1530_n;
  wire g1531_p;
  wire g1531_n;
  wire g1532_p;
  wire g1532_n;
  wire g1533_p;
  wire g1533_n;
  wire g1534_p;
  wire g1534_n;
  wire g1535_p;
  wire g1535_n;
  wire g1536_p;
  wire g1536_n;
  wire g1537_p;
  wire g1537_n;
  wire g1538_p;
  wire g1538_n;
  wire g1539_p;
  wire g1539_n;
  wire g1540_p;
  wire g1540_n;
  wire g1541_p;
  wire g1541_n;
  wire g1542_p;
  wire g1542_n;
  wire g1543_p;
  wire g1543_n;
  wire g1544_p;
  wire g1544_n;
  wire g1545_p;
  wire g1545_n;
  wire G153_n_spl_;
  wire G156_n_spl_;
  wire G66_p_spl_;
  wire G66_p_spl_0;
  wire G66_p_spl_00;
  wire G66_p_spl_01;
  wire G66_p_spl_1;
  wire G1_p_spl_;
  wire G165_n_spl_;
  wire G11_n_spl_;
  wire g185_n_spl_;
  wire g185_n_spl_0;
  wire g185_n_spl_00;
  wire g185_n_spl_000;
  wire g185_n_spl_01;
  wire g185_n_spl_1;
  wire g185_n_spl_10;
  wire g185_n_spl_11;
  wire G163_n_spl_;
  wire G163_n_spl_0;
  wire G163_n_spl_00;
  wire G163_n_spl_01;
  wire G163_n_spl_1;
  wire G163_p_spl_;
  wire G163_p_spl_0;
  wire G163_p_spl_00;
  wire G163_p_spl_01;
  wire G163_p_spl_1;
  wire G128_p_spl_;
  wire G128_p_spl_0;
  wire G128_p_spl_00;
  wire G128_p_spl_000;
  wire G128_p_spl_01;
  wire G128_p_spl_1;
  wire G128_p_spl_10;
  wire G128_p_spl_11;
  wire G168_p_spl_;
  wire G168_p_spl_0;
  wire G168_p_spl_00;
  wire G168_p_spl_000;
  wire G168_p_spl_001;
  wire G168_p_spl_01;
  wire G168_p_spl_010;
  wire G168_p_spl_1;
  wire G168_p_spl_10;
  wire G168_p_spl_11;
  wire G128_n_spl_;
  wire G128_n_spl_0;
  wire G128_n_spl_00;
  wire G128_n_spl_000;
  wire G128_n_spl_01;
  wire G128_n_spl_1;
  wire G128_n_spl_10;
  wire G128_n_spl_11;
  wire G169_p_spl_;
  wire G169_p_spl_0;
  wire G169_p_spl_00;
  wire G169_p_spl_000;
  wire G169_p_spl_001;
  wire G169_p_spl_01;
  wire G169_p_spl_010;
  wire G169_p_spl_011;
  wire G169_p_spl_1;
  wire G169_p_spl_10;
  wire G169_p_spl_11;
  wire G150_p_spl_;
  wire G150_p_spl_0;
  wire G150_p_spl_00;
  wire G150_p_spl_1;
  wire G167_n_spl_;
  wire G167_n_spl_0;
  wire G167_n_spl_00;
  wire G167_n_spl_000;
  wire G167_n_spl_001;
  wire G167_n_spl_01;
  wire G167_n_spl_010;
  wire G167_n_spl_1;
  wire G167_n_spl_10;
  wire G167_n_spl_11;
  wire G166_n_spl_;
  wire G166_n_spl_0;
  wire G166_n_spl_00;
  wire G166_n_spl_000;
  wire G166_n_spl_001;
  wire G166_n_spl_01;
  wire G166_n_spl_010;
  wire G166_n_spl_011;
  wire G166_n_spl_1;
  wire G166_n_spl_10;
  wire G166_n_spl_11;
  wire G150_n_spl_;
  wire G150_n_spl_0;
  wire G150_n_spl_00;
  wire G150_n_spl_1;
  wire G126_p_spl_;
  wire G126_p_spl_0;
  wire G126_p_spl_00;
  wire G126_p_spl_000;
  wire G126_p_spl_01;
  wire G126_p_spl_1;
  wire G126_p_spl_10;
  wire G126_p_spl_11;
  wire G126_n_spl_;
  wire G126_n_spl_0;
  wire G126_n_spl_00;
  wire G126_n_spl_000;
  wire G126_n_spl_01;
  wire G126_n_spl_1;
  wire G126_n_spl_10;
  wire G126_n_spl_11;
  wire G149_p_spl_;
  wire G149_p_spl_0;
  wire G149_p_spl_00;
  wire G149_p_spl_1;
  wire G149_n_spl_;
  wire G149_n_spl_0;
  wire G149_n_spl_00;
  wire G149_n_spl_1;
  wire g224_n_spl_;
  wire g233_n_spl_;
  wire G102_p_spl_;
  wire G102_p_spl_0;
  wire G102_p_spl_00;
  wire G102_p_spl_000;
  wire G102_p_spl_001;
  wire G102_p_spl_01;
  wire G102_p_spl_010;
  wire G102_p_spl_011;
  wire G102_p_spl_1;
  wire G102_p_spl_10;
  wire G102_p_spl_100;
  wire G102_p_spl_101;
  wire G102_p_spl_11;
  wire G102_p_spl_110;
  wire G113_p_spl_;
  wire G113_p_spl_0;
  wire G113_p_spl_00;
  wire G113_p_spl_1;
  wire G102_n_spl_;
  wire G102_n_spl_0;
  wire G102_n_spl_00;
  wire G102_n_spl_000;
  wire G102_n_spl_001;
  wire G102_n_spl_01;
  wire G102_n_spl_010;
  wire G102_n_spl_011;
  wire G102_n_spl_1;
  wire G102_n_spl_10;
  wire G102_n_spl_100;
  wire G102_n_spl_101;
  wire G102_n_spl_11;
  wire G102_n_spl_110;
  wire G113_n_spl_;
  wire G113_n_spl_0;
  wire G113_n_spl_00;
  wire G113_n_spl_01;
  wire G113_n_spl_1;
  wire G98_p_spl_;
  wire G98_p_spl_0;
  wire G98_p_spl_00;
  wire G98_p_spl_000;
  wire G98_p_spl_001;
  wire G98_p_spl_01;
  wire G98_p_spl_010;
  wire G98_p_spl_011;
  wire G98_p_spl_1;
  wire G98_p_spl_10;
  wire G98_p_spl_100;
  wire G98_p_spl_101;
  wire G98_p_spl_11;
  wire G98_p_spl_110;
  wire G98_p_spl_111;
  wire G98_n_spl_;
  wire G98_n_spl_0;
  wire G98_n_spl_00;
  wire G98_n_spl_000;
  wire G98_n_spl_001;
  wire G98_n_spl_01;
  wire G98_n_spl_010;
  wire G98_n_spl_011;
  wire G98_n_spl_1;
  wire G98_n_spl_10;
  wire G98_n_spl_100;
  wire G98_n_spl_101;
  wire G98_n_spl_11;
  wire G98_n_spl_110;
  wire G98_n_spl_111;
  wire G101_p_spl_;
  wire G101_p_spl_0;
  wire G101_p_spl_00;
  wire G101_p_spl_000;
  wire G101_p_spl_001;
  wire G101_p_spl_01;
  wire G101_p_spl_010;
  wire G101_p_spl_011;
  wire G101_p_spl_1;
  wire G101_p_spl_10;
  wire G101_p_spl_100;
  wire G101_p_spl_101;
  wire G101_p_spl_11;
  wire G101_p_spl_110;
  wire G101_p_spl_111;
  wire G115_p_spl_;
  wire G115_p_spl_0;
  wire G115_p_spl_00;
  wire G115_p_spl_1;
  wire G101_n_spl_;
  wire G101_n_spl_0;
  wire G101_n_spl_00;
  wire G101_n_spl_000;
  wire G101_n_spl_001;
  wire G101_n_spl_01;
  wire G101_n_spl_010;
  wire G101_n_spl_011;
  wire G101_n_spl_1;
  wire G101_n_spl_10;
  wire G101_n_spl_100;
  wire G101_n_spl_101;
  wire G101_n_spl_11;
  wire G101_n_spl_110;
  wire G101_n_spl_111;
  wire G115_n_spl_;
  wire G115_n_spl_0;
  wire G115_n_spl_00;
  wire G115_n_spl_1;
  wire G100_p_spl_;
  wire G100_p_spl_0;
  wire G100_p_spl_00;
  wire G100_p_spl_000;
  wire G100_p_spl_0000;
  wire G100_p_spl_001;
  wire G100_p_spl_01;
  wire G100_p_spl_010;
  wire G100_p_spl_011;
  wire G100_p_spl_1;
  wire G100_p_spl_10;
  wire G100_p_spl_100;
  wire G100_p_spl_101;
  wire G100_p_spl_11;
  wire G100_p_spl_110;
  wire G100_p_spl_111;
  wire G100_n_spl_;
  wire G100_n_spl_0;
  wire G100_n_spl_00;
  wire G100_n_spl_000;
  wire G100_n_spl_0000;
  wire G100_n_spl_001;
  wire G100_n_spl_01;
  wire G100_n_spl_010;
  wire G100_n_spl_011;
  wire G100_n_spl_1;
  wire G100_n_spl_10;
  wire G100_n_spl_100;
  wire G100_n_spl_101;
  wire G100_n_spl_11;
  wire G100_n_spl_110;
  wire G100_n_spl_111;
  wire g237_n_spl_;
  wire g237_n_spl_0;
  wire g237_n_spl_1;
  wire g240_p_spl_;
  wire g237_p_spl_;
  wire g240_n_spl_;
  wire g240_n_spl_0;
  wire g241_n_spl_;
  wire G130_p_spl_;
  wire G130_p_spl_0;
  wire G130_p_spl_00;
  wire G130_p_spl_1;
  wire G130_n_spl_;
  wire G130_n_spl_0;
  wire G130_n_spl_00;
  wire G130_n_spl_1;
  wire G148_n_spl_;
  wire G148_n_spl_0;
  wire G148_n_spl_00;
  wire G148_n_spl_1;
  wire G148_p_spl_;
  wire G148_p_spl_0;
  wire G148_p_spl_00;
  wire G148_p_spl_1;
  wire g245_n_spl_;
  wire g245_n_spl_0;
  wire g245_n_spl_1;
  wire g248_n_spl_;
  wire G119_p_spl_;
  wire G119_p_spl_0;
  wire G119_p_spl_00;
  wire G119_p_spl_01;
  wire G119_p_spl_1;
  wire G119_p_spl_10;
  wire G119_n_spl_;
  wire G119_n_spl_0;
  wire G119_n_spl_00;
  wire G119_n_spl_01;
  wire G119_n_spl_1;
  wire G119_n_spl_10;
  wire G146_p_spl_;
  wire G146_p_spl_0;
  wire G146_p_spl_1;
  wire G146_n_spl_;
  wire G146_n_spl_0;
  wire G146_n_spl_1;
  wire G117_p_spl_;
  wire G117_p_spl_0;
  wire G117_p_spl_00;
  wire G117_p_spl_01;
  wire G117_p_spl_1;
  wire G117_p_spl_10;
  wire G117_n_spl_;
  wire G117_n_spl_0;
  wire G117_n_spl_00;
  wire G117_n_spl_01;
  wire G117_n_spl_1;
  wire G117_n_spl_10;
  wire G145_p_spl_;
  wire G145_p_spl_0;
  wire G145_p_spl_1;
  wire G145_n_spl_;
  wire G145_n_spl_0;
  wire G145_n_spl_1;
  wire g258_p_spl_;
  wire g267_p_spl_;
  wire g258_n_spl_;
  wire g258_n_spl_0;
  wire g267_n_spl_;
  wire g267_n_spl_0;
  wire G121_p_spl_;
  wire G121_p_spl_0;
  wire G121_p_spl_00;
  wire G121_p_spl_000;
  wire G121_p_spl_01;
  wire G121_p_spl_1;
  wire G121_p_spl_10;
  wire G121_p_spl_11;
  wire G121_n_spl_;
  wire G121_n_spl_0;
  wire G121_n_spl_00;
  wire G121_n_spl_000;
  wire G121_n_spl_01;
  wire G121_n_spl_1;
  wire G121_n_spl_10;
  wire G121_n_spl_11;
  wire G147_p_spl_;
  wire G147_p_spl_0;
  wire G147_p_spl_00;
  wire G147_p_spl_1;
  wire G147_n_spl_;
  wire G147_n_spl_0;
  wire G147_n_spl_00;
  wire G147_n_spl_1;
  wire g268_n_spl_;
  wire g277_n_spl_;
  wire G107_p_spl_;
  wire G107_p_spl_0;
  wire G107_p_spl_00;
  wire G107_p_spl_000;
  wire G107_p_spl_01;
  wire G107_p_spl_1;
  wire G107_p_spl_10;
  wire G107_p_spl_11;
  wire G107_n_spl_;
  wire G107_n_spl_0;
  wire G107_n_spl_00;
  wire G107_n_spl_000;
  wire G107_n_spl_01;
  wire G107_n_spl_1;
  wire G107_n_spl_10;
  wire G107_n_spl_11;
  wire G139_p_spl_;
  wire G139_p_spl_0;
  wire G139_p_spl_00;
  wire G139_p_spl_1;
  wire G139_n_spl_;
  wire G139_n_spl_0;
  wire G139_n_spl_00;
  wire G139_n_spl_1;
  wire G105_p_spl_;
  wire G105_p_spl_0;
  wire G105_p_spl_00;
  wire G105_p_spl_000;
  wire G105_p_spl_01;
  wire G105_p_spl_1;
  wire G105_p_spl_10;
  wire G105_p_spl_11;
  wire G105_n_spl_;
  wire G105_n_spl_0;
  wire G105_n_spl_00;
  wire G105_n_spl_000;
  wire G105_n_spl_01;
  wire G105_n_spl_1;
  wire G105_n_spl_10;
  wire G105_n_spl_11;
  wire G138_p_spl_;
  wire G138_p_spl_0;
  wire G138_p_spl_00;
  wire G138_p_spl_1;
  wire G138_n_spl_;
  wire G138_n_spl_0;
  wire G138_n_spl_00;
  wire G138_n_spl_1;
  wire g289_n_spl_;
  wire g298_n_spl_;
  wire G109_p_spl_;
  wire G109_p_spl_0;
  wire G109_p_spl_00;
  wire G109_p_spl_000;
  wire G109_p_spl_01;
  wire G109_p_spl_1;
  wire G109_p_spl_10;
  wire G109_p_spl_11;
  wire G109_n_spl_;
  wire G109_n_spl_0;
  wire G109_n_spl_00;
  wire G109_n_spl_000;
  wire G109_n_spl_01;
  wire G109_n_spl_1;
  wire G109_n_spl_10;
  wire G109_n_spl_11;
  wire G135_p_spl_;
  wire G135_p_spl_0;
  wire G135_p_spl_00;
  wire G135_p_spl_1;
  wire G135_n_spl_;
  wire G135_n_spl_0;
  wire G135_n_spl_00;
  wire G135_n_spl_1;
  wire G88_p_spl_;
  wire G88_p_spl_0;
  wire G88_p_spl_00;
  wire G88_p_spl_01;
  wire G88_p_spl_1;
  wire G88_p_spl_10;
  wire G88_n_spl_;
  wire G88_n_spl_0;
  wire G88_n_spl_00;
  wire G88_n_spl_01;
  wire G88_n_spl_1;
  wire G88_n_spl_10;
  wire G142_p_spl_;
  wire G142_p_spl_0;
  wire G142_p_spl_1;
  wire G142_n_spl_;
  wire G142_n_spl_0;
  wire G142_n_spl_1;
  wire g308_n_spl_;
  wire g317_n_spl_;
  wire g317_n_spl_0;
  wire g317_n_spl_1;
  wire G90_p_spl_;
  wire G90_p_spl_0;
  wire G90_p_spl_00;
  wire G90_p_spl_000;
  wire G90_p_spl_01;
  wire G90_p_spl_1;
  wire G90_p_spl_10;
  wire G90_p_spl_11;
  wire G90_n_spl_;
  wire G90_n_spl_0;
  wire G90_n_spl_00;
  wire G90_n_spl_000;
  wire G90_n_spl_01;
  wire G90_n_spl_1;
  wire G90_n_spl_10;
  wire G90_n_spl_11;
  wire G143_p_spl_;
  wire G143_p_spl_0;
  wire G143_p_spl_00;
  wire G143_p_spl_1;
  wire G143_n_spl_;
  wire G143_n_spl_0;
  wire G143_n_spl_00;
  wire G143_n_spl_1;
  wire G92_p_spl_;
  wire G92_p_spl_0;
  wire G92_p_spl_00;
  wire G92_p_spl_000;
  wire G92_p_spl_01;
  wire G92_p_spl_1;
  wire G92_p_spl_10;
  wire G92_p_spl_11;
  wire G92_n_spl_;
  wire G92_n_spl_0;
  wire G92_n_spl_00;
  wire G92_n_spl_000;
  wire G92_n_spl_01;
  wire G92_n_spl_1;
  wire G92_n_spl_10;
  wire G92_n_spl_11;
  wire G144_p_spl_;
  wire G144_p_spl_0;
  wire G144_p_spl_00;
  wire G144_p_spl_1;
  wire G144_n_spl_;
  wire G144_n_spl_0;
  wire G144_n_spl_00;
  wire G144_n_spl_1;
  wire g328_n_spl_;
  wire g337_n_spl_;
  wire G94_p_spl_;
  wire G94_p_spl_0;
  wire G94_p_spl_00;
  wire G94_p_spl_000;
  wire G94_p_spl_01;
  wire G94_p_spl_1;
  wire G94_p_spl_10;
  wire G94_p_spl_11;
  wire G94_n_spl_;
  wire G94_n_spl_0;
  wire G94_n_spl_00;
  wire G94_n_spl_000;
  wire G94_n_spl_01;
  wire G94_n_spl_1;
  wire G94_n_spl_10;
  wire G94_n_spl_11;
  wire G140_p_spl_;
  wire G140_p_spl_0;
  wire G140_p_spl_00;
  wire G140_p_spl_1;
  wire G140_n_spl_;
  wire G140_n_spl_0;
  wire G140_n_spl_00;
  wire G140_n_spl_1;
  wire G96_p_spl_;
  wire G96_p_spl_0;
  wire G96_p_spl_00;
  wire G96_p_spl_000;
  wire G96_p_spl_01;
  wire G96_p_spl_1;
  wire G96_p_spl_10;
  wire G96_p_spl_11;
  wire G96_n_spl_;
  wire G96_n_spl_0;
  wire G96_n_spl_00;
  wire G96_n_spl_000;
  wire G96_n_spl_01;
  wire G96_n_spl_1;
  wire G96_n_spl_10;
  wire G96_n_spl_11;
  wire G141_p_spl_;
  wire G141_p_spl_0;
  wire G141_p_spl_00;
  wire G141_p_spl_1;
  wire G141_n_spl_;
  wire G141_n_spl_0;
  wire G141_n_spl_00;
  wire G141_n_spl_1;
  wire G103_p_spl_;
  wire G103_p_spl_0;
  wire G103_p_spl_00;
  wire G103_p_spl_000;
  wire G103_p_spl_01;
  wire G103_p_spl_1;
  wire G103_p_spl_10;
  wire G103_p_spl_11;
  wire G103_n_spl_;
  wire G103_n_spl_0;
  wire G103_n_spl_00;
  wire G103_n_spl_000;
  wire G103_n_spl_01;
  wire G103_n_spl_1;
  wire G103_n_spl_10;
  wire G103_n_spl_11;
  wire G137_p_spl_;
  wire G137_p_spl_0;
  wire G137_p_spl_00;
  wire G137_p_spl_1;
  wire G137_n_spl_;
  wire G137_n_spl_0;
  wire G137_n_spl_00;
  wire G137_n_spl_1;
  wire g356_n_spl_;
  wire g365_n_spl_;
  wire g347_n_spl_;
  wire G124_n_spl_;
  wire G124_n_spl_0;
  wire G124_n_spl_00;
  wire G124_n_spl_000;
  wire G124_n_spl_0000;
  wire G124_n_spl_0001;
  wire G124_n_spl_001;
  wire G124_n_spl_0010;
  wire G124_n_spl_0011;
  wire G124_n_spl_01;
  wire G124_n_spl_010;
  wire G124_n_spl_011;
  wire G124_n_spl_1;
  wire G124_n_spl_10;
  wire G124_n_spl_100;
  wire G124_n_spl_101;
  wire G124_n_spl_11;
  wire G124_n_spl_110;
  wire G124_n_spl_111;
  wire G124_p_spl_;
  wire G124_p_spl_0;
  wire G124_p_spl_00;
  wire G124_p_spl_000;
  wire G124_p_spl_0000;
  wire G124_p_spl_0001;
  wire G124_p_spl_001;
  wire G124_p_spl_0010;
  wire G124_p_spl_0011;
  wire G124_p_spl_01;
  wire G124_p_spl_010;
  wire G124_p_spl_011;
  wire G124_p_spl_1;
  wire G124_p_spl_10;
  wire G124_p_spl_100;
  wire G124_p_spl_101;
  wire G124_p_spl_11;
  wire G124_p_spl_110;
  wire G124_p_spl_111;
  wire g372_p_spl_;
  wire g372_p_spl_0;
  wire g372_p_spl_1;
  wire g372_n_spl_;
  wire g372_n_spl_0;
  wire g372_n_spl_1;
  wire g373_n_spl_;
  wire g373_n_spl_0;
  wire g374_n_spl_;
  wire g374_n_spl_0;
  wire g374_n_spl_1;
  wire g373_p_spl_;
  wire g373_p_spl_0;
  wire g374_p_spl_;
  wire g374_p_spl_0;
  wire g374_p_spl_1;
  wire g378_p_spl_;
  wire g378_p_spl_0;
  wire g378_p_spl_1;
  wire g378_n_spl_;
  wire g378_n_spl_0;
  wire g378_n_spl_1;
  wire g379_n_spl_;
  wire g380_n_spl_;
  wire g379_p_spl_;
  wire g380_p_spl_;
  wire g375_p_spl_;
  wire g375_p_spl_0;
  wire g375_p_spl_00;
  wire g375_p_spl_1;
  wire g381_p_spl_;
  wire g381_p_spl_0;
  wire g381_p_spl_00;
  wire g381_p_spl_01;
  wire g381_p_spl_1;
  wire g381_p_spl_10;
  wire g375_n_spl_;
  wire g375_n_spl_0;
  wire g375_n_spl_00;
  wire g375_n_spl_1;
  wire g381_n_spl_;
  wire g381_n_spl_0;
  wire g381_n_spl_00;
  wire g381_n_spl_01;
  wire g381_n_spl_1;
  wire g381_n_spl_10;
  wire g385_p_spl_;
  wire g385_p_spl_0;
  wire g385_p_spl_1;
  wire g385_n_spl_;
  wire g385_n_spl_0;
  wire g385_n_spl_1;
  wire g386_n_spl_;
  wire g387_n_spl_;
  wire g386_p_spl_;
  wire g387_p_spl_;
  wire g382_p_spl_;
  wire g388_p_spl_;
  wire g388_p_spl_0;
  wire g388_p_spl_00;
  wire g388_p_spl_01;
  wire g388_p_spl_1;
  wire g382_n_spl_;
  wire g388_n_spl_;
  wire g388_n_spl_0;
  wire g388_n_spl_00;
  wire g388_n_spl_01;
  wire g388_n_spl_1;
  wire g392_p_spl_;
  wire g392_p_spl_0;
  wire g392_p_spl_1;
  wire g392_n_spl_;
  wire g392_n_spl_0;
  wire g392_n_spl_1;
  wire g393_n_spl_;
  wire g389_n_spl_;
  wire g389_n_spl_0;
  wire g395_n_spl_;
  wire g395_n_spl_0;
  wire g395_n_spl_00;
  wire g395_n_spl_01;
  wire g395_n_spl_1;
  wire g395_n_spl_10;
  wire g399_p_spl_;
  wire g399_p_spl_0;
  wire g399_p_spl_1;
  wire g399_n_spl_;
  wire g399_n_spl_0;
  wire g399_n_spl_1;
  wire g400_n_spl_;
  wire g400_n_spl_0;
  wire g400_n_spl_00;
  wire g400_n_spl_1;
  wire g401_n_spl_;
  wire g401_n_spl_0;
  wire g400_p_spl_;
  wire g400_p_spl_0;
  wire g400_p_spl_00;
  wire g400_p_spl_1;
  wire g401_p_spl_;
  wire g401_p_spl_0;
  wire g405_p_spl_;
  wire g405_p_spl_0;
  wire g405_p_spl_1;
  wire g405_n_spl_;
  wire g405_n_spl_0;
  wire g405_n_spl_1;
  wire g406_n_spl_;
  wire g406_n_spl_0;
  wire g406_p_spl_;
  wire g406_p_spl_0;
  wire g402_p_spl_;
  wire g402_p_spl_0;
  wire g402_p_spl_1;
  wire g408_p_spl_;
  wire g408_p_spl_0;
  wire g408_p_spl_1;
  wire g402_n_spl_;
  wire g402_n_spl_0;
  wire g408_n_spl_;
  wire g408_n_spl_0;
  wire g408_n_spl_00;
  wire g408_n_spl_1;
  wire g412_p_spl_;
  wire g412_p_spl_0;
  wire g412_p_spl_1;
  wire g412_n_spl_;
  wire g412_n_spl_0;
  wire g412_n_spl_1;
  wire g413_n_spl_;
  wire g413_p_spl_;
  wire g409_p_spl_;
  wire g409_p_spl_0;
  wire g415_p_spl_;
  wire g415_p_spl_0;
  wire g415_p_spl_00;
  wire g415_p_spl_1;
  wire g409_n_spl_;
  wire g409_n_spl_0;
  wire g415_n_spl_;
  wire g415_n_spl_0;
  wire g415_n_spl_00;
  wire g415_n_spl_1;
  wire g419_p_spl_;
  wire g419_p_spl_0;
  wire g419_p_spl_1;
  wire g419_n_spl_;
  wire g419_n_spl_0;
  wire g419_n_spl_1;
  wire g420_n_spl_;
  wire g420_n_spl_0;
  wire g420_p_spl_;
  wire g420_p_spl_0;
  wire g416_p_spl_;
  wire g416_p_spl_0;
  wire g422_p_spl_;
  wire g422_p_spl_0;
  wire g422_p_spl_00;
  wire g422_p_spl_1;
  wire g416_n_spl_;
  wire g416_n_spl_0;
  wire g422_n_spl_;
  wire g422_n_spl_0;
  wire g422_n_spl_00;
  wire g422_n_spl_01;
  wire g422_n_spl_1;
  wire g426_p_spl_;
  wire g426_p_spl_0;
  wire g426_p_spl_1;
  wire g426_n_spl_;
  wire g426_n_spl_0;
  wire g426_n_spl_1;
  wire g427_n_spl_;
  wire g427_p_spl_;
  wire g423_p_spl_;
  wire g429_p_spl_;
  wire g429_p_spl_0;
  wire g429_p_spl_00;
  wire g429_p_spl_01;
  wire g429_p_spl_1;
  wire g429_p_spl_10;
  wire g423_n_spl_;
  wire g429_n_spl_;
  wire g429_n_spl_0;
  wire g429_n_spl_00;
  wire g429_n_spl_01;
  wire g429_n_spl_1;
  wire g429_n_spl_10;
  wire g396_n_spl_;
  wire g430_n_spl_;
  wire g430_n_spl_0;
  wire g430_n_spl_1;
  wire G123_n_spl_;
  wire G123_n_spl_0;
  wire G123_n_spl_00;
  wire G123_n_spl_000;
  wire G123_n_spl_0000;
  wire G123_n_spl_0001;
  wire G123_n_spl_001;
  wire G123_n_spl_0010;
  wire G123_n_spl_01;
  wire G123_n_spl_010;
  wire G123_n_spl_011;
  wire G123_n_spl_1;
  wire G123_n_spl_10;
  wire G123_n_spl_100;
  wire G123_n_spl_101;
  wire G123_n_spl_11;
  wire G123_n_spl_110;
  wire G123_n_spl_111;
  wire G123_p_spl_;
  wire G123_p_spl_0;
  wire G123_p_spl_00;
  wire G123_p_spl_000;
  wire G123_p_spl_0000;
  wire G123_p_spl_0001;
  wire G123_p_spl_001;
  wire G123_p_spl_0010;
  wire G123_p_spl_01;
  wire G123_p_spl_010;
  wire G123_p_spl_011;
  wire G123_p_spl_1;
  wire G123_p_spl_10;
  wire G123_p_spl_100;
  wire G123_p_spl_101;
  wire G123_p_spl_11;
  wire G123_p_spl_110;
  wire G123_p_spl_111;
  wire g434_p_spl_;
  wire g434_p_spl_0;
  wire g434_p_spl_1;
  wire g434_n_spl_;
  wire g434_n_spl_0;
  wire g434_n_spl_1;
  wire g435_n_spl_;
  wire g435_p_spl_;
  wire g440_p_spl_;
  wire g440_p_spl_0;
  wire g440_p_spl_1;
  wire g440_n_spl_;
  wire g440_n_spl_0;
  wire g440_n_spl_1;
  wire g441_n_spl_;
  wire g441_n_spl_0;
  wire g441_n_spl_00;
  wire g441_n_spl_1;
  wire g442_n_spl_;
  wire g442_n_spl_0;
  wire g442_n_spl_1;
  wire g441_p_spl_;
  wire g441_p_spl_0;
  wire g441_p_spl_00;
  wire g441_p_spl_1;
  wire g442_p_spl_;
  wire g442_p_spl_0;
  wire g442_p_spl_1;
  wire g437_p_spl_;
  wire g437_p_spl_0;
  wire g437_p_spl_00;
  wire g437_p_spl_01;
  wire g437_p_spl_1;
  wire g443_p_spl_;
  wire g443_p_spl_0;
  wire g443_p_spl_00;
  wire g443_p_spl_1;
  wire g437_n_spl_;
  wire g437_n_spl_0;
  wire g437_n_spl_00;
  wire g437_n_spl_01;
  wire g437_n_spl_1;
  wire g443_n_spl_;
  wire g443_n_spl_0;
  wire g443_n_spl_00;
  wire g443_n_spl_1;
  wire g447_p_spl_;
  wire g447_p_spl_0;
  wire g447_p_spl_1;
  wire g447_n_spl_;
  wire g447_n_spl_0;
  wire g447_n_spl_1;
  wire g448_n_spl_;
  wire g448_p_spl_;
  wire G125_n_spl_;
  wire g451_n_spl_;
  wire g451_n_spl_0;
  wire g451_n_spl_1;
  wire g451_p_spl_;
  wire g451_p_spl_0;
  wire g451_p_spl_1;
  wire g452_n_spl_;
  wire g452_n_spl_0;
  wire g452_p_spl_;
  wire g452_p_spl_0;
  wire g450_p_spl_;
  wire g450_p_spl_0;
  wire g450_p_spl_1;
  wire g454_p_spl_;
  wire g454_p_spl_0;
  wire g454_p_spl_1;
  wire g450_n_spl_;
  wire g450_n_spl_0;
  wire g450_n_spl_1;
  wire g454_n_spl_;
  wire g454_n_spl_0;
  wire g454_n_spl_00;
  wire g454_n_spl_1;
  wire G129_n_spl_;
  wire g458_p_spl_;
  wire g458_p_spl_0;
  wire g458_p_spl_1;
  wire g458_n_spl_;
  wire g458_n_spl_0;
  wire g458_n_spl_1;
  wire g459_n_spl_;
  wire g459_n_spl_0;
  wire g459_p_spl_;
  wire g459_p_spl_0;
  wire G131_n_spl_;
  wire g461_p_spl_;
  wire g461_p_spl_0;
  wire g464_n_spl_;
  wire g464_n_spl_0;
  wire g464_n_spl_00;
  wire g464_n_spl_01;
  wire g464_n_spl_1;
  wire g464_n_spl_10;
  wire g461_n_spl_;
  wire g461_n_spl_0;
  wire g464_p_spl_;
  wire g464_p_spl_0;
  wire g464_p_spl_00;
  wire g464_p_spl_01;
  wire g464_p_spl_1;
  wire g464_p_spl_10;
  wire G127_n_spl_;
  wire g468_p_spl_;
  wire g468_p_spl_0;
  wire g468_p_spl_1;
  wire g468_n_spl_;
  wire g468_n_spl_0;
  wire g468_n_spl_1;
  wire g469_n_spl_;
  wire g469_n_spl_0;
  wire g469_p_spl_;
  wire g469_p_spl_0;
  wire g465_p_spl_;
  wire g465_p_spl_0;
  wire g471_p_spl_;
  wire g471_p_spl_0;
  wire g471_p_spl_1;
  wire g465_n_spl_;
  wire g465_n_spl_0;
  wire g471_n_spl_;
  wire g471_n_spl_0;
  wire g471_n_spl_00;
  wire g471_n_spl_1;
  wire g455_p_spl_;
  wire g472_p_spl_;
  wire g455_n_spl_;
  wire g472_n_spl_;
  wire G114_n_spl_;
  wire G114_n_spl_0;
  wire G114_p_spl_;
  wire g476_n_spl_;
  wire g476_n_spl_0;
  wire g476_n_spl_1;
  wire g479_n_spl_;
  wire g479_n_spl_0;
  wire g479_n_spl_00;
  wire g479_n_spl_01;
  wire g479_n_spl_1;
  wire g479_n_spl_10;
  wire g476_p_spl_;
  wire g476_p_spl_0;
  wire g476_p_spl_00;
  wire g476_p_spl_1;
  wire g479_p_spl_;
  wire g479_p_spl_0;
  wire g479_p_spl_00;
  wire g479_p_spl_01;
  wire g479_p_spl_1;
  wire g479_p_spl_10;
  wire g473_p_spl_;
  wire g480_p_spl_;
  wire g480_p_spl_0;
  wire g444_p_spl_;
  wire g444_p_spl_0;
  wire g485_p_spl_;
  wire g488_n_spl_;
  wire g485_n_spl_;
  wire g488_p_spl_;
  wire G132_n_spl_;
  wire G132_n_spl_0;
  wire G132_p_spl_;
  wire G132_p_spl_0;
  wire g494_n_spl_;
  wire g494_p_spl_;
  wire g497_n_spl_;
  wire g500_n_spl_;
  wire g497_p_spl_;
  wire g500_p_spl_;
  wire g509_p_spl_;
  wire g512_n_spl_;
  wire g509_n_spl_;
  wire g512_p_spl_;
  wire G111_n_spl_;
  wire G111_n_spl_0;
  wire G111_p_spl_;
  wire G111_p_spl_0;
  wire g518_n_spl_;
  wire g521_n_spl_;
  wire g518_p_spl_;
  wire g521_p_spl_;
  wire g524_n_spl_;
  wire g527_n_spl_;
  wire g524_p_spl_;
  wire g527_p_spl_;
  wire g535_n_spl_;
  wire g535_n_spl_0;
  wire g535_n_spl_1;
  wire g535_p_spl_;
  wire g535_p_spl_0;
  wire g535_p_spl_1;
  wire g537_n_spl_;
  wire g537_n_spl_0;
  wire g537_n_spl_00;
  wire g537_n_spl_1;
  wire g537_p_spl_;
  wire g537_p_spl_0;
  wire g537_p_spl_00;
  wire g537_p_spl_1;
  wire g539_n_spl_;
  wire g539_n_spl_0;
  wire g539_n_spl_1;
  wire g539_p_spl_;
  wire g539_p_spl_0;
  wire g539_p_spl_1;
  wire g541_p_spl_;
  wire g541_p_spl_0;
  wire g541_p_spl_00;
  wire g541_p_spl_1;
  wire g544_n_spl_;
  wire g544_n_spl_0;
  wire g544_n_spl_1;
  wire g544_p_spl_;
  wire g544_p_spl_0;
  wire g544_p_spl_1;
  wire g545_n_spl_;
  wire g545_p_spl_;
  wire g546_p_spl_;
  wire g546_p_spl_0;
  wire g546_p_spl_1;
  wire G177_p_spl_;
  wire G177_p_spl_0;
  wire G177_p_spl_00;
  wire G177_p_spl_000;
  wire G177_p_spl_0000;
  wire G177_p_spl_0001;
  wire G177_p_spl_001;
  wire G177_p_spl_0010;
  wire G177_p_spl_0011;
  wire G177_p_spl_01;
  wire G177_p_spl_010;
  wire G177_p_spl_0100;
  wire G177_p_spl_0101;
  wire G177_p_spl_011;
  wire G177_p_spl_0110;
  wire G177_p_spl_0111;
  wire G177_p_spl_1;
  wire G177_p_spl_10;
  wire G177_p_spl_100;
  wire G177_p_spl_1000;
  wire G177_p_spl_1001;
  wire G177_p_spl_101;
  wire G177_p_spl_11;
  wire G177_p_spl_110;
  wire G177_p_spl_111;
  wire g553_p_spl_;
  wire G176_p_spl_;
  wire G176_p_spl_0;
  wire G176_p_spl_00;
  wire G176_p_spl_000;
  wire G176_p_spl_0000;
  wire G176_p_spl_00000;
  wire G176_p_spl_00001;
  wire G176_p_spl_0001;
  wire G176_p_spl_001;
  wire G176_p_spl_0010;
  wire G176_p_spl_0011;
  wire G176_p_spl_01;
  wire G176_p_spl_010;
  wire G176_p_spl_0100;
  wire G176_p_spl_0101;
  wire G176_p_spl_011;
  wire G176_p_spl_0110;
  wire G176_p_spl_0111;
  wire G176_p_spl_1;
  wire G176_p_spl_10;
  wire G176_p_spl_100;
  wire G176_p_spl_1000;
  wire G176_p_spl_1001;
  wire G176_p_spl_101;
  wire G176_p_spl_1010;
  wire G176_p_spl_1011;
  wire G176_p_spl_11;
  wire G176_p_spl_110;
  wire G176_p_spl_1100;
  wire G176_p_spl_1101;
  wire G176_p_spl_111;
  wire G176_p_spl_1110;
  wire G176_p_spl_1111;
  wire G177_n_spl_;
  wire G177_n_spl_0;
  wire G177_n_spl_00;
  wire G177_n_spl_000;
  wire G177_n_spl_0000;
  wire G177_n_spl_0001;
  wire G177_n_spl_001;
  wire G177_n_spl_0010;
  wire G177_n_spl_0011;
  wire G177_n_spl_01;
  wire G177_n_spl_010;
  wire G177_n_spl_011;
  wire G177_n_spl_1;
  wire G177_n_spl_10;
  wire G177_n_spl_100;
  wire G177_n_spl_101;
  wire G177_n_spl_11;
  wire G177_n_spl_110;
  wire G177_n_spl_111;
  wire G176_n_spl_;
  wire G176_n_spl_0;
  wire G176_n_spl_00;
  wire G176_n_spl_000;
  wire G176_n_spl_0000;
  wire G176_n_spl_0001;
  wire G176_n_spl_001;
  wire G176_n_spl_0010;
  wire G176_n_spl_0011;
  wire G176_n_spl_01;
  wire G176_n_spl_010;
  wire G176_n_spl_0100;
  wire G176_n_spl_0101;
  wire G176_n_spl_011;
  wire G176_n_spl_1;
  wire G176_n_spl_10;
  wire G176_n_spl_100;
  wire G176_n_spl_101;
  wire G176_n_spl_11;
  wire G176_n_spl_110;
  wire G176_n_spl_111;
  wire g562_n_spl_;
  wire g562_n_spl_0;
  wire G2_p_spl_;
  wire G2_p_spl_0;
  wire G2_p_spl_1;
  wire G2_n_spl_;
  wire G2_n_spl_0;
  wire g570_n_spl_;
  wire g572_p_spl_;
  wire G22_p_spl_;
  wire G173_n_spl_;
  wire G173_n_spl_0;
  wire G173_n_spl_00;
  wire G173_n_spl_000;
  wire G173_n_spl_0000;
  wire G173_n_spl_0001;
  wire G173_n_spl_001;
  wire G173_n_spl_0010;
  wire G173_n_spl_0011;
  wire G173_n_spl_01;
  wire G173_n_spl_010;
  wire G173_n_spl_011;
  wire G173_n_spl_1;
  wire G173_n_spl_10;
  wire G173_n_spl_100;
  wire G173_n_spl_101;
  wire G173_n_spl_11;
  wire G173_n_spl_110;
  wire G173_n_spl_111;
  wire G3_p_spl_;
  wire G173_p_spl_;
  wire G173_p_spl_0;
  wire G173_p_spl_00;
  wire G173_p_spl_000;
  wire G173_p_spl_0000;
  wire G173_p_spl_0001;
  wire G173_p_spl_001;
  wire G173_p_spl_0010;
  wire G173_p_spl_0011;
  wire G173_p_spl_01;
  wire G173_p_spl_010;
  wire G173_p_spl_011;
  wire G173_p_spl_1;
  wire G173_p_spl_10;
  wire G173_p_spl_100;
  wire G173_p_spl_101;
  wire G173_p_spl_11;
  wire G173_p_spl_110;
  wire G173_p_spl_111;
  wire G172_n_spl_;
  wire G172_n_spl_0;
  wire G172_n_spl_00;
  wire G172_n_spl_000;
  wire G172_n_spl_001;
  wire G172_n_spl_01;
  wire G172_n_spl_1;
  wire G172_n_spl_10;
  wire G172_n_spl_11;
  wire g579_p_spl_;
  wire g579_p_spl_0;
  wire g579_p_spl_00;
  wire g579_p_spl_1;
  wire g560_p_spl_;
  wire g560_p_spl_0;
  wire g560_p_spl_00;
  wire g560_p_spl_1;
  wire G172_p_spl_;
  wire G172_p_spl_0;
  wire G172_p_spl_00;
  wire G172_p_spl_000;
  wire G172_p_spl_001;
  wire G172_p_spl_01;
  wire G172_p_spl_1;
  wire G172_p_spl_10;
  wire G172_p_spl_11;
  wire g594_n_spl_;
  wire g594_p_spl_;
  wire g595_n_spl_;
  wire g596_n_spl_;
  wire g596_n_spl_0;
  wire g596_p_spl_;
  wire g596_p_spl_0;
  wire g596_p_spl_1;
  wire g597_p_spl_;
  wire g598_p_spl_;
  wire g598_p_spl_0;
  wire g598_n_spl_;
  wire g598_n_spl_0;
  wire g601_p_spl_;
  wire g610_n_spl_;
  wire g617_p_spl_;
  wire g617_p_spl_0;
  wire g619_n_spl_;
  wire G174_n_spl_;
  wire G174_n_spl_0;
  wire G174_n_spl_00;
  wire G174_n_spl_000;
  wire G174_n_spl_0000;
  wire G174_n_spl_0001;
  wire G174_n_spl_001;
  wire G174_n_spl_0010;
  wire G174_n_spl_0011;
  wire G174_n_spl_01;
  wire G174_n_spl_010;
  wire G174_n_spl_011;
  wire G174_n_spl_1;
  wire G174_n_spl_10;
  wire G174_n_spl_100;
  wire G174_n_spl_101;
  wire G174_n_spl_11;
  wire G174_n_spl_110;
  wire G174_n_spl_111;
  wire G174_p_spl_;
  wire G174_p_spl_0;
  wire G174_p_spl_00;
  wire G174_p_spl_000;
  wire G174_p_spl_0000;
  wire G174_p_spl_0001;
  wire G174_p_spl_001;
  wire G174_p_spl_0010;
  wire G174_p_spl_0011;
  wire G174_p_spl_01;
  wire G174_p_spl_010;
  wire G174_p_spl_011;
  wire G174_p_spl_1;
  wire G174_p_spl_10;
  wire G174_p_spl_100;
  wire G174_p_spl_101;
  wire G174_p_spl_11;
  wire G174_p_spl_110;
  wire G174_p_spl_111;
  wire G175_n_spl_;
  wire G175_n_spl_0;
  wire G175_n_spl_00;
  wire G175_n_spl_000;
  wire G175_n_spl_001;
  wire G175_n_spl_01;
  wire G175_n_spl_1;
  wire G175_n_spl_10;
  wire G175_n_spl_11;
  wire G175_p_spl_;
  wire G175_p_spl_0;
  wire G175_p_spl_00;
  wire G175_p_spl_000;
  wire G175_p_spl_001;
  wire G175_p_spl_01;
  wire G175_p_spl_1;
  wire G175_p_spl_10;
  wire G175_p_spl_11;
  wire g638_p_spl_;
  wire g639_p_spl_;
  wire g643_n_spl_;
  wire g652_n_spl_;
  wire g659_p_spl_;
  wire g660_p_spl_;
  wire g664_n_spl_;
  wire g673_n_spl_;
  wire g581_n_spl_;
  wire g581_n_spl_0;
  wire g581_n_spl_00;
  wire g581_n_spl_01;
  wire g581_n_spl_1;
  wire g581_n_spl_10;
  wire g581_n_spl_11;
  wire g681_p_spl_;
  wire g581_p_spl_;
  wire g581_p_spl_0;
  wire g581_p_spl_00;
  wire g581_p_spl_01;
  wire g581_p_spl_1;
  wire g681_n_spl_;
  wire g687_n_spl_;
  wire g687_p_spl_;
  wire g693_n_spl_;
  wire g696_n_spl_;
  wire g693_p_spl_;
  wire g696_p_spl_;
  wire g690_p_spl_;
  wire g699_n_spl_;
  wire g690_n_spl_;
  wire g699_p_spl_;
  wire g708_p_spl_;
  wire g711_n_spl_;
  wire g708_n_spl_;
  wire g711_p_spl_;
  wire g717_n_spl_;
  wire g717_p_spl_;
  wire g720_p_spl_;
  wire g723_n_spl_;
  wire g720_n_spl_;
  wire g723_p_spl_;
  wire g726_n_spl_;
  wire g729_n_spl_;
  wire g726_p_spl_;
  wire g729_p_spl_;
  wire g430_p_spl_;
  wire g430_p_spl_0;
  wire g541_n_spl_;
  wire g541_n_spl_0;
  wire g541_n_spl_1;
  wire g737_p_spl_;
  wire g737_p_spl_0;
  wire g737_p_spl_00;
  wire g737_p_spl_1;
  wire g737_n_spl_;
  wire g737_n_spl_0;
  wire g737_n_spl_00;
  wire g737_n_spl_1;
  wire g743_p_spl_;
  wire g747_p_spl_;
  wire g389_p_spl_;
  wire g546_n_spl_;
  wire g546_n_spl_0;
  wire g395_p_spl_;
  wire g395_p_spl_0;
  wire g395_p_spl_00;
  wire g395_p_spl_1;
  wire g755_p_spl_;
  wire g760_p_spl_;
  wire g774_p_spl_;
  wire g774_p_spl_0;
  wire g774_p_spl_00;
  wire g774_p_spl_01;
  wire g774_p_spl_1;
  wire g774_n_spl_;
  wire g774_n_spl_0;
  wire g774_n_spl_00;
  wire g774_n_spl_01;
  wire g774_n_spl_1;
  wire g777_p_spl_;
  wire g444_n_spl_;
  wire g780_p_spl_;
  wire g780_p_spl_0;
  wire g780_p_spl_1;
  wire g780_n_spl_;
  wire g780_n_spl_0;
  wire g780_n_spl_1;
  wire g785_p_spl_;
  wire g791_p_spl_;
  wire G81_p_spl_;
  wire G158_n_spl_;
  wire G158_n_spl_0;
  wire G158_n_spl_00;
  wire G158_n_spl_000;
  wire G158_n_spl_0000;
  wire G158_n_spl_0001;
  wire G158_n_spl_001;
  wire G158_n_spl_0010;
  wire G158_n_spl_0011;
  wire G158_n_spl_01;
  wire G158_n_spl_010;
  wire G158_n_spl_011;
  wire G158_n_spl_1;
  wire G158_n_spl_10;
  wire G158_n_spl_100;
  wire G158_n_spl_101;
  wire G158_n_spl_11;
  wire G158_n_spl_110;
  wire G158_n_spl_111;
  wire G80_p_spl_;
  wire G158_p_spl_;
  wire G158_p_spl_0;
  wire G158_p_spl_00;
  wire G158_p_spl_000;
  wire G158_p_spl_0000;
  wire G158_p_spl_0001;
  wire G158_p_spl_001;
  wire G158_p_spl_0010;
  wire G158_p_spl_0011;
  wire G158_p_spl_01;
  wire G158_p_spl_010;
  wire G158_p_spl_011;
  wire G158_p_spl_1;
  wire G158_p_spl_10;
  wire G158_p_spl_100;
  wire G158_p_spl_101;
  wire G158_p_spl_11;
  wire G158_p_spl_110;
  wire G158_p_spl_111;
  wire G159_n_spl_;
  wire G159_n_spl_0;
  wire G159_n_spl_00;
  wire G159_n_spl_000;
  wire G159_n_spl_001;
  wire G159_n_spl_01;
  wire G159_n_spl_1;
  wire G159_n_spl_10;
  wire G159_n_spl_11;
  wire G159_p_spl_;
  wire G159_p_spl_0;
  wire G159_p_spl_00;
  wire G159_p_spl_000;
  wire G159_p_spl_001;
  wire G159_p_spl_01;
  wire G159_p_spl_1;
  wire G159_p_spl_10;
  wire G159_p_spl_11;
  wire G64_p_spl_;
  wire G64_p_spl_0;
  wire G64_p_spl_00;
  wire G64_p_spl_000;
  wire G64_p_spl_0000;
  wire G64_p_spl_0001;
  wire G64_p_spl_001;
  wire G64_p_spl_0010;
  wire G64_p_spl_01;
  wire G64_p_spl_010;
  wire G64_p_spl_011;
  wire G64_p_spl_1;
  wire G64_p_spl_10;
  wire G64_p_spl_100;
  wire G64_p_spl_101;
  wire G64_p_spl_11;
  wire G64_p_spl_110;
  wire G64_p_spl_111;
  wire G160_n_spl_;
  wire G160_n_spl_0;
  wire G160_n_spl_00;
  wire G160_n_spl_000;
  wire G160_n_spl_0000;
  wire G160_n_spl_0001;
  wire G160_n_spl_001;
  wire G160_n_spl_0010;
  wire G160_n_spl_0011;
  wire G160_n_spl_01;
  wire G160_n_spl_010;
  wire G160_n_spl_011;
  wire G160_n_spl_1;
  wire G160_n_spl_10;
  wire G160_n_spl_100;
  wire G160_n_spl_101;
  wire G160_n_spl_11;
  wire G160_n_spl_110;
  wire G160_n_spl_111;
  wire G160_p_spl_;
  wire G160_p_spl_0;
  wire G160_p_spl_00;
  wire G160_p_spl_000;
  wire G160_p_spl_0000;
  wire G160_p_spl_0001;
  wire G160_p_spl_001;
  wire G160_p_spl_0010;
  wire G160_p_spl_0011;
  wire G160_p_spl_01;
  wire G160_p_spl_010;
  wire G160_p_spl_011;
  wire G160_p_spl_1;
  wire G160_p_spl_10;
  wire G160_p_spl_100;
  wire G160_p_spl_101;
  wire G160_p_spl_11;
  wire G160_p_spl_110;
  wire G160_p_spl_111;
  wire G161_n_spl_;
  wire G161_n_spl_0;
  wire G161_n_spl_00;
  wire G161_n_spl_000;
  wire G161_n_spl_001;
  wire G161_n_spl_01;
  wire G161_n_spl_1;
  wire G161_n_spl_10;
  wire G161_n_spl_11;
  wire G161_p_spl_;
  wire G161_p_spl_0;
  wire G161_p_spl_00;
  wire G161_p_spl_000;
  wire G161_p_spl_001;
  wire G161_p_spl_01;
  wire G161_p_spl_1;
  wire G161_p_spl_10;
  wire G161_p_spl_11;
  wire G14_p_spl_;
  wire G16_p_spl_;
  wire g647_n_spl_;
  wire g647_n_spl_0;
  wire g647_n_spl_00;
  wire g647_n_spl_1;
  wire g605_n_spl_;
  wire g605_n_spl_0;
  wire g605_n_spl_00;
  wire g605_n_spl_1;
  wire G6_p_spl_;
  wire G27_p_spl_;
  wire g656_n_spl_;
  wire g656_n_spl_0;
  wire g656_n_spl_00;
  wire g656_n_spl_1;
  wire g614_n_spl_;
  wire g614_n_spl_0;
  wire g614_n_spl_00;
  wire g614_n_spl_1;
  wire G5_p_spl_;
  wire G26_p_spl_;
  wire g669_n_spl_;
  wire g669_n_spl_0;
  wire g669_n_spl_00;
  wire g669_n_spl_1;
  wire g624_n_spl_;
  wire g624_n_spl_0;
  wire g624_n_spl_00;
  wire g624_n_spl_1;
  wire G25_p_spl_;
  wire G24_p_spl_;
  wire g678_n_spl_;
  wire g678_n_spl_0;
  wire g678_n_spl_00;
  wire g678_n_spl_1;
  wire g569_p_spl_;
  wire g569_p_spl_0;
  wire g569_p_spl_00;
  wire g569_p_spl_1;
  wire G76_p_spl_;
  wire G86_p_spl_;
  wire G72_p_spl_;
  wire G82_p_spl_;
  wire G70_p_spl_;
  wire G71_p_spl_;
  wire G68_p_spl_;
  wire G69_p_spl_;
  wire G171_p_spl_;
  wire G54_p_spl_;
  wire G171_n_spl_;
  wire G61_n_spl_;
  wire G61_p_spl_;
  wire g975_p_spl_;
  wire G99_n_spl_;
  wire g533_n_spl_;
  wire g735_n_spl_;
  wire G155_n_spl_;
  wire g184_n_spl_;
  wire g179_n_spl_;
  wire g705_n_spl_;
  wire g506_n_spl_;
  wire g1025_n_spl_;
  wire g1025_n_spl_0;
  wire g1025_n_spl_00;
  wire g1025_n_spl_1;
  wire g990_p_spl_;
  wire g990_p_spl_0;
  wire g990_p_spl_00;
  wire g990_p_spl_1;
  wire G41_p_spl_;
  wire G42_p_spl_;
  wire G18_p_spl_;
  wire G17_p_spl_;
  wire g1032_n_spl_;
  wire g1032_n_spl_0;
  wire g1032_n_spl_00;
  wire g1032_n_spl_1;
  wire g997_n_spl_;
  wire g997_n_spl_0;
  wire g997_n_spl_00;
  wire g997_n_spl_1;
  wire G40_p_spl_;
  wire G39_p_spl_;
  wire g1039_n_spl_;
  wire g1039_n_spl_0;
  wire g1039_n_spl_00;
  wire g1039_n_spl_1;
  wire g1004_n_spl_;
  wire g1004_n_spl_0;
  wire g1004_n_spl_00;
  wire g1004_n_spl_1;
  wire G15_p_spl_;
  wire G36_p_spl_;
  wire g1046_n_spl_;
  wire g1046_n_spl_0;
  wire g1046_n_spl_00;
  wire g1046_n_spl_1;
  wire g1011_n_spl_;
  wire g1011_n_spl_0;
  wire g1011_n_spl_00;
  wire g1011_n_spl_1;
  wire G77_p_spl_;
  wire G87_p_spl_;
  wire G75_p_spl_;
  wire G85_p_spl_;
  wire G74_p_spl_;
  wire G84_p_spl_;
  wire G73_p_spl_;
  wire G83_p_spl_;
  wire g1200_p_spl_;
  wire g1202_n_spl_;
  wire g1200_n_spl_;
  wire g1202_p_spl_;
  wire g1214_n_spl_;
  wire g1223_p_spl_;
  wire g1214_p_spl_;
  wire g1223_n_spl_;
  wire g1229_n_spl_;
  wire g1238_p_spl_;
  wire g1229_p_spl_;
  wire g1238_n_spl_;
  wire g1241_p_spl_;
  wire g245_p_spl_;
  wire g1241_n_spl_;
  wire g1226_p_spl_;
  wire g1244_n_spl_;
  wire g1226_n_spl_;
  wire g1244_p_spl_;
  wire g1254_n_spl_;
  wire g617_n_spl_;
  wire g1254_p_spl_;
  wire g1257_p_spl_;
  wire g1257_n_spl_;
  wire G162_n_spl_;
  wire G162_p_spl_;
  wire g1260_p_spl_;
  wire g1263_p_spl_;
  wire g1260_n_spl_;
  wire g1263_n_spl_;
  wire g1268_n_spl_;
  wire g1268_p_spl_;
  wire g1266_n_spl_;
  wire g1271_n_spl_;
  wire g1266_p_spl_;
  wire g1271_p_spl_;
  wire g1275_n_spl_;
  wire g1275_p_spl_;
  wire g1278_p_spl_;
  wire g1278_n_spl_;
  wire g1281_p_spl_;
  wire g1281_n_spl_;
  wire g1282_n_spl_;
  wire g1282_p_spl_;
  wire g1284_n_spl_;
  wire g1284_p_spl_;
  wire g1288_n_spl_;
  wire g1288_p_spl_;
  wire g1299_p_spl_;
  wire g1299_n_spl_;
  wire g1308_n_spl_;
  wire g1320_n_spl_;
  wire g1329_p_spl_;
  wire g1320_p_spl_;
  wire g1329_n_spl_;
  wire g1341_n_spl_;
  wire g317_p_spl_;
  wire g1341_p_spl_;
  wire g1332_n_spl_;
  wire g1344_p_spl_;
  wire g1332_p_spl_;
  wire g1344_n_spl_;
  wire g1356_n_spl_;
  wire g1365_p_spl_;
  wire g1356_p_spl_;
  wire g1365_n_spl_;
  wire g1377_n_spl_;
  wire g1386_p_spl_;
  wire g1377_p_spl_;
  wire g1386_n_spl_;
  wire g1389_p_spl_;
  wire g1398_n_spl_;
  wire g1389_n_spl_;
  wire g1398_p_spl_;
  wire g1368_p_spl_;
  wire g1401_n_spl_;
  wire g1368_n_spl_;
  wire g1401_p_spl_;
  wire g1409_n_spl_;
  wire g1412_n_spl_;
  wire g1409_p_spl_;
  wire g1412_p_spl_;
  wire g1415_p_spl_;
  wire g1415_n_spl_;
  wire g1416_n_spl_;
  wire g1416_p_spl_;
  wire g1420_p_spl_;
  wire g1420_n_spl_;
  wire g1423_p_spl_;
  wire g1423_n_spl_;
  wire g1426_p_spl_;
  wire g1426_n_spl_;
  wire g1432_p_spl_;
  wire g1432_n_spl_;
  wire g1435_p_spl_;
  wire g1435_n_spl_;
  wire g1438_p_spl_;
  wire g1438_n_spl_;
  wire g1441_n_spl_;
  wire g1441_p_spl_;
  wire g1430_n_spl_;
  wire g1430_p_spl_;
  wire G157_n_spl_;
  wire G157_n_spl_0;
  wire G157_n_spl_1;
  wire G157_p_spl_;
  wire G157_p_spl_0;
  wire G157_p_spl_1;
  wire g1453_n_spl_;
  wire g1453_p_spl_;
  wire g1458_n_spl_;
  wire g1458_n_spl_0;
  wire g1458_n_spl_1;
  wire g1458_p_spl_;
  wire g1458_p_spl_0;
  wire g1458_p_spl_1;
  wire g1456_n_spl_;
  wire g1461_p_spl_;
  wire g1456_p_spl_;
  wire g1461_n_spl_;
  wire g1464_n_spl_;
  wire g1464_p_spl_;
  wire g1471_n_spl_;
  wire g1471_p_spl_;
  wire g1470_n_spl_;
  wire g1474_p_spl_;
  wire g1470_p_spl_;
  wire g1474_n_spl_;
  wire g1469_n_spl_;
  wire g1477_p_spl_;
  wire g1469_p_spl_;
  wire g1477_n_spl_;
  wire g1480_n_spl_;
  wire g1483_p_spl_;
  wire g1480_p_spl_;
  wire g1483_n_spl_;
  wire g1488_p_spl_;
  wire g1488_n_spl_;
  wire g1491_n_spl_;
  wire g1491_p_spl_;
  wire g1500_n_spl_;
  wire G23_n_spl_;
  wire G4_n_spl_;
  wire g1509_p_spl_;
  wire g1509_p_spl_0;
  wire g1509_p_spl_1;
  wire g1512_p_spl_;
  wire g1512_p_spl_0;
  wire g1512_p_spl_1;
  wire G79_n_spl_;
  wire G78_n_spl_;
  wire G64_n_spl_;
  wire G151_n_spl_;
  wire G151_n_spl_0;
  wire G152_p_spl_;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire G1_n_spl_1;
  wire g194_n_spl_;
  wire g431_n_spl_;
  wire g482_p_spl_;
  wire g549_p_spl_;
  wire g550_n_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  buf

  (
    G42_p,
    G42
  );


  not

  (
    G42_n,
    G42
  );


  buf

  (
    G43_p,
    G43
  );


  not

  (
    G43_n,
    G43
  );


  buf

  (
    G44_p,
    G44
  );


  not

  (
    G44_n,
    G44
  );


  buf

  (
    G45_p,
    G45
  );


  not

  (
    G45_n,
    G45
  );


  buf

  (
    G46_p,
    G46
  );


  not

  (
    G46_n,
    G46
  );


  buf

  (
    G47_p,
    G47
  );


  not

  (
    G47_n,
    G47
  );


  buf

  (
    G48_p,
    G48
  );


  not

  (
    G48_n,
    G48
  );


  buf

  (
    G49_p,
    G49
  );


  not

  (
    G49_n,
    G49
  );


  buf

  (
    G50_p,
    G50
  );


  not

  (
    G50_n,
    G50
  );


  buf

  (
    G51_p,
    G51
  );


  not

  (
    G51_n,
    G51
  );


  buf

  (
    G52_p,
    G52
  );


  not

  (
    G52_n,
    G52
  );


  buf

  (
    G53_p,
    G53
  );


  not

  (
    G53_n,
    G53
  );


  buf

  (
    G54_p,
    G54
  );


  not

  (
    G54_n,
    G54
  );


  buf

  (
    G55_p,
    G55
  );


  not

  (
    G55_n,
    G55
  );


  buf

  (
    G56_p,
    G56
  );


  not

  (
    G56_n,
    G56
  );


  buf

  (
    G57_p,
    G57
  );


  not

  (
    G57_n,
    G57
  );


  buf

  (
    G58_p,
    G58
  );


  not

  (
    G58_n,
    G58
  );


  buf

  (
    G59_p,
    G59
  );


  not

  (
    G59_n,
    G59
  );


  buf

  (
    G60_p,
    G60
  );


  not

  (
    G60_n,
    G60
  );


  buf

  (
    G61_p,
    G61
  );


  not

  (
    G61_n,
    G61
  );


  buf

  (
    G62_p,
    G62
  );


  not

  (
    G62_n,
    G62
  );


  buf

  (
    G63_p,
    G63
  );


  not

  (
    G63_n,
    G63
  );


  buf

  (
    G64_p,
    G64
  );


  not

  (
    G64_n,
    G64
  );


  buf

  (
    G65_p,
    G65
  );


  not

  (
    G65_n,
    G65
  );


  buf

  (
    G66_p,
    G66
  );


  not

  (
    G66_n,
    G66
  );


  buf

  (
    G67_p,
    G67
  );


  not

  (
    G67_n,
    G67
  );


  buf

  (
    G68_p,
    G68
  );


  not

  (
    G68_n,
    G68
  );


  buf

  (
    G69_p,
    G69
  );


  not

  (
    G69_n,
    G69
  );


  buf

  (
    G70_p,
    G70
  );


  not

  (
    G70_n,
    G70
  );


  buf

  (
    G71_p,
    G71
  );


  not

  (
    G71_n,
    G71
  );


  buf

  (
    G72_p,
    G72
  );


  not

  (
    G72_n,
    G72
  );


  buf

  (
    G73_p,
    G73
  );


  not

  (
    G73_n,
    G73
  );


  buf

  (
    G74_p,
    G74
  );


  not

  (
    G74_n,
    G74
  );


  buf

  (
    G75_p,
    G75
  );


  not

  (
    G75_n,
    G75
  );


  buf

  (
    G76_p,
    G76
  );


  not

  (
    G76_n,
    G76
  );


  buf

  (
    G77_p,
    G77
  );


  not

  (
    G77_n,
    G77
  );


  buf

  (
    G78_p,
    G78
  );


  not

  (
    G78_n,
    G78
  );


  buf

  (
    G79_p,
    G79
  );


  not

  (
    G79_n,
    G79
  );


  buf

  (
    G80_p,
    G80
  );


  not

  (
    G80_n,
    G80
  );


  buf

  (
    G81_p,
    G81
  );


  not

  (
    G81_n,
    G81
  );


  buf

  (
    G82_p,
    G82
  );


  not

  (
    G82_n,
    G82
  );


  buf

  (
    G83_p,
    G83
  );


  not

  (
    G83_n,
    G83
  );


  buf

  (
    G84_p,
    G84
  );


  not

  (
    G84_n,
    G84
  );


  buf

  (
    G85_p,
    G85
  );


  not

  (
    G85_n,
    G85
  );


  buf

  (
    G86_p,
    G86
  );


  not

  (
    G86_n,
    G86
  );


  buf

  (
    G87_p,
    G87
  );


  not

  (
    G87_n,
    G87
  );


  buf

  (
    G88_p,
    G88
  );


  not

  (
    G88_n,
    G88
  );


  buf

  (
    G89_p,
    G89
  );


  not

  (
    G89_n,
    G89
  );


  buf

  (
    G90_p,
    G90
  );


  not

  (
    G90_n,
    G90
  );


  buf

  (
    G91_p,
    G91
  );


  not

  (
    G91_n,
    G91
  );


  buf

  (
    G92_p,
    G92
  );


  not

  (
    G92_n,
    G92
  );


  buf

  (
    G93_p,
    G93
  );


  not

  (
    G93_n,
    G93
  );


  buf

  (
    G94_p,
    G94
  );


  not

  (
    G94_n,
    G94
  );


  buf

  (
    G95_p,
    G95
  );


  not

  (
    G95_n,
    G95
  );


  buf

  (
    G96_p,
    G96
  );


  not

  (
    G96_n,
    G96
  );


  buf

  (
    G97_p,
    G97
  );


  not

  (
    G97_n,
    G97
  );


  buf

  (
    G98_p,
    G98
  );


  not

  (
    G98_n,
    G98
  );


  buf

  (
    G99_p,
    G99
  );


  not

  (
    G99_n,
    G99
  );


  buf

  (
    G100_p,
    G100
  );


  not

  (
    G100_n,
    G100
  );


  buf

  (
    G101_p,
    G101
  );


  not

  (
    G101_n,
    G101
  );


  buf

  (
    G102_p,
    G102
  );


  not

  (
    G102_n,
    G102
  );


  buf

  (
    G103_p,
    G103
  );


  not

  (
    G103_n,
    G103
  );


  buf

  (
    G104_p,
    G104
  );


  not

  (
    G104_n,
    G104
  );


  buf

  (
    G105_p,
    G105
  );


  not

  (
    G105_n,
    G105
  );


  buf

  (
    G106_p,
    G106
  );


  not

  (
    G106_n,
    G106
  );


  buf

  (
    G107_p,
    G107
  );


  not

  (
    G107_n,
    G107
  );


  buf

  (
    G108_p,
    G108
  );


  not

  (
    G108_n,
    G108
  );


  buf

  (
    G109_p,
    G109
  );


  not

  (
    G109_n,
    G109
  );


  buf

  (
    G110_p,
    G110
  );


  not

  (
    G110_n,
    G110
  );


  buf

  (
    G111_p,
    G111
  );


  not

  (
    G111_n,
    G111
  );


  buf

  (
    G112_p,
    G112
  );


  not

  (
    G112_n,
    G112
  );


  buf

  (
    G113_p,
    G113
  );


  not

  (
    G113_n,
    G113
  );


  buf

  (
    G114_p,
    G114
  );


  not

  (
    G114_n,
    G114
  );


  buf

  (
    G115_p,
    G115
  );


  not

  (
    G115_n,
    G115
  );


  buf

  (
    G116_p,
    G116
  );


  not

  (
    G116_n,
    G116
  );


  buf

  (
    G117_p,
    G117
  );


  not

  (
    G117_n,
    G117
  );


  buf

  (
    G118_p,
    G118
  );


  not

  (
    G118_n,
    G118
  );


  buf

  (
    G119_p,
    G119
  );


  not

  (
    G119_n,
    G119
  );


  buf

  (
    G120_p,
    G120
  );


  not

  (
    G120_n,
    G120
  );


  buf

  (
    G121_p,
    G121
  );


  not

  (
    G121_n,
    G121
  );


  buf

  (
    G122_p,
    G122
  );


  not

  (
    G122_n,
    G122
  );


  buf

  (
    G123_p,
    G123
  );


  not

  (
    G123_n,
    G123
  );


  buf

  (
    G124_p,
    G124
  );


  not

  (
    G124_n,
    G124
  );


  buf

  (
    G125_p,
    G125
  );


  not

  (
    G125_n,
    G125
  );


  buf

  (
    G126_p,
    G126
  );


  not

  (
    G126_n,
    G126
  );


  buf

  (
    G127_p,
    G127
  );


  not

  (
    G127_n,
    G127
  );


  buf

  (
    G128_p,
    G128
  );


  not

  (
    G128_n,
    G128
  );


  buf

  (
    G129_p,
    G129
  );


  not

  (
    G129_n,
    G129
  );


  buf

  (
    G130_p,
    G130
  );


  not

  (
    G130_n,
    G130
  );


  buf

  (
    G131_p,
    G131
  );


  not

  (
    G131_n,
    G131
  );


  buf

  (
    G132_p,
    G132
  );


  not

  (
    G132_n,
    G132
  );


  buf

  (
    G133_p,
    G133
  );


  not

  (
    G133_n,
    G133
  );


  buf

  (
    G134_p,
    G134
  );


  not

  (
    G134_n,
    G134
  );


  buf

  (
    G135_p,
    G135
  );


  not

  (
    G135_n,
    G135
  );


  buf

  (
    G136_p,
    G136
  );


  not

  (
    G136_n,
    G136
  );


  buf

  (
    G137_p,
    G137
  );


  not

  (
    G137_n,
    G137
  );


  buf

  (
    G138_p,
    G138
  );


  not

  (
    G138_n,
    G138
  );


  buf

  (
    G139_p,
    G139
  );


  not

  (
    G139_n,
    G139
  );


  buf

  (
    G140_p,
    G140
  );


  not

  (
    G140_n,
    G140
  );


  buf

  (
    G141_p,
    G141
  );


  not

  (
    G141_n,
    G141
  );


  buf

  (
    G142_p,
    G142
  );


  not

  (
    G142_n,
    G142
  );


  buf

  (
    G143_p,
    G143
  );


  not

  (
    G143_n,
    G143
  );


  buf

  (
    G144_p,
    G144
  );


  not

  (
    G144_n,
    G144
  );


  buf

  (
    G145_p,
    G145
  );


  not

  (
    G145_n,
    G145
  );


  buf

  (
    G146_p,
    G146
  );


  not

  (
    G146_n,
    G146
  );


  buf

  (
    G147_p,
    G147
  );


  not

  (
    G147_n,
    G147
  );


  buf

  (
    G148_p,
    G148
  );


  not

  (
    G148_n,
    G148
  );


  buf

  (
    G149_p,
    G149
  );


  not

  (
    G149_n,
    G149
  );


  buf

  (
    G150_p,
    G150
  );


  not

  (
    G150_n,
    G150
  );


  buf

  (
    G151_p,
    G151
  );


  not

  (
    G151_n,
    G151
  );


  buf

  (
    G152_p,
    G152
  );


  not

  (
    G152_n,
    G152
  );


  buf

  (
    G153_p,
    G153
  );


  not

  (
    G153_n,
    G153
  );


  buf

  (
    G154_p,
    G154
  );


  not

  (
    G154_n,
    G154
  );


  buf

  (
    G155_p,
    G155
  );


  not

  (
    G155_n,
    G155
  );


  buf

  (
    G156_p,
    G156
  );


  not

  (
    G156_n,
    G156
  );


  buf

  (
    G157_p,
    G157
  );


  not

  (
    G157_n,
    G157
  );


  buf

  (
    G158_p,
    G158
  );


  not

  (
    G158_n,
    G158
  );


  buf

  (
    G159_p,
    G159
  );


  not

  (
    G159_n,
    G159
  );


  buf

  (
    G160_p,
    G160
  );


  not

  (
    G160_n,
    G160
  );


  buf

  (
    G161_p,
    G161
  );


  not

  (
    G161_n,
    G161
  );


  buf

  (
    G162_p,
    G162
  );


  not

  (
    G162_n,
    G162
  );


  buf

  (
    G163_p,
    G163
  );


  not

  (
    G163_n,
    G163
  );


  buf

  (
    G164_p,
    G164
  );


  not

  (
    G164_n,
    G164
  );


  buf

  (
    G165_p,
    G165
  );


  not

  (
    G165_n,
    G165
  );


  buf

  (
    G166_p,
    G166
  );


  not

  (
    G166_n,
    G166
  );


  buf

  (
    G167_p,
    G167
  );


  not

  (
    G167_n,
    G167
  );


  buf

  (
    G168_p,
    G168
  );


  not

  (
    G168_n,
    G168
  );


  buf

  (
    G169_p,
    G169
  );


  not

  (
    G169_n,
    G169
  );


  buf

  (
    G170_p,
    G170
  );


  not

  (
    G170_n,
    G170
  );


  buf

  (
    G171_p,
    G171
  );


  not

  (
    G171_n,
    G171
  );


  buf

  (
    G172_p,
    G172
  );


  not

  (
    G172_n,
    G172
  );


  buf

  (
    G173_p,
    G173
  );


  not

  (
    G173_n,
    G173
  );


  buf

  (
    G174_p,
    G174
  );


  not

  (
    G174_n,
    G174
  );


  buf

  (
    G175_p,
    G175
  );


  not

  (
    G175_n,
    G175
  );


  buf

  (
    G176_p,
    G176
  );


  not

  (
    G176_n,
    G176
  );


  buf

  (
    G177_p,
    G177
  );


  not

  (
    G177_n,
    G177
  );


  buf

  (
    G178_p,
    G178
  );


  not

  (
    G178_n,
    G178
  );


  or

  (
    g179_n,
    G153_n_spl_,
    G156_n_spl_
  );


  and

  (
    g180_p,
    G66_p_spl_00,
    G67_p
  );


  and

  (
    g181_p,
    G1_p_spl_,
    G134_p
  );


  and

  (
    g182_p,
    G63_p,
    G165_n_spl_
  );


  or

  (
    g183_n,
    G11_n_spl_,
    G164_p
  );


  or

  (
    g184_n,
    G136_n,
    G154_n
  );


  or

  (
    g185_n,
    G11_n_spl_,
    G12_n
  );


  or

  (
    g186_n,
    G65_n,
    g185_n_spl_000
  );


  or

  (
    g187_n,
    G34_n,
    G163_n_spl_00
  );


  or

  (
    g188_n,
    G33_n,
    G163_p_spl_00
  );


  and

  (
    g189_p,
    g187_n,
    g188_n
  );


  or

  (
    g190_n,
    g185_n_spl_000,
    g189_p
  );


  or

  (
    g191_n,
    G13_n,
    G163_n_spl_00
  );


  or

  (
    g192_n,
    G35_n,
    G163_p_spl_00
  );


  and

  (
    g193_p,
    g191_n,
    g192_n
  );


  or

  (
    g194_n,
    g185_n_spl_00,
    g193_p
  );


  or

  (
    g195_n,
    G32_n,
    g185_n_spl_01
  );


  and

  (
    g196_p,
    G8_p,
    G163_p_spl_01
  );


  and

  (
    g197_p,
    G9_p,
    G163_n_spl_01
  );


  or

  (
    g198_n,
    g185_n_spl_01,
    g197_p
  );


  or

  (
    g199_n,
    g196_p,
    g198_n
  );


  and

  (
    g200_p,
    G66_p_spl_00,
    g199_n
  );


  and

  (
    g201_p,
    G10_p,
    G163_p_spl_01
  );


  and

  (
    g202_p,
    G30_p,
    G163_n_spl_01
  );


  or

  (
    g203_n,
    g185_n_spl_10,
    g202_p
  );


  or

  (
    g204_n,
    g201_p,
    g203_n
  );


  and

  (
    g205_p,
    G66_p_spl_01,
    g204_n
  );


  and

  (
    g206_p,
    G28_p,
    G163_p_spl_1
  );


  and

  (
    g207_p,
    G7_p,
    G163_n_spl_1
  );


  or

  (
    g208_n,
    g185_n_spl_10,
    g207_p
  );


  or

  (
    g209_n,
    g206_p,
    g208_n
  );


  and

  (
    g210_p,
    G66_p_spl_01,
    g209_n
  );


  and

  (
    g211_p,
    G31_p,
    G163_p_spl_1
  );


  and

  (
    g212_p,
    G29_p,
    G163_n_spl_1
  );


  or

  (
    g213_n,
    g185_n_spl_11,
    g212_p
  );


  or

  (
    g214_n,
    g211_p,
    g213_n
  );


  and

  (
    g215_p,
    G66_p_spl_1,
    g214_n
  );


  and

  (
    g216_p,
    G128_p_spl_000,
    G168_p_spl_000
  );


  and

  (
    g217_p,
    G128_n_spl_000,
    G169_p_spl_000
  );


  or

  (
    g218_n,
    g216_p,
    g217_p
  );


  and

  (
    g219_p,
    G150_p_spl_00,
    g218_n
  );


  and

  (
    g220_p,
    G128_p_spl_000,
    G167_n_spl_000
  );


  and

  (
    g221_p,
    G128_n_spl_000,
    G166_n_spl_000
  );


  or

  (
    g222_n,
    g220_p,
    g221_p
  );


  and

  (
    g223_p,
    G150_n_spl_00,
    g222_n
  );


  or

  (
    g224_n,
    g219_p,
    g223_p
  );


  and

  (
    g225_p,
    G126_p_spl_000,
    G168_p_spl_000
  );


  and

  (
    g226_p,
    G126_n_spl_000,
    G169_p_spl_000
  );


  or

  (
    g227_n,
    g225_p,
    g226_p
  );


  and

  (
    g228_p,
    G149_p_spl_00,
    g227_n
  );


  and

  (
    g229_p,
    G126_p_spl_000,
    G167_n_spl_000
  );


  and

  (
    g230_p,
    G126_n_spl_000,
    G166_n_spl_000
  );


  or

  (
    g231_n,
    g229_p,
    g230_p
  );


  and

  (
    g232_p,
    G149_n_spl_00,
    g231_n
  );


  or

  (
    g233_n,
    g228_p,
    g232_p
  );


  or

  (
    g234_n,
    g224_n_spl_,
    g233_n_spl_
  );


  and

  (
    g235_p,
    G102_p_spl_000,
    G113_p_spl_00
  );


  or

  (
    g235_n,
    G102_n_spl_000,
    G113_n_spl_00
  );


  and

  (
    g236_p,
    G98_p_spl_000,
    G113_n_spl_00
  );


  or

  (
    g236_n,
    G98_n_spl_000,
    G113_p_spl_00
  );


  and

  (
    g237_p,
    g235_n,
    g236_n
  );


  or

  (
    g237_n,
    g235_p,
    g236_p
  );


  and

  (
    g238_p,
    G101_p_spl_000,
    G115_p_spl_00
  );


  or

  (
    g238_n,
    G101_n_spl_000,
    G115_n_spl_00
  );


  and

  (
    g239_p,
    G100_p_spl_0000,
    G115_n_spl_00
  );


  or

  (
    g239_n,
    G100_n_spl_0000,
    G115_p_spl_00
  );


  and

  (
    g240_p,
    g238_n,
    g239_n
  );


  or

  (
    g240_n,
    g238_p,
    g239_p
  );


  and

  (
    g241_p,
    g237_n_spl_0,
    g240_p_spl_
  );


  or

  (
    g241_n,
    g237_p_spl_,
    g240_n_spl_0
  );


  or

  (
    g242_n,
    g234_n,
    g241_n_spl_
  );


  and

  (
    g243_p,
    G101_p_spl_000,
    G130_p_spl_00
  );


  or

  (
    g243_n,
    G101_n_spl_000,
    G130_n_spl_00
  );


  and

  (
    g244_p,
    G100_p_spl_0000,
    G130_n_spl_00
  );


  or

  (
    g244_n,
    G100_n_spl_0000,
    G130_p_spl_00
  );


  and

  (
    g245_p,
    g243_n,
    g244_n
  );


  or

  (
    g245_n,
    g243_p,
    g244_p
  );


  and

  (
    g246_p,
    G148_n_spl_00,
    G166_n_spl_001
  );


  and

  (
    g247_p,
    G148_p_spl_00,
    G169_p_spl_001
  );


  or

  (
    g248_n,
    g246_p,
    g247_p
  );


  or

  (
    g249_n,
    g245_n_spl_0,
    g248_n_spl_
  );


  and

  (
    g250_p,
    G101_p_spl_001,
    G119_p_spl_00
  );


  or

  (
    g250_n,
    G101_n_spl_001,
    G119_n_spl_00
  );


  and

  (
    g251_p,
    G100_p_spl_000,
    G119_n_spl_00
  );


  or

  (
    g251_n,
    G100_n_spl_000,
    G119_p_spl_00
  );


  and

  (
    g252_p,
    g250_n,
    g251_n
  );


  or

  (
    g252_n,
    g250_p,
    g251_p
  );


  and

  (
    g253_p,
    G146_p_spl_0,
    g252_n
  );


  or

  (
    g253_n,
    G146_n_spl_0,
    g252_p
  );


  and

  (
    g254_p,
    G102_n_spl_000,
    G119_p_spl_01
  );


  or

  (
    g254_n,
    G102_p_spl_000,
    G119_n_spl_01
  );


  and

  (
    g255_p,
    G98_n_spl_000,
    G119_n_spl_01
  );


  or

  (
    g255_n,
    G98_p_spl_000,
    G119_p_spl_01
  );


  and

  (
    g256_p,
    g254_n,
    g255_n
  );


  or

  (
    g256_n,
    g254_p,
    g255_p
  );


  and

  (
    g257_p,
    G146_n_spl_0,
    g256_n
  );


  or

  (
    g257_n,
    G146_p_spl_0,
    g256_p
  );


  and

  (
    g258_p,
    g253_n,
    g257_n
  );


  or

  (
    g258_n,
    g253_p,
    g257_p
  );


  and

  (
    g259_p,
    G101_p_spl_001,
    G117_p_spl_00
  );


  or

  (
    g259_n,
    G101_n_spl_001,
    G117_n_spl_00
  );


  and

  (
    g260_p,
    G100_p_spl_001,
    G117_n_spl_00
  );


  or

  (
    g260_n,
    G100_n_spl_001,
    G117_p_spl_00
  );


  and

  (
    g261_p,
    g259_n,
    g260_n
  );


  or

  (
    g261_n,
    g259_p,
    g260_p
  );


  and

  (
    g262_p,
    G145_p_spl_0,
    g261_n
  );


  or

  (
    g262_n,
    G145_n_spl_0,
    g261_p
  );


  and

  (
    g263_p,
    G102_n_spl_001,
    G117_p_spl_01
  );


  or

  (
    g263_n,
    G102_p_spl_001,
    G117_n_spl_01
  );


  and

  (
    g264_p,
    G98_n_spl_001,
    G117_n_spl_01
  );


  or

  (
    g264_n,
    G98_p_spl_001,
    G117_p_spl_01
  );


  and

  (
    g265_p,
    g263_n,
    g264_n
  );


  or

  (
    g265_n,
    g263_p,
    g264_p
  );


  and

  (
    g266_p,
    G145_n_spl_0,
    g265_n
  );


  or

  (
    g266_n,
    G145_p_spl_0,
    g265_p
  );


  and

  (
    g267_p,
    g262_n,
    g266_n
  );


  or

  (
    g267_n,
    g262_p,
    g266_p
  );


  and

  (
    g268_p,
    g258_p_spl_,
    g267_p_spl_
  );


  or

  (
    g268_n,
    g258_n_spl_0,
    g267_n_spl_0
  );


  and

  (
    g269_p,
    G121_p_spl_000,
    G168_p_spl_001
  );


  and

  (
    g270_p,
    G121_n_spl_000,
    G169_p_spl_001
  );


  or

  (
    g271_n,
    g269_p,
    g270_p
  );


  and

  (
    g272_p,
    G147_p_spl_00,
    g271_n
  );


  and

  (
    g273_p,
    G121_p_spl_000,
    G167_n_spl_001
  );


  and

  (
    g274_p,
    G121_n_spl_000,
    G166_n_spl_001
  );


  or

  (
    g275_n,
    g273_p,
    g274_p
  );


  and

  (
    g276_p,
    G147_n_spl_00,
    g275_n
  );


  or

  (
    g277_n,
    g272_p,
    g276_p
  );


  or

  (
    g278_n,
    g268_n_spl_,
    g277_n_spl_
  );


  or

  (
    g279_n,
    g249_n,
    g278_n
  );


  or

  (
    g280_n,
    g242_n,
    g279_n
  );


  and

  (
    g281_p,
    G107_p_spl_000,
    G168_p_spl_001
  );


  and

  (
    g282_p,
    G107_n_spl_000,
    G169_p_spl_010
  );


  or

  (
    g283_n,
    g281_p,
    g282_p
  );


  and

  (
    g284_p,
    G139_p_spl_00,
    g283_n
  );


  and

  (
    g285_p,
    G107_p_spl_000,
    G167_n_spl_001
  );


  and

  (
    g286_p,
    G107_n_spl_000,
    G166_n_spl_010
  );


  or

  (
    g287_n,
    g285_p,
    g286_p
  );


  and

  (
    g288_p,
    G139_n_spl_00,
    g287_n
  );


  or

  (
    g289_n,
    g284_p,
    g288_p
  );


  and

  (
    g290_p,
    G105_p_spl_000,
    G168_p_spl_010
  );


  and

  (
    g291_p,
    G105_n_spl_000,
    G169_p_spl_010
  );


  or

  (
    g292_n,
    g290_p,
    g291_p
  );


  and

  (
    g293_p,
    G138_p_spl_00,
    g292_n
  );


  and

  (
    g294_p,
    G105_p_spl_000,
    G167_n_spl_010
  );


  and

  (
    g295_p,
    G105_n_spl_000,
    G166_n_spl_010
  );


  or

  (
    g296_n,
    g294_p,
    g295_p
  );


  and

  (
    g297_p,
    G138_n_spl_00,
    g296_n
  );


  or

  (
    g298_n,
    g293_p,
    g297_p
  );


  or

  (
    g299_n,
    g289_n_spl_,
    g298_n_spl_
  );


  and

  (
    g300_p,
    G109_p_spl_000,
    G168_p_spl_010
  );


  and

  (
    g301_p,
    G109_n_spl_000,
    G169_p_spl_011
  );


  or

  (
    g302_n,
    g300_p,
    g301_p
  );


  and

  (
    g303_p,
    G135_p_spl_00,
    g302_n
  );


  and

  (
    g304_p,
    G109_p_spl_000,
    G167_n_spl_010
  );


  and

  (
    g305_p,
    G109_n_spl_000,
    G166_n_spl_011
  );


  or

  (
    g306_n,
    g304_p,
    g305_p
  );


  and

  (
    g307_p,
    G135_n_spl_00,
    g306_n
  );


  or

  (
    g308_n,
    g303_p,
    g307_p
  );


  and

  (
    g309_p,
    G88_p_spl_00,
    G100_p_spl_001
  );


  or

  (
    g309_n,
    G88_n_spl_00,
    G100_n_spl_001
  );


  and

  (
    g310_p,
    G88_n_spl_00,
    G101_p_spl_010
  );


  or

  (
    g310_n,
    G88_p_spl_00,
    G101_n_spl_010
  );


  and

  (
    g311_p,
    g309_n,
    g310_n
  );


  or

  (
    g311_n,
    g309_p,
    g310_p
  );


  and

  (
    g312_p,
    G142_p_spl_0,
    g311_n
  );


  or

  (
    g312_n,
    G142_n_spl_0,
    g311_p
  );


  and

  (
    g313_p,
    G88_n_spl_01,
    G102_n_spl_001
  );


  or

  (
    g313_n,
    G88_p_spl_01,
    G102_p_spl_001
  );


  and

  (
    g314_p,
    G88_p_spl_01,
    G98_n_spl_001
  );


  or

  (
    g314_n,
    G88_n_spl_01,
    G98_p_spl_001
  );


  and

  (
    g315_p,
    g313_n,
    g314_n
  );


  or

  (
    g315_n,
    g313_p,
    g314_p
  );


  and

  (
    g316_p,
    G142_n_spl_0,
    g315_n
  );


  or

  (
    g316_n,
    G142_p_spl_0,
    g315_p
  );


  and

  (
    g317_p,
    g312_n,
    g316_n
  );


  or

  (
    g317_n,
    g312_p,
    g316_p
  );


  or

  (
    g318_n,
    g308_n_spl_,
    g317_n_spl_0
  );


  or

  (
    g319_n,
    g299_n,
    g318_n
  );


  and

  (
    g320_p,
    G90_p_spl_000,
    G168_p_spl_01
  );


  and

  (
    g321_p,
    G90_n_spl_000,
    G169_p_spl_011
  );


  or

  (
    g322_n,
    g320_p,
    g321_p
  );


  and

  (
    g323_p,
    G143_p_spl_00,
    g322_n
  );


  and

  (
    g324_p,
    G90_p_spl_000,
    G167_n_spl_01
  );


  and

  (
    g325_p,
    G90_n_spl_000,
    G166_n_spl_011
  );


  or

  (
    g326_n,
    g324_p,
    g325_p
  );


  and

  (
    g327_p,
    G143_n_spl_00,
    g326_n
  );


  or

  (
    g328_n,
    g323_p,
    g327_p
  );


  and

  (
    g329_p,
    G92_p_spl_000,
    G168_p_spl_10
  );


  and

  (
    g330_p,
    G92_n_spl_000,
    G169_p_spl_10
  );


  or

  (
    g331_n,
    g329_p,
    g330_p
  );


  and

  (
    g332_p,
    G144_p_spl_00,
    g331_n
  );


  and

  (
    g333_p,
    G92_p_spl_000,
    G167_n_spl_10
  );


  and

  (
    g334_p,
    G92_n_spl_000,
    G166_n_spl_10
  );


  or

  (
    g335_n,
    g333_p,
    g334_p
  );


  and

  (
    g336_p,
    G144_n_spl_00,
    g335_n
  );


  or

  (
    g337_n,
    g332_p,
    g336_p
  );


  or

  (
    g338_n,
    g328_n_spl_,
    g337_n_spl_
  );


  and

  (
    g339_p,
    G94_p_spl_000,
    G168_p_spl_10
  );


  and

  (
    g340_p,
    G94_n_spl_000,
    G169_p_spl_10
  );


  or

  (
    g341_n,
    g339_p,
    g340_p
  );


  and

  (
    g342_p,
    G140_p_spl_00,
    g341_n
  );


  and

  (
    g343_p,
    G94_p_spl_000,
    G167_n_spl_10
  );


  and

  (
    g344_p,
    G94_n_spl_000,
    G166_n_spl_10
  );


  or

  (
    g345_n,
    g343_p,
    g344_p
  );


  and

  (
    g346_p,
    G140_n_spl_00,
    g345_n
  );


  or

  (
    g347_n,
    g342_p,
    g346_p
  );


  and

  (
    g348_p,
    G96_p_spl_000,
    G168_p_spl_11
  );


  and

  (
    g349_p,
    G96_n_spl_000,
    G169_p_spl_11
  );


  or

  (
    g350_n,
    g348_p,
    g349_p
  );


  and

  (
    g351_p,
    G141_p_spl_00,
    g350_n
  );


  and

  (
    g352_p,
    G96_p_spl_000,
    G167_n_spl_11
  );


  and

  (
    g353_p,
    G96_n_spl_000,
    G166_n_spl_11
  );


  or

  (
    g354_n,
    g352_p,
    g353_p
  );


  and

  (
    g355_p,
    G141_n_spl_00,
    g354_n
  );


  or

  (
    g356_n,
    g351_p,
    g355_p
  );


  and

  (
    g357_p,
    G103_p_spl_000,
    G168_p_spl_11
  );


  and

  (
    g358_p,
    G103_n_spl_000,
    G169_p_spl_11
  );


  or

  (
    g359_n,
    g357_p,
    g358_p
  );


  and

  (
    g360_p,
    G137_p_spl_00,
    g359_n
  );


  and

  (
    g361_p,
    G103_p_spl_000,
    G167_n_spl_11
  );


  and

  (
    g362_p,
    G103_n_spl_000,
    G166_n_spl_11
  );


  or

  (
    g363_n,
    g361_p,
    g362_p
  );


  and

  (
    g364_p,
    G137_n_spl_00,
    g363_n
  );


  or

  (
    g365_n,
    g360_p,
    g364_p
  );


  or

  (
    g366_n,
    g356_n_spl_,
    g365_n_spl_
  );


  or

  (
    g367_n,
    g347_n_spl_,
    g366_n
  );


  or

  (
    g368_n,
    g338_n,
    g367_n
  );


  or

  (
    g369_n,
    g319_n,
    g368_n
  );


  and

  (
    g370_p,
    G95_n,
    G124_n_spl_0000
  );


  or

  (
    g370_n,
    G95_p,
    G124_p_spl_0000
  );


  and

  (
    g371_p,
    G94_n_spl_00,
    G124_p_spl_0000
  );


  or

  (
    g371_n,
    G94_p_spl_00,
    G124_n_spl_0000
  );


  and

  (
    g372_p,
    g370_n,
    g371_n
  );


  or

  (
    g372_n,
    g370_p,
    g371_p
  );


  and

  (
    g373_p,
    G140_p_spl_00,
    g372_p_spl_0
  );


  or

  (
    g373_n,
    G140_n_spl_00,
    g372_n_spl_0
  );


  and

  (
    g374_p,
    G140_n_spl_0,
    g372_n_spl_0
  );


  or

  (
    g374_n,
    G140_p_spl_0,
    g372_p_spl_0
  );


  and

  (
    g375_p,
    g373_n_spl_0,
    g374_n_spl_0
  );


  or

  (
    g375_n,
    g373_p_spl_0,
    g374_p_spl_0
  );


  and

  (
    g376_p,
    G93_n,
    G124_n_spl_0001
  );


  or

  (
    g376_n,
    G93_p,
    G124_p_spl_0001
  );


  and

  (
    g377_p,
    G92_n_spl_00,
    G124_p_spl_0001
  );


  or

  (
    g377_n,
    G92_p_spl_00,
    G124_n_spl_0001
  );


  and

  (
    g378_p,
    g376_n,
    g377_n
  );


  or

  (
    g378_n,
    g376_p,
    g377_p
  );


  and

  (
    g379_p,
    G144_p_spl_00,
    g378_p_spl_0
  );


  or

  (
    g379_n,
    G144_n_spl_00,
    g378_n_spl_0
  );


  and

  (
    g380_p,
    G144_n_spl_0,
    g378_n_spl_0
  );


  or

  (
    g380_n,
    G144_p_spl_0,
    g378_p_spl_0
  );


  and

  (
    g381_p,
    g379_n_spl_,
    g380_n_spl_
  );


  or

  (
    g381_n,
    g379_p_spl_,
    g380_p_spl_
  );


  and

  (
    g382_p,
    g375_p_spl_00,
    g381_p_spl_00
  );


  or

  (
    g382_n,
    g375_n_spl_00,
    g381_n_spl_00
  );


  and

  (
    g383_p,
    G91_n,
    G124_n_spl_0010
  );


  or

  (
    g383_n,
    G91_p,
    G124_p_spl_0010
  );


  and

  (
    g384_p,
    G90_n_spl_00,
    G124_p_spl_0010
  );


  or

  (
    g384_n,
    G90_p_spl_00,
    G124_n_spl_0010
  );


  and

  (
    g385_p,
    g383_n,
    g384_n
  );


  or

  (
    g385_n,
    g383_p,
    g384_p
  );


  and

  (
    g386_p,
    G143_p_spl_00,
    g385_p_spl_0
  );


  or

  (
    g386_n,
    G143_n_spl_00,
    g385_n_spl_0
  );


  and

  (
    g387_p,
    G143_n_spl_0,
    g385_n_spl_0
  );


  or

  (
    g387_n,
    G143_p_spl_0,
    g385_p_spl_0
  );


  and

  (
    g388_p,
    g386_n_spl_,
    g387_n_spl_
  );


  or

  (
    g388_n,
    g386_p_spl_,
    g387_p_spl_
  );


  and

  (
    g389_p,
    g382_p_spl_,
    g388_p_spl_00
  );


  or

  (
    g389_n,
    g382_n_spl_,
    g388_n_spl_00
  );


  and

  (
    g390_p,
    G89_n,
    G124_n_spl_0011
  );


  or

  (
    g390_n,
    G89_p,
    G124_p_spl_0011
  );


  and

  (
    g391_p,
    G88_n_spl_10,
    G124_p_spl_0011
  );


  or

  (
    g391_n,
    G88_p_spl_10,
    G124_n_spl_0011
  );


  and

  (
    g392_p,
    g390_n,
    g391_n
  );


  or

  (
    g392_n,
    g390_p,
    g391_p
  );


  and

  (
    g393_p,
    G142_p_spl_1,
    g392_p_spl_0
  );


  or

  (
    g393_n,
    G142_n_spl_1,
    g392_n_spl_0
  );


  and

  (
    g394_p,
    G142_n_spl_1,
    g392_n_spl_0
  );


  or

  (
    g394_n,
    G142_p_spl_1,
    g392_p_spl_0
  );


  and

  (
    g395_p,
    g393_n_spl_,
    g394_n
  );


  or

  (
    g395_n,
    g393_p,
    g394_p
  );


  or

  (
    g396_n,
    g389_n_spl_0,
    g395_n_spl_00
  );


  and

  (
    g397_p,
    G110_n,
    G124_n_spl_010
  );


  or

  (
    g397_n,
    G110_p,
    G124_p_spl_010
  );


  and

  (
    g398_p,
    G109_n_spl_00,
    G124_p_spl_010
  );


  or

  (
    g398_n,
    G109_p_spl_00,
    G124_n_spl_010
  );


  and

  (
    g399_p,
    g397_n,
    g398_n
  );


  or

  (
    g399_n,
    g397_p,
    g398_p
  );


  and

  (
    g400_p,
    G135_p_spl_00,
    g399_p_spl_0
  );


  or

  (
    g400_n,
    G135_n_spl_00,
    g399_n_spl_0
  );


  and

  (
    g401_p,
    G135_n_spl_0,
    g399_n_spl_0
  );


  or

  (
    g401_n,
    G135_p_spl_0,
    g399_p_spl_0
  );


  and

  (
    g402_p,
    g400_n_spl_00,
    g401_n_spl_0
  );


  or

  (
    g402_n,
    g400_p_spl_00,
    g401_p_spl_0
  );


  and

  (
    g403_p,
    G108_n,
    G124_n_spl_011
  );


  or

  (
    g403_n,
    G108_p,
    G124_p_spl_011
  );


  and

  (
    g404_p,
    G107_n_spl_00,
    G124_p_spl_011
  );


  or

  (
    g404_n,
    G107_p_spl_00,
    G124_n_spl_011
  );


  and

  (
    g405_p,
    g403_n,
    g404_n
  );


  or

  (
    g405_n,
    g403_p,
    g404_p
  );


  and

  (
    g406_p,
    G139_p_spl_00,
    g405_p_spl_0
  );


  or

  (
    g406_n,
    G139_n_spl_00,
    g405_n_spl_0
  );


  and

  (
    g407_p,
    G139_n_spl_0,
    g405_n_spl_0
  );


  or

  (
    g407_n,
    G139_p_spl_0,
    g405_p_spl_0
  );


  and

  (
    g408_p,
    g406_n_spl_0,
    g407_n
  );


  or

  (
    g408_n,
    g406_p_spl_0,
    g407_p
  );


  and

  (
    g409_p,
    g402_p_spl_0,
    g408_p_spl_0
  );


  or

  (
    g409_n,
    g402_n_spl_0,
    g408_n_spl_00
  );


  and

  (
    g410_p,
    G106_n,
    G124_n_spl_100
  );


  or

  (
    g410_n,
    G106_p,
    G124_p_spl_100
  );


  and

  (
    g411_p,
    G105_n_spl_00,
    G124_p_spl_100
  );


  or

  (
    g411_n,
    G105_p_spl_00,
    G124_n_spl_100
  );


  and

  (
    g412_p,
    g410_n,
    g411_n
  );


  or

  (
    g412_n,
    g410_p,
    g411_p
  );


  and

  (
    g413_p,
    G138_p_spl_00,
    g412_p_spl_0
  );


  or

  (
    g413_n,
    G138_n_spl_00,
    g412_n_spl_0
  );


  and

  (
    g414_p,
    G138_n_spl_0,
    g412_n_spl_0
  );


  or

  (
    g414_n,
    G138_p_spl_0,
    g412_p_spl_0
  );


  and

  (
    g415_p,
    g413_n_spl_,
    g414_n
  );


  or

  (
    g415_n,
    g413_p_spl_,
    g414_p
  );


  and

  (
    g416_p,
    g409_p_spl_0,
    g415_p_spl_00
  );


  or

  (
    g416_n,
    g409_n_spl_0,
    g415_n_spl_00
  );


  and

  (
    g417_p,
    G104_n,
    G124_n_spl_101
  );


  or

  (
    g417_n,
    G104_p,
    G124_p_spl_101
  );


  and

  (
    g418_p,
    G103_n_spl_00,
    G124_p_spl_101
  );


  or

  (
    g418_n,
    G103_p_spl_00,
    G124_n_spl_101
  );


  and

  (
    g419_p,
    g417_n,
    g418_n
  );


  or

  (
    g419_n,
    g417_p,
    g418_p
  );


  and

  (
    g420_p,
    G137_p_spl_00,
    g419_p_spl_0
  );


  or

  (
    g420_n,
    G137_n_spl_00,
    g419_n_spl_0
  );


  and

  (
    g421_p,
    G137_n_spl_0,
    g419_n_spl_0
  );


  or

  (
    g421_n,
    G137_p_spl_0,
    g419_p_spl_0
  );


  and

  (
    g422_p,
    g420_n_spl_0,
    g421_n
  );


  or

  (
    g422_n,
    g420_p_spl_0,
    g421_p
  );


  and

  (
    g423_p,
    g416_p_spl_0,
    g422_p_spl_00
  );


  or

  (
    g423_n,
    g416_n_spl_0,
    g422_n_spl_00
  );


  and

  (
    g424_p,
    G97_n,
    G124_n_spl_110
  );


  or

  (
    g424_n,
    G97_p,
    G124_p_spl_110
  );


  and

  (
    g425_p,
    G96_n_spl_00,
    G124_p_spl_110
  );


  or

  (
    g425_n,
    G96_p_spl_00,
    G124_n_spl_110
  );


  and

  (
    g426_p,
    g424_n,
    g425_n
  );


  or

  (
    g426_n,
    g424_p,
    g425_p
  );


  and

  (
    g427_p,
    G141_p_spl_00,
    g426_p_spl_0
  );


  or

  (
    g427_n,
    G141_n_spl_00,
    g426_n_spl_0
  );


  and

  (
    g428_p,
    G141_n_spl_0,
    g426_n_spl_0
  );


  or

  (
    g428_n,
    G141_p_spl_0,
    g426_p_spl_0
  );


  and

  (
    g429_p,
    g427_n_spl_,
    g428_n
  );


  or

  (
    g429_n,
    g427_p_spl_,
    g428_p
  );


  and

  (
    g430_p,
    g423_p_spl_,
    g429_p_spl_00
  );


  or

  (
    g430_n,
    g423_n_spl_,
    g429_n_spl_00
  );


  or

  (
    g431_n,
    g396_n_spl_,
    g430_n_spl_0
  );


  and

  (
    g432_p,
    G118_n,
    G123_n_spl_0000
  );


  or

  (
    g432_n,
    G118_p,
    G123_p_spl_0000
  );


  and

  (
    g433_p,
    G117_n_spl_10,
    G123_p_spl_0000
  );


  or

  (
    g433_n,
    G117_p_spl_10,
    G123_n_spl_0000
  );


  and

  (
    g434_p,
    g432_n,
    g433_n
  );


  or

  (
    g434_n,
    g432_p,
    g433_p
  );


  and

  (
    g435_p,
    G145_p_spl_1,
    g434_p_spl_0
  );


  or

  (
    g435_n,
    G145_n_spl_1,
    g434_n_spl_0
  );


  and

  (
    g436_p,
    G145_n_spl_1,
    g434_n_spl_0
  );


  or

  (
    g436_n,
    G145_p_spl_1,
    g434_p_spl_0
  );


  and

  (
    g437_p,
    g435_n_spl_,
    g436_n
  );


  or

  (
    g437_n,
    g435_p_spl_,
    g436_p
  );


  and

  (
    g438_p,
    G120_n,
    G123_n_spl_0001
  );


  or

  (
    g438_n,
    G120_p,
    G123_p_spl_0001
  );


  and

  (
    g439_p,
    G119_n_spl_10,
    G123_p_spl_0001
  );


  or

  (
    g439_n,
    G119_p_spl_10,
    G123_n_spl_0001
  );


  and

  (
    g440_p,
    g438_n,
    g439_n
  );


  or

  (
    g440_n,
    g438_p,
    g439_p
  );


  and

  (
    g441_p,
    G146_p_spl_1,
    g440_p_spl_0
  );


  or

  (
    g441_n,
    G146_n_spl_1,
    g440_n_spl_0
  );


  and

  (
    g442_p,
    G146_n_spl_1,
    g440_n_spl_0
  );


  or

  (
    g442_n,
    G146_p_spl_1,
    g440_p_spl_0
  );


  and

  (
    g443_p,
    g441_n_spl_00,
    g442_n_spl_0
  );


  or

  (
    g443_n,
    g441_p_spl_00,
    g442_p_spl_0
  );


  and

  (
    g444_p,
    g437_p_spl_00,
    g443_p_spl_00
  );


  or

  (
    g444_n,
    g437_n_spl_00,
    g443_n_spl_00
  );


  and

  (
    g445_p,
    G122_n,
    G123_n_spl_0010
  );


  or

  (
    g445_n,
    G122_p,
    G123_p_spl_0010
  );


  and

  (
    g446_p,
    G121_n_spl_00,
    G123_p_spl_0010
  );


  or

  (
    g446_n,
    G121_p_spl_00,
    G123_n_spl_0010
  );


  and

  (
    g447_p,
    g445_n,
    g446_n
  );


  or

  (
    g447_n,
    g445_p,
    g446_p
  );


  and

  (
    g448_p,
    G147_p_spl_00,
    g447_p_spl_0
  );


  or

  (
    g448_n,
    G147_n_spl_00,
    g447_n_spl_0
  );


  and

  (
    g449_p,
    G147_n_spl_0,
    g447_n_spl_0
  );


  or

  (
    g449_n,
    G147_p_spl_0,
    g447_p_spl_0
  );


  and

  (
    g450_p,
    g448_n_spl_,
    g449_n
  );


  or

  (
    g450_n,
    g448_p_spl_,
    g449_p
  );


  and

  (
    g451_p,
    G123_n_spl_001,
    G125_n_spl_
  );


  or

  (
    g451_n,
    G123_p_spl_001,
    G125_p
  );


  and

  (
    g452_p,
    G148_p_spl_00,
    g451_n_spl_0
  );


  or

  (
    g452_n,
    G148_n_spl_00,
    g451_p_spl_0
  );


  and

  (
    g453_p,
    G148_n_spl_0,
    g451_p_spl_0
  );


  or

  (
    g453_n,
    G148_p_spl_0,
    g451_n_spl_0
  );


  and

  (
    g454_p,
    g452_n_spl_0,
    g453_n
  );


  or

  (
    g454_n,
    g452_p_spl_0,
    g453_p
  );


  and

  (
    g455_p,
    g450_p_spl_0,
    g454_p_spl_0
  );


  or

  (
    g455_n,
    g450_n_spl_0,
    g454_n_spl_00
  );


  and

  (
    g456_p,
    G123_n_spl_010,
    G129_n_spl_
  );


  or

  (
    g456_n,
    G123_p_spl_010,
    G129_p
  );


  and

  (
    g457_p,
    G123_p_spl_010,
    G128_n_spl_00
  );


  or

  (
    g457_n,
    G123_n_spl_010,
    G128_p_spl_00
  );


  and

  (
    g458_p,
    g456_n,
    g457_n
  );


  or

  (
    g458_n,
    g456_p,
    g457_p
  );


  and

  (
    g459_p,
    G150_p_spl_00,
    g458_p_spl_0
  );


  or

  (
    g459_n,
    G150_n_spl_00,
    g458_n_spl_0
  );


  and

  (
    g460_p,
    G150_n_spl_0,
    g458_n_spl_0
  );


  or

  (
    g460_n,
    G150_p_spl_0,
    g458_p_spl_0
  );


  and

  (
    g461_p,
    g459_n_spl_0,
    g460_n
  );


  or

  (
    g461_n,
    g459_p_spl_0,
    g460_p
  );


  and

  (
    g462_p,
    G123_n_spl_011,
    G131_n_spl_
  );


  or

  (
    g462_n,
    G123_p_spl_011,
    G131_p
  );


  and

  (
    g463_p,
    G123_p_spl_011,
    G130_n_spl_0
  );


  or

  (
    g463_n,
    G123_n_spl_011,
    G130_p_spl_0
  );


  and

  (
    g464_p,
    g462_n,
    g463_n
  );


  or

  (
    g464_n,
    g462_p,
    g463_p
  );


  and

  (
    g465_p,
    g461_p_spl_0,
    g464_n_spl_00
  );


  or

  (
    g465_n,
    g461_n_spl_0,
    g464_p_spl_00
  );


  and

  (
    g466_p,
    G123_n_spl_100,
    G127_n_spl_
  );


  or

  (
    g466_n,
    G123_p_spl_100,
    G127_p
  );


  and

  (
    g467_p,
    G123_p_spl_100,
    G126_n_spl_00
  );


  or

  (
    g467_n,
    G123_n_spl_100,
    G126_p_spl_00
  );


  and

  (
    g468_p,
    g466_n,
    g467_n
  );


  or

  (
    g468_n,
    g466_p,
    g467_p
  );


  and

  (
    g469_p,
    G149_p_spl_00,
    g468_p_spl_0
  );


  or

  (
    g469_n,
    G149_n_spl_00,
    g468_n_spl_0
  );


  and

  (
    g470_p,
    G149_n_spl_0,
    g468_n_spl_0
  );


  or

  (
    g470_n,
    G149_p_spl_0,
    g468_p_spl_0
  );


  and

  (
    g471_p,
    g469_n_spl_0,
    g470_n
  );


  or

  (
    g471_n,
    g469_p_spl_0,
    g470_p
  );


  and

  (
    g472_p,
    g465_p_spl_0,
    g471_p_spl_0
  );


  or

  (
    g472_n,
    g465_n_spl_0,
    g471_n_spl_00
  );


  and

  (
    g473_p,
    g455_p_spl_,
    g472_p_spl_
  );


  or

  (
    g473_n,
    g455_n_spl_,
    g472_n_spl_
  );


  and

  (
    g474_p,
    G114_n_spl_0,
    G123_n_spl_101
  );


  or

  (
    g474_n,
    G114_p_spl_,
    G123_p_spl_101
  );


  and

  (
    g475_p,
    G113_n_spl_01,
    G123_p_spl_101
  );


  or

  (
    g475_n,
    G113_p_spl_0,
    G123_n_spl_101
  );


  and

  (
    g476_p,
    g474_n,
    g475_n
  );


  or

  (
    g476_n,
    g474_p,
    g475_p
  );


  and

  (
    g477_p,
    G116_n,
    G123_n_spl_110
  );


  or

  (
    g477_n,
    G116_p,
    G123_p_spl_110
  );


  and

  (
    g478_p,
    G115_n_spl_0,
    G123_p_spl_110
  );


  or

  (
    g478_n,
    G115_p_spl_0,
    G123_n_spl_110
  );


  and

  (
    g479_p,
    g477_n,
    g478_n
  );


  or

  (
    g479_n,
    g477_p,
    g478_p
  );


  and

  (
    g480_p,
    g476_n_spl_0,
    g479_n_spl_00
  );


  or

  (
    g480_n,
    g476_p_spl_00,
    g479_p_spl_00
  );


  and

  (
    g481_p,
    g473_p_spl_,
    g480_p_spl_0
  );


  and

  (
    g482_p,
    g444_p_spl_0,
    g481_p
  );


  and

  (
    g483_p,
    G117_n_spl_10,
    G119_n_spl_10
  );


  or

  (
    g483_n,
    G117_p_spl_10,
    G119_p_spl_10
  );


  and

  (
    g484_p,
    G117_p_spl_1,
    G119_p_spl_1
  );


  or

  (
    g484_n,
    G117_n_spl_1,
    G119_n_spl_1
  );


  and

  (
    g485_p,
    g483_n,
    g484_n
  );


  or

  (
    g485_n,
    g483_p,
    g484_p
  );


  and

  (
    g486_p,
    G113_n_spl_01,
    G115_n_spl_1
  );


  or

  (
    g486_n,
    G113_p_spl_1,
    G115_p_spl_1
  );


  and

  (
    g487_p,
    G113_p_spl_1,
    G115_p_spl_1
  );


  or

  (
    g487_n,
    G113_n_spl_1,
    G115_n_spl_1
  );


  and

  (
    g488_p,
    g486_n,
    g487_n
  );


  or

  (
    g488_n,
    g486_p,
    g487_p
  );


  and

  (
    g489_p,
    g485_p_spl_,
    g488_n_spl_
  );


  or

  (
    g489_n,
    g485_n_spl_,
    g488_p_spl_
  );


  and

  (
    g490_p,
    g485_n_spl_,
    g488_p_spl_
  );


  or

  (
    g490_n,
    g485_p_spl_,
    g488_n_spl_
  );


  and

  (
    g491_p,
    g489_n,
    g490_n
  );


  or

  (
    g491_n,
    g489_p,
    g490_p
  );


  and

  (
    g492_p,
    G130_n_spl_1,
    G132_n_spl_0
  );


  or

  (
    g492_n,
    G130_p_spl_1,
    G132_p_spl_0
  );


  and

  (
    g493_p,
    G130_p_spl_1,
    G132_p_spl_0
  );


  or

  (
    g493_n,
    G130_n_spl_1,
    G132_n_spl_0
  );


  and

  (
    g494_p,
    g492_n,
    g493_n
  );


  or

  (
    g494_n,
    g492_p,
    g493_p
  );


  and

  (
    g495_p,
    G121_p_spl_01,
    g494_n_spl_
  );


  or

  (
    g495_n,
    G121_n_spl_01,
    g494_p_spl_
  );


  and

  (
    g496_p,
    G121_n_spl_01,
    g494_p_spl_
  );


  or

  (
    g496_n,
    G121_p_spl_01,
    g494_n_spl_
  );


  and

  (
    g497_p,
    g495_n,
    g496_n
  );


  or

  (
    g497_n,
    g495_p,
    g496_p
  );


  and

  (
    g498_p,
    G126_n_spl_01,
    G128_n_spl_01
  );


  or

  (
    g498_n,
    G126_p_spl_01,
    G128_p_spl_01
  );


  and

  (
    g499_p,
    G126_p_spl_01,
    G128_p_spl_01
  );


  or

  (
    g499_n,
    G126_n_spl_01,
    G128_n_spl_01
  );


  and

  (
    g500_p,
    g498_n,
    g499_n
  );


  or

  (
    g500_n,
    g498_p,
    g499_p
  );


  and

  (
    g501_p,
    g497_n_spl_,
    g500_n_spl_
  );


  or

  (
    g501_n,
    g497_p_spl_,
    g500_p_spl_
  );


  and

  (
    g502_p,
    g497_p_spl_,
    g500_p_spl_
  );


  or

  (
    g502_n,
    g497_n_spl_,
    g500_n_spl_
  );


  and

  (
    g503_p,
    g501_n,
    g502_n
  );


  or

  (
    g503_n,
    g501_p,
    g502_p
  );


  and

  (
    g504_p,
    g491_n,
    g503_p
  );


  and

  (
    g505_p,
    g491_p,
    g503_n
  );


  or

  (
    g506_n,
    g504_p,
    g505_p
  );


  and

  (
    g507_p,
    G92_n_spl_01,
    G94_n_spl_01
  );


  or

  (
    g507_n,
    G92_p_spl_01,
    G94_p_spl_01
  );


  and

  (
    g508_p,
    G92_p_spl_01,
    G94_p_spl_01
  );


  or

  (
    g508_n,
    G92_n_spl_01,
    G94_n_spl_01
  );


  and

  (
    g509_p,
    g507_n,
    g508_n
  );


  or

  (
    g509_n,
    g507_p,
    g508_p
  );


  and

  (
    g510_p,
    G88_p_spl_10,
    G90_n_spl_01
  );


  or

  (
    g510_n,
    G88_n_spl_10,
    G90_p_spl_01
  );


  and

  (
    g511_p,
    G88_n_spl_1,
    G90_p_spl_01
  );


  or

  (
    g511_n,
    G88_p_spl_1,
    G90_n_spl_01
  );


  and

  (
    g512_p,
    g510_n,
    g511_n
  );


  or

  (
    g512_n,
    g510_p,
    g511_p
  );


  and

  (
    g513_p,
    g509_p_spl_,
    g512_n_spl_
  );


  or

  (
    g513_n,
    g509_n_spl_,
    g512_p_spl_
  );


  and

  (
    g514_p,
    g509_n_spl_,
    g512_p_spl_
  );


  or

  (
    g514_n,
    g509_p_spl_,
    g512_n_spl_
  );


  and

  (
    g515_p,
    g513_n,
    g514_n
  );


  or

  (
    g515_n,
    g513_p,
    g514_p
  );


  and

  (
    g516_p,
    G96_n_spl_01,
    G103_n_spl_01
  );


  or

  (
    g516_n,
    G96_p_spl_01,
    G103_p_spl_01
  );


  and

  (
    g517_p,
    G96_p_spl_01,
    G103_p_spl_01
  );


  or

  (
    g517_n,
    G96_n_spl_01,
    G103_n_spl_01
  );


  and

  (
    g518_p,
    g516_n,
    g517_n
  );


  or

  (
    g518_n,
    g516_p,
    g517_p
  );


  and

  (
    g519_p,
    G109_n_spl_01,
    G111_n_spl_0
  );


  or

  (
    g519_n,
    G109_p_spl_01,
    G111_p_spl_0
  );


  and

  (
    g520_p,
    G109_p_spl_01,
    G111_p_spl_0
  );


  or

  (
    g520_n,
    G109_n_spl_01,
    G111_n_spl_0
  );


  and

  (
    g521_p,
    g519_n,
    g520_n
  );


  or

  (
    g521_n,
    g519_p,
    g520_p
  );


  and

  (
    g522_p,
    g518_n_spl_,
    g521_n_spl_
  );


  or

  (
    g522_n,
    g518_p_spl_,
    g521_p_spl_
  );


  and

  (
    g523_p,
    g518_p_spl_,
    g521_p_spl_
  );


  or

  (
    g523_n,
    g518_n_spl_,
    g521_n_spl_
  );


  and

  (
    g524_p,
    g522_n,
    g523_n
  );


  or

  (
    g524_n,
    g522_p,
    g523_p
  );


  and

  (
    g525_p,
    G105_n_spl_01,
    G107_n_spl_01
  );


  or

  (
    g525_n,
    G105_p_spl_01,
    G107_p_spl_01
  );


  and

  (
    g526_p,
    G105_p_spl_01,
    G107_p_spl_01
  );


  or

  (
    g526_n,
    G105_n_spl_01,
    G107_n_spl_01
  );


  and

  (
    g527_p,
    g525_n,
    g526_n
  );


  or

  (
    g527_n,
    g525_p,
    g526_p
  );


  and

  (
    g528_p,
    g524_n_spl_,
    g527_n_spl_
  );


  or

  (
    g528_n,
    g524_p_spl_,
    g527_p_spl_
  );


  and

  (
    g529_p,
    g524_p_spl_,
    g527_p_spl_
  );


  or

  (
    g529_n,
    g524_n_spl_,
    g527_n_spl_
  );


  and

  (
    g530_p,
    g528_n,
    g529_n
  );


  or

  (
    g530_n,
    g528_p,
    g529_p
  );


  and

  (
    g531_p,
    g515_n,
    g530_p
  );


  and

  (
    g532_p,
    g515_p,
    g530_n
  );


  or

  (
    g533_n,
    g531_p,
    g532_p
  );


  and

  (
    g534_p,
    g400_p_spl_00,
    g408_p_spl_0
  );


  or

  (
    g534_n,
    g400_n_spl_00,
    g408_n_spl_00
  );


  and

  (
    g535_p,
    g406_n_spl_0,
    g534_n
  );


  or

  (
    g535_n,
    g406_p_spl_0,
    g534_p
  );


  and

  (
    g536_p,
    g415_p_spl_00,
    g535_n_spl_0
  );


  or

  (
    g536_n,
    g415_n_spl_00,
    g535_p_spl_0
  );


  and

  (
    g537_p,
    g413_n_spl_,
    g536_n
  );


  or

  (
    g537_n,
    g413_p_spl_,
    g536_p
  );


  and

  (
    g538_p,
    g422_p_spl_00,
    g537_n_spl_00
  );


  or

  (
    g538_n,
    g422_n_spl_00,
    g537_p_spl_00
  );


  and

  (
    g539_p,
    g420_n_spl_0,
    g538_n
  );


  or

  (
    g539_n,
    g420_p_spl_0,
    g538_p
  );


  and

  (
    g540_p,
    g429_p_spl_00,
    g539_n_spl_0
  );


  or

  (
    g540_n,
    g429_n_spl_00,
    g539_p_spl_0
  );


  and

  (
    g541_p,
    g427_n_spl_,
    g540_n
  );


  or

  (
    g541_n,
    g427_p_spl_,
    g540_p
  );


  or

  (
    g542_n,
    g396_n_spl_,
    g541_p_spl_00
  );


  and

  (
    g543_p,
    g373_p_spl_0,
    g381_p_spl_00
  );


  or

  (
    g543_n,
    g373_n_spl_0,
    g381_n_spl_00
  );


  and

  (
    g544_p,
    g379_n_spl_,
    g543_n
  );


  or

  (
    g544_n,
    g379_p_spl_,
    g543_p
  );


  and

  (
    g545_p,
    g387_n_spl_,
    g544_n_spl_0
  );


  or

  (
    g545_n,
    g387_p_spl_,
    g544_p_spl_0
  );


  and

  (
    g546_p,
    g386_n_spl_,
    g545_n_spl_
  );


  or

  (
    g546_n,
    g386_p_spl_,
    g545_p_spl_
  );


  or

  (
    g547_n,
    g395_n_spl_00,
    g546_p_spl_0
  );


  and

  (
    g548_p,
    g542_n,
    g547_n
  );


  and

  (
    g549_p,
    g393_n_spl_,
    g548_p
  );


  or

  (
    g550_n,
    g476_p_spl_00,
    g480_p_spl_0
  );


  or

  (
    g551_n,
    G21_n,
    g464_p_spl_00
  );


  or

  (
    g552_n,
    G21_p,
    g464_n_spl_00
  );


  and

  (
    g553_p,
    g551_n,
    g552_n
  );


  and

  (
    g554_p,
    G177_p_spl_0000,
    g553_p_spl_
  );


  or

  (
    g555_n,
    G176_p_spl_00000,
    g554_p
  );


  or

  (
    g556_n,
    G177_n_spl_0000,
    g245_n_spl_0
  );


  or

  (
    g557_n,
    G176_n_spl_0000,
    g556_n
  );


  or

  (
    g558_n,
    G60_p,
    G177_p_spl_0000
  );


  and

  (
    g559_p,
    g557_n,
    g558_n
  );


  and

  (
    g560_p,
    g555_n,
    g559_p
  );


  and

  (
    g561_p,
    g461_n_spl_0,
    g464_p_spl_01
  );


  or

  (
    g561_n,
    g461_p_spl_0,
    g464_n_spl_01
  );


  and

  (
    g562_p,
    g465_n_spl_0,
    g561_n
  );


  or

  (
    g562_n,
    g465_p_spl_0,
    g561_p
  );


  and

  (
    g563_p,
    G177_p_spl_0001,
    g562_n_spl_0
  );


  or

  (
    g564_n,
    G176_p_spl_00000,
    g563_p
  );


  or

  (
    g565_n,
    G177_n_spl_0000,
    g224_n_spl_
  );


  or

  (
    g566_n,
    G176_n_spl_0000,
    g565_n
  );


  or

  (
    g567_n,
    G58_p,
    G177_p_spl_0001
  );


  and

  (
    g568_p,
    g566_n,
    g567_n
  );


  and

  (
    g569_p,
    g564_n,
    g568_p
  );


  and

  (
    g570_p,
    G2_p_spl_0,
    g402_p_spl_0
  );


  or

  (
    g570_n,
    G2_n_spl_0,
    g402_n_spl_0
  );


  or

  (
    g571_n,
    G2_p_spl_0,
    g402_p_spl_1
  );


  and

  (
    g572_p,
    g570_n_spl_,
    g571_n
  );


  and

  (
    g573_p,
    G177_p_spl_0010,
    g572_p_spl_
  );


  or

  (
    g574_n,
    G176_p_spl_00001,
    g573_p
  );


  or

  (
    g575_n,
    G177_n_spl_0001,
    g308_n_spl_
  );


  or

  (
    g576_n,
    G176_n_spl_0001,
    g575_n
  );


  or

  (
    g577_n,
    G48_p,
    G177_p_spl_0010
  );


  and

  (
    g578_p,
    g576_n,
    g577_n
  );


  and

  (
    g579_p,
    g574_n,
    g578_p
  );


  and

  (
    g580_p,
    g476_p_spl_0,
    g479_p_spl_00
  );


  or

  (
    g580_n,
    g476_n_spl_0,
    g479_n_spl_00
  );


  and

  (
    g581_p,
    g480_n,
    g580_n
  );


  or

  (
    g581_n,
    g480_p_spl_,
    g580_p
  );


  and

  (
    g582_p,
    G22_p_spl_,
    G173_n_spl_0000
  );


  and

  (
    g583_p,
    G3_p_spl_,
    G173_p_spl_0000
  );


  or

  (
    g584_n,
    g582_p,
    g583_p
  );


  and

  (
    g585_p,
    G172_n_spl_000,
    g584_n
  );


  or

  (
    g586_n,
    G173_p_spl_0000,
    g579_p_spl_00
  );


  or

  (
    g587_n,
    G173_n_spl_0000,
    g560_p_spl_00
  );


  and

  (
    g588_p,
    G172_p_spl_000,
    g587_n
  );


  and

  (
    g589_p,
    g586_n,
    g588_p
  );


  or

  (
    g590_n,
    g585_p,
    g589_p
  );


  and

  (
    g591_p,
    G19_p,
    G177_n_spl_0001
  );


  and

  (
    g592_p,
    G176_p_spl_00001,
    g591_p
  );


  and

  (
    g593_p,
    G176_p_spl_0001,
    g277_n_spl_
  );


  and

  (
    g594_p,
    g459_p_spl_0,
    g471_p_spl_0
  );


  or

  (
    g594_n,
    g459_n_spl_0,
    g471_n_spl_00
  );


  and

  (
    g595_p,
    g472_n_spl_,
    g594_n_spl_
  );


  or

  (
    g595_n,
    g472_p_spl_,
    g594_p_spl_
  );


  and

  (
    g596_p,
    g469_n_spl_0,
    g595_p
  );


  or

  (
    g596_n,
    g469_p_spl_0,
    g595_n_spl_
  );


  and

  (
    g597_p,
    g454_p_spl_0,
    g596_n_spl_0
  );


  or

  (
    g597_n,
    g454_n_spl_00,
    g596_p_spl_0
  );


  and

  (
    g598_p,
    g452_n_spl_0,
    g597_n
  );


  or

  (
    g598_n,
    g452_p_spl_0,
    g597_p_spl_
  );


  or

  (
    g599_n,
    g450_p_spl_0,
    g598_p_spl_0
  );


  or

  (
    g600_n,
    g450_n_spl_0,
    g598_n_spl_0
  );


  and

  (
    g601_p,
    g599_n,
    g600_n
  );


  and

  (
    g602_p,
    G176_n_spl_0001,
    g601_p_spl_
  );


  or

  (
    g603_n,
    g593_p,
    g602_p
  );


  and

  (
    g604_p,
    G177_p_spl_0011,
    g603_n
  );


  or

  (
    g605_n,
    g592_p,
    g604_p
  );


  and

  (
    g606_p,
    G59_p,
    G177_n_spl_0010
  );


  and

  (
    g607_p,
    G176_p_spl_0001,
    g606_p
  );


  and

  (
    g608_p,
    G176_p_spl_0010,
    g248_n_spl_
  );


  and

  (
    g609_p,
    g454_n_spl_0,
    g596_p_spl_0
  );


  or

  (
    g610_n,
    g597_p_spl_,
    g609_p
  );


  and

  (
    g611_p,
    G176_n_spl_0010,
    g610_n_spl_
  );


  or

  (
    g612_n,
    g608_p,
    g611_p
  );


  and

  (
    g613_p,
    G177_p_spl_0011,
    g612_n
  );


  or

  (
    g614_n,
    g607_p,
    g613_p
  );


  and

  (
    g615_p,
    G50_p,
    G177_n_spl_0010
  );


  and

  (
    g616_p,
    G176_p_spl_0010,
    g615_p
  );


  and

  (
    g617_p,
    g459_n_spl_,
    g465_n_spl_
  );


  or

  (
    g617_n,
    g459_p_spl_,
    g465_p_spl_
  );


  and

  (
    g618_p,
    g471_n_spl_0,
    g617_p_spl_0
  );


  or

  (
    g619_n,
    g595_n_spl_,
    g618_p
  );


  or

  (
    g620_n,
    G176_p_spl_0011,
    g619_n_spl_
  );


  or

  (
    g621_n,
    G176_n_spl_0010,
    g233_n_spl_
  );


  and

  (
    g622_p,
    G177_p_spl_0100,
    g621_n
  );


  and

  (
    g623_p,
    g620_n,
    g622_p
  );


  or

  (
    g624_n,
    g616_p,
    g623_p
  );


  and

  (
    g625_p,
    G22_p_spl_,
    G174_n_spl_0000
  );


  and

  (
    g626_p,
    G3_p_spl_,
    G174_p_spl_0000
  );


  or

  (
    g627_n,
    g625_p,
    g626_p
  );


  and

  (
    g628_p,
    G175_n_spl_000,
    g627_n
  );


  or

  (
    g629_n,
    G174_p_spl_0000,
    g579_p_spl_00
  );


  or

  (
    g630_n,
    G174_n_spl_0000,
    g560_p_spl_00
  );


  and

  (
    g631_p,
    G175_p_spl_000,
    g630_n
  );


  and

  (
    g632_p,
    g629_n,
    g631_p
  );


  or

  (
    g633_n,
    g628_p,
    g632_p
  );


  and

  (
    g634_p,
    G53_p,
    G177_n_spl_0011
  );


  and

  (
    g635_p,
    G176_p_spl_0011,
    g634_p
  );


  or

  (
    g636_n,
    G176_n_spl_0011,
    g356_n_spl_
  );


  and

  (
    g637_p,
    G2_p_spl_1,
    g416_p_spl_0
  );


  or

  (
    g637_n,
    G2_n_spl_0,
    g416_n_spl_0
  );


  and

  (
    g638_p,
    g537_p_spl_00,
    g637_n
  );


  or

  (
    g638_n,
    g537_n_spl_00,
    g637_p
  );


  and

  (
    g639_p,
    g422_p_spl_0,
    g638_n
  );


  or

  (
    g639_n,
    g422_n_spl_01,
    g638_p_spl_
  );


  and

  (
    g640_p,
    g420_n_spl_,
    g639_n
  );


  or

  (
    g640_n,
    g420_p_spl_,
    g639_p_spl_
  );


  and

  (
    g641_p,
    g429_n_spl_01,
    g640_p
  );


  and

  (
    g642_p,
    g429_p_spl_01,
    g640_n
  );


  or

  (
    g643_n,
    g641_p,
    g642_p
  );


  or

  (
    g644_n,
    G176_p_spl_0100,
    g643_n_spl_
  );


  and

  (
    g645_p,
    G177_p_spl_0100,
    g644_n
  );


  and

  (
    g646_p,
    g636_n,
    g645_p
  );


  or

  (
    g647_n,
    g635_p,
    g646_p
  );


  and

  (
    g648_p,
    G57_p,
    G177_n_spl_0011
  );


  and

  (
    g649_p,
    G176_p_spl_0100,
    g648_p
  );


  and

  (
    g650_p,
    G176_p_spl_0101,
    g365_n_spl_
  );


  and

  (
    g651_p,
    g422_n_spl_01,
    g638_p_spl_
  );


  or

  (
    g652_n,
    g639_p_spl_,
    g651_p
  );


  and

  (
    g653_p,
    G176_n_spl_0011,
    g652_n_spl_
  );


  or

  (
    g654_n,
    g650_p,
    g653_p
  );


  and

  (
    g655_p,
    G177_p_spl_0101,
    g654_n
  );


  or

  (
    g656_n,
    g649_p,
    g655_p
  );


  and

  (
    g657_p,
    G56_p,
    G177_n_spl_010
  );


  and

  (
    g658_p,
    G176_p_spl_0101,
    g657_p
  );


  and

  (
    g659_p,
    g400_n_spl_0,
    g570_n_spl_
  );


  or

  (
    g659_n,
    g400_p_spl_0,
    g570_p
  );


  and

  (
    g660_p,
    g408_p_spl_1,
    g659_n
  );


  or

  (
    g660_n,
    g408_n_spl_0,
    g659_p_spl_
  );


  and

  (
    g661_p,
    g406_n_spl_,
    g660_n
  );


  or

  (
    g661_n,
    g406_p_spl_,
    g660_p_spl_
  );


  and

  (
    g662_p,
    g415_n_spl_0,
    g661_p
  );


  and

  (
    g663_p,
    g415_p_spl_0,
    g661_n
  );


  or

  (
    g664_n,
    g662_p,
    g663_p
  );


  or

  (
    g665_n,
    G176_p_spl_0110,
    g664_n_spl_
  );


  or

  (
    g666_n,
    G176_n_spl_0100,
    g298_n_spl_
  );


  and

  (
    g667_p,
    G177_p_spl_0101,
    g666_n
  );


  and

  (
    g668_p,
    g665_n,
    g667_p
  );


  or

  (
    g669_n,
    g658_p,
    g668_p
  );


  and

  (
    g670_p,
    G55_p,
    G177_n_spl_010
  );


  and

  (
    g671_p,
    G176_p_spl_0110,
    g670_p
  );


  and

  (
    g672_p,
    g408_n_spl_1,
    g659_p_spl_
  );


  or

  (
    g673_n,
    g660_p_spl_,
    g672_p
  );


  or

  (
    g674_n,
    G176_p_spl_0111,
    g673_n_spl_
  );


  or

  (
    g675_n,
    G176_n_spl_0100,
    g289_n_spl_
  );


  and

  (
    g676_p,
    G177_p_spl_0110,
    g675_n
  );


  and

  (
    g677_p,
    g674_n,
    g676_p
  );


  or

  (
    g678_n,
    g671_p,
    g677_p
  );


  and

  (
    g679_p,
    g434_n_spl_1,
    g440_n_spl_1
  );


  or

  (
    g679_n,
    g434_p_spl_1,
    g440_p_spl_1
  );


  and

  (
    g680_p,
    g434_p_spl_1,
    g440_p_spl_1
  );


  or

  (
    g680_n,
    g434_n_spl_1,
    g440_n_spl_1
  );


  and

  (
    g681_p,
    g679_n,
    g680_n
  );


  or

  (
    g681_n,
    g679_p,
    g680_p
  );


  and

  (
    g682_p,
    g581_n_spl_00,
    g681_p_spl_
  );


  or

  (
    g682_n,
    g581_p_spl_00,
    g681_n_spl_
  );


  and

  (
    g683_p,
    g581_p_spl_00,
    g681_n_spl_
  );


  or

  (
    g683_n,
    g581_n_spl_00,
    g681_p_spl_
  );


  and

  (
    g684_p,
    g682_n,
    g683_n
  );


  or

  (
    g684_n,
    g682_p,
    g683_p
  );


  and

  (
    g685_p,
    G123_n_spl_111,
    G133_n
  );


  or

  (
    g685_n,
    G123_p_spl_111,
    G133_p
  );


  and

  (
    g686_p,
    G123_p_spl_111,
    G132_n_spl_
  );


  or

  (
    g686_n,
    G123_n_spl_111,
    G132_p_spl_
  );


  and

  (
    g687_p,
    g685_n,
    g686_n
  );


  or

  (
    g687_n,
    g685_p,
    g686_p
  );


  and

  (
    g688_p,
    g464_n_spl_01,
    g687_n_spl_
  );


  or

  (
    g688_n,
    g464_p_spl_01,
    g687_p_spl_
  );


  and

  (
    g689_p,
    g464_p_spl_10,
    g687_p_spl_
  );


  or

  (
    g689_n,
    g464_n_spl_10,
    g687_n_spl_
  );


  and

  (
    g690_p,
    g688_n,
    g689_n
  );


  or

  (
    g690_n,
    g688_p,
    g689_p
  );


  and

  (
    g691_p,
    g447_n_spl_1,
    g451_p_spl_1
  );


  or

  (
    g691_n,
    g447_p_spl_1,
    g451_n_spl_1
  );


  and

  (
    g692_p,
    g447_p_spl_1,
    g451_n_spl_1
  );


  or

  (
    g692_n,
    g447_n_spl_1,
    g451_p_spl_1
  );


  and

  (
    g693_p,
    g691_n,
    g692_n
  );


  or

  (
    g693_n,
    g691_p,
    g692_p
  );


  and

  (
    g694_p,
    g458_n_spl_1,
    g468_n_spl_1
  );


  or

  (
    g694_n,
    g458_p_spl_1,
    g468_p_spl_1
  );


  and

  (
    g695_p,
    g458_p_spl_1,
    g468_p_spl_1
  );


  or

  (
    g695_n,
    g458_n_spl_1,
    g468_n_spl_1
  );


  and

  (
    g696_p,
    g694_n,
    g695_n
  );


  or

  (
    g696_n,
    g694_p,
    g695_p
  );


  and

  (
    g697_p,
    g693_n_spl_,
    g696_n_spl_
  );


  or

  (
    g697_n,
    g693_p_spl_,
    g696_p_spl_
  );


  and

  (
    g698_p,
    g693_p_spl_,
    g696_p_spl_
  );


  or

  (
    g698_n,
    g693_n_spl_,
    g696_n_spl_
  );


  and

  (
    g699_p,
    g697_n,
    g698_n
  );


  or

  (
    g699_n,
    g697_p,
    g698_p
  );


  and

  (
    g700_p,
    g690_p_spl_,
    g699_n_spl_
  );


  or

  (
    g700_n,
    g690_n_spl_,
    g699_p_spl_
  );


  and

  (
    g701_p,
    g690_n_spl_,
    g699_p_spl_
  );


  or

  (
    g701_n,
    g690_p_spl_,
    g699_n_spl_
  );


  and

  (
    g702_p,
    g700_n,
    g701_n
  );


  or

  (
    g702_n,
    g700_p,
    g701_p
  );


  and

  (
    g703_p,
    g684_n,
    g702_p
  );


  and

  (
    g704_p,
    g684_p,
    g702_n
  );


  or

  (
    g705_n,
    g703_p,
    g704_p
  );


  and

  (
    g706_p,
    g399_n_spl_1,
    g405_n_spl_1
  );


  or

  (
    g706_n,
    g399_p_spl_1,
    g405_p_spl_1
  );


  and

  (
    g707_p,
    g399_p_spl_1,
    g405_p_spl_1
  );


  or

  (
    g707_n,
    g399_n_spl_1,
    g405_n_spl_1
  );


  and

  (
    g708_p,
    g706_n,
    g707_n
  );


  or

  (
    g708_n,
    g706_p,
    g707_p
  );


  and

  (
    g709_p,
    g412_n_spl_1,
    g419_n_spl_1
  );


  or

  (
    g709_n,
    g412_p_spl_1,
    g419_p_spl_1
  );


  and

  (
    g710_p,
    g412_p_spl_1,
    g419_p_spl_1
  );


  or

  (
    g710_n,
    g412_n_spl_1,
    g419_n_spl_1
  );


  and

  (
    g711_p,
    g709_n,
    g710_n
  );


  or

  (
    g711_n,
    g709_p,
    g710_p
  );


  and

  (
    g712_p,
    g708_p_spl_,
    g711_n_spl_
  );


  or

  (
    g712_n,
    g708_n_spl_,
    g711_p_spl_
  );


  and

  (
    g713_p,
    g708_n_spl_,
    g711_p_spl_
  );


  or

  (
    g713_n,
    g708_p_spl_,
    g711_n_spl_
  );


  and

  (
    g714_p,
    g712_n,
    g713_n
  );


  or

  (
    g714_n,
    g712_p,
    g713_p
  );


  and

  (
    g715_p,
    G112_n,
    G124_n_spl_111
  );


  or

  (
    g715_n,
    G112_p,
    G124_p_spl_111
  );


  and

  (
    g716_p,
    G111_n_spl_,
    G124_p_spl_111
  );


  or

  (
    g716_n,
    G111_p_spl_,
    G124_n_spl_111
  );


  and

  (
    g717_p,
    g715_n,
    g716_n
  );


  or

  (
    g717_n,
    g715_p,
    g716_p
  );


  and

  (
    g718_p,
    g392_n_spl_1,
    g717_n_spl_
  );


  or

  (
    g718_n,
    g392_p_spl_1,
    g717_p_spl_
  );


  and

  (
    g719_p,
    g392_p_spl_1,
    g717_p_spl_
  );


  or

  (
    g719_n,
    g392_n_spl_1,
    g717_n_spl_
  );


  and

  (
    g720_p,
    g718_n,
    g719_n
  );


  or

  (
    g720_n,
    g718_p,
    g719_p
  );


  and

  (
    g721_p,
    g372_n_spl_1,
    g426_n_spl_1
  );


  or

  (
    g721_n,
    g372_p_spl_1,
    g426_p_spl_1
  );


  and

  (
    g722_p,
    g372_p_spl_1,
    g426_p_spl_1
  );


  or

  (
    g722_n,
    g372_n_spl_1,
    g426_n_spl_1
  );


  and

  (
    g723_p,
    g721_n,
    g722_n
  );


  or

  (
    g723_n,
    g721_p,
    g722_p
  );


  and

  (
    g724_p,
    g720_p_spl_,
    g723_n_spl_
  );


  or

  (
    g724_n,
    g720_n_spl_,
    g723_p_spl_
  );


  and

  (
    g725_p,
    g720_n_spl_,
    g723_p_spl_
  );


  or

  (
    g725_n,
    g720_p_spl_,
    g723_n_spl_
  );


  and

  (
    g726_p,
    g724_n,
    g725_n
  );


  or

  (
    g726_n,
    g724_p,
    g725_p
  );


  and

  (
    g727_p,
    g378_n_spl_1,
    g385_n_spl_1
  );


  or

  (
    g727_n,
    g378_p_spl_1,
    g385_p_spl_1
  );


  and

  (
    g728_p,
    g378_p_spl_1,
    g385_p_spl_1
  );


  or

  (
    g728_n,
    g378_n_spl_1,
    g385_n_spl_1
  );


  and

  (
    g729_p,
    g727_n,
    g728_n
  );


  or

  (
    g729_n,
    g727_p,
    g728_p
  );


  and

  (
    g730_p,
    g726_n_spl_,
    g729_n_spl_
  );


  or

  (
    g730_n,
    g726_p_spl_,
    g729_p_spl_
  );


  and

  (
    g731_p,
    g726_p_spl_,
    g729_p_spl_
  );


  or

  (
    g731_n,
    g726_n_spl_,
    g729_n_spl_
  );


  and

  (
    g732_p,
    g730_n,
    g731_n
  );


  or

  (
    g732_n,
    g730_p,
    g731_p
  );


  and

  (
    g733_p,
    g714_n,
    g732_p
  );


  and

  (
    g734_p,
    g714_p,
    g732_n
  );


  or

  (
    g735_n,
    g733_p,
    g734_p
  );


  and

  (
    g736_p,
    G2_p_spl_1,
    g430_p_spl_0
  );


  or

  (
    g736_n,
    G2_n_spl_,
    g430_n_spl_0
  );


  and

  (
    g737_p,
    g541_p_spl_00,
    g736_n
  );


  or

  (
    g737_n,
    g541_n_spl_0,
    g736_p
  );


  and

  (
    g738_p,
    g373_p_spl_,
    g737_p_spl_00
  );


  or

  (
    g738_n,
    g373_n_spl_,
    g737_n_spl_00
  );


  and

  (
    g739_p,
    g374_p_spl_0,
    g737_n_spl_00
  );


  or

  (
    g739_n,
    g374_n_spl_0,
    g737_p_spl_00
  );


  and

  (
    g740_p,
    g738_n,
    g739_n
  );


  or

  (
    g740_n,
    g738_p,
    g739_p
  );


  or

  (
    g741_n,
    g381_n_spl_01,
    g740_p
  );


  or

  (
    g742_n,
    g381_p_spl_01,
    g740_n
  );


  and

  (
    g743_p,
    g741_n,
    g742_n
  );


  or

  (
    g744_n,
    g664_n_spl_,
    g743_p_spl_
  );


  or

  (
    g745_n,
    g375_n_spl_00,
    g737_p_spl_0
  );


  or

  (
    g746_n,
    g375_p_spl_00,
    g737_n_spl_0
  );


  and

  (
    g747_p,
    g745_n,
    g746_n
  );


  or

  (
    g748_n,
    g572_p_spl_,
    g747_p_spl_
  );


  or

  (
    g749_n,
    g744_n,
    g748_n
  );


  or

  (
    g750_n,
    g643_n_spl_,
    g652_n_spl_
  );


  and

  (
    g751_p,
    g382_p_spl_,
    g737_n_spl_1
  );


  or

  (
    g751_n,
    g382_n_spl_,
    g737_p_spl_1
  );


  and

  (
    g752_p,
    g544_p_spl_0,
    g751_n
  );


  or

  (
    g752_n,
    g544_n_spl_0,
    g751_p
  );


  or

  (
    g753_n,
    g388_n_spl_00,
    g752_n
  );


  or

  (
    g754_n,
    g388_p_spl_00,
    g752_p
  );


  and

  (
    g755_p,
    g753_n,
    g754_n
  );


  and

  (
    g756_p,
    g389_p_spl_,
    g737_n_spl_1
  );


  or

  (
    g756_n,
    g389_n_spl_0,
    g737_p_spl_1
  );


  and

  (
    g757_p,
    g546_p_spl_0,
    g756_n
  );


  or

  (
    g757_n,
    g546_n_spl_0,
    g756_p
  );


  or

  (
    g758_n,
    g395_n_spl_01,
    g757_n
  );


  or

  (
    g759_n,
    g395_p_spl_00,
    g757_p
  );


  and

  (
    g760_p,
    g758_n,
    g759_n
  );


  or

  (
    g761_n,
    g755_p_spl_,
    g760_p_spl_
  );


  or

  (
    g762_n,
    g673_n_spl_,
    g761_n
  );


  or

  (
    g763_n,
    g750_n,
    g762_n
  );


  or

  (
    g764_n,
    g749_n,
    g763_n
  );


  or

  (
    g765_n,
    g601_p_spl_,
    g619_n_spl_
  );


  or

  (
    g766_n,
    g553_p_spl_,
    g581_n_spl_01
  );


  or

  (
    g767_n,
    g610_n_spl_,
    g766_n
  );


  or

  (
    g768_n,
    g765_n,
    g767_n
  );


  and

  (
    g769_p,
    g469_n_spl_,
    g594_n_spl_
  );


  or

  (
    g769_n,
    g469_p_spl_,
    g594_p_spl_
  );


  and

  (
    g770_p,
    g454_p_spl_1,
    g769_n
  );


  or

  (
    g770_n,
    g454_n_spl_1,
    g769_p
  );


  and

  (
    g771_p,
    g452_n_spl_,
    g770_n
  );


  or

  (
    g771_n,
    g452_p_spl_,
    g770_p
  );


  and

  (
    g772_p,
    g450_p_spl_1,
    g771_n
  );


  or

  (
    g772_n,
    g450_n_spl_1,
    g771_p
  );


  and

  (
    g773_p,
    g473_n,
    g772_n
  );


  or

  (
    g773_n,
    g473_p_spl_,
    g772_p
  );


  and

  (
    g774_p,
    g448_n_spl_,
    g773_p
  );


  or

  (
    g774_n,
    g448_p_spl_,
    g773_n
  );


  or

  (
    g775_n,
    g443_n_spl_00,
    g774_p_spl_00
  );


  or

  (
    g776_n,
    g443_p_spl_00,
    g774_n_spl_00
  );


  and

  (
    g777_p,
    g775_n,
    g776_n
  );


  or

  (
    g778_n,
    g562_n_spl_0,
    g777_p_spl_
  );


  and

  (
    g779_p,
    g437_p_spl_00,
    g441_p_spl_00
  );


  or

  (
    g779_n,
    g437_n_spl_00,
    g441_n_spl_00
  );


  and

  (
    g780_p,
    g435_n_spl_,
    g779_n
  );


  or

  (
    g780_n,
    g435_p_spl_,
    g779_p
  );


  and

  (
    g781_p,
    g444_p_spl_0,
    g774_n_spl_00
  );


  or

  (
    g781_n,
    g444_n_spl_,
    g774_p_spl_00
  );


  and

  (
    g782_p,
    g780_p_spl_0,
    g781_n
  );


  or

  (
    g782_n,
    g780_n_spl_0,
    g781_p
  );


  or

  (
    g783_n,
    g479_p_spl_01,
    g782_n
  );


  or

  (
    g784_n,
    g479_n_spl_01,
    g782_p
  );


  and

  (
    g785_p,
    g783_n,
    g784_n
  );


  and

  (
    g786_p,
    g441_p_spl_0,
    g774_p_spl_01
  );


  or

  (
    g786_n,
    g441_n_spl_0,
    g774_n_spl_01
  );


  and

  (
    g787_p,
    g442_p_spl_0,
    g774_n_spl_01
  );


  or

  (
    g787_n,
    g442_n_spl_0,
    g774_p_spl_01
  );


  and

  (
    g788_p,
    g786_n,
    g787_n
  );


  or

  (
    g788_n,
    g786_p,
    g787_p
  );


  or

  (
    g789_n,
    g437_n_spl_01,
    g788_p
  );


  or

  (
    g790_n,
    g437_p_spl_01,
    g788_n
  );


  and

  (
    g791_p,
    g789_n,
    g790_n
  );


  or

  (
    g792_n,
    g785_p_spl_,
    g791_p_spl_
  );


  or

  (
    g793_n,
    g778_n,
    g792_n
  );


  or

  (
    g794_n,
    g768_n,
    g793_n
  );


  and

  (
    g795_p,
    G81_p_spl_,
    G158_n_spl_0000
  );


  and

  (
    g796_p,
    G80_p_spl_,
    G158_p_spl_0000
  );


  or

  (
    g797_n,
    g795_p,
    g796_p
  );


  and

  (
    g798_p,
    G159_n_spl_000,
    g797_n
  );


  and

  (
    g799_p,
    G158_p_spl_0000,
    g560_p_spl_0
  );


  and

  (
    g800_p,
    G158_n_spl_0000,
    g579_p_spl_0
  );


  or

  (
    g801_n,
    g799_p,
    g800_p
  );


  and

  (
    g802_p,
    G159_p_spl_000,
    g801_n
  );


  or

  (
    g803_n,
    g798_p,
    g802_p
  );


  and

  (
    g804_p,
    G64_p_spl_0000,
    g803_n
  );


  and

  (
    g805_p,
    G81_p_spl_,
    G160_n_spl_0000
  );


  and

  (
    g806_p,
    G80_p_spl_,
    G160_p_spl_0000
  );


  or

  (
    g807_n,
    g805_p,
    g806_p
  );


  and

  (
    g808_p,
    G161_n_spl_000,
    g807_n
  );


  and

  (
    g809_p,
    G160_p_spl_0000,
    g560_p_spl_1
  );


  and

  (
    g810_p,
    G160_n_spl_0000,
    g579_p_spl_1
  );


  or

  (
    g811_n,
    g809_p,
    g810_p
  );


  and

  (
    g812_p,
    G161_p_spl_000,
    g811_n
  );


  or

  (
    g813_n,
    g808_p,
    g812_p
  );


  and

  (
    g814_p,
    G64_p_spl_0000,
    g813_n
  );


  and

  (
    g815_p,
    G14_p_spl_,
    G173_n_spl_0001
  );


  and

  (
    g816_p,
    G16_p_spl_,
    G173_p_spl_0001
  );


  or

  (
    g817_n,
    g815_p,
    g816_p
  );


  and

  (
    g818_p,
    G172_n_spl_000,
    g817_n
  );


  or

  (
    g819_n,
    G173_p_spl_0001,
    g647_n_spl_00
  );


  or

  (
    g820_n,
    G173_n_spl_0001,
    g605_n_spl_00
  );


  and

  (
    g821_p,
    G172_p_spl_000,
    g820_n
  );


  and

  (
    g822_p,
    g819_n,
    g821_p
  );


  or

  (
    g823_n,
    g818_p,
    g822_p
  );


  and

  (
    g824_p,
    G6_p_spl_,
    G173_n_spl_0010
  );


  and

  (
    g825_p,
    G27_p_spl_,
    G173_p_spl_0010
  );


  or

  (
    g826_n,
    g824_p,
    g825_p
  );


  and

  (
    g827_p,
    G172_n_spl_001,
    g826_n
  );


  or

  (
    g828_n,
    G173_p_spl_0010,
    g656_n_spl_00
  );


  or

  (
    g829_n,
    G173_n_spl_0010,
    g614_n_spl_00
  );


  and

  (
    g830_p,
    G172_p_spl_001,
    g829_n
  );


  and

  (
    g831_p,
    g828_n,
    g830_p
  );


  or

  (
    g832_n,
    g827_p,
    g831_p
  );


  and

  (
    g833_p,
    G5_p_spl_,
    G173_n_spl_0011
  );


  and

  (
    g834_p,
    G26_p_spl_,
    G173_p_spl_0011
  );


  or

  (
    g835_n,
    g833_p,
    g834_p
  );


  and

  (
    g836_p,
    G172_n_spl_001,
    g835_n
  );


  or

  (
    g837_n,
    G173_p_spl_0011,
    g669_n_spl_00
  );


  or

  (
    g838_n,
    G173_n_spl_0011,
    g624_n_spl_00
  );


  and

  (
    g839_p,
    G172_p_spl_001,
    g838_n
  );


  and

  (
    g840_p,
    g837_n,
    g839_p
  );


  or

  (
    g841_n,
    g836_p,
    g840_p
  );


  and

  (
    g842_p,
    G25_p_spl_,
    G173_n_spl_010
  );


  and

  (
    g843_p,
    G24_p_spl_,
    G173_p_spl_010
  );


  or

  (
    g844_n,
    g842_p,
    g843_p
  );


  and

  (
    g845_p,
    G172_n_spl_01,
    g844_n
  );


  or

  (
    g846_n,
    G173_p_spl_010,
    g678_n_spl_00
  );


  or

  (
    g847_n,
    G173_n_spl_010,
    g569_p_spl_00
  );


  and

  (
    g848_p,
    G172_p_spl_01,
    g847_n
  );


  and

  (
    g849_p,
    g846_n,
    g848_p
  );


  or

  (
    g850_n,
    g845_p,
    g849_p
  );


  and

  (
    g851_p,
    G14_p_spl_,
    G174_n_spl_0001
  );


  and

  (
    g852_p,
    G16_p_spl_,
    G174_p_spl_0001
  );


  or

  (
    g853_n,
    g851_p,
    g852_p
  );


  and

  (
    g854_p,
    G175_n_spl_000,
    g853_n
  );


  or

  (
    g855_n,
    G174_p_spl_0001,
    g647_n_spl_00
  );


  or

  (
    g856_n,
    G174_n_spl_0001,
    g605_n_spl_00
  );


  and

  (
    g857_p,
    G175_p_spl_000,
    g856_n
  );


  and

  (
    g858_p,
    g855_n,
    g857_p
  );


  or

  (
    g859_n,
    g854_p,
    g858_p
  );


  and

  (
    g860_p,
    G6_p_spl_,
    G174_n_spl_0010
  );


  and

  (
    g861_p,
    G27_p_spl_,
    G174_p_spl_0010
  );


  or

  (
    g862_n,
    g860_p,
    g861_p
  );


  and

  (
    g863_p,
    G175_n_spl_001,
    g862_n
  );


  or

  (
    g864_n,
    G174_p_spl_0010,
    g656_n_spl_00
  );


  or

  (
    g865_n,
    G174_n_spl_0010,
    g614_n_spl_00
  );


  and

  (
    g866_p,
    G175_p_spl_001,
    g865_n
  );


  and

  (
    g867_p,
    g864_n,
    g866_p
  );


  or

  (
    g868_n,
    g863_p,
    g867_p
  );


  and

  (
    g869_p,
    G5_p_spl_,
    G174_n_spl_0011
  );


  and

  (
    g870_p,
    G26_p_spl_,
    G174_p_spl_0011
  );


  or

  (
    g871_n,
    g869_p,
    g870_p
  );


  and

  (
    g872_p,
    G175_n_spl_001,
    g871_n
  );


  or

  (
    g873_n,
    G174_p_spl_0011,
    g669_n_spl_00
  );


  or

  (
    g874_n,
    G174_n_spl_0011,
    g624_n_spl_00
  );


  and

  (
    g875_p,
    G175_p_spl_001,
    g874_n
  );


  and

  (
    g876_p,
    g873_n,
    g875_p
  );


  or

  (
    g877_n,
    g872_p,
    g876_p
  );


  and

  (
    g878_p,
    G25_p_spl_,
    G174_n_spl_010
  );


  and

  (
    g879_p,
    G24_p_spl_,
    G174_p_spl_010
  );


  or

  (
    g880_n,
    g878_p,
    g879_p
  );


  and

  (
    g881_p,
    G175_n_spl_01,
    g880_n
  );


  or

  (
    g882_n,
    G174_p_spl_010,
    g678_n_spl_00
  );


  or

  (
    g883_n,
    G174_n_spl_010,
    g569_p_spl_00
  );


  and

  (
    g884_p,
    G175_p_spl_01,
    g883_n
  );


  and

  (
    g885_p,
    g882_n,
    g884_p
  );


  or

  (
    g886_n,
    g881_p,
    g885_p
  );


  and

  (
    g887_p,
    G76_p_spl_,
    G158_n_spl_0001
  );


  and

  (
    g888_p,
    G86_p_spl_,
    G158_p_spl_0001
  );


  or

  (
    g889_n,
    g887_p,
    g888_p
  );


  and

  (
    g890_p,
    G159_n_spl_000,
    g889_n
  );


  and

  (
    g891_p,
    G158_p_spl_0001,
    g605_n_spl_0
  );


  and

  (
    g892_p,
    G158_n_spl_0001,
    g647_n_spl_0
  );


  or

  (
    g893_n,
    g891_p,
    g892_p
  );


  and

  (
    g894_p,
    G159_p_spl_000,
    g893_n
  );


  or

  (
    g895_n,
    g890_p,
    g894_p
  );


  and

  (
    g896_p,
    G64_p_spl_0001,
    g895_n
  );


  and

  (
    g897_p,
    G72_p_spl_,
    G158_n_spl_0010
  );


  and

  (
    g898_p,
    G82_p_spl_,
    G158_p_spl_0010
  );


  or

  (
    g899_n,
    g897_p,
    g898_p
  );


  and

  (
    g900_p,
    G159_n_spl_001,
    g899_n
  );


  and

  (
    g901_p,
    G158_p_spl_0010,
    g569_p_spl_0
  );


  and

  (
    g902_p,
    G158_n_spl_0010,
    g678_n_spl_0
  );


  or

  (
    g903_n,
    g901_p,
    g902_p
  );


  and

  (
    g904_p,
    G159_p_spl_001,
    g903_n
  );


  or

  (
    g905_n,
    g900_p,
    g904_p
  );


  and

  (
    g906_p,
    G64_p_spl_0001,
    g905_n
  );


  and

  (
    g907_p,
    G70_p_spl_,
    G158_n_spl_0011
  );


  and

  (
    g908_p,
    G71_p_spl_,
    G158_p_spl_0011
  );


  or

  (
    g909_n,
    g907_p,
    g908_p
  );


  and

  (
    g910_p,
    G159_n_spl_001,
    g909_n
  );


  and

  (
    g911_p,
    G158_p_spl_0011,
    g624_n_spl_0
  );


  and

  (
    g912_p,
    G158_n_spl_0011,
    g669_n_spl_0
  );


  or

  (
    g913_n,
    g911_p,
    g912_p
  );


  and

  (
    g914_p,
    G159_p_spl_001,
    g913_n
  );


  or

  (
    g915_n,
    g910_p,
    g914_p
  );


  and

  (
    g916_p,
    G64_p_spl_0010,
    g915_n
  );


  and

  (
    g917_p,
    G68_p_spl_,
    G158_n_spl_010
  );


  and

  (
    g918_p,
    G69_p_spl_,
    G158_p_spl_010
  );


  or

  (
    g919_n,
    g917_p,
    g918_p
  );


  and

  (
    g920_p,
    G159_n_spl_01,
    g919_n
  );


  and

  (
    g921_p,
    G158_p_spl_010,
    g614_n_spl_0
  );


  and

  (
    g922_p,
    G158_n_spl_010,
    g656_n_spl_0
  );


  or

  (
    g923_n,
    g921_p,
    g922_p
  );


  and

  (
    g924_p,
    G159_p_spl_01,
    g923_n
  );


  or

  (
    g925_n,
    g920_p,
    g924_p
  );


  and

  (
    g926_p,
    G64_p_spl_0010,
    g925_n
  );


  and

  (
    g927_p,
    G76_p_spl_,
    G160_n_spl_0001
  );


  and

  (
    g928_p,
    G86_p_spl_,
    G160_p_spl_0001
  );


  or

  (
    g929_n,
    g927_p,
    g928_p
  );


  and

  (
    g930_p,
    G161_n_spl_000,
    g929_n
  );


  and

  (
    g931_p,
    G160_p_spl_0001,
    g605_n_spl_1
  );


  and

  (
    g932_p,
    G160_n_spl_0001,
    g647_n_spl_1
  );


  or

  (
    g933_n,
    g931_p,
    g932_p
  );


  and

  (
    g934_p,
    G161_p_spl_000,
    g933_n
  );


  or

  (
    g935_n,
    g930_p,
    g934_p
  );


  and

  (
    g936_p,
    G64_p_spl_001,
    g935_n
  );


  and

  (
    g937_p,
    G72_p_spl_,
    G160_n_spl_0010
  );


  and

  (
    g938_p,
    G82_p_spl_,
    G160_p_spl_0010
  );


  or

  (
    g939_n,
    g937_p,
    g938_p
  );


  and

  (
    g940_p,
    G161_n_spl_001,
    g939_n
  );


  and

  (
    g941_p,
    G160_p_spl_0010,
    g569_p_spl_1
  );


  and

  (
    g942_p,
    G160_n_spl_0010,
    g678_n_spl_1
  );


  or

  (
    g943_n,
    g941_p,
    g942_p
  );


  and

  (
    g944_p,
    G161_p_spl_001,
    g943_n
  );


  or

  (
    g945_n,
    g940_p,
    g944_p
  );


  and

  (
    g946_p,
    G64_p_spl_010,
    g945_n
  );


  and

  (
    g947_p,
    G70_p_spl_,
    G160_n_spl_0011
  );


  and

  (
    g948_p,
    G71_p_spl_,
    G160_p_spl_0011
  );


  or

  (
    g949_n,
    g947_p,
    g948_p
  );


  and

  (
    g950_p,
    G161_n_spl_001,
    g949_n
  );


  and

  (
    g951_p,
    G160_p_spl_0011,
    g624_n_spl_1
  );


  and

  (
    g952_p,
    G160_n_spl_0011,
    g669_n_spl_1
  );


  or

  (
    g953_n,
    g951_p,
    g952_p
  );


  and

  (
    g954_p,
    G161_p_spl_001,
    g953_n
  );


  or

  (
    g955_n,
    g950_p,
    g954_p
  );


  and

  (
    g956_p,
    G64_p_spl_010,
    g955_n
  );


  and

  (
    g957_p,
    G68_p_spl_,
    G160_n_spl_010
  );


  and

  (
    g958_p,
    G69_p_spl_,
    G160_p_spl_010
  );


  or

  (
    g959_n,
    g957_p,
    g958_p
  );


  and

  (
    g960_p,
    G161_n_spl_01,
    g959_n
  );


  and

  (
    g961_p,
    G160_p_spl_010,
    g614_n_spl_1
  );


  and

  (
    g962_p,
    G160_n_spl_010,
    g656_n_spl_1
  );


  or

  (
    g963_n,
    g961_p,
    g962_p
  );


  and

  (
    g964_p,
    G161_p_spl_01,
    g963_n
  );


  or

  (
    g965_n,
    g960_p,
    g964_p
  );


  and

  (
    g966_p,
    G64_p_spl_011,
    g965_n
  );


  or

  (
    g967_n,
    G62_n,
    G178_n
  );


  and

  (
    g968_p,
    G171_p_spl_,
    g581_n_spl_01
  );


  and

  (
    g969_p,
    G54_p_spl_,
    G171_n_spl_
  );


  or

  (
    g970_n,
    g968_p,
    g969_p
  );


  and

  (
    g971_p,
    G170_p,
    g970_n
  );


  and

  (
    g972_p,
    G171_n_spl_,
    g237_n_spl_0
  );


  and

  (
    g973_p,
    G61_n_spl_,
    g476_n_spl_1
  );


  or

  (
    g973_n,
    G61_p_spl_,
    g476_p_spl_1
  );


  and

  (
    g974_p,
    G61_p_spl_,
    g476_p_spl_1
  );


  or

  (
    g974_n,
    G61_n_spl_,
    g476_n_spl_1
  );


  and

  (
    g975_p,
    g973_n,
    g974_n
  );


  or

  (
    g975_n,
    g973_p,
    g974_p
  );


  and

  (
    g976_p,
    G171_p_spl_,
    g975_p_spl_
  );


  or

  (
    g977_n,
    g972_p,
    g976_p
  );


  and

  (
    g978_p,
    G170_n,
    g977_n
  );


  or

  (
    g979_n,
    g971_p,
    g978_p
  );


  and

  (
    g980_p,
    g967_n,
    g979_n
  );


  and

  (
    g981_p,
    g581_n_spl_10,
    g975_n
  );


  and

  (
    g982_p,
    g581_p_spl_01,
    g975_p_spl_
  );


  or

  (
    g983_n,
    g981_p,
    g982_p
  );


  and

  (
    g984_p,
    G177_p_spl_0110,
    g581_n_spl_10
  );


  or

  (
    g985_n,
    G176_p_spl_0111,
    g984_p
  );


  or

  (
    g986_n,
    G177_n_spl_011,
    g237_n_spl_1
  );


  or

  (
    g987_n,
    G176_n_spl_0101,
    g986_n
  );


  or

  (
    g988_n,
    G54_p_spl_,
    G177_p_spl_0111
  );


  and

  (
    g989_p,
    g987_n,
    g988_n
  );


  and

  (
    g990_p,
    g985_n,
    g989_p
  );


  and

  (
    g991_p,
    G52_p,
    G177_n_spl_011
  );


  and

  (
    g992_p,
    G176_p_spl_1000,
    g991_p
  );


  or

  (
    g993_n,
    G176_p_spl_1000,
    g785_p_spl_
  );


  or

  (
    g994_n,
    G176_n_spl_0101,
    g240_n_spl_0
  );


  and

  (
    g995_p,
    G177_p_spl_0111,
    g994_n
  );


  and

  (
    g996_p,
    g993_n,
    g995_p
  );


  or

  (
    g997_n,
    g992_p,
    g996_p
  );


  and

  (
    g998_p,
    G47_p,
    G177_n_spl_100
  );


  and

  (
    g999_p,
    G176_p_spl_1001,
    g998_p
  );


  or

  (
    g1000_n,
    G176_p_spl_1001,
    g791_p_spl_
  );


  or

  (
    g1001_n,
    G176_n_spl_011,
    g267_n_spl_0
  );


  and

  (
    g1002_p,
    G177_p_spl_1000,
    g1001_n
  );


  and

  (
    g1003_p,
    g1000_n,
    g1002_p
  );


  or

  (
    g1004_n,
    g999_p,
    g1003_p
  );


  and

  (
    g1005_p,
    G43_p,
    G177_n_spl_100
  );


  and

  (
    g1006_p,
    G176_p_spl_1010,
    g1005_p
  );


  or

  (
    g1007_n,
    G176_n_spl_011,
    g258_n_spl_0
  );


  or

  (
    g1008_n,
    G176_p_spl_1010,
    g777_p_spl_
  );


  and

  (
    g1009_p,
    G177_p_spl_1000,
    g1008_n
  );


  and

  (
    g1010_p,
    g1007_n,
    g1009_p
  );


  or

  (
    g1011_n,
    g1006_p,
    g1010_p
  );


  or

  (
    g1012_n,
    G99_n_spl_,
    g533_n_spl_
  );


  or

  (
    g1013_n,
    g735_n_spl_,
    g1012_n
  );


  or

  (
    g1014_n,
    G155_n_spl_,
    g184_n_spl_
  );


  or

  (
    g1015_n,
    g179_n_spl_,
    g1014_n
  );


  or

  (
    g1016_n,
    g705_n_spl_,
    g1015_n
  );


  or

  (
    g1017_n,
    g506_n_spl_,
    g1016_n
  );


  or

  (
    g1018_n,
    g1013_n,
    g1017_n
  );


  and

  (
    g1019_p,
    G46_p,
    G177_n_spl_101
  );


  and

  (
    g1020_p,
    G176_p_spl_1011,
    g1019_p
  );


  or

  (
    g1021_n,
    G176_p_spl_1011,
    g760_p_spl_
  );


  or

  (
    g1022_n,
    G176_n_spl_100,
    g317_n_spl_0
  );


  and

  (
    g1023_p,
    G177_p_spl_1001,
    g1022_n
  );


  and

  (
    g1024_p,
    g1021_n,
    g1023_p
  );


  or

  (
    g1025_n,
    g1020_p,
    g1024_p
  );


  and

  (
    g1026_p,
    G45_p,
    G177_n_spl_101
  );


  and

  (
    g1027_p,
    G176_p_spl_1100,
    g1026_p
  );


  or

  (
    g1028_n,
    G176_p_spl_1100,
    g755_p_spl_
  );


  or

  (
    g1029_n,
    G176_n_spl_100,
    g328_n_spl_
  );


  and

  (
    g1030_p,
    G177_p_spl_1001,
    g1029_n
  );


  and

  (
    g1031_p,
    g1028_n,
    g1030_p
  );


  or

  (
    g1032_n,
    g1027_p,
    g1031_p
  );


  and

  (
    g1033_p,
    G20_p,
    G177_n_spl_110
  );


  and

  (
    g1034_p,
    G176_p_spl_1101,
    g1033_p
  );


  or

  (
    g1035_n,
    G176_p_spl_1101,
    g743_p_spl_
  );


  or

  (
    g1036_n,
    G176_n_spl_101,
    g337_n_spl_
  );


  and

  (
    g1037_p,
    G177_p_spl_101,
    g1036_n
  );


  and

  (
    g1038_p,
    g1035_n,
    g1037_p
  );


  or

  (
    g1039_n,
    g1034_p,
    g1038_p
  );


  and

  (
    g1040_p,
    G44_p,
    G177_n_spl_110
  );


  and

  (
    g1041_p,
    G176_p_spl_1110,
    g1040_p
  );


  or

  (
    g1042_n,
    G176_p_spl_1110,
    g747_p_spl_
  );


  or

  (
    g1043_n,
    G176_n_spl_101,
    g347_n_spl_
  );


  and

  (
    g1044_p,
    G177_p_spl_101,
    g1043_n
  );


  and

  (
    g1045_p,
    g1042_n,
    g1044_p
  );


  or

  (
    g1046_n,
    g1041_p,
    g1045_p
  );


  or

  (
    g1047_n,
    G174_p_spl_011,
    g1025_n_spl_00
  );


  or

  (
    g1048_n,
    G174_n_spl_011,
    g990_p_spl_00
  );


  and

  (
    g1049_p,
    G175_p_spl_01,
    g1048_n
  );


  and

  (
    g1050_p,
    g1047_n,
    g1049_p
  );


  and

  (
    g1051_p,
    G41_p_spl_,
    G174_n_spl_011
  );


  and

  (
    g1052_p,
    G42_p_spl_,
    G174_p_spl_011
  );


  or

  (
    g1053_n,
    g1051_p,
    g1052_p
  );


  and

  (
    g1054_p,
    G175_n_spl_01,
    g1053_n
  );


  or

  (
    g1055_n,
    g1050_p,
    g1054_p
  );


  or

  (
    g1056_n,
    G173_p_spl_011,
    g1025_n_spl_00
  );


  or

  (
    g1057_n,
    G173_n_spl_011,
    g990_p_spl_00
  );


  and

  (
    g1058_p,
    G172_p_spl_01,
    g1057_n
  );


  and

  (
    g1059_p,
    g1056_n,
    g1058_p
  );


  and

  (
    g1060_p,
    G41_p_spl_,
    G173_n_spl_011
  );


  and

  (
    g1061_p,
    G42_p_spl_,
    G173_p_spl_011
  );


  or

  (
    g1062_n,
    g1060_p,
    g1061_p
  );


  and

  (
    g1063_p,
    G172_n_spl_01,
    g1062_n
  );


  or

  (
    g1064_n,
    g1059_p,
    g1063_p
  );


  and

  (
    g1065_p,
    G18_p_spl_,
    G173_n_spl_100
  );


  and

  (
    g1066_p,
    G17_p_spl_,
    G173_p_spl_100
  );


  or

  (
    g1067_n,
    g1065_p,
    g1066_p
  );


  and

  (
    g1068_p,
    G172_n_spl_10,
    g1067_n
  );


  or

  (
    g1069_n,
    G173_p_spl_100,
    g1032_n_spl_00
  );


  or

  (
    g1070_n,
    G173_n_spl_100,
    g997_n_spl_00
  );


  and

  (
    g1071_p,
    G172_p_spl_10,
    g1070_n
  );


  and

  (
    g1072_p,
    g1069_n,
    g1071_p
  );


  or

  (
    g1073_n,
    g1068_p,
    g1072_p
  );


  and

  (
    g1074_p,
    G40_p_spl_,
    G173_n_spl_101
  );


  and

  (
    g1075_p,
    G39_p_spl_,
    G173_p_spl_101
  );


  or

  (
    g1076_n,
    g1074_p,
    g1075_p
  );


  and

  (
    g1077_p,
    G172_n_spl_10,
    g1076_n
  );


  or

  (
    g1078_n,
    G173_p_spl_101,
    g1039_n_spl_00
  );


  or

  (
    g1079_n,
    G173_n_spl_101,
    g1004_n_spl_00
  );


  and

  (
    g1080_p,
    G172_p_spl_10,
    g1079_n
  );


  and

  (
    g1081_p,
    g1078_n,
    g1080_p
  );


  or

  (
    g1082_n,
    g1077_p,
    g1081_p
  );


  and

  (
    g1083_p,
    G15_p_spl_,
    G173_n_spl_110
  );


  and

  (
    g1084_p,
    G36_p_spl_,
    G173_p_spl_110
  );


  or

  (
    g1085_n,
    g1083_p,
    g1084_p
  );


  and

  (
    g1086_p,
    G172_n_spl_11,
    g1085_n
  );


  or

  (
    g1087_n,
    G173_p_spl_110,
    g1046_n_spl_00
  );


  or

  (
    g1088_n,
    G173_n_spl_110,
    g1011_n_spl_00
  );


  and

  (
    g1089_p,
    G172_p_spl_11,
    g1088_n
  );


  and

  (
    g1090_p,
    g1087_n,
    g1089_p
  );


  or

  (
    g1091_n,
    g1086_p,
    g1090_p
  );


  and

  (
    g1092_p,
    G18_p_spl_,
    G174_n_spl_100
  );


  and

  (
    g1093_p,
    G17_p_spl_,
    G174_p_spl_100
  );


  or

  (
    g1094_n,
    g1092_p,
    g1093_p
  );


  and

  (
    g1095_p,
    G175_n_spl_10,
    g1094_n
  );


  or

  (
    g1096_n,
    G174_p_spl_100,
    g1032_n_spl_00
  );


  or

  (
    g1097_n,
    G174_n_spl_100,
    g997_n_spl_00
  );


  and

  (
    g1098_p,
    G175_p_spl_10,
    g1097_n
  );


  and

  (
    g1099_p,
    g1096_n,
    g1098_p
  );


  or

  (
    g1100_n,
    g1095_p,
    g1099_p
  );


  and

  (
    g1101_p,
    G40_p_spl_,
    G174_n_spl_101
  );


  and

  (
    g1102_p,
    G39_p_spl_,
    G174_p_spl_101
  );


  or

  (
    g1103_n,
    g1101_p,
    g1102_p
  );


  and

  (
    g1104_p,
    G175_n_spl_10,
    g1103_n
  );


  or

  (
    g1105_n,
    G174_p_spl_101,
    g1039_n_spl_00
  );


  or

  (
    g1106_n,
    G174_n_spl_101,
    g1004_n_spl_00
  );


  and

  (
    g1107_p,
    G175_p_spl_10,
    g1106_n
  );


  and

  (
    g1108_p,
    g1105_n,
    g1107_p
  );


  or

  (
    g1109_n,
    g1104_p,
    g1108_p
  );


  and

  (
    g1110_p,
    G15_p_spl_,
    G174_n_spl_110
  );


  and

  (
    g1111_p,
    G36_p_spl_,
    G174_p_spl_110
  );


  or

  (
    g1112_n,
    g1110_p,
    g1111_p
  );


  and

  (
    g1113_p,
    G175_n_spl_11,
    g1112_n
  );


  or

  (
    g1114_n,
    G174_p_spl_110,
    g1046_n_spl_00
  );


  or

  (
    g1115_n,
    G174_n_spl_110,
    g1011_n_spl_00
  );


  and

  (
    g1116_p,
    G175_p_spl_11,
    g1115_n
  );


  and

  (
    g1117_p,
    g1114_n,
    g1116_p
  );


  or

  (
    g1118_n,
    g1113_p,
    g1117_p
  );


  and

  (
    g1119_p,
    G77_p_spl_,
    G158_n_spl_011
  );


  and

  (
    g1120_p,
    G87_p_spl_,
    G158_p_spl_011
  );


  or

  (
    g1121_n,
    g1119_p,
    g1120_p
  );


  and

  (
    g1122_p,
    G159_n_spl_01,
    g1121_n
  );


  and

  (
    g1123_p,
    G158_p_spl_011,
    g1011_n_spl_0
  );


  and

  (
    g1124_p,
    G158_n_spl_011,
    g1046_n_spl_0
  );


  or

  (
    g1125_n,
    g1123_p,
    g1124_p
  );


  and

  (
    g1126_p,
    G159_p_spl_01,
    g1125_n
  );


  or

  (
    g1127_n,
    g1122_p,
    g1126_p
  );


  and

  (
    g1128_p,
    G64_p_spl_011,
    g1127_n
  );


  and

  (
    g1129_p,
    G75_p_spl_,
    G158_n_spl_100
  );


  and

  (
    g1130_p,
    G85_p_spl_,
    G158_p_spl_100
  );


  or

  (
    g1131_n,
    g1129_p,
    g1130_p
  );


  and

  (
    g1132_p,
    G159_n_spl_10,
    g1131_n
  );


  and

  (
    g1133_p,
    G158_p_spl_100,
    g1004_n_spl_0
  );


  and

  (
    g1134_p,
    G158_n_spl_100,
    g1039_n_spl_0
  );


  or

  (
    g1135_n,
    g1133_p,
    g1134_p
  );


  and

  (
    g1136_p,
    G159_p_spl_10,
    g1135_n
  );


  or

  (
    g1137_n,
    g1132_p,
    g1136_p
  );


  and

  (
    g1138_p,
    G64_p_spl_100,
    g1137_n
  );


  and

  (
    g1139_p,
    G74_p_spl_,
    G158_n_spl_101
  );


  and

  (
    g1140_p,
    G84_p_spl_,
    G158_p_spl_101
  );


  or

  (
    g1141_n,
    g1139_p,
    g1140_p
  );


  and

  (
    g1142_p,
    G159_n_spl_10,
    g1141_n
  );


  and

  (
    g1143_p,
    G158_p_spl_101,
    g997_n_spl_0
  );


  and

  (
    g1144_p,
    G158_n_spl_101,
    g1032_n_spl_0
  );


  or

  (
    g1145_n,
    g1143_p,
    g1144_p
  );


  and

  (
    g1146_p,
    G159_p_spl_10,
    g1145_n
  );


  or

  (
    g1147_n,
    g1142_p,
    g1146_p
  );


  and

  (
    g1148_p,
    G64_p_spl_100,
    g1147_n
  );


  or

  (
    g1149_n,
    G158_p_spl_110,
    g1025_n_spl_0
  );


  or

  (
    g1150_n,
    G158_n_spl_110,
    g990_p_spl_0
  );


  and

  (
    g1151_p,
    G159_p_spl_11,
    g1150_n
  );


  and

  (
    g1152_p,
    g1149_n,
    g1151_p
  );


  and

  (
    g1153_p,
    G73_p_spl_,
    G158_n_spl_110
  );


  and

  (
    g1154_p,
    G83_p_spl_,
    G158_p_spl_110
  );


  or

  (
    g1155_n,
    g1153_p,
    g1154_p
  );


  and

  (
    g1156_p,
    G159_n_spl_11,
    g1155_n
  );


  or

  (
    g1157_n,
    g1152_p,
    g1156_p
  );


  and

  (
    g1158_p,
    G64_p_spl_101,
    g1157_n
  );


  and

  (
    g1159_p,
    G77_p_spl_,
    G160_n_spl_011
  );


  and

  (
    g1160_p,
    G87_p_spl_,
    G160_p_spl_011
  );


  or

  (
    g1161_n,
    g1159_p,
    g1160_p
  );


  and

  (
    g1162_p,
    G161_n_spl_01,
    g1161_n
  );


  and

  (
    g1163_p,
    G160_p_spl_011,
    g1011_n_spl_1
  );


  and

  (
    g1164_p,
    G160_n_spl_011,
    g1046_n_spl_1
  );


  or

  (
    g1165_n,
    g1163_p,
    g1164_p
  );


  and

  (
    g1166_p,
    G161_p_spl_01,
    g1165_n
  );


  or

  (
    g1167_n,
    g1162_p,
    g1166_p
  );


  and

  (
    g1168_p,
    G64_p_spl_101,
    g1167_n
  );


  and

  (
    g1169_p,
    G75_p_spl_,
    G160_n_spl_100
  );


  and

  (
    g1170_p,
    G85_p_spl_,
    G160_p_spl_100
  );


  or

  (
    g1171_n,
    g1169_p,
    g1170_p
  );


  and

  (
    g1172_p,
    G161_n_spl_10,
    g1171_n
  );


  and

  (
    g1173_p,
    G160_p_spl_100,
    g1004_n_spl_1
  );


  and

  (
    g1174_p,
    G160_n_spl_100,
    g1039_n_spl_1
  );


  or

  (
    g1175_n,
    g1173_p,
    g1174_p
  );


  and

  (
    g1176_p,
    G161_p_spl_10,
    g1175_n
  );


  or

  (
    g1177_n,
    g1172_p,
    g1176_p
  );


  and

  (
    g1178_p,
    G64_p_spl_110,
    g1177_n
  );


  and

  (
    g1179_p,
    G74_p_spl_,
    G160_n_spl_101
  );


  and

  (
    g1180_p,
    G84_p_spl_,
    G160_p_spl_101
  );


  or

  (
    g1181_n,
    g1179_p,
    g1180_p
  );


  and

  (
    g1182_p,
    G161_n_spl_10,
    g1181_n
  );


  and

  (
    g1183_p,
    G160_p_spl_101,
    g997_n_spl_1
  );


  and

  (
    g1184_p,
    G160_n_spl_101,
    g1032_n_spl_1
  );


  or

  (
    g1185_n,
    g1183_p,
    g1184_p
  );


  and

  (
    g1186_p,
    G161_p_spl_10,
    g1185_n
  );


  or

  (
    g1187_n,
    g1182_p,
    g1186_p
  );


  and

  (
    g1188_p,
    G64_p_spl_110,
    g1187_n
  );


  or

  (
    g1189_n,
    G160_p_spl_110,
    g1025_n_spl_1
  );


  or

  (
    g1190_n,
    G160_n_spl_110,
    g990_p_spl_1
  );


  and

  (
    g1191_p,
    G161_p_spl_11,
    g1190_n
  );


  and

  (
    g1192_p,
    g1189_n,
    g1191_p
  );


  and

  (
    g1193_p,
    G73_p_spl_,
    G160_n_spl_110
  );


  and

  (
    g1194_p,
    G83_p_spl_,
    G160_p_spl_110
  );


  or

  (
    g1195_n,
    g1193_p,
    g1194_p
  );


  and

  (
    g1196_p,
    G161_n_spl_11,
    g1195_n
  );


  or

  (
    g1197_n,
    g1192_p,
    g1196_p
  );


  and

  (
    g1198_p,
    G64_p_spl_111,
    g1197_n
  );


  and

  (
    g1199_p,
    g258_n_spl_,
    g267_n_spl_
  );


  or

  (
    g1199_n,
    g258_p_spl_,
    g267_p_spl_
  );


  and

  (
    g1200_p,
    g268_n_spl_,
    g1199_n
  );


  or

  (
    g1200_n,
    g268_p,
    g1199_p
  );


  and

  (
    g1201_p,
    g237_p_spl_,
    g240_n_spl_
  );


  or

  (
    g1201_n,
    g237_n_spl_1,
    g240_p_spl_
  );


  and

  (
    g1202_p,
    g241_n_spl_,
    g1201_n
  );


  or

  (
    g1202_n,
    g241_p,
    g1201_p
  );


  and

  (
    g1203_p,
    g1200_p_spl_,
    g1202_n_spl_
  );


  or

  (
    g1203_n,
    g1200_n_spl_,
    g1202_p_spl_
  );


  and

  (
    g1204_p,
    g1200_n_spl_,
    g1202_p_spl_
  );


  or

  (
    g1204_n,
    g1200_p_spl_,
    g1202_n_spl_
  );


  and

  (
    g1205_p,
    g1203_n,
    g1204_n
  );


  or

  (
    g1205_n,
    g1203_p,
    g1204_p
  );


  and

  (
    g1206_p,
    G101_p_spl_010,
    G128_p_spl_10
  );


  or

  (
    g1206_n,
    G101_n_spl_010,
    G128_n_spl_10
  );


  and

  (
    g1207_p,
    G100_p_spl_010,
    G128_n_spl_10
  );


  or

  (
    g1207_n,
    G100_n_spl_010,
    G128_p_spl_10
  );


  and

  (
    g1208_p,
    g1206_n,
    g1207_n
  );


  or

  (
    g1208_n,
    g1206_p,
    g1207_p
  );


  and

  (
    g1209_p,
    G150_p_spl_1,
    g1208_n
  );


  or

  (
    g1209_n,
    G150_n_spl_1,
    g1208_p
  );


  and

  (
    g1210_p,
    G102_n_spl_010,
    G128_p_spl_11
  );


  or

  (
    g1210_n,
    G102_p_spl_010,
    G128_n_spl_11
  );


  and

  (
    g1211_p,
    G98_n_spl_010,
    G128_n_spl_11
  );


  or

  (
    g1211_n,
    G98_p_spl_010,
    G128_p_spl_11
  );


  and

  (
    g1212_p,
    g1210_n,
    g1211_n
  );


  or

  (
    g1212_n,
    g1210_p,
    g1211_p
  );


  and

  (
    g1213_p,
    G150_n_spl_1,
    g1212_n
  );


  or

  (
    g1213_n,
    G150_p_spl_1,
    g1212_p
  );


  and

  (
    g1214_p,
    g1209_n,
    g1213_n
  );


  or

  (
    g1214_n,
    g1209_p,
    g1213_p
  );


  and

  (
    g1215_p,
    G101_p_spl_011,
    G126_p_spl_10
  );


  or

  (
    g1215_n,
    G101_n_spl_011,
    G126_n_spl_10
  );


  and

  (
    g1216_p,
    G100_p_spl_010,
    G126_n_spl_10
  );


  or

  (
    g1216_n,
    G100_n_spl_010,
    G126_p_spl_10
  );


  and

  (
    g1217_p,
    g1215_n,
    g1216_n
  );


  or

  (
    g1217_n,
    g1215_p,
    g1216_p
  );


  and

  (
    g1218_p,
    G149_p_spl_1,
    g1217_n
  );


  or

  (
    g1218_n,
    G149_n_spl_1,
    g1217_p
  );


  and

  (
    g1219_p,
    G102_n_spl_010,
    G126_p_spl_11
  );


  or

  (
    g1219_n,
    G102_p_spl_010,
    G126_n_spl_11
  );


  and

  (
    g1220_p,
    G98_n_spl_010,
    G126_n_spl_11
  );


  or

  (
    g1220_n,
    G98_p_spl_010,
    G126_p_spl_11
  );


  and

  (
    g1221_p,
    g1219_n,
    g1220_n
  );


  or

  (
    g1221_n,
    g1219_p,
    g1220_p
  );


  and

  (
    g1222_p,
    G149_n_spl_1,
    g1221_n
  );


  or

  (
    g1222_n,
    G149_p_spl_1,
    g1221_p
  );


  and

  (
    g1223_p,
    g1218_n,
    g1222_n
  );


  or

  (
    g1223_n,
    g1218_p,
    g1222_p
  );


  and

  (
    g1224_p,
    g1214_n_spl_,
    g1223_p_spl_
  );


  or

  (
    g1224_n,
    g1214_p_spl_,
    g1223_n_spl_
  );


  and

  (
    g1225_p,
    g1214_p_spl_,
    g1223_n_spl_
  );


  or

  (
    g1225_n,
    g1214_n_spl_,
    g1223_p_spl_
  );


  and

  (
    g1226_p,
    g1224_n,
    g1225_n
  );


  or

  (
    g1226_n,
    g1224_p,
    g1225_p
  );


  and

  (
    g1227_p,
    G98_n_spl_011,
    G148_n_spl_1
  );


  or

  (
    g1227_n,
    G98_p_spl_011,
    G148_p_spl_1
  );


  and

  (
    g1228_p,
    G100_p_spl_011,
    G148_p_spl_1
  );


  or

  (
    g1228_n,
    G100_n_spl_011,
    G148_n_spl_1
  );


  and

  (
    g1229_p,
    g1227_n,
    g1228_n
  );


  or

  (
    g1229_n,
    g1227_p,
    g1228_p
  );


  and

  (
    g1230_p,
    G101_p_spl_011,
    G121_p_spl_10
  );


  or

  (
    g1230_n,
    G101_n_spl_011,
    G121_n_spl_10
  );


  and

  (
    g1231_p,
    G100_p_spl_011,
    G121_n_spl_10
  );


  or

  (
    g1231_n,
    G100_n_spl_011,
    G121_p_spl_10
  );


  and

  (
    g1232_p,
    g1230_n,
    g1231_n
  );


  or

  (
    g1232_n,
    g1230_p,
    g1231_p
  );


  and

  (
    g1233_p,
    G147_p_spl_1,
    g1232_n
  );


  or

  (
    g1233_n,
    G147_n_spl_1,
    g1232_p
  );


  and

  (
    g1234_p,
    G102_n_spl_011,
    G121_p_spl_11
  );


  or

  (
    g1234_n,
    G102_p_spl_011,
    G121_n_spl_11
  );


  and

  (
    g1235_p,
    G98_n_spl_011,
    G121_n_spl_11
  );


  or

  (
    g1235_n,
    G98_p_spl_011,
    G121_p_spl_11
  );


  and

  (
    g1236_p,
    g1234_n,
    g1235_n
  );


  or

  (
    g1236_n,
    g1234_p,
    g1235_p
  );


  and

  (
    g1237_p,
    G147_n_spl_1,
    g1236_n
  );


  or

  (
    g1237_n,
    G147_p_spl_1,
    g1236_p
  );


  and

  (
    g1238_p,
    g1233_n,
    g1237_n
  );


  or

  (
    g1238_n,
    g1233_p,
    g1237_p
  );


  and

  (
    g1239_p,
    g1229_n_spl_,
    g1238_p_spl_
  );


  or

  (
    g1239_n,
    g1229_p_spl_,
    g1238_n_spl_
  );


  and

  (
    g1240_p,
    g1229_p_spl_,
    g1238_n_spl_
  );


  or

  (
    g1240_n,
    g1229_n_spl_,
    g1238_p_spl_
  );


  and

  (
    g1241_p,
    g1239_n,
    g1240_n
  );


  or

  (
    g1241_n,
    g1239_p,
    g1240_p
  );


  and

  (
    g1242_p,
    g245_n_spl_1,
    g1241_p_spl_
  );


  or

  (
    g1242_n,
    g245_p_spl_,
    g1241_n_spl_
  );


  and

  (
    g1243_p,
    g245_p_spl_,
    g1241_n_spl_
  );


  or

  (
    g1243_n,
    g245_n_spl_1,
    g1241_p_spl_
  );


  and

  (
    g1244_p,
    g1242_n,
    g1243_n
  );


  or

  (
    g1244_n,
    g1242_p,
    g1243_p
  );


  and

  (
    g1245_p,
    g1226_p_spl_,
    g1244_n_spl_
  );


  or

  (
    g1245_n,
    g1226_n_spl_,
    g1244_p_spl_
  );


  and

  (
    g1246_p,
    g1226_n_spl_,
    g1244_p_spl_
  );


  or

  (
    g1246_n,
    g1226_p_spl_,
    g1244_n_spl_
  );


  and

  (
    g1247_p,
    g1245_n,
    g1246_n
  );


  or

  (
    g1247_n,
    g1245_p,
    g1246_p
  );


  or

  (
    g1248_n,
    g1205_p,
    g1247_n
  );


  or

  (
    g1249_n,
    g1205_n,
    g1247_p
  );


  and

  (
    g1250_p,
    g1248_n,
    g1249_n
  );


  or

  (
    g1251_n,
    G176_n_spl_110,
    g1250_p
  );


  and

  (
    g1252_p,
    g464_n_spl_10,
    g596_n_spl_0
  );


  or

  (
    g1252_n,
    g464_p_spl_10,
    g596_p_spl_1
  );


  and

  (
    g1253_p,
    g464_p_spl_1,
    g596_p_spl_1
  );


  or

  (
    g1253_n,
    g464_n_spl_1,
    g596_n_spl_
  );


  and

  (
    g1254_p,
    g1252_n,
    g1253_n
  );


  or

  (
    g1254_n,
    g1252_p,
    g1253_p
  );


  and

  (
    g1255_p,
    g617_p_spl_0,
    g1254_n_spl_
  );


  or

  (
    g1255_n,
    g617_n_spl_,
    g1254_p_spl_
  );


  and

  (
    g1256_p,
    g617_n_spl_,
    g1254_p_spl_
  );


  or

  (
    g1256_n,
    g617_p_spl_,
    g1254_n_spl_
  );


  and

  (
    g1257_p,
    g1255_n,
    g1256_n
  );


  or

  (
    g1257_n,
    g1255_p,
    g1256_p
  );


  and

  (
    g1258_p,
    g598_p_spl_0,
    g1257_p_spl_
  );


  or

  (
    g1258_n,
    g598_n_spl_0,
    g1257_n_spl_
  );


  and

  (
    g1259_p,
    g598_n_spl_,
    g1257_n_spl_
  );


  or

  (
    g1259_n,
    g598_p_spl_,
    g1257_p_spl_
  );


  and

  (
    g1260_p,
    g1258_n,
    g1259_n
  );


  or

  (
    g1260_n,
    g1258_p,
    g1259_p
  );


  and

  (
    g1261_p,
    G162_n_spl_,
    g562_p
  );


  or

  (
    g1261_n,
    G162_p_spl_,
    g562_n_spl_
  );


  and

  (
    g1262_p,
    G162_p_spl_,
    g461_n_spl_
  );


  or

  (
    g1262_n,
    G162_n_spl_,
    g461_p_spl_
  );


  and

  (
    g1263_p,
    g1261_n,
    g1262_n
  );


  or

  (
    g1263_n,
    g1261_p,
    g1262_p
  );


  and

  (
    g1264_p,
    g1260_p_spl_,
    g1263_p_spl_
  );


  or

  (
    g1264_n,
    g1260_n_spl_,
    g1263_n_spl_
  );


  and

  (
    g1265_p,
    g1260_n_spl_,
    g1263_n_spl_
  );


  or

  (
    g1265_n,
    g1260_p_spl_,
    g1263_p_spl_
  );


  and

  (
    g1266_p,
    g1264_n,
    g1265_n
  );


  or

  (
    g1266_n,
    g1264_p,
    g1265_p
  );


  and

  (
    g1267_p,
    g450_n_spl_1,
    g454_n_spl_1
  );


  or

  (
    g1267_n,
    g450_p_spl_1,
    g454_p_spl_1
  );


  and

  (
    g1268_p,
    g455_n_spl_,
    g1267_n
  );


  or

  (
    g1268_n,
    g455_p_spl_,
    g1267_p
  );


  and

  (
    g1269_p,
    g471_p_spl_1,
    g1268_n_spl_
  );


  or

  (
    g1269_n,
    g471_n_spl_1,
    g1268_p_spl_
  );


  and

  (
    g1270_p,
    g471_n_spl_1,
    g1268_p_spl_
  );


  or

  (
    g1270_n,
    g471_p_spl_1,
    g1268_n_spl_
  );


  and

  (
    g1271_p,
    g1269_n,
    g1270_n
  );


  or

  (
    g1271_n,
    g1269_p,
    g1270_p
  );


  and

  (
    g1272_p,
    g1266_n_spl_,
    g1271_n_spl_
  );


  or

  (
    g1272_n,
    g1266_p_spl_,
    g1271_p_spl_
  );


  and

  (
    g1273_p,
    g1266_p_spl_,
    g1271_p_spl_
  );


  or

  (
    g1273_n,
    g1266_n_spl_,
    g1271_n_spl_
  );


  and

  (
    g1274_p,
    g1272_n,
    g1273_n
  );


  or

  (
    g1274_n,
    g1272_p,
    g1273_p
  );


  and

  (
    g1275_p,
    g444_n_spl_,
    g780_p_spl_0
  );


  or

  (
    g1275_n,
    g444_p_spl_,
    g780_n_spl_0
  );


  and

  (
    g1276_p,
    g442_n_spl_1,
    g1275_n_spl_
  );


  or

  (
    g1276_n,
    g442_p_spl_1,
    g1275_p_spl_
  );


  and

  (
    g1277_p,
    g442_p_spl_1,
    g1275_p_spl_
  );


  or

  (
    g1277_n,
    g442_n_spl_1,
    g1275_n_spl_
  );


  and

  (
    g1278_p,
    g1276_n,
    g1277_n
  );


  or

  (
    g1278_n,
    g1276_p,
    g1277_p
  );


  and

  (
    g1279_p,
    g479_n_spl_01,
    g1278_p_spl_
  );


  or

  (
    g1279_n,
    g479_p_spl_01,
    g1278_n_spl_
  );


  and

  (
    g1280_p,
    g479_p_spl_10,
    g1278_n_spl_
  );


  or

  (
    g1280_n,
    g479_n_spl_10,
    g1278_p_spl_
  );


  and

  (
    g1281_p,
    g1279_n,
    g1280_n
  );


  or

  (
    g1281_n,
    g1279_p,
    g1280_p
  );


  and

  (
    g1282_p,
    g443_n_spl_0,
    g1281_p_spl_
  );


  or

  (
    g1282_n,
    g443_p_spl_0,
    g1281_n_spl_
  );


  and

  (
    g1283_p,
    g443_p_spl_1,
    g1281_n_spl_
  );


  or

  (
    g1283_n,
    g443_n_spl_1,
    g1281_p_spl_
  );


  and

  (
    g1284_p,
    g1282_n_spl_,
    g1283_n
  );


  or

  (
    g1284_n,
    g1282_p_spl_,
    g1283_p
  );


  and

  (
    g1285_p,
    g437_p_spl_01,
    g1284_n_spl_
  );


  or

  (
    g1285_n,
    g437_n_spl_01,
    g1284_p_spl_
  );


  and

  (
    g1286_p,
    g441_p_spl_1,
    g780_n_spl_1
  );


  or

  (
    g1286_n,
    g441_n_spl_1,
    g780_p_spl_1
  );


  and

  (
    g1287_p,
    g441_n_spl_1,
    g780_p_spl_1
  );


  or

  (
    g1287_n,
    g441_p_spl_1,
    g780_n_spl_1
  );


  and

  (
    g1288_p,
    g1286_n,
    g1287_n
  );


  or

  (
    g1288_n,
    g1286_p,
    g1287_p
  );


  and

  (
    g1289_p,
    g479_p_spl_10,
    g1288_n_spl_
  );


  or

  (
    g1289_n,
    g479_n_spl_10,
    g1288_p_spl_
  );


  and

  (
    g1290_p,
    g479_n_spl_1,
    g1288_p_spl_
  );


  or

  (
    g1290_n,
    g479_p_spl_1,
    g1288_n_spl_
  );


  and

  (
    g1291_p,
    g1289_n,
    g1290_n
  );


  or

  (
    g1291_n,
    g1289_p,
    g1290_p
  );


  and

  (
    g1292_p,
    g443_p_spl_1,
    g1291_n
  );


  or

  (
    g1292_n,
    g443_n_spl_1,
    g1291_p
  );


  and

  (
    g1293_p,
    g437_n_spl_1,
    g1292_n
  );


  or

  (
    g1293_n,
    g437_p_spl_1,
    g1292_p
  );


  and

  (
    g1294_p,
    g1282_n_spl_,
    g1293_p
  );


  or

  (
    g1294_n,
    g1282_p_spl_,
    g1293_n
  );


  and

  (
    g1295_p,
    g774_p_spl_1,
    g1294_p
  );


  or

  (
    g1295_n,
    g774_n_spl_1,
    g1294_n
  );


  and

  (
    g1296_p,
    g1285_n,
    g1295_n
  );


  or

  (
    g1296_n,
    g1285_p,
    g1295_p
  );


  and

  (
    g1297_p,
    g437_n_spl_1,
    g774_n_spl_1
  );


  or

  (
    g1297_n,
    g437_p_spl_1,
    g774_p_spl_1
  );


  and

  (
    g1298_p,
    g1284_p_spl_,
    g1297_p
  );


  or

  (
    g1298_n,
    g1284_n_spl_,
    g1297_n
  );


  and

  (
    g1299_p,
    g1296_p,
    g1298_n
  );


  or

  (
    g1299_n,
    g1296_n,
    g1298_p
  );


  and

  (
    g1300_p,
    g581_p_spl_01,
    g1299_p_spl_
  );


  or

  (
    g1300_n,
    g581_n_spl_11,
    g1299_n_spl_
  );


  and

  (
    g1301_p,
    g581_n_spl_11,
    g1299_n_spl_
  );


  or

  (
    g1301_n,
    g581_p_spl_1,
    g1299_p_spl_
  );


  and

  (
    g1302_p,
    g1300_n,
    g1301_n
  );


  or

  (
    g1302_n,
    g1300_p,
    g1301_p
  );


  and

  (
    g1303_p,
    g1274_p,
    g1302_n
  );


  and

  (
    g1304_p,
    g1274_n,
    g1302_p
  );


  or

  (
    g1305_n,
    G176_p_spl_1111,
    g1304_p
  );


  or

  (
    g1306_n,
    g1303_p,
    g1305_n
  );


  and

  (
    g1307_p,
    g1251_n,
    g1306_n
  );


  or

  (
    g1308_n,
    G177_n_spl_111,
    g1307_p
  );


  or

  (
    g1309_n,
    G51_p,
    G177_p_spl_110
  );


  or

  (
    g1310_n,
    G176_n_spl_110,
    g1309_n
  );


  and

  (
    g1311_p,
    g1308_n_spl_,
    g1310_n
  );


  and

  (
    g1312_p,
    G94_p_spl_10,
    G101_p_spl_100
  );


  or

  (
    g1312_n,
    G94_n_spl_10,
    G101_n_spl_100
  );


  and

  (
    g1313_p,
    G94_n_spl_10,
    G100_p_spl_100
  );


  or

  (
    g1313_n,
    G94_p_spl_10,
    G100_n_spl_100
  );


  and

  (
    g1314_p,
    g1312_n,
    g1313_n
  );


  or

  (
    g1314_n,
    g1312_p,
    g1313_p
  );


  and

  (
    g1315_p,
    G140_p_spl_1,
    g1314_n
  );


  or

  (
    g1315_n,
    G140_n_spl_1,
    g1314_p
  );


  and

  (
    g1316_p,
    G94_p_spl_11,
    G102_n_spl_011
  );


  or

  (
    g1316_n,
    G94_n_spl_11,
    G102_p_spl_011
  );


  and

  (
    g1317_p,
    G94_n_spl_11,
    G98_n_spl_100
  );


  or

  (
    g1317_n,
    G94_p_spl_11,
    G98_p_spl_100
  );


  and

  (
    g1318_p,
    g1316_n,
    g1317_n
  );


  or

  (
    g1318_n,
    g1316_p,
    g1317_p
  );


  and

  (
    g1319_p,
    G140_n_spl_1,
    g1318_n
  );


  or

  (
    g1319_n,
    G140_p_spl_1,
    g1318_p
  );


  and

  (
    g1320_p,
    g1315_n,
    g1319_n
  );


  or

  (
    g1320_n,
    g1315_p,
    g1319_p
  );


  and

  (
    g1321_p,
    G92_p_spl_10,
    G101_p_spl_100
  );


  or

  (
    g1321_n,
    G92_n_spl_10,
    G101_n_spl_100
  );


  and

  (
    g1322_p,
    G92_n_spl_10,
    G100_p_spl_100
  );


  or

  (
    g1322_n,
    G92_p_spl_10,
    G100_n_spl_100
  );


  and

  (
    g1323_p,
    g1321_n,
    g1322_n
  );


  or

  (
    g1323_n,
    g1321_p,
    g1322_p
  );


  and

  (
    g1324_p,
    G144_p_spl_1,
    g1323_n
  );


  or

  (
    g1324_n,
    G144_n_spl_1,
    g1323_p
  );


  and

  (
    g1325_p,
    G92_p_spl_11,
    G102_n_spl_100
  );


  or

  (
    g1325_n,
    G92_n_spl_11,
    G102_p_spl_100
  );


  and

  (
    g1326_p,
    G92_n_spl_11,
    G98_n_spl_100
  );


  or

  (
    g1326_n,
    G92_p_spl_11,
    G98_p_spl_100
  );


  and

  (
    g1327_p,
    g1325_n,
    g1326_n
  );


  or

  (
    g1327_n,
    g1325_p,
    g1326_p
  );


  and

  (
    g1328_p,
    G144_n_spl_1,
    g1327_n
  );


  or

  (
    g1328_n,
    G144_p_spl_1,
    g1327_p
  );


  and

  (
    g1329_p,
    g1324_n,
    g1328_n
  );


  or

  (
    g1329_n,
    g1324_p,
    g1328_p
  );


  and

  (
    g1330_p,
    g1320_n_spl_,
    g1329_p_spl_
  );


  or

  (
    g1330_n,
    g1320_p_spl_,
    g1329_n_spl_
  );


  and

  (
    g1331_p,
    g1320_p_spl_,
    g1329_n_spl_
  );


  or

  (
    g1331_n,
    g1320_n_spl_,
    g1329_p_spl_
  );


  and

  (
    g1332_p,
    g1330_n,
    g1331_n
  );


  or

  (
    g1332_n,
    g1330_p,
    g1331_p
  );


  and

  (
    g1333_p,
    G90_p_spl_10,
    G101_p_spl_101
  );


  or

  (
    g1333_n,
    G90_n_spl_10,
    G101_n_spl_101
  );


  and

  (
    g1334_p,
    G90_n_spl_10,
    G100_p_spl_101
  );


  or

  (
    g1334_n,
    G90_p_spl_10,
    G100_n_spl_101
  );


  and

  (
    g1335_p,
    g1333_n,
    g1334_n
  );


  or

  (
    g1335_n,
    g1333_p,
    g1334_p
  );


  and

  (
    g1336_p,
    G143_p_spl_1,
    g1335_n
  );


  or

  (
    g1336_n,
    G143_n_spl_1,
    g1335_p
  );


  and

  (
    g1337_p,
    G90_p_spl_11,
    G102_n_spl_100
  );


  or

  (
    g1337_n,
    G90_n_spl_11,
    G102_p_spl_100
  );


  and

  (
    g1338_p,
    G90_n_spl_11,
    G98_n_spl_101
  );


  or

  (
    g1338_n,
    G90_p_spl_11,
    G98_p_spl_101
  );


  and

  (
    g1339_p,
    g1337_n,
    g1338_n
  );


  or

  (
    g1339_n,
    g1337_p,
    g1338_p
  );


  and

  (
    g1340_p,
    G143_n_spl_1,
    g1339_n
  );


  or

  (
    g1340_n,
    G143_p_spl_1,
    g1339_p
  );


  and

  (
    g1341_p,
    g1336_n,
    g1340_n
  );


  or

  (
    g1341_n,
    g1336_p,
    g1340_p
  );


  and

  (
    g1342_p,
    g317_n_spl_1,
    g1341_n_spl_
  );


  or

  (
    g1342_n,
    g317_p_spl_,
    g1341_p_spl_
  );


  and

  (
    g1343_p,
    g317_p_spl_,
    g1341_p_spl_
  );


  or

  (
    g1343_n,
    g317_n_spl_1,
    g1341_n_spl_
  );


  and

  (
    g1344_p,
    g1342_n,
    g1343_n
  );


  or

  (
    g1344_n,
    g1342_p,
    g1343_p
  );


  and

  (
    g1345_p,
    g1332_n_spl_,
    g1344_p_spl_
  );


  or

  (
    g1345_n,
    g1332_p_spl_,
    g1344_n_spl_
  );


  and

  (
    g1346_p,
    g1332_p_spl_,
    g1344_n_spl_
  );


  or

  (
    g1346_n,
    g1332_n_spl_,
    g1344_p_spl_
  );


  and

  (
    g1347_p,
    g1345_n,
    g1346_n
  );


  or

  (
    g1347_n,
    g1345_p,
    g1346_p
  );


  and

  (
    g1348_p,
    G101_p_spl_101,
    G107_p_spl_10
  );


  or

  (
    g1348_n,
    G101_n_spl_101,
    G107_n_spl_10
  );


  and

  (
    g1349_p,
    G100_p_spl_101,
    G107_n_spl_10
  );


  or

  (
    g1349_n,
    G100_n_spl_101,
    G107_p_spl_10
  );


  and

  (
    g1350_p,
    g1348_n,
    g1349_n
  );


  or

  (
    g1350_n,
    g1348_p,
    g1349_p
  );


  and

  (
    g1351_p,
    G139_p_spl_1,
    g1350_n
  );


  or

  (
    g1351_n,
    G139_n_spl_1,
    g1350_p
  );


  and

  (
    g1352_p,
    G102_n_spl_101,
    G107_p_spl_11
  );


  or

  (
    g1352_n,
    G102_p_spl_101,
    G107_n_spl_11
  );


  and

  (
    g1353_p,
    G98_n_spl_101,
    G107_n_spl_11
  );


  or

  (
    g1353_n,
    G98_p_spl_101,
    G107_p_spl_11
  );


  and

  (
    g1354_p,
    g1352_n,
    g1353_n
  );


  or

  (
    g1354_n,
    g1352_p,
    g1353_p
  );


  and

  (
    g1355_p,
    G139_n_spl_1,
    g1354_n
  );


  or

  (
    g1355_n,
    G139_p_spl_1,
    g1354_p
  );


  and

  (
    g1356_p,
    g1351_n,
    g1355_n
  );


  or

  (
    g1356_n,
    g1351_p,
    g1355_p
  );


  and

  (
    g1357_p,
    G101_p_spl_110,
    G105_p_spl_10
  );


  or

  (
    g1357_n,
    G101_n_spl_110,
    G105_n_spl_10
  );


  and

  (
    g1358_p,
    G100_p_spl_110,
    G105_n_spl_10
  );


  or

  (
    g1358_n,
    G100_n_spl_110,
    G105_p_spl_10
  );


  and

  (
    g1359_p,
    g1357_n,
    g1358_n
  );


  or

  (
    g1359_n,
    g1357_p,
    g1358_p
  );


  and

  (
    g1360_p,
    G138_p_spl_1,
    g1359_n
  );


  or

  (
    g1360_n,
    G138_n_spl_1,
    g1359_p
  );


  and

  (
    g1361_p,
    G102_n_spl_101,
    G105_p_spl_11
  );


  or

  (
    g1361_n,
    G102_p_spl_101,
    G105_n_spl_11
  );


  and

  (
    g1362_p,
    G98_n_spl_110,
    G105_n_spl_11
  );


  or

  (
    g1362_n,
    G98_p_spl_110,
    G105_p_spl_11
  );


  and

  (
    g1363_p,
    g1361_n,
    g1362_n
  );


  or

  (
    g1363_n,
    g1361_p,
    g1362_p
  );


  and

  (
    g1364_p,
    G138_n_spl_1,
    g1363_n
  );


  or

  (
    g1364_n,
    G138_p_spl_1,
    g1363_p
  );


  and

  (
    g1365_p,
    g1360_n,
    g1364_n
  );


  or

  (
    g1365_n,
    g1360_p,
    g1364_p
  );


  and

  (
    g1366_p,
    g1356_n_spl_,
    g1365_p_spl_
  );


  or

  (
    g1366_n,
    g1356_p_spl_,
    g1365_n_spl_
  );


  and

  (
    g1367_p,
    g1356_p_spl_,
    g1365_n_spl_
  );


  or

  (
    g1367_n,
    g1356_n_spl_,
    g1365_p_spl_
  );


  and

  (
    g1368_p,
    g1366_n,
    g1367_n
  );


  or

  (
    g1368_n,
    g1366_p,
    g1367_p
  );


  and

  (
    g1369_p,
    G101_p_spl_110,
    G103_p_spl_10
  );


  or

  (
    g1369_n,
    G101_n_spl_110,
    G103_n_spl_10
  );


  and

  (
    g1370_p,
    G100_p_spl_110,
    G103_n_spl_10
  );


  or

  (
    g1370_n,
    G100_n_spl_110,
    G103_p_spl_10
  );


  and

  (
    g1371_p,
    g1369_n,
    g1370_n
  );


  or

  (
    g1371_n,
    g1369_p,
    g1370_p
  );


  and

  (
    g1372_p,
    G137_p_spl_1,
    g1371_n
  );


  or

  (
    g1372_n,
    G137_n_spl_1,
    g1371_p
  );


  and

  (
    g1373_p,
    G102_n_spl_110,
    G103_p_spl_11
  );


  or

  (
    g1373_n,
    G102_p_spl_110,
    G103_n_spl_11
  );


  and

  (
    g1374_p,
    G98_n_spl_110,
    G103_n_spl_11
  );


  or

  (
    g1374_n,
    G98_p_spl_110,
    G103_p_spl_11
  );


  and

  (
    g1375_p,
    g1373_n,
    g1374_n
  );


  or

  (
    g1375_n,
    g1373_p,
    g1374_p
  );


  and

  (
    g1376_p,
    G137_n_spl_1,
    g1375_n
  );


  or

  (
    g1376_n,
    G137_p_spl_1,
    g1375_p
  );


  and

  (
    g1377_p,
    g1372_n,
    g1376_n
  );


  or

  (
    g1377_n,
    g1372_p,
    g1376_p
  );


  and

  (
    g1378_p,
    G96_p_spl_10,
    G101_p_spl_111
  );


  or

  (
    g1378_n,
    G96_n_spl_10,
    G101_n_spl_111
  );


  and

  (
    g1379_p,
    G96_n_spl_10,
    G100_p_spl_111
  );


  or

  (
    g1379_n,
    G96_p_spl_10,
    G100_n_spl_111
  );


  and

  (
    g1380_p,
    g1378_n,
    g1379_n
  );


  or

  (
    g1380_n,
    g1378_p,
    g1379_p
  );


  and

  (
    g1381_p,
    G141_p_spl_1,
    g1380_n
  );


  or

  (
    g1381_n,
    G141_n_spl_1,
    g1380_p
  );


  and

  (
    g1382_p,
    G96_p_spl_11,
    G102_n_spl_110
  );


  or

  (
    g1382_n,
    G96_n_spl_11,
    G102_p_spl_110
  );


  and

  (
    g1383_p,
    G96_n_spl_11,
    G98_n_spl_111
  );


  or

  (
    g1383_n,
    G96_p_spl_11,
    G98_p_spl_111
  );


  and

  (
    g1384_p,
    g1382_n,
    g1383_n
  );


  or

  (
    g1384_n,
    g1382_p,
    g1383_p
  );


  and

  (
    g1385_p,
    G141_n_spl_1,
    g1384_n
  );


  or

  (
    g1385_n,
    G141_p_spl_1,
    g1384_p
  );


  and

  (
    g1386_p,
    g1381_n,
    g1385_n
  );


  or

  (
    g1386_n,
    g1381_p,
    g1385_p
  );


  and

  (
    g1387_p,
    g1377_n_spl_,
    g1386_p_spl_
  );


  or

  (
    g1387_n,
    g1377_p_spl_,
    g1386_n_spl_
  );


  and

  (
    g1388_p,
    g1377_p_spl_,
    g1386_n_spl_
  );


  or

  (
    g1388_n,
    g1377_n_spl_,
    g1386_p_spl_
  );


  and

  (
    g1389_p,
    g1387_n,
    g1388_n
  );


  or

  (
    g1389_n,
    g1387_p,
    g1388_p
  );


  and

  (
    g1390_p,
    G101_p_spl_111,
    G109_p_spl_10
  );


  or

  (
    g1390_n,
    G101_n_spl_111,
    G109_n_spl_10
  );


  and

  (
    g1391_p,
    G100_p_spl_111,
    G109_n_spl_10
  );


  or

  (
    g1391_n,
    G100_n_spl_111,
    G109_p_spl_10
  );


  and

  (
    g1392_p,
    g1390_n,
    g1391_n
  );


  or

  (
    g1392_n,
    g1390_p,
    g1391_p
  );


  and

  (
    g1393_p,
    G135_p_spl_1,
    g1392_n
  );


  or

  (
    g1393_n,
    G135_n_spl_1,
    g1392_p
  );


  and

  (
    g1394_p,
    G102_n_spl_11,
    G109_p_spl_11
  );


  or

  (
    g1394_n,
    G102_p_spl_11,
    G109_n_spl_11
  );


  and

  (
    g1395_p,
    G98_n_spl_111,
    G109_n_spl_11
  );


  or

  (
    g1395_n,
    G98_p_spl_111,
    G109_p_spl_11
  );


  and

  (
    g1396_p,
    g1394_n,
    g1395_n
  );


  or

  (
    g1396_n,
    g1394_p,
    g1395_p
  );


  and

  (
    g1397_p,
    G135_n_spl_1,
    g1396_n
  );


  or

  (
    g1397_n,
    G135_p_spl_1,
    g1396_p
  );


  and

  (
    g1398_p,
    g1393_n,
    g1397_n
  );


  or

  (
    g1398_n,
    g1393_p,
    g1397_p
  );


  and

  (
    g1399_p,
    g1389_p_spl_,
    g1398_n_spl_
  );


  or

  (
    g1399_n,
    g1389_n_spl_,
    g1398_p_spl_
  );


  and

  (
    g1400_p,
    g1389_n_spl_,
    g1398_p_spl_
  );


  or

  (
    g1400_n,
    g1389_p_spl_,
    g1398_n_spl_
  );


  and

  (
    g1401_p,
    g1399_n,
    g1400_n
  );


  or

  (
    g1401_n,
    g1399_p,
    g1400_p
  );


  and

  (
    g1402_p,
    g1368_p_spl_,
    g1401_n_spl_
  );


  or

  (
    g1402_n,
    g1368_n_spl_,
    g1401_p_spl_
  );


  and

  (
    g1403_p,
    g1368_n_spl_,
    g1401_p_spl_
  );


  or

  (
    g1403_n,
    g1368_p_spl_,
    g1401_n_spl_
  );


  and

  (
    g1404_p,
    g1402_n,
    g1403_n
  );


  or

  (
    g1404_n,
    g1402_p,
    g1403_p
  );


  or

  (
    g1405_n,
    g1347_p,
    g1404_n
  );


  or

  (
    g1406_n,
    g1347_n,
    g1404_p
  );


  and

  (
    g1407_p,
    g1405_n,
    g1406_n
  );


  or

  (
    g1408_n,
    G176_n_spl_111,
    g1407_p
  );


  and

  (
    g1409_p,
    g389_n_spl_,
    g546_p_spl_1
  );


  or

  (
    g1409_n,
    g389_p_spl_,
    g546_n_spl_0
  );


  and

  (
    g1410_p,
    g374_p_spl_1,
    g544_n_spl_1
  );


  or

  (
    g1410_n,
    g374_n_spl_1,
    g544_p_spl_1
  );


  and

  (
    g1411_p,
    g374_n_spl_1,
    g380_p_spl_
  );


  or

  (
    g1411_n,
    g374_p_spl_1,
    g380_n_spl_
  );


  and

  (
    g1412_p,
    g1410_n,
    g1411_n
  );


  or

  (
    g1412_n,
    g1410_p,
    g1411_p
  );


  and

  (
    g1413_p,
    g1409_n_spl_,
    g1412_n_spl_
  );


  or

  (
    g1413_n,
    g1409_p_spl_,
    g1412_p_spl_
  );


  and

  (
    g1414_p,
    g1409_p_spl_,
    g1412_p_spl_
  );


  or

  (
    g1414_n,
    g1409_n_spl_,
    g1412_n_spl_
  );


  and

  (
    g1415_p,
    g1413_n,
    g1414_n
  );


  or

  (
    g1415_n,
    g1413_p,
    g1414_p
  );


  and

  (
    g1416_p,
    g375_n_spl_0,
    g1415_p_spl_
  );


  or

  (
    g1416_n,
    g375_p_spl_0,
    g1415_n_spl_
  );


  and

  (
    g1417_p,
    g544_p_spl_1,
    g546_p_spl_1
  );


  or

  (
    g1417_n,
    g544_n_spl_1,
    g546_n_spl_
  );


  and

  (
    g1418_p,
    g545_n_spl_,
    g1417_n
  );


  or

  (
    g1418_n,
    g545_p_spl_,
    g1417_p
  );


  and

  (
    g1419_p,
    g375_p_spl_1,
    g1418_n
  );


  or

  (
    g1419_n,
    g375_n_spl_1,
    g1418_p
  );


  and

  (
    g1420_p,
    g1416_n_spl_,
    g1419_n
  );


  or

  (
    g1420_n,
    g1416_p_spl_,
    g1419_p
  );


  and

  (
    g1421_p,
    g381_n_spl_01,
    g1420_p_spl_
  );


  or

  (
    g1421_n,
    g381_p_spl_01,
    g1420_n_spl_
  );


  and

  (
    g1422_p,
    g381_p_spl_10,
    g1420_n_spl_
  );


  or

  (
    g1422_n,
    g381_n_spl_10,
    g1420_p_spl_
  );


  and

  (
    g1423_p,
    g1421_n,
    g1422_n
  );


  or

  (
    g1423_n,
    g1421_p,
    g1422_p
  );


  and

  (
    g1424_p,
    g395_n_spl_01,
    g1423_p_spl_
  );


  or

  (
    g1424_n,
    g395_p_spl_00,
    g1423_n_spl_
  );


  and

  (
    g1425_p,
    g395_p_spl_0,
    g1423_n_spl_
  );


  or

  (
    g1425_n,
    g395_n_spl_10,
    g1423_p_spl_
  );


  and

  (
    g1426_p,
    g1424_n,
    g1425_n
  );


  or

  (
    g1426_n,
    g1424_p,
    g1425_p
  );


  and

  (
    g1427_p,
    g388_n_spl_01,
    g1426_p_spl_
  );


  or

  (
    g1427_n,
    g388_p_spl_01,
    g1426_n_spl_
  );


  and

  (
    g1428_p,
    g388_p_spl_01,
    g1426_n_spl_
  );


  or

  (
    g1428_n,
    g388_n_spl_01,
    g1426_p_spl_
  );


  and

  (
    g1429_p,
    g1427_n,
    g1428_n
  );


  or

  (
    g1429_n,
    g1427_p,
    g1428_p
  );


  and

  (
    g1430_p,
    g541_p_spl_0,
    g1429_n
  );


  or

  (
    g1430_n,
    g541_n_spl_0,
    g1429_p
  );


  and

  (
    g1431_p,
    g375_p_spl_1,
    g1415_n_spl_
  );


  or

  (
    g1431_n,
    g375_n_spl_1,
    g1415_p_spl_
  );


  and

  (
    g1432_p,
    g1416_n_spl_,
    g1431_n
  );


  or

  (
    g1432_n,
    g1416_p_spl_,
    g1431_p
  );


  and

  (
    g1433_p,
    g381_n_spl_10,
    g1432_p_spl_
  );


  or

  (
    g1433_n,
    g381_p_spl_10,
    g1432_n_spl_
  );


  and

  (
    g1434_p,
    g381_p_spl_1,
    g1432_n_spl_
  );


  or

  (
    g1434_n,
    g381_n_spl_1,
    g1432_p_spl_
  );


  and

  (
    g1435_p,
    g1433_n,
    g1434_n
  );


  or

  (
    g1435_n,
    g1433_p,
    g1434_p
  );


  and

  (
    g1436_p,
    g395_n_spl_10,
    g1435_p_spl_
  );


  or

  (
    g1436_n,
    g395_p_spl_1,
    g1435_n_spl_
  );


  and

  (
    g1437_p,
    g395_p_spl_1,
    g1435_n_spl_
  );


  or

  (
    g1437_n,
    g395_n_spl_1,
    g1435_p_spl_
  );


  and

  (
    g1438_p,
    g1436_n,
    g1437_n
  );


  or

  (
    g1438_n,
    g1436_p,
    g1437_p
  );


  and

  (
    g1439_p,
    g388_n_spl_1,
    g1438_p_spl_
  );


  or

  (
    g1439_n,
    g388_p_spl_1,
    g1438_n_spl_
  );


  and

  (
    g1440_p,
    g388_p_spl_1,
    g1438_n_spl_
  );


  or

  (
    g1440_n,
    g388_n_spl_1,
    g1438_p_spl_
  );


  and

  (
    g1441_p,
    g1439_n,
    g1440_n
  );


  or

  (
    g1441_n,
    g1439_p,
    g1440_p
  );


  and

  (
    g1442_p,
    g541_n_spl_1,
    g1441_n_spl_
  );


  or

  (
    g1442_n,
    g541_p_spl_1,
    g1441_p_spl_
  );


  and

  (
    g1443_p,
    g1430_n_spl_,
    g1442_n
  );


  or

  (
    g1443_n,
    g1430_p_spl_,
    g1442_p
  );


  and

  (
    g1444_p,
    G157_n_spl_0,
    g1443_n
  );


  or

  (
    g1444_n,
    G157_p_spl_0,
    g1443_p
  );


  and

  (
    g1445_p,
    g430_n_spl_1,
    g541_p_spl_1
  );


  or

  (
    g1445_n,
    g430_p_spl_0,
    g541_n_spl_1
  );


  and

  (
    g1446_p,
    g1441_n_spl_,
    g1445_n
  );


  or

  (
    g1446_n,
    g1441_p_spl_,
    g1445_p
  );


  and

  (
    g1447_p,
    g430_n_spl_1,
    g1430_p_spl_
  );


  or

  (
    g1447_n,
    g430_p_spl_,
    g1430_n_spl_
  );


  and

  (
    g1448_p,
    g1446_n,
    g1447_n
  );


  or

  (
    g1448_n,
    g1446_p,
    g1447_p
  );


  and

  (
    g1449_p,
    G157_p_spl_0,
    g1448_n
  );


  or

  (
    g1449_n,
    G157_n_spl_0,
    g1448_p
  );


  and

  (
    g1450_p,
    g1444_n,
    g1449_n
  );


  or

  (
    g1450_n,
    g1444_p,
    g1449_p
  );


  and

  (
    g1451_p,
    g400_p_spl_1,
    g537_n_spl_0
  );


  or

  (
    g1451_n,
    g400_n_spl_1,
    g537_p_spl_0
  );


  and

  (
    g1452_p,
    g400_n_spl_1,
    g537_p_spl_1
  );


  or

  (
    g1452_n,
    g400_p_spl_1,
    g537_n_spl_1
  );


  and

  (
    g1453_p,
    g1451_n,
    g1452_n
  );


  or

  (
    g1453_n,
    g1451_p,
    g1452_p
  );


  and

  (
    g1454_p,
    g535_p_spl_0,
    g1453_n_spl_
  );


  or

  (
    g1454_n,
    g535_n_spl_0,
    g1453_p_spl_
  );


  and

  (
    g1455_p,
    g535_n_spl_1,
    g1453_p_spl_
  );


  or

  (
    g1455_n,
    g535_p_spl_1,
    g1453_n_spl_
  );


  and

  (
    g1456_p,
    g1454_n,
    g1455_n
  );


  or

  (
    g1456_n,
    g1454_p,
    g1455_p
  );


  and

  (
    g1457_p,
    g402_n_spl_,
    g408_n_spl_1
  );


  or

  (
    g1457_n,
    g402_p_spl_1,
    g408_p_spl_1
  );


  and

  (
    g1458_p,
    g409_n_spl_0,
    g1457_n
  );


  or

  (
    g1458_n,
    g409_p_spl_0,
    g1457_p
  );


  and

  (
    g1459_p,
    g539_n_spl_0,
    g1458_n_spl_0
  );


  or

  (
    g1459_n,
    g539_p_spl_0,
    g1458_p_spl_0
  );


  and

  (
    g1460_p,
    g539_p_spl_1,
    g1458_p_spl_0
  );


  or

  (
    g1460_n,
    g539_n_spl_1,
    g1458_n_spl_0
  );


  and

  (
    g1461_p,
    g1459_n,
    g1460_n
  );


  or

  (
    g1461_n,
    g1459_p,
    g1460_p
  );


  and

  (
    g1462_p,
    g1456_n_spl_,
    g1461_p_spl_
  );


  or

  (
    g1462_n,
    g1456_p_spl_,
    g1461_n_spl_
  );


  and

  (
    g1463_p,
    g1456_p_spl_,
    g1461_n_spl_
  );


  or

  (
    g1463_n,
    g1456_n_spl_,
    g1461_p_spl_
  );


  and

  (
    g1464_p,
    g1462_n,
    g1463_n
  );


  or

  (
    g1464_n,
    g1462_p,
    g1463_p
  );


  and

  (
    g1465_p,
    g429_n_spl_01,
    g1464_n_spl_
  );


  or

  (
    g1465_n,
    g429_p_spl_01,
    g1464_p_spl_
  );


  and

  (
    g1466_p,
    g429_p_spl_10,
    g1464_p_spl_
  );


  or

  (
    g1466_n,
    g429_n_spl_10,
    g1464_n_spl_
  );


  and

  (
    g1467_p,
    g1465_n,
    g1466_n
  );


  or

  (
    g1467_n,
    g1465_p,
    g1466_p
  );


  and

  (
    g1468_p,
    G157_n_spl_1,
    g1467_p
  );


  or

  (
    g1468_n,
    G157_p_spl_1,
    g1467_n
  );


  and

  (
    g1469_p,
    g423_n_spl_,
    g539_p_spl_1
  );


  or

  (
    g1469_n,
    g423_p_spl_,
    g539_n_spl_1
  );


  and

  (
    g1470_p,
    g409_n_spl_,
    g535_p_spl_1
  );


  or

  (
    g1470_n,
    g409_p_spl_,
    g535_n_spl_1
  );


  and

  (
    g1471_p,
    g416_n_spl_,
    g537_p_spl_1
  );


  or

  (
    g1471_n,
    g416_p_spl_,
    g537_n_spl_1
  );


  and

  (
    g1472_p,
    g401_n_spl_0,
    g1471_n_spl_
  );


  or

  (
    g1472_n,
    g401_p_spl_0,
    g1471_p_spl_
  );


  and

  (
    g1473_p,
    g401_p_spl_,
    g1471_p_spl_
  );


  or

  (
    g1473_n,
    g401_n_spl_,
    g1471_n_spl_
  );


  and

  (
    g1474_p,
    g1472_n,
    g1473_n
  );


  or

  (
    g1474_n,
    g1472_p,
    g1473_p
  );


  and

  (
    g1475_p,
    g1470_n_spl_,
    g1474_p_spl_
  );


  or

  (
    g1475_n,
    g1470_p_spl_,
    g1474_n_spl_
  );


  and

  (
    g1476_p,
    g1470_p_spl_,
    g1474_n_spl_
  );


  or

  (
    g1476_n,
    g1470_n_spl_,
    g1474_p_spl_
  );


  and

  (
    g1477_p,
    g1475_n,
    g1476_n
  );


  or

  (
    g1477_n,
    g1475_p,
    g1476_p
  );


  and

  (
    g1478_p,
    g1469_n_spl_,
    g1477_p_spl_
  );


  or

  (
    g1478_n,
    g1469_p_spl_,
    g1477_n_spl_
  );


  and

  (
    g1479_p,
    g1469_p_spl_,
    g1477_n_spl_
  );


  or

  (
    g1479_n,
    g1469_n_spl_,
    g1477_p_spl_
  );


  and

  (
    g1480_p,
    g1478_n,
    g1479_n
  );


  or

  (
    g1480_n,
    g1478_p,
    g1479_p
  );


  and

  (
    g1481_p,
    g429_n_spl_10,
    g1458_n_spl_1
  );


  or

  (
    g1481_n,
    g429_p_spl_10,
    g1458_p_spl_1
  );


  and

  (
    g1482_p,
    g429_p_spl_1,
    g1458_p_spl_1
  );


  or

  (
    g1482_n,
    g429_n_spl_1,
    g1458_n_spl_1
  );


  and

  (
    g1483_p,
    g1481_n,
    g1482_n
  );


  or

  (
    g1483_n,
    g1481_p,
    g1482_p
  );


  and

  (
    g1484_p,
    g1480_n_spl_,
    g1483_p_spl_
  );


  or

  (
    g1484_n,
    g1480_p_spl_,
    g1483_n_spl_
  );


  and

  (
    g1485_p,
    g1480_p_spl_,
    g1483_n_spl_
  );


  or

  (
    g1485_n,
    g1480_n_spl_,
    g1483_p_spl_
  );


  and

  (
    g1486_p,
    g1484_n,
    g1485_n
  );


  or

  (
    g1486_n,
    g1484_p,
    g1485_p
  );


  and

  (
    g1487_p,
    G157_p_spl_1,
    g1486_n
  );


  or

  (
    g1487_n,
    G157_n_spl_1,
    g1486_p
  );


  and

  (
    g1488_p,
    g1468_n,
    g1487_n
  );


  or

  (
    g1488_n,
    g1468_p,
    g1487_p
  );


  and

  (
    g1489_p,
    g415_p_spl_1,
    g1488_p_spl_
  );


  or

  (
    g1489_n,
    g415_n_spl_1,
    g1488_n_spl_
  );


  and

  (
    g1490_p,
    g415_n_spl_1,
    g1488_n_spl_
  );


  or

  (
    g1490_n,
    g415_p_spl_1,
    g1488_p_spl_
  );


  and

  (
    g1491_p,
    g1489_n,
    g1490_n
  );


  or

  (
    g1491_n,
    g1489_p,
    g1490_p
  );


  and

  (
    g1492_p,
    g422_p_spl_1,
    g1491_n_spl_
  );


  or

  (
    g1492_n,
    g422_n_spl_1,
    g1491_p_spl_
  );


  and

  (
    g1493_p,
    g422_n_spl_1,
    g1491_p_spl_
  );


  or

  (
    g1493_n,
    g422_p_spl_1,
    g1491_n_spl_
  );


  and

  (
    g1494_p,
    g1492_n,
    g1493_n
  );


  or

  (
    g1494_n,
    g1492_p,
    g1493_p
  );


  and

  (
    g1495_p,
    g1450_n,
    g1494_n
  );


  and

  (
    g1496_p,
    g1450_p,
    g1494_p
  );


  or

  (
    g1497_n,
    G176_p_spl_1111,
    g1496_p
  );


  or

  (
    g1498_n,
    g1495_p,
    g1497_n
  );


  and

  (
    g1499_p,
    g1408_n,
    g1498_n
  );


  or

  (
    g1500_n,
    G177_n_spl_111,
    g1499_p
  );


  or

  (
    g1501_n,
    G49_p,
    G177_p_spl_110
  );


  or

  (
    g1502_n,
    G176_n_spl_111,
    g1501_n
  );


  and

  (
    g1503_p,
    g1500_n_spl_,
    g1502_n
  );


  or

  (
    g1504_n,
    G23_n_spl_,
    G173_p_spl_111
  );


  or

  (
    g1505_n,
    G4_n_spl_,
    G173_n_spl_111
  );


  and

  (
    g1506_p,
    g1504_n,
    g1505_n
  );


  or

  (
    g1507_n,
    G172_p_spl_11,
    g1506_p
  );


  or

  (
    g1508_n,
    G38_n,
    G177_p_spl_111
  );


  and

  (
    g1509_p,
    g1500_n_spl_,
    g1508_n
  );


  and

  (
    g1510_p,
    G173_n_spl_111,
    g1509_p_spl_0
  );


  or

  (
    g1511_n,
    G37_n,
    G177_p_spl_111
  );


  and

  (
    g1512_p,
    g1308_n_spl_,
    g1511_n
  );


  and

  (
    g1513_p,
    G173_p_spl_111,
    g1512_p_spl_0
  );


  or

  (
    g1514_n,
    G172_n_spl_11,
    g1513_p
  );


  or

  (
    g1515_n,
    g1510_p,
    g1514_n
  );


  and

  (
    g1516_p,
    g1507_n,
    g1515_n
  );


  or

  (
    g1517_n,
    G23_n_spl_,
    G174_p_spl_111
  );


  or

  (
    g1518_n,
    G4_n_spl_,
    G174_n_spl_111
  );


  and

  (
    g1519_p,
    g1517_n,
    g1518_n
  );


  or

  (
    g1520_n,
    G175_p_spl_11,
    g1519_p
  );


  and

  (
    g1521_p,
    G174_n_spl_111,
    g1509_p_spl_0
  );


  and

  (
    g1522_p,
    G174_p_spl_111,
    g1512_p_spl_0
  );


  or

  (
    g1523_n,
    G175_n_spl_11,
    g1522_p
  );


  or

  (
    g1524_n,
    g1521_p,
    g1523_n
  );


  and

  (
    g1525_p,
    g1520_n,
    g1524_n
  );


  or

  (
    g1526_n,
    G79_n_spl_,
    G158_p_spl_111
  );


  or

  (
    g1527_n,
    G78_n_spl_,
    G158_n_spl_111
  );


  and

  (
    g1528_p,
    g1526_n,
    g1527_n
  );


  or

  (
    g1529_n,
    G159_p_spl_11,
    g1528_p
  );


  or

  (
    g1530_n,
    G158_n_spl_111,
    g1512_p_spl_1
  );


  or

  (
    g1531_n,
    G158_p_spl_111,
    g1509_p_spl_1
  );


  and

  (
    g1532_p,
    g1530_n,
    g1531_n
  );


  or

  (
    g1533_n,
    G159_n_spl_11,
    g1532_p
  );


  and

  (
    g1534_p,
    g1529_n,
    g1533_n
  );


  or

  (
    g1535_n,
    G64_n_spl_,
    g1534_p
  );


  or

  (
    g1536_n,
    G79_n_spl_,
    G160_p_spl_111
  );


  or

  (
    g1537_n,
    G78_n_spl_,
    G160_n_spl_111
  );


  and

  (
    g1538_p,
    g1536_n,
    g1537_n
  );


  or

  (
    g1539_n,
    G161_p_spl_11,
    g1538_p
  );


  or

  (
    g1540_n,
    G160_n_spl_111,
    g1512_p_spl_1
  );


  or

  (
    g1541_n,
    G160_p_spl_111,
    g1509_p_spl_1
  );


  and

  (
    g1542_p,
    g1540_n,
    g1541_n
  );


  or

  (
    g1543_n,
    G161_n_spl_11,
    g1542_p
  );


  and

  (
    g1544_p,
    g1539_n,
    g1543_n
  );


  or

  (
    g1545_n,
    G64_n_spl_,
    g1544_p
  );


  buf

  (
    G5193,
    G66_n
  );


  buf

  (
    G5194,
    G113_n_spl_1
  );


  buf

  (
    G5195,
    G165_n_spl_
  );


  buf

  (
    G5196,
    G151_n_spl_0
  );


  buf

  (
    G5197,
    G127_n_spl_
  );


  buf

  (
    G5198,
    G131_n_spl_
  );


  not

  (
    G5199,
    g179_n_spl_
  );


  buf

  (
    G5200,
    G152_n
  );


  buf

  (
    G5201,
    G151_n_spl_0
  );


  buf

  (
    G5202,
    G151_n_spl_
  );


  buf

  (
    G5203,
    G125_n_spl_
  );


  buf

  (
    G5204,
    G129_n_spl_
  );


  buf

  (
    G5205,
    g180_p
  );


  buf

  (
    G5206,
    G99_n_spl_
  );


  buf

  (
    G5207,
    G153_n_spl_
  );


  buf

  (
    G5208,
    G156_n_spl_
  );


  buf

  (
    G5209,
    G155_n_spl_
  );


  buf

  (
    G5210,
    g181_p
  );


  buf

  (
    G5211,
    g182_p
  );


  buf

  (
    G5212,
    g183_n
  );


  buf

  (
    G5213,
    g184_n_spl_
  );


  buf

  (
    G5214,
    G64_p_spl_111
  );


  buf

  (
    G5215,
    G66_p_spl_1
  );


  buf

  (
    G5216,
    G1_p_spl_
  );


  buf

  (
    G5217,
    G152_p_spl_
  );


  buf

  (
    G5218,
    G114_p_spl_
  );


  buf

  (
    G5219,
    G152_p_spl_
  );


  buf

  (
    G5220,
    g186_n
  );


  buf

  (
    G5221,
    g185_n_spl_11
  );


  buf

  (
    G5222,
    G1_n_spl_0
  );


  buf

  (
    G5223,
    G1_n_spl_0
  );


  buf

  (
    G5224,
    G1_n_spl_1
  );


  buf

  (
    G5225,
    G1_n_spl_1
  );


  buf

  (
    G5226,
    G114_n_spl_0
  );


  buf

  (
    G5227,
    G114_n_spl_
  );


  buf

  (
    G5228,
    g190_n
  );


  buf

  (
    G5229,
    g194_n_spl_
  );


  buf

  (
    G5230,
    g194_n_spl_
  );


  buf

  (
    G5231,
    g195_n
  );


  buf

  (
    G5232,
    g200_p
  );


  buf

  (
    G5233,
    g205_p
  );


  buf

  (
    G5234,
    g210_p
  );


  buf

  (
    G5235,
    g215_p
  );


  not

  (
    G5236,
    g280_n
  );


  not

  (
    G5237,
    g369_n
  );


  not

  (
    G5238,
    g431_n_spl_
  );


  buf

  (
    G5239,
    g482_p_spl_
  );


  buf

  (
    G5240,
    g482_p_spl_
  );


  not

  (
    G5241,
    g431_n_spl_
  );


  not

  (
    G5242,
    g506_n_spl_
  );


  not

  (
    G5243,
    g533_n_spl_
  );


  not

  (
    G5244,
    g549_p_spl_
  );


  buf

  (
    G5245,
    g550_n_spl_
  );


  not

  (
    G5246,
    g549_p_spl_
  );


  buf

  (
    G5247,
    g550_n_spl_
  );


  not

  (
    G5248,
    g560_p_spl_1
  );


  not

  (
    G5249,
    g569_p_spl_1
  );


  not

  (
    G5250,
    g579_p_spl_1
  );


  buf

  (
    G5251,
    g581_p_spl_1
  );


  buf

  (
    G5252,
    g590_n
  );


  not

  (
    G5253,
    g605_n_spl_1
  );


  not

  (
    G5254,
    g614_n_spl_1
  );


  not

  (
    G5255,
    g624_n_spl_1
  );


  buf

  (
    G5256,
    g633_n
  );


  not

  (
    G5257,
    g647_n_spl_1
  );


  not

  (
    G5258,
    g656_n_spl_1
  );


  not

  (
    G5259,
    g669_n_spl_1
  );


  not

  (
    G5260,
    g678_n_spl_1
  );


  not

  (
    G5261,
    g705_n_spl_
  );


  not

  (
    G5262,
    g735_n_spl_
  );


  not

  (
    G5263,
    g764_n
  );


  not

  (
    G5264,
    g794_n
  );


  buf

  (
    G5265,
    g804_p
  );


  buf

  (
    G5266,
    g814_p
  );


  buf

  (
    G5267,
    g823_n
  );


  buf

  (
    G5268,
    g832_n
  );


  buf

  (
    G5269,
    g841_n
  );


  buf

  (
    G5270,
    g850_n
  );


  buf

  (
    G5271,
    g859_n
  );


  buf

  (
    G5272,
    g868_n
  );


  buf

  (
    G5273,
    g877_n
  );


  buf

  (
    G5274,
    g886_n
  );


  buf

  (
    G5275,
    g896_p
  );


  buf

  (
    G5276,
    g906_p
  );


  buf

  (
    G5277,
    g916_p
  );


  buf

  (
    G5278,
    g926_p
  );


  buf

  (
    G5279,
    g936_p
  );


  buf

  (
    G5280,
    g946_p
  );


  buf

  (
    G5281,
    g956_p
  );


  buf

  (
    G5282,
    g966_p
  );


  buf

  (
    G5283,
    g980_p
  );


  buf

  (
    G5284,
    g983_n
  );


  not

  (
    G5285,
    g990_p_spl_1
  );


  not

  (
    G5286,
    g997_n_spl_1
  );


  not

  (
    G5287,
    g1004_n_spl_1
  );


  not

  (
    G5288,
    g1011_n_spl_1
  );


  not

  (
    G5289,
    g1018_n
  );


  not

  (
    G5290,
    g1025_n_spl_1
  );


  not

  (
    G5291,
    g1032_n_spl_1
  );


  not

  (
    G5292,
    g1039_n_spl_1
  );


  not

  (
    G5293,
    g1046_n_spl_1
  );


  buf

  (
    G5294,
    g1055_n
  );


  buf

  (
    G5295,
    g1064_n
  );


  buf

  (
    G5296,
    g1073_n
  );


  buf

  (
    G5297,
    g1082_n
  );


  buf

  (
    G5298,
    g1091_n
  );


  buf

  (
    G5299,
    g1100_n
  );


  buf

  (
    G5300,
    g1109_n
  );


  buf

  (
    G5301,
    g1118_n
  );


  buf

  (
    G5302,
    g1128_p
  );


  buf

  (
    G5303,
    g1138_p
  );


  buf

  (
    G5304,
    g1148_p
  );


  buf

  (
    G5305,
    g1158_p
  );


  buf

  (
    G5306,
    g1168_p
  );


  buf

  (
    G5307,
    g1178_p
  );


  buf

  (
    G5308,
    g1188_p
  );


  buf

  (
    G5309,
    g1198_p
  );


  buf

  (
    G5310,
    g1311_p
  );


  buf

  (
    G5311,
    g1503_p
  );


  not

  (
    G5312,
    g1516_p
  );


  not

  (
    G5313,
    g1525_p
  );


  buf

  (
    G5314,
    g1535_n
  );


  buf

  (
    G5315,
    g1545_n
  );


  buf

  (
    G153_n_spl_,
    G153_n
  );


  buf

  (
    G156_n_spl_,
    G156_n
  );


  buf

  (
    G66_p_spl_,
    G66_p
  );


  buf

  (
    G66_p_spl_0,
    G66_p_spl_
  );


  buf

  (
    G66_p_spl_00,
    G66_p_spl_0
  );


  buf

  (
    G66_p_spl_01,
    G66_p_spl_0
  );


  buf

  (
    G66_p_spl_1,
    G66_p_spl_
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G165_n_spl_,
    G165_n
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    g185_n_spl_,
    g185_n
  );


  buf

  (
    g185_n_spl_0,
    g185_n_spl_
  );


  buf

  (
    g185_n_spl_00,
    g185_n_spl_0
  );


  buf

  (
    g185_n_spl_000,
    g185_n_spl_00
  );


  buf

  (
    g185_n_spl_01,
    g185_n_spl_0
  );


  buf

  (
    g185_n_spl_1,
    g185_n_spl_
  );


  buf

  (
    g185_n_spl_10,
    g185_n_spl_1
  );


  buf

  (
    g185_n_spl_11,
    g185_n_spl_1
  );


  buf

  (
    G163_n_spl_,
    G163_n
  );


  buf

  (
    G163_n_spl_0,
    G163_n_spl_
  );


  buf

  (
    G163_n_spl_00,
    G163_n_spl_0
  );


  buf

  (
    G163_n_spl_01,
    G163_n_spl_0
  );


  buf

  (
    G163_n_spl_1,
    G163_n_spl_
  );


  buf

  (
    G163_p_spl_,
    G163_p
  );


  buf

  (
    G163_p_spl_0,
    G163_p_spl_
  );


  buf

  (
    G163_p_spl_00,
    G163_p_spl_0
  );


  buf

  (
    G163_p_spl_01,
    G163_p_spl_0
  );


  buf

  (
    G163_p_spl_1,
    G163_p_spl_
  );


  buf

  (
    G128_p_spl_,
    G128_p
  );


  buf

  (
    G128_p_spl_0,
    G128_p_spl_
  );


  buf

  (
    G128_p_spl_00,
    G128_p_spl_0
  );


  buf

  (
    G128_p_spl_000,
    G128_p_spl_00
  );


  buf

  (
    G128_p_spl_01,
    G128_p_spl_0
  );


  buf

  (
    G128_p_spl_1,
    G128_p_spl_
  );


  buf

  (
    G128_p_spl_10,
    G128_p_spl_1
  );


  buf

  (
    G128_p_spl_11,
    G128_p_spl_1
  );


  buf

  (
    G168_p_spl_,
    G168_p
  );


  buf

  (
    G168_p_spl_0,
    G168_p_spl_
  );


  buf

  (
    G168_p_spl_00,
    G168_p_spl_0
  );


  buf

  (
    G168_p_spl_000,
    G168_p_spl_00
  );


  buf

  (
    G168_p_spl_001,
    G168_p_spl_00
  );


  buf

  (
    G168_p_spl_01,
    G168_p_spl_0
  );


  buf

  (
    G168_p_spl_010,
    G168_p_spl_01
  );


  buf

  (
    G168_p_spl_1,
    G168_p_spl_
  );


  buf

  (
    G168_p_spl_10,
    G168_p_spl_1
  );


  buf

  (
    G168_p_spl_11,
    G168_p_spl_1
  );


  buf

  (
    G128_n_spl_,
    G128_n
  );


  buf

  (
    G128_n_spl_0,
    G128_n_spl_
  );


  buf

  (
    G128_n_spl_00,
    G128_n_spl_0
  );


  buf

  (
    G128_n_spl_000,
    G128_n_spl_00
  );


  buf

  (
    G128_n_spl_01,
    G128_n_spl_0
  );


  buf

  (
    G128_n_spl_1,
    G128_n_spl_
  );


  buf

  (
    G128_n_spl_10,
    G128_n_spl_1
  );


  buf

  (
    G128_n_spl_11,
    G128_n_spl_1
  );


  buf

  (
    G169_p_spl_,
    G169_p
  );


  buf

  (
    G169_p_spl_0,
    G169_p_spl_
  );


  buf

  (
    G169_p_spl_00,
    G169_p_spl_0
  );


  buf

  (
    G169_p_spl_000,
    G169_p_spl_00
  );


  buf

  (
    G169_p_spl_001,
    G169_p_spl_00
  );


  buf

  (
    G169_p_spl_01,
    G169_p_spl_0
  );


  buf

  (
    G169_p_spl_010,
    G169_p_spl_01
  );


  buf

  (
    G169_p_spl_011,
    G169_p_spl_01
  );


  buf

  (
    G169_p_spl_1,
    G169_p_spl_
  );


  buf

  (
    G169_p_spl_10,
    G169_p_spl_1
  );


  buf

  (
    G169_p_spl_11,
    G169_p_spl_1
  );


  buf

  (
    G150_p_spl_,
    G150_p
  );


  buf

  (
    G150_p_spl_0,
    G150_p_spl_
  );


  buf

  (
    G150_p_spl_00,
    G150_p_spl_0
  );


  buf

  (
    G150_p_spl_1,
    G150_p_spl_
  );


  buf

  (
    G167_n_spl_,
    G167_n
  );


  buf

  (
    G167_n_spl_0,
    G167_n_spl_
  );


  buf

  (
    G167_n_spl_00,
    G167_n_spl_0
  );


  buf

  (
    G167_n_spl_000,
    G167_n_spl_00
  );


  buf

  (
    G167_n_spl_001,
    G167_n_spl_00
  );


  buf

  (
    G167_n_spl_01,
    G167_n_spl_0
  );


  buf

  (
    G167_n_spl_010,
    G167_n_spl_01
  );


  buf

  (
    G167_n_spl_1,
    G167_n_spl_
  );


  buf

  (
    G167_n_spl_10,
    G167_n_spl_1
  );


  buf

  (
    G167_n_spl_11,
    G167_n_spl_1
  );


  buf

  (
    G166_n_spl_,
    G166_n
  );


  buf

  (
    G166_n_spl_0,
    G166_n_spl_
  );


  buf

  (
    G166_n_spl_00,
    G166_n_spl_0
  );


  buf

  (
    G166_n_spl_000,
    G166_n_spl_00
  );


  buf

  (
    G166_n_spl_001,
    G166_n_spl_00
  );


  buf

  (
    G166_n_spl_01,
    G166_n_spl_0
  );


  buf

  (
    G166_n_spl_010,
    G166_n_spl_01
  );


  buf

  (
    G166_n_spl_011,
    G166_n_spl_01
  );


  buf

  (
    G166_n_spl_1,
    G166_n_spl_
  );


  buf

  (
    G166_n_spl_10,
    G166_n_spl_1
  );


  buf

  (
    G166_n_spl_11,
    G166_n_spl_1
  );


  buf

  (
    G150_n_spl_,
    G150_n
  );


  buf

  (
    G150_n_spl_0,
    G150_n_spl_
  );


  buf

  (
    G150_n_spl_00,
    G150_n_spl_0
  );


  buf

  (
    G150_n_spl_1,
    G150_n_spl_
  );


  buf

  (
    G126_p_spl_,
    G126_p
  );


  buf

  (
    G126_p_spl_0,
    G126_p_spl_
  );


  buf

  (
    G126_p_spl_00,
    G126_p_spl_0
  );


  buf

  (
    G126_p_spl_000,
    G126_p_spl_00
  );


  buf

  (
    G126_p_spl_01,
    G126_p_spl_0
  );


  buf

  (
    G126_p_spl_1,
    G126_p_spl_
  );


  buf

  (
    G126_p_spl_10,
    G126_p_spl_1
  );


  buf

  (
    G126_p_spl_11,
    G126_p_spl_1
  );


  buf

  (
    G126_n_spl_,
    G126_n
  );


  buf

  (
    G126_n_spl_0,
    G126_n_spl_
  );


  buf

  (
    G126_n_spl_00,
    G126_n_spl_0
  );


  buf

  (
    G126_n_spl_000,
    G126_n_spl_00
  );


  buf

  (
    G126_n_spl_01,
    G126_n_spl_0
  );


  buf

  (
    G126_n_spl_1,
    G126_n_spl_
  );


  buf

  (
    G126_n_spl_10,
    G126_n_spl_1
  );


  buf

  (
    G126_n_spl_11,
    G126_n_spl_1
  );


  buf

  (
    G149_p_spl_,
    G149_p
  );


  buf

  (
    G149_p_spl_0,
    G149_p_spl_
  );


  buf

  (
    G149_p_spl_00,
    G149_p_spl_0
  );


  buf

  (
    G149_p_spl_1,
    G149_p_spl_
  );


  buf

  (
    G149_n_spl_,
    G149_n
  );


  buf

  (
    G149_n_spl_0,
    G149_n_spl_
  );


  buf

  (
    G149_n_spl_00,
    G149_n_spl_0
  );


  buf

  (
    G149_n_spl_1,
    G149_n_spl_
  );


  buf

  (
    g224_n_spl_,
    g224_n
  );


  buf

  (
    g233_n_spl_,
    g233_n
  );


  buf

  (
    G102_p_spl_,
    G102_p
  );


  buf

  (
    G102_p_spl_0,
    G102_p_spl_
  );


  buf

  (
    G102_p_spl_00,
    G102_p_spl_0
  );


  buf

  (
    G102_p_spl_000,
    G102_p_spl_00
  );


  buf

  (
    G102_p_spl_001,
    G102_p_spl_00
  );


  buf

  (
    G102_p_spl_01,
    G102_p_spl_0
  );


  buf

  (
    G102_p_spl_010,
    G102_p_spl_01
  );


  buf

  (
    G102_p_spl_011,
    G102_p_spl_01
  );


  buf

  (
    G102_p_spl_1,
    G102_p_spl_
  );


  buf

  (
    G102_p_spl_10,
    G102_p_spl_1
  );


  buf

  (
    G102_p_spl_100,
    G102_p_spl_10
  );


  buf

  (
    G102_p_spl_101,
    G102_p_spl_10
  );


  buf

  (
    G102_p_spl_11,
    G102_p_spl_1
  );


  buf

  (
    G102_p_spl_110,
    G102_p_spl_11
  );


  buf

  (
    G113_p_spl_,
    G113_p
  );


  buf

  (
    G113_p_spl_0,
    G113_p_spl_
  );


  buf

  (
    G113_p_spl_00,
    G113_p_spl_0
  );


  buf

  (
    G113_p_spl_1,
    G113_p_spl_
  );


  buf

  (
    G102_n_spl_,
    G102_n
  );


  buf

  (
    G102_n_spl_0,
    G102_n_spl_
  );


  buf

  (
    G102_n_spl_00,
    G102_n_spl_0
  );


  buf

  (
    G102_n_spl_000,
    G102_n_spl_00
  );


  buf

  (
    G102_n_spl_001,
    G102_n_spl_00
  );


  buf

  (
    G102_n_spl_01,
    G102_n_spl_0
  );


  buf

  (
    G102_n_spl_010,
    G102_n_spl_01
  );


  buf

  (
    G102_n_spl_011,
    G102_n_spl_01
  );


  buf

  (
    G102_n_spl_1,
    G102_n_spl_
  );


  buf

  (
    G102_n_spl_10,
    G102_n_spl_1
  );


  buf

  (
    G102_n_spl_100,
    G102_n_spl_10
  );


  buf

  (
    G102_n_spl_101,
    G102_n_spl_10
  );


  buf

  (
    G102_n_spl_11,
    G102_n_spl_1
  );


  buf

  (
    G102_n_spl_110,
    G102_n_spl_11
  );


  buf

  (
    G113_n_spl_,
    G113_n
  );


  buf

  (
    G113_n_spl_0,
    G113_n_spl_
  );


  buf

  (
    G113_n_spl_00,
    G113_n_spl_0
  );


  buf

  (
    G113_n_spl_01,
    G113_n_spl_0
  );


  buf

  (
    G113_n_spl_1,
    G113_n_spl_
  );


  buf

  (
    G98_p_spl_,
    G98_p
  );


  buf

  (
    G98_p_spl_0,
    G98_p_spl_
  );


  buf

  (
    G98_p_spl_00,
    G98_p_spl_0
  );


  buf

  (
    G98_p_spl_000,
    G98_p_spl_00
  );


  buf

  (
    G98_p_spl_001,
    G98_p_spl_00
  );


  buf

  (
    G98_p_spl_01,
    G98_p_spl_0
  );


  buf

  (
    G98_p_spl_010,
    G98_p_spl_01
  );


  buf

  (
    G98_p_spl_011,
    G98_p_spl_01
  );


  buf

  (
    G98_p_spl_1,
    G98_p_spl_
  );


  buf

  (
    G98_p_spl_10,
    G98_p_spl_1
  );


  buf

  (
    G98_p_spl_100,
    G98_p_spl_10
  );


  buf

  (
    G98_p_spl_101,
    G98_p_spl_10
  );


  buf

  (
    G98_p_spl_11,
    G98_p_spl_1
  );


  buf

  (
    G98_p_spl_110,
    G98_p_spl_11
  );


  buf

  (
    G98_p_spl_111,
    G98_p_spl_11
  );


  buf

  (
    G98_n_spl_,
    G98_n
  );


  buf

  (
    G98_n_spl_0,
    G98_n_spl_
  );


  buf

  (
    G98_n_spl_00,
    G98_n_spl_0
  );


  buf

  (
    G98_n_spl_000,
    G98_n_spl_00
  );


  buf

  (
    G98_n_spl_001,
    G98_n_spl_00
  );


  buf

  (
    G98_n_spl_01,
    G98_n_spl_0
  );


  buf

  (
    G98_n_spl_010,
    G98_n_spl_01
  );


  buf

  (
    G98_n_spl_011,
    G98_n_spl_01
  );


  buf

  (
    G98_n_spl_1,
    G98_n_spl_
  );


  buf

  (
    G98_n_spl_10,
    G98_n_spl_1
  );


  buf

  (
    G98_n_spl_100,
    G98_n_spl_10
  );


  buf

  (
    G98_n_spl_101,
    G98_n_spl_10
  );


  buf

  (
    G98_n_spl_11,
    G98_n_spl_1
  );


  buf

  (
    G98_n_spl_110,
    G98_n_spl_11
  );


  buf

  (
    G98_n_spl_111,
    G98_n_spl_11
  );


  buf

  (
    G101_p_spl_,
    G101_p
  );


  buf

  (
    G101_p_spl_0,
    G101_p_spl_
  );


  buf

  (
    G101_p_spl_00,
    G101_p_spl_0
  );


  buf

  (
    G101_p_spl_000,
    G101_p_spl_00
  );


  buf

  (
    G101_p_spl_001,
    G101_p_spl_00
  );


  buf

  (
    G101_p_spl_01,
    G101_p_spl_0
  );


  buf

  (
    G101_p_spl_010,
    G101_p_spl_01
  );


  buf

  (
    G101_p_spl_011,
    G101_p_spl_01
  );


  buf

  (
    G101_p_spl_1,
    G101_p_spl_
  );


  buf

  (
    G101_p_spl_10,
    G101_p_spl_1
  );


  buf

  (
    G101_p_spl_100,
    G101_p_spl_10
  );


  buf

  (
    G101_p_spl_101,
    G101_p_spl_10
  );


  buf

  (
    G101_p_spl_11,
    G101_p_spl_1
  );


  buf

  (
    G101_p_spl_110,
    G101_p_spl_11
  );


  buf

  (
    G101_p_spl_111,
    G101_p_spl_11
  );


  buf

  (
    G115_p_spl_,
    G115_p
  );


  buf

  (
    G115_p_spl_0,
    G115_p_spl_
  );


  buf

  (
    G115_p_spl_00,
    G115_p_spl_0
  );


  buf

  (
    G115_p_spl_1,
    G115_p_spl_
  );


  buf

  (
    G101_n_spl_,
    G101_n
  );


  buf

  (
    G101_n_spl_0,
    G101_n_spl_
  );


  buf

  (
    G101_n_spl_00,
    G101_n_spl_0
  );


  buf

  (
    G101_n_spl_000,
    G101_n_spl_00
  );


  buf

  (
    G101_n_spl_001,
    G101_n_spl_00
  );


  buf

  (
    G101_n_spl_01,
    G101_n_spl_0
  );


  buf

  (
    G101_n_spl_010,
    G101_n_spl_01
  );


  buf

  (
    G101_n_spl_011,
    G101_n_spl_01
  );


  buf

  (
    G101_n_spl_1,
    G101_n_spl_
  );


  buf

  (
    G101_n_spl_10,
    G101_n_spl_1
  );


  buf

  (
    G101_n_spl_100,
    G101_n_spl_10
  );


  buf

  (
    G101_n_spl_101,
    G101_n_spl_10
  );


  buf

  (
    G101_n_spl_11,
    G101_n_spl_1
  );


  buf

  (
    G101_n_spl_110,
    G101_n_spl_11
  );


  buf

  (
    G101_n_spl_111,
    G101_n_spl_11
  );


  buf

  (
    G115_n_spl_,
    G115_n
  );


  buf

  (
    G115_n_spl_0,
    G115_n_spl_
  );


  buf

  (
    G115_n_spl_00,
    G115_n_spl_0
  );


  buf

  (
    G115_n_spl_1,
    G115_n_spl_
  );


  buf

  (
    G100_p_spl_,
    G100_p
  );


  buf

  (
    G100_p_spl_0,
    G100_p_spl_
  );


  buf

  (
    G100_p_spl_00,
    G100_p_spl_0
  );


  buf

  (
    G100_p_spl_000,
    G100_p_spl_00
  );


  buf

  (
    G100_p_spl_0000,
    G100_p_spl_000
  );


  buf

  (
    G100_p_spl_001,
    G100_p_spl_00
  );


  buf

  (
    G100_p_spl_01,
    G100_p_spl_0
  );


  buf

  (
    G100_p_spl_010,
    G100_p_spl_01
  );


  buf

  (
    G100_p_spl_011,
    G100_p_spl_01
  );


  buf

  (
    G100_p_spl_1,
    G100_p_spl_
  );


  buf

  (
    G100_p_spl_10,
    G100_p_spl_1
  );


  buf

  (
    G100_p_spl_100,
    G100_p_spl_10
  );


  buf

  (
    G100_p_spl_101,
    G100_p_spl_10
  );


  buf

  (
    G100_p_spl_11,
    G100_p_spl_1
  );


  buf

  (
    G100_p_spl_110,
    G100_p_spl_11
  );


  buf

  (
    G100_p_spl_111,
    G100_p_spl_11
  );


  buf

  (
    G100_n_spl_,
    G100_n
  );


  buf

  (
    G100_n_spl_0,
    G100_n_spl_
  );


  buf

  (
    G100_n_spl_00,
    G100_n_spl_0
  );


  buf

  (
    G100_n_spl_000,
    G100_n_spl_00
  );


  buf

  (
    G100_n_spl_0000,
    G100_n_spl_000
  );


  buf

  (
    G100_n_spl_001,
    G100_n_spl_00
  );


  buf

  (
    G100_n_spl_01,
    G100_n_spl_0
  );


  buf

  (
    G100_n_spl_010,
    G100_n_spl_01
  );


  buf

  (
    G100_n_spl_011,
    G100_n_spl_01
  );


  buf

  (
    G100_n_spl_1,
    G100_n_spl_
  );


  buf

  (
    G100_n_spl_10,
    G100_n_spl_1
  );


  buf

  (
    G100_n_spl_100,
    G100_n_spl_10
  );


  buf

  (
    G100_n_spl_101,
    G100_n_spl_10
  );


  buf

  (
    G100_n_spl_11,
    G100_n_spl_1
  );


  buf

  (
    G100_n_spl_110,
    G100_n_spl_11
  );


  buf

  (
    G100_n_spl_111,
    G100_n_spl_11
  );


  buf

  (
    g237_n_spl_,
    g237_n
  );


  buf

  (
    g237_n_spl_0,
    g237_n_spl_
  );


  buf

  (
    g237_n_spl_1,
    g237_n_spl_
  );


  buf

  (
    g240_p_spl_,
    g240_p
  );


  buf

  (
    g237_p_spl_,
    g237_p
  );


  buf

  (
    g240_n_spl_,
    g240_n
  );


  buf

  (
    g240_n_spl_0,
    g240_n_spl_
  );


  buf

  (
    g241_n_spl_,
    g241_n
  );


  buf

  (
    G130_p_spl_,
    G130_p
  );


  buf

  (
    G130_p_spl_0,
    G130_p_spl_
  );


  buf

  (
    G130_p_spl_00,
    G130_p_spl_0
  );


  buf

  (
    G130_p_spl_1,
    G130_p_spl_
  );


  buf

  (
    G130_n_spl_,
    G130_n
  );


  buf

  (
    G130_n_spl_0,
    G130_n_spl_
  );


  buf

  (
    G130_n_spl_00,
    G130_n_spl_0
  );


  buf

  (
    G130_n_spl_1,
    G130_n_spl_
  );


  buf

  (
    G148_n_spl_,
    G148_n
  );


  buf

  (
    G148_n_spl_0,
    G148_n_spl_
  );


  buf

  (
    G148_n_spl_00,
    G148_n_spl_0
  );


  buf

  (
    G148_n_spl_1,
    G148_n_spl_
  );


  buf

  (
    G148_p_spl_,
    G148_p
  );


  buf

  (
    G148_p_spl_0,
    G148_p_spl_
  );


  buf

  (
    G148_p_spl_00,
    G148_p_spl_0
  );


  buf

  (
    G148_p_spl_1,
    G148_p_spl_
  );


  buf

  (
    g245_n_spl_,
    g245_n
  );


  buf

  (
    g245_n_spl_0,
    g245_n_spl_
  );


  buf

  (
    g245_n_spl_1,
    g245_n_spl_
  );


  buf

  (
    g248_n_spl_,
    g248_n
  );


  buf

  (
    G119_p_spl_,
    G119_p
  );


  buf

  (
    G119_p_spl_0,
    G119_p_spl_
  );


  buf

  (
    G119_p_spl_00,
    G119_p_spl_0
  );


  buf

  (
    G119_p_spl_01,
    G119_p_spl_0
  );


  buf

  (
    G119_p_spl_1,
    G119_p_spl_
  );


  buf

  (
    G119_p_spl_10,
    G119_p_spl_1
  );


  buf

  (
    G119_n_spl_,
    G119_n
  );


  buf

  (
    G119_n_spl_0,
    G119_n_spl_
  );


  buf

  (
    G119_n_spl_00,
    G119_n_spl_0
  );


  buf

  (
    G119_n_spl_01,
    G119_n_spl_0
  );


  buf

  (
    G119_n_spl_1,
    G119_n_spl_
  );


  buf

  (
    G119_n_spl_10,
    G119_n_spl_1
  );


  buf

  (
    G146_p_spl_,
    G146_p
  );


  buf

  (
    G146_p_spl_0,
    G146_p_spl_
  );


  buf

  (
    G146_p_spl_1,
    G146_p_spl_
  );


  buf

  (
    G146_n_spl_,
    G146_n
  );


  buf

  (
    G146_n_spl_0,
    G146_n_spl_
  );


  buf

  (
    G146_n_spl_1,
    G146_n_spl_
  );


  buf

  (
    G117_p_spl_,
    G117_p
  );


  buf

  (
    G117_p_spl_0,
    G117_p_spl_
  );


  buf

  (
    G117_p_spl_00,
    G117_p_spl_0
  );


  buf

  (
    G117_p_spl_01,
    G117_p_spl_0
  );


  buf

  (
    G117_p_spl_1,
    G117_p_spl_
  );


  buf

  (
    G117_p_spl_10,
    G117_p_spl_1
  );


  buf

  (
    G117_n_spl_,
    G117_n
  );


  buf

  (
    G117_n_spl_0,
    G117_n_spl_
  );


  buf

  (
    G117_n_spl_00,
    G117_n_spl_0
  );


  buf

  (
    G117_n_spl_01,
    G117_n_spl_0
  );


  buf

  (
    G117_n_spl_1,
    G117_n_spl_
  );


  buf

  (
    G117_n_spl_10,
    G117_n_spl_1
  );


  buf

  (
    G145_p_spl_,
    G145_p
  );


  buf

  (
    G145_p_spl_0,
    G145_p_spl_
  );


  buf

  (
    G145_p_spl_1,
    G145_p_spl_
  );


  buf

  (
    G145_n_spl_,
    G145_n
  );


  buf

  (
    G145_n_spl_0,
    G145_n_spl_
  );


  buf

  (
    G145_n_spl_1,
    G145_n_spl_
  );


  buf

  (
    g258_p_spl_,
    g258_p
  );


  buf

  (
    g267_p_spl_,
    g267_p
  );


  buf

  (
    g258_n_spl_,
    g258_n
  );


  buf

  (
    g258_n_spl_0,
    g258_n_spl_
  );


  buf

  (
    g267_n_spl_,
    g267_n
  );


  buf

  (
    g267_n_spl_0,
    g267_n_spl_
  );


  buf

  (
    G121_p_spl_,
    G121_p
  );


  buf

  (
    G121_p_spl_0,
    G121_p_spl_
  );


  buf

  (
    G121_p_spl_00,
    G121_p_spl_0
  );


  buf

  (
    G121_p_spl_000,
    G121_p_spl_00
  );


  buf

  (
    G121_p_spl_01,
    G121_p_spl_0
  );


  buf

  (
    G121_p_spl_1,
    G121_p_spl_
  );


  buf

  (
    G121_p_spl_10,
    G121_p_spl_1
  );


  buf

  (
    G121_p_spl_11,
    G121_p_spl_1
  );


  buf

  (
    G121_n_spl_,
    G121_n
  );


  buf

  (
    G121_n_spl_0,
    G121_n_spl_
  );


  buf

  (
    G121_n_spl_00,
    G121_n_spl_0
  );


  buf

  (
    G121_n_spl_000,
    G121_n_spl_00
  );


  buf

  (
    G121_n_spl_01,
    G121_n_spl_0
  );


  buf

  (
    G121_n_spl_1,
    G121_n_spl_
  );


  buf

  (
    G121_n_spl_10,
    G121_n_spl_1
  );


  buf

  (
    G121_n_spl_11,
    G121_n_spl_1
  );


  buf

  (
    G147_p_spl_,
    G147_p
  );


  buf

  (
    G147_p_spl_0,
    G147_p_spl_
  );


  buf

  (
    G147_p_spl_00,
    G147_p_spl_0
  );


  buf

  (
    G147_p_spl_1,
    G147_p_spl_
  );


  buf

  (
    G147_n_spl_,
    G147_n
  );


  buf

  (
    G147_n_spl_0,
    G147_n_spl_
  );


  buf

  (
    G147_n_spl_00,
    G147_n_spl_0
  );


  buf

  (
    G147_n_spl_1,
    G147_n_spl_
  );


  buf

  (
    g268_n_spl_,
    g268_n
  );


  buf

  (
    g277_n_spl_,
    g277_n
  );


  buf

  (
    G107_p_spl_,
    G107_p
  );


  buf

  (
    G107_p_spl_0,
    G107_p_spl_
  );


  buf

  (
    G107_p_spl_00,
    G107_p_spl_0
  );


  buf

  (
    G107_p_spl_000,
    G107_p_spl_00
  );


  buf

  (
    G107_p_spl_01,
    G107_p_spl_0
  );


  buf

  (
    G107_p_spl_1,
    G107_p_spl_
  );


  buf

  (
    G107_p_spl_10,
    G107_p_spl_1
  );


  buf

  (
    G107_p_spl_11,
    G107_p_spl_1
  );


  buf

  (
    G107_n_spl_,
    G107_n
  );


  buf

  (
    G107_n_spl_0,
    G107_n_spl_
  );


  buf

  (
    G107_n_spl_00,
    G107_n_spl_0
  );


  buf

  (
    G107_n_spl_000,
    G107_n_spl_00
  );


  buf

  (
    G107_n_spl_01,
    G107_n_spl_0
  );


  buf

  (
    G107_n_spl_1,
    G107_n_spl_
  );


  buf

  (
    G107_n_spl_10,
    G107_n_spl_1
  );


  buf

  (
    G107_n_spl_11,
    G107_n_spl_1
  );


  buf

  (
    G139_p_spl_,
    G139_p
  );


  buf

  (
    G139_p_spl_0,
    G139_p_spl_
  );


  buf

  (
    G139_p_spl_00,
    G139_p_spl_0
  );


  buf

  (
    G139_p_spl_1,
    G139_p_spl_
  );


  buf

  (
    G139_n_spl_,
    G139_n
  );


  buf

  (
    G139_n_spl_0,
    G139_n_spl_
  );


  buf

  (
    G139_n_spl_00,
    G139_n_spl_0
  );


  buf

  (
    G139_n_spl_1,
    G139_n_spl_
  );


  buf

  (
    G105_p_spl_,
    G105_p
  );


  buf

  (
    G105_p_spl_0,
    G105_p_spl_
  );


  buf

  (
    G105_p_spl_00,
    G105_p_spl_0
  );


  buf

  (
    G105_p_spl_000,
    G105_p_spl_00
  );


  buf

  (
    G105_p_spl_01,
    G105_p_spl_0
  );


  buf

  (
    G105_p_spl_1,
    G105_p_spl_
  );


  buf

  (
    G105_p_spl_10,
    G105_p_spl_1
  );


  buf

  (
    G105_p_spl_11,
    G105_p_spl_1
  );


  buf

  (
    G105_n_spl_,
    G105_n
  );


  buf

  (
    G105_n_spl_0,
    G105_n_spl_
  );


  buf

  (
    G105_n_spl_00,
    G105_n_spl_0
  );


  buf

  (
    G105_n_spl_000,
    G105_n_spl_00
  );


  buf

  (
    G105_n_spl_01,
    G105_n_spl_0
  );


  buf

  (
    G105_n_spl_1,
    G105_n_spl_
  );


  buf

  (
    G105_n_spl_10,
    G105_n_spl_1
  );


  buf

  (
    G105_n_spl_11,
    G105_n_spl_1
  );


  buf

  (
    G138_p_spl_,
    G138_p
  );


  buf

  (
    G138_p_spl_0,
    G138_p_spl_
  );


  buf

  (
    G138_p_spl_00,
    G138_p_spl_0
  );


  buf

  (
    G138_p_spl_1,
    G138_p_spl_
  );


  buf

  (
    G138_n_spl_,
    G138_n
  );


  buf

  (
    G138_n_spl_0,
    G138_n_spl_
  );


  buf

  (
    G138_n_spl_00,
    G138_n_spl_0
  );


  buf

  (
    G138_n_spl_1,
    G138_n_spl_
  );


  buf

  (
    g289_n_spl_,
    g289_n
  );


  buf

  (
    g298_n_spl_,
    g298_n
  );


  buf

  (
    G109_p_spl_,
    G109_p
  );


  buf

  (
    G109_p_spl_0,
    G109_p_spl_
  );


  buf

  (
    G109_p_spl_00,
    G109_p_spl_0
  );


  buf

  (
    G109_p_spl_000,
    G109_p_spl_00
  );


  buf

  (
    G109_p_spl_01,
    G109_p_spl_0
  );


  buf

  (
    G109_p_spl_1,
    G109_p_spl_
  );


  buf

  (
    G109_p_spl_10,
    G109_p_spl_1
  );


  buf

  (
    G109_p_spl_11,
    G109_p_spl_1
  );


  buf

  (
    G109_n_spl_,
    G109_n
  );


  buf

  (
    G109_n_spl_0,
    G109_n_spl_
  );


  buf

  (
    G109_n_spl_00,
    G109_n_spl_0
  );


  buf

  (
    G109_n_spl_000,
    G109_n_spl_00
  );


  buf

  (
    G109_n_spl_01,
    G109_n_spl_0
  );


  buf

  (
    G109_n_spl_1,
    G109_n_spl_
  );


  buf

  (
    G109_n_spl_10,
    G109_n_spl_1
  );


  buf

  (
    G109_n_spl_11,
    G109_n_spl_1
  );


  buf

  (
    G135_p_spl_,
    G135_p
  );


  buf

  (
    G135_p_spl_0,
    G135_p_spl_
  );


  buf

  (
    G135_p_spl_00,
    G135_p_spl_0
  );


  buf

  (
    G135_p_spl_1,
    G135_p_spl_
  );


  buf

  (
    G135_n_spl_,
    G135_n
  );


  buf

  (
    G135_n_spl_0,
    G135_n_spl_
  );


  buf

  (
    G135_n_spl_00,
    G135_n_spl_0
  );


  buf

  (
    G135_n_spl_1,
    G135_n_spl_
  );


  buf

  (
    G88_p_spl_,
    G88_p
  );


  buf

  (
    G88_p_spl_0,
    G88_p_spl_
  );


  buf

  (
    G88_p_spl_00,
    G88_p_spl_0
  );


  buf

  (
    G88_p_spl_01,
    G88_p_spl_0
  );


  buf

  (
    G88_p_spl_1,
    G88_p_spl_
  );


  buf

  (
    G88_p_spl_10,
    G88_p_spl_1
  );


  buf

  (
    G88_n_spl_,
    G88_n
  );


  buf

  (
    G88_n_spl_0,
    G88_n_spl_
  );


  buf

  (
    G88_n_spl_00,
    G88_n_spl_0
  );


  buf

  (
    G88_n_spl_01,
    G88_n_spl_0
  );


  buf

  (
    G88_n_spl_1,
    G88_n_spl_
  );


  buf

  (
    G88_n_spl_10,
    G88_n_spl_1
  );


  buf

  (
    G142_p_spl_,
    G142_p
  );


  buf

  (
    G142_p_spl_0,
    G142_p_spl_
  );


  buf

  (
    G142_p_spl_1,
    G142_p_spl_
  );


  buf

  (
    G142_n_spl_,
    G142_n
  );


  buf

  (
    G142_n_spl_0,
    G142_n_spl_
  );


  buf

  (
    G142_n_spl_1,
    G142_n_spl_
  );


  buf

  (
    g308_n_spl_,
    g308_n
  );


  buf

  (
    g317_n_spl_,
    g317_n
  );


  buf

  (
    g317_n_spl_0,
    g317_n_spl_
  );


  buf

  (
    g317_n_spl_1,
    g317_n_spl_
  );


  buf

  (
    G90_p_spl_,
    G90_p
  );


  buf

  (
    G90_p_spl_0,
    G90_p_spl_
  );


  buf

  (
    G90_p_spl_00,
    G90_p_spl_0
  );


  buf

  (
    G90_p_spl_000,
    G90_p_spl_00
  );


  buf

  (
    G90_p_spl_01,
    G90_p_spl_0
  );


  buf

  (
    G90_p_spl_1,
    G90_p_spl_
  );


  buf

  (
    G90_p_spl_10,
    G90_p_spl_1
  );


  buf

  (
    G90_p_spl_11,
    G90_p_spl_1
  );


  buf

  (
    G90_n_spl_,
    G90_n
  );


  buf

  (
    G90_n_spl_0,
    G90_n_spl_
  );


  buf

  (
    G90_n_spl_00,
    G90_n_spl_0
  );


  buf

  (
    G90_n_spl_000,
    G90_n_spl_00
  );


  buf

  (
    G90_n_spl_01,
    G90_n_spl_0
  );


  buf

  (
    G90_n_spl_1,
    G90_n_spl_
  );


  buf

  (
    G90_n_spl_10,
    G90_n_spl_1
  );


  buf

  (
    G90_n_spl_11,
    G90_n_spl_1
  );


  buf

  (
    G143_p_spl_,
    G143_p
  );


  buf

  (
    G143_p_spl_0,
    G143_p_spl_
  );


  buf

  (
    G143_p_spl_00,
    G143_p_spl_0
  );


  buf

  (
    G143_p_spl_1,
    G143_p_spl_
  );


  buf

  (
    G143_n_spl_,
    G143_n
  );


  buf

  (
    G143_n_spl_0,
    G143_n_spl_
  );


  buf

  (
    G143_n_spl_00,
    G143_n_spl_0
  );


  buf

  (
    G143_n_spl_1,
    G143_n_spl_
  );


  buf

  (
    G92_p_spl_,
    G92_p
  );


  buf

  (
    G92_p_spl_0,
    G92_p_spl_
  );


  buf

  (
    G92_p_spl_00,
    G92_p_spl_0
  );


  buf

  (
    G92_p_spl_000,
    G92_p_spl_00
  );


  buf

  (
    G92_p_spl_01,
    G92_p_spl_0
  );


  buf

  (
    G92_p_spl_1,
    G92_p_spl_
  );


  buf

  (
    G92_p_spl_10,
    G92_p_spl_1
  );


  buf

  (
    G92_p_spl_11,
    G92_p_spl_1
  );


  buf

  (
    G92_n_spl_,
    G92_n
  );


  buf

  (
    G92_n_spl_0,
    G92_n_spl_
  );


  buf

  (
    G92_n_spl_00,
    G92_n_spl_0
  );


  buf

  (
    G92_n_spl_000,
    G92_n_spl_00
  );


  buf

  (
    G92_n_spl_01,
    G92_n_spl_0
  );


  buf

  (
    G92_n_spl_1,
    G92_n_spl_
  );


  buf

  (
    G92_n_spl_10,
    G92_n_spl_1
  );


  buf

  (
    G92_n_spl_11,
    G92_n_spl_1
  );


  buf

  (
    G144_p_spl_,
    G144_p
  );


  buf

  (
    G144_p_spl_0,
    G144_p_spl_
  );


  buf

  (
    G144_p_spl_00,
    G144_p_spl_0
  );


  buf

  (
    G144_p_spl_1,
    G144_p_spl_
  );


  buf

  (
    G144_n_spl_,
    G144_n
  );


  buf

  (
    G144_n_spl_0,
    G144_n_spl_
  );


  buf

  (
    G144_n_spl_00,
    G144_n_spl_0
  );


  buf

  (
    G144_n_spl_1,
    G144_n_spl_
  );


  buf

  (
    g328_n_spl_,
    g328_n
  );


  buf

  (
    g337_n_spl_,
    g337_n
  );


  buf

  (
    G94_p_spl_,
    G94_p
  );


  buf

  (
    G94_p_spl_0,
    G94_p_spl_
  );


  buf

  (
    G94_p_spl_00,
    G94_p_spl_0
  );


  buf

  (
    G94_p_spl_000,
    G94_p_spl_00
  );


  buf

  (
    G94_p_spl_01,
    G94_p_spl_0
  );


  buf

  (
    G94_p_spl_1,
    G94_p_spl_
  );


  buf

  (
    G94_p_spl_10,
    G94_p_spl_1
  );


  buf

  (
    G94_p_spl_11,
    G94_p_spl_1
  );


  buf

  (
    G94_n_spl_,
    G94_n
  );


  buf

  (
    G94_n_spl_0,
    G94_n_spl_
  );


  buf

  (
    G94_n_spl_00,
    G94_n_spl_0
  );


  buf

  (
    G94_n_spl_000,
    G94_n_spl_00
  );


  buf

  (
    G94_n_spl_01,
    G94_n_spl_0
  );


  buf

  (
    G94_n_spl_1,
    G94_n_spl_
  );


  buf

  (
    G94_n_spl_10,
    G94_n_spl_1
  );


  buf

  (
    G94_n_spl_11,
    G94_n_spl_1
  );


  buf

  (
    G140_p_spl_,
    G140_p
  );


  buf

  (
    G140_p_spl_0,
    G140_p_spl_
  );


  buf

  (
    G140_p_spl_00,
    G140_p_spl_0
  );


  buf

  (
    G140_p_spl_1,
    G140_p_spl_
  );


  buf

  (
    G140_n_spl_,
    G140_n
  );


  buf

  (
    G140_n_spl_0,
    G140_n_spl_
  );


  buf

  (
    G140_n_spl_00,
    G140_n_spl_0
  );


  buf

  (
    G140_n_spl_1,
    G140_n_spl_
  );


  buf

  (
    G96_p_spl_,
    G96_p
  );


  buf

  (
    G96_p_spl_0,
    G96_p_spl_
  );


  buf

  (
    G96_p_spl_00,
    G96_p_spl_0
  );


  buf

  (
    G96_p_spl_000,
    G96_p_spl_00
  );


  buf

  (
    G96_p_spl_01,
    G96_p_spl_0
  );


  buf

  (
    G96_p_spl_1,
    G96_p_spl_
  );


  buf

  (
    G96_p_spl_10,
    G96_p_spl_1
  );


  buf

  (
    G96_p_spl_11,
    G96_p_spl_1
  );


  buf

  (
    G96_n_spl_,
    G96_n
  );


  buf

  (
    G96_n_spl_0,
    G96_n_spl_
  );


  buf

  (
    G96_n_spl_00,
    G96_n_spl_0
  );


  buf

  (
    G96_n_spl_000,
    G96_n_spl_00
  );


  buf

  (
    G96_n_spl_01,
    G96_n_spl_0
  );


  buf

  (
    G96_n_spl_1,
    G96_n_spl_
  );


  buf

  (
    G96_n_spl_10,
    G96_n_spl_1
  );


  buf

  (
    G96_n_spl_11,
    G96_n_spl_1
  );


  buf

  (
    G141_p_spl_,
    G141_p
  );


  buf

  (
    G141_p_spl_0,
    G141_p_spl_
  );


  buf

  (
    G141_p_spl_00,
    G141_p_spl_0
  );


  buf

  (
    G141_p_spl_1,
    G141_p_spl_
  );


  buf

  (
    G141_n_spl_,
    G141_n
  );


  buf

  (
    G141_n_spl_0,
    G141_n_spl_
  );


  buf

  (
    G141_n_spl_00,
    G141_n_spl_0
  );


  buf

  (
    G141_n_spl_1,
    G141_n_spl_
  );


  buf

  (
    G103_p_spl_,
    G103_p
  );


  buf

  (
    G103_p_spl_0,
    G103_p_spl_
  );


  buf

  (
    G103_p_spl_00,
    G103_p_spl_0
  );


  buf

  (
    G103_p_spl_000,
    G103_p_spl_00
  );


  buf

  (
    G103_p_spl_01,
    G103_p_spl_0
  );


  buf

  (
    G103_p_spl_1,
    G103_p_spl_
  );


  buf

  (
    G103_p_spl_10,
    G103_p_spl_1
  );


  buf

  (
    G103_p_spl_11,
    G103_p_spl_1
  );


  buf

  (
    G103_n_spl_,
    G103_n
  );


  buf

  (
    G103_n_spl_0,
    G103_n_spl_
  );


  buf

  (
    G103_n_spl_00,
    G103_n_spl_0
  );


  buf

  (
    G103_n_spl_000,
    G103_n_spl_00
  );


  buf

  (
    G103_n_spl_01,
    G103_n_spl_0
  );


  buf

  (
    G103_n_spl_1,
    G103_n_spl_
  );


  buf

  (
    G103_n_spl_10,
    G103_n_spl_1
  );


  buf

  (
    G103_n_spl_11,
    G103_n_spl_1
  );


  buf

  (
    G137_p_spl_,
    G137_p
  );


  buf

  (
    G137_p_spl_0,
    G137_p_spl_
  );


  buf

  (
    G137_p_spl_00,
    G137_p_spl_0
  );


  buf

  (
    G137_p_spl_1,
    G137_p_spl_
  );


  buf

  (
    G137_n_spl_,
    G137_n
  );


  buf

  (
    G137_n_spl_0,
    G137_n_spl_
  );


  buf

  (
    G137_n_spl_00,
    G137_n_spl_0
  );


  buf

  (
    G137_n_spl_1,
    G137_n_spl_
  );


  buf

  (
    g356_n_spl_,
    g356_n
  );


  buf

  (
    g365_n_spl_,
    g365_n
  );


  buf

  (
    g347_n_spl_,
    g347_n
  );


  buf

  (
    G124_n_spl_,
    G124_n
  );


  buf

  (
    G124_n_spl_0,
    G124_n_spl_
  );


  buf

  (
    G124_n_spl_00,
    G124_n_spl_0
  );


  buf

  (
    G124_n_spl_000,
    G124_n_spl_00
  );


  buf

  (
    G124_n_spl_0000,
    G124_n_spl_000
  );


  buf

  (
    G124_n_spl_0001,
    G124_n_spl_000
  );


  buf

  (
    G124_n_spl_001,
    G124_n_spl_00
  );


  buf

  (
    G124_n_spl_0010,
    G124_n_spl_001
  );


  buf

  (
    G124_n_spl_0011,
    G124_n_spl_001
  );


  buf

  (
    G124_n_spl_01,
    G124_n_spl_0
  );


  buf

  (
    G124_n_spl_010,
    G124_n_spl_01
  );


  buf

  (
    G124_n_spl_011,
    G124_n_spl_01
  );


  buf

  (
    G124_n_spl_1,
    G124_n_spl_
  );


  buf

  (
    G124_n_spl_10,
    G124_n_spl_1
  );


  buf

  (
    G124_n_spl_100,
    G124_n_spl_10
  );


  buf

  (
    G124_n_spl_101,
    G124_n_spl_10
  );


  buf

  (
    G124_n_spl_11,
    G124_n_spl_1
  );


  buf

  (
    G124_n_spl_110,
    G124_n_spl_11
  );


  buf

  (
    G124_n_spl_111,
    G124_n_spl_11
  );


  buf

  (
    G124_p_spl_,
    G124_p
  );


  buf

  (
    G124_p_spl_0,
    G124_p_spl_
  );


  buf

  (
    G124_p_spl_00,
    G124_p_spl_0
  );


  buf

  (
    G124_p_spl_000,
    G124_p_spl_00
  );


  buf

  (
    G124_p_spl_0000,
    G124_p_spl_000
  );


  buf

  (
    G124_p_spl_0001,
    G124_p_spl_000
  );


  buf

  (
    G124_p_spl_001,
    G124_p_spl_00
  );


  buf

  (
    G124_p_spl_0010,
    G124_p_spl_001
  );


  buf

  (
    G124_p_spl_0011,
    G124_p_spl_001
  );


  buf

  (
    G124_p_spl_01,
    G124_p_spl_0
  );


  buf

  (
    G124_p_spl_010,
    G124_p_spl_01
  );


  buf

  (
    G124_p_spl_011,
    G124_p_spl_01
  );


  buf

  (
    G124_p_spl_1,
    G124_p_spl_
  );


  buf

  (
    G124_p_spl_10,
    G124_p_spl_1
  );


  buf

  (
    G124_p_spl_100,
    G124_p_spl_10
  );


  buf

  (
    G124_p_spl_101,
    G124_p_spl_10
  );


  buf

  (
    G124_p_spl_11,
    G124_p_spl_1
  );


  buf

  (
    G124_p_spl_110,
    G124_p_spl_11
  );


  buf

  (
    G124_p_spl_111,
    G124_p_spl_11
  );


  buf

  (
    g372_p_spl_,
    g372_p
  );


  buf

  (
    g372_p_spl_0,
    g372_p_spl_
  );


  buf

  (
    g372_p_spl_1,
    g372_p_spl_
  );


  buf

  (
    g372_n_spl_,
    g372_n
  );


  buf

  (
    g372_n_spl_0,
    g372_n_spl_
  );


  buf

  (
    g372_n_spl_1,
    g372_n_spl_
  );


  buf

  (
    g373_n_spl_,
    g373_n
  );


  buf

  (
    g373_n_spl_0,
    g373_n_spl_
  );


  buf

  (
    g374_n_spl_,
    g374_n
  );


  buf

  (
    g374_n_spl_0,
    g374_n_spl_
  );


  buf

  (
    g374_n_spl_1,
    g374_n_spl_
  );


  buf

  (
    g373_p_spl_,
    g373_p
  );


  buf

  (
    g373_p_spl_0,
    g373_p_spl_
  );


  buf

  (
    g374_p_spl_,
    g374_p
  );


  buf

  (
    g374_p_spl_0,
    g374_p_spl_
  );


  buf

  (
    g374_p_spl_1,
    g374_p_spl_
  );


  buf

  (
    g378_p_spl_,
    g378_p
  );


  buf

  (
    g378_p_spl_0,
    g378_p_spl_
  );


  buf

  (
    g378_p_spl_1,
    g378_p_spl_
  );


  buf

  (
    g378_n_spl_,
    g378_n
  );


  buf

  (
    g378_n_spl_0,
    g378_n_spl_
  );


  buf

  (
    g378_n_spl_1,
    g378_n_spl_
  );


  buf

  (
    g379_n_spl_,
    g379_n
  );


  buf

  (
    g380_n_spl_,
    g380_n
  );


  buf

  (
    g379_p_spl_,
    g379_p
  );


  buf

  (
    g380_p_spl_,
    g380_p
  );


  buf

  (
    g375_p_spl_,
    g375_p
  );


  buf

  (
    g375_p_spl_0,
    g375_p_spl_
  );


  buf

  (
    g375_p_spl_00,
    g375_p_spl_0
  );


  buf

  (
    g375_p_spl_1,
    g375_p_spl_
  );


  buf

  (
    g381_p_spl_,
    g381_p
  );


  buf

  (
    g381_p_spl_0,
    g381_p_spl_
  );


  buf

  (
    g381_p_spl_00,
    g381_p_spl_0
  );


  buf

  (
    g381_p_spl_01,
    g381_p_spl_0
  );


  buf

  (
    g381_p_spl_1,
    g381_p_spl_
  );


  buf

  (
    g381_p_spl_10,
    g381_p_spl_1
  );


  buf

  (
    g375_n_spl_,
    g375_n
  );


  buf

  (
    g375_n_spl_0,
    g375_n_spl_
  );


  buf

  (
    g375_n_spl_00,
    g375_n_spl_0
  );


  buf

  (
    g375_n_spl_1,
    g375_n_spl_
  );


  buf

  (
    g381_n_spl_,
    g381_n
  );


  buf

  (
    g381_n_spl_0,
    g381_n_spl_
  );


  buf

  (
    g381_n_spl_00,
    g381_n_spl_0
  );


  buf

  (
    g381_n_spl_01,
    g381_n_spl_0
  );


  buf

  (
    g381_n_spl_1,
    g381_n_spl_
  );


  buf

  (
    g381_n_spl_10,
    g381_n_spl_1
  );


  buf

  (
    g385_p_spl_,
    g385_p
  );


  buf

  (
    g385_p_spl_0,
    g385_p_spl_
  );


  buf

  (
    g385_p_spl_1,
    g385_p_spl_
  );


  buf

  (
    g385_n_spl_,
    g385_n
  );


  buf

  (
    g385_n_spl_0,
    g385_n_spl_
  );


  buf

  (
    g385_n_spl_1,
    g385_n_spl_
  );


  buf

  (
    g386_n_spl_,
    g386_n
  );


  buf

  (
    g387_n_spl_,
    g387_n
  );


  buf

  (
    g386_p_spl_,
    g386_p
  );


  buf

  (
    g387_p_spl_,
    g387_p
  );


  buf

  (
    g382_p_spl_,
    g382_p
  );


  buf

  (
    g388_p_spl_,
    g388_p
  );


  buf

  (
    g388_p_spl_0,
    g388_p_spl_
  );


  buf

  (
    g388_p_spl_00,
    g388_p_spl_0
  );


  buf

  (
    g388_p_spl_01,
    g388_p_spl_0
  );


  buf

  (
    g388_p_spl_1,
    g388_p_spl_
  );


  buf

  (
    g382_n_spl_,
    g382_n
  );


  buf

  (
    g388_n_spl_,
    g388_n
  );


  buf

  (
    g388_n_spl_0,
    g388_n_spl_
  );


  buf

  (
    g388_n_spl_00,
    g388_n_spl_0
  );


  buf

  (
    g388_n_spl_01,
    g388_n_spl_0
  );


  buf

  (
    g388_n_spl_1,
    g388_n_spl_
  );


  buf

  (
    g392_p_spl_,
    g392_p
  );


  buf

  (
    g392_p_spl_0,
    g392_p_spl_
  );


  buf

  (
    g392_p_spl_1,
    g392_p_spl_
  );


  buf

  (
    g392_n_spl_,
    g392_n
  );


  buf

  (
    g392_n_spl_0,
    g392_n_spl_
  );


  buf

  (
    g392_n_spl_1,
    g392_n_spl_
  );


  buf

  (
    g393_n_spl_,
    g393_n
  );


  buf

  (
    g389_n_spl_,
    g389_n
  );


  buf

  (
    g389_n_spl_0,
    g389_n_spl_
  );


  buf

  (
    g395_n_spl_,
    g395_n
  );


  buf

  (
    g395_n_spl_0,
    g395_n_spl_
  );


  buf

  (
    g395_n_spl_00,
    g395_n_spl_0
  );


  buf

  (
    g395_n_spl_01,
    g395_n_spl_0
  );


  buf

  (
    g395_n_spl_1,
    g395_n_spl_
  );


  buf

  (
    g395_n_spl_10,
    g395_n_spl_1
  );


  buf

  (
    g399_p_spl_,
    g399_p
  );


  buf

  (
    g399_p_spl_0,
    g399_p_spl_
  );


  buf

  (
    g399_p_spl_1,
    g399_p_spl_
  );


  buf

  (
    g399_n_spl_,
    g399_n
  );


  buf

  (
    g399_n_spl_0,
    g399_n_spl_
  );


  buf

  (
    g399_n_spl_1,
    g399_n_spl_
  );


  buf

  (
    g400_n_spl_,
    g400_n
  );


  buf

  (
    g400_n_spl_0,
    g400_n_spl_
  );


  buf

  (
    g400_n_spl_00,
    g400_n_spl_0
  );


  buf

  (
    g400_n_spl_1,
    g400_n_spl_
  );


  buf

  (
    g401_n_spl_,
    g401_n
  );


  buf

  (
    g401_n_spl_0,
    g401_n_spl_
  );


  buf

  (
    g400_p_spl_,
    g400_p
  );


  buf

  (
    g400_p_spl_0,
    g400_p_spl_
  );


  buf

  (
    g400_p_spl_00,
    g400_p_spl_0
  );


  buf

  (
    g400_p_spl_1,
    g400_p_spl_
  );


  buf

  (
    g401_p_spl_,
    g401_p
  );


  buf

  (
    g401_p_spl_0,
    g401_p_spl_
  );


  buf

  (
    g405_p_spl_,
    g405_p
  );


  buf

  (
    g405_p_spl_0,
    g405_p_spl_
  );


  buf

  (
    g405_p_spl_1,
    g405_p_spl_
  );


  buf

  (
    g405_n_spl_,
    g405_n
  );


  buf

  (
    g405_n_spl_0,
    g405_n_spl_
  );


  buf

  (
    g405_n_spl_1,
    g405_n_spl_
  );


  buf

  (
    g406_n_spl_,
    g406_n
  );


  buf

  (
    g406_n_spl_0,
    g406_n_spl_
  );


  buf

  (
    g406_p_spl_,
    g406_p
  );


  buf

  (
    g406_p_spl_0,
    g406_p_spl_
  );


  buf

  (
    g402_p_spl_,
    g402_p
  );


  buf

  (
    g402_p_spl_0,
    g402_p_spl_
  );


  buf

  (
    g402_p_spl_1,
    g402_p_spl_
  );


  buf

  (
    g408_p_spl_,
    g408_p
  );


  buf

  (
    g408_p_spl_0,
    g408_p_spl_
  );


  buf

  (
    g408_p_spl_1,
    g408_p_spl_
  );


  buf

  (
    g402_n_spl_,
    g402_n
  );


  buf

  (
    g402_n_spl_0,
    g402_n_spl_
  );


  buf

  (
    g408_n_spl_,
    g408_n
  );


  buf

  (
    g408_n_spl_0,
    g408_n_spl_
  );


  buf

  (
    g408_n_spl_00,
    g408_n_spl_0
  );


  buf

  (
    g408_n_spl_1,
    g408_n_spl_
  );


  buf

  (
    g412_p_spl_,
    g412_p
  );


  buf

  (
    g412_p_spl_0,
    g412_p_spl_
  );


  buf

  (
    g412_p_spl_1,
    g412_p_spl_
  );


  buf

  (
    g412_n_spl_,
    g412_n
  );


  buf

  (
    g412_n_spl_0,
    g412_n_spl_
  );


  buf

  (
    g412_n_spl_1,
    g412_n_spl_
  );


  buf

  (
    g413_n_spl_,
    g413_n
  );


  buf

  (
    g413_p_spl_,
    g413_p
  );


  buf

  (
    g409_p_spl_,
    g409_p
  );


  buf

  (
    g409_p_spl_0,
    g409_p_spl_
  );


  buf

  (
    g415_p_spl_,
    g415_p
  );


  buf

  (
    g415_p_spl_0,
    g415_p_spl_
  );


  buf

  (
    g415_p_spl_00,
    g415_p_spl_0
  );


  buf

  (
    g415_p_spl_1,
    g415_p_spl_
  );


  buf

  (
    g409_n_spl_,
    g409_n
  );


  buf

  (
    g409_n_spl_0,
    g409_n_spl_
  );


  buf

  (
    g415_n_spl_,
    g415_n
  );


  buf

  (
    g415_n_spl_0,
    g415_n_spl_
  );


  buf

  (
    g415_n_spl_00,
    g415_n_spl_0
  );


  buf

  (
    g415_n_spl_1,
    g415_n_spl_
  );


  buf

  (
    g419_p_spl_,
    g419_p
  );


  buf

  (
    g419_p_spl_0,
    g419_p_spl_
  );


  buf

  (
    g419_p_spl_1,
    g419_p_spl_
  );


  buf

  (
    g419_n_spl_,
    g419_n
  );


  buf

  (
    g419_n_spl_0,
    g419_n_spl_
  );


  buf

  (
    g419_n_spl_1,
    g419_n_spl_
  );


  buf

  (
    g420_n_spl_,
    g420_n
  );


  buf

  (
    g420_n_spl_0,
    g420_n_spl_
  );


  buf

  (
    g420_p_spl_,
    g420_p
  );


  buf

  (
    g420_p_spl_0,
    g420_p_spl_
  );


  buf

  (
    g416_p_spl_,
    g416_p
  );


  buf

  (
    g416_p_spl_0,
    g416_p_spl_
  );


  buf

  (
    g422_p_spl_,
    g422_p
  );


  buf

  (
    g422_p_spl_0,
    g422_p_spl_
  );


  buf

  (
    g422_p_spl_00,
    g422_p_spl_0
  );


  buf

  (
    g422_p_spl_1,
    g422_p_spl_
  );


  buf

  (
    g416_n_spl_,
    g416_n
  );


  buf

  (
    g416_n_spl_0,
    g416_n_spl_
  );


  buf

  (
    g422_n_spl_,
    g422_n
  );


  buf

  (
    g422_n_spl_0,
    g422_n_spl_
  );


  buf

  (
    g422_n_spl_00,
    g422_n_spl_0
  );


  buf

  (
    g422_n_spl_01,
    g422_n_spl_0
  );


  buf

  (
    g422_n_spl_1,
    g422_n_spl_
  );


  buf

  (
    g426_p_spl_,
    g426_p
  );


  buf

  (
    g426_p_spl_0,
    g426_p_spl_
  );


  buf

  (
    g426_p_spl_1,
    g426_p_spl_
  );


  buf

  (
    g426_n_spl_,
    g426_n
  );


  buf

  (
    g426_n_spl_0,
    g426_n_spl_
  );


  buf

  (
    g426_n_spl_1,
    g426_n_spl_
  );


  buf

  (
    g427_n_spl_,
    g427_n
  );


  buf

  (
    g427_p_spl_,
    g427_p
  );


  buf

  (
    g423_p_spl_,
    g423_p
  );


  buf

  (
    g429_p_spl_,
    g429_p
  );


  buf

  (
    g429_p_spl_0,
    g429_p_spl_
  );


  buf

  (
    g429_p_spl_00,
    g429_p_spl_0
  );


  buf

  (
    g429_p_spl_01,
    g429_p_spl_0
  );


  buf

  (
    g429_p_spl_1,
    g429_p_spl_
  );


  buf

  (
    g429_p_spl_10,
    g429_p_spl_1
  );


  buf

  (
    g423_n_spl_,
    g423_n
  );


  buf

  (
    g429_n_spl_,
    g429_n
  );


  buf

  (
    g429_n_spl_0,
    g429_n_spl_
  );


  buf

  (
    g429_n_spl_00,
    g429_n_spl_0
  );


  buf

  (
    g429_n_spl_01,
    g429_n_spl_0
  );


  buf

  (
    g429_n_spl_1,
    g429_n_spl_
  );


  buf

  (
    g429_n_spl_10,
    g429_n_spl_1
  );


  buf

  (
    g396_n_spl_,
    g396_n
  );


  buf

  (
    g430_n_spl_,
    g430_n
  );


  buf

  (
    g430_n_spl_0,
    g430_n_spl_
  );


  buf

  (
    g430_n_spl_1,
    g430_n_spl_
  );


  buf

  (
    G123_n_spl_,
    G123_n
  );


  buf

  (
    G123_n_spl_0,
    G123_n_spl_
  );


  buf

  (
    G123_n_spl_00,
    G123_n_spl_0
  );


  buf

  (
    G123_n_spl_000,
    G123_n_spl_00
  );


  buf

  (
    G123_n_spl_0000,
    G123_n_spl_000
  );


  buf

  (
    G123_n_spl_0001,
    G123_n_spl_000
  );


  buf

  (
    G123_n_spl_001,
    G123_n_spl_00
  );


  buf

  (
    G123_n_spl_0010,
    G123_n_spl_001
  );


  buf

  (
    G123_n_spl_01,
    G123_n_spl_0
  );


  buf

  (
    G123_n_spl_010,
    G123_n_spl_01
  );


  buf

  (
    G123_n_spl_011,
    G123_n_spl_01
  );


  buf

  (
    G123_n_spl_1,
    G123_n_spl_
  );


  buf

  (
    G123_n_spl_10,
    G123_n_spl_1
  );


  buf

  (
    G123_n_spl_100,
    G123_n_spl_10
  );


  buf

  (
    G123_n_spl_101,
    G123_n_spl_10
  );


  buf

  (
    G123_n_spl_11,
    G123_n_spl_1
  );


  buf

  (
    G123_n_spl_110,
    G123_n_spl_11
  );


  buf

  (
    G123_n_spl_111,
    G123_n_spl_11
  );


  buf

  (
    G123_p_spl_,
    G123_p
  );


  buf

  (
    G123_p_spl_0,
    G123_p_spl_
  );


  buf

  (
    G123_p_spl_00,
    G123_p_spl_0
  );


  buf

  (
    G123_p_spl_000,
    G123_p_spl_00
  );


  buf

  (
    G123_p_spl_0000,
    G123_p_spl_000
  );


  buf

  (
    G123_p_spl_0001,
    G123_p_spl_000
  );


  buf

  (
    G123_p_spl_001,
    G123_p_spl_00
  );


  buf

  (
    G123_p_spl_0010,
    G123_p_spl_001
  );


  buf

  (
    G123_p_spl_01,
    G123_p_spl_0
  );


  buf

  (
    G123_p_spl_010,
    G123_p_spl_01
  );


  buf

  (
    G123_p_spl_011,
    G123_p_spl_01
  );


  buf

  (
    G123_p_spl_1,
    G123_p_spl_
  );


  buf

  (
    G123_p_spl_10,
    G123_p_spl_1
  );


  buf

  (
    G123_p_spl_100,
    G123_p_spl_10
  );


  buf

  (
    G123_p_spl_101,
    G123_p_spl_10
  );


  buf

  (
    G123_p_spl_11,
    G123_p_spl_1
  );


  buf

  (
    G123_p_spl_110,
    G123_p_spl_11
  );


  buf

  (
    G123_p_spl_111,
    G123_p_spl_11
  );


  buf

  (
    g434_p_spl_,
    g434_p
  );


  buf

  (
    g434_p_spl_0,
    g434_p_spl_
  );


  buf

  (
    g434_p_spl_1,
    g434_p_spl_
  );


  buf

  (
    g434_n_spl_,
    g434_n
  );


  buf

  (
    g434_n_spl_0,
    g434_n_spl_
  );


  buf

  (
    g434_n_spl_1,
    g434_n_spl_
  );


  buf

  (
    g435_n_spl_,
    g435_n
  );


  buf

  (
    g435_p_spl_,
    g435_p
  );


  buf

  (
    g440_p_spl_,
    g440_p
  );


  buf

  (
    g440_p_spl_0,
    g440_p_spl_
  );


  buf

  (
    g440_p_spl_1,
    g440_p_spl_
  );


  buf

  (
    g440_n_spl_,
    g440_n
  );


  buf

  (
    g440_n_spl_0,
    g440_n_spl_
  );


  buf

  (
    g440_n_spl_1,
    g440_n_spl_
  );


  buf

  (
    g441_n_spl_,
    g441_n
  );


  buf

  (
    g441_n_spl_0,
    g441_n_spl_
  );


  buf

  (
    g441_n_spl_00,
    g441_n_spl_0
  );


  buf

  (
    g441_n_spl_1,
    g441_n_spl_
  );


  buf

  (
    g442_n_spl_,
    g442_n
  );


  buf

  (
    g442_n_spl_0,
    g442_n_spl_
  );


  buf

  (
    g442_n_spl_1,
    g442_n_spl_
  );


  buf

  (
    g441_p_spl_,
    g441_p
  );


  buf

  (
    g441_p_spl_0,
    g441_p_spl_
  );


  buf

  (
    g441_p_spl_00,
    g441_p_spl_0
  );


  buf

  (
    g441_p_spl_1,
    g441_p_spl_
  );


  buf

  (
    g442_p_spl_,
    g442_p
  );


  buf

  (
    g442_p_spl_0,
    g442_p_spl_
  );


  buf

  (
    g442_p_spl_1,
    g442_p_spl_
  );


  buf

  (
    g437_p_spl_,
    g437_p
  );


  buf

  (
    g437_p_spl_0,
    g437_p_spl_
  );


  buf

  (
    g437_p_spl_00,
    g437_p_spl_0
  );


  buf

  (
    g437_p_spl_01,
    g437_p_spl_0
  );


  buf

  (
    g437_p_spl_1,
    g437_p_spl_
  );


  buf

  (
    g443_p_spl_,
    g443_p
  );


  buf

  (
    g443_p_spl_0,
    g443_p_spl_
  );


  buf

  (
    g443_p_spl_00,
    g443_p_spl_0
  );


  buf

  (
    g443_p_spl_1,
    g443_p_spl_
  );


  buf

  (
    g437_n_spl_,
    g437_n
  );


  buf

  (
    g437_n_spl_0,
    g437_n_spl_
  );


  buf

  (
    g437_n_spl_00,
    g437_n_spl_0
  );


  buf

  (
    g437_n_spl_01,
    g437_n_spl_0
  );


  buf

  (
    g437_n_spl_1,
    g437_n_spl_
  );


  buf

  (
    g443_n_spl_,
    g443_n
  );


  buf

  (
    g443_n_spl_0,
    g443_n_spl_
  );


  buf

  (
    g443_n_spl_00,
    g443_n_spl_0
  );


  buf

  (
    g443_n_spl_1,
    g443_n_spl_
  );


  buf

  (
    g447_p_spl_,
    g447_p
  );


  buf

  (
    g447_p_spl_0,
    g447_p_spl_
  );


  buf

  (
    g447_p_spl_1,
    g447_p_spl_
  );


  buf

  (
    g447_n_spl_,
    g447_n
  );


  buf

  (
    g447_n_spl_0,
    g447_n_spl_
  );


  buf

  (
    g447_n_spl_1,
    g447_n_spl_
  );


  buf

  (
    g448_n_spl_,
    g448_n
  );


  buf

  (
    g448_p_spl_,
    g448_p
  );


  buf

  (
    G125_n_spl_,
    G125_n
  );


  buf

  (
    g451_n_spl_,
    g451_n
  );


  buf

  (
    g451_n_spl_0,
    g451_n_spl_
  );


  buf

  (
    g451_n_spl_1,
    g451_n_spl_
  );


  buf

  (
    g451_p_spl_,
    g451_p
  );


  buf

  (
    g451_p_spl_0,
    g451_p_spl_
  );


  buf

  (
    g451_p_spl_1,
    g451_p_spl_
  );


  buf

  (
    g452_n_spl_,
    g452_n
  );


  buf

  (
    g452_n_spl_0,
    g452_n_spl_
  );


  buf

  (
    g452_p_spl_,
    g452_p
  );


  buf

  (
    g452_p_spl_0,
    g452_p_spl_
  );


  buf

  (
    g450_p_spl_,
    g450_p
  );


  buf

  (
    g450_p_spl_0,
    g450_p_spl_
  );


  buf

  (
    g450_p_spl_1,
    g450_p_spl_
  );


  buf

  (
    g454_p_spl_,
    g454_p
  );


  buf

  (
    g454_p_spl_0,
    g454_p_spl_
  );


  buf

  (
    g454_p_spl_1,
    g454_p_spl_
  );


  buf

  (
    g450_n_spl_,
    g450_n
  );


  buf

  (
    g450_n_spl_0,
    g450_n_spl_
  );


  buf

  (
    g450_n_spl_1,
    g450_n_spl_
  );


  buf

  (
    g454_n_spl_,
    g454_n
  );


  buf

  (
    g454_n_spl_0,
    g454_n_spl_
  );


  buf

  (
    g454_n_spl_00,
    g454_n_spl_0
  );


  buf

  (
    g454_n_spl_1,
    g454_n_spl_
  );


  buf

  (
    G129_n_spl_,
    G129_n
  );


  buf

  (
    g458_p_spl_,
    g458_p
  );


  buf

  (
    g458_p_spl_0,
    g458_p_spl_
  );


  buf

  (
    g458_p_spl_1,
    g458_p_spl_
  );


  buf

  (
    g458_n_spl_,
    g458_n
  );


  buf

  (
    g458_n_spl_0,
    g458_n_spl_
  );


  buf

  (
    g458_n_spl_1,
    g458_n_spl_
  );


  buf

  (
    g459_n_spl_,
    g459_n
  );


  buf

  (
    g459_n_spl_0,
    g459_n_spl_
  );


  buf

  (
    g459_p_spl_,
    g459_p
  );


  buf

  (
    g459_p_spl_0,
    g459_p_spl_
  );


  buf

  (
    G131_n_spl_,
    G131_n
  );


  buf

  (
    g461_p_spl_,
    g461_p
  );


  buf

  (
    g461_p_spl_0,
    g461_p_spl_
  );


  buf

  (
    g464_n_spl_,
    g464_n
  );


  buf

  (
    g464_n_spl_0,
    g464_n_spl_
  );


  buf

  (
    g464_n_spl_00,
    g464_n_spl_0
  );


  buf

  (
    g464_n_spl_01,
    g464_n_spl_0
  );


  buf

  (
    g464_n_spl_1,
    g464_n_spl_
  );


  buf

  (
    g464_n_spl_10,
    g464_n_spl_1
  );


  buf

  (
    g461_n_spl_,
    g461_n
  );


  buf

  (
    g461_n_spl_0,
    g461_n_spl_
  );


  buf

  (
    g464_p_spl_,
    g464_p
  );


  buf

  (
    g464_p_spl_0,
    g464_p_spl_
  );


  buf

  (
    g464_p_spl_00,
    g464_p_spl_0
  );


  buf

  (
    g464_p_spl_01,
    g464_p_spl_0
  );


  buf

  (
    g464_p_spl_1,
    g464_p_spl_
  );


  buf

  (
    g464_p_spl_10,
    g464_p_spl_1
  );


  buf

  (
    G127_n_spl_,
    G127_n
  );


  buf

  (
    g468_p_spl_,
    g468_p
  );


  buf

  (
    g468_p_spl_0,
    g468_p_spl_
  );


  buf

  (
    g468_p_spl_1,
    g468_p_spl_
  );


  buf

  (
    g468_n_spl_,
    g468_n
  );


  buf

  (
    g468_n_spl_0,
    g468_n_spl_
  );


  buf

  (
    g468_n_spl_1,
    g468_n_spl_
  );


  buf

  (
    g469_n_spl_,
    g469_n
  );


  buf

  (
    g469_n_spl_0,
    g469_n_spl_
  );


  buf

  (
    g469_p_spl_,
    g469_p
  );


  buf

  (
    g469_p_spl_0,
    g469_p_spl_
  );


  buf

  (
    g465_p_spl_,
    g465_p
  );


  buf

  (
    g465_p_spl_0,
    g465_p_spl_
  );


  buf

  (
    g471_p_spl_,
    g471_p
  );


  buf

  (
    g471_p_spl_0,
    g471_p_spl_
  );


  buf

  (
    g471_p_spl_1,
    g471_p_spl_
  );


  buf

  (
    g465_n_spl_,
    g465_n
  );


  buf

  (
    g465_n_spl_0,
    g465_n_spl_
  );


  buf

  (
    g471_n_spl_,
    g471_n
  );


  buf

  (
    g471_n_spl_0,
    g471_n_spl_
  );


  buf

  (
    g471_n_spl_00,
    g471_n_spl_0
  );


  buf

  (
    g471_n_spl_1,
    g471_n_spl_
  );


  buf

  (
    g455_p_spl_,
    g455_p
  );


  buf

  (
    g472_p_spl_,
    g472_p
  );


  buf

  (
    g455_n_spl_,
    g455_n
  );


  buf

  (
    g472_n_spl_,
    g472_n
  );


  buf

  (
    G114_n_spl_,
    G114_n
  );


  buf

  (
    G114_n_spl_0,
    G114_n_spl_
  );


  buf

  (
    G114_p_spl_,
    G114_p
  );


  buf

  (
    g476_n_spl_,
    g476_n
  );


  buf

  (
    g476_n_spl_0,
    g476_n_spl_
  );


  buf

  (
    g476_n_spl_1,
    g476_n_spl_
  );


  buf

  (
    g479_n_spl_,
    g479_n
  );


  buf

  (
    g479_n_spl_0,
    g479_n_spl_
  );


  buf

  (
    g479_n_spl_00,
    g479_n_spl_0
  );


  buf

  (
    g479_n_spl_01,
    g479_n_spl_0
  );


  buf

  (
    g479_n_spl_1,
    g479_n_spl_
  );


  buf

  (
    g479_n_spl_10,
    g479_n_spl_1
  );


  buf

  (
    g476_p_spl_,
    g476_p
  );


  buf

  (
    g476_p_spl_0,
    g476_p_spl_
  );


  buf

  (
    g476_p_spl_00,
    g476_p_spl_0
  );


  buf

  (
    g476_p_spl_1,
    g476_p_spl_
  );


  buf

  (
    g479_p_spl_,
    g479_p
  );


  buf

  (
    g479_p_spl_0,
    g479_p_spl_
  );


  buf

  (
    g479_p_spl_00,
    g479_p_spl_0
  );


  buf

  (
    g479_p_spl_01,
    g479_p_spl_0
  );


  buf

  (
    g479_p_spl_1,
    g479_p_spl_
  );


  buf

  (
    g479_p_spl_10,
    g479_p_spl_1
  );


  buf

  (
    g473_p_spl_,
    g473_p
  );


  buf

  (
    g480_p_spl_,
    g480_p
  );


  buf

  (
    g480_p_spl_0,
    g480_p_spl_
  );


  buf

  (
    g444_p_spl_,
    g444_p
  );


  buf

  (
    g444_p_spl_0,
    g444_p_spl_
  );


  buf

  (
    g485_p_spl_,
    g485_p
  );


  buf

  (
    g488_n_spl_,
    g488_n
  );


  buf

  (
    g485_n_spl_,
    g485_n
  );


  buf

  (
    g488_p_spl_,
    g488_p
  );


  buf

  (
    G132_n_spl_,
    G132_n
  );


  buf

  (
    G132_n_spl_0,
    G132_n_spl_
  );


  buf

  (
    G132_p_spl_,
    G132_p
  );


  buf

  (
    G132_p_spl_0,
    G132_p_spl_
  );


  buf

  (
    g494_n_spl_,
    g494_n
  );


  buf

  (
    g494_p_spl_,
    g494_p
  );


  buf

  (
    g497_n_spl_,
    g497_n
  );


  buf

  (
    g500_n_spl_,
    g500_n
  );


  buf

  (
    g497_p_spl_,
    g497_p
  );


  buf

  (
    g500_p_spl_,
    g500_p
  );


  buf

  (
    g509_p_spl_,
    g509_p
  );


  buf

  (
    g512_n_spl_,
    g512_n
  );


  buf

  (
    g509_n_spl_,
    g509_n
  );


  buf

  (
    g512_p_spl_,
    g512_p
  );


  buf

  (
    G111_n_spl_,
    G111_n
  );


  buf

  (
    G111_n_spl_0,
    G111_n_spl_
  );


  buf

  (
    G111_p_spl_,
    G111_p
  );


  buf

  (
    G111_p_spl_0,
    G111_p_spl_
  );


  buf

  (
    g518_n_spl_,
    g518_n
  );


  buf

  (
    g521_n_spl_,
    g521_n
  );


  buf

  (
    g518_p_spl_,
    g518_p
  );


  buf

  (
    g521_p_spl_,
    g521_p
  );


  buf

  (
    g524_n_spl_,
    g524_n
  );


  buf

  (
    g527_n_spl_,
    g527_n
  );


  buf

  (
    g524_p_spl_,
    g524_p
  );


  buf

  (
    g527_p_spl_,
    g527_p
  );


  buf

  (
    g535_n_spl_,
    g535_n
  );


  buf

  (
    g535_n_spl_0,
    g535_n_spl_
  );


  buf

  (
    g535_n_spl_1,
    g535_n_spl_
  );


  buf

  (
    g535_p_spl_,
    g535_p
  );


  buf

  (
    g535_p_spl_0,
    g535_p_spl_
  );


  buf

  (
    g535_p_spl_1,
    g535_p_spl_
  );


  buf

  (
    g537_n_spl_,
    g537_n
  );


  buf

  (
    g537_n_spl_0,
    g537_n_spl_
  );


  buf

  (
    g537_n_spl_00,
    g537_n_spl_0
  );


  buf

  (
    g537_n_spl_1,
    g537_n_spl_
  );


  buf

  (
    g537_p_spl_,
    g537_p
  );


  buf

  (
    g537_p_spl_0,
    g537_p_spl_
  );


  buf

  (
    g537_p_spl_00,
    g537_p_spl_0
  );


  buf

  (
    g537_p_spl_1,
    g537_p_spl_
  );


  buf

  (
    g539_n_spl_,
    g539_n
  );


  buf

  (
    g539_n_spl_0,
    g539_n_spl_
  );


  buf

  (
    g539_n_spl_1,
    g539_n_spl_
  );


  buf

  (
    g539_p_spl_,
    g539_p
  );


  buf

  (
    g539_p_spl_0,
    g539_p_spl_
  );


  buf

  (
    g539_p_spl_1,
    g539_p_spl_
  );


  buf

  (
    g541_p_spl_,
    g541_p
  );


  buf

  (
    g541_p_spl_0,
    g541_p_spl_
  );


  buf

  (
    g541_p_spl_00,
    g541_p_spl_0
  );


  buf

  (
    g541_p_spl_1,
    g541_p_spl_
  );


  buf

  (
    g544_n_spl_,
    g544_n
  );


  buf

  (
    g544_n_spl_0,
    g544_n_spl_
  );


  buf

  (
    g544_n_spl_1,
    g544_n_spl_
  );


  buf

  (
    g544_p_spl_,
    g544_p
  );


  buf

  (
    g544_p_spl_0,
    g544_p_spl_
  );


  buf

  (
    g544_p_spl_1,
    g544_p_spl_
  );


  buf

  (
    g545_n_spl_,
    g545_n
  );


  buf

  (
    g545_p_spl_,
    g545_p
  );


  buf

  (
    g546_p_spl_,
    g546_p
  );


  buf

  (
    g546_p_spl_0,
    g546_p_spl_
  );


  buf

  (
    g546_p_spl_1,
    g546_p_spl_
  );


  buf

  (
    G177_p_spl_,
    G177_p
  );


  buf

  (
    G177_p_spl_0,
    G177_p_spl_
  );


  buf

  (
    G177_p_spl_00,
    G177_p_spl_0
  );


  buf

  (
    G177_p_spl_000,
    G177_p_spl_00
  );


  buf

  (
    G177_p_spl_0000,
    G177_p_spl_000
  );


  buf

  (
    G177_p_spl_0001,
    G177_p_spl_000
  );


  buf

  (
    G177_p_spl_001,
    G177_p_spl_00
  );


  buf

  (
    G177_p_spl_0010,
    G177_p_spl_001
  );


  buf

  (
    G177_p_spl_0011,
    G177_p_spl_001
  );


  buf

  (
    G177_p_spl_01,
    G177_p_spl_0
  );


  buf

  (
    G177_p_spl_010,
    G177_p_spl_01
  );


  buf

  (
    G177_p_spl_0100,
    G177_p_spl_010
  );


  buf

  (
    G177_p_spl_0101,
    G177_p_spl_010
  );


  buf

  (
    G177_p_spl_011,
    G177_p_spl_01
  );


  buf

  (
    G177_p_spl_0110,
    G177_p_spl_011
  );


  buf

  (
    G177_p_spl_0111,
    G177_p_spl_011
  );


  buf

  (
    G177_p_spl_1,
    G177_p_spl_
  );


  buf

  (
    G177_p_spl_10,
    G177_p_spl_1
  );


  buf

  (
    G177_p_spl_100,
    G177_p_spl_10
  );


  buf

  (
    G177_p_spl_1000,
    G177_p_spl_100
  );


  buf

  (
    G177_p_spl_1001,
    G177_p_spl_100
  );


  buf

  (
    G177_p_spl_101,
    G177_p_spl_10
  );


  buf

  (
    G177_p_spl_11,
    G177_p_spl_1
  );


  buf

  (
    G177_p_spl_110,
    G177_p_spl_11
  );


  buf

  (
    G177_p_spl_111,
    G177_p_spl_11
  );


  buf

  (
    g553_p_spl_,
    g553_p
  );


  buf

  (
    G176_p_spl_,
    G176_p
  );


  buf

  (
    G176_p_spl_0,
    G176_p_spl_
  );


  buf

  (
    G176_p_spl_00,
    G176_p_spl_0
  );


  buf

  (
    G176_p_spl_000,
    G176_p_spl_00
  );


  buf

  (
    G176_p_spl_0000,
    G176_p_spl_000
  );


  buf

  (
    G176_p_spl_00000,
    G176_p_spl_0000
  );


  buf

  (
    G176_p_spl_00001,
    G176_p_spl_0000
  );


  buf

  (
    G176_p_spl_0001,
    G176_p_spl_000
  );


  buf

  (
    G176_p_spl_001,
    G176_p_spl_00
  );


  buf

  (
    G176_p_spl_0010,
    G176_p_spl_001
  );


  buf

  (
    G176_p_spl_0011,
    G176_p_spl_001
  );


  buf

  (
    G176_p_spl_01,
    G176_p_spl_0
  );


  buf

  (
    G176_p_spl_010,
    G176_p_spl_01
  );


  buf

  (
    G176_p_spl_0100,
    G176_p_spl_010
  );


  buf

  (
    G176_p_spl_0101,
    G176_p_spl_010
  );


  buf

  (
    G176_p_spl_011,
    G176_p_spl_01
  );


  buf

  (
    G176_p_spl_0110,
    G176_p_spl_011
  );


  buf

  (
    G176_p_spl_0111,
    G176_p_spl_011
  );


  buf

  (
    G176_p_spl_1,
    G176_p_spl_
  );


  buf

  (
    G176_p_spl_10,
    G176_p_spl_1
  );


  buf

  (
    G176_p_spl_100,
    G176_p_spl_10
  );


  buf

  (
    G176_p_spl_1000,
    G176_p_spl_100
  );


  buf

  (
    G176_p_spl_1001,
    G176_p_spl_100
  );


  buf

  (
    G176_p_spl_101,
    G176_p_spl_10
  );


  buf

  (
    G176_p_spl_1010,
    G176_p_spl_101
  );


  buf

  (
    G176_p_spl_1011,
    G176_p_spl_101
  );


  buf

  (
    G176_p_spl_11,
    G176_p_spl_1
  );


  buf

  (
    G176_p_spl_110,
    G176_p_spl_11
  );


  buf

  (
    G176_p_spl_1100,
    G176_p_spl_110
  );


  buf

  (
    G176_p_spl_1101,
    G176_p_spl_110
  );


  buf

  (
    G176_p_spl_111,
    G176_p_spl_11
  );


  buf

  (
    G176_p_spl_1110,
    G176_p_spl_111
  );


  buf

  (
    G176_p_spl_1111,
    G176_p_spl_111
  );


  buf

  (
    G177_n_spl_,
    G177_n
  );


  buf

  (
    G177_n_spl_0,
    G177_n_spl_
  );


  buf

  (
    G177_n_spl_00,
    G177_n_spl_0
  );


  buf

  (
    G177_n_spl_000,
    G177_n_spl_00
  );


  buf

  (
    G177_n_spl_0000,
    G177_n_spl_000
  );


  buf

  (
    G177_n_spl_0001,
    G177_n_spl_000
  );


  buf

  (
    G177_n_spl_001,
    G177_n_spl_00
  );


  buf

  (
    G177_n_spl_0010,
    G177_n_spl_001
  );


  buf

  (
    G177_n_spl_0011,
    G177_n_spl_001
  );


  buf

  (
    G177_n_spl_01,
    G177_n_spl_0
  );


  buf

  (
    G177_n_spl_010,
    G177_n_spl_01
  );


  buf

  (
    G177_n_spl_011,
    G177_n_spl_01
  );


  buf

  (
    G177_n_spl_1,
    G177_n_spl_
  );


  buf

  (
    G177_n_spl_10,
    G177_n_spl_1
  );


  buf

  (
    G177_n_spl_100,
    G177_n_spl_10
  );


  buf

  (
    G177_n_spl_101,
    G177_n_spl_10
  );


  buf

  (
    G177_n_spl_11,
    G177_n_spl_1
  );


  buf

  (
    G177_n_spl_110,
    G177_n_spl_11
  );


  buf

  (
    G177_n_spl_111,
    G177_n_spl_11
  );


  buf

  (
    G176_n_spl_,
    G176_n
  );


  buf

  (
    G176_n_spl_0,
    G176_n_spl_
  );


  buf

  (
    G176_n_spl_00,
    G176_n_spl_0
  );


  buf

  (
    G176_n_spl_000,
    G176_n_spl_00
  );


  buf

  (
    G176_n_spl_0000,
    G176_n_spl_000
  );


  buf

  (
    G176_n_spl_0001,
    G176_n_spl_000
  );


  buf

  (
    G176_n_spl_001,
    G176_n_spl_00
  );


  buf

  (
    G176_n_spl_0010,
    G176_n_spl_001
  );


  buf

  (
    G176_n_spl_0011,
    G176_n_spl_001
  );


  buf

  (
    G176_n_spl_01,
    G176_n_spl_0
  );


  buf

  (
    G176_n_spl_010,
    G176_n_spl_01
  );


  buf

  (
    G176_n_spl_0100,
    G176_n_spl_010
  );


  buf

  (
    G176_n_spl_0101,
    G176_n_spl_010
  );


  buf

  (
    G176_n_spl_011,
    G176_n_spl_01
  );


  buf

  (
    G176_n_spl_1,
    G176_n_spl_
  );


  buf

  (
    G176_n_spl_10,
    G176_n_spl_1
  );


  buf

  (
    G176_n_spl_100,
    G176_n_spl_10
  );


  buf

  (
    G176_n_spl_101,
    G176_n_spl_10
  );


  buf

  (
    G176_n_spl_11,
    G176_n_spl_1
  );


  buf

  (
    G176_n_spl_110,
    G176_n_spl_11
  );


  buf

  (
    G176_n_spl_111,
    G176_n_spl_11
  );


  buf

  (
    g562_n_spl_,
    g562_n
  );


  buf

  (
    g562_n_spl_0,
    g562_n_spl_
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G2_p_spl_0,
    G2_p_spl_
  );


  buf

  (
    G2_p_spl_1,
    G2_p_spl_
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G2_n_spl_0,
    G2_n_spl_
  );


  buf

  (
    g570_n_spl_,
    g570_n
  );


  buf

  (
    g572_p_spl_,
    g572_p
  );


  buf

  (
    G22_p_spl_,
    G22_p
  );


  buf

  (
    G173_n_spl_,
    G173_n
  );


  buf

  (
    G173_n_spl_0,
    G173_n_spl_
  );


  buf

  (
    G173_n_spl_00,
    G173_n_spl_0
  );


  buf

  (
    G173_n_spl_000,
    G173_n_spl_00
  );


  buf

  (
    G173_n_spl_0000,
    G173_n_spl_000
  );


  buf

  (
    G173_n_spl_0001,
    G173_n_spl_000
  );


  buf

  (
    G173_n_spl_001,
    G173_n_spl_00
  );


  buf

  (
    G173_n_spl_0010,
    G173_n_spl_001
  );


  buf

  (
    G173_n_spl_0011,
    G173_n_spl_001
  );


  buf

  (
    G173_n_spl_01,
    G173_n_spl_0
  );


  buf

  (
    G173_n_spl_010,
    G173_n_spl_01
  );


  buf

  (
    G173_n_spl_011,
    G173_n_spl_01
  );


  buf

  (
    G173_n_spl_1,
    G173_n_spl_
  );


  buf

  (
    G173_n_spl_10,
    G173_n_spl_1
  );


  buf

  (
    G173_n_spl_100,
    G173_n_spl_10
  );


  buf

  (
    G173_n_spl_101,
    G173_n_spl_10
  );


  buf

  (
    G173_n_spl_11,
    G173_n_spl_1
  );


  buf

  (
    G173_n_spl_110,
    G173_n_spl_11
  );


  buf

  (
    G173_n_spl_111,
    G173_n_spl_11
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G173_p_spl_,
    G173_p
  );


  buf

  (
    G173_p_spl_0,
    G173_p_spl_
  );


  buf

  (
    G173_p_spl_00,
    G173_p_spl_0
  );


  buf

  (
    G173_p_spl_000,
    G173_p_spl_00
  );


  buf

  (
    G173_p_spl_0000,
    G173_p_spl_000
  );


  buf

  (
    G173_p_spl_0001,
    G173_p_spl_000
  );


  buf

  (
    G173_p_spl_001,
    G173_p_spl_00
  );


  buf

  (
    G173_p_spl_0010,
    G173_p_spl_001
  );


  buf

  (
    G173_p_spl_0011,
    G173_p_spl_001
  );


  buf

  (
    G173_p_spl_01,
    G173_p_spl_0
  );


  buf

  (
    G173_p_spl_010,
    G173_p_spl_01
  );


  buf

  (
    G173_p_spl_011,
    G173_p_spl_01
  );


  buf

  (
    G173_p_spl_1,
    G173_p_spl_
  );


  buf

  (
    G173_p_spl_10,
    G173_p_spl_1
  );


  buf

  (
    G173_p_spl_100,
    G173_p_spl_10
  );


  buf

  (
    G173_p_spl_101,
    G173_p_spl_10
  );


  buf

  (
    G173_p_spl_11,
    G173_p_spl_1
  );


  buf

  (
    G173_p_spl_110,
    G173_p_spl_11
  );


  buf

  (
    G173_p_spl_111,
    G173_p_spl_11
  );


  buf

  (
    G172_n_spl_,
    G172_n
  );


  buf

  (
    G172_n_spl_0,
    G172_n_spl_
  );


  buf

  (
    G172_n_spl_00,
    G172_n_spl_0
  );


  buf

  (
    G172_n_spl_000,
    G172_n_spl_00
  );


  buf

  (
    G172_n_spl_001,
    G172_n_spl_00
  );


  buf

  (
    G172_n_spl_01,
    G172_n_spl_0
  );


  buf

  (
    G172_n_spl_1,
    G172_n_spl_
  );


  buf

  (
    G172_n_spl_10,
    G172_n_spl_1
  );


  buf

  (
    G172_n_spl_11,
    G172_n_spl_1
  );


  buf

  (
    g579_p_spl_,
    g579_p
  );


  buf

  (
    g579_p_spl_0,
    g579_p_spl_
  );


  buf

  (
    g579_p_spl_00,
    g579_p_spl_0
  );


  buf

  (
    g579_p_spl_1,
    g579_p_spl_
  );


  buf

  (
    g560_p_spl_,
    g560_p
  );


  buf

  (
    g560_p_spl_0,
    g560_p_spl_
  );


  buf

  (
    g560_p_spl_00,
    g560_p_spl_0
  );


  buf

  (
    g560_p_spl_1,
    g560_p_spl_
  );


  buf

  (
    G172_p_spl_,
    G172_p
  );


  buf

  (
    G172_p_spl_0,
    G172_p_spl_
  );


  buf

  (
    G172_p_spl_00,
    G172_p_spl_0
  );


  buf

  (
    G172_p_spl_000,
    G172_p_spl_00
  );


  buf

  (
    G172_p_spl_001,
    G172_p_spl_00
  );


  buf

  (
    G172_p_spl_01,
    G172_p_spl_0
  );


  buf

  (
    G172_p_spl_1,
    G172_p_spl_
  );


  buf

  (
    G172_p_spl_10,
    G172_p_spl_1
  );


  buf

  (
    G172_p_spl_11,
    G172_p_spl_1
  );


  buf

  (
    g594_n_spl_,
    g594_n
  );


  buf

  (
    g594_p_spl_,
    g594_p
  );


  buf

  (
    g595_n_spl_,
    g595_n
  );


  buf

  (
    g596_n_spl_,
    g596_n
  );


  buf

  (
    g596_n_spl_0,
    g596_n_spl_
  );


  buf

  (
    g596_p_spl_,
    g596_p
  );


  buf

  (
    g596_p_spl_0,
    g596_p_spl_
  );


  buf

  (
    g596_p_spl_1,
    g596_p_spl_
  );


  buf

  (
    g597_p_spl_,
    g597_p
  );


  buf

  (
    g598_p_spl_,
    g598_p
  );


  buf

  (
    g598_p_spl_0,
    g598_p_spl_
  );


  buf

  (
    g598_n_spl_,
    g598_n
  );


  buf

  (
    g598_n_spl_0,
    g598_n_spl_
  );


  buf

  (
    g601_p_spl_,
    g601_p
  );


  buf

  (
    g610_n_spl_,
    g610_n
  );


  buf

  (
    g617_p_spl_,
    g617_p
  );


  buf

  (
    g617_p_spl_0,
    g617_p_spl_
  );


  buf

  (
    g619_n_spl_,
    g619_n
  );


  buf

  (
    G174_n_spl_,
    G174_n
  );


  buf

  (
    G174_n_spl_0,
    G174_n_spl_
  );


  buf

  (
    G174_n_spl_00,
    G174_n_spl_0
  );


  buf

  (
    G174_n_spl_000,
    G174_n_spl_00
  );


  buf

  (
    G174_n_spl_0000,
    G174_n_spl_000
  );


  buf

  (
    G174_n_spl_0001,
    G174_n_spl_000
  );


  buf

  (
    G174_n_spl_001,
    G174_n_spl_00
  );


  buf

  (
    G174_n_spl_0010,
    G174_n_spl_001
  );


  buf

  (
    G174_n_spl_0011,
    G174_n_spl_001
  );


  buf

  (
    G174_n_spl_01,
    G174_n_spl_0
  );


  buf

  (
    G174_n_spl_010,
    G174_n_spl_01
  );


  buf

  (
    G174_n_spl_011,
    G174_n_spl_01
  );


  buf

  (
    G174_n_spl_1,
    G174_n_spl_
  );


  buf

  (
    G174_n_spl_10,
    G174_n_spl_1
  );


  buf

  (
    G174_n_spl_100,
    G174_n_spl_10
  );


  buf

  (
    G174_n_spl_101,
    G174_n_spl_10
  );


  buf

  (
    G174_n_spl_11,
    G174_n_spl_1
  );


  buf

  (
    G174_n_spl_110,
    G174_n_spl_11
  );


  buf

  (
    G174_n_spl_111,
    G174_n_spl_11
  );


  buf

  (
    G174_p_spl_,
    G174_p
  );


  buf

  (
    G174_p_spl_0,
    G174_p_spl_
  );


  buf

  (
    G174_p_spl_00,
    G174_p_spl_0
  );


  buf

  (
    G174_p_spl_000,
    G174_p_spl_00
  );


  buf

  (
    G174_p_spl_0000,
    G174_p_spl_000
  );


  buf

  (
    G174_p_spl_0001,
    G174_p_spl_000
  );


  buf

  (
    G174_p_spl_001,
    G174_p_spl_00
  );


  buf

  (
    G174_p_spl_0010,
    G174_p_spl_001
  );


  buf

  (
    G174_p_spl_0011,
    G174_p_spl_001
  );


  buf

  (
    G174_p_spl_01,
    G174_p_spl_0
  );


  buf

  (
    G174_p_spl_010,
    G174_p_spl_01
  );


  buf

  (
    G174_p_spl_011,
    G174_p_spl_01
  );


  buf

  (
    G174_p_spl_1,
    G174_p_spl_
  );


  buf

  (
    G174_p_spl_10,
    G174_p_spl_1
  );


  buf

  (
    G174_p_spl_100,
    G174_p_spl_10
  );


  buf

  (
    G174_p_spl_101,
    G174_p_spl_10
  );


  buf

  (
    G174_p_spl_11,
    G174_p_spl_1
  );


  buf

  (
    G174_p_spl_110,
    G174_p_spl_11
  );


  buf

  (
    G174_p_spl_111,
    G174_p_spl_11
  );


  buf

  (
    G175_n_spl_,
    G175_n
  );


  buf

  (
    G175_n_spl_0,
    G175_n_spl_
  );


  buf

  (
    G175_n_spl_00,
    G175_n_spl_0
  );


  buf

  (
    G175_n_spl_000,
    G175_n_spl_00
  );


  buf

  (
    G175_n_spl_001,
    G175_n_spl_00
  );


  buf

  (
    G175_n_spl_01,
    G175_n_spl_0
  );


  buf

  (
    G175_n_spl_1,
    G175_n_spl_
  );


  buf

  (
    G175_n_spl_10,
    G175_n_spl_1
  );


  buf

  (
    G175_n_spl_11,
    G175_n_spl_1
  );


  buf

  (
    G175_p_spl_,
    G175_p
  );


  buf

  (
    G175_p_spl_0,
    G175_p_spl_
  );


  buf

  (
    G175_p_spl_00,
    G175_p_spl_0
  );


  buf

  (
    G175_p_spl_000,
    G175_p_spl_00
  );


  buf

  (
    G175_p_spl_001,
    G175_p_spl_00
  );


  buf

  (
    G175_p_spl_01,
    G175_p_spl_0
  );


  buf

  (
    G175_p_spl_1,
    G175_p_spl_
  );


  buf

  (
    G175_p_spl_10,
    G175_p_spl_1
  );


  buf

  (
    G175_p_spl_11,
    G175_p_spl_1
  );


  buf

  (
    g638_p_spl_,
    g638_p
  );


  buf

  (
    g639_p_spl_,
    g639_p
  );


  buf

  (
    g643_n_spl_,
    g643_n
  );


  buf

  (
    g652_n_spl_,
    g652_n
  );


  buf

  (
    g659_p_spl_,
    g659_p
  );


  buf

  (
    g660_p_spl_,
    g660_p
  );


  buf

  (
    g664_n_spl_,
    g664_n
  );


  buf

  (
    g673_n_spl_,
    g673_n
  );


  buf

  (
    g581_n_spl_,
    g581_n
  );


  buf

  (
    g581_n_spl_0,
    g581_n_spl_
  );


  buf

  (
    g581_n_spl_00,
    g581_n_spl_0
  );


  buf

  (
    g581_n_spl_01,
    g581_n_spl_0
  );


  buf

  (
    g581_n_spl_1,
    g581_n_spl_
  );


  buf

  (
    g581_n_spl_10,
    g581_n_spl_1
  );


  buf

  (
    g581_n_spl_11,
    g581_n_spl_1
  );


  buf

  (
    g681_p_spl_,
    g681_p
  );


  buf

  (
    g581_p_spl_,
    g581_p
  );


  buf

  (
    g581_p_spl_0,
    g581_p_spl_
  );


  buf

  (
    g581_p_spl_00,
    g581_p_spl_0
  );


  buf

  (
    g581_p_spl_01,
    g581_p_spl_0
  );


  buf

  (
    g581_p_spl_1,
    g581_p_spl_
  );


  buf

  (
    g681_n_spl_,
    g681_n
  );


  buf

  (
    g687_n_spl_,
    g687_n
  );


  buf

  (
    g687_p_spl_,
    g687_p
  );


  buf

  (
    g693_n_spl_,
    g693_n
  );


  buf

  (
    g696_n_spl_,
    g696_n
  );


  buf

  (
    g693_p_spl_,
    g693_p
  );


  buf

  (
    g696_p_spl_,
    g696_p
  );


  buf

  (
    g690_p_spl_,
    g690_p
  );


  buf

  (
    g699_n_spl_,
    g699_n
  );


  buf

  (
    g690_n_spl_,
    g690_n
  );


  buf

  (
    g699_p_spl_,
    g699_p
  );


  buf

  (
    g708_p_spl_,
    g708_p
  );


  buf

  (
    g711_n_spl_,
    g711_n
  );


  buf

  (
    g708_n_spl_,
    g708_n
  );


  buf

  (
    g711_p_spl_,
    g711_p
  );


  buf

  (
    g717_n_spl_,
    g717_n
  );


  buf

  (
    g717_p_spl_,
    g717_p
  );


  buf

  (
    g720_p_spl_,
    g720_p
  );


  buf

  (
    g723_n_spl_,
    g723_n
  );


  buf

  (
    g720_n_spl_,
    g720_n
  );


  buf

  (
    g723_p_spl_,
    g723_p
  );


  buf

  (
    g726_n_spl_,
    g726_n
  );


  buf

  (
    g729_n_spl_,
    g729_n
  );


  buf

  (
    g726_p_spl_,
    g726_p
  );


  buf

  (
    g729_p_spl_,
    g729_p
  );


  buf

  (
    g430_p_spl_,
    g430_p
  );


  buf

  (
    g430_p_spl_0,
    g430_p_spl_
  );


  buf

  (
    g541_n_spl_,
    g541_n
  );


  buf

  (
    g541_n_spl_0,
    g541_n_spl_
  );


  buf

  (
    g541_n_spl_1,
    g541_n_spl_
  );


  buf

  (
    g737_p_spl_,
    g737_p
  );


  buf

  (
    g737_p_spl_0,
    g737_p_spl_
  );


  buf

  (
    g737_p_spl_00,
    g737_p_spl_0
  );


  buf

  (
    g737_p_spl_1,
    g737_p_spl_
  );


  buf

  (
    g737_n_spl_,
    g737_n
  );


  buf

  (
    g737_n_spl_0,
    g737_n_spl_
  );


  buf

  (
    g737_n_spl_00,
    g737_n_spl_0
  );


  buf

  (
    g737_n_spl_1,
    g737_n_spl_
  );


  buf

  (
    g743_p_spl_,
    g743_p
  );


  buf

  (
    g747_p_spl_,
    g747_p
  );


  buf

  (
    g389_p_spl_,
    g389_p
  );


  buf

  (
    g546_n_spl_,
    g546_n
  );


  buf

  (
    g546_n_spl_0,
    g546_n_spl_
  );


  buf

  (
    g395_p_spl_,
    g395_p
  );


  buf

  (
    g395_p_spl_0,
    g395_p_spl_
  );


  buf

  (
    g395_p_spl_00,
    g395_p_spl_0
  );


  buf

  (
    g395_p_spl_1,
    g395_p_spl_
  );


  buf

  (
    g755_p_spl_,
    g755_p
  );


  buf

  (
    g760_p_spl_,
    g760_p
  );


  buf

  (
    g774_p_spl_,
    g774_p
  );


  buf

  (
    g774_p_spl_0,
    g774_p_spl_
  );


  buf

  (
    g774_p_spl_00,
    g774_p_spl_0
  );


  buf

  (
    g774_p_spl_01,
    g774_p_spl_0
  );


  buf

  (
    g774_p_spl_1,
    g774_p_spl_
  );


  buf

  (
    g774_n_spl_,
    g774_n
  );


  buf

  (
    g774_n_spl_0,
    g774_n_spl_
  );


  buf

  (
    g774_n_spl_00,
    g774_n_spl_0
  );


  buf

  (
    g774_n_spl_01,
    g774_n_spl_0
  );


  buf

  (
    g774_n_spl_1,
    g774_n_spl_
  );


  buf

  (
    g777_p_spl_,
    g777_p
  );


  buf

  (
    g444_n_spl_,
    g444_n
  );


  buf

  (
    g780_p_spl_,
    g780_p
  );


  buf

  (
    g780_p_spl_0,
    g780_p_spl_
  );


  buf

  (
    g780_p_spl_1,
    g780_p_spl_
  );


  buf

  (
    g780_n_spl_,
    g780_n
  );


  buf

  (
    g780_n_spl_0,
    g780_n_spl_
  );


  buf

  (
    g780_n_spl_1,
    g780_n_spl_
  );


  buf

  (
    g785_p_spl_,
    g785_p
  );


  buf

  (
    g791_p_spl_,
    g791_p
  );


  buf

  (
    G81_p_spl_,
    G81_p
  );


  buf

  (
    G158_n_spl_,
    G158_n
  );


  buf

  (
    G158_n_spl_0,
    G158_n_spl_
  );


  buf

  (
    G158_n_spl_00,
    G158_n_spl_0
  );


  buf

  (
    G158_n_spl_000,
    G158_n_spl_00
  );


  buf

  (
    G158_n_spl_0000,
    G158_n_spl_000
  );


  buf

  (
    G158_n_spl_0001,
    G158_n_spl_000
  );


  buf

  (
    G158_n_spl_001,
    G158_n_spl_00
  );


  buf

  (
    G158_n_spl_0010,
    G158_n_spl_001
  );


  buf

  (
    G158_n_spl_0011,
    G158_n_spl_001
  );


  buf

  (
    G158_n_spl_01,
    G158_n_spl_0
  );


  buf

  (
    G158_n_spl_010,
    G158_n_spl_01
  );


  buf

  (
    G158_n_spl_011,
    G158_n_spl_01
  );


  buf

  (
    G158_n_spl_1,
    G158_n_spl_
  );


  buf

  (
    G158_n_spl_10,
    G158_n_spl_1
  );


  buf

  (
    G158_n_spl_100,
    G158_n_spl_10
  );


  buf

  (
    G158_n_spl_101,
    G158_n_spl_10
  );


  buf

  (
    G158_n_spl_11,
    G158_n_spl_1
  );


  buf

  (
    G158_n_spl_110,
    G158_n_spl_11
  );


  buf

  (
    G158_n_spl_111,
    G158_n_spl_11
  );


  buf

  (
    G80_p_spl_,
    G80_p
  );


  buf

  (
    G158_p_spl_,
    G158_p
  );


  buf

  (
    G158_p_spl_0,
    G158_p_spl_
  );


  buf

  (
    G158_p_spl_00,
    G158_p_spl_0
  );


  buf

  (
    G158_p_spl_000,
    G158_p_spl_00
  );


  buf

  (
    G158_p_spl_0000,
    G158_p_spl_000
  );


  buf

  (
    G158_p_spl_0001,
    G158_p_spl_000
  );


  buf

  (
    G158_p_spl_001,
    G158_p_spl_00
  );


  buf

  (
    G158_p_spl_0010,
    G158_p_spl_001
  );


  buf

  (
    G158_p_spl_0011,
    G158_p_spl_001
  );


  buf

  (
    G158_p_spl_01,
    G158_p_spl_0
  );


  buf

  (
    G158_p_spl_010,
    G158_p_spl_01
  );


  buf

  (
    G158_p_spl_011,
    G158_p_spl_01
  );


  buf

  (
    G158_p_spl_1,
    G158_p_spl_
  );


  buf

  (
    G158_p_spl_10,
    G158_p_spl_1
  );


  buf

  (
    G158_p_spl_100,
    G158_p_spl_10
  );


  buf

  (
    G158_p_spl_101,
    G158_p_spl_10
  );


  buf

  (
    G158_p_spl_11,
    G158_p_spl_1
  );


  buf

  (
    G158_p_spl_110,
    G158_p_spl_11
  );


  buf

  (
    G158_p_spl_111,
    G158_p_spl_11
  );


  buf

  (
    G159_n_spl_,
    G159_n
  );


  buf

  (
    G159_n_spl_0,
    G159_n_spl_
  );


  buf

  (
    G159_n_spl_00,
    G159_n_spl_0
  );


  buf

  (
    G159_n_spl_000,
    G159_n_spl_00
  );


  buf

  (
    G159_n_spl_001,
    G159_n_spl_00
  );


  buf

  (
    G159_n_spl_01,
    G159_n_spl_0
  );


  buf

  (
    G159_n_spl_1,
    G159_n_spl_
  );


  buf

  (
    G159_n_spl_10,
    G159_n_spl_1
  );


  buf

  (
    G159_n_spl_11,
    G159_n_spl_1
  );


  buf

  (
    G159_p_spl_,
    G159_p
  );


  buf

  (
    G159_p_spl_0,
    G159_p_spl_
  );


  buf

  (
    G159_p_spl_00,
    G159_p_spl_0
  );


  buf

  (
    G159_p_spl_000,
    G159_p_spl_00
  );


  buf

  (
    G159_p_spl_001,
    G159_p_spl_00
  );


  buf

  (
    G159_p_spl_01,
    G159_p_spl_0
  );


  buf

  (
    G159_p_spl_1,
    G159_p_spl_
  );


  buf

  (
    G159_p_spl_10,
    G159_p_spl_1
  );


  buf

  (
    G159_p_spl_11,
    G159_p_spl_1
  );


  buf

  (
    G64_p_spl_,
    G64_p
  );


  buf

  (
    G64_p_spl_0,
    G64_p_spl_
  );


  buf

  (
    G64_p_spl_00,
    G64_p_spl_0
  );


  buf

  (
    G64_p_spl_000,
    G64_p_spl_00
  );


  buf

  (
    G64_p_spl_0000,
    G64_p_spl_000
  );


  buf

  (
    G64_p_spl_0001,
    G64_p_spl_000
  );


  buf

  (
    G64_p_spl_001,
    G64_p_spl_00
  );


  buf

  (
    G64_p_spl_0010,
    G64_p_spl_001
  );


  buf

  (
    G64_p_spl_01,
    G64_p_spl_0
  );


  buf

  (
    G64_p_spl_010,
    G64_p_spl_01
  );


  buf

  (
    G64_p_spl_011,
    G64_p_spl_01
  );


  buf

  (
    G64_p_spl_1,
    G64_p_spl_
  );


  buf

  (
    G64_p_spl_10,
    G64_p_spl_1
  );


  buf

  (
    G64_p_spl_100,
    G64_p_spl_10
  );


  buf

  (
    G64_p_spl_101,
    G64_p_spl_10
  );


  buf

  (
    G64_p_spl_11,
    G64_p_spl_1
  );


  buf

  (
    G64_p_spl_110,
    G64_p_spl_11
  );


  buf

  (
    G64_p_spl_111,
    G64_p_spl_11
  );


  buf

  (
    G160_n_spl_,
    G160_n
  );


  buf

  (
    G160_n_spl_0,
    G160_n_spl_
  );


  buf

  (
    G160_n_spl_00,
    G160_n_spl_0
  );


  buf

  (
    G160_n_spl_000,
    G160_n_spl_00
  );


  buf

  (
    G160_n_spl_0000,
    G160_n_spl_000
  );


  buf

  (
    G160_n_spl_0001,
    G160_n_spl_000
  );


  buf

  (
    G160_n_spl_001,
    G160_n_spl_00
  );


  buf

  (
    G160_n_spl_0010,
    G160_n_spl_001
  );


  buf

  (
    G160_n_spl_0011,
    G160_n_spl_001
  );


  buf

  (
    G160_n_spl_01,
    G160_n_spl_0
  );


  buf

  (
    G160_n_spl_010,
    G160_n_spl_01
  );


  buf

  (
    G160_n_spl_011,
    G160_n_spl_01
  );


  buf

  (
    G160_n_spl_1,
    G160_n_spl_
  );


  buf

  (
    G160_n_spl_10,
    G160_n_spl_1
  );


  buf

  (
    G160_n_spl_100,
    G160_n_spl_10
  );


  buf

  (
    G160_n_spl_101,
    G160_n_spl_10
  );


  buf

  (
    G160_n_spl_11,
    G160_n_spl_1
  );


  buf

  (
    G160_n_spl_110,
    G160_n_spl_11
  );


  buf

  (
    G160_n_spl_111,
    G160_n_spl_11
  );


  buf

  (
    G160_p_spl_,
    G160_p
  );


  buf

  (
    G160_p_spl_0,
    G160_p_spl_
  );


  buf

  (
    G160_p_spl_00,
    G160_p_spl_0
  );


  buf

  (
    G160_p_spl_000,
    G160_p_spl_00
  );


  buf

  (
    G160_p_spl_0000,
    G160_p_spl_000
  );


  buf

  (
    G160_p_spl_0001,
    G160_p_spl_000
  );


  buf

  (
    G160_p_spl_001,
    G160_p_spl_00
  );


  buf

  (
    G160_p_spl_0010,
    G160_p_spl_001
  );


  buf

  (
    G160_p_spl_0011,
    G160_p_spl_001
  );


  buf

  (
    G160_p_spl_01,
    G160_p_spl_0
  );


  buf

  (
    G160_p_spl_010,
    G160_p_spl_01
  );


  buf

  (
    G160_p_spl_011,
    G160_p_spl_01
  );


  buf

  (
    G160_p_spl_1,
    G160_p_spl_
  );


  buf

  (
    G160_p_spl_10,
    G160_p_spl_1
  );


  buf

  (
    G160_p_spl_100,
    G160_p_spl_10
  );


  buf

  (
    G160_p_spl_101,
    G160_p_spl_10
  );


  buf

  (
    G160_p_spl_11,
    G160_p_spl_1
  );


  buf

  (
    G160_p_spl_110,
    G160_p_spl_11
  );


  buf

  (
    G160_p_spl_111,
    G160_p_spl_11
  );


  buf

  (
    G161_n_spl_,
    G161_n
  );


  buf

  (
    G161_n_spl_0,
    G161_n_spl_
  );


  buf

  (
    G161_n_spl_00,
    G161_n_spl_0
  );


  buf

  (
    G161_n_spl_000,
    G161_n_spl_00
  );


  buf

  (
    G161_n_spl_001,
    G161_n_spl_00
  );


  buf

  (
    G161_n_spl_01,
    G161_n_spl_0
  );


  buf

  (
    G161_n_spl_1,
    G161_n_spl_
  );


  buf

  (
    G161_n_spl_10,
    G161_n_spl_1
  );


  buf

  (
    G161_n_spl_11,
    G161_n_spl_1
  );


  buf

  (
    G161_p_spl_,
    G161_p
  );


  buf

  (
    G161_p_spl_0,
    G161_p_spl_
  );


  buf

  (
    G161_p_spl_00,
    G161_p_spl_0
  );


  buf

  (
    G161_p_spl_000,
    G161_p_spl_00
  );


  buf

  (
    G161_p_spl_001,
    G161_p_spl_00
  );


  buf

  (
    G161_p_spl_01,
    G161_p_spl_0
  );


  buf

  (
    G161_p_spl_1,
    G161_p_spl_
  );


  buf

  (
    G161_p_spl_10,
    G161_p_spl_1
  );


  buf

  (
    G161_p_spl_11,
    G161_p_spl_1
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    g647_n_spl_,
    g647_n
  );


  buf

  (
    g647_n_spl_0,
    g647_n_spl_
  );


  buf

  (
    g647_n_spl_00,
    g647_n_spl_0
  );


  buf

  (
    g647_n_spl_1,
    g647_n_spl_
  );


  buf

  (
    g605_n_spl_,
    g605_n
  );


  buf

  (
    g605_n_spl_0,
    g605_n_spl_
  );


  buf

  (
    g605_n_spl_00,
    g605_n_spl_0
  );


  buf

  (
    g605_n_spl_1,
    g605_n_spl_
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G27_p_spl_,
    G27_p
  );


  buf

  (
    g656_n_spl_,
    g656_n
  );


  buf

  (
    g656_n_spl_0,
    g656_n_spl_
  );


  buf

  (
    g656_n_spl_00,
    g656_n_spl_0
  );


  buf

  (
    g656_n_spl_1,
    g656_n_spl_
  );


  buf

  (
    g614_n_spl_,
    g614_n
  );


  buf

  (
    g614_n_spl_0,
    g614_n_spl_
  );


  buf

  (
    g614_n_spl_00,
    g614_n_spl_0
  );


  buf

  (
    g614_n_spl_1,
    g614_n_spl_
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G26_p_spl_,
    G26_p
  );


  buf

  (
    g669_n_spl_,
    g669_n
  );


  buf

  (
    g669_n_spl_0,
    g669_n_spl_
  );


  buf

  (
    g669_n_spl_00,
    g669_n_spl_0
  );


  buf

  (
    g669_n_spl_1,
    g669_n_spl_
  );


  buf

  (
    g624_n_spl_,
    g624_n
  );


  buf

  (
    g624_n_spl_0,
    g624_n_spl_
  );


  buf

  (
    g624_n_spl_00,
    g624_n_spl_0
  );


  buf

  (
    g624_n_spl_1,
    g624_n_spl_
  );


  buf

  (
    G25_p_spl_,
    G25_p
  );


  buf

  (
    G24_p_spl_,
    G24_p
  );


  buf

  (
    g678_n_spl_,
    g678_n
  );


  buf

  (
    g678_n_spl_0,
    g678_n_spl_
  );


  buf

  (
    g678_n_spl_00,
    g678_n_spl_0
  );


  buf

  (
    g678_n_spl_1,
    g678_n_spl_
  );


  buf

  (
    g569_p_spl_,
    g569_p
  );


  buf

  (
    g569_p_spl_0,
    g569_p_spl_
  );


  buf

  (
    g569_p_spl_00,
    g569_p_spl_0
  );


  buf

  (
    g569_p_spl_1,
    g569_p_spl_
  );


  buf

  (
    G76_p_spl_,
    G76_p
  );


  buf

  (
    G86_p_spl_,
    G86_p
  );


  buf

  (
    G72_p_spl_,
    G72_p
  );


  buf

  (
    G82_p_spl_,
    G82_p
  );


  buf

  (
    G70_p_spl_,
    G70_p
  );


  buf

  (
    G71_p_spl_,
    G71_p
  );


  buf

  (
    G68_p_spl_,
    G68_p
  );


  buf

  (
    G69_p_spl_,
    G69_p
  );


  buf

  (
    G171_p_spl_,
    G171_p
  );


  buf

  (
    G54_p_spl_,
    G54_p
  );


  buf

  (
    G171_n_spl_,
    G171_n
  );


  buf

  (
    G61_n_spl_,
    G61_n
  );


  buf

  (
    G61_p_spl_,
    G61_p
  );


  buf

  (
    g975_p_spl_,
    g975_p
  );


  buf

  (
    G99_n_spl_,
    G99_n
  );


  buf

  (
    g533_n_spl_,
    g533_n
  );


  buf

  (
    g735_n_spl_,
    g735_n
  );


  buf

  (
    G155_n_spl_,
    G155_n
  );


  buf

  (
    g184_n_spl_,
    g184_n
  );


  buf

  (
    g179_n_spl_,
    g179_n
  );


  buf

  (
    g705_n_spl_,
    g705_n
  );


  buf

  (
    g506_n_spl_,
    g506_n
  );


  buf

  (
    g1025_n_spl_,
    g1025_n
  );


  buf

  (
    g1025_n_spl_0,
    g1025_n_spl_
  );


  buf

  (
    g1025_n_spl_00,
    g1025_n_spl_0
  );


  buf

  (
    g1025_n_spl_1,
    g1025_n_spl_
  );


  buf

  (
    g990_p_spl_,
    g990_p
  );


  buf

  (
    g990_p_spl_0,
    g990_p_spl_
  );


  buf

  (
    g990_p_spl_00,
    g990_p_spl_0
  );


  buf

  (
    g990_p_spl_1,
    g990_p_spl_
  );


  buf

  (
    G41_p_spl_,
    G41_p
  );


  buf

  (
    G42_p_spl_,
    G42_p
  );


  buf

  (
    G18_p_spl_,
    G18_p
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    g1032_n_spl_,
    g1032_n
  );


  buf

  (
    g1032_n_spl_0,
    g1032_n_spl_
  );


  buf

  (
    g1032_n_spl_00,
    g1032_n_spl_0
  );


  buf

  (
    g1032_n_spl_1,
    g1032_n_spl_
  );


  buf

  (
    g997_n_spl_,
    g997_n
  );


  buf

  (
    g997_n_spl_0,
    g997_n_spl_
  );


  buf

  (
    g997_n_spl_00,
    g997_n_spl_0
  );


  buf

  (
    g997_n_spl_1,
    g997_n_spl_
  );


  buf

  (
    G40_p_spl_,
    G40_p
  );


  buf

  (
    G39_p_spl_,
    G39_p
  );


  buf

  (
    g1039_n_spl_,
    g1039_n
  );


  buf

  (
    g1039_n_spl_0,
    g1039_n_spl_
  );


  buf

  (
    g1039_n_spl_00,
    g1039_n_spl_0
  );


  buf

  (
    g1039_n_spl_1,
    g1039_n_spl_
  );


  buf

  (
    g1004_n_spl_,
    g1004_n
  );


  buf

  (
    g1004_n_spl_0,
    g1004_n_spl_
  );


  buf

  (
    g1004_n_spl_00,
    g1004_n_spl_0
  );


  buf

  (
    g1004_n_spl_1,
    g1004_n_spl_
  );


  buf

  (
    G15_p_spl_,
    G15_p
  );


  buf

  (
    G36_p_spl_,
    G36_p
  );


  buf

  (
    g1046_n_spl_,
    g1046_n
  );


  buf

  (
    g1046_n_spl_0,
    g1046_n_spl_
  );


  buf

  (
    g1046_n_spl_00,
    g1046_n_spl_0
  );


  buf

  (
    g1046_n_spl_1,
    g1046_n_spl_
  );


  buf

  (
    g1011_n_spl_,
    g1011_n
  );


  buf

  (
    g1011_n_spl_0,
    g1011_n_spl_
  );


  buf

  (
    g1011_n_spl_00,
    g1011_n_spl_0
  );


  buf

  (
    g1011_n_spl_1,
    g1011_n_spl_
  );


  buf

  (
    G77_p_spl_,
    G77_p
  );


  buf

  (
    G87_p_spl_,
    G87_p
  );


  buf

  (
    G75_p_spl_,
    G75_p
  );


  buf

  (
    G85_p_spl_,
    G85_p
  );


  buf

  (
    G74_p_spl_,
    G74_p
  );


  buf

  (
    G84_p_spl_,
    G84_p
  );


  buf

  (
    G73_p_spl_,
    G73_p
  );


  buf

  (
    G83_p_spl_,
    G83_p
  );


  buf

  (
    g1200_p_spl_,
    g1200_p
  );


  buf

  (
    g1202_n_spl_,
    g1202_n
  );


  buf

  (
    g1200_n_spl_,
    g1200_n
  );


  buf

  (
    g1202_p_spl_,
    g1202_p
  );


  buf

  (
    g1214_n_spl_,
    g1214_n
  );


  buf

  (
    g1223_p_spl_,
    g1223_p
  );


  buf

  (
    g1214_p_spl_,
    g1214_p
  );


  buf

  (
    g1223_n_spl_,
    g1223_n
  );


  buf

  (
    g1229_n_spl_,
    g1229_n
  );


  buf

  (
    g1238_p_spl_,
    g1238_p
  );


  buf

  (
    g1229_p_spl_,
    g1229_p
  );


  buf

  (
    g1238_n_spl_,
    g1238_n
  );


  buf

  (
    g1241_p_spl_,
    g1241_p
  );


  buf

  (
    g245_p_spl_,
    g245_p
  );


  buf

  (
    g1241_n_spl_,
    g1241_n
  );


  buf

  (
    g1226_p_spl_,
    g1226_p
  );


  buf

  (
    g1244_n_spl_,
    g1244_n
  );


  buf

  (
    g1226_n_spl_,
    g1226_n
  );


  buf

  (
    g1244_p_spl_,
    g1244_p
  );


  buf

  (
    g1254_n_spl_,
    g1254_n
  );


  buf

  (
    g617_n_spl_,
    g617_n
  );


  buf

  (
    g1254_p_spl_,
    g1254_p
  );


  buf

  (
    g1257_p_spl_,
    g1257_p
  );


  buf

  (
    g1257_n_spl_,
    g1257_n
  );


  buf

  (
    G162_n_spl_,
    G162_n
  );


  buf

  (
    G162_p_spl_,
    G162_p
  );


  buf

  (
    g1260_p_spl_,
    g1260_p
  );


  buf

  (
    g1263_p_spl_,
    g1263_p
  );


  buf

  (
    g1260_n_spl_,
    g1260_n
  );


  buf

  (
    g1263_n_spl_,
    g1263_n
  );


  buf

  (
    g1268_n_spl_,
    g1268_n
  );


  buf

  (
    g1268_p_spl_,
    g1268_p
  );


  buf

  (
    g1266_n_spl_,
    g1266_n
  );


  buf

  (
    g1271_n_spl_,
    g1271_n
  );


  buf

  (
    g1266_p_spl_,
    g1266_p
  );


  buf

  (
    g1271_p_spl_,
    g1271_p
  );


  buf

  (
    g1275_n_spl_,
    g1275_n
  );


  buf

  (
    g1275_p_spl_,
    g1275_p
  );


  buf

  (
    g1278_p_spl_,
    g1278_p
  );


  buf

  (
    g1278_n_spl_,
    g1278_n
  );


  buf

  (
    g1281_p_spl_,
    g1281_p
  );


  buf

  (
    g1281_n_spl_,
    g1281_n
  );


  buf

  (
    g1282_n_spl_,
    g1282_n
  );


  buf

  (
    g1282_p_spl_,
    g1282_p
  );


  buf

  (
    g1284_n_spl_,
    g1284_n
  );


  buf

  (
    g1284_p_spl_,
    g1284_p
  );


  buf

  (
    g1288_n_spl_,
    g1288_n
  );


  buf

  (
    g1288_p_spl_,
    g1288_p
  );


  buf

  (
    g1299_p_spl_,
    g1299_p
  );


  buf

  (
    g1299_n_spl_,
    g1299_n
  );


  buf

  (
    g1308_n_spl_,
    g1308_n
  );


  buf

  (
    g1320_n_spl_,
    g1320_n
  );


  buf

  (
    g1329_p_spl_,
    g1329_p
  );


  buf

  (
    g1320_p_spl_,
    g1320_p
  );


  buf

  (
    g1329_n_spl_,
    g1329_n
  );


  buf

  (
    g1341_n_spl_,
    g1341_n
  );


  buf

  (
    g317_p_spl_,
    g317_p
  );


  buf

  (
    g1341_p_spl_,
    g1341_p
  );


  buf

  (
    g1332_n_spl_,
    g1332_n
  );


  buf

  (
    g1344_p_spl_,
    g1344_p
  );


  buf

  (
    g1332_p_spl_,
    g1332_p
  );


  buf

  (
    g1344_n_spl_,
    g1344_n
  );


  buf

  (
    g1356_n_spl_,
    g1356_n
  );


  buf

  (
    g1365_p_spl_,
    g1365_p
  );


  buf

  (
    g1356_p_spl_,
    g1356_p
  );


  buf

  (
    g1365_n_spl_,
    g1365_n
  );


  buf

  (
    g1377_n_spl_,
    g1377_n
  );


  buf

  (
    g1386_p_spl_,
    g1386_p
  );


  buf

  (
    g1377_p_spl_,
    g1377_p
  );


  buf

  (
    g1386_n_spl_,
    g1386_n
  );


  buf

  (
    g1389_p_spl_,
    g1389_p
  );


  buf

  (
    g1398_n_spl_,
    g1398_n
  );


  buf

  (
    g1389_n_spl_,
    g1389_n
  );


  buf

  (
    g1398_p_spl_,
    g1398_p
  );


  buf

  (
    g1368_p_spl_,
    g1368_p
  );


  buf

  (
    g1401_n_spl_,
    g1401_n
  );


  buf

  (
    g1368_n_spl_,
    g1368_n
  );


  buf

  (
    g1401_p_spl_,
    g1401_p
  );


  buf

  (
    g1409_n_spl_,
    g1409_n
  );


  buf

  (
    g1412_n_spl_,
    g1412_n
  );


  buf

  (
    g1409_p_spl_,
    g1409_p
  );


  buf

  (
    g1412_p_spl_,
    g1412_p
  );


  buf

  (
    g1415_p_spl_,
    g1415_p
  );


  buf

  (
    g1415_n_spl_,
    g1415_n
  );


  buf

  (
    g1416_n_spl_,
    g1416_n
  );


  buf

  (
    g1416_p_spl_,
    g1416_p
  );


  buf

  (
    g1420_p_spl_,
    g1420_p
  );


  buf

  (
    g1420_n_spl_,
    g1420_n
  );


  buf

  (
    g1423_p_spl_,
    g1423_p
  );


  buf

  (
    g1423_n_spl_,
    g1423_n
  );


  buf

  (
    g1426_p_spl_,
    g1426_p
  );


  buf

  (
    g1426_n_spl_,
    g1426_n
  );


  buf

  (
    g1432_p_spl_,
    g1432_p
  );


  buf

  (
    g1432_n_spl_,
    g1432_n
  );


  buf

  (
    g1435_p_spl_,
    g1435_p
  );


  buf

  (
    g1435_n_spl_,
    g1435_n
  );


  buf

  (
    g1438_p_spl_,
    g1438_p
  );


  buf

  (
    g1438_n_spl_,
    g1438_n
  );


  buf

  (
    g1441_n_spl_,
    g1441_n
  );


  buf

  (
    g1441_p_spl_,
    g1441_p
  );


  buf

  (
    g1430_n_spl_,
    g1430_n
  );


  buf

  (
    g1430_p_spl_,
    g1430_p
  );


  buf

  (
    G157_n_spl_,
    G157_n
  );


  buf

  (
    G157_n_spl_0,
    G157_n_spl_
  );


  buf

  (
    G157_n_spl_1,
    G157_n_spl_
  );


  buf

  (
    G157_p_spl_,
    G157_p
  );


  buf

  (
    G157_p_spl_0,
    G157_p_spl_
  );


  buf

  (
    G157_p_spl_1,
    G157_p_spl_
  );


  buf

  (
    g1453_n_spl_,
    g1453_n
  );


  buf

  (
    g1453_p_spl_,
    g1453_p
  );


  buf

  (
    g1458_n_spl_,
    g1458_n
  );


  buf

  (
    g1458_n_spl_0,
    g1458_n_spl_
  );


  buf

  (
    g1458_n_spl_1,
    g1458_n_spl_
  );


  buf

  (
    g1458_p_spl_,
    g1458_p
  );


  buf

  (
    g1458_p_spl_0,
    g1458_p_spl_
  );


  buf

  (
    g1458_p_spl_1,
    g1458_p_spl_
  );


  buf

  (
    g1456_n_spl_,
    g1456_n
  );


  buf

  (
    g1461_p_spl_,
    g1461_p
  );


  buf

  (
    g1456_p_spl_,
    g1456_p
  );


  buf

  (
    g1461_n_spl_,
    g1461_n
  );


  buf

  (
    g1464_n_spl_,
    g1464_n
  );


  buf

  (
    g1464_p_spl_,
    g1464_p
  );


  buf

  (
    g1471_n_spl_,
    g1471_n
  );


  buf

  (
    g1471_p_spl_,
    g1471_p
  );


  buf

  (
    g1470_n_spl_,
    g1470_n
  );


  buf

  (
    g1474_p_spl_,
    g1474_p
  );


  buf

  (
    g1470_p_spl_,
    g1470_p
  );


  buf

  (
    g1474_n_spl_,
    g1474_n
  );


  buf

  (
    g1469_n_spl_,
    g1469_n
  );


  buf

  (
    g1477_p_spl_,
    g1477_p
  );


  buf

  (
    g1469_p_spl_,
    g1469_p
  );


  buf

  (
    g1477_n_spl_,
    g1477_n
  );


  buf

  (
    g1480_n_spl_,
    g1480_n
  );


  buf

  (
    g1483_p_spl_,
    g1483_p
  );


  buf

  (
    g1480_p_spl_,
    g1480_p
  );


  buf

  (
    g1483_n_spl_,
    g1483_n
  );


  buf

  (
    g1488_p_spl_,
    g1488_p
  );


  buf

  (
    g1488_n_spl_,
    g1488_n
  );


  buf

  (
    g1491_n_spl_,
    g1491_n
  );


  buf

  (
    g1491_p_spl_,
    g1491_p
  );


  buf

  (
    g1500_n_spl_,
    g1500_n
  );


  buf

  (
    G23_n_spl_,
    G23_n
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    g1509_p_spl_,
    g1509_p
  );


  buf

  (
    g1509_p_spl_0,
    g1509_p_spl_
  );


  buf

  (
    g1509_p_spl_1,
    g1509_p_spl_
  );


  buf

  (
    g1512_p_spl_,
    g1512_p
  );


  buf

  (
    g1512_p_spl_0,
    g1512_p_spl_
  );


  buf

  (
    g1512_p_spl_1,
    g1512_p_spl_
  );


  buf

  (
    G79_n_spl_,
    G79_n
  );


  buf

  (
    G78_n_spl_,
    G78_n
  );


  buf

  (
    G64_n_spl_,
    G64_n
  );


  buf

  (
    G151_n_spl_,
    G151_n
  );


  buf

  (
    G151_n_spl_0,
    G151_n_spl_
  );


  buf

  (
    G152_p_spl_,
    G152_p
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    G1_n_spl_1,
    G1_n_spl_
  );


  buf

  (
    g194_n_spl_,
    g194_n
  );


  buf

  (
    g431_n_spl_,
    g431_n
  );


  buf

  (
    g482_p_spl_,
    g482_p
  );


  buf

  (
    g549_p_spl_,
    g549_p
  );


  buf

  (
    g550_n_spl_,
    g550_n
  );


endmodule
