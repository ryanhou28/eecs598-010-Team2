module c432(G1,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,
  G24,G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G34,G35,G36,G4,G426,G427,G428,
  G429,G430,G431,G432,G5,G6,G7,G8,G9);
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
  G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36;
output G426,G427,G428,G429,G430,G431,G432;

  wire G118,G119,G122,G123,G126,G127,G130,G131,G134,G135,G138,G139,G142,G143,
    G146,G147,G150,G151,G154,G157,G158,G159,G162,G165,G168,G171,G174,G177,G180,
    G183,G184,G185,G186,G187,G188,G189,G190,G191,G192,G193,G194,G195,G196,G197,
    G198,G199,G203,G213,G223,G226,G229,G232,G235,G238,G241,G242,G245,G246,G249,
    G250,G253,G254,G255,G256,G257,G258,G259,G262,G263,G266,G269,G272,G275,G278,
    G281,G284,G287,G288,G289,G290,G291,G292,G293,G294,G295,G299,G300,G301,G302,
    G303,G304,G305,G306,G307,G308,G318,G328,G329,G330,G331,G332,G333,G334,G335,
    G336,G337,G338,G339,G340,G341,G342,G343,G344,G345,G346,G347,G348,G349,G350,
    G351,G352,G353,G354,G355,G358,G368,G369,G370,G371,G372,G373,G374,G375,G376,
    G377,G378,G383,G390,G396,G401,G404,G408,G411,G412,G413,G414,G415,G416,G417,
    G418,G421,G424,G425;

  not (G118,G1);
  not (G119,G2);
  not (G122,G4);
  not (G123,G6);
  not (G126,G8);
  not (G127,G10);
  not (G130,G12);
  not (G131,G14);
  not (G134,G16);
  not (G135,G18);
  not (G138,G20);
  not (G139,G22);
  not (G142,G24);
  not (G143,G26);
  not (G146,G28);
  not (G147,G30);
  not (G150,G32);
  not (G151,G34);
  nand (G154,G118,G2);
  nor (G157,G3,G119);
  nor (G158,G5,G119);
  nand (G159,G122,G6);
  nand (G162,G126,G10);
  nand (G165,G130,G14);
  nand (G168,G134,G18);
  nand (G171,G138,G22);
  nand (G174,G142,G26);
  nand (G177,G146,G30);
  nand (G180,G150,G34);
  nor (G183,G7,G123);
  nor (G184,G9,G123);
  nor (G185,G11,G127);
  nor (G186,G13,G127);
  nor (G187,G15,G131);
  nor (G188,G17,G131);
  nor (G189,G19,G135);
  nor (G190,G21,G135);
  nor (G191,G23,G139);
  nor (G192,G25,G139);
  nor (G193,G27,G143);
  nor (G194,G29,G143);
  nor (G195,G31,G147);
  nor (G196,G33,G147);
  nor (G197,G35,G151);
  nor (G198,G36,G151);
  and (G199,G154,G159,G162,G165,G168,G171,G174,G177,G180);
  not (G203,G199);
  not (G213,G199);
  xor (G223,G203,G154);
  xor (G226,G203,G159);
  xor (G229,G203,G162);
  xor (G232,G203,G165);
  xor (G235,G203,G168);
  xor (G238,G203,G171);
  nand (G241,G1,G213);
  xor (G242,G203,G174);
  nand (G245,G213,G4);
  xor (G246,G203,G177);
  nand (G249,G213,G8);
  xor (G250,G203,G180);
  nand (G253,G213,G12);
  nand (G254,G213,G16);
  nand (G255,G213,G20);
  nand (G256,G213,G24);
  nand (G257,G213,G28);
  nand (G258,G213,G32);
  nand (G259,G223,G157);
  nand (G262,G223,G158);
  nand (G263,G226,G183);
  nand (G266,G229,G185);
  nand (G269,G232,G187);
  nand (G272,G235,G189);
  nand (G275,G238,G191);
  nand (G278,G242,G193);
  nand (G281,G246,G195);
  nand (G284,G250,G197);
  nand (G287,G226,G184);
  nand (G288,G229,G186);
  nand (G289,G232,G188);
  nand (G290,G235,G190);
  nand (G291,G238,G192);
  nand (G292,G242,G194);
  nand (G293,G246,G196);
  nand (G294,G250,G198);
  and (G295,G259,G263,G266,G269,G272,G275,G278,G281,G284);
  not (G299,G262);
  not (G300,G287);
  not (G301,G288);
  not (G302,G289);
  not (G303,G290);
  not (G304,G291);
  not (G305,G292);
  not (G306,G293);
  not (G307,G294);
  not (G308,G295);
  not (G318,G295);
  xor (G328,G308,G259);
  xor (G329,G308,G263);
  xor (G330,G308,G266);
  xor (G331,G308,G269);
  nand (G332,G3,G318);
  xor (G333,G308,G272);
  nand (G334,G318,G7);
  xor (G335,G308,G275);
  nand (G336,G318,G11);
  xor (G337,G308,G278);
  nand (G338,G318,G15);
  xor (G339,G308,G281);
  nand (G340,G318,G19);
  xor (G341,G308,G284);
  nand (G342,G318,G23);
  nand (G343,G318,G27);
  nand (G344,G318,G31);
  nand (G345,G318,G35);
  nand (G346,G328,G299);
  nand (G347,G329,G300);
  nand (G348,G330,G301);
  nand (G349,G331,G302);
  nand (G350,G333,G303);
  nand (G351,G335,G304);
  nand (G352,G337,G305);
  nand (G353,G339,G306);
  nand (G354,G341,G307);
  and (G355,G346,G347,G348,G349,G350,G351,G352,G353,G354);
  not (G358,G355);
  nand (G368,G5,G358);
  nand (G369,G358,G9);
  nand (G370,G358,G13);
  nand (G371,G358,G17);
  nand (G372,G358,G21);
  nand (G373,G358,G25);
  nand (G374,G358,G29);
  nand (G375,G358,G33);
  nand (G376,G358,G36);
  nand (G377,G2,G241,G332,G368);
  nand (G378,G245,G334,G369,G6);
  nand (G383,G249,G336,G370,G10);
  nand (G390,G253,G338,G371,G14);
  nand (G396,G254,G340,G372,G18);
  nand (G401,G255,G342,G373,G22);
  nand (G404,G256,G343,G374,G26);
  nand (G408,G257,G344,G375,G30);
  nand (G411,G258,G345,G376,G34);
  not (G412,G377);
  and (G413,G378,G383,G390,G396,G401,G404,G408,G411);
  not (G414,G390);
  not (G415,G401);
  not (G416,G404);
  not (G417,G408);
  nand (G418,G383,G414);
  nand (G421,G383,G390,G415,G396);
  nand (G424,G396,G390,G416);
  nand (G425,G383,G390,G404,G417);
  not (G426,G199);
  not (G427,G295);
  not (G428,G355);
  nor (G429,G412,G413);
  nand (G430,G378,G383,G418,G396);
  nand (G431,G378,G383,G421,G424);
  nand (G432,G378,G418,G421,G425);

endmodule
