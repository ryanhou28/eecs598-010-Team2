// Benchmark "mymod" written by ABC on Wed Nov  1 23:37:42 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58,
    G59, G60,
    G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, G865, G866,
    G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, G877, G878,
    G879, G880  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G58, G59, G60;
  output G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, G865,
    G866, G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, G877,
    G878, G879, G880;
  reg n492_lo, n495_lo, n498_lo, n501_lo, n516_lo, n528_lo, n540_lo,
    n543_lo, n546_lo, n549_lo, n552_lo, n564_lo, n600_lo, n603_lo, n606_lo,
    n609_lo, n615_lo, n618_lo, n621_lo, n627_lo, n630_lo, n633_lo, n639_lo,
    n642_lo, n645_lo, n648_lo, n660_lo, n672_lo, n675_lo, n678_lo, n681_lo,
    n684_lo, n687_lo, n690_lo, n693_lo, n696_lo, n699_lo, n702_lo, n705_lo,
    n708_lo, n711_lo, n714_lo, n717_lo, n720_lo, n723_lo, n726_lo, n729_lo,
    n732_lo, n735_lo, n738_lo, n741_lo, n744_lo, n747_lo, n750_lo, n753_lo,
    n756_lo, n759_lo, n762_lo, n765_lo, n768_lo, n771_lo, n774_lo, n777_lo,
    n780_lo, n783_lo, n786_lo, n792_lo, n795_lo, n798_lo, n807_lo, n816_lo,
    n819_lo, n828_lo, n831_lo, n843_lo, n846_lo, n849_lo, n852_lo, n855_lo,
    n858_lo, n861_lo, n864_lo, n867_lo, n870_lo, n879_lo, n882_lo, n891_lo,
    n903_lo, n915_lo, n918_lo, n951_lo, n954_lo, n957_lo, n960_lo, n963_lo,
    n966_lo, n969_lo, n972_lo, n975_lo, n978_lo, n981_lo, n984_lo, n987_lo,
    n990_lo, n993_lo, n996_lo, n999_lo, n1002_lo, n1008_lo, n1011_lo,
    n1014_lo, n1020_lo, n1023_lo, n1032_lo, n1035_lo, n1044_lo, n1047_lo,
    n1050_lo, n1053_lo, n1056_lo, n1059_lo, n1062_lo, n1065_lo, n1068_lo,
    n1071_lo, n1074_lo, n1077_lo, n1080_lo, n1083_lo, n1086_lo, n1089_lo,
    n1092_lo, n1095_lo, n1098_lo, n1101_lo, n1104_lo, n1107_lo, n1110_lo,
    n1113_lo, n1116_lo, n1119_lo, n1122_lo, n1125_lo, n1128_lo, n1131_lo,
    n1134_lo, n1137_lo, n1143_lo, n1146_lo, n1149_lo, n1152_lo, n1155_lo,
    n1164_lo, n1167_lo, n1170_lo, n1173_lo, n1176_lo, n1188_lo, n563_inv,
    n1429_o2, n1427_o2, n1471_o2, n1476_o2, n1499_o2, n1500_o2, n1501_o2,
    n1516_o2, n1517_o2, n1562_o2, n1563_o2, n1564_o2, n1582_o2, n1583_o2,
    n1618_o2, n1622_o2, n1502_o2, n1503_o2, n1504_o2, n1505_o2, n1506_o2,
    n1512_o2, n1513_o2, n1514_o2, n1515_o2, n1644_o2, n1647_o2, n1527_o2,
    n650_inv, n653_inv, n656_inv, n1567_o2, n955_o2, n1568_o2, n1037_o2,
    n960_o2, n1587_o2, n1040_o2, n1039_o2, n1589_o2, n1624_o2, n1643_o2,
    n1038_o2, n1645_o2, n1029_o2, n701_inv, n1662_o2, n1663_o2, n710_inv,
    n813_o2, lo114_buf_o2, n1031_o2, lo186_buf_o2, n1042_o2, n728_inv,
    n917_o2, n734_inv, n1649_o2, n1650_o2, n1651_o2, n1652_o2, n1653_o2,
    lo138_buf_o2, n1664_o2, n1665_o2, n1666_o2, n1667_o2, n944_o2,
    n770_inv, n1672_o2, n776_inv, n1679_o2, n782_inv, n785_inv,
    lo110_buf_o2, lo134_buf_o2, n1030_o2, lo182_buf_o2, n830_o2, n1021_o2,
    n806_inv, n809_inv, n946_o2, lo038_buf_o2, lo238_buf_o2, n1010_o2,
    n1006_o2, n907_o2, n902_o2, lo154_buf_o2, n836_inv, n839_inv,
    lo122_buf_o2, n845_inv, n904_o2, lo106_buf_o2, n980_o2, n1023_o2,
    lo178_buf_o2, n981_o2, n837_o2, n1013_o2, n840_o2, n849_o2, n852_o2,
    n864_o2, n867_o2, n1044_o2, n876_o2, n893_inv, n879_o2, n925_o2,
    n902_inv, lo146_buf_o2, n1026_o2, n1032_o2, lo118_buf_o2, n917_inv,
    lo190_buf_o2, n1036_o2, n926_inv, n929_inv, lo002_buf_o2, lo014_buf_o2,
    lo030_buf_o2, lo034_buf_o2, lo042_buf_o2, lo113_buf_o2, lo185_buf_o2,
    n939_o2, n941_o2, lo142_buf_o2, lo230_buf_o2, lo006_buf_o2,
    lo018_buf_o2, lo022_buf_o2, lo066_buf_o2, n977_inv, n826_o2, n892_o2,
    lo152_buf_o2, n896_o2, n905_o2, n995_inv, lo037_buf_o2, lo237_buf_o2,
    lo062_buf_o2, n1007_inv, n1010_inv, n891_o2;
  wire new_n705_, new_n706_, new_n707_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n731_, new_n733_, new_n735_, new_n737_, new_n739_,
    new_n741_, new_n743_, new_n745_, new_n747_, new_n749_, new_n751_,
    new_n753_, new_n755_, new_n757_, new_n759_, new_n761_, new_n763_,
    new_n765_, new_n767_, new_n769_, new_n771_, new_n773_, new_n775_,
    new_n777_, new_n779_, new_n781_, new_n784_, new_n785_, new_n787_,
    new_n789_, new_n791_, new_n793_, new_n795_, new_n797_, new_n799_,
    new_n801_, new_n803_, new_n805_, new_n807_, new_n809_, new_n811_,
    new_n813_, new_n815_, new_n817_, new_n819_, new_n821_, new_n823_,
    new_n826_, new_n827_, new_n829_, new_n832_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n850_, new_n851_, new_n853_,
    new_n856_, new_n857_, new_n859_, new_n862_, new_n863_, new_n865_,
    new_n868_, new_n869_, new_n871_, new_n873_, new_n876_, new_n878_,
    new_n880_, new_n881_, new_n883_, new_n885_, new_n888_, new_n889_,
    new_n891_, new_n893_, new_n896_, new_n897_, new_n899_, new_n901_,
    new_n903_, new_n905_, new_n907_, new_n909_, new_n911_, new_n913_,
    new_n915_, new_n917_, new_n919_, new_n921_, new_n923_, new_n925_,
    new_n927_, new_n929_, new_n931_, new_n933_, new_n934_, new_n936_,
    new_n937_, new_n939_, new_n941_, new_n942_, new_n944_, new_n945_,
    new_n947_, new_n949_, new_n950_, new_n952_, new_n953_, new_n955_,
    new_n958_, new_n959_, new_n961_, new_n963_, new_n966_, new_n967_,
    new_n970_, new_n971_, new_n973_, new_n975_, new_n977_, new_n979_,
    new_n980_, new_n981_, new_n983_, new_n985_, new_n987_, new_n988_,
    new_n989_, new_n991_, new_n992_, new_n993_, new_n995_, new_n997_,
    new_n999_, new_n1001_, new_n1004_, new_n1005_, new_n1007_, new_n1009_,
    new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1015_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1023_, new_n1025_,
    new_n1026_, new_n1028_, new_n1029_, new_n1031_, new_n1033_, new_n1034_,
    new_n1036_, new_n1037_, new_n1039_, new_n1042_, new_n1043_, new_n1045_,
    new_n1046_, new_n1048_, new_n1049_, new_n1052_, new_n1053_, new_n1056_,
    new_n1057_, new_n1059_, new_n1061_, new_n1063_, new_n1064_, new_n1065_,
    new_n1067_, new_n1069_, new_n1072_, new_n1073_, new_n1075_, new_n1077_,
    new_n1080_, new_n1081_, new_n1083_, new_n1085_, new_n1088_, new_n1089_,
    new_n1091_, new_n1093_, new_n1096_, new_n1097_, new_n1099_, new_n1101_,
    new_n1104_, new_n1105_, new_n1107_, new_n1109_, new_n1112_, new_n1113_,
    new_n1115_, new_n1117_, new_n1119_, new_n1121_, new_n1123_, new_n1126_,
    new_n1127_, new_n1130_, new_n1131_, new_n1133_, new_n1135_, new_n1138_,
    new_n1140_, new_n1142_, new_n1144_, new_n1145_, new_n1148_, new_n1150_,
    new_n1151_, new_n1152_, new_n1153_, new_n1156_, new_n1158_, new_n1160_,
    new_n1161_, new_n1162_, new_n1164_, new_n1165_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1174_, new_n1176_,
    new_n1177_, new_n1179_, new_n1181_, new_n1183_, new_n1185_, new_n1186_,
    new_n1187_, new_n1189_, new_n1191_, new_n1194_, new_n1196_, new_n1197_,
    new_n1199_, new_n1200_, new_n1201_, new_n1203_, new_n1206_, new_n1207_,
    new_n1208_, new_n1209_, new_n1212_, new_n1213_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1232_, new_n1233_, new_n1235_, new_n1237_, new_n1239_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1253_, new_n1255_,
    new_n1257_, new_n1259_, new_n1260_, new_n1261_, new_n1263_, new_n1265_,
    new_n1267_, new_n1269_, new_n1271_, new_n1273_, new_n1275_, new_n1277_,
    new_n1279_, new_n1281_, new_n1283_, new_n1285_, new_n1287_, new_n1288_,
    new_n1289_, new_n1291_, new_n1292_, new_n1293_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1300_, new_n1301_, new_n1302_, new_n1303_,
    new_n1305_, new_n1307_, new_n1309_, new_n1310_, new_n1311_, new_n1313_,
    new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1320_,
    new_n1322_, new_n1323_, new_n1325_, new_n1327_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1336_, new_n1337_,
    new_n1338_, new_n1339_, new_n1340_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1363_,
    new_n1364_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1372_,
    new_n1374_, new_n1375_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1391_, new_n1393_, new_n1395_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1402_, new_n1404_, new_n1405_,
    new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1411_, new_n1413_,
    new_n1415_, new_n1417_, new_n1418_, new_n1419_, new_n1421_, new_n1423_,
    new_n1425_, new_n1427_, new_n1429_, new_n1430_, new_n1431_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1439_, new_n1441_,
    new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_,
    new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_,
    new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_,
    new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_,
    new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_,
    new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_,
    new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_,
    new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_,
    new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_,
    new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_,
    new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_,
    new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_,
    new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_,
    new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_,
    new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_,
    new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_,
    new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_,
    new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_,
    new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_,
    new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_,
    new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_,
    new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_,
    new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_,
    new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_,
    new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_,
    new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_,
    new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_,
    new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_,
    new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_,
    new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_,
    new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_,
    new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_,
    new_n1779_, new_n1780_, new_n2116_, new_n2117_, new_n2118_, new_n2119_,
    new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_,
    new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_,
    new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_,
    new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_,
    new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_,
    new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_,
    new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_,
    new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_,
    new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_,
    new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_,
    new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_,
    new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_,
    new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_,
    new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_,
    new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_,
    new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_,
    new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_,
    new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_,
    new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_,
    new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_,
    new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_,
    new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_,
    new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_,
    new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_,
    new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_,
    new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_,
    new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_,
    new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_,
    new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_,
    new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_,
    new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_,
    new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_,
    new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_,
    new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_,
    new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_,
    new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_,
    new_n2336_, new_n2337_, new_n2338_, n1654_li007_li007,
    n1657_li008_li008, n1660_li009_li009, n1663_li010_li010,
    n1678_li015_li015, n1690_li019_li019, n1702_li023_li023,
    n1705_li024_li024, n1708_li025_li025, n1711_li026_li026,
    n1714_li027_li027, n1726_li031_li031, n1762_li043_li043,
    n1765_li044_li044, n1768_li045_li045, n1771_li046_li046,
    n1777_li048_li048, n1780_li049_li049, n1783_li050_li050,
    n1789_li052_li052, n1792_li053_li053, n1795_li054_li054,
    n1801_li056_li056, n1804_li057_li057, n1807_li058_li058,
    n1810_li059_li059, n1822_li063_li063, n1834_li067_li067,
    n1837_li068_li068, n1840_li069_li069, n1843_li070_li070,
    n1846_li071_li071, n1849_li072_li072, n1852_li073_li073,
    n1855_li074_li074, n1858_li075_li075, n1861_li076_li076,
    n1864_li077_li077, n1867_li078_li078, n1870_li079_li079,
    n1873_li080_li080, n1876_li081_li081, n1879_li082_li082,
    n1882_li083_li083, n1885_li084_li084, n1888_li085_li085,
    n1891_li086_li086, n1894_li087_li087, n1897_li088_li088,
    n1900_li089_li089, n1903_li090_li090, n1906_li091_li091,
    n1909_li092_li092, n1912_li093_li093, n1915_li094_li094,
    n1918_li095_li095, n1921_li096_li096, n1924_li097_li097,
    n1927_li098_li098, n1930_li099_li099, n1933_li100_li100,
    n1936_li101_li101, n1939_li102_li102, n1942_li103_li103,
    n1945_li104_li104, n1948_li105_li105, n1954_li107_li107,
    n1957_li108_li108, n1960_li109_li109, n1969_li112_li112,
    n1978_li115_li115, n1981_li116_li116, n1990_li119_li119,
    n1993_li120_li120, n2005_li124_li124, n2008_li125_li125,
    n2011_li126_li126, n2014_li127_li127, n2017_li128_li128,
    n2020_li129_li129, n2023_li130_li130, n2026_li131_li131,
    n2029_li132_li132, n2032_li133_li133, n2041_li136_li136,
    n2044_li137_li137, n2053_li140_li140, n2065_li144_li144,
    n2077_li148_li148, n2080_li149_li149, n2113_li160_li160,
    n2116_li161_li161, n2119_li162_li162, n2122_li163_li163,
    n2125_li164_li164, n2128_li165_li165, n2131_li166_li166,
    n2134_li167_li167, n2137_li168_li168, n2140_li169_li169,
    n2143_li170_li170, n2146_li171_li171, n2149_li172_li172,
    n2152_li173_li173, n2155_li174_li174, n2158_li175_li175,
    n2161_li176_li176, n2164_li177_li177, n2170_li179_li179,
    n2173_li180_li180, n2176_li181_li181, n2182_li183_li183,
    n2185_li184_li184, n2194_li187_li187, n2197_li188_li188,
    n2206_li191_li191, n2209_li192_li192, n2212_li193_li193,
    n2215_li194_li194, n2218_li195_li195, n2221_li196_li196,
    n2224_li197_li197, n2227_li198_li198, n2230_li199_li199,
    n2233_li200_li200, n2236_li201_li201, n2239_li202_li202,
    n2242_li203_li203, n2245_li204_li204, n2248_li205_li205,
    n2251_li206_li206, n2254_li207_li207, n2257_li208_li208,
    n2260_li209_li209, n2263_li210_li210, n2266_li211_li211,
    n2269_li212_li212, n2272_li213_li213, n2275_li214_li214,
    n2278_li215_li215, n2281_li216_li216, n2284_li217_li217,
    n2287_li218_li218, n2290_li219_li219, n2293_li220_li220,
    n2296_li221_li221, n2299_li222_li222, n2305_li224_li224,
    n2308_li225_li225, n2311_li226_li226, n2314_li227_li227,
    n2317_li228_li228, n2326_li231_li231, n2329_li232_li232,
    n2332_li233_li233, n2335_li234_li234, n2338_li235_li235,
    n2350_li239_li239, n1428_i2, n1429_i2, n1427_i2, n1471_i2, n1476_i2,
    n1499_i2, n1500_i2, n1501_i2, n1516_i2, n1517_i2, n1562_i2, n1563_i2,
    n1564_i2, n1582_i2, n1583_i2, n1618_i2, n1622_i2, n1502_i2, n1503_i2,
    n1504_i2, n1505_i2, n1506_i2, n1512_i2, n1513_i2, n1514_i2, n1515_i2,
    n1644_i2, n1647_i2, n1527_i2, n1526_i2, n1528_i2, n1529_i2, n1567_i2,
    n955_i2, n1568_i2, n1037_i2, n960_i2, n1587_i2, n1040_i2, n1039_i2,
    n1589_i2, n1624_i2, n1643_i2, n1038_i2, n1645_i2, n1029_i2, n1648_i2,
    n1662_i2, n1663_i2, n1668_i2, n813_i2, lo114_buf_i2, n1031_i2,
    lo186_buf_i2, n1042_i2, n911_i2, n917_i2, n942_i2, n1649_i2, n1650_i2,
    n1651_i2, n1652_i2, n1653_i2, lo138_buf_i2, n1664_i2, n1665_i2,
    n1666_i2, n1667_i2, n944_i2, n945_i2, n1672_i2, n1676_i2, n1679_i2,
    n1680_i2, n1681_i2, lo110_buf_i2, lo134_buf_i2, n1030_i2, lo182_buf_i2,
    n830_i2, n1021_i2, n943_i2, n936_i2, n946_i2, lo038_buf_i2,
    lo238_buf_i2, n1010_i2, n1006_i2, n907_i2, n902_i2, lo154_buf_i2,
    n938_i2, n947_i2, lo122_buf_i2, n899_i2, n904_i2, lo106_buf_i2,
    n980_i2, n1023_i2, lo178_buf_i2, n981_i2, n837_i2, n1013_i2, n840_i2,
    n849_i2, n852_i2, n864_i2, n867_i2, n1044_i2, n876_i2, n937_i2,
    n879_i2, n925_i2, n954_i2, lo146_buf_i2, n1026_i2, n1032_i2,
    lo118_buf_i2, n957_i2, lo190_buf_i2, n1036_i2, n949_i2, n910_i2,
    lo002_buf_i2, lo014_buf_i2, lo030_buf_i2, lo034_buf_i2, lo042_buf_i2,
    lo113_buf_i2, lo185_buf_i2, n939_i2, n941_i2, lo142_buf_i2,
    lo230_buf_i2, lo006_buf_i2, lo018_buf_i2, lo022_buf_i2, lo066_buf_i2,
    n913_i2, n826_i2, n892_i2, lo152_buf_i2, n896_i2, n905_i2, n821_i2,
    lo037_buf_i2, lo237_buf_i2, lo062_buf_i2, n827_i2, n809_i2, n891_i2;
  assign new_n705_ = G1;
  assign new_n706_ = ~G1;
  assign new_n707_ = G2;
  assign new_n709_ = G3;
  assign new_n711_ = G4;
  assign new_n712_ = ~G4;
  assign new_n713_ = G5;
  assign new_n714_ = ~G5;
  assign new_n715_ = G6;
  assign new_n717_ = G7;
  assign new_n719_ = G8;
  assign new_n720_ = ~G8;
  assign new_n721_ = G9;
  assign new_n722_ = ~G9;
  assign new_n723_ = G10;
  assign new_n725_ = G11;
  assign new_n726_ = ~G11;
  assign new_n727_ = G12;
  assign new_n729_ = G13;
  assign new_n731_ = G14;
  assign new_n733_ = G15;
  assign new_n735_ = G16;
  assign new_n737_ = G17;
  assign new_n739_ = G18;
  assign new_n741_ = G19;
  assign new_n743_ = G20;
  assign new_n745_ = G21;
  assign new_n747_ = G22;
  assign new_n749_ = G23;
  assign new_n751_ = G24;
  assign new_n753_ = G25;
  assign new_n755_ = G26;
  assign new_n757_ = G27;
  assign new_n759_ = G28;
  assign new_n761_ = G29;
  assign new_n763_ = G30;
  assign new_n765_ = G31;
  assign new_n767_ = G32;
  assign new_n769_ = G33;
  assign new_n771_ = G34;
  assign new_n773_ = G35;
  assign new_n775_ = G36;
  assign new_n777_ = G37;
  assign new_n779_ = G38;
  assign new_n781_ = G39;
  assign new_n784_ = ~G40;
  assign new_n785_ = G41;
  assign new_n787_ = G42;
  assign new_n789_ = G43;
  assign new_n791_ = G44;
  assign new_n793_ = G45;
  assign new_n795_ = G46;
  assign new_n797_ = G47;
  assign new_n799_ = G48;
  assign new_n801_ = G49;
  assign new_n803_ = G50;
  assign new_n805_ = G51;
  assign new_n807_ = G52;
  assign new_n809_ = G53;
  assign new_n811_ = G54;
  assign new_n813_ = G55;
  assign new_n815_ = G56;
  assign new_n817_ = G57;
  assign new_n819_ = G58;
  assign new_n821_ = G59;
  assign new_n823_ = G60;
  assign new_n826_ = ~n492_lo;
  assign new_n827_ = n495_lo;
  assign new_n829_ = n498_lo;
  assign new_n832_ = ~n501_lo;
  assign new_n834_ = ~n516_lo;
  assign new_n836_ = ~n528_lo;
  assign new_n837_ = n540_lo;
  assign new_n838_ = ~n540_lo;
  assign new_n839_ = n543_lo;
  assign new_n841_ = n546_lo;
  assign new_n843_ = n549_lo;
  assign new_n845_ = n552_lo;
  assign new_n846_ = ~n552_lo;
  assign new_n847_ = n564_lo;
  assign new_n848_ = ~n564_lo;
  assign new_n850_ = ~n600_lo;
  assign new_n851_ = n603_lo;
  assign new_n853_ = n606_lo;
  assign new_n856_ = ~n609_lo;
  assign new_n857_ = n615_lo;
  assign new_n859_ = n618_lo;
  assign new_n862_ = ~n621_lo;
  assign new_n863_ = n627_lo;
  assign new_n865_ = n630_lo;
  assign new_n868_ = ~n633_lo;
  assign new_n869_ = n639_lo;
  assign new_n871_ = n642_lo;
  assign new_n873_ = n645_lo;
  assign new_n876_ = ~n648_lo;
  assign new_n878_ = ~n660_lo;
  assign new_n880_ = ~n672_lo;
  assign new_n881_ = n675_lo;
  assign new_n883_ = n678_lo;
  assign new_n885_ = n681_lo;
  assign new_n888_ = ~n684_lo;
  assign new_n889_ = n687_lo;
  assign new_n891_ = n690_lo;
  assign new_n893_ = n693_lo;
  assign new_n896_ = ~n696_lo;
  assign new_n897_ = n699_lo;
  assign new_n899_ = n702_lo;
  assign new_n901_ = n705_lo;
  assign new_n903_ = n708_lo;
  assign new_n905_ = n711_lo;
  assign new_n907_ = n714_lo;
  assign new_n909_ = n717_lo;
  assign new_n911_ = n720_lo;
  assign new_n913_ = n723_lo;
  assign new_n915_ = n726_lo;
  assign new_n917_ = n729_lo;
  assign new_n919_ = n732_lo;
  assign new_n921_ = n735_lo;
  assign new_n923_ = n738_lo;
  assign new_n925_ = n741_lo;
  assign new_n927_ = n744_lo;
  assign new_n929_ = n747_lo;
  assign new_n931_ = n750_lo;
  assign new_n933_ = n753_lo;
  assign new_n934_ = ~n753_lo;
  assign new_n936_ = ~n756_lo;
  assign new_n937_ = n759_lo;
  assign new_n939_ = n762_lo;
  assign new_n941_ = n765_lo;
  assign new_n942_ = ~n765_lo;
  assign new_n944_ = ~n768_lo;
  assign new_n945_ = n771_lo;
  assign new_n947_ = n774_lo;
  assign new_n949_ = n777_lo;
  assign new_n950_ = ~n777_lo;
  assign new_n952_ = ~n780_lo;
  assign new_n953_ = n783_lo;
  assign new_n955_ = n786_lo;
  assign new_n958_ = ~n792_lo;
  assign new_n959_ = n795_lo;
  assign new_n961_ = n798_lo;
  assign new_n963_ = n807_lo;
  assign new_n966_ = ~n816_lo;
  assign new_n967_ = n819_lo;
  assign new_n970_ = ~n828_lo;
  assign new_n971_ = n831_lo;
  assign new_n973_ = n843_lo;
  assign new_n975_ = n846_lo;
  assign new_n977_ = n849_lo;
  assign new_n979_ = n852_lo;
  assign new_n980_ = ~n852_lo;
  assign new_n981_ = n855_lo;
  assign new_n983_ = n858_lo;
  assign new_n985_ = n861_lo;
  assign new_n987_ = n864_lo;
  assign new_n988_ = ~n864_lo;
  assign new_n989_ = n867_lo;
  assign new_n991_ = n870_lo;
  assign new_n992_ = ~n870_lo;
  assign new_n993_ = n879_lo;
  assign new_n995_ = n882_lo;
  assign new_n997_ = n891_lo;
  assign new_n999_ = n903_lo;
  assign new_n1001_ = n915_lo;
  assign new_n1004_ = ~n918_lo;
  assign new_n1005_ = n951_lo;
  assign new_n1007_ = n954_lo;
  assign new_n1009_ = n957_lo;
  assign new_n1010_ = ~n957_lo;
  assign new_n1011_ = n960_lo;
  assign new_n1012_ = ~n960_lo;
  assign new_n1013_ = n963_lo;
  assign new_n1015_ = n966_lo;
  assign new_n1017_ = n969_lo;
  assign new_n1018_ = ~n969_lo;
  assign new_n1019_ = n972_lo;
  assign new_n1020_ = ~n972_lo;
  assign new_n1021_ = n975_lo;
  assign new_n1023_ = n978_lo;
  assign new_n1025_ = n981_lo;
  assign new_n1026_ = ~n981_lo;
  assign new_n1028_ = ~n984_lo;
  assign new_n1029_ = n987_lo;
  assign new_n1031_ = n990_lo;
  assign new_n1033_ = n993_lo;
  assign new_n1034_ = ~n993_lo;
  assign new_n1036_ = ~n996_lo;
  assign new_n1037_ = n999_lo;
  assign new_n1039_ = n1002_lo;
  assign new_n1042_ = ~n1008_lo;
  assign new_n1043_ = n1011_lo;
  assign new_n1045_ = n1014_lo;
  assign new_n1046_ = ~n1014_lo;
  assign new_n1048_ = ~n1020_lo;
  assign new_n1049_ = n1023_lo;
  assign new_n1052_ = ~n1032_lo;
  assign new_n1053_ = n1035_lo;
  assign new_n1056_ = ~n1044_lo;
  assign new_n1057_ = n1047_lo;
  assign new_n1059_ = n1050_lo;
  assign new_n1061_ = n1053_lo;
  assign new_n1063_ = n1056_lo;
  assign new_n1064_ = ~n1056_lo;
  assign new_n1065_ = n1059_lo;
  assign new_n1067_ = n1062_lo;
  assign new_n1069_ = n1065_lo;
  assign new_n1072_ = ~n1068_lo;
  assign new_n1073_ = n1071_lo;
  assign new_n1075_ = n1074_lo;
  assign new_n1077_ = n1077_lo;
  assign new_n1080_ = ~n1080_lo;
  assign new_n1081_ = n1083_lo;
  assign new_n1083_ = n1086_lo;
  assign new_n1085_ = n1089_lo;
  assign new_n1088_ = ~n1092_lo;
  assign new_n1089_ = n1095_lo;
  assign new_n1091_ = n1098_lo;
  assign new_n1093_ = n1101_lo;
  assign new_n1096_ = ~n1104_lo;
  assign new_n1097_ = n1107_lo;
  assign new_n1099_ = n1110_lo;
  assign new_n1101_ = n1113_lo;
  assign new_n1104_ = ~n1116_lo;
  assign new_n1105_ = n1119_lo;
  assign new_n1107_ = n1122_lo;
  assign new_n1109_ = n1125_lo;
  assign new_n1112_ = ~n1128_lo;
  assign new_n1113_ = n1131_lo;
  assign new_n1115_ = n1134_lo;
  assign new_n1117_ = n1137_lo;
  assign new_n1119_ = n1143_lo;
  assign new_n1121_ = n1146_lo;
  assign new_n1123_ = n1149_lo;
  assign new_n1126_ = ~n1152_lo;
  assign new_n1127_ = n1155_lo;
  assign new_n1130_ = ~n1164_lo;
  assign new_n1131_ = n1167_lo;
  assign new_n1133_ = n1170_lo;
  assign new_n1135_ = n1173_lo;
  assign new_n1138_ = ~n1176_lo;
  assign new_n1140_ = ~n1188_lo;
  assign new_n1142_ = ~n563_inv;
  assign new_n1144_ = ~n1429_o2;
  assign new_n1145_ = n1427_o2;
  assign new_n1148_ = ~n1471_o2;
  assign new_n1150_ = ~n1476_o2;
  assign new_n1151_ = n1499_o2;
  assign new_n1152_ = ~n1499_o2;
  assign new_n1153_ = n1500_o2;
  assign new_n1156_ = ~n1501_o2;
  assign new_n1158_ = ~n1516_o2;
  assign new_n1160_ = ~n1517_o2;
  assign new_n1161_ = n1562_o2;
  assign new_n1162_ = ~n1562_o2;
  assign new_n1164_ = ~n1563_o2;
  assign new_n1165_ = n1564_o2;
  assign new_n1167_ = n1582_o2;
  assign new_n1168_ = ~n1582_o2;
  assign new_n1169_ = n1583_o2;
  assign new_n1170_ = ~n1583_o2;
  assign new_n1171_ = n1618_o2;
  assign new_n1172_ = ~n1618_o2;
  assign new_n1174_ = ~n1622_o2;
  assign new_n1176_ = ~n1502_o2;
  assign new_n1177_ = n1503_o2;
  assign new_n1179_ = n1504_o2;
  assign new_n1181_ = n1505_o2;
  assign new_n1183_ = n1506_o2;
  assign new_n1185_ = n1512_o2;
  assign new_n1186_ = ~n1512_o2;
  assign new_n1187_ = n1513_o2;
  assign new_n1189_ = n1514_o2;
  assign new_n1191_ = n1515_o2;
  assign new_n1194_ = ~n1644_o2;
  assign new_n1196_ = ~n1647_o2;
  assign new_n1197_ = n1527_o2;
  assign new_n1199_ = n650_inv;
  assign new_n1200_ = ~n650_inv;
  assign new_n1201_ = n653_inv;
  assign new_n1203_ = n656_inv;
  assign new_n1206_ = ~n1567_o2;
  assign new_n1207_ = n955_o2;
  assign new_n1208_ = ~n955_o2;
  assign new_n1209_ = n1568_o2;
  assign new_n1212_ = ~n1037_o2;
  assign new_n1213_ = n960_o2;
  assign new_n1215_ = n1587_o2;
  assign new_n1216_ = ~n1587_o2;
  assign new_n1217_ = n1040_o2;
  assign new_n1218_ = ~n1040_o2;
  assign new_n1219_ = n1039_o2;
  assign new_n1220_ = ~n1039_o2;
  assign new_n1221_ = n1589_o2;
  assign new_n1222_ = ~n1589_o2;
  assign new_n1224_ = ~n1624_o2;
  assign new_n1225_ = n1643_o2;
  assign new_n1226_ = ~n1643_o2;
  assign new_n1227_ = n1038_o2;
  assign new_n1228_ = ~n1038_o2;
  assign new_n1229_ = n1645_o2;
  assign new_n1230_ = ~n1645_o2;
  assign new_n1232_ = ~n1029_o2;
  assign new_n1233_ = n701_inv;
  assign new_n1235_ = n1662_o2;
  assign new_n1237_ = n1663_o2;
  assign new_n1239_ = n710_inv;
  assign new_n1242_ = ~n813_o2;
  assign new_n1243_ = lo114_buf_o2;
  assign new_n1244_ = ~lo114_buf_o2;
  assign new_n1245_ = n1031_o2;
  assign new_n1246_ = ~n1031_o2;
  assign new_n1247_ = lo186_buf_o2;
  assign new_n1248_ = ~lo186_buf_o2;
  assign new_n1249_ = n1042_o2;
  assign new_n1250_ = ~n1042_o2;
  assign new_n1251_ = n728_inv;
  assign new_n1253_ = n917_o2;
  assign new_n1255_ = n734_inv;
  assign new_n1257_ = n1649_o2;
  assign new_n1259_ = n1650_o2;
  assign new_n1260_ = ~n1650_o2;
  assign new_n1261_ = n1651_o2;
  assign new_n1263_ = n1652_o2;
  assign new_n1265_ = n1653_o2;
  assign new_n1267_ = lo138_buf_o2;
  assign new_n1269_ = n1664_o2;
  assign new_n1271_ = n1665_o2;
  assign new_n1273_ = n1666_o2;
  assign new_n1275_ = n1667_o2;
  assign new_n1277_ = n944_o2;
  assign new_n1279_ = n770_inv;
  assign new_n1281_ = n1672_o2;
  assign new_n1283_ = n776_inv;
  assign new_n1285_ = n1679_o2;
  assign new_n1287_ = n782_inv;
  assign new_n1288_ = ~n782_inv;
  assign new_n1289_ = n785_inv;
  assign new_n1291_ = lo110_buf_o2;
  assign new_n1292_ = ~lo110_buf_o2;
  assign new_n1293_ = lo134_buf_o2;
  assign new_n1295_ = n1030_o2;
  assign new_n1296_ = ~n1030_o2;
  assign new_n1297_ = lo182_buf_o2;
  assign new_n1298_ = ~lo182_buf_o2;
  assign new_n1300_ = ~n830_o2;
  assign new_n1301_ = n1021_o2;
  assign new_n1302_ = ~n1021_o2;
  assign new_n1303_ = n806_inv;
  assign new_n1305_ = n809_inv;
  assign new_n1307_ = n946_o2;
  assign new_n1309_ = lo038_buf_o2;
  assign new_n1310_ = ~lo038_buf_o2;
  assign new_n1311_ = lo238_buf_o2;
  assign new_n1313_ = n1010_o2;
  assign new_n1314_ = ~n1010_o2;
  assign new_n1315_ = n1006_o2;
  assign new_n1316_ = ~n1006_o2;
  assign new_n1317_ = n907_o2;
  assign new_n1318_ = ~n907_o2;
  assign new_n1320_ = ~n902_o2;
  assign new_n1322_ = ~lo154_buf_o2;
  assign new_n1323_ = n836_inv;
  assign new_n1325_ = n839_inv;
  assign new_n1327_ = lo122_buf_o2;
  assign new_n1329_ = n845_inv;
  assign new_n1330_ = ~n845_inv;
  assign new_n1331_ = n904_o2;
  assign new_n1332_ = ~n904_o2;
  assign new_n1333_ = lo106_buf_o2;
  assign new_n1334_ = ~lo106_buf_o2;
  assign new_n1336_ = ~n980_o2;
  assign new_n1337_ = n1023_o2;
  assign new_n1338_ = ~n1023_o2;
  assign new_n1339_ = lo178_buf_o2;
  assign new_n1340_ = ~lo178_buf_o2;
  assign new_n1342_ = ~n981_o2;
  assign new_n1343_ = n837_o2;
  assign new_n1344_ = ~n837_o2;
  assign new_n1345_ = n1013_o2;
  assign new_n1346_ = ~n1013_o2;
  assign new_n1347_ = n840_o2;
  assign new_n1348_ = ~n840_o2;
  assign new_n1349_ = n849_o2;
  assign new_n1350_ = ~n849_o2;
  assign new_n1351_ = n852_o2;
  assign new_n1352_ = ~n852_o2;
  assign new_n1353_ = n864_o2;
  assign new_n1354_ = ~n864_o2;
  assign new_n1355_ = n867_o2;
  assign new_n1356_ = ~n867_o2;
  assign new_n1357_ = n1044_o2;
  assign new_n1358_ = ~n1044_o2;
  assign new_n1359_ = n876_o2;
  assign new_n1360_ = ~n876_o2;
  assign new_n1361_ = n893_inv;
  assign new_n1363_ = n879_o2;
  assign new_n1364_ = ~n879_o2;
  assign new_n1366_ = ~n925_o2;
  assign new_n1367_ = n902_inv;
  assign new_n1368_ = ~n902_inv;
  assign new_n1369_ = lo146_buf_o2;
  assign new_n1372_ = ~n1026_o2;
  assign new_n1374_ = ~n1032_o2;
  assign new_n1375_ = lo118_buf_o2;
  assign new_n1377_ = n917_inv;
  assign new_n1378_ = ~n917_inv;
  assign new_n1379_ = lo190_buf_o2;
  assign new_n1380_ = ~lo190_buf_o2;
  assign new_n1382_ = ~n1036_o2;
  assign new_n1383_ = n926_inv;
  assign new_n1384_ = ~n926_inv;
  assign new_n1385_ = n929_inv;
  assign new_n1386_ = ~n929_inv;
  assign new_n1387_ = lo002_buf_o2;
  assign new_n1388_ = ~lo002_buf_o2;
  assign new_n1389_ = lo014_buf_o2;
  assign new_n1391_ = lo030_buf_o2;
  assign new_n1393_ = lo034_buf_o2;
  assign new_n1395_ = lo042_buf_o2;
  assign new_n1397_ = lo113_buf_o2;
  assign new_n1398_ = ~lo113_buf_o2;
  assign new_n1399_ = lo185_buf_o2;
  assign new_n1400_ = ~lo185_buf_o2;
  assign new_n1402_ = ~n939_o2;
  assign new_n1404_ = ~n941_o2;
  assign new_n1405_ = lo142_buf_o2;
  assign new_n1406_ = ~lo142_buf_o2;
  assign new_n1407_ = lo230_buf_o2;
  assign new_n1408_ = ~lo230_buf_o2;
  assign new_n1409_ = lo006_buf_o2;
  assign new_n1411_ = lo018_buf_o2;
  assign new_n1413_ = lo022_buf_o2;
  assign new_n1415_ = lo066_buf_o2;
  assign new_n1417_ = n977_inv;
  assign new_n1418_ = ~n977_inv;
  assign new_n1419_ = n826_o2;
  assign new_n1421_ = n892_o2;
  assign new_n1423_ = lo152_buf_o2;
  assign new_n1425_ = n896_o2;
  assign new_n1427_ = n905_o2;
  assign new_n1429_ = n995_inv;
  assign new_n1430_ = ~n995_inv;
  assign new_n1431_ = lo037_buf_o2;
  assign new_n1433_ = lo237_buf_o2;
  assign new_n1434_ = ~lo237_buf_o2;
  assign new_n1435_ = lo062_buf_o2;
  assign new_n1436_ = ~lo062_buf_o2;
  assign new_n1437_ = n1007_inv;
  assign new_n1439_ = n1010_inv;
  assign new_n1441_ = n891_o2;
  assign new_n1443_ = new_n837_ & new_n847_;
  assign new_n1444_ = new_n2116_ | new_n848_;
  assign new_n1445_ = new_n2117_ | new_n2118_;
  assign new_n1446_ = new_n2120_ | new_n1144_;
  assign new_n1447_ = new_n2121_ & new_n1443_;
  assign new_n1448_ = new_n2120_ | new_n2118_;
  assign new_n1449_ = new_n888_ | new_n896_;
  assign new_n1450_ = new_n834_ | new_n1242_;
  assign new_n1451_ = new_n826_ | new_n2122_;
  assign new_n1452_ = new_n836_ | new_n2122_;
  assign new_n1453_ = new_n1447_ | new_n2123_;
  assign new_n1454_ = new_n2124_ | new_n880_;
  assign new_n1455_ = new_n2117_ | new_n2125_;
  assign new_n1456_ = new_n2119_ | new_n2125_;
  assign new_n1457_ = new_n2121_ & new_n1145_;
  assign new_n1458_ = new_n903_ | new_n911_;
  assign new_n1459_ = new_n927_ & new_n2126_;
  assign new_n1460_ = new_n2127_ | new_n2123_;
  assign new_n1461_ = new_n2116_ | new_n2128_;
  assign new_n1462_ = new_n2124_ | new_n876_;
  assign new_n1463_ = new_n2128_ | new_n1462_;
  assign new_n1464_ = new_n919_ & new_n2126_;
  assign new_n1465_ = new_n2129_ & new_n2130_;
  assign new_n1466_ = new_n2131_ | new_n2132_;
  assign new_n1467_ = new_n2131_ & new_n2132_;
  assign new_n1468_ = new_n2129_ | new_n2130_;
  assign new_n1469_ = new_n1466_ & new_n1468_;
  assign new_n1470_ = new_n1465_ | new_n1467_;
  assign new_n1471_ = new_n2134_ & new_n2136_;
  assign new_n1472_ = new_n2138_ | new_n2140_;
  assign new_n1473_ = new_n2138_ & new_n2140_;
  assign new_n1474_ = new_n2134_ | new_n2136_;
  assign new_n1475_ = new_n1472_ & new_n1474_;
  assign new_n1476_ = new_n1471_ | new_n1473_;
  assign new_n1477_ = new_n2141_ & new_n2142_;
  assign new_n1478_ = new_n2143_ | new_n2144_;
  assign new_n1479_ = new_n2143_ & new_n2144_;
  assign new_n1480_ = new_n2141_ | new_n2142_;
  assign new_n1481_ = new_n1478_ & new_n1480_;
  assign new_n1482_ = new_n1477_ | new_n1479_;
  assign new_n1483_ = new_n2145_ & new_n2146_;
  assign new_n1484_ = new_n2147_ | new_n2148_;
  assign new_n1485_ = new_n2147_ & new_n2148_;
  assign new_n1486_ = new_n2145_ | new_n2146_;
  assign new_n1487_ = new_n1484_ & new_n1486_;
  assign new_n1488_ = new_n1483_ | new_n1485_;
  assign new_n1489_ = new_n1476_ & new_n1488_;
  assign new_n1490_ = new_n1475_ & new_n1487_;
  assign new_n1491_ = new_n1489_ | new_n1490_;
  assign new_n1492_ = new_n2149_ & new_n2150_;
  assign new_n1493_ = new_n2151_ | new_n2152_;
  assign new_n1494_ = new_n2151_ & new_n2152_;
  assign new_n1495_ = new_n2149_ | new_n2150_;
  assign new_n1496_ = new_n1493_ & new_n1495_;
  assign new_n1497_ = new_n1492_ | new_n1494_;
  assign new_n1498_ = new_n2135_ & new_n2153_;
  assign new_n1499_ = new_n2139_ | new_n2154_;
  assign new_n1500_ = new_n2139_ & new_n2154_;
  assign new_n1501_ = new_n2135_ | new_n2153_;
  assign new_n1502_ = new_n1499_ & new_n1501_;
  assign new_n1503_ = new_n1498_ | new_n1500_;
  assign new_n1504_ = new_n2155_ & new_n2156_;
  assign new_n1505_ = new_n2157_ | new_n2158_;
  assign new_n1506_ = new_n2157_ & new_n2158_;
  assign new_n1507_ = new_n2155_ | new_n2156_;
  assign new_n1508_ = new_n1505_ & new_n1507_;
  assign new_n1509_ = new_n1504_ | new_n1506_;
  assign new_n1510_ = new_n2159_ & new_n2160_;
  assign new_n1511_ = new_n2161_ | new_n2162_;
  assign new_n1512_ = new_n2161_ & new_n2162_;
  assign new_n1513_ = new_n2159_ | new_n2160_;
  assign new_n1514_ = new_n1511_ & new_n1513_;
  assign new_n1515_ = new_n1510_ | new_n1512_;
  assign new_n1516_ = new_n1503_ & new_n1515_;
  assign new_n1517_ = new_n1502_ & new_n1514_;
  assign new_n1518_ = new_n1516_ | new_n1517_;
  assign new_n1519_ = new_n2165_ & new_n1151_;
  assign new_n1520_ = new_n1150_ | new_n1519_;
  assign new_n1521_ = new_n2173_ | new_n1130_;
  assign new_n1522_ = new_n1520_ & new_n1521_;
  assign new_n1523_ = new_n2173_ | new_n1153_;
  assign new_n1524_ = new_n2182_ & new_n1152_;
  assign new_n1525_ = new_n1523_ & new_n1524_;
  assign new_n1526_ = new_n1522_ | new_n1525_;
  assign new_n1527_ = new_n2189_ | new_n1148_;
  assign new_n1528_ = new_n1056_ | new_n2196_;
  assign new_n1529_ = new_n970_ | new_n2203_;
  assign new_n1530_ = new_n2207_ | new_n1138_;
  assign new_n1531_ = new_n1529_ & new_n1530_;
  assign new_n1532_ = new_n1528_ & new_n1531_;
  assign new_n1533_ = new_n1527_ & new_n1532_;
  assign new_n1534_ = new_n1526_ & new_n1533_;
  assign new_n1535_ = new_n2174_ | new_n1196_;
  assign new_n1536_ = new_n2165_ & new_n1207_;
  assign new_n1537_ = new_n1194_ | new_n1536_;
  assign new_n1538_ = new_n1535_ & new_n1537_;
  assign new_n1539_ = new_n2174_ | new_n1213_;
  assign new_n1540_ = new_n2182_ & new_n1208_;
  assign new_n1541_ = new_n1539_ & new_n1540_;
  assign new_n1542_ = new_n1538_ | new_n1541_;
  assign new_n1543_ = new_n2189_ | new_n1174_;
  assign new_n1544_ = new_n958_ | new_n2203_;
  assign new_n1545_ = new_n1042_ | new_n2196_;
  assign new_n1546_ = new_n1544_ & new_n1545_;
  assign new_n1547_ = new_n1543_ & new_n1546_;
  assign new_n1548_ = new_n1542_ & new_n1547_;
  assign new_n1549_ = new_n2208_ & new_n1171_;
  assign new_n1550_ = new_n1167_ | new_n1172_;
  assign new_n1551_ = new_n1170_ | new_n1549_;
  assign new_n1552_ = new_n1169_ | new_n2209_;
  assign new_n1553_ = new_n1551_ & new_n1552_;
  assign new_n1554_ = new_n2176_ | new_n1553_;
  assign new_n1555_ = new_n2183_ | new_n2209_;
  assign new_n1556_ = new_n2166_ | new_n2208_;
  assign new_n1557_ = new_n2190_ | new_n1164_;
  assign new_n1558_ = new_n1048_ | new_n2197_;
  assign new_n1559_ = new_n1336_ & new_n1342_;
  assign new_n1560_ = new_n1558_ & new_n1559_;
  assign new_n1561_ = new_n1557_ & new_n1560_;
  assign new_n1562_ = new_n1556_ & new_n1561_;
  assign new_n1563_ = new_n1555_ & new_n1562_;
  assign new_n1564_ = new_n1554_ & new_n1563_;
  assign new_n1565_ = new_n2166_ & new_n1161_;
  assign new_n1566_ = new_n1158_ | new_n1565_;
  assign new_n1567_ = new_n2176_ | new_n1160_;
  assign new_n1568_ = new_n1566_ & new_n1567_;
  assign new_n1569_ = new_n2175_ | new_n1165_;
  assign new_n1570_ = new_n2183_ & new_n1162_;
  assign new_n1571_ = new_n1569_ & new_n1570_;
  assign new_n1572_ = new_n1568_ | new_n1571_;
  assign new_n1573_ = new_n2190_ | new_n1156_;
  assign new_n1574_ = new_n1052_ | new_n2197_;
  assign new_n1575_ = new_n966_ | new_n2204_;
  assign new_n1576_ = new_n2207_ | new_n1126_;
  assign new_n1577_ = new_n1575_ & new_n1576_;
  assign new_n1578_ = new_n1574_ & new_n1577_;
  assign new_n1579_ = new_n1573_ & new_n1578_;
  assign new_n1580_ = new_n1572_ & new_n1579_;
  assign new_n1581_ = new_n2210_ & new_n2211_;
  assign new_n1582_ = new_n2213_ | new_n2215_;
  assign new_n1583_ = new_n2213_ & new_n2215_;
  assign new_n1584_ = new_n2210_ | new_n2211_;
  assign new_n1585_ = new_n2216_ & new_n2217_;
  assign new_n1586_ = new_n1019_ | new_n1301_;
  assign new_n1587_ = new_n2219_ & new_n2220_;
  assign new_n1588_ = new_n2221_ | new_n2222_;
  assign new_n1589_ = new_n2223_ & new_n1588_;
  assign new_n1590_ = new_n2224_ | new_n1587_;
  assign new_n1591_ = new_n2225_ | new_n2226_;
  assign new_n1592_ = new_n2228_ & new_n1591_;
  assign new_n1593_ = new_n1217_ & new_n2229_;
  assign new_n1594_ = new_n1218_ | new_n1227_;
  assign new_n1595_ = new_n1220_ | new_n1593_;
  assign new_n1596_ = new_n1219_ | new_n2230_;
  assign new_n1597_ = new_n1595_ & new_n1596_;
  assign new_n1598_ = new_n2178_ | new_n1597_;
  assign new_n1599_ = new_n2185_ | new_n2230_;
  assign new_n1600_ = new_n2168_ | new_n2229_;
  assign new_n1601_ = new_n2192_ | new_n1212_;
  assign new_n1602_ = new_n1036_ | new_n2199_;
  assign new_n1603_ = new_n952_ | new_n2204_;
  assign new_n1604_ = new_n1602_ & new_n1603_;
  assign new_n1605_ = new_n1601_ & new_n1604_;
  assign new_n1606_ = new_n1600_ & new_n1605_;
  assign new_n1607_ = new_n1599_ & new_n1606_;
  assign new_n1608_ = new_n1598_ & new_n1607_;
  assign new_n1609_ = new_n2228_ & new_n1584_;
  assign new_n1610_ = new_n1581_ | new_n2225_;
  assign new_n1611_ = new_n1589_ & new_n1609_;
  assign new_n1612_ = new_n2226_ & new_n2231_;
  assign new_n1613_ = new_n2178_ | new_n1612_;
  assign new_n1614_ = new_n1611_ | new_n1613_;
  assign new_n1615_ = new_n2185_ | new_n2231_;
  assign new_n1616_ = new_n2168_ | new_n2227_;
  assign new_n1617_ = new_n2192_ | new_n2214_;
  assign new_n1618_ = new_n2206_ | new_n1140_;
  assign new_n1619_ = new_n2212_ | new_n2199_;
  assign new_n1620_ = new_n1618_ & new_n1619_;
  assign new_n1621_ = new_n1617_ & new_n1620_;
  assign new_n1622_ = new_n1616_ & new_n1621_;
  assign new_n1623_ = new_n1615_ & new_n1622_;
  assign new_n1624_ = new_n1614_ & new_n1623_;
  assign new_n1625_ = new_n2219_ & new_n2223_;
  assign new_n1626_ = new_n2221_ | new_n2224_;
  assign new_n1627_ = new_n2222_ & new_n1625_;
  assign new_n1628_ = new_n2220_ & new_n2232_;
  assign new_n1629_ = new_n2179_ | new_n1628_;
  assign new_n1630_ = new_n1627_ | new_n1629_;
  assign new_n1631_ = new_n2186_ | new_n2232_;
  assign new_n1632_ = new_n2169_ | new_n2218_;
  assign new_n1633_ = new_n2193_ | new_n2217_;
  assign new_n1634_ = new_n936_ | new_n2206_;
  assign new_n1635_ = new_n2216_ | new_n2200_;
  assign new_n1636_ = new_n1634_ & new_n1635_;
  assign new_n1637_ = new_n1633_ & new_n1636_;
  assign new_n1638_ = new_n1632_ & new_n1637_;
  assign new_n1639_ = new_n1631_ & new_n1638_;
  assign new_n1640_ = new_n1630_ & new_n1639_;
  assign new_n1641_ = new_n1245_ & new_n2233_;
  assign new_n1642_ = new_n1246_ | new_n1295_;
  assign new_n1643_ = new_n1250_ & new_n2234_;
  assign new_n1644_ = new_n1249_ & new_n1641_;
  assign new_n1645_ = new_n2179_ | new_n1644_;
  assign new_n1646_ = new_n1643_ | new_n1645_;
  assign new_n1647_ = new_n2186_ | new_n2234_;
  assign new_n1648_ = new_n2169_ | new_n2233_;
  assign new_n1649_ = new_n2193_ | new_n1232_;
  assign new_n1650_ = new_n944_ | new_n2205_;
  assign new_n1651_ = new_n1028_ | new_n2200_;
  assign new_n1652_ = new_n1650_ & new_n1651_;
  assign new_n1653_ = new_n1649_ & new_n1652_;
  assign new_n1654_ = new_n1648_ & new_n1653_;
  assign new_n1655_ = new_n1647_ & new_n1654_;
  assign new_n1656_ = new_n1646_ & new_n1655_;
  assign new_n1657_ = new_n2235_ | new_n1368_;
  assign new_n1658_ = new_n1374_ & new_n1382_;
  assign new_n1659_ = new_n1378_ | new_n1384_;
  assign new_n1660_ = new_n2237_ & new_n2239_;
  assign new_n1661_ = new_n2240_ & new_n2241_;
  assign new_n1662_ = new_n2237_ | new_n2239_;
  assign new_n1663_ = new_n2242_ | new_n1222_;
  assign new_n1664_ = new_n1224_ | new_n1314_;
  assign new_n1665_ = new_n1316_ & new_n1372_;
  assign new_n1666_ = new_n1664_ & new_n1665_;
  assign new_n1667_ = new_n1663_ & new_n1666_;
  assign new_n1668_ = new_n832_ | new_n1176_;
  assign new_n1669_ = new_n2244_ & new_n2246_;
  assign new_n1670_ = new_n2247_ | new_n2248_;
  assign new_n1671_ = new_n2249_ & new_n1670_;
  assign new_n1672_ = new_n1380_ | new_n1386_;
  assign new_n1673_ = new_n1408_ | new_n1418_;
  assign new_n1674_ = new_n1402_ & new_n1404_;
  assign new_n1675_ = new_n2250_ & new_n2252_;
  assign new_n1676_ = new_n2253_ & new_n2254_;
  assign new_n1677_ = new_n2244_ | new_n2246_;
  assign new_n1678_ = new_n1186_ | new_n1206_;
  assign new_n1679_ = new_n856_ | new_n1678_;
  assign new_n1680_ = new_n2255_ | new_n1679_;
  assign new_n1681_ = new_n2257_ & new_n2258_;
  assign new_n1682_ = new_n1235_ & new_n2259_;
  assign new_n1683_ = new_n1181_ & new_n2260_;
  assign new_n1684_ = new_n2261_ | new_n1683_;
  assign new_n1685_ = new_n1682_ | new_n1684_;
  assign new_n1686_ = new_n1681_ | new_n1685_;
  assign new_n1687_ = new_n2250_ | new_n2252_;
  assign new_n1688_ = new_n1330_ | new_n1398_;
  assign new_n1689_ = new_n1317_ | new_n1406_;
  assign new_n1690_ = new_n1332_ & new_n1689_;
  assign new_n1691_ = new_n1688_ & new_n1690_;
  assign new_n1692_ = new_n2262_ | new_n2263_;
  assign new_n1693_ = new_n1281_ | new_n1310_;
  assign new_n1694_ = new_n1288_ | new_n1693_;
  assign new_n1695_ = new_n1260_ | new_n2264_;
  assign new_n1696_ = new_n1320_ | new_n1695_;
  assign new_n1697_ = new_n1427_ & new_n2266_;
  assign new_n1698_ = new_n1388_ | new_n1697_;
  assign new_n1699_ = new_n2268_ & new_n2269_;
  assign new_n1700_ = new_n2266_ & new_n1699_;
  assign new_n1701_ = new_n2270_ | new_n2272_;
  assign new_n1702_ = new_n2273_ & new_n2274_;
  assign new_n1703_ = new_n2275_ & new_n1441_;
  assign new_n1704_ = new_n2267_ & new_n1703_;
  assign new_n1705_ = new_n1430_ | new_n1436_;
  assign new_n1706_ = new_n1419_ & new_n1425_;
  assign new_n1707_ = new_n1705_ & new_n1706_;
  assign new_n1708_ = new_n1704_ | new_n1707_;
  assign new_n1709_ = new_n2276_ & new_n1434_;
  assign new_n1710_ = new_n2277_ & new_n1709_;
  assign new_n1711_ = new_n2278_ & new_n2279_;
  assign new_n1712_ = new_n2281_ & new_n2282_;
  assign new_n1713_ = new_n2283_ & new_n1117_;
  assign new_n1714_ = new_n2285_ | new_n2257_;
  assign new_n1715_ = new_n934_ | new_n942_;
  assign new_n1716_ = new_n1714_ & new_n1715_;
  assign new_n1717_ = new_n2285_ & new_n2258_;
  assign new_n1718_ = new_n2286_ & new_n2260_;
  assign new_n1719_ = new_n2261_ | new_n1718_;
  assign new_n1720_ = new_n1267_ & new_n2259_;
  assign new_n1721_ = new_n1719_ | new_n1720_;
  assign new_n1722_ = new_n1717_ | new_n1721_;
  assign new_n1723_ = new_n2287_ | new_n2288_;
  assign new_n1724_ = new_n2242_ | new_n1334_;
  assign new_n1725_ = new_n1723_ & new_n1724_;
  assign new_n1726_ = new_n2289_ | new_n2279_;
  assign new_n1727_ = new_n1244_ | new_n1292_;
  assign new_n1728_ = new_n1726_ & new_n1727_;
  assign new_n1729_ = new_n1215_ | new_n2290_;
  assign new_n1730_ = new_n1216_ | new_n1226_;
  assign new_n1731_ = new_n1729_ & new_n1730_;
  assign new_n1732_ = new_n2291_ | new_n2281_;
  assign new_n1733_ = new_n1010_ | new_n1018_;
  assign new_n1734_ = new_n1732_ & new_n1733_;
  assign new_n1735_ = new_n2292_ | new_n2293_;
  assign new_n1736_ = new_n2243_ | new_n2236_;
  assign new_n1737_ = new_n1735_ & new_n1736_;
  assign new_n1738_ = new_n2294_ | new_n2295_;
  assign new_n1739_ = new_n2296_ & new_n1738_;
  assign new_n1740_ = new_n2297_ | new_n2298_;
  assign new_n1741_ = new_n1298_ | new_n2235_;
  assign new_n1742_ = new_n1740_ & new_n1741_;
  assign new_n1743_ = new_n2270_ & new_n2272_;
  assign new_n1744_ = new_n2299_ | new_n2300_;
  assign new_n1745_ = new_n1230_ | new_n1248_;
  assign new_n1746_ = new_n1744_ & new_n1745_;
  assign new_n1747_ = new_n862_ | new_n868_;
  assign new_n1748_ = new_n1200_ | new_n1747_;
  assign new_n1749_ = new_n2301_ | new_n1748_;
  assign new_n1750_ = new_n2302_ & new_n2304_;
  assign new_n1751_ = new_n2305_ & new_n1318_;
  assign new_n1752_ = new_n1331_ | new_n1751_;
  assign new_n1753_ = new_n1750_ | new_n1752_;
  assign new_n1754_ = new_n2306_ & new_n2307_;
  assign new_n1755_ = new_n2308_ & new_n2304_;
  assign new_n1756_ = new_n2309_ | new_n2310_;
  assign new_n1757_ = new_n1322_ | new_n2311_;
  assign new_n1758_ = new_n992_ | new_n1004_;
  assign new_n1759_ = new_n2312_ & new_n1758_;
  assign new_n1760_ = new_n1757_ & new_n1759_;
  assign new_n1761_ = new_n2313_ & new_n2314_;
  assign new_n1762_ = new_n2315_ | new_n1761_;
  assign new_n1763_ = new_n2316_ & new_n2318_;
  assign new_n1764_ = new_n2319_ & new_n2321_;
  assign new_n1765_ = new_n2323_ | new_n1764_;
  assign new_n1766_ = new_n1763_ | new_n1765_;
  assign new_n1767_ = new_n2324_ & new_n2318_;
  assign new_n1768_ = new_n2325_ & new_n2321_;
  assign new_n1769_ = new_n2323_ | new_n1768_;
  assign new_n1770_ = new_n2326_ | new_n2327_;
  assign new_n1771_ = new_n706_ | new_n722_;
  assign new_n1772_ = new_n726_ | new_n784_;
  assign new_n1773_ = new_n2328_ & new_n2330_;
  assign new_n1774_ = new_n2330_ & new_n2332_;
  assign new_n1775_ = new_n2334_ & new_n2335_;
  assign new_n1776_ = new_n714_ | new_n2336_;
  assign new_n1777_ = new_n2337_ & new_n2338_;
  assign new_n1778_ = new_n2331_ & new_n720_;
  assign new_n1779_ = new_n712_ & new_n2334_;
  assign new_n1780_ = new_n1778_ | new_n1779_;
  assign G855 = new_n1445_;
  assign G856 = new_n1446_;
  assign G857 = new_n2127_;
  assign G858 = new_n1449_;
  assign G859 = new_n1451_;
  assign G860 = ~new_n1453_;
  assign G861 = ~new_n1455_;
  assign G862 = ~new_n1456_;
  assign G863 = new_n1457_;
  assign G864 = ~new_n1459_;
  assign G865 = ~new_n1460_;
  assign G866 = new_n1142_;
  assign G867 = new_n1461_;
  assign G868 = new_n1463_;
  assign G869 = ~new_n1464_;
  assign G870 = new_n1491_;
  assign G871 = new_n1518_;
  assign G872 = new_n1534_;
  assign G873 = new_n1548_;
  assign G874 = new_n1564_;
  assign G875 = new_n1580_;
  assign G876 = new_n1592_;
  assign G877 = new_n1608_;
  assign G878 = new_n1624_;
  assign G879 = new_n1640_;
  assign G880 = new_n1656_;
  assign n1654_li007_li007 = new_n2286_;
  assign n1657_li008_li008 = new_n709_;
  assign n1660_li009_li009 = new_n827_;
  assign n1663_li010_li010 = new_n829_;
  assign n1678_li015_li015 = new_n1177_;
  assign n1690_li019_li019 = new_n1187_;
  assign n1702_li023_li023 = new_n1189_;
  assign n1705_li024_li024 = new_n717_;
  assign n1708_li025_li025 = new_n839_;
  assign n1711_li026_li026 = new_n841_;
  assign n1714_li027_li027 = new_n843_;
  assign n1726_li031_li031 = new_n1179_;
  assign n1762_li043_li043 = new_n1183_;
  assign n1765_li044_li044 = new_n727_;
  assign n1768_li045_li045 = new_n851_;
  assign n1771_li046_li046 = new_n853_;
  assign n1777_li048_li048 = new_n729_;
  assign n1780_li049_li049 = new_n857_;
  assign n1783_li050_li050 = new_n859_;
  assign n1789_li052_li052 = new_n731_;
  assign n1792_li053_li053 = new_n863_;
  assign n1795_li054_li054 = new_n865_;
  assign n1801_li056_li056 = new_n733_;
  assign n1804_li057_li057 = new_n869_;
  assign n1807_li058_li058 = new_n871_;
  assign n1810_li059_li059 = new_n873_;
  assign n1822_li063_li063 = new_n1197_;
  assign n1834_li067_li067 = new_n1191_;
  assign n1837_li068_li068 = new_n739_;
  assign n1840_li069_li069 = new_n881_;
  assign n1843_li070_li070 = new_n883_;
  assign n1846_li071_li071 = new_n885_;
  assign n1849_li072_li072 = new_n741_;
  assign n1852_li073_li073 = new_n889_;
  assign n1855_li074_li074 = new_n891_;
  assign n1858_li075_li075 = new_n893_;
  assign n1861_li076_li076 = new_n743_;
  assign n1864_li077_li077 = new_n897_;
  assign n1867_li078_li078 = new_n899_;
  assign n1870_li079_li079 = new_n901_;
  assign n1873_li080_li080 = new_n745_;
  assign n1876_li081_li081 = new_n905_;
  assign n1879_li082_li082 = new_n907_;
  assign n1882_li083_li083 = new_n909_;
  assign n1885_li084_li084 = new_n747_;
  assign n1888_li085_li085 = new_n913_;
  assign n1891_li086_li086 = new_n915_;
  assign n1894_li087_li087 = new_n917_;
  assign n1897_li088_li088 = new_n749_;
  assign n1900_li089_li089 = new_n921_;
  assign n1903_li090_li090 = new_n923_;
  assign n1906_li091_li091 = new_n925_;
  assign n1909_li092_li092 = new_n751_;
  assign n1912_li093_li093 = new_n929_;
  assign n1915_li094_li094 = new_n931_;
  assign n1918_li095_li095 = new_n2284_;
  assign n1921_li096_li096 = new_n753_;
  assign n1924_li097_li097 = new_n937_;
  assign n1927_li098_li098 = new_n939_;
  assign n1930_li099_li099 = new_n2256_;
  assign n1933_li100_li100 = new_n755_;
  assign n1936_li101_li101 = new_n945_;
  assign n1939_li102_li102 = new_n947_;
  assign n1942_li103_li103 = new_n2287_;
  assign n1945_li104_li104 = new_n757_;
  assign n1948_li105_li105 = new_n953_;
  assign n1954_li107_li107 = new_n2288_;
  assign n1957_li108_li108 = new_n759_;
  assign n1960_li109_li109 = new_n959_;
  assign n1969_li112_li112 = new_n761_;
  assign n1978_li115_li115 = new_n2289_;
  assign n1981_li116_li116 = new_n763_;
  assign n1990_li119_li119 = new_n2290_;
  assign n1993_li120_li120 = new_n765_;
  assign n2005_li124_li124 = new_n767_;
  assign n2008_li125_li125 = new_n973_;
  assign n2011_li126_li126 = new_n975_;
  assign n2014_li127_li127 = new_n977_;
  assign n2017_li128_li128 = new_n769_;
  assign n2020_li129_li129 = new_n981_;
  assign n2023_li130_li130 = new_n983_;
  assign n2026_li131_li131 = new_n985_;
  assign n2029_li132_li132 = new_n771_;
  assign n2032_li133_li133 = new_n989_;
  assign n2041_li136_li136 = new_n773_;
  assign n2044_li137_li137 = new_n993_;
  assign n2053_li140_li140 = new_n775_;
  assign n2065_li144_li144 = new_n777_;
  assign n2077_li148_li148 = new_n779_;
  assign n2080_li149_li149 = new_n1001_;
  assign n2113_li160_li160 = new_n785_;
  assign n2116_li161_li161 = new_n1005_;
  assign n2119_li162_li162 = new_n1007_;
  assign n2122_li163_li163 = new_n2291_;
  assign n2125_li164_li164 = new_n787_;
  assign n2128_li165_li165 = new_n1013_;
  assign n2131_li166_li166 = new_n1015_;
  assign n2134_li167_li167 = new_n2280_;
  assign n2137_li168_li168 = new_n789_;
  assign n2140_li169_li169 = new_n1021_;
  assign n2143_li170_li170 = new_n1023_;
  assign n2146_li171_li171 = new_n2292_;
  assign n2149_li172_li172 = new_n791_;
  assign n2152_li173_li173 = new_n1029_;
  assign n2155_li174_li174 = new_n1031_;
  assign n2158_li175_li175 = new_n2293_;
  assign n2161_li176_li176 = new_n793_;
  assign n2164_li177_li177 = new_n1037_;
  assign n2170_li179_li179 = new_n2298_;
  assign n2173_li180_li180 = new_n795_;
  assign n2176_li181_li181 = new_n1043_;
  assign n2182_li183_li183 = new_n2297_;
  assign n2185_li184_li184 = new_n797_;
  assign n2194_li187_li187 = new_n2300_;
  assign n2197_li188_li188 = new_n799_;
  assign n2206_li191_li191 = new_n2299_;
  assign n2209_li192_li192 = new_n801_;
  assign n2212_li193_li193 = new_n1057_;
  assign n2215_li194_li194 = new_n1059_;
  assign n2218_li195_li195 = new_n1061_;
  assign n2221_li196_li196 = new_n803_;
  assign n2224_li197_li197 = new_n1065_;
  assign n2227_li198_li198 = new_n1067_;
  assign n2230_li199_li199 = new_n2278_;
  assign n2233_li200_li200 = new_n805_;
  assign n2236_li201_li201 = new_n1073_;
  assign n2239_li202_li202 = new_n1075_;
  assign n2242_li203_li203 = new_n1077_;
  assign n2245_li204_li204 = new_n807_;
  assign n2248_li205_li205 = new_n1081_;
  assign n2251_li206_li206 = new_n1083_;
  assign n2254_li207_li207 = new_n1085_;
  assign n2257_li208_li208 = new_n809_;
  assign n2260_li209_li209 = new_n1089_;
  assign n2263_li210_li210 = new_n1091_;
  assign n2266_li211_li211 = new_n1093_;
  assign n2269_li212_li212 = new_n811_;
  assign n2272_li213_li213 = new_n1097_;
  assign n2275_li214_li214 = new_n1099_;
  assign n2278_li215_li215 = new_n1101_;
  assign n2281_li216_li216 = new_n813_;
  assign n2284_li217_li217 = new_n1105_;
  assign n2287_li218_li218 = new_n1107_;
  assign n2290_li219_li219 = new_n2283_;
  assign n2293_li220_li220 = new_n815_;
  assign n2296_li221_li221 = new_n1113_;
  assign n2299_li222_li222 = new_n1115_;
  assign n2305_li224_li224 = new_n817_;
  assign n2308_li225_li225 = new_n1119_;
  assign n2311_li226_li226 = new_n1121_;
  assign n2314_li227_li227 = new_n1123_;
  assign n2317_li228_li228 = new_n819_;
  assign n2326_li231_li231 = new_n1237_;
  assign n2329_li232_li232 = new_n821_;
  assign n2332_li233_li233 = new_n1131_;
  assign n2335_li234_li234 = new_n1133_;
  assign n2338_li235_li235 = new_n1135_;
  assign n2350_li239_li239 = new_n1209_;
  assign n1428_i2 = new_n1201_;
  assign n1429_i2 = new_n1203_;
  assign n1427_i2 = new_n1199_;
  assign n1471_i2 = new_n1233_;
  assign n1476_i2 = new_n1239_;
  assign n1499_i2 = new_n1251_;
  assign n1500_i2 = new_n1253_;
  assign n1501_i2 = new_n1255_;
  assign n1516_i2 = new_n1277_;
  assign n1517_i2 = new_n1279_;
  assign n1562_i2 = new_n1303_;
  assign n1563_i2 = new_n1305_;
  assign n1564_i2 = new_n1307_;
  assign n1582_i2 = new_n1323_;
  assign n1583_i2 = new_n1325_;
  assign n1618_i2 = new_n1361_;
  assign n1622_i2 = new_n1367_;
  assign n1502_i2 = new_n1257_;
  assign n1503_i2 = new_n2307_;
  assign n1504_i2 = new_n1261_;
  assign n1505_i2 = new_n1263_;
  assign n1506_i2 = new_n1265_;
  assign n1512_i2 = new_n1269_;
  assign n1513_i2 = new_n1271_;
  assign n1514_i2 = new_n1273_;
  assign n1515_i2 = new_n1275_;
  assign n1644_i2 = new_n1377_;
  assign n1647_i2 = new_n1383_;
  assign n1527_i2 = new_n1285_;
  assign n1526_i2 = new_n1283_;
  assign n1528_i2 = new_n1287_;
  assign n1529_i2 = new_n1289_;
  assign n1567_i2 = new_n1309_;
  assign n955_i2 = ~new_n2240_;
  assign n1568_i2 = new_n2264_;
  assign n1037_i2 = ~new_n2238_;
  assign n960_i2 = ~new_n2241_;
  assign n1587_i2 = new_n1327_;
  assign n1040_i2 = ~new_n2247_;
  assign n1039_i2 = ~new_n2248_;
  assign n1589_i2 = new_n2303_;
  assign n1624_i2 = new_n1369_;
  assign n1643_i2 = new_n1375_;
  assign n1038_i2 = ~new_n2249_;
  assign n1645_i2 = new_n1379_;
  assign n1029_i2 = ~new_n2245_;
  assign n1648_i2 = new_n1385_;
  assign n1662_i2 = new_n1405_;
  assign n1663_i2 = new_n1407_;
  assign n1668_i2 = new_n1417_;
  assign n813_i2 = ~new_n2255_;
  assign lo114_buf_i2 = new_n1397_;
  assign n1031_i2 = ~new_n2294_;
  assign lo186_buf_i2 = new_n1399_;
  assign n1042_i2 = ~new_n2295_;
  assign n911_i2 = ~new_n2253_;
  assign n917_i2 = ~new_n2254_;
  assign n942_i2 = ~new_n2251_;
  assign n1649_i2 = new_n1387_;
  assign n1650_i2 = new_n1389_;
  assign n1651_i2 = new_n1391_;
  assign n1652_i2 = new_n1393_;
  assign n1653_i2 = new_n1395_;
  assign lo138_buf_i2 = new_n2305_;
  assign n1664_i2 = new_n1409_;
  assign n1665_i2 = new_n1411_;
  assign n1666_i2 = new_n1413_;
  assign n1667_i2 = new_n1415_;
  assign n944_i2 = ~new_n2262_;
  assign n945_i2 = ~new_n2263_;
  assign n1672_i2 = new_n2275_;
  assign n1676_i2 = new_n1429_;
  assign n1679_i2 = new_n2268_;
  assign n1680_i2 = new_n2267_;
  assign n1681_i2 = new_n2269_;
  assign lo110_buf_i2 = new_n2302_;
  assign lo134_buf_i2 = new_n2306_;
  assign n1030_i2 = ~new_n2296_;
  assign lo182_buf_i2 = new_n1045_;
  assign n830_i2 = ~new_n2301_;
  assign n1021_i2 = new_n2282_;
  assign n943_i2 = ~new_n2273_;
  assign n936_i2 = ~new_n2271_;
  assign n946_i2 = ~new_n2274_;
  assign lo038_buf_i2 = new_n2276_;
  assign lo238_buf_i2 = new_n1433_;
  assign n1010_i2 = ~new_n2311_;
  assign n1006_i2 = ~new_n2312_;
  assign n907_i2 = ~new_n2320_;
  assign n902_i2 = new_n2277_;
  assign lo154_buf_i2 = new_n2319_;
  assign n938_i2 = ~new_n2313_;
  assign n947_i2 = ~new_n2314_;
  assign lo122_buf_i2 = new_n2316_;
  assign n899_i2 = new_n2317_;
  assign n904_i2 = new_n2322_;
  assign lo106_buf_i2 = new_n2308_;
  assign n980_i2 = new_n1711_;
  assign n1023_i2 = new_n1712_;
  assign lo178_buf_i2 = new_n2309_;
  assign n981_i2 = new_n1713_;
  assign n837_i2 = new_n1716_;
  assign n1013_i2 = new_n1722_;
  assign n840_i2 = new_n1725_;
  assign n849_i2 = new_n1728_;
  assign n852_i2 = new_n1731_;
  assign n864_i2 = new_n1734_;
  assign n867_i2 = new_n1737_;
  assign n1044_i2 = ~new_n1739_;
  assign n876_i2 = new_n1742_;
  assign n937_i2 = ~new_n2315_;
  assign n879_i2 = new_n1746_;
  assign n925_i2 = ~new_n1749_;
  assign n954_i2 = new_n2310_;
  assign lo146_buf_i2 = new_n2325_;
  assign n1026_i2 = new_n1754_;
  assign n1032_i2 = new_n1755_;
  assign lo118_buf_i2 = new_n2324_;
  assign n957_i2 = new_n1756_;
  assign lo190_buf_i2 = new_n2326_;
  assign n1036_i2 = ~new_n1760_;
  assign n949_i2 = ~new_n1762_;
  assign n910_i2 = new_n2327_;
  assign lo002_buf_i2 = new_n705_;
  assign lo014_buf_i2 = new_n2331_;
  assign lo030_buf_i2 = new_n2333_;
  assign lo034_buf_i2 = new_n721_;
  assign lo042_buf_i2 = new_n2335_;
  assign lo113_buf_i2 = new_n963_;
  assign lo185_buf_i2 = new_n1049_;
  assign n939_i2 = new_n1767_;
  assign n941_i2 = new_n1769_;
  assign lo142_buf_i2 = new_n997_;
  assign lo230_buf_i2 = new_n1127_;
  assign lo006_buf_i2 = new_n2328_;
  assign lo018_buf_i2 = new_n713_;
  assign lo022_buf_i2 = new_n2337_;
  assign lo066_buf_i2 = new_n2338_;
  assign n913_i2 = new_n1770_;
  assign n826_i2 = ~new_n2336_;
  assign n892_i2 = ~new_n2332_;
  assign lo152_buf_i2 = new_n781_;
  assign n896_i2 = new_n1773_;
  assign n905_i2 = new_n1774_;
  assign n821_i2 = new_n1775_;
  assign lo037_buf_i2 = new_n723_;
  assign lo237_buf_i2 = new_n823_;
  assign lo062_buf_i2 = new_n735_;
  assign n827_i2 = ~new_n1776_;
  assign n809_i2 = new_n1777_;
  assign n891_i2 = new_n1780_;
  assign new_n2116_ = new_n838_;
  assign new_n2117_ = new_n878_;
  assign new_n2118_ = new_n1444_;
  assign new_n2119_ = new_n846_;
  assign new_n2120_ = new_n2119_;
  assign new_n2121_ = new_n845_;
  assign new_n2122_ = new_n1450_;
  assign new_n2123_ = new_n1452_;
  assign new_n2124_ = new_n850_;
  assign new_n2125_ = new_n1454_;
  assign new_n2126_ = new_n1458_;
  assign new_n2127_ = new_n1448_;
  assign new_n2128_ = new_n1300_;
  assign new_n2129_ = new_n1344_;
  assign new_n2130_ = new_n1348_;
  assign new_n2131_ = new_n1343_;
  assign new_n2132_ = new_n1347_;
  assign new_n2133_ = new_n979_;
  assign new_n2134_ = new_n2133_;
  assign new_n2135_ = new_n2133_;
  assign new_n2136_ = new_n1469_;
  assign new_n2137_ = new_n980_;
  assign new_n2138_ = new_n2137_;
  assign new_n2139_ = new_n2137_;
  assign new_n2140_ = new_n1470_;
  assign new_n2141_ = new_n1350_;
  assign new_n2142_ = new_n1352_;
  assign new_n2143_ = new_n1349_;
  assign new_n2144_ = new_n1351_;
  assign new_n2145_ = new_n987_;
  assign new_n2146_ = new_n1481_;
  assign new_n2147_ = new_n988_;
  assign new_n2148_ = new_n1482_;
  assign new_n2149_ = new_n1354_;
  assign new_n2150_ = new_n1356_;
  assign new_n2151_ = new_n1353_;
  assign new_n2152_ = new_n1355_;
  assign new_n2153_ = new_n1496_;
  assign new_n2154_ = new_n1497_;
  assign new_n2155_ = new_n1360_;
  assign new_n2156_ = new_n1364_;
  assign new_n2157_ = new_n1359_;
  assign new_n2158_ = new_n1363_;
  assign new_n2159_ = new_n1063_;
  assign new_n2160_ = new_n1508_;
  assign new_n2161_ = new_n1064_;
  assign new_n2162_ = new_n1509_;
  assign new_n2163_ = new_n1096_;
  assign new_n2164_ = new_n2163_;
  assign new_n2165_ = new_n2164_;
  assign new_n2166_ = new_n2164_;
  assign new_n2167_ = new_n2163_;
  assign new_n2168_ = new_n2167_;
  assign new_n2169_ = new_n2167_;
  assign new_n2170_ = new_n1080_;
  assign new_n2171_ = new_n2170_;
  assign new_n2172_ = new_n2171_;
  assign new_n2173_ = new_n2172_;
  assign new_n2174_ = new_n2172_;
  assign new_n2175_ = new_n2171_;
  assign new_n2176_ = new_n2175_;
  assign new_n2177_ = new_n2170_;
  assign new_n2178_ = new_n2177_;
  assign new_n2179_ = new_n2177_;
  assign new_n2180_ = new_n1088_;
  assign new_n2181_ = new_n2180_;
  assign new_n2182_ = new_n2181_;
  assign new_n2183_ = new_n2181_;
  assign new_n2184_ = new_n2180_;
  assign new_n2185_ = new_n2184_;
  assign new_n2186_ = new_n2184_;
  assign new_n2187_ = new_n1104_;
  assign new_n2188_ = new_n2187_;
  assign new_n2189_ = new_n2188_;
  assign new_n2190_ = new_n2188_;
  assign new_n2191_ = new_n2187_;
  assign new_n2192_ = new_n2191_;
  assign new_n2193_ = new_n2191_;
  assign new_n2194_ = new_n1366_;
  assign new_n2195_ = new_n2194_;
  assign new_n2196_ = new_n2195_;
  assign new_n2197_ = new_n2195_;
  assign new_n2198_ = new_n2194_;
  assign new_n2199_ = new_n2198_;
  assign new_n2200_ = new_n2198_;
  assign new_n2201_ = new_n1072_;
  assign new_n2202_ = new_n2201_;
  assign new_n2203_ = new_n2202_;
  assign new_n2204_ = new_n2202_;
  assign new_n2205_ = new_n2201_;
  assign new_n2206_ = new_n2205_;
  assign new_n2207_ = new_n1112_;
  assign new_n2208_ = new_n1168_;
  assign new_n2209_ = new_n1550_;
  assign new_n2210_ = new_n1011_;
  assign new_n2211_ = new_n1345_;
  assign new_n2212_ = new_n1012_;
  assign new_n2213_ = new_n2212_;
  assign new_n2214_ = new_n1346_;
  assign new_n2215_ = new_n2214_;
  assign new_n2216_ = new_n1020_;
  assign new_n2217_ = new_n1302_;
  assign new_n2218_ = new_n1338_;
  assign new_n2219_ = new_n2218_;
  assign new_n2220_ = new_n1358_;
  assign new_n2221_ = new_n1337_;
  assign new_n2222_ = new_n1357_;
  assign new_n2223_ = new_n1586_;
  assign new_n2224_ = new_n1585_;
  assign new_n2225_ = new_n1583_;
  assign new_n2226_ = new_n1590_;
  assign new_n2227_ = new_n1582_;
  assign new_n2228_ = new_n2227_;
  assign new_n2229_ = new_n1228_;
  assign new_n2230_ = new_n1594_;
  assign new_n2231_ = new_n1610_;
  assign new_n2232_ = new_n1626_;
  assign new_n2233_ = new_n1296_;
  assign new_n2234_ = new_n1642_;
  assign new_n2235_ = new_n1340_;
  assign new_n2236_ = new_n1034_;
  assign new_n2237_ = new_n2236_;
  assign new_n2238_ = new_n1658_;
  assign new_n2239_ = new_n2238_;
  assign new_n2240_ = new_n1657_;
  assign new_n2241_ = new_n1659_;
  assign new_n2242_ = new_n950_;
  assign new_n2243_ = new_n1026_;
  assign new_n2244_ = new_n2243_;
  assign new_n2245_ = new_n1667_;
  assign new_n2246_ = new_n2245_;
  assign new_n2247_ = new_n1660_;
  assign new_n2248_ = new_n1661_;
  assign new_n2249_ = new_n1662_;
  assign new_n2250_ = new_n1400_;
  assign new_n2251_ = new_n1674_;
  assign new_n2252_ = new_n2251_;
  assign new_n2253_ = new_n1672_;
  assign new_n2254_ = new_n1673_;
  assign new_n2255_ = new_n1668_;
  assign new_n2256_ = new_n941_;
  assign new_n2257_ = new_n2256_;
  assign new_n2258_ = new_n1221_;
  assign new_n2259_ = new_n1313_;
  assign new_n2260_ = new_n1293_;
  assign new_n2261_ = new_n1315_;
  assign new_n2262_ = new_n1675_;
  assign new_n2263_ = new_n1676_;
  assign new_n2264_ = new_n1311_;
  assign new_n2265_ = new_n1437_;
  assign new_n2266_ = new_n2265_;
  assign new_n2267_ = new_n2265_;
  assign new_n2268_ = new_n1435_;
  assign new_n2269_ = new_n1439_;
  assign new_n2270_ = new_n1046_;
  assign new_n2271_ = new_n1691_;
  assign new_n2272_ = new_n2271_;
  assign new_n2273_ = new_n1687_;
  assign new_n2274_ = new_n1692_;
  assign new_n2275_ = new_n1421_;
  assign new_n2276_ = new_n1431_;
  assign new_n2277_ = new_n1700_;
  assign new_n2278_ = new_n1069_;
  assign new_n2279_ = new_n1291_;
  assign new_n2280_ = new_n1017_;
  assign new_n2281_ = new_n2280_;
  assign new_n2282_ = new_n1686_;
  assign new_n2283_ = new_n1109_;
  assign new_n2284_ = new_n933_;
  assign new_n2285_ = new_n2284_;
  assign new_n2286_ = new_n1185_;
  assign new_n2287_ = new_n949_;
  assign new_n2288_ = new_n1333_;
  assign new_n2289_ = new_n1243_;
  assign new_n2290_ = new_n1225_;
  assign new_n2291_ = new_n1009_;
  assign new_n2292_ = new_n1025_;
  assign new_n2293_ = new_n1033_;
  assign new_n2294_ = new_n1669_;
  assign new_n2295_ = new_n1671_;
  assign new_n2296_ = new_n1677_;
  assign new_n2297_ = new_n1297_;
  assign new_n2298_ = new_n1339_;
  assign new_n2299_ = new_n1229_;
  assign new_n2300_ = new_n1247_;
  assign new_n2301_ = new_n1680_;
  assign new_n2302_ = new_n961_;
  assign new_n2303_ = new_n1329_;
  assign new_n2304_ = new_n2303_;
  assign new_n2305_ = new_n995_;
  assign new_n2306_ = new_n991_;
  assign new_n2307_ = new_n1259_;
  assign new_n2308_ = new_n955_;
  assign new_n2309_ = new_n1039_;
  assign new_n2310_ = new_n1753_;
  assign new_n2311_ = new_n1694_;
  assign new_n2312_ = new_n1696_;
  assign new_n2313_ = new_n1701_;
  assign new_n2314_ = new_n1702_;
  assign new_n2315_ = new_n1743_;
  assign new_n2316_ = new_n971_;
  assign new_n2317_ = new_n1708_;
  assign new_n2318_ = new_n2317_;
  assign new_n2319_ = new_n1423_;
  assign new_n2320_ = new_n1698_;
  assign new_n2321_ = new_n2320_;
  assign new_n2322_ = new_n1710_;
  assign new_n2323_ = new_n2322_;
  assign new_n2324_ = new_n967_;
  assign new_n2325_ = new_n999_;
  assign new_n2326_ = new_n1053_;
  assign new_n2327_ = new_n1766_;
  assign new_n2328_ = new_n707_;
  assign new_n2329_ = new_n711_;
  assign new_n2330_ = new_n2329_;
  assign new_n2331_ = new_n2329_;
  assign new_n2332_ = new_n1772_;
  assign new_n2333_ = new_n719_;
  assign new_n2334_ = new_n2333_;
  assign new_n2335_ = new_n725_;
  assign new_n2336_ = new_n1771_;
  assign new_n2337_ = new_n715_;
  assign new_n2338_ = new_n737_;
  always @ (posedge clock) begin
    n492_lo <= n1654_li007_li007;
    n495_lo <= n1657_li008_li008;
    n498_lo <= n1660_li009_li009;
    n501_lo <= n1663_li010_li010;
    n516_lo <= n1678_li015_li015;
    n528_lo <= n1690_li019_li019;
    n540_lo <= n1702_li023_li023;
    n543_lo <= n1705_li024_li024;
    n546_lo <= n1708_li025_li025;
    n549_lo <= n1711_li026_li026;
    n552_lo <= n1714_li027_li027;
    n564_lo <= n1726_li031_li031;
    n600_lo <= n1762_li043_li043;
    n603_lo <= n1765_li044_li044;
    n606_lo <= n1768_li045_li045;
    n609_lo <= n1771_li046_li046;
    n615_lo <= n1777_li048_li048;
    n618_lo <= n1780_li049_li049;
    n621_lo <= n1783_li050_li050;
    n627_lo <= n1789_li052_li052;
    n630_lo <= n1792_li053_li053;
    n633_lo <= n1795_li054_li054;
    n639_lo <= n1801_li056_li056;
    n642_lo <= n1804_li057_li057;
    n645_lo <= n1807_li058_li058;
    n648_lo <= n1810_li059_li059;
    n660_lo <= n1822_li063_li063;
    n672_lo <= n1834_li067_li067;
    n675_lo <= n1837_li068_li068;
    n678_lo <= n1840_li069_li069;
    n681_lo <= n1843_li070_li070;
    n684_lo <= n1846_li071_li071;
    n687_lo <= n1849_li072_li072;
    n690_lo <= n1852_li073_li073;
    n693_lo <= n1855_li074_li074;
    n696_lo <= n1858_li075_li075;
    n699_lo <= n1861_li076_li076;
    n702_lo <= n1864_li077_li077;
    n705_lo <= n1867_li078_li078;
    n708_lo <= n1870_li079_li079;
    n711_lo <= n1873_li080_li080;
    n714_lo <= n1876_li081_li081;
    n717_lo <= n1879_li082_li082;
    n720_lo <= n1882_li083_li083;
    n723_lo <= n1885_li084_li084;
    n726_lo <= n1888_li085_li085;
    n729_lo <= n1891_li086_li086;
    n732_lo <= n1894_li087_li087;
    n735_lo <= n1897_li088_li088;
    n738_lo <= n1900_li089_li089;
    n741_lo <= n1903_li090_li090;
    n744_lo <= n1906_li091_li091;
    n747_lo <= n1909_li092_li092;
    n750_lo <= n1912_li093_li093;
    n753_lo <= n1915_li094_li094;
    n756_lo <= n1918_li095_li095;
    n759_lo <= n1921_li096_li096;
    n762_lo <= n1924_li097_li097;
    n765_lo <= n1927_li098_li098;
    n768_lo <= n1930_li099_li099;
    n771_lo <= n1933_li100_li100;
    n774_lo <= n1936_li101_li101;
    n777_lo <= n1939_li102_li102;
    n780_lo <= n1942_li103_li103;
    n783_lo <= n1945_li104_li104;
    n786_lo <= n1948_li105_li105;
    n792_lo <= n1954_li107_li107;
    n795_lo <= n1957_li108_li108;
    n798_lo <= n1960_li109_li109;
    n807_lo <= n1969_li112_li112;
    n816_lo <= n1978_li115_li115;
    n819_lo <= n1981_li116_li116;
    n828_lo <= n1990_li119_li119;
    n831_lo <= n1993_li120_li120;
    n843_lo <= n2005_li124_li124;
    n846_lo <= n2008_li125_li125;
    n849_lo <= n2011_li126_li126;
    n852_lo <= n2014_li127_li127;
    n855_lo <= n2017_li128_li128;
    n858_lo <= n2020_li129_li129;
    n861_lo <= n2023_li130_li130;
    n864_lo <= n2026_li131_li131;
    n867_lo <= n2029_li132_li132;
    n870_lo <= n2032_li133_li133;
    n879_lo <= n2041_li136_li136;
    n882_lo <= n2044_li137_li137;
    n891_lo <= n2053_li140_li140;
    n903_lo <= n2065_li144_li144;
    n915_lo <= n2077_li148_li148;
    n918_lo <= n2080_li149_li149;
    n951_lo <= n2113_li160_li160;
    n954_lo <= n2116_li161_li161;
    n957_lo <= n2119_li162_li162;
    n960_lo <= n2122_li163_li163;
    n963_lo <= n2125_li164_li164;
    n966_lo <= n2128_li165_li165;
    n969_lo <= n2131_li166_li166;
    n972_lo <= n2134_li167_li167;
    n975_lo <= n2137_li168_li168;
    n978_lo <= n2140_li169_li169;
    n981_lo <= n2143_li170_li170;
    n984_lo <= n2146_li171_li171;
    n987_lo <= n2149_li172_li172;
    n990_lo <= n2152_li173_li173;
    n993_lo <= n2155_li174_li174;
    n996_lo <= n2158_li175_li175;
    n999_lo <= n2161_li176_li176;
    n1002_lo <= n2164_li177_li177;
    n1008_lo <= n2170_li179_li179;
    n1011_lo <= n2173_li180_li180;
    n1014_lo <= n2176_li181_li181;
    n1020_lo <= n2182_li183_li183;
    n1023_lo <= n2185_li184_li184;
    n1032_lo <= n2194_li187_li187;
    n1035_lo <= n2197_li188_li188;
    n1044_lo <= n2206_li191_li191;
    n1047_lo <= n2209_li192_li192;
    n1050_lo <= n2212_li193_li193;
    n1053_lo <= n2215_li194_li194;
    n1056_lo <= n2218_li195_li195;
    n1059_lo <= n2221_li196_li196;
    n1062_lo <= n2224_li197_li197;
    n1065_lo <= n2227_li198_li198;
    n1068_lo <= n2230_li199_li199;
    n1071_lo <= n2233_li200_li200;
    n1074_lo <= n2236_li201_li201;
    n1077_lo <= n2239_li202_li202;
    n1080_lo <= n2242_li203_li203;
    n1083_lo <= n2245_li204_li204;
    n1086_lo <= n2248_li205_li205;
    n1089_lo <= n2251_li206_li206;
    n1092_lo <= n2254_li207_li207;
    n1095_lo <= n2257_li208_li208;
    n1098_lo <= n2260_li209_li209;
    n1101_lo <= n2263_li210_li210;
    n1104_lo <= n2266_li211_li211;
    n1107_lo <= n2269_li212_li212;
    n1110_lo <= n2272_li213_li213;
    n1113_lo <= n2275_li214_li214;
    n1116_lo <= n2278_li215_li215;
    n1119_lo <= n2281_li216_li216;
    n1122_lo <= n2284_li217_li217;
    n1125_lo <= n2287_li218_li218;
    n1128_lo <= n2290_li219_li219;
    n1131_lo <= n2293_li220_li220;
    n1134_lo <= n2296_li221_li221;
    n1137_lo <= n2299_li222_li222;
    n1143_lo <= n2305_li224_li224;
    n1146_lo <= n2308_li225_li225;
    n1149_lo <= n2311_li226_li226;
    n1152_lo <= n2314_li227_li227;
    n1155_lo <= n2317_li228_li228;
    n1164_lo <= n2326_li231_li231;
    n1167_lo <= n2329_li232_li232;
    n1170_lo <= n2332_li233_li233;
    n1173_lo <= n2335_li234_li234;
    n1176_lo <= n2338_li235_li235;
    n1188_lo <= n2350_li239_li239;
    n563_inv <= n1428_i2;
    n1429_o2 <= n1429_i2;
    n1427_o2 <= n1427_i2;
    n1471_o2 <= n1471_i2;
    n1476_o2 <= n1476_i2;
    n1499_o2 <= n1499_i2;
    n1500_o2 <= n1500_i2;
    n1501_o2 <= n1501_i2;
    n1516_o2 <= n1516_i2;
    n1517_o2 <= n1517_i2;
    n1562_o2 <= n1562_i2;
    n1563_o2 <= n1563_i2;
    n1564_o2 <= n1564_i2;
    n1582_o2 <= n1582_i2;
    n1583_o2 <= n1583_i2;
    n1618_o2 <= n1618_i2;
    n1622_o2 <= n1622_i2;
    n1502_o2 <= n1502_i2;
    n1503_o2 <= n1503_i2;
    n1504_o2 <= n1504_i2;
    n1505_o2 <= n1505_i2;
    n1506_o2 <= n1506_i2;
    n1512_o2 <= n1512_i2;
    n1513_o2 <= n1513_i2;
    n1514_o2 <= n1514_i2;
    n1515_o2 <= n1515_i2;
    n1644_o2 <= n1644_i2;
    n1647_o2 <= n1647_i2;
    n1527_o2 <= n1527_i2;
    n650_inv <= n1526_i2;
    n653_inv <= n1528_i2;
    n656_inv <= n1529_i2;
    n1567_o2 <= n1567_i2;
    n955_o2 <= n955_i2;
    n1568_o2 <= n1568_i2;
    n1037_o2 <= n1037_i2;
    n960_o2 <= n960_i2;
    n1587_o2 <= n1587_i2;
    n1040_o2 <= n1040_i2;
    n1039_o2 <= n1039_i2;
    n1589_o2 <= n1589_i2;
    n1624_o2 <= n1624_i2;
    n1643_o2 <= n1643_i2;
    n1038_o2 <= n1038_i2;
    n1645_o2 <= n1645_i2;
    n1029_o2 <= n1029_i2;
    n701_inv <= n1648_i2;
    n1662_o2 <= n1662_i2;
    n1663_o2 <= n1663_i2;
    n710_inv <= n1668_i2;
    n813_o2 <= n813_i2;
    lo114_buf_o2 <= lo114_buf_i2;
    n1031_o2 <= n1031_i2;
    lo186_buf_o2 <= lo186_buf_i2;
    n1042_o2 <= n1042_i2;
    n728_inv <= n911_i2;
    n917_o2 <= n917_i2;
    n734_inv <= n942_i2;
    n1649_o2 <= n1649_i2;
    n1650_o2 <= n1650_i2;
    n1651_o2 <= n1651_i2;
    n1652_o2 <= n1652_i2;
    n1653_o2 <= n1653_i2;
    lo138_buf_o2 <= lo138_buf_i2;
    n1664_o2 <= n1664_i2;
    n1665_o2 <= n1665_i2;
    n1666_o2 <= n1666_i2;
    n1667_o2 <= n1667_i2;
    n944_o2 <= n944_i2;
    n770_inv <= n945_i2;
    n1672_o2 <= n1672_i2;
    n776_inv <= n1676_i2;
    n1679_o2 <= n1679_i2;
    n782_inv <= n1680_i2;
    n785_inv <= n1681_i2;
    lo110_buf_o2 <= lo110_buf_i2;
    lo134_buf_o2 <= lo134_buf_i2;
    n1030_o2 <= n1030_i2;
    lo182_buf_o2 <= lo182_buf_i2;
    n830_o2 <= n830_i2;
    n1021_o2 <= n1021_i2;
    n806_inv <= n943_i2;
    n809_inv <= n936_i2;
    n946_o2 <= n946_i2;
    lo038_buf_o2 <= lo038_buf_i2;
    lo238_buf_o2 <= lo238_buf_i2;
    n1010_o2 <= n1010_i2;
    n1006_o2 <= n1006_i2;
    n907_o2 <= n907_i2;
    n902_o2 <= n902_i2;
    lo154_buf_o2 <= lo154_buf_i2;
    n836_inv <= n938_i2;
    n839_inv <= n947_i2;
    lo122_buf_o2 <= lo122_buf_i2;
    n845_inv <= n899_i2;
    n904_o2 <= n904_i2;
    lo106_buf_o2 <= lo106_buf_i2;
    n980_o2 <= n980_i2;
    n1023_o2 <= n1023_i2;
    lo178_buf_o2 <= lo178_buf_i2;
    n981_o2 <= n981_i2;
    n837_o2 <= n837_i2;
    n1013_o2 <= n1013_i2;
    n840_o2 <= n840_i2;
    n849_o2 <= n849_i2;
    n852_o2 <= n852_i2;
    n864_o2 <= n864_i2;
    n867_o2 <= n867_i2;
    n1044_o2 <= n1044_i2;
    n876_o2 <= n876_i2;
    n893_inv <= n937_i2;
    n879_o2 <= n879_i2;
    n925_o2 <= n925_i2;
    n902_inv <= n954_i2;
    lo146_buf_o2 <= lo146_buf_i2;
    n1026_o2 <= n1026_i2;
    n1032_o2 <= n1032_i2;
    lo118_buf_o2 <= lo118_buf_i2;
    n917_inv <= n957_i2;
    lo190_buf_o2 <= lo190_buf_i2;
    n1036_o2 <= n1036_i2;
    n926_inv <= n949_i2;
    n929_inv <= n910_i2;
    lo002_buf_o2 <= lo002_buf_i2;
    lo014_buf_o2 <= lo014_buf_i2;
    lo030_buf_o2 <= lo030_buf_i2;
    lo034_buf_o2 <= lo034_buf_i2;
    lo042_buf_o2 <= lo042_buf_i2;
    lo113_buf_o2 <= lo113_buf_i2;
    lo185_buf_o2 <= lo185_buf_i2;
    n939_o2 <= n939_i2;
    n941_o2 <= n941_i2;
    lo142_buf_o2 <= lo142_buf_i2;
    lo230_buf_o2 <= lo230_buf_i2;
    lo006_buf_o2 <= lo006_buf_i2;
    lo018_buf_o2 <= lo018_buf_i2;
    lo022_buf_o2 <= lo022_buf_i2;
    lo066_buf_o2 <= lo066_buf_i2;
    n977_inv <= n913_i2;
    n826_o2 <= n826_i2;
    n892_o2 <= n892_i2;
    lo152_buf_o2 <= lo152_buf_i2;
    n896_o2 <= n896_i2;
    n905_o2 <= n905_i2;
    n995_inv <= n821_i2;
    lo037_buf_o2 <= lo037_buf_i2;
    lo237_buf_o2 <= lo237_buf_i2;
    lo062_buf_o2 <= lo062_buf_i2;
    n1007_inv <= n827_i2;
    n1010_inv <= n809_i2;
    n891_o2 <= n891_i2;
  end
  initial begin
    n492_lo <= 1'b0;
    n495_lo <= 1'b0;
    n498_lo <= 1'b0;
    n501_lo <= 1'b0;
    n516_lo <= 1'b0;
    n528_lo <= 1'b0;
    n540_lo <= 1'b0;
    n543_lo <= 1'b0;
    n546_lo <= 1'b0;
    n549_lo <= 1'b0;
    n552_lo <= 1'b0;
    n564_lo <= 1'b0;
    n600_lo <= 1'b0;
    n603_lo <= 1'b0;
    n606_lo <= 1'b0;
    n609_lo <= 1'b0;
    n615_lo <= 1'b0;
    n618_lo <= 1'b0;
    n621_lo <= 1'b0;
    n627_lo <= 1'b0;
    n630_lo <= 1'b0;
    n633_lo <= 1'b0;
    n639_lo <= 1'b0;
    n642_lo <= 1'b0;
    n645_lo <= 1'b0;
    n648_lo <= 1'b0;
    n660_lo <= 1'b0;
    n672_lo <= 1'b0;
    n675_lo <= 1'b0;
    n678_lo <= 1'b0;
    n681_lo <= 1'b0;
    n684_lo <= 1'b0;
    n687_lo <= 1'b0;
    n690_lo <= 1'b0;
    n693_lo <= 1'b0;
    n696_lo <= 1'b0;
    n699_lo <= 1'b0;
    n702_lo <= 1'b0;
    n705_lo <= 1'b0;
    n708_lo <= 1'b0;
    n711_lo <= 1'b0;
    n714_lo <= 1'b0;
    n717_lo <= 1'b0;
    n720_lo <= 1'b0;
    n723_lo <= 1'b0;
    n726_lo <= 1'b0;
    n729_lo <= 1'b0;
    n732_lo <= 1'b0;
    n735_lo <= 1'b0;
    n738_lo <= 1'b0;
    n741_lo <= 1'b0;
    n744_lo <= 1'b0;
    n747_lo <= 1'b0;
    n750_lo <= 1'b0;
    n753_lo <= 1'b0;
    n756_lo <= 1'b0;
    n759_lo <= 1'b0;
    n762_lo <= 1'b0;
    n765_lo <= 1'b0;
    n768_lo <= 1'b0;
    n771_lo <= 1'b0;
    n774_lo <= 1'b0;
    n777_lo <= 1'b0;
    n780_lo <= 1'b0;
    n783_lo <= 1'b0;
    n786_lo <= 1'b0;
    n792_lo <= 1'b0;
    n795_lo <= 1'b0;
    n798_lo <= 1'b0;
    n807_lo <= 1'b0;
    n816_lo <= 1'b0;
    n819_lo <= 1'b0;
    n828_lo <= 1'b0;
    n831_lo <= 1'b0;
    n843_lo <= 1'b0;
    n846_lo <= 1'b0;
    n849_lo <= 1'b0;
    n852_lo <= 1'b0;
    n855_lo <= 1'b0;
    n858_lo <= 1'b0;
    n861_lo <= 1'b0;
    n864_lo <= 1'b0;
    n867_lo <= 1'b0;
    n870_lo <= 1'b0;
    n879_lo <= 1'b0;
    n882_lo <= 1'b0;
    n891_lo <= 1'b0;
    n903_lo <= 1'b0;
    n915_lo <= 1'b0;
    n918_lo <= 1'b0;
    n951_lo <= 1'b0;
    n954_lo <= 1'b0;
    n957_lo <= 1'b0;
    n960_lo <= 1'b0;
    n963_lo <= 1'b0;
    n966_lo <= 1'b0;
    n969_lo <= 1'b0;
    n972_lo <= 1'b0;
    n975_lo <= 1'b0;
    n978_lo <= 1'b0;
    n981_lo <= 1'b0;
    n984_lo <= 1'b0;
    n987_lo <= 1'b0;
    n990_lo <= 1'b0;
    n993_lo <= 1'b0;
    n996_lo <= 1'b0;
    n999_lo <= 1'b0;
    n1002_lo <= 1'b0;
    n1008_lo <= 1'b0;
    n1011_lo <= 1'b0;
    n1014_lo <= 1'b0;
    n1020_lo <= 1'b0;
    n1023_lo <= 1'b0;
    n1032_lo <= 1'b0;
    n1035_lo <= 1'b0;
    n1044_lo <= 1'b0;
    n1047_lo <= 1'b0;
    n1050_lo <= 1'b0;
    n1053_lo <= 1'b0;
    n1056_lo <= 1'b0;
    n1059_lo <= 1'b0;
    n1062_lo <= 1'b0;
    n1065_lo <= 1'b0;
    n1068_lo <= 1'b0;
    n1071_lo <= 1'b0;
    n1074_lo <= 1'b0;
    n1077_lo <= 1'b0;
    n1080_lo <= 1'b0;
    n1083_lo <= 1'b0;
    n1086_lo <= 1'b0;
    n1089_lo <= 1'b0;
    n1092_lo <= 1'b0;
    n1095_lo <= 1'b0;
    n1098_lo <= 1'b0;
    n1101_lo <= 1'b0;
    n1104_lo <= 1'b0;
    n1107_lo <= 1'b0;
    n1110_lo <= 1'b0;
    n1113_lo <= 1'b0;
    n1116_lo <= 1'b0;
    n1119_lo <= 1'b0;
    n1122_lo <= 1'b0;
    n1125_lo <= 1'b0;
    n1128_lo <= 1'b0;
    n1131_lo <= 1'b0;
    n1134_lo <= 1'b0;
    n1137_lo <= 1'b0;
    n1143_lo <= 1'b0;
    n1146_lo <= 1'b0;
    n1149_lo <= 1'b0;
    n1152_lo <= 1'b0;
    n1155_lo <= 1'b0;
    n1164_lo <= 1'b0;
    n1167_lo <= 1'b0;
    n1170_lo <= 1'b0;
    n1173_lo <= 1'b0;
    n1176_lo <= 1'b0;
    n1188_lo <= 1'b0;
    n563_inv <= 1'b0;
    n1429_o2 <= 1'b0;
    n1427_o2 <= 1'b0;
    n1471_o2 <= 1'b0;
    n1476_o2 <= 1'b0;
    n1499_o2 <= 1'b0;
    n1500_o2 <= 1'b0;
    n1501_o2 <= 1'b0;
    n1516_o2 <= 1'b0;
    n1517_o2 <= 1'b0;
    n1562_o2 <= 1'b0;
    n1563_o2 <= 1'b0;
    n1564_o2 <= 1'b0;
    n1582_o2 <= 1'b0;
    n1583_o2 <= 1'b0;
    n1618_o2 <= 1'b0;
    n1622_o2 <= 1'b0;
    n1502_o2 <= 1'b0;
    n1503_o2 <= 1'b0;
    n1504_o2 <= 1'b0;
    n1505_o2 <= 1'b0;
    n1506_o2 <= 1'b0;
    n1512_o2 <= 1'b0;
    n1513_o2 <= 1'b0;
    n1514_o2 <= 1'b0;
    n1515_o2 <= 1'b0;
    n1644_o2 <= 1'b0;
    n1647_o2 <= 1'b0;
    n1527_o2 <= 1'b0;
    n650_inv <= 1'b0;
    n653_inv <= 1'b0;
    n656_inv <= 1'b0;
    n1567_o2 <= 1'b0;
    n955_o2 <= 1'b0;
    n1568_o2 <= 1'b0;
    n1037_o2 <= 1'b0;
    n960_o2 <= 1'b0;
    n1587_o2 <= 1'b0;
    n1040_o2 <= 1'b0;
    n1039_o2 <= 1'b0;
    n1589_o2 <= 1'b0;
    n1624_o2 <= 1'b0;
    n1643_o2 <= 1'b0;
    n1038_o2 <= 1'b0;
    n1645_o2 <= 1'b0;
    n1029_o2 <= 1'b0;
    n701_inv <= 1'b0;
    n1662_o2 <= 1'b0;
    n1663_o2 <= 1'b0;
    n710_inv <= 1'b0;
    n813_o2 <= 1'b0;
    lo114_buf_o2 <= 1'b0;
    n1031_o2 <= 1'b0;
    lo186_buf_o2 <= 1'b0;
    n1042_o2 <= 1'b0;
    n728_inv <= 1'b0;
    n917_o2 <= 1'b0;
    n734_inv <= 1'b0;
    n1649_o2 <= 1'b0;
    n1650_o2 <= 1'b0;
    n1651_o2 <= 1'b0;
    n1652_o2 <= 1'b0;
    n1653_o2 <= 1'b0;
    lo138_buf_o2 <= 1'b0;
    n1664_o2 <= 1'b0;
    n1665_o2 <= 1'b0;
    n1666_o2 <= 1'b0;
    n1667_o2 <= 1'b0;
    n944_o2 <= 1'b0;
    n770_inv <= 1'b0;
    n1672_o2 <= 1'b0;
    n776_inv <= 1'b0;
    n1679_o2 <= 1'b0;
    n782_inv <= 1'b0;
    n785_inv <= 1'b0;
    lo110_buf_o2 <= 1'b0;
    lo134_buf_o2 <= 1'b0;
    n1030_o2 <= 1'b0;
    lo182_buf_o2 <= 1'b0;
    n830_o2 <= 1'b0;
    n1021_o2 <= 1'b0;
    n806_inv <= 1'b0;
    n809_inv <= 1'b0;
    n946_o2 <= 1'b0;
    lo038_buf_o2 <= 1'b0;
    lo238_buf_o2 <= 1'b0;
    n1010_o2 <= 1'b0;
    n1006_o2 <= 1'b0;
    n907_o2 <= 1'b0;
    n902_o2 <= 1'b0;
    lo154_buf_o2 <= 1'b0;
    n836_inv <= 1'b0;
    n839_inv <= 1'b0;
    lo122_buf_o2 <= 1'b0;
    n845_inv <= 1'b0;
    n904_o2 <= 1'b0;
    lo106_buf_o2 <= 1'b0;
    n980_o2 <= 1'b0;
    n1023_o2 <= 1'b0;
    lo178_buf_o2 <= 1'b0;
    n981_o2 <= 1'b0;
    n837_o2 <= 1'b0;
    n1013_o2 <= 1'b0;
    n840_o2 <= 1'b0;
    n849_o2 <= 1'b0;
    n852_o2 <= 1'b0;
    n864_o2 <= 1'b0;
    n867_o2 <= 1'b0;
    n1044_o2 <= 1'b0;
    n876_o2 <= 1'b0;
    n893_inv <= 1'b0;
    n879_o2 <= 1'b0;
    n925_o2 <= 1'b0;
    n902_inv <= 1'b0;
    lo146_buf_o2 <= 1'b0;
    n1026_o2 <= 1'b0;
    n1032_o2 <= 1'b0;
    lo118_buf_o2 <= 1'b0;
    n917_inv <= 1'b0;
    lo190_buf_o2 <= 1'b0;
    n1036_o2 <= 1'b0;
    n926_inv <= 1'b0;
    n929_inv <= 1'b0;
    lo002_buf_o2 <= 1'b0;
    lo014_buf_o2 <= 1'b0;
    lo030_buf_o2 <= 1'b0;
    lo034_buf_o2 <= 1'b0;
    lo042_buf_o2 <= 1'b0;
    lo113_buf_o2 <= 1'b0;
    lo185_buf_o2 <= 1'b0;
    n939_o2 <= 1'b0;
    n941_o2 <= 1'b0;
    lo142_buf_o2 <= 1'b0;
    lo230_buf_o2 <= 1'b0;
    lo006_buf_o2 <= 1'b0;
    lo018_buf_o2 <= 1'b0;
    lo022_buf_o2 <= 1'b0;
    lo066_buf_o2 <= 1'b0;
    n977_inv <= 1'b0;
    n826_o2 <= 1'b0;
    n892_o2 <= 1'b0;
    lo152_buf_o2 <= 1'b0;
    n896_o2 <= 1'b0;
    n905_o2 <= 1'b0;
    n995_inv <= 1'b0;
    lo037_buf_o2 <= 1'b0;
    lo237_buf_o2 <= 1'b0;
    lo062_buf_o2 <= 1'b0;
    n1007_inv <= 1'b0;
    n1010_inv <= 1'b0;
    n891_o2 <= 1'b0;
  end
endmodule


