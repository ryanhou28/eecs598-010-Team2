// Benchmark "mymod" written by ABC on Sun Oct 29 23:44:46 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50,
    G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528,
    G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538,
    G3539, G3540  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50;
  output G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528,
    G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538,
    G3539, G3540;
  reg n1752_lo, n1776_lo, n1824_lo, n1836_lo, n1848_lo, n1860_lo, n1872_lo,
    n1884_lo, n1896_lo, n1908_lo, n1911_lo, n1914_lo, n1923_lo, n1926_lo,
    n1935_lo, n1938_lo, n1947_lo, n1950_lo, n1959_lo, n1962_lo, n1971_lo,
    n1974_lo, n1983_lo, n1995_lo, n2055_lo, n2064_lo, n2067_lo, n2079_lo,
    n2100_lo, n2112_lo, n2124_lo, n2136_lo, n2148_lo, n2160_lo, n2172_lo,
    n2184_lo, n2235_lo, n2238_lo, n2247_lo, n2250_lo, n2259_lo, n2262_lo,
    n2271_lo, n2274_lo, n2283_lo, n2286_lo, n2289_lo, n2295_lo, n2298_lo,
    n2304_lo, n2307_lo, n2316_lo, n2331_lo, n2334_lo, n2337_lo, n2340_lo,
    n2071_o2, n2080_o2, n2137_o2, n2368_o2, n2383_o2, n2405_o2, n2471_o2,
    n2617_o2, n2765_o2, n2775_o2, n2829_o2, n2579_o2, n2580_o2, n2618_o2,
    n2619_o2, n2620_o2, n2621_o2, n2622_o2, n2623_o2, n2624_o2, n2625_o2,
    n2626_o2, n2627_o2, n3029_o2, n3035_o2, n2643_o2, n2644_o2, n2645_o2,
    n327_inv, n2658_o2, n2659_o2, n2674_o2, n2675_o2, n2676_o2, n3119_o2,
    n3153_o2, n351_inv, n2729_o2, n2730_o2, n2731_o2, n698_o2, n366_inv,
    n2757_o2, n2758_o2, n1000_o2, n1160_o2, n1153_o2, n2793_o2, n2794_o2,
    n2795_o2, n1001_o2, n2859_o2, n744_o2, n402_inv, n2926_o2, n408_inv,
    n2966_o2, n2967_o2, n2947_o2, n1010_o2, n2976_o2, n3069_o2, n3028_o2,
    n3081_o2, n3082_o2, n3142_o2, n3214_o2, n2992_o2, n2993_o2, n870_o2,
    n3086_o2, n3087_o2, n3088_o2, n3089_o2, n3090_o2, n3091_o2, n3092_o2,
    n3093_o2, n3094_o2, n3095_o2, n483_inv, n3170_o2, n3171_o2, n3172_o2,
    n3179_o2, n498_inv, n3193_o2, n3211_o2, n3212_o2, n3213_o2, n513_inv,
    n1125_o2, n1081_o2, n1139_o2, n3245_o2, n3246_o2, n3247_o2,
    lo074_buf_o2, lo078_buf_o2, lo186_buf_o2, lo118_buf_o2, lo146_buf_o2,
    n1038_o2, n1044_o2, n555_inv, n558_inv, lo026_buf_o2, lo030_buf_o2,
    lo090_buf_o2, lo094_buf_o2, lo098_buf_o2, lo102_buf_o2, lo066_buf_o2,
    lo070_buf_o2, n1202_o2, n1003_o2, n1031_o2, n1034_o2, n1040_o2,
    n1046_o2, n1380_o2, n1425_o2, n697_o2, n1143_o2, n673_o2, n789_o2,
    n786_o2, n1047_o2, n1036_o2, n1307_o2, n1035_o2, n1297_o2, n1099_o2,
    n1128_o2, n645_inv, n826_o2, n853_o2, n654_inv, n700_o2, n884_o2,
    lo082_buf_o2, lo086_buf_o2, n801_o2, n840_o2, n675_inv, lo002_buf_o2,
    lo010_buf_o2, lo166_buf_o2, lo170_buf_o2, n1426_o2, n1082_o2, n1310_o2,
    n1015_o2, n1206_o2, n1262_o2, n1456_o2, n1244_o2, n1280_o2, n1290_o2,
    n1012_o2, n1074_o2, n1112_o2, n1212_o2, n1454_o2, n1182_o2, n1220_o2,
    n701_o2, n744_inv, n1282_o2, n1144_o2, n1278_o2, n1459_o2, n1324_o2,
    n1288_o2, n1271_o2, n1132_o2, n1231_o2, n1462_o2, n1482_o2, n994_o2,
    n998_o2, lo106_buf_o2, n769_o2, n814_o2, n841_o2, n867_o2,
    lo006_buf_o2, lo014_buf_o2, lo022_buf_o2, lo042_buf_o2, lo046_buf_o2,
    lo050_buf_o2, lo054_buf_o2, lo130_buf_o2, lo134_buf_o2, lo154_buf_o2,
    lo174_buf_o2, lo178_buf_o2, n1007_o2, n1294_o2, n1084_o2, n1399_o2,
    n1311_o2, n1392_o2, n1102_o2, n1041_o2, n1298_o2, n738_o2, n1214_o2,
    n1222_o2, n1155_o2, n1147_o2, n1393_o2, n999_o2, n1306_o2, n1312_o2,
    n1382_o2, n1383_o2, n1152_o2, n1334_o2, n1335_o2, n906_inv, n773_o2,
    lo190_buf_o2, n1368_o2, n1362_o2, n1406_o2, n1403_o2, n741_o2,
    n1407_o2, n1395_o2, n1359_o2, n1159_o2, n1221_o2, n945_inv, n989_o2,
    n881_o2, n1340_o2, n1341_o2, n906_o2, n1388_o2, n791_o2, n1372_o2,
    n815_o2, n868_o2, lo018_buf_o2, lo138_buf_o2, lo158_buf_o2, n780_o2,
    n728_o2, n993_inv, n929_o2, n955_o2, n938_o2, n1117_o2, n1121_o2,
    n965_o2, n752_o2, n753_o2, n760_o2, n770_o2, n923_o2, n947_o2, n897_o2,
    n919_o2, n895_o2, n917_o2, n751_o2, n774_o2, lo126_buf_o2,
    lo142_buf_o2, lo162_buf_o2, n1059_inv, n792_o2, n869_o2, n1068_inv,
    lo024_buf_o2, lo028_buf_o2, lo088_buf_o2, lo092_buf_o2, lo096_buf_o2,
    lo100_buf_o2, n763_o2, n754_o2, n755_o2, n822_o2, n849_o2, n777_o2,
    n778_o2, n820_o2, n846_o2, n806_o2, n771_o2, n854_o2, n828_o2,
    lo117_buf_o2, lo145_buf_o2, n762_o2, n805_o2, n859_o2, n833_o2,
    lo034_buf_o2, lo038_buf_o2, lo122_buf_o2, lo150_buf_o2;
  wire new_new_n795__, new_new_n796__, new_new_n797__, new_new_n798__,
    new_new_n799__, new_new_n800__, new_new_n801__, new_new_n802__,
    new_new_n803__, new_new_n805__, new_new_n807__, new_new_n809__,
    new_new_n811__, new_new_n813__, new_new_n815__, new_new_n817__,
    new_new_n818__, new_new_n819__, new_new_n820__, new_new_n821__,
    new_new_n823__, new_new_n825__, new_new_n827__, new_new_n829__,
    new_new_n831__, new_new_n833__, new_new_n835__, new_new_n837__,
    new_new_n839__, new_new_n841__, new_new_n843__, new_new_n845__,
    new_new_n847__, new_new_n849__, new_new_n851__, new_new_n853__,
    new_new_n855__, new_new_n857__, new_new_n858__, new_new_n859__,
    new_new_n860__, new_new_n861__, new_new_n862__, new_new_n863__,
    new_new_n865__, new_new_n866__, new_new_n867__, new_new_n869__,
    new_new_n871__, new_new_n872__, new_new_n873__, new_new_n875__,
    new_new_n877__, new_new_n879__, new_new_n881__, new_new_n883__,
    new_new_n885__, new_new_n887__, new_new_n889__, new_new_n891__,
    new_new_n893__, new_new_n896__, new_new_n897__, new_new_n898__,
    new_new_n899__, new_new_n900__, new_new_n901__, new_new_n903__,
    new_new_n904__, new_new_n905__, new_new_n906__, new_new_n907__,
    new_new_n908__, new_new_n909__, new_new_n910__, new_new_n911__,
    new_new_n912__, new_new_n913__, new_new_n914__, new_new_n915__,
    new_new_n917__, new_new_n919__, new_new_n921__, new_new_n923__,
    new_new_n925__, new_new_n927__, new_new_n929__, new_new_n931__,
    new_new_n933__, new_new_n935__, new_new_n937__, new_new_n938__,
    new_new_n939__, new_new_n941__, new_new_n943__, new_new_n944__,
    new_new_n945__, new_new_n946__, new_new_n947__, new_new_n949__,
    new_new_n951__, new_new_n952__, new_new_n953__, new_new_n954__,
    new_new_n955__, new_new_n956__, new_new_n957__, new_new_n958__,
    new_new_n959__, new_new_n960__, new_new_n961__, new_new_n962__,
    new_new_n963__, new_new_n964__, new_new_n965__, new_new_n966__,
    new_new_n967__, new_new_n969__, new_new_n970__, new_new_n971__,
    new_new_n973__, new_new_n975__, new_new_n977__, new_new_n979__,
    new_new_n981__, new_new_n983__, new_new_n985__, new_new_n988__,
    new_new_n989__, new_new_n991__, new_new_n992__, new_new_n993__,
    new_new_n994__, new_new_n995__, new_new_n996__, new_new_n997__,
    new_new_n998__, new_new_n999__, new_new_n1001__, new_new_n1003__,
    new_new_n1005__, new_new_n1006__, new_new_n1007__, new_new_n1008__,
    new_new_n1009__, new_new_n1010__, new_new_n1012__, new_new_n1014__,
    new_new_n1016__, new_new_n1017__, new_new_n1018__, new_new_n1019__,
    new_new_n1021__, new_new_n1023__, new_new_n1025__, new_new_n1026__,
    new_new_n1027__, new_new_n1029__, new_new_n1030__, new_new_n1031__,
    new_new_n1032__, new_new_n1033__, new_new_n1035__, new_new_n1036__,
    new_new_n1037__, new_new_n1038__, new_new_n1039__, new_new_n1040__,
    new_new_n1041__, new_new_n1042__, new_new_n1043__, new_new_n1044__,
    new_new_n1045__, new_new_n1046__, new_new_n1047__, new_new_n1049__,
    new_new_n1051__, new_new_n1052__, new_new_n1053__, new_new_n1055__,
    new_new_n1056__, new_new_n1057__, new_new_n1058__, new_new_n1059__,
    new_new_n1061__, new_new_n1062__, new_new_n1063__, new_new_n1064__,
    new_new_n1065__, new_new_n1068__, new_new_n1069__, new_new_n1071__,
    new_new_n1073__, new_new_n1074__, new_new_n1075__, new_new_n1076__,
    new_new_n1077__, new_new_n1079__, new_new_n1081__, new_new_n1082__,
    new_new_n1083__, new_new_n1084__, new_new_n1085__, new_new_n1087__,
    new_new_n1088__, new_new_n1090__, new_new_n1091__, new_new_n1093__,
    new_new_n1095__, new_new_n1097__, new_new_n1098__, new_new_n1099__,
    new_new_n1100__, new_new_n1101__, new_new_n1102__, new_new_n1103__,
    new_new_n1104__, new_new_n1105__, new_new_n1106__, new_new_n1107__,
    new_new_n1108__, new_new_n1110__, new_new_n1111__, new_new_n1112__,
    new_new_n1113__, new_new_n1115__, new_new_n1116__, new_new_n1117__,
    new_new_n1119__, new_new_n1121__, new_new_n1123__, new_new_n1125__,
    new_new_n1126__, new_new_n1127__, new_new_n1128__, new_new_n1129__,
    new_new_n1131__, new_new_n1132__, new_new_n1133__, new_new_n1134__,
    new_new_n1135__, new_new_n1136__, new_new_n1137__, new_new_n1139__,
    new_new_n1140__, new_new_n1141__, new_new_n1143__, new_new_n1144__,
    new_new_n1145__, new_new_n1147__, new_new_n1149__, new_new_n1150__,
    new_new_n1151__, new_new_n1153__, new_new_n1154__, new_new_n1155__,
    new_new_n1156__, new_new_n1157__, new_new_n1158__, new_new_n1159__,
    new_new_n1160__, new_new_n1161__, new_new_n1163__, new_new_n1165__,
    new_new_n1167__, new_new_n1169__, new_new_n1171__, new_new_n1173__,
    new_new_n1174__, new_new_n1175__, new_new_n1177__, new_new_n1180__,
    new_new_n1181__, new_new_n1183__, new_new_n1185__, new_new_n1187__,
    new_new_n1189__, new_new_n1190__, new_new_n1191__, new_new_n1192__,
    new_new_n1194__, new_new_n1195__, new_new_n1196__, new_new_n1197__,
    new_new_n1198__, new_new_n1199__, new_new_n1201__, new_new_n1202__,
    new_new_n1203__, new_new_n1204__, new_new_n1205__, new_new_n1206__,
    new_new_n1207__, new_new_n1209__, new_new_n1211__, new_new_n1212__,
    new_new_n1213__, new_new_n1214__, new_new_n1215__, new_new_n1217__,
    new_new_n1219__, new_new_n1220__, new_new_n1221__, new_new_n1222__,
    new_new_n1223__, new_new_n1225__, new_new_n1226__, new_new_n1227__,
    new_new_n1228__, new_new_n1229__, new_new_n1230__, new_new_n1231__,
    new_new_n1233__, new_new_n1236__, new_new_n1237__, new_new_n1238__,
    new_new_n1239__, new_new_n1240__, new_new_n1241__, new_new_n1242__,
    new_new_n1243__, new_new_n1244__, new_new_n1245__, new_new_n1246__,
    new_new_n1247__, new_new_n1249__, new_new_n1251__, new_new_n1254__,
    new_new_n1255__, new_new_n1257__, new_new_n1258__, new_new_n1259__,
    new_new_n1260__, new_new_n1261__, new_new_n1263__, new_new_n1265__,
    new_new_n1267__, new_new_n1269__, new_new_n1272__, new_new_n1273__,
    new_new_n1274__, new_new_n1275__, new_new_n1277__, new_new_n1279__,
    new_new_n1281__, new_new_n1283__, new_new_n1285__, new_new_n1286__,
    new_new_n1287__, new_new_n1288__, new_new_n1289__, new_new_n1290__,
    new_new_n1291__, new_new_n1292__, new_new_n1293__, new_new_n1294__,
    new_new_n1295__, new_new_n1296__, new_new_n1297__, new_new_n1298__,
    new_new_n1299__, new_new_n1300__, new_new_n1301__, new_new_n1302__,
    new_new_n1303__, new_new_n1304__, new_new_n1305__, new_new_n1306__,
    new_new_n1307__, new_new_n1308__, new_new_n1310__, new_new_n1311__,
    new_new_n1312__, new_new_n1313__, new_new_n1316__, new_new_n1317__,
    new_new_n1318__, new_new_n1319__, new_new_n1320__, new_new_n1321__,
    new_new_n1322__, new_new_n1323__, new_new_n1324__, new_new_n1325__,
    new_new_n1326__, new_new_n1327__, new_new_n1328__, new_new_n1329__,
    new_new_n1330__, new_new_n1331__, new_new_n1332__, new_new_n1333__,
    new_new_n1334__, new_new_n1335__, new_new_n1336__, new_new_n1337__,
    new_new_n1338__, new_new_n1339__, new_new_n1341__, new_new_n1343__,
    new_new_n1344__, new_new_n1345__, new_new_n1347__, new_new_n1348__,
    new_new_n1349__, new_new_n1350__, new_new_n1351__, new_new_n1352__,
    new_new_n1353__, new_new_n1354__, new_new_n1356__, new_new_n1357__,
    new_new_n1358__, new_new_n1359__, new_new_n1360__, new_new_n1361__,
    new_new_n1362__, new_new_n1363__, new_new_n1364__, new_new_n1365__,
    new_new_n1366__, new_new_n1367__, new_new_n1368__, new_new_n1369__,
    new_new_n1371__, new_new_n1372__, new_new_n1373__, new_new_n1374__,
    new_new_n1375__, new_new_n1376__, new_new_n1377__, new_new_n1379__,
    new_new_n1381__, new_new_n1382__, new_new_n1383__, new_new_n1384__,
    new_new_n1385__, new_new_n1386__, new_new_n1387__, new_new_n1388__,
    new_new_n1389__, new_new_n1390__, new_new_n1391__, new_new_n1392__,
    new_new_n1393__, new_new_n1394__, new_new_n1395__, new_new_n1397__,
    new_new_n1398__, new_new_n1399__, new_new_n1400__, new_new_n1401__,
    new_new_n1402__, new_new_n1403__, new_new_n1404__, new_new_n1406__,
    new_new_n1408__, new_new_n1410__, new_new_n1411__, new_new_n1414__,
    new_new_n1415__, new_new_n1416__, new_new_n1417__, new_new_n1418__,
    new_new_n1420__, new_new_n1421__, new_new_n1422__, new_new_n1423__,
    new_new_n1424__, new_new_n1425__, new_new_n1426__, new_new_n1427__,
    new_new_n1428__, new_new_n1429__, new_new_n1430__, new_new_n1431__,
    new_new_n1433__, new_new_n1434__, new_new_n1435__, new_new_n1437__,
    new_new_n1439__, new_new_n1440__, new_new_n1441__, new_new_n1442__,
    new_new_n1443__, new_new_n1444__, new_new_n1445__, new_new_n1446__,
    new_new_n1447__, new_new_n1448__, new_new_n1449__, new_new_n1451__,
    new_new_n1452__, new_new_n1453__, new_new_n1456__, new_new_n1458__,
    new_new_n1460__, new_new_n1462__, new_new_n1463__, new_new_n1464__,
    new_new_n1466__, new_new_n1467__, new_new_n1469__, new_new_n1471__,
    new_new_n1472__, new_new_n1473__, new_new_n1474__, new_new_n1475__,
    new_new_n1476__, new_new_n1477__, new_new_n1478__, new_new_n1479__,
    new_new_n1480__, new_new_n1481__, new_new_n1482__, new_new_n1483__,
    new_new_n1484__, new_new_n1485__, new_new_n1486__, new_new_n1487__,
    new_new_n1489__, new_new_n1490__, new_new_n1492__, new_new_n1493__,
    new_new_n1494__, new_new_n1495__, new_new_n1496__, new_new_n1497__,
    new_new_n1498__, new_new_n1499__, new_new_n1500__, new_new_n1501__,
    new_new_n1503__, new_new_n1504__, new_new_n1505__, new_new_n1507__,
    new_new_n1509__, new_new_n1510__, new_new_n1511__, new_new_n1512__,
    new_new_n1513__, new_new_n1514__, new_new_n1515__, new_new_n1516__,
    new_new_n1517__, new_new_n1518__, new_new_n1519__, new_new_n1520__,
    new_new_n1521__, new_new_n1523__, new_new_n1524__, new_new_n1525__,
    new_new_n1526__, new_new_n1527__, new_new_n1529__, new_new_n1530__,
    new_new_n1531__, new_new_n1532__, new_new_n1533__, new_new_n1534__,
    new_new_n1535__, new_new_n1536__, new_new_n1537__, new_new_n1538__,
    new_new_n1539__, new_new_n1540__, new_new_n1541__, new_new_n1542__,
    new_new_n1543__, new_new_n1544__, new_new_n1545__, new_new_n1546__,
    new_new_n1547__, new_new_n1548__, new_new_n1549__, new_new_n1551__,
    new_new_n1552__, new_new_n1553__, new_new_n1554__, new_new_n1555__,
    new_new_n1556__, new_new_n1557__, new_new_n1559__, new_new_n1560__,
    new_new_n1561__, new_new_n1562__, new_new_n1563__, new_new_n1564__,
    new_new_n1565__, new_new_n1566__, new_new_n1567__, new_new_n1569__,
    new_new_n1571__, new_new_n1572__, new_new_n1573__, new_new_n1574__,
    new_new_n1575__, new_new_n1576__, new_new_n1577__, new_new_n1578__,
    new_new_n1579__, new_new_n1580__, new_new_n1581__, new_new_n1582__,
    new_new_n1583__, new_new_n1584__, new_new_n1585__, new_new_n1586__,
    new_new_n1587__, new_new_n1588__, new_new_n1589__, new_new_n1590__,
    new_new_n1591__, new_new_n1592__, new_new_n1593__, new_new_n1594__,
    new_new_n1595__, new_new_n1596__, new_new_n1597__, new_new_n1598__,
    new_new_n1599__, new_new_n1600__, new_new_n1601__, new_new_n1602__,
    new_new_n1603__, new_new_n1604__, new_new_n1605__, new_new_n1606__,
    new_new_n1607__, new_new_n1608__, new_new_n1609__, new_new_n1610__,
    new_new_n1611__, new_new_n1612__, new_new_n1613__, new_new_n1614__,
    new_new_n1615__, new_new_n1616__, new_new_n1617__, new_new_n1618__,
    new_new_n1619__, new_new_n1620__, new_new_n1621__, new_new_n1622__,
    new_new_n1623__, new_new_n1624__, new_new_n1625__, new_new_n1626__,
    new_new_n1627__, new_new_n1628__, new_new_n1629__, new_new_n1630__,
    new_new_n1631__, new_new_n1632__, new_new_n1633__, new_new_n1634__,
    new_new_n1635__, new_new_n1636__, new_new_n1637__, new_new_n1638__,
    new_new_n1639__, new_new_n1640__, new_new_n1641__, new_new_n1642__,
    new_new_n1643__, new_new_n1644__, new_new_n1645__, new_new_n1646__,
    new_new_n1647__, new_new_n1648__, new_new_n1649__, new_new_n1650__,
    new_new_n1651__, new_new_n1652__, new_new_n1653__, new_new_n1654__,
    new_new_n1655__, new_new_n1656__, new_new_n1657__, new_new_n1658__,
    new_new_n1659__, new_new_n1660__, new_new_n1661__, new_new_n1662__,
    new_new_n1663__, new_new_n1664__, new_new_n1665__, new_new_n1666__,
    new_new_n1667__, new_new_n1668__, new_new_n1669__, new_new_n1670__,
    new_new_n1671__, new_new_n1672__, new_new_n1673__, new_new_n1674__,
    new_new_n1675__, new_new_n1676__, new_new_n1677__, new_new_n1678__,
    new_new_n1679__, new_new_n1680__, new_new_n1681__, new_new_n1682__,
    new_new_n1683__, new_new_n1684__, new_new_n1685__, new_new_n1686__,
    new_new_n1687__, new_new_n1688__, new_new_n1689__, new_new_n1690__,
    new_new_n1691__, new_new_n1692__, new_new_n1693__, new_new_n1694__,
    new_new_n1695__, new_new_n1696__, new_new_n1697__, new_new_n1698__,
    new_new_n1699__, new_new_n1700__, new_new_n1701__, new_new_n1702__,
    new_new_n1703__, new_new_n1704__, new_new_n1705__, new_new_n1706__,
    new_new_n1707__, new_new_n1708__, new_new_n1709__, new_new_n1710__,
    new_new_n1711__, new_new_n1712__, new_new_n1713__, new_new_n1714__,
    new_new_n1715__, new_new_n1716__, new_new_n1717__, new_new_n1718__,
    new_new_n1719__, new_new_n1720__, new_new_n1721__, new_new_n1722__,
    new_new_n1723__, new_new_n1724__, new_new_n1725__, new_new_n1726__,
    new_new_n1727__, new_new_n1728__, new_new_n1729__, new_new_n1730__,
    new_new_n1731__, new_new_n1732__, new_new_n1733__, new_new_n1734__,
    new_new_n1735__, new_new_n1736__, new_new_n1737__, new_new_n1738__,
    new_new_n1739__, new_new_n1740__, new_new_n1741__, new_new_n1742__,
    new_new_n1743__, new_new_n1744__, new_new_n1745__, new_new_n1746__,
    new_new_n1747__, new_new_n1748__, new_new_n1749__, new_new_n1750__,
    new_new_n1751__, new_new_n1752__, new_new_n1753__, new_new_n1754__,
    new_new_n1755__, new_new_n1756__, new_new_n1757__, new_new_n1758__,
    new_new_n1759__, new_new_n1760__, new_new_n1761__, new_new_n1762__,
    new_new_n1763__, new_new_n1764__, new_new_n1765__, new_new_n1766__,
    new_new_n1767__, new_new_n1768__, new_new_n1769__, new_new_n1770__,
    new_new_n1771__, new_new_n1772__, new_new_n1773__, new_new_n1774__,
    new_new_n1775__, new_new_n1776__, new_new_n1777__, new_new_n1778__,
    new_new_n1779__, new_new_n1780__, new_new_n1781__, new_new_n1782__,
    new_new_n1783__, new_new_n1784__, new_new_n1785__, new_new_n1786__,
    new_new_n1787__, new_new_n1788__, new_new_n1789__, new_new_n1790__,
    new_new_n1791__, new_new_n1792__, new_new_n1793__, new_new_n1794__,
    new_new_n1795__, new_new_n1796__, new_new_n1797__, new_new_n1798__,
    new_new_n1799__, new_new_n1800__, new_new_n1801__, new_new_n1802__,
    new_new_n1803__, new_new_n1804__, new_new_n1805__, new_new_n1806__,
    new_new_n1807__, new_new_n1808__, new_new_n1809__, new_new_n1810__,
    new_new_n1811__, new_new_n1812__, new_new_n1813__, new_new_n1814__,
    new_new_n1815__, new_new_n1816__, new_new_n1817__, new_new_n1818__,
    new_new_n1819__, new_new_n1820__, new_new_n1821__, new_new_n1822__,
    new_new_n1823__, new_new_n1824__, new_new_n1825__, new_new_n1826__,
    new_new_n1827__, new_new_n1828__, new_new_n1829__, new_new_n1830__,
    new_new_n1831__, new_new_n1832__, new_new_n1833__, new_new_n1834__,
    new_new_n1835__, new_new_n1836__, new_new_n1837__, new_new_n1838__,
    new_new_n1839__, new_new_n1840__, new_new_n1841__, new_new_n1842__,
    new_new_n1843__, new_new_n1844__, new_new_n1845__, new_new_n1846__,
    new_new_n1847__, new_new_n1848__, new_new_n1849__, new_new_n1850__,
    new_new_n1851__, new_new_n1852__, new_new_n1853__, new_new_n1854__,
    new_new_n1855__, new_new_n1856__, new_new_n1857__, new_new_n1858__,
    new_new_n1859__, new_new_n1860__, new_new_n1861__, new_new_n1862__,
    new_new_n1863__, new_new_n1864__, new_new_n1865__, new_new_n1866__,
    new_new_n1867__, new_new_n1868__, new_new_n1869__, new_new_n1870__,
    new_new_n1871__, new_new_n1872__, new_new_n1873__, new_new_n1874__,
    new_new_n1875__, new_new_n1876__, new_new_n1877__, new_new_n1878__,
    new_new_n1879__, new_new_n1880__, new_new_n1881__, new_new_n1882__,
    new_new_n1883__, new_new_n1884__, new_new_n1885__, new_new_n1886__,
    new_new_n1887__, new_new_n1888__, new_new_n1889__, new_new_n1890__,
    new_new_n1891__, new_new_n1892__, new_new_n1893__, new_new_n1894__,
    new_new_n1895__, new_new_n1896__, new_new_n1897__, new_new_n1898__,
    new_new_n1899__, new_new_n1900__, new_new_n1901__, new_new_n1902__,
    new_new_n1903__, new_new_n1904__, new_new_n1905__, new_new_n1906__,
    new_new_n1907__, new_new_n1908__, new_new_n1909__, new_new_n1910__,
    new_new_n1911__, new_new_n1912__, new_new_n1913__, new_new_n1914__,
    new_new_n1915__, new_new_n1916__, new_new_n1917__, new_new_n1918__,
    new_new_n1919__, new_new_n1920__, new_new_n1921__, new_new_n1922__,
    new_new_n1923__, new_new_n1924__, new_new_n1925__, new_new_n1926__,
    new_new_n1927__, new_new_n1928__, new_new_n1929__, new_new_n1930__,
    new_new_n1931__, new_new_n1932__, new_new_n1933__, new_new_n1934__,
    new_new_n1935__, new_new_n1936__, new_new_n1937__, new_new_n1938__,
    new_new_n1939__, new_new_n1940__, new_new_n1941__, new_new_n1942__,
    new_new_n1943__, new_new_n1944__, new_new_n1945__, new_new_n1946__,
    new_new_n1947__, new_new_n1948__, new_new_n1949__, new_new_n1950__,
    new_new_n1951__, new_new_n1952__, new_new_n1953__, new_new_n1954__,
    new_new_n1955__, new_new_n1956__, new_new_n1957__, new_new_n1958__,
    new_new_n1959__, new_new_n1960__, new_new_n1961__, new_new_n1962__,
    new_new_n1963__, new_new_n1964__, new_new_n1965__, new_new_n1966__,
    new_new_n1967__, new_new_n1968__, new_new_n1969__, new_new_n1970__,
    new_new_n1971__, new_new_n1972__, new_new_n1973__, new_new_n1974__,
    new_new_n1975__, new_new_n1976__, new_new_n1977__, new_new_n1978__,
    new_new_n1979__, new_new_n1980__, new_new_n1981__, new_new_n1982__,
    new_new_n1983__, new_new_n1984__, new_new_n1985__, new_new_n1986__,
    new_new_n1987__, new_new_n1988__, new_new_n1989__, new_new_n1990__,
    new_new_n1991__, new_new_n1992__, new_new_n1993__, new_new_n1994__,
    new_new_n1995__, new_new_n1996__, new_new_n1997__, new_new_n1998__,
    new_new_n1999__, new_new_n2000__, new_new_n2001__, new_new_n2002__,
    new_new_n2003__, new_new_n2004__, new_new_n2005__, new_new_n2006__,
    new_new_n2007__, new_new_n2008__, new_new_n2009__, new_new_n2010__,
    new_new_n2011__, new_new_n2012__, new_new_n2013__, new_new_n2014__,
    new_new_n2015__, new_new_n2016__, new_new_n2017__, new_new_n2018__,
    new_new_n2019__, new_new_n2020__, new_new_n2021__, new_new_n2022__,
    new_new_n2023__, new_new_n2024__, new_new_n2025__, new_new_n2026__,
    new_new_n2027__, new_new_n2028__, new_new_n2029__, new_new_n2030__,
    new_new_n2031__, new_new_n2032__, new_new_n2033__, new_new_n2034__,
    new_new_n2035__, new_new_n2036__, new_new_n2037__, new_new_n2038__,
    new_new_n2039__, new_new_n2040__, new_new_n2041__, new_new_n2042__,
    new_new_n2043__, new_new_n2044__, new_new_n2045__, new_new_n2046__,
    new_new_n2047__, new_new_n2048__, new_new_n2049__, new_new_n2050__,
    new_new_n2051__, new_new_n2052__, new_new_n2053__, new_new_n2054__,
    new_new_n2055__, new_new_n2056__, new_new_n2057__, new_new_n2058__,
    new_new_n2059__, new_new_n2060__, new_new_n2061__, new_new_n2062__,
    new_new_n2063__, new_new_n2064__, new_new_n2065__, new_new_n2066__,
    new_new_n2067__, new_new_n2068__, new_new_n2069__, new_new_n2070__,
    new_new_n2071__, new_new_n2072__, new_new_n2073__, new_new_n2074__,
    new_new_n2075__, new_new_n2076__, new_new_n2077__, new_new_n2078__,
    new_new_n2079__, new_new_n2080__, new_new_n2081__, new_new_n2082__,
    new_new_n2083__, new_new_n2084__, new_new_n2085__, new_new_n2086__,
    new_new_n2087__, new_new_n2088__, new_new_n2089__, new_new_n2090__,
    new_new_n2091__, new_new_n2092__, new_new_n2093__, new_new_n2094__,
    new_new_n2095__, new_new_n2096__, new_new_n2097__, new_new_n2098__,
    new_new_n2099__, new_new_n2100__, new_new_n2101__, new_new_n2102__,
    new_new_n2103__, new_new_n2104__, new_new_n2105__, new_new_n2106__,
    new_new_n2107__, new_new_n2108__, new_new_n2109__, new_new_n2110__,
    new_new_n2111__, new_new_n2112__, new_new_n2113__, new_new_n2114__,
    new_new_n2115__, new_new_n2116__, new_new_n2117__, new_new_n2118__,
    new_new_n2119__, new_new_n2120__, new_new_n2121__, new_new_n2122__,
    new_new_n2123__, new_new_n2124__, new_new_n2125__, new_new_n2126__,
    new_new_n2127__, new_new_n2128__, new_new_n2129__, new_new_n2130__,
    new_new_n2131__, new_new_n2132__, new_new_n2133__, new_new_n2134__,
    new_new_n2135__, new_new_n2136__, new_new_n2137__, new_new_n2138__,
    new_new_n2139__, new_new_n2140__, new_new_n2141__, new_new_n2142__,
    new_new_n2143__, new_new_n2144__, new_new_n2145__, new_new_n2146__,
    new_new_n2147__, new_new_n2148__, new_new_n2149__, new_new_n2150__,
    new_new_n2151__, new_new_n2152__, new_new_n2153__, new_new_n2154__,
    new_new_n2155__, new_new_n2156__, new_new_n2157__, new_new_n2158__,
    new_new_n2159__, new_new_n2160__, new_new_n2161__, new_new_n2162__,
    new_new_n2163__, new_new_n2164__, new_new_n2165__, new_new_n2166__,
    new_new_n2167__, new_new_n2168__, new_new_n2169__, new_new_n2170__,
    new_new_n2171__, new_new_n2172__, new_new_n2173__, new_new_n2174__,
    new_new_n2175__, new_new_n2176__, new_new_n2177__, new_new_n2178__,
    new_new_n2179__, new_new_n2180__, new_new_n2181__, new_new_n2182__,
    new_new_n2183__, new_new_n2184__, new_new_n2185__, new_new_n2186__,
    new_new_n2187__, new_new_n2188__, new_new_n2189__, new_new_n2190__,
    new_new_n2191__, new_new_n2192__, new_new_n2193__, new_new_n2194__,
    new_new_n2195__, new_new_n2196__, new_new_n2197__, new_new_n2198__,
    new_new_n2199__, new_new_n2200__, new_new_n2201__, new_new_n2202__,
    new_new_n2203__, new_new_n2204__, new_new_n2205__, new_new_n2206__,
    new_new_n2207__, new_new_n2208__, new_new_n2209__, new_new_n2210__,
    new_new_n2211__, new_new_n2212__, new_new_n2213__, new_new_n2214__,
    new_new_n2215__, new_new_n2216__, new_new_n2217__, new_new_n2218__,
    new_new_n2219__, new_new_n2220__, new_new_n2221__, new_new_n2222__,
    new_new_n2223__, new_new_n2224__, new_new_n2225__, new_new_n2226__,
    new_new_n2227__, new_new_n2228__, new_new_n2229__, new_new_n2230__,
    new_new_n2231__, new_new_n2232__, new_new_n2233__, new_new_n2234__,
    new_new_n2235__, new_new_n2236__, new_new_n2237__, new_new_n2238__,
    new_new_n2239__, new_new_n2240__, new_new_n2241__, new_new_n2242__,
    new_new_n2243__, new_new_n2244__, new_new_n2245__, new_new_n2246__,
    new_new_n2247__, new_new_n2248__, new_new_n2249__, new_new_n2250__,
    new_new_n2251__, new_new_n2252__, new_new_n2253__, new_new_n2254__,
    new_new_n2255__, new_new_n2256__, new_new_n2257__, new_new_n2258__,
    new_new_n2259__, new_new_n2260__, new_new_n2261__, new_new_n2262__,
    new_new_n2263__, new_new_n2264__, new_new_n2265__, new_new_n2266__,
    new_new_n2267__, new_new_n2268__, new_new_n2269__, new_new_n2270__,
    new_new_n2271__, new_new_n2272__, new_new_n2273__, new_new_n2274__,
    new_new_n2275__, new_new_n2276__, new_new_n2277__, new_new_n2278__,
    new_new_n2279__, new_new_n2280__, new_new_n2281__, new_new_n2282__,
    new_new_n2283__, new_new_n2284__, new_new_n2285__, new_new_n2286__,
    new_new_n2287__, new_new_n2288__, new_new_n2289__, new_new_n2290__,
    new_new_n2291__, new_new_n2292__, new_new_n2293__, new_new_n2294__,
    new_new_n2295__, new_new_n2296__, new_new_n2297__, new_new_n2298__,
    new_new_n2299__, new_new_n2300__, new_new_n2301__, new_new_n2302__,
    new_new_n2303__, new_new_n2304__, new_new_n2305__, new_new_n2306__,
    new_new_n2307__, new_new_n2308__, new_new_n2309__, new_new_n2310__,
    new_new_n2311__, new_new_n2312__, new_new_n2313__, new_new_n2314__,
    new_new_n2315__, new_new_n2316__, new_new_n2317__, new_new_n2318__,
    new_new_n2319__, new_new_n2320__, new_new_n2321__, new_new_n2322__,
    new_new_n2323__, new_new_n2324__, new_new_n2325__, new_new_n2326__,
    new_new_n2327__, new_new_n2328__, new_new_n2329__, new_new_n2330__,
    new_new_n2331__, new_new_n2332__, new_new_n2333__, new_new_n2334__,
    new_new_n2335__, new_new_n2336__, new_new_n2337__, new_new_n2338__,
    new_new_n2339__, new_new_n2340__, new_new_n2341__, new_new_n2342__,
    new_new_n2343__, new_new_n2344__, new_new_n2345__, new_new_n2346__,
    new_new_n2347__, new_new_n2348__, new_new_n2349__, new_new_n2350__,
    new_new_n2351__, new_new_n2352__, new_new_n2353__, new_new_n2354__,
    new_new_n2355__, new_new_n2356__, new_new_n2357__, new_new_n2358__,
    new_new_n2359__, new_new_n2360__, new_new_n2361__, new_new_n2362__,
    new_new_n2363__, new_new_n2364__, new_new_n2365__, new_new_n2366__,
    new_new_n2367__, new_new_n2368__, new_new_n2369__, new_new_n2370__,
    new_new_n2371__, new_new_n2372__, new_new_n2373__, new_new_n2374__,
    new_new_n2375__, new_new_n2376__, new_new_n2377__, new_new_n2378__,
    new_new_n2379__, new_new_n2380__, new_new_n2381__, new_new_n2382__,
    new_new_n2383__, new_new_n2384__, new_new_n2385__, new_new_n2386__,
    new_new_n2387__, new_new_n2388__, new_new_n2389__, new_new_n2390__,
    new_new_n2391__, new_new_n2392__, new_new_n2393__, new_new_n2394__,
    new_new_n2395__, new_new_n2396__, new_new_n2397__, new_new_n2398__,
    new_new_n2399__, new_new_n2400__, new_new_n2401__, new_new_n2402__,
    new_new_n2403__, new_new_n2404__, new_new_n2405__, new_new_n2406__,
    new_new_n2407__, new_new_n2408__, new_new_n2409__, new_new_n2410__,
    new_new_n2411__, new_new_n2412__, new_new_n2413__, new_new_n2414__,
    new_new_n2415__, new_new_n2416__, new_new_n2417__, new_new_n2418__,
    new_new_n2419__, new_new_n2420__, new_new_n2421__, new_new_n2422__,
    new_new_n2423__, new_new_n2424__, new_new_n2425__, new_new_n2426__,
    new_new_n2427__, new_new_n2428__, new_new_n2429__, new_new_n2430__,
    new_new_n2431__, new_new_n2432__, new_new_n2433__, new_new_n2434__,
    new_new_n2435__, new_new_n2436__, new_new_n2437__, new_new_n2438__,
    new_new_n2439__, new_new_n2440__, new_new_n2441__, new_new_n2442__,
    new_new_n2443__, new_new_n2444__, new_new_n2445__, new_new_n2446__,
    new_new_n2447__, new_new_n2448__, new_new_n2449__, new_new_n2450__,
    new_new_n2451__, new_new_n2452__, new_new_n2453__, new_new_n2454__,
    new_new_n2455__, new_new_n2456__, new_new_n2457__, new_new_n2458__,
    new_new_n2459__, new_new_n2460__, new_new_n2461__, new_new_n2462__,
    new_new_n2463__, new_new_n2464__, new_new_n2465__, new_new_n2466__,
    new_new_n2467__, new_new_n2468__, new_new_n2469__, new_new_n2470__,
    new_new_n2471__, new_new_n2472__, new_new_n2473__, new_new_n2474__,
    new_new_n2475__, new_new_n2476__, new_new_n2477__, new_new_n2478__,
    new_new_n2479__, new_new_n2480__, new_new_n2481__, new_new_n2482__,
    new_new_n2483__, new_new_n2484__, new_new_n2485__, new_new_n2486__,
    new_new_n2487__, new_new_n2488__, new_new_n2489__, new_new_n2490__,
    new_new_n2491__, new_new_n2492__, new_new_n2493__, new_new_n2494__,
    new_new_n2495__, new_new_n2496__, new_new_n2497__, new_new_n2498__,
    new_new_n2499__, new_new_n2500__, new_new_n2501__, new_new_n2502__,
    new_new_n2503__, new_new_n2504__, new_new_n2505__, new_new_n2506__,
    new_new_n2507__, new_new_n2508__, new_new_n2509__, new_new_n2510__,
    new_new_n2511__, new_new_n2512__, new_new_n2513__, new_new_n2514__,
    new_new_n2515__, new_new_n2516__, new_new_n2517__, new_new_n2518__,
    new_new_n2519__, new_new_n2520__, new_new_n2521__, new_new_n2522__,
    new_new_n2523__, new_new_n2524__, new_new_n2525__, new_new_n2526__,
    new_new_n2527__, new_new_n2528__, new_new_n2529__, new_new_n2530__,
    new_new_n2531__, new_new_n2532__, new_new_n2533__, new_new_n2534__,
    new_new_n2535__, new_new_n2536__, new_new_n2537__, new_new_n2538__,
    new_new_n2539__, new_new_n2540__, new_new_n2541__, new_new_n2542__,
    new_new_n2543__, new_new_n2544__, new_new_n2545__, new_new_n2546__,
    new_new_n2547__, new_new_n2548__, new_new_n2549__, new_new_n2550__,
    new_new_n2551__, new_new_n2552__, new_new_n2553__, new_new_n2554__,
    new_new_n2555__, new_new_n2556__, new_new_n2557__, new_new_n2558__,
    new_new_n2559__, new_new_n2560__, new_new_n2561__, new_new_n2562__,
    new_new_n2563__, new_new_n2564__, new_new_n2565__, new_new_n2566__,
    new_new_n2567__, new_new_n2568__, new_new_n2569__, new_new_n2570__,
    new_new_n2571__, new_new_n2572__, new_new_n2573__, new_new_n2574__,
    new_new_n2575__, new_new_n2576__, new_new_n2577__, new_new_n2578__,
    new_new_n2579__, new_new_n2580__, new_new_n2581__, new_new_n2582__,
    new_new_n2583__, new_new_n2584__, new_new_n2585__, new_new_n2586__,
    new_new_n2587__, new_new_n2588__, new_new_n2589__, new_new_n2590__,
    new_new_n2591__, new_new_n2592__, new_new_n2593__, new_new_n2594__,
    new_new_n2595__, new_new_n2596__, new_new_n2597__, new_new_n2598__,
    new_new_n2599__, new_new_n2600__, new_new_n2601__, new_new_n2602__,
    new_new_n2603__, new_new_n2604__, new_new_n2605__, new_new_n2606__,
    new_new_n2607__, new_new_n2608__, new_new_n2609__, new_new_n2610__,
    new_new_n2611__, new_new_n2612__, new_new_n2613__, new_new_n2614__,
    new_new_n2615__, new_new_n2616__, new_new_n2617__, new_new_n2618__,
    new_new_n2619__, new_new_n2620__, new_new_n2621__, new_new_n2622__,
    new_new_n2623__, new_new_n2624__, new_new_n2625__, new_new_n2626__,
    new_new_n2627__, new_new_n2628__, new_new_n2629__, new_new_n2630__,
    new_new_n2631__, new_new_n2632__, new_new_n2633__, new_new_n2634__,
    new_new_n2635__, new_new_n2636__, new_new_n2637__, new_new_n2638__,
    new_new_n2639__, new_new_n2640__, new_new_n2641__, new_new_n2642__,
    new_new_n2643__, new_new_n2644__, new_new_n2645__, new_new_n2646__,
    new_new_n2647__, new_new_n2648__, new_new_n2649__, new_new_n2650__,
    new_new_n2651__, new_new_n2652__, new_new_n2653__, new_new_n2654__,
    new_new_n2655__, new_new_n2656__, new_new_n2657__, new_new_n2658__,
    new_new_n2659__, new_new_n2660__, new_new_n2661__, new_new_n2662__,
    new_new_n2663__, new_new_n2664__, new_new_n2665__, new_new_n2666__,
    new_new_n2667__, new_new_n2668__, new_new_n2669__, new_new_n2670__,
    new_new_n2671__, new_new_n2672__, new_new_n2673__, new_new_n2674__,
    new_new_n2675__, new_new_n2676__, new_new_n2677__, new_new_n2678__,
    new_new_n2679__, new_new_n3063__, new_new_n3064__, new_new_n3065__,
    new_new_n3066__, new_new_n3067__, new_new_n3068__, new_new_n3069__,
    new_new_n3070__, new_new_n3071__, new_new_n3072__, new_new_n3073__,
    new_new_n3074__, new_new_n3075__, new_new_n3076__, new_new_n3077__,
    new_new_n3078__, new_new_n3079__, new_new_n3080__, new_new_n3081__,
    new_new_n3082__, new_new_n3083__, new_new_n3084__, new_new_n3085__,
    new_new_n3086__, new_new_n3087__, new_new_n3088__, new_new_n3089__,
    new_new_n3090__, new_new_n3091__, new_new_n3092__, new_new_n3093__,
    new_new_n3094__, new_new_n3095__, new_new_n3096__, new_new_n3097__,
    new_new_n3098__, new_new_n3099__, new_new_n3100__, new_new_n3101__,
    new_new_n3102__, new_new_n3103__, new_new_n3104__, new_new_n3105__,
    new_new_n3106__, new_new_n3107__, new_new_n3108__, new_new_n3109__,
    new_new_n3110__, new_new_n3111__, new_new_n3112__, new_new_n3113__,
    new_new_n3114__, new_new_n3115__, new_new_n3116__, new_new_n3117__,
    new_new_n3118__, new_new_n3119__, new_new_n3120__, new_new_n3121__,
    new_new_n3122__, new_new_n3123__, new_new_n3124__, new_new_n3125__,
    new_new_n3126__, new_new_n3127__, new_new_n3128__, new_new_n3129__,
    new_new_n3130__, new_new_n3131__, new_new_n3132__, new_new_n3133__,
    new_new_n3134__, new_new_n3135__, new_new_n3136__, new_new_n3137__,
    new_new_n3138__, new_new_n3139__, new_new_n3140__, new_new_n3141__,
    new_new_n3142__, new_new_n3143__, new_new_n3144__, new_new_n3145__,
    new_new_n3146__, new_new_n3147__, new_new_n3148__, new_new_n3149__,
    new_new_n3150__, new_new_n3151__, new_new_n3152__, new_new_n3153__,
    new_new_n3154__, new_new_n3155__, new_new_n3156__, new_new_n3157__,
    new_new_n3158__, new_new_n3159__, new_new_n3160__, new_new_n3161__,
    new_new_n3162__, new_new_n3163__, new_new_n3164__, new_new_n3165__,
    new_new_n3166__, new_new_n3167__, new_new_n3168__, new_new_n3169__,
    new_new_n3170__, new_new_n3171__, new_new_n3172__, new_new_n3173__,
    new_new_n3174__, new_new_n3175__, new_new_n3176__, new_new_n3177__,
    new_new_n3178__, new_new_n3179__, new_new_n3180__, new_new_n3181__,
    new_new_n3182__, new_new_n3183__, new_new_n3184__, new_new_n3185__,
    new_new_n3186__, new_new_n3187__, new_new_n3188__, new_new_n3189__,
    new_new_n3190__, new_new_n3191__, new_new_n3192__, new_new_n3193__,
    new_new_n3194__, new_new_n3195__, new_new_n3196__, new_new_n3197__,
    new_new_n3198__, new_new_n3199__, new_new_n3200__, new_new_n3201__,
    new_new_n3202__, new_new_n3203__, new_new_n3204__, new_new_n3205__,
    new_new_n3206__, new_new_n3207__, new_new_n3208__, new_new_n3209__,
    new_new_n3210__, new_new_n3211__, new_new_n3212__, new_new_n3213__,
    new_new_n3214__, new_new_n3215__, new_new_n3216__, new_new_n3217__,
    new_new_n3218__, new_new_n3219__, new_new_n3220__, new_new_n3221__,
    new_new_n3222__, new_new_n3223__, new_new_n3224__, new_new_n3225__,
    new_new_n3226__, new_new_n3227__, new_new_n3228__, new_new_n3229__,
    new_new_n3230__, new_new_n3231__, new_new_n3232__, new_new_n3233__,
    new_new_n3234__, new_new_n3235__, new_new_n3236__, new_new_n3237__,
    new_new_n3238__, new_new_n3239__, new_new_n3240__, new_new_n3241__,
    new_new_n3242__, new_new_n3243__, new_new_n3244__, new_new_n3245__,
    new_new_n3246__, new_new_n3247__, new_new_n3248__, new_new_n3249__,
    new_new_n3250__, new_new_n3251__, new_new_n3252__, new_new_n3253__,
    new_new_n3254__, new_new_n3255__, new_new_n3256__, new_new_n3257__,
    new_new_n3258__, new_new_n3259__, new_new_n3260__, new_new_n3261__,
    new_new_n3262__, new_new_n3263__, new_new_n3264__, new_new_n3265__,
    new_new_n3266__, new_new_n3267__, new_new_n3268__, new_new_n3269__,
    new_new_n3270__, new_new_n3271__, new_new_n3272__, new_new_n3273__,
    new_new_n3274__, new_new_n3275__, new_new_n3276__, new_new_n3277__,
    new_new_n3278__, new_new_n3279__, new_new_n3280__, new_new_n3281__,
    new_new_n3282__, new_new_n3283__, new_new_n3284__, new_new_n3285__,
    new_new_n3286__, new_new_n3287__, new_new_n3288__, new_new_n3289__,
    new_new_n3290__, new_new_n3291__, new_new_n3292__, new_new_n3293__,
    new_new_n3294__, new_new_n3295__, new_new_n3296__, new_new_n3297__,
    new_new_n3298__, new_new_n3299__, new_new_n3300__, new_new_n3301__,
    new_new_n3302__, new_new_n3303__, new_new_n3304__, new_new_n3305__,
    new_new_n3306__, new_new_n3307__, new_new_n3308__, new_new_n3309__,
    new_new_n3310__, new_new_n3311__, new_new_n3312__, new_new_n3313__,
    new_new_n3314__, new_new_n3315__, new_new_n3316__, new_new_n3317__,
    new_new_n3318__, new_new_n3319__, new_new_n3320__, new_new_n3321__,
    new_new_n3322__, new_new_n3323__, new_new_n3324__, new_new_n3325__,
    new_new_n3326__, new_new_n3327__, new_new_n3328__, new_new_n3329__,
    new_new_n3330__, new_new_n3331__, new_new_n3332__, new_new_n3333__,
    new_new_n3334__, new_new_n3335__, new_new_n3336__, new_new_n3337__,
    new_new_n3338__, new_new_n3339__, new_new_n3340__, new_new_n3341__,
    new_new_n3342__, new_new_n3343__, new_new_n3344__, new_new_n3345__,
    new_new_n3346__, new_new_n3347__, new_new_n3348__, new_new_n3349__,
    new_new_n3350__, new_new_n3351__, new_new_n3352__, new_new_n3353__,
    new_new_n3354__, new_new_n3355__, new_new_n3356__, new_new_n3357__,
    new_new_n3358__, new_new_n3359__, new_new_n3360__, new_new_n3361__,
    new_new_n3362__, new_new_n3363__, new_new_n3364__, new_new_n3365__,
    new_new_n3366__, new_new_n3367__, new_new_n3368__, new_new_n3369__,
    new_new_n3370__, new_new_n3371__, new_new_n3372__, new_new_n3373__,
    new_new_n3374__, new_new_n3375__, new_new_n3376__, new_new_n3377__,
    new_new_n3378__, new_new_n3379__, new_new_n3380__, new_new_n3381__,
    new_new_n3382__, new_new_n3383__, new_new_n3384__, new_new_n3385__,
    new_new_n3386__, new_new_n3387__, new_new_n3388__, new_new_n3389__,
    new_new_n3390__, new_new_n3391__, new_new_n3392__, new_new_n3393__,
    new_new_n3394__, new_new_n3395__, new_new_n3396__, new_new_n3397__,
    new_new_n3398__, new_new_n3399__, new_new_n3400__, new_new_n3401__,
    new_new_n3402__, new_new_n3403__, new_new_n3404__, new_new_n3405__,
    new_new_n3406__, new_new_n3407__, new_new_n3408__, new_new_n3409__,
    new_new_n3410__, new_new_n3411__, new_new_n3412__, new_new_n3413__,
    new_new_n3414__, new_new_n3415__, new_new_n3416__, new_new_n3417__,
    new_new_n3418__, new_new_n3419__, new_new_n3420__, new_new_n3421__,
    new_new_n3422__, new_new_n3423__, new_new_n3424__, new_new_n3425__,
    new_new_n3426__, new_new_n3427__, new_new_n3428__, new_new_n3429__,
    new_new_n3430__, new_new_n3431__, new_new_n3432__, new_new_n3433__,
    new_new_n3434__, new_new_n3435__, new_new_n3436__, new_new_n3437__,
    new_new_n3438__, new_new_n3439__, new_new_n3440__, new_new_n3441__,
    new_new_n3442__, new_new_n3443__, new_new_n3444__, new_new_n3445__,
    new_new_n3446__, new_new_n3447__, new_new_n3448__, new_new_n3449__,
    new_new_n3450__, new_new_n3451__, new_new_n3452__, new_new_n3453__,
    new_new_n3454__, new_new_n3455__, new_new_n3456__, new_new_n3457__,
    new_new_n3458__, new_new_n3459__, new_new_n3460__, new_new_n3461__,
    new_new_n3462__, new_new_n3463__, new_new_n3464__, new_new_n3465__,
    new_new_n3466__, new_new_n3467__, new_new_n3468__, new_new_n3469__,
    new_new_n3470__, new_new_n3471__, new_new_n3472__, new_new_n3473__,
    new_new_n3474__, new_new_n3475__, new_new_n3476__, new_new_n3477__,
    new_new_n3478__, new_new_n3479__, new_new_n3480__, new_new_n3481__,
    new_new_n3482__, new_new_n3483__, new_new_n3484__, new_new_n3485__,
    new_new_n3486__, new_new_n3487__, new_new_n3488__, new_new_n3489__,
    new_new_n3490__, new_new_n3491__, new_new_n3492__, new_new_n3493__,
    new_new_n3494__, new_new_n3495__, new_new_n3496__, new_new_n3497__,
    new_new_n3498__, new_new_n3499__, new_new_n3500__, new_new_n3501__,
    new_new_n3502__, new_new_n3503__, new_new_n3504__, new_new_n3505__,
    new_new_n3506__, new_new_n3507__, new_new_n3508__, new_new_n3509__,
    new_new_n3510__, new_new_n3511__, new_new_n3512__, new_new_n3513__,
    new_new_n3514__, new_new_n3515__, new_new_n3516__, new_new_n3517__,
    new_new_n3518__, new_new_n3519__, new_new_n3520__, new_new_n3521__,
    new_new_n3522__, new_new_n3523__, new_new_n3524__, new_new_n3525__,
    new_new_n3526__, new_new_n3527__, new_new_n3528__, new_new_n3529__,
    new_new_n3530__, new_new_n3531__, new_new_n3532__, new_new_n3533__,
    new_new_n3534__, new_new_n3535__, new_new_n3536__, new_new_n3537__,
    new_new_n3538__, new_new_n3539__, new_new_n3540__, new_new_n3541__,
    new_new_n3542__, new_new_n3543__, new_new_n3544__, new_new_n3545__,
    new_new_n3546__, new_new_n3547__, new_new_n3548__, new_new_n3549__,
    new_new_n3550__, new_new_n3551__, new_new_n3552__, new_new_n3553__,
    new_new_n3554__, new_new_n3555__, new_new_n3556__, new_new_n3557__,
    new_new_n3558__, new_new_n3559__, new_new_n3560__, new_new_n3561__,
    new_new_n3562__, new_new_n3563__, new_new_n3564__, new_new_n3565__,
    new_new_n3566__, new_new_n3567__, new_new_n3568__, new_new_n3569__,
    new_new_n3570__, new_new_n3571__, new_new_n3572__, new_new_n3573__,
    new_new_n3574__, new_new_n3575__, new_new_n3576__, new_new_n3577__,
    new_new_n3578__, new_new_n3579__, new_new_n3580__, new_new_n3581__,
    new_new_n3582__, new_new_n3583__, new_new_n3584__, new_new_n3585__,
    new_new_n3586__, new_new_n3587__, new_new_n3588__, new_new_n3589__,
    new_new_n3590__, new_new_n3591__, new_new_n3592__, new_new_n3593__,
    new_new_n3594__, new_new_n3595__, new_new_n3596__, new_new_n3597__,
    new_new_n3598__, new_new_n3599__, new_new_n3600__, new_new_n3601__,
    new_new_n3602__, new_new_n3603__, new_new_n3604__, new_new_n3605__,
    new_new_n3606__, new_new_n3607__, new_new_n3608__, new_new_n3609__,
    new_new_n3610__, new_new_n3611__, new_new_n3612__, new_new_n3613__,
    new_new_n3614__, new_new_n3615__, new_new_n3616__, new_new_n3617__,
    new_new_n3618__, new_new_n3619__, new_new_n3620__, new_new_n3621__,
    new_new_n3622__, new_new_n3623__, new_new_n3624__, new_new_n3625__,
    new_new_n3626__, new_new_n3627__, new_new_n3628__, new_new_n3629__,
    new_new_n3630__, new_new_n3631__, new_new_n3632__, new_new_n3633__,
    new_new_n3634__, new_new_n3635__, new_new_n3636__, new_new_n3637__,
    new_new_n3638__, new_new_n3639__, new_new_n3640__, new_new_n3641__,
    new_new_n3642__, new_new_n3643__, new_new_n3644__, new_new_n3645__,
    new_new_n3646__, new_new_n3647__, new_new_n3648__, new_new_n3649__,
    new_new_n3650__, new_new_n3651__, new_new_n3652__, new_new_n3653__,
    new_new_n3654__, new_new_n3655__, new_new_n3656__, new_new_n3657__,
    new_new_n3658__, new_new_n3659__, new_new_n3660__, new_new_n3661__,
    new_new_n3662__, new_new_n3663__, new_new_n3664__, new_new_n3665__,
    new_new_n3666__, new_new_n3667__, new_new_n3668__, new_new_n3669__,
    new_new_n3670__, new_new_n3671__, new_new_n3672__, new_new_n3673__,
    new_new_n3674__, new_new_n3675__, new_new_n3676__, new_new_n3677__,
    new_new_n3678__, new_new_n3679__, new_new_n3680__, new_new_n3681__,
    new_new_n3682__, new_new_n3683__, new_new_n3684__, new_new_n3685__,
    new_new_n3686__, new_new_n3687__, new_new_n3688__, new_new_n3689__,
    new_new_n3690__, new_new_n3691__, new_new_n3692__, new_new_n3693__,
    new_new_n3694__, new_new_n3695__, new_new_n3696__, new_new_n3697__,
    new_new_n3698__, new_new_n3699__, new_new_n3700__, new_new_n3701__,
    new_new_n3702__, new_new_n3703__, new_new_n3704__, new_new_n3705__,
    new_new_n3706__, new_new_n3707__, new_new_n3708__, new_new_n3709__,
    new_new_n3710__, new_new_n3711__, new_new_n3712__, new_new_n3713__,
    new_new_n3714__, new_new_n3715__, new_new_n3716__, new_new_n3717__,
    new_new_n3718__, new_new_n3719__, new_new_n3720__, new_new_n3721__,
    new_new_n3722__, new_new_n3723__, new_new_n3724__, new_new_n3725__,
    new_new_n3726__, new_new_n3727__, new_new_n3728__, new_new_n3729__,
    new_new_n3730__, new_new_n3731__, new_new_n3732__, new_new_n3733__,
    new_new_n3734__, new_new_n3735__, new_new_n3736__, new_new_n3737__,
    new_new_n3738__, new_new_n3739__, new_new_n3740__, new_new_n3741__,
    new_new_n3742__, new_new_n3743__, new_new_n3744__, new_new_n3745__,
    new_new_n3746__, new_new_n3747__, new_new_n3748__, new_new_n3749__,
    new_new_n3750__, new_new_n3751__, new_new_n3752__, new_new_n3753__,
    new_new_n3754__, new_new_n3755__, new_new_n3756__, new_new_n3757__,
    new_new_n3758__, new_new_n3759__, new_new_n3760__, new_new_n3761__,
    new_new_n3762__, new_new_n3763__, new_new_n3764__, new_new_n3765__,
    new_new_n3766__, new_new_n3767__, new_new_n3768__, new_new_n3769__,
    new_new_n3770__, new_new_n3771__, new_new_n3772__, new_new_n3773__,
    new_new_n3774__, new_new_n3775__, new_new_n3776__, new_new_n3777__,
    new_new_n3778__, new_new_n3779__, new_new_n3780__, new_new_n3781__,
    new_new_n3782__, new_new_n3783__, new_new_n3784__, new_new_n3785__,
    new_new_n3786__, new_new_n3787__, new_new_n3788__, new_new_n3789__,
    new_new_n3790__, new_new_n3791__, new_new_n3792__, new_new_n3793__,
    new_new_n3794__, new_new_n3795__, new_new_n3796__, new_new_n3797__,
    new_new_n3798__, new_new_n3799__, new_new_n3800__, new_new_n3801__,
    new_new_n3802__, new_new_n3803__, new_new_n3804__, new_new_n3805__,
    new_new_n3806__, new_new_n3807__, new_new_n3808__, new_new_n3809__,
    new_new_n3810__, new_new_n3811__, new_new_n3812__, new_new_n3813__,
    new_new_n3814__, new_new_n3815__, new_new_n3816__, new_new_n3817__,
    new_new_n3818__, new_new_n3819__, new_new_n3820__, new_new_n3821__,
    new_new_n3822__, new_new_n3823__, new_new_n3824__, new_new_n3825__,
    new_new_n3826__, new_new_n3827__, new_new_n3828__, new_new_n3829__,
    new_new_n3830__, new_new_n3831__, new_new_n3832__, new_new_n3833__,
    new_new_n3834__, new_new_n3835__, new_new_n3836__, new_new_n3837__,
    new_new_n3838__, new_new_n3839__, new_new_n3840__, new_new_n3841__,
    new_new_n3842__, new_new_n3843__, new_new_n3844__, new_new_n3845__,
    new_new_n3846__, new_new_n3847__, new_new_n3848__, new_new_n3849__,
    new_new_n3850__, new_new_n3851__, new_new_n3852__, new_new_n3853__,
    new_new_n3854__, new_new_n3855__, new_new_n3856__, new_new_n3857__,
    new_new_n3858__, new_new_n3859__, new_new_n3860__, new_new_n3861__,
    new_new_n3862__, new_new_n3863__, new_new_n3864__, new_new_n3865__,
    new_new_n3866__, new_new_n3867__, new_new_n3868__, new_new_n3869__,
    new_new_n3870__, n6268, n6271, n6274, n6277, n6280, n6283, n6286,
    n6289, n6292, n6295, n6298, n6301, n6304, n6307, n6310, n6313, n6316,
    n6319, n6322, n6325, n6328, n6331, n6334, n6337, n6340, n6343, n6346,
    n6349, n6352, n6355, n6358, n6361, n6364, n6367, n6370, n6373, n6376,
    n6379, n6382, n6385, n6388, n6391, n6394, n6397, n6400, n6403, n6406,
    n6409, n6412, n6415, n6418, n6421, n6424, n6427, n6430, n6433, n6436,
    n6439, n6442, n6445, n6448, n6451, n6454, n6457, n6460, n6463, n6466,
    n6469, n6472, n6475, n6478, n6481, n6484, n6487, n6490, n6493, n6496,
    n6499, n6502, n6505, n6508, n6511, n6514, n6517, n6520, n6523, n6526,
    n6529, n6532, n6535, n6538, n6541, n6544, n6547, n6550, n6553, n6556,
    n6559, n6562, n6565, n6568, n6571, n6574, n6577, n6580, n6583, n6586,
    n6589, n6592, n6595, n6598, n6601, n6604, n6607, n6610, n6613, n6616,
    n6619, n6622, n6625, n6628, n6631, n6634, n6637, n6640, n6643, n6646,
    n6649, n6652, n6655, n6658, n6661, n6664, n6667, n6670, n6673, n6676,
    n6679, n6682, n6685, n6688, n6691, n6694, n6697, n6700, n6703, n6706,
    n6709, n6712, n6715, n6718, n6721, n6724, n6727, n6730, n6733, n6736,
    n6739, n6742, n6745, n6748, n6751, n6754, n6757, n6760, n6763, n6766,
    n6769, n6772, n6775, n6778, n6781, n6784, n6787, n6790, n6793, n6796,
    n6799, n6802, n6805, n6808, n6811, n6814, n6817, n6820, n6823, n6826,
    n6829, n6832, n6835, n6838, n6841, n6844, n6847, n6850, n6853, n6856,
    n6859, n6862, n6865, n6868, n6871, n6874, n6877, n6880, n6883, n6886,
    n6889, n6892, n6895, n6898, n6901, n6904, n6907, n6910, n6913, n6916,
    n6919, n6922, n6925, n6928, n6931, n6934, n6937, n6940, n6943, n6946,
    n6949, n6952, n6955, n6958, n6961, n6964, n6967, n6970, n6973, n6976,
    n6979, n6982, n6985, n6988, n6991, n6994, n6997, n7000, n7003, n7006,
    n7009, n7012, n7015, n7018, n7021, n7024, n7027, n7030, n7033, n7036,
    n7039, n7042, n7045, n7048, n7051, n7054, n7057, n7060, n7063, n7066,
    n7069, n7072, n7075, n7078, n7081, n7084, n7087, n7090, n7093, n7096,
    n7099, n7102, n7105, n7108, n7111, n7114, n7117, n7120, n7123, n7126,
    n7129, n7132, n7135, n7138, n7141, n7144, n7147, n7150, n7153, n7156,
    n7159, n7162, n7165, n7168, n7171, n7174, n7177, n7180, n7183, n7186,
    n7189, n7192, n7195, n7198, n7201, n7204, n7207, n7210, n7213, n7216,
    n7219, n7222, n7225, n7228, n7231, n7234, n7237, n7240, n7243, n7246,
    n7249, n7252, n7255, n7258, n7261, n7264, n7267, n7270, n7273, n7276,
    n7279, n7282, n7285, n7288, n7291, n7294, n7297, n7300, n7303, n7306,
    n7309, n7312, n7315, n7318, n7321, n7324, n7327, n7330, n7333, n7336,
    n7339, n7342, n7345, n7348;
  buf1  g0000(.din(G1), .dout(new_new_n795__));
  not1  g0001(.din(G1), .dout(new_new_n796__));
  buf1  g0002(.din(G2), .dout(new_new_n797__));
  not1  g0003(.din(G2), .dout(new_new_n798__));
  buf1  g0004(.din(G3), .dout(new_new_n799__));
  not1  g0005(.din(G3), .dout(new_new_n800__));
  buf1  g0006(.din(G4), .dout(new_new_n801__));
  not1  g0007(.din(G4), .dout(new_new_n802__));
  buf1  g0008(.din(G5), .dout(new_new_n803__));
  buf1  g0009(.din(G6), .dout(new_new_n805__));
  buf1  g0010(.din(G7), .dout(new_new_n807__));
  buf1  g0011(.din(G8), .dout(new_new_n809__));
  buf1  g0012(.din(G9), .dout(new_new_n811__));
  buf1  g0013(.din(G10), .dout(new_new_n813__));
  buf1  g0014(.din(G11), .dout(new_new_n815__));
  buf1  g0015(.din(G12), .dout(new_new_n817__));
  not1  g0016(.din(G12), .dout(new_new_n818__));
  buf1  g0017(.din(G13), .dout(new_new_n819__));
  not1  g0018(.din(G13), .dout(new_new_n820__));
  buf1  g0019(.din(G14), .dout(new_new_n821__));
  buf1  g0020(.din(G15), .dout(new_new_n823__));
  buf1  g0021(.din(G16), .dout(new_new_n825__));
  buf1  g0022(.din(G17), .dout(new_new_n827__));
  buf1  g0023(.din(G18), .dout(new_new_n829__));
  buf1  g0024(.din(G19), .dout(new_new_n831__));
  buf1  g0025(.din(G20), .dout(new_new_n833__));
  buf1  g0026(.din(G21), .dout(new_new_n835__));
  buf1  g0027(.din(G22), .dout(new_new_n837__));
  buf1  g0028(.din(G23), .dout(new_new_n839__));
  buf1  g0029(.din(G24), .dout(new_new_n841__));
  buf1  g0030(.din(G25), .dout(new_new_n843__));
  buf1  g0031(.din(G26), .dout(new_new_n845__));
  buf1  g0032(.din(G27), .dout(new_new_n847__));
  buf1  g0033(.din(G28), .dout(new_new_n849__));
  buf1  g0034(.din(G29), .dout(new_new_n851__));
  buf1  g0035(.din(G30), .dout(new_new_n853__));
  buf1  g0036(.din(G31), .dout(new_new_n855__));
  buf1  g0037(.din(G32), .dout(new_new_n857__));
  not1  g0038(.din(G32), .dout(new_new_n858__));
  buf1  g0039(.din(G33), .dout(new_new_n859__));
  not1  g0040(.din(G33), .dout(new_new_n860__));
  buf1  g0041(.din(G34), .dout(new_new_n861__));
  not1  g0042(.din(G34), .dout(new_new_n862__));
  buf1  g0043(.din(G35), .dout(new_new_n863__));
  buf1  g0044(.din(G36), .dout(new_new_n865__));
  not1  g0045(.din(G36), .dout(new_new_n866__));
  buf1  g0046(.din(G37), .dout(new_new_n867__));
  buf1  g0047(.din(G38), .dout(new_new_n869__));
  buf1  g0048(.din(G39), .dout(new_new_n871__));
  not1  g0049(.din(G39), .dout(new_new_n872__));
  buf1  g0050(.din(G40), .dout(new_new_n873__));
  buf1  g0051(.din(G41), .dout(new_new_n875__));
  buf1  g0052(.din(G42), .dout(new_new_n877__));
  buf1  g0053(.din(G43), .dout(new_new_n879__));
  buf1  g0054(.din(G44), .dout(new_new_n881__));
  buf1  g0055(.din(G45), .dout(new_new_n883__));
  buf1  g0056(.din(G46), .dout(new_new_n885__));
  buf1  g0057(.din(G47), .dout(new_new_n887__));
  buf1  g0058(.din(G48), .dout(new_new_n889__));
  buf1  g0059(.din(G49), .dout(new_new_n891__));
  buf1  g0060(.din(G50), .dout(new_new_n893__));
  not1  g0061(.din(n1752_lo), .dout(new_new_n896__));
  buf1  g0062(.din(n1776_lo), .dout(new_new_n897__));
  not1  g0063(.din(n1776_lo), .dout(new_new_n898__));
  buf1  g0064(.din(n1824_lo), .dout(new_new_n899__));
  not1  g0065(.din(n1824_lo), .dout(new_new_n900__));
  buf1  g0066(.din(n1836_lo), .dout(new_new_n901__));
  buf1  g0067(.din(n1848_lo), .dout(new_new_n903__));
  not1  g0068(.din(n1848_lo), .dout(new_new_n904__));
  buf1  g0069(.din(n1860_lo), .dout(new_new_n905__));
  not1  g0070(.din(n1860_lo), .dout(new_new_n906__));
  buf1  g0071(.din(n1872_lo), .dout(new_new_n907__));
  not1  g0072(.din(n1872_lo), .dout(new_new_n908__));
  buf1  g0073(.din(n1884_lo), .dout(new_new_n909__));
  not1  g0074(.din(n1884_lo), .dout(new_new_n910__));
  buf1  g0075(.din(n1896_lo), .dout(new_new_n911__));
  not1  g0076(.din(n1896_lo), .dout(new_new_n912__));
  buf1  g0077(.din(n1908_lo), .dout(new_new_n913__));
  not1  g0078(.din(n1908_lo), .dout(new_new_n914__));
  buf1  g0079(.din(n1911_lo), .dout(new_new_n915__));
  buf1  g0080(.din(n1914_lo), .dout(new_new_n917__));
  buf1  g0081(.din(n1923_lo), .dout(new_new_n919__));
  buf1  g0082(.din(n1926_lo), .dout(new_new_n921__));
  buf1  g0083(.din(n1935_lo), .dout(new_new_n923__));
  buf1  g0084(.din(n1938_lo), .dout(new_new_n925__));
  buf1  g0085(.din(n1947_lo), .dout(new_new_n927__));
  buf1  g0086(.din(n1950_lo), .dout(new_new_n929__));
  buf1  g0087(.din(n1959_lo), .dout(new_new_n931__));
  buf1  g0088(.din(n1962_lo), .dout(new_new_n933__));
  buf1  g0089(.din(n1971_lo), .dout(new_new_n935__));
  buf1  g0090(.din(n1974_lo), .dout(new_new_n937__));
  not1  g0091(.din(n1974_lo), .dout(new_new_n938__));
  buf1  g0092(.din(n1983_lo), .dout(new_new_n939__));
  buf1  g0093(.din(n1995_lo), .dout(new_new_n941__));
  buf1  g0094(.din(n2055_lo), .dout(new_new_n943__));
  not1  g0095(.din(n2055_lo), .dout(new_new_n944__));
  buf1  g0096(.din(n2064_lo), .dout(new_new_n945__));
  not1  g0097(.din(n2064_lo), .dout(new_new_n946__));
  buf1  g0098(.din(n2067_lo), .dout(new_new_n947__));
  buf1  g0099(.din(n2079_lo), .dout(new_new_n949__));
  buf1  g0100(.din(n2100_lo), .dout(new_new_n951__));
  not1  g0101(.din(n2100_lo), .dout(new_new_n952__));
  buf1  g0102(.din(n2112_lo), .dout(new_new_n953__));
  not1  g0103(.din(n2112_lo), .dout(new_new_n954__));
  buf1  g0104(.din(n2124_lo), .dout(new_new_n955__));
  not1  g0105(.din(n2124_lo), .dout(new_new_n956__));
  buf1  g0106(.din(n2136_lo), .dout(new_new_n957__));
  not1  g0107(.din(n2136_lo), .dout(new_new_n958__));
  buf1  g0108(.din(n2148_lo), .dout(new_new_n959__));
  not1  g0109(.din(n2148_lo), .dout(new_new_n960__));
  buf1  g0110(.din(n2160_lo), .dout(new_new_n961__));
  not1  g0111(.din(n2160_lo), .dout(new_new_n962__));
  buf1  g0112(.din(n2172_lo), .dout(new_new_n963__));
  not1  g0113(.din(n2172_lo), .dout(new_new_n964__));
  buf1  g0114(.din(n2184_lo), .dout(new_new_n965__));
  not1  g0115(.din(n2184_lo), .dout(new_new_n966__));
  buf1  g0116(.din(n2235_lo), .dout(new_new_n967__));
  buf1  g0117(.din(n2238_lo), .dout(new_new_n969__));
  not1  g0118(.din(n2238_lo), .dout(new_new_n970__));
  buf1  g0119(.din(n2247_lo), .dout(new_new_n971__));
  buf1  g0120(.din(n2250_lo), .dout(new_new_n973__));
  buf1  g0121(.din(n2259_lo), .dout(new_new_n975__));
  buf1  g0122(.din(n2262_lo), .dout(new_new_n977__));
  buf1  g0123(.din(n2271_lo), .dout(new_new_n979__));
  buf1  g0124(.din(n2274_lo), .dout(new_new_n981__));
  buf1  g0125(.din(n2283_lo), .dout(new_new_n983__));
  buf1  g0126(.din(n2286_lo), .dout(new_new_n985__));
  not1  g0127(.din(n2289_lo), .dout(new_new_n988__));
  buf1  g0128(.din(n2295_lo), .dout(new_new_n989__));
  buf1  g0129(.din(n2298_lo), .dout(new_new_n991__));
  not1  g0130(.din(n2298_lo), .dout(new_new_n992__));
  buf1  g0131(.din(n2304_lo), .dout(new_new_n993__));
  not1  g0132(.din(n2304_lo), .dout(new_new_n994__));
  buf1  g0133(.din(n2307_lo), .dout(new_new_n995__));
  not1  g0134(.din(n2307_lo), .dout(new_new_n996__));
  buf1  g0135(.din(n2316_lo), .dout(new_new_n997__));
  not1  g0136(.din(n2316_lo), .dout(new_new_n998__));
  buf1  g0137(.din(n2331_lo), .dout(new_new_n999__));
  buf1  g0138(.din(n2334_lo), .dout(new_new_n1001__));
  buf1  g0139(.din(n2337_lo), .dout(new_new_n1003__));
  buf1  g0140(.din(n2340_lo), .dout(new_new_n1005__));
  not1  g0141(.din(n2340_lo), .dout(new_new_n1006__));
  buf1  g0142(.din(n2071_o2), .dout(new_new_n1007__));
  not1  g0143(.din(n2071_o2), .dout(new_new_n1008__));
  buf1  g0144(.din(n2080_o2), .dout(new_new_n1009__));
  not1  g0145(.din(n2080_o2), .dout(new_new_n1010__));
  not1  g0146(.din(n2137_o2), .dout(new_new_n1012__));
  not1  g0147(.din(n2368_o2), .dout(new_new_n1014__));
  not1  g0148(.din(n2383_o2), .dout(new_new_n1016__));
  buf1  g0149(.din(n2405_o2), .dout(new_new_n1017__));
  not1  g0150(.din(n2405_o2), .dout(new_new_n1018__));
  buf1  g0151(.din(n2471_o2), .dout(new_new_n1019__));
  buf1  g0152(.din(n2617_o2), .dout(new_new_n1021__));
  buf1  g0153(.din(n2765_o2), .dout(new_new_n1023__));
  buf1  g0154(.din(n2775_o2), .dout(new_new_n1025__));
  not1  g0155(.din(n2775_o2), .dout(new_new_n1026__));
  buf1  g0156(.din(n2829_o2), .dout(new_new_n1027__));
  buf1  g0157(.din(n2579_o2), .dout(new_new_n1029__));
  not1  g0158(.din(n2579_o2), .dout(new_new_n1030__));
  buf1  g0159(.din(n2580_o2), .dout(new_new_n1031__));
  not1  g0160(.din(n2580_o2), .dout(new_new_n1032__));
  buf1  g0161(.din(n2618_o2), .dout(new_new_n1033__));
  buf1  g0162(.din(n2619_o2), .dout(new_new_n1035__));
  not1  g0163(.din(n2619_o2), .dout(new_new_n1036__));
  buf1  g0164(.din(n2620_o2), .dout(new_new_n1037__));
  not1  g0165(.din(n2620_o2), .dout(new_new_n1038__));
  buf1  g0166(.din(n2621_o2), .dout(new_new_n1039__));
  not1  g0167(.din(n2621_o2), .dout(new_new_n1040__));
  buf1  g0168(.din(n2622_o2), .dout(new_new_n1041__));
  not1  g0169(.din(n2622_o2), .dout(new_new_n1042__));
  buf1  g0170(.din(n2623_o2), .dout(new_new_n1043__));
  not1  g0171(.din(n2623_o2), .dout(new_new_n1044__));
  buf1  g0172(.din(n2624_o2), .dout(new_new_n1045__));
  not1  g0173(.din(n2624_o2), .dout(new_new_n1046__));
  buf1  g0174(.din(n2625_o2), .dout(new_new_n1047__));
  buf1  g0175(.din(n2626_o2), .dout(new_new_n1049__));
  buf1  g0176(.din(n2627_o2), .dout(new_new_n1051__));
  not1  g0177(.din(n2627_o2), .dout(new_new_n1052__));
  buf1  g0178(.din(n3029_o2), .dout(new_new_n1053__));
  buf1  g0179(.din(n3035_o2), .dout(new_new_n1055__));
  not1  g0180(.din(n3035_o2), .dout(new_new_n1056__));
  buf1  g0181(.din(n2643_o2), .dout(new_new_n1057__));
  not1  g0182(.din(n2643_o2), .dout(new_new_n1058__));
  buf1  g0183(.din(n2644_o2), .dout(new_new_n1059__));
  buf1  g0184(.din(n2645_o2), .dout(new_new_n1061__));
  not1  g0185(.din(n2645_o2), .dout(new_new_n1062__));
  buf1  g0186(.din(n327_inv), .dout(new_new_n1063__));
  not1  g0187(.din(n327_inv), .dout(new_new_n1064__));
  buf1  g0188(.din(n2658_o2), .dout(new_new_n1065__));
  not1  g0189(.din(n2659_o2), .dout(new_new_n1068__));
  buf1  g0190(.din(n2674_o2), .dout(new_new_n1069__));
  buf1  g0191(.din(n2675_o2), .dout(new_new_n1071__));
  buf1  g0192(.din(n2676_o2), .dout(new_new_n1073__));
  not1  g0193(.din(n2676_o2), .dout(new_new_n1074__));
  buf1  g0194(.din(n3119_o2), .dout(new_new_n1075__));
  not1  g0195(.din(n3119_o2), .dout(new_new_n1076__));
  buf1  g0196(.din(n3153_o2), .dout(new_new_n1077__));
  buf1  g0197(.din(n351_inv), .dout(new_new_n1079__));
  buf1  g0198(.din(n2729_o2), .dout(new_new_n1081__));
  not1  g0199(.din(n2729_o2), .dout(new_new_n1082__));
  buf1  g0200(.din(n2730_o2), .dout(new_new_n1083__));
  not1  g0201(.din(n2730_o2), .dout(new_new_n1084__));
  buf1  g0202(.din(n2731_o2), .dout(new_new_n1085__));
  buf1  g0203(.din(n698_o2), .dout(new_new_n1087__));
  not1  g0204(.din(n698_o2), .dout(new_new_n1088__));
  not1  g0205(.din(n366_inv), .dout(new_new_n1090__));
  buf1  g0206(.din(n2757_o2), .dout(new_new_n1091__));
  buf1  g0207(.din(n2758_o2), .dout(new_new_n1093__));
  buf1  g0208(.din(n1000_o2), .dout(new_new_n1095__));
  buf1  g0209(.din(n1160_o2), .dout(new_new_n1097__));
  not1  g0210(.din(n1160_o2), .dout(new_new_n1098__));
  buf1  g0211(.din(n1153_o2), .dout(new_new_n1099__));
  not1  g0212(.din(n1153_o2), .dout(new_new_n1100__));
  buf1  g0213(.din(n2793_o2), .dout(new_new_n1101__));
  not1  g0214(.din(n2793_o2), .dout(new_new_n1102__));
  buf1  g0215(.din(n2794_o2), .dout(new_new_n1103__));
  not1  g0216(.din(n2794_o2), .dout(new_new_n1104__));
  buf1  g0217(.din(n2795_o2), .dout(new_new_n1105__));
  not1  g0218(.din(n2795_o2), .dout(new_new_n1106__));
  buf1  g0219(.din(n1001_o2), .dout(new_new_n1107__));
  not1  g0220(.din(n1001_o2), .dout(new_new_n1108__));
  not1  g0221(.din(n2859_o2), .dout(new_new_n1110__));
  buf1  g0222(.din(n744_o2), .dout(new_new_n1111__));
  not1  g0223(.din(n744_o2), .dout(new_new_n1112__));
  buf1  g0224(.din(n402_inv), .dout(new_new_n1113__));
  buf1  g0225(.din(n2926_o2), .dout(new_new_n1115__));
  not1  g0226(.din(n2926_o2), .dout(new_new_n1116__));
  buf1  g0227(.din(n408_inv), .dout(new_new_n1117__));
  buf1  g0228(.din(n2966_o2), .dout(new_new_n1119__));
  buf1  g0229(.din(n2967_o2), .dout(new_new_n1121__));
  buf1  g0230(.din(n2947_o2), .dout(new_new_n1123__));
  buf1  g0231(.din(n1010_o2), .dout(new_new_n1125__));
  not1  g0232(.din(n1010_o2), .dout(new_new_n1126__));
  buf1  g0233(.din(n2976_o2), .dout(new_new_n1127__));
  not1  g0234(.din(n2976_o2), .dout(new_new_n1128__));
  buf1  g0235(.din(n3069_o2), .dout(new_new_n1129__));
  buf1  g0236(.din(n3028_o2), .dout(new_new_n1131__));
  not1  g0237(.din(n3028_o2), .dout(new_new_n1132__));
  buf1  g0238(.din(n3081_o2), .dout(new_new_n1133__));
  not1  g0239(.din(n3081_o2), .dout(new_new_n1134__));
  buf1  g0240(.din(n3082_o2), .dout(new_new_n1135__));
  not1  g0241(.din(n3082_o2), .dout(new_new_n1136__));
  buf1  g0242(.din(n3142_o2), .dout(new_new_n1137__));
  buf1  g0243(.din(n3214_o2), .dout(new_new_n1139__));
  not1  g0244(.din(n3214_o2), .dout(new_new_n1140__));
  buf1  g0245(.din(n2992_o2), .dout(new_new_n1141__));
  buf1  g0246(.din(n2993_o2), .dout(new_new_n1143__));
  not1  g0247(.din(n2993_o2), .dout(new_new_n1144__));
  buf1  g0248(.din(n870_o2), .dout(new_new_n1145__));
  buf1  g0249(.din(n3086_o2), .dout(new_new_n1147__));
  buf1  g0250(.din(n3087_o2), .dout(new_new_n1149__));
  not1  g0251(.din(n3087_o2), .dout(new_new_n1150__));
  buf1  g0252(.din(n3088_o2), .dout(new_new_n1151__));
  buf1  g0253(.din(n3089_o2), .dout(new_new_n1153__));
  not1  g0254(.din(n3089_o2), .dout(new_new_n1154__));
  buf1  g0255(.din(n3090_o2), .dout(new_new_n1155__));
  not1  g0256(.din(n3090_o2), .dout(new_new_n1156__));
  buf1  g0257(.din(n3091_o2), .dout(new_new_n1157__));
  not1  g0258(.din(n3091_o2), .dout(new_new_n1158__));
  buf1  g0259(.din(n3092_o2), .dout(new_new_n1159__));
  not1  g0260(.din(n3092_o2), .dout(new_new_n1160__));
  buf1  g0261(.din(n3093_o2), .dout(new_new_n1161__));
  buf1  g0262(.din(n3094_o2), .dout(new_new_n1163__));
  buf1  g0263(.din(n3095_o2), .dout(new_new_n1165__));
  buf1  g0264(.din(n483_inv), .dout(new_new_n1167__));
  buf1  g0265(.din(n3170_o2), .dout(new_new_n1169__));
  buf1  g0266(.din(n3171_o2), .dout(new_new_n1171__));
  buf1  g0267(.din(n3172_o2), .dout(new_new_n1173__));
  not1  g0268(.din(n3172_o2), .dout(new_new_n1174__));
  buf1  g0269(.din(n3179_o2), .dout(new_new_n1175__));
  buf1  g0270(.din(n498_inv), .dout(new_new_n1177__));
  not1  g0271(.din(n3193_o2), .dout(new_new_n1180__));
  buf1  g0272(.din(n3211_o2), .dout(new_new_n1181__));
  buf1  g0273(.din(n3212_o2), .dout(new_new_n1183__));
  buf1  g0274(.din(n3213_o2), .dout(new_new_n1185__));
  buf1  g0275(.din(n513_inv), .dout(new_new_n1187__));
  buf1  g0276(.din(n1125_o2), .dout(new_new_n1189__));
  not1  g0277(.din(n1125_o2), .dout(new_new_n1190__));
  buf1  g0278(.din(n1081_o2), .dout(new_new_n1191__));
  not1  g0279(.din(n1081_o2), .dout(new_new_n1192__));
  not1  g0280(.din(n1139_o2), .dout(new_new_n1194__));
  buf1  g0281(.din(n3245_o2), .dout(new_new_n1195__));
  not1  g0282(.din(n3245_o2), .dout(new_new_n1196__));
  buf1  g0283(.din(n3246_o2), .dout(new_new_n1197__));
  not1  g0284(.din(n3246_o2), .dout(new_new_n1198__));
  buf1  g0285(.din(n3247_o2), .dout(new_new_n1199__));
  buf1  g0286(.din(lo074_buf_o2), .dout(new_new_n1201__));
  not1  g0287(.din(lo074_buf_o2), .dout(new_new_n1202__));
  buf1  g0288(.din(lo078_buf_o2), .dout(new_new_n1203__));
  not1  g0289(.din(lo078_buf_o2), .dout(new_new_n1204__));
  buf1  g0290(.din(lo186_buf_o2), .dout(new_new_n1205__));
  not1  g0291(.din(lo186_buf_o2), .dout(new_new_n1206__));
  buf1  g0292(.din(lo118_buf_o2), .dout(new_new_n1207__));
  buf1  g0293(.din(lo146_buf_o2), .dout(new_new_n1209__));
  buf1  g0294(.din(n1038_o2), .dout(new_new_n1211__));
  not1  g0295(.din(n1038_o2), .dout(new_new_n1212__));
  buf1  g0296(.din(n1044_o2), .dout(new_new_n1213__));
  not1  g0297(.din(n1044_o2), .dout(new_new_n1214__));
  buf1  g0298(.din(n555_inv), .dout(new_new_n1215__));
  buf1  g0299(.din(n558_inv), .dout(new_new_n1217__));
  buf1  g0300(.din(lo026_buf_o2), .dout(new_new_n1219__));
  not1  g0301(.din(lo026_buf_o2), .dout(new_new_n1220__));
  buf1  g0302(.din(lo030_buf_o2), .dout(new_new_n1221__));
  not1  g0303(.din(lo030_buf_o2), .dout(new_new_n1222__));
  buf1  g0304(.din(lo090_buf_o2), .dout(new_new_n1223__));
  buf1  g0305(.din(lo094_buf_o2), .dout(new_new_n1225__));
  not1  g0306(.din(lo094_buf_o2), .dout(new_new_n1226__));
  buf1  g0307(.din(lo098_buf_o2), .dout(new_new_n1227__));
  not1  g0308(.din(lo098_buf_o2), .dout(new_new_n1228__));
  buf1  g0309(.din(lo102_buf_o2), .dout(new_new_n1229__));
  not1  g0310(.din(lo102_buf_o2), .dout(new_new_n1230__));
  buf1  g0311(.din(lo066_buf_o2), .dout(new_new_n1231__));
  buf1  g0312(.din(lo070_buf_o2), .dout(new_new_n1233__));
  not1  g0313(.din(n1202_o2), .dout(new_new_n1236__));
  buf1  g0314(.din(n1003_o2), .dout(new_new_n1237__));
  not1  g0315(.din(n1003_o2), .dout(new_new_n1238__));
  buf1  g0316(.din(n1031_o2), .dout(new_new_n1239__));
  not1  g0317(.din(n1031_o2), .dout(new_new_n1240__));
  buf1  g0318(.din(n1034_o2), .dout(new_new_n1241__));
  not1  g0319(.din(n1034_o2), .dout(new_new_n1242__));
  buf1  g0320(.din(n1040_o2), .dout(new_new_n1243__));
  not1  g0321(.din(n1040_o2), .dout(new_new_n1244__));
  buf1  g0322(.din(n1046_o2), .dout(new_new_n1245__));
  not1  g0323(.din(n1046_o2), .dout(new_new_n1246__));
  buf1  g0324(.din(n1380_o2), .dout(new_new_n1247__));
  buf1  g0325(.din(n1425_o2), .dout(new_new_n1249__));
  buf1  g0326(.din(n697_o2), .dout(new_new_n1251__));
  not1  g0327(.din(n1143_o2), .dout(new_new_n1254__));
  buf1  g0328(.din(n673_o2), .dout(new_new_n1255__));
  buf1  g0329(.din(n789_o2), .dout(new_new_n1257__));
  not1  g0330(.din(n789_o2), .dout(new_new_n1258__));
  buf1  g0331(.din(n786_o2), .dout(new_new_n1259__));
  not1  g0332(.din(n786_o2), .dout(new_new_n1260__));
  buf1  g0333(.din(n1047_o2), .dout(new_new_n1261__));
  buf1  g0334(.din(n1036_o2), .dout(new_new_n1263__));
  buf1  g0335(.din(n1307_o2), .dout(new_new_n1265__));
  buf1  g0336(.din(n1035_o2), .dout(new_new_n1267__));
  buf1  g0337(.din(n1297_o2), .dout(new_new_n1269__));
  not1  g0338(.din(n1099_o2), .dout(new_new_n1272__));
  buf1  g0339(.din(n1128_o2), .dout(new_new_n1273__));
  not1  g0340(.din(n1128_o2), .dout(new_new_n1274__));
  buf1  g0341(.din(n645_inv), .dout(new_new_n1275__));
  buf1  g0342(.din(n826_o2), .dout(new_new_n1277__));
  buf1  g0343(.din(n853_o2), .dout(new_new_n1279__));
  buf1  g0344(.din(n654_inv), .dout(new_new_n1281__));
  buf1  g0345(.din(n700_o2), .dout(new_new_n1283__));
  buf1  g0346(.din(n884_o2), .dout(new_new_n1285__));
  not1  g0347(.din(n884_o2), .dout(new_new_n1286__));
  buf1  g0348(.din(lo082_buf_o2), .dout(new_new_n1287__));
  not1  g0349(.din(lo082_buf_o2), .dout(new_new_n1288__));
  buf1  g0350(.din(lo086_buf_o2), .dout(new_new_n1289__));
  not1  g0351(.din(lo086_buf_o2), .dout(new_new_n1290__));
  buf1  g0352(.din(n801_o2), .dout(new_new_n1291__));
  not1  g0353(.din(n801_o2), .dout(new_new_n1292__));
  buf1  g0354(.din(n840_o2), .dout(new_new_n1293__));
  not1  g0355(.din(n840_o2), .dout(new_new_n1294__));
  buf1  g0356(.din(n675_inv), .dout(new_new_n1295__));
  not1  g0357(.din(n675_inv), .dout(new_new_n1296__));
  buf1  g0358(.din(lo002_buf_o2), .dout(new_new_n1297__));
  not1  g0359(.din(lo002_buf_o2), .dout(new_new_n1298__));
  buf1  g0360(.din(lo010_buf_o2), .dout(new_new_n1299__));
  not1  g0361(.din(lo010_buf_o2), .dout(new_new_n1300__));
  buf1  g0362(.din(lo166_buf_o2), .dout(new_new_n1301__));
  not1  g0363(.din(lo166_buf_o2), .dout(new_new_n1302__));
  buf1  g0364(.din(lo170_buf_o2), .dout(new_new_n1303__));
  not1  g0365(.din(lo170_buf_o2), .dout(new_new_n1304__));
  buf1  g0366(.din(n1426_o2), .dout(new_new_n1305__));
  not1  g0367(.din(n1426_o2), .dout(new_new_n1306__));
  buf1  g0368(.din(n1082_o2), .dout(new_new_n1307__));
  not1  g0369(.din(n1082_o2), .dout(new_new_n1308__));
  not1  g0370(.din(n1310_o2), .dout(new_new_n1310__));
  buf1  g0371(.din(n1015_o2), .dout(new_new_n1311__));
  not1  g0372(.din(n1015_o2), .dout(new_new_n1312__));
  buf1  g0373(.din(n1206_o2), .dout(new_new_n1313__));
  not1  g0374(.din(n1262_o2), .dout(new_new_n1316__));
  buf1  g0375(.din(n1456_o2), .dout(new_new_n1317__));
  not1  g0376(.din(n1456_o2), .dout(new_new_n1318__));
  buf1  g0377(.din(n1244_o2), .dout(new_new_n1319__));
  not1  g0378(.din(n1244_o2), .dout(new_new_n1320__));
  buf1  g0379(.din(n1280_o2), .dout(new_new_n1321__));
  not1  g0380(.din(n1280_o2), .dout(new_new_n1322__));
  buf1  g0381(.din(n1290_o2), .dout(new_new_n1323__));
  not1  g0382(.din(n1290_o2), .dout(new_new_n1324__));
  buf1  g0383(.din(n1012_o2), .dout(new_new_n1325__));
  not1  g0384(.din(n1012_o2), .dout(new_new_n1326__));
  buf1  g0385(.din(n1074_o2), .dout(new_new_n1327__));
  not1  g0386(.din(n1074_o2), .dout(new_new_n1328__));
  buf1  g0387(.din(n1112_o2), .dout(new_new_n1329__));
  not1  g0388(.din(n1112_o2), .dout(new_new_n1330__));
  buf1  g0389(.din(n1212_o2), .dout(new_new_n1331__));
  not1  g0390(.din(n1212_o2), .dout(new_new_n1332__));
  buf1  g0391(.din(n1454_o2), .dout(new_new_n1333__));
  not1  g0392(.din(n1454_o2), .dout(new_new_n1334__));
  buf1  g0393(.din(n1182_o2), .dout(new_new_n1335__));
  not1  g0394(.din(n1182_o2), .dout(new_new_n1336__));
  buf1  g0395(.din(n1220_o2), .dout(new_new_n1337__));
  not1  g0396(.din(n1220_o2), .dout(new_new_n1338__));
  buf1  g0397(.din(n701_o2), .dout(new_new_n1339__));
  buf1  g0398(.din(n744_inv), .dout(new_new_n1341__));
  buf1  g0399(.din(n1282_o2), .dout(new_new_n1343__));
  not1  g0400(.din(n1282_o2), .dout(new_new_n1344__));
  buf1  g0401(.din(n1144_o2), .dout(new_new_n1345__));
  buf1  g0402(.din(n1278_o2), .dout(new_new_n1347__));
  not1  g0403(.din(n1278_o2), .dout(new_new_n1348__));
  buf1  g0404(.din(n1459_o2), .dout(new_new_n1349__));
  not1  g0405(.din(n1459_o2), .dout(new_new_n1350__));
  buf1  g0406(.din(n1324_o2), .dout(new_new_n1351__));
  not1  g0407(.din(n1324_o2), .dout(new_new_n1352__));
  buf1  g0408(.din(n1288_o2), .dout(new_new_n1353__));
  not1  g0409(.din(n1288_o2), .dout(new_new_n1354__));
  not1  g0410(.din(n1271_o2), .dout(new_new_n1356__));
  buf1  g0411(.din(n1132_o2), .dout(new_new_n1357__));
  not1  g0412(.din(n1132_o2), .dout(new_new_n1358__));
  buf1  g0413(.din(n1231_o2), .dout(new_new_n1359__));
  not1  g0414(.din(n1231_o2), .dout(new_new_n1360__));
  buf1  g0415(.din(n1462_o2), .dout(new_new_n1361__));
  not1  g0416(.din(n1462_o2), .dout(new_new_n1362__));
  buf1  g0417(.din(n1482_o2), .dout(new_new_n1363__));
  not1  g0418(.din(n1482_o2), .dout(new_new_n1364__));
  buf1  g0419(.din(n994_o2), .dout(new_new_n1365__));
  not1  g0420(.din(n994_o2), .dout(new_new_n1366__));
  buf1  g0421(.din(n998_o2), .dout(new_new_n1367__));
  not1  g0422(.din(n998_o2), .dout(new_new_n1368__));
  buf1  g0423(.din(lo106_buf_o2), .dout(new_new_n1369__));
  buf1  g0424(.din(n769_o2), .dout(new_new_n1371__));
  not1  g0425(.din(n769_o2), .dout(new_new_n1372__));
  buf1  g0426(.din(n814_o2), .dout(new_new_n1373__));
  not1  g0427(.din(n814_o2), .dout(new_new_n1374__));
  buf1  g0428(.din(n841_o2), .dout(new_new_n1375__));
  not1  g0429(.din(n841_o2), .dout(new_new_n1376__));
  buf1  g0430(.din(n867_o2), .dout(new_new_n1377__));
  buf1  g0431(.din(lo006_buf_o2), .dout(new_new_n1379__));
  buf1  g0432(.din(lo014_buf_o2), .dout(new_new_n1381__));
  not1  g0433(.din(lo014_buf_o2), .dout(new_new_n1382__));
  buf1  g0434(.din(lo022_buf_o2), .dout(new_new_n1383__));
  not1  g0435(.din(lo022_buf_o2), .dout(new_new_n1384__));
  buf1  g0436(.din(lo042_buf_o2), .dout(new_new_n1385__));
  not1  g0437(.din(lo042_buf_o2), .dout(new_new_n1386__));
  buf1  g0438(.din(lo046_buf_o2), .dout(new_new_n1387__));
  not1  g0439(.din(lo046_buf_o2), .dout(new_new_n1388__));
  buf1  g0440(.din(lo050_buf_o2), .dout(new_new_n1389__));
  not1  g0441(.din(lo050_buf_o2), .dout(new_new_n1390__));
  buf1  g0442(.din(lo054_buf_o2), .dout(new_new_n1391__));
  not1  g0443(.din(lo054_buf_o2), .dout(new_new_n1392__));
  buf1  g0444(.din(lo130_buf_o2), .dout(new_new_n1393__));
  not1  g0445(.din(lo130_buf_o2), .dout(new_new_n1394__));
  buf1  g0446(.din(lo134_buf_o2), .dout(new_new_n1395__));
  buf1  g0447(.din(lo154_buf_o2), .dout(new_new_n1397__));
  not1  g0448(.din(lo154_buf_o2), .dout(new_new_n1398__));
  buf1  g0449(.din(lo174_buf_o2), .dout(new_new_n1399__));
  not1  g0450(.din(lo174_buf_o2), .dout(new_new_n1400__));
  buf1  g0451(.din(lo178_buf_o2), .dout(new_new_n1401__));
  not1  g0452(.din(lo178_buf_o2), .dout(new_new_n1402__));
  buf1  g0453(.din(n1007_o2), .dout(new_new_n1403__));
  not1  g0454(.din(n1007_o2), .dout(new_new_n1404__));
  not1  g0455(.din(n1294_o2), .dout(new_new_n1406__));
  not1  g0456(.din(n1084_o2), .dout(new_new_n1408__));
  not1  g0457(.din(n1399_o2), .dout(new_new_n1410__));
  buf1  g0458(.din(n1311_o2), .dout(new_new_n1411__));
  not1  g0459(.din(n1392_o2), .dout(new_new_n1414__));
  buf1  g0460(.din(n1102_o2), .dout(new_new_n1415__));
  not1  g0461(.din(n1102_o2), .dout(new_new_n1416__));
  buf1  g0462(.din(n1041_o2), .dout(new_new_n1417__));
  not1  g0463(.din(n1041_o2), .dout(new_new_n1418__));
  not1  g0464(.din(n1298_o2), .dout(new_new_n1420__));
  buf1  g0465(.din(n738_o2), .dout(new_new_n1421__));
  not1  g0466(.din(n738_o2), .dout(new_new_n1422__));
  buf1  g0467(.din(n1214_o2), .dout(new_new_n1423__));
  not1  g0468(.din(n1214_o2), .dout(new_new_n1424__));
  buf1  g0469(.din(n1222_o2), .dout(new_new_n1425__));
  not1  g0470(.din(n1222_o2), .dout(new_new_n1426__));
  buf1  g0471(.din(n1155_o2), .dout(new_new_n1427__));
  not1  g0472(.din(n1155_o2), .dout(new_new_n1428__));
  buf1  g0473(.din(n1147_o2), .dout(new_new_n1429__));
  not1  g0474(.din(n1147_o2), .dout(new_new_n1430__));
  buf1  g0475(.din(n1393_o2), .dout(new_new_n1431__));
  buf1  g0476(.din(n999_o2), .dout(new_new_n1433__));
  not1  g0477(.din(n999_o2), .dout(new_new_n1434__));
  buf1  g0478(.din(n1306_o2), .dout(new_new_n1435__));
  buf1  g0479(.din(n1312_o2), .dout(new_new_n1437__));
  buf1  g0480(.din(n1382_o2), .dout(new_new_n1439__));
  not1  g0481(.din(n1382_o2), .dout(new_new_n1440__));
  buf1  g0482(.din(n1383_o2), .dout(new_new_n1441__));
  not1  g0483(.din(n1383_o2), .dout(new_new_n1442__));
  buf1  g0484(.din(n1152_o2), .dout(new_new_n1443__));
  not1  g0485(.din(n1152_o2), .dout(new_new_n1444__));
  buf1  g0486(.din(n1334_o2), .dout(new_new_n1445__));
  not1  g0487(.din(n1334_o2), .dout(new_new_n1446__));
  buf1  g0488(.din(n1335_o2), .dout(new_new_n1447__));
  not1  g0489(.din(n1335_o2), .dout(new_new_n1448__));
  buf1  g0490(.din(n906_inv), .dout(new_new_n1449__));
  buf1  g0491(.din(n773_o2), .dout(new_new_n1451__));
  not1  g0492(.din(n773_o2), .dout(new_new_n1452__));
  buf1  g0493(.din(lo190_buf_o2), .dout(new_new_n1453__));
  not1  g0494(.din(n1368_o2), .dout(new_new_n1456__));
  not1  g0495(.din(n1362_o2), .dout(new_new_n1458__));
  not1  g0496(.din(n1406_o2), .dout(new_new_n1460__));
  not1  g0497(.din(n1403_o2), .dout(new_new_n1462__));
  buf1  g0498(.din(n741_o2), .dout(new_new_n1463__));
  not1  g0499(.din(n741_o2), .dout(new_new_n1464__));
  not1  g0500(.din(n1407_o2), .dout(new_new_n1466__));
  buf1  g0501(.din(n1395_o2), .dout(new_new_n1467__));
  buf1  g0502(.din(n1359_o2), .dout(new_new_n1469__));
  buf1  g0503(.din(n1159_o2), .dout(new_new_n1471__));
  not1  g0504(.din(n1159_o2), .dout(new_new_n1472__));
  buf1  g0505(.din(n1221_o2), .dout(new_new_n1473__));
  not1  g0506(.din(n1221_o2), .dout(new_new_n1474__));
  buf1  g0507(.din(n945_inv), .dout(new_new_n1475__));
  not1  g0508(.din(n945_inv), .dout(new_new_n1476__));
  buf1  g0509(.din(n989_o2), .dout(new_new_n1477__));
  not1  g0510(.din(n989_o2), .dout(new_new_n1478__));
  buf1  g0511(.din(n881_o2), .dout(new_new_n1479__));
  not1  g0512(.din(n881_o2), .dout(new_new_n1480__));
  buf1  g0513(.din(n1340_o2), .dout(new_new_n1481__));
  not1  g0514(.din(n1340_o2), .dout(new_new_n1482__));
  buf1  g0515(.din(n1341_o2), .dout(new_new_n1483__));
  not1  g0516(.din(n1341_o2), .dout(new_new_n1484__));
  buf1  g0517(.din(n906_o2), .dout(new_new_n1485__));
  not1  g0518(.din(n906_o2), .dout(new_new_n1486__));
  buf1  g0519(.din(n1388_o2), .dout(new_new_n1487__));
  buf1  g0520(.din(n791_o2), .dout(new_new_n1489__));
  not1  g0521(.din(n791_o2), .dout(new_new_n1490__));
  not1  g0522(.din(n1372_o2), .dout(new_new_n1492__));
  buf1  g0523(.din(n815_o2), .dout(new_new_n1493__));
  not1  g0524(.din(n815_o2), .dout(new_new_n1494__));
  buf1  g0525(.din(n868_o2), .dout(new_new_n1495__));
  not1  g0526(.din(n868_o2), .dout(new_new_n1496__));
  buf1  g0527(.din(lo018_buf_o2), .dout(new_new_n1497__));
  not1  g0528(.din(lo018_buf_o2), .dout(new_new_n1498__));
  buf1  g0529(.din(lo138_buf_o2), .dout(new_new_n1499__));
  not1  g0530(.din(lo138_buf_o2), .dout(new_new_n1500__));
  buf1  g0531(.din(lo158_buf_o2), .dout(new_new_n1501__));
  buf1  g0532(.din(n780_o2), .dout(new_new_n1503__));
  not1  g0533(.din(n780_o2), .dout(new_new_n1504__));
  buf1  g0534(.din(n728_o2), .dout(new_new_n1505__));
  buf1  g0535(.din(n993_inv), .dout(new_new_n1507__));
  buf1  g0536(.din(n929_o2), .dout(new_new_n1509__));
  not1  g0537(.din(n929_o2), .dout(new_new_n1510__));
  buf1  g0538(.din(n955_o2), .dout(new_new_n1511__));
  not1  g0539(.din(n955_o2), .dout(new_new_n1512__));
  buf1  g0540(.din(n938_o2), .dout(new_new_n1513__));
  not1  g0541(.din(n938_o2), .dout(new_new_n1514__));
  buf1  g0542(.din(n1117_o2), .dout(new_new_n1515__));
  not1  g0543(.din(n1117_o2), .dout(new_new_n1516__));
  buf1  g0544(.din(n1121_o2), .dout(new_new_n1517__));
  not1  g0545(.din(n1121_o2), .dout(new_new_n1518__));
  buf1  g0546(.din(n965_o2), .dout(new_new_n1519__));
  not1  g0547(.din(n965_o2), .dout(new_new_n1520__));
  buf1  g0548(.din(n752_o2), .dout(new_new_n1521__));
  buf1  g0549(.din(n753_o2), .dout(new_new_n1523__));
  not1  g0550(.din(n753_o2), .dout(new_new_n1524__));
  buf1  g0551(.din(n760_o2), .dout(new_new_n1525__));
  not1  g0552(.din(n760_o2), .dout(new_new_n1526__));
  buf1  g0553(.din(n770_o2), .dout(new_new_n1527__));
  buf1  g0554(.din(n923_o2), .dout(new_new_n1529__));
  not1  g0555(.din(n923_o2), .dout(new_new_n1530__));
  buf1  g0556(.din(n947_o2), .dout(new_new_n1531__));
  not1  g0557(.din(n947_o2), .dout(new_new_n1532__));
  buf1  g0558(.din(n897_o2), .dout(new_new_n1533__));
  not1  g0559(.din(n897_o2), .dout(new_new_n1534__));
  buf1  g0560(.din(n919_o2), .dout(new_new_n1535__));
  not1  g0561(.din(n919_o2), .dout(new_new_n1536__));
  buf1  g0562(.din(n895_o2), .dout(new_new_n1537__));
  not1  g0563(.din(n895_o2), .dout(new_new_n1538__));
  buf1  g0564(.din(n917_o2), .dout(new_new_n1539__));
  not1  g0565(.din(n917_o2), .dout(new_new_n1540__));
  buf1  g0566(.din(n751_o2), .dout(new_new_n1541__));
  not1  g0567(.din(n751_o2), .dout(new_new_n1542__));
  buf1  g0568(.din(n774_o2), .dout(new_new_n1543__));
  not1  g0569(.din(n774_o2), .dout(new_new_n1544__));
  buf1  g0570(.din(lo126_buf_o2), .dout(new_new_n1545__));
  not1  g0571(.din(lo126_buf_o2), .dout(new_new_n1546__));
  buf1  g0572(.din(lo142_buf_o2), .dout(new_new_n1547__));
  not1  g0573(.din(lo142_buf_o2), .dout(new_new_n1548__));
  buf1  g0574(.din(lo162_buf_o2), .dout(new_new_n1549__));
  buf1  g0575(.din(n1059_inv), .dout(new_new_n1551__));
  not1  g0576(.din(n1059_inv), .dout(new_new_n1552__));
  buf1  g0577(.din(n792_o2), .dout(new_new_n1553__));
  not1  g0578(.din(n792_o2), .dout(new_new_n1554__));
  buf1  g0579(.din(n869_o2), .dout(new_new_n1555__));
  not1  g0580(.din(n869_o2), .dout(new_new_n1556__));
  buf1  g0581(.din(n1068_inv), .dout(new_new_n1557__));
  buf1  g0582(.din(lo024_buf_o2), .dout(new_new_n1559__));
  not1  g0583(.din(lo024_buf_o2), .dout(new_new_n1560__));
  buf1  g0584(.din(lo028_buf_o2), .dout(new_new_n1561__));
  not1  g0585(.din(lo028_buf_o2), .dout(new_new_n1562__));
  buf1  g0586(.din(lo088_buf_o2), .dout(new_new_n1563__));
  not1  g0587(.din(lo088_buf_o2), .dout(new_new_n1564__));
  buf1  g0588(.din(lo092_buf_o2), .dout(new_new_n1565__));
  not1  g0589(.din(lo092_buf_o2), .dout(new_new_n1566__));
  buf1  g0590(.din(lo096_buf_o2), .dout(new_new_n1567__));
  buf1  g0591(.din(lo100_buf_o2), .dout(new_new_n1569__));
  buf1  g0592(.din(n763_o2), .dout(new_new_n1571__));
  not1  g0593(.din(n763_o2), .dout(new_new_n1572__));
  buf1  g0594(.din(n754_o2), .dout(new_new_n1573__));
  not1  g0595(.din(n754_o2), .dout(new_new_n1574__));
  buf1  g0596(.din(n755_o2), .dout(new_new_n1575__));
  not1  g0597(.din(n755_o2), .dout(new_new_n1576__));
  buf1  g0598(.din(n822_o2), .dout(new_new_n1577__));
  not1  g0599(.din(n822_o2), .dout(new_new_n1578__));
  buf1  g0600(.din(n849_o2), .dout(new_new_n1579__));
  not1  g0601(.din(n849_o2), .dout(new_new_n1580__));
  buf1  g0602(.din(n777_o2), .dout(new_new_n1581__));
  not1  g0603(.din(n777_o2), .dout(new_new_n1582__));
  buf1  g0604(.din(n778_o2), .dout(new_new_n1583__));
  not1  g0605(.din(n778_o2), .dout(new_new_n1584__));
  buf1  g0606(.din(n820_o2), .dout(new_new_n1585__));
  not1  g0607(.din(n820_o2), .dout(new_new_n1586__));
  buf1  g0608(.din(n846_o2), .dout(new_new_n1587__));
  not1  g0609(.din(n846_o2), .dout(new_new_n1588__));
  buf1  g0610(.din(n806_o2), .dout(new_new_n1589__));
  not1  g0611(.din(n806_o2), .dout(new_new_n1590__));
  buf1  g0612(.din(n771_o2), .dout(new_new_n1591__));
  not1  g0613(.din(n771_o2), .dout(new_new_n1592__));
  buf1  g0614(.din(n854_o2), .dout(new_new_n1593__));
  not1  g0615(.din(n854_o2), .dout(new_new_n1594__));
  buf1  g0616(.din(n828_o2), .dout(new_new_n1595__));
  not1  g0617(.din(n828_o2), .dout(new_new_n1596__));
  buf1  g0618(.din(lo117_buf_o2), .dout(new_new_n1597__));
  not1  g0619(.din(lo117_buf_o2), .dout(new_new_n1598__));
  buf1  g0620(.din(lo145_buf_o2), .dout(new_new_n1599__));
  not1  g0621(.din(lo145_buf_o2), .dout(new_new_n1600__));
  buf1  g0622(.din(n762_o2), .dout(new_new_n1601__));
  not1  g0623(.din(n762_o2), .dout(new_new_n1602__));
  buf1  g0624(.din(n805_o2), .dout(new_new_n1603__));
  not1  g0625(.din(n805_o2), .dout(new_new_n1604__));
  buf1  g0626(.din(n859_o2), .dout(new_new_n1605__));
  not1  g0627(.din(n859_o2), .dout(new_new_n1606__));
  buf1  g0628(.din(n833_o2), .dout(new_new_n1607__));
  not1  g0629(.din(n833_o2), .dout(new_new_n1608__));
  buf1  g0630(.din(lo034_buf_o2), .dout(new_new_n1609__));
  not1  g0631(.din(lo034_buf_o2), .dout(new_new_n1610__));
  buf1  g0632(.din(lo038_buf_o2), .dout(new_new_n1611__));
  not1  g0633(.din(lo038_buf_o2), .dout(new_new_n1612__));
  buf1  g0634(.din(lo122_buf_o2), .dout(new_new_n1613__));
  not1  g0635(.din(lo122_buf_o2), .dout(new_new_n1614__));
  buf1  g0636(.din(lo150_buf_o2), .dout(new_new_n1615__));
  not1  g0637(.din(lo150_buf_o2), .dout(new_new_n1616__));
  and1  g0638(.dina(new_new_n1014__), .dinb(new_new_n3063__), .dout(new_new_n1617__));
  and1  g0639(.dina(new_new_n3064__), .dinb(new_new_n3065__), .dout(new_new_n1618__));
  or1   g0640(.dina(new_new_n3067__), .dinb(new_new_n3069__), .dout(new_new_n1619__));
  or1   g0641(.dina(new_new_n3071__), .dinb(new_new_n903__), .dout(new_new_n1620__));
  and1  g0642(.dina(new_new_n1620__), .dinb(new_new_n1619__), .dout(new_new_n1621__));
  or1   g0643(.dina(new_new_n3073__), .dinb(new_new_n3074__), .dout(new_new_n1622__));
  or1   g0644(.dina(new_new_n3076__), .dinb(new_new_n905__), .dout(new_new_n1623__));
  and1  g0645(.dina(new_new_n1623__), .dinb(new_new_n1622__), .dout(new_new_n1624__));
  and1  g0646(.dina(new_new_n1624__), .dinb(new_new_n1621__), .dout(new_new_n1625__));
  or1   g0647(.dina(new_new_n3078__), .dinb(new_new_n3080__), .dout(new_new_n1626__));
  or1   g0648(.dina(new_new_n3082__), .dinb(new_new_n901__), .dout(new_new_n1627__));
  and1  g0649(.dina(new_new_n1627__), .dinb(new_new_n1626__), .dout(new_new_n1628__));
  or1   g0650(.dina(new_new_n3084__), .dinb(new_new_n3086__), .dout(new_new_n1629__));
  or1   g0651(.dina(new_new_n3088__), .dinb(new_new_n3091__), .dout(new_new_n1630__));
  and1  g0652(.dina(new_new_n1630__), .dinb(new_new_n1629__), .dout(new_new_n1631__));
  and1  g0653(.dina(new_new_n1631__), .dinb(new_new_n1628__), .dout(new_new_n1632__));
  and1  g0654(.dina(new_new_n1632__), .dinb(new_new_n1625__), .dout(new_new_n1633__));
  or1   g0655(.dina(new_new_n1633__), .dinb(new_new_n1618__), .dout(new_new_n1634__));
  and1  g0656(.dina(new_new_n1007__), .dinb(new_new_n3064__), .dout(new_new_n1635__));
  or1   g0657(.dina(new_new_n1008__), .dinb(new_new_n897__), .dout(new_new_n1636__));
  or1   g0658(.dina(new_new_n3092__), .dinb(new_new_n1088__), .dout(new_new_n1637__));
  and1  g0659(.dina(new_new_n3088__), .dinb(new_new_n3084__), .dout(new_new_n1638__));
  or1   g0660(.dina(new_new_n1638__), .dinb(new_new_n3067__), .dout(new_new_n1639__));
  or1   g0661(.dina(new_new_n1639__), .dinb(new_new_n1019__), .dout(new_new_n1640__));
  and1  g0662(.dina(new_new_n1640__), .dinb(new_new_n1637__), .dout(new_new_n1641__));
  and1  g0663(.dina(new_new_n1641__), .dinb(new_new_n1634__), .dout(new_new_n1642__));
  and1  g0664(.dina(new_new_n3078__), .dinb(new_new_n3093__), .dout(new_new_n1643__));
  or1   g0665(.dina(new_new_n3094__), .dinb(new_new_n3089__), .dout(new_new_n1644__));
  and1  g0666(.dina(new_new_n3094__), .dinb(new_new_n3089__), .dout(new_new_n1645__));
  or1   g0667(.dina(new_new_n3077__), .dinb(new_new_n3093__), .dout(new_new_n1646__));
  and1  g0668(.dina(new_new_n1646__), .dinb(new_new_n1644__), .dout(new_new_n1647__));
  or1   g0669(.dina(new_new_n1645__), .dinb(new_new_n1643__), .dout(new_new_n1648__));
  and1  g0670(.dina(new_new_n3085__), .dinb(new_new_n3095__), .dout(new_new_n1649__));
  or1   g0671(.dina(new_new_n3096__), .dinb(new_new_n3068__), .dout(new_new_n1650__));
  and1  g0672(.dina(new_new_n3096__), .dinb(new_new_n3068__), .dout(new_new_n1651__));
  or1   g0673(.dina(new_new_n3085__), .dinb(new_new_n3095__), .dout(new_new_n1652__));
  and1  g0674(.dina(new_new_n1652__), .dinb(new_new_n1650__), .dout(new_new_n1653__));
  or1   g0675(.dina(new_new_n1651__), .dinb(new_new_n1649__), .dout(new_new_n1654__));
  and1  g0676(.dina(new_new_n3097__), .dinb(new_new_n3098__), .dout(new_new_n1655__));
  or1   g0677(.dina(new_new_n3099__), .dinb(new_new_n3100__), .dout(new_new_n1656__));
  and1  g0678(.dina(new_new_n3099__), .dinb(new_new_n3100__), .dout(new_new_n1657__));
  or1   g0679(.dina(new_new_n3097__), .dinb(new_new_n3098__), .dout(new_new_n1658__));
  and1  g0680(.dina(new_new_n1658__), .dinb(new_new_n1656__), .dout(new_new_n1659__));
  or1   g0681(.dina(new_new_n1657__), .dinb(new_new_n1655__), .dout(new_new_n1660__));
  and1  g0682(.dina(new_new_n3076__), .dinb(new_new_n3101__), .dout(new_new_n1661__));
  or1   g0683(.dina(new_new_n3102__), .dinb(new_new_n3071__), .dout(new_new_n1662__));
  and1  g0684(.dina(new_new_n3102__), .dinb(new_new_n3070__), .dout(new_new_n1663__));
  or1   g0685(.dina(new_new_n3075__), .dinb(new_new_n3101__), .dout(new_new_n1664__));
  and1  g0686(.dina(new_new_n1664__), .dinb(new_new_n1662__), .dout(new_new_n1665__));
  or1   g0687(.dina(new_new_n1663__), .dinb(new_new_n1661__), .dout(new_new_n1666__));
  and1  g0688(.dina(new_new_n3082__), .dinb(new_new_n3103__), .dout(new_new_n1667__));
  or1   g0689(.dina(new_new_n3104__), .dinb(new_new_n3073__), .dout(new_new_n1668__));
  and1  g0690(.dina(new_new_n3104__), .dinb(new_new_n3072__), .dout(new_new_n1669__));
  or1   g0691(.dina(new_new_n3081__), .dinb(new_new_n3103__), .dout(new_new_n1670__));
  and1  g0692(.dina(new_new_n1670__), .dinb(new_new_n1668__), .dout(new_new_n1671__));
  or1   g0693(.dina(new_new_n1669__), .dinb(new_new_n1667__), .dout(new_new_n1672__));
  and1  g0694(.dina(new_new_n3105__), .dinb(new_new_n3106__), .dout(new_new_n1673__));
  or1   g0695(.dina(new_new_n3107__), .dinb(new_new_n3108__), .dout(new_new_n1674__));
  and1  g0696(.dina(new_new_n3107__), .dinb(new_new_n3108__), .dout(new_new_n1675__));
  or1   g0697(.dina(new_new_n3105__), .dinb(new_new_n3106__), .dout(new_new_n1676__));
  and1  g0698(.dina(new_new_n1676__), .dinb(new_new_n1674__), .dout(new_new_n1677__));
  or1   g0699(.dina(new_new_n1675__), .dinb(new_new_n1673__), .dout(new_new_n1678__));
  or1   g0700(.dina(new_new_n1677__), .dinb(new_new_n1659__), .dout(new_new_n1679__));
  or1   g0701(.dina(new_new_n1678__), .dinb(new_new_n1660__), .dout(new_new_n1680__));
  and1  g0702(.dina(new_new_n1680__), .dinb(new_new_n1679__), .dout(new_new_n1681__));
  and1  g0703(.dina(new_new_n3086__), .dinb(new_new_n3069__), .dout(new_new_n1682__));
  or1   g0704(.dina(new_new_n910__), .dinb(new_new_n908__), .dout(new_new_n1683__));
  and1  g0705(.dina(new_new_n1683__), .dinb(new_new_n1009__), .dout(new_new_n1684__));
  or1   g0706(.dina(new_new_n1682__), .dinb(new_new_n1010__), .dout(new_new_n1685__));
  and1  g0707(.dina(new_new_n3110__), .dinb(new_new_n3091__), .dout(new_new_n1686__));
  or1   g0708(.dina(new_new_n3080__), .dinb(new_new_n3111__), .dout(new_new_n1687__));
  and1  g0709(.dina(new_new_n3079__), .dinb(new_new_n3111__), .dout(new_new_n1688__));
  or1   g0710(.dina(new_new_n3110__), .dinb(new_new_n3090__), .dout(new_new_n1689__));
  and1  g0711(.dina(new_new_n1689__), .dinb(new_new_n1687__), .dout(new_new_n1690__));
  or1   g0712(.dina(new_new_n1688__), .dinb(new_new_n1686__), .dout(new_new_n1691__));
  and1  g0713(.dina(new_new_n3112__), .dinb(new_new_n3113__), .dout(new_new_n1692__));
  or1   g0714(.dina(new_new_n3114__), .dinb(new_new_n3115__), .dout(new_new_n1693__));
  and1  g0715(.dina(new_new_n3114__), .dinb(new_new_n3115__), .dout(new_new_n1694__));
  or1   g0716(.dina(new_new_n3112__), .dinb(new_new_n3113__), .dout(new_new_n1695__));
  and1  g0717(.dina(new_new_n1695__), .dinb(new_new_n1693__), .dout(new_new_n1696__));
  or1   g0718(.dina(new_new_n1694__), .dinb(new_new_n1692__), .dout(new_new_n1697__));
  and1  g0719(.dina(new_new_n1697__), .dinb(new_new_n1112__), .dout(new_new_n1698__));
  and1  g0720(.dina(new_new_n1696__), .dinb(new_new_n1111__), .dout(new_new_n1699__));
  or1   g0721(.dina(new_new_n1699__), .dinb(new_new_n1698__), .dout(new_new_n1700__));
  and1  g0722(.dina(new_new_n3116__), .dinb(new_new_n1021__), .dout(new_new_n1701__));
  and1  g0723(.dina(new_new_n3116__), .dinb(new_new_n1023__), .dout(new_new_n1702__));
  or1   g0724(.dina(new_new_n1702__), .dinb(new_new_n1077__), .dout(new_new_n1703__));
  and1  g0725(.dina(new_new_n3118__), .dinb(new_new_n1087__), .dout(new_new_n1704__));
  and1  g0726(.dina(new_new_n1027__), .dinb(new_new_n3065__), .dout(new_new_n1705__));
  or1   g0727(.dina(new_new_n1705__), .dinb(new_new_n1704__), .dout(new_new_n1706__));
  and1  g0728(.dina(new_new_n1326__), .dinb(new_new_n3119__), .dout(new_new_n1707__));
  or1   g0729(.dina(new_new_n1325__), .dinb(new_new_n3120__), .dout(new_new_n1708__));
  and1  g0730(.dina(new_new_n1327__), .dinb(new_new_n1312__), .dout(new_new_n1709__));
  or1   g0731(.dina(new_new_n1328__), .dinb(new_new_n1311__), .dout(new_new_n1710__));
  and1  g0732(.dina(new_new_n1710__), .dinb(new_new_n1708__), .dout(new_new_n1711__));
  or1   g0733(.dina(new_new_n1709__), .dinb(new_new_n1707__), .dout(new_new_n1712__));
  and1  g0734(.dina(new_new_n1329__), .dinb(new_new_n1308__), .dout(new_new_n1713__));
  or1   g0735(.dina(new_new_n1330__), .dinb(new_new_n1307__), .dout(new_new_n1714__));
  and1  g0736(.dina(new_new_n1357__), .dinb(new_new_n3119__), .dout(new_new_n1715__));
  or1   g0737(.dina(new_new_n1358__), .dinb(new_new_n3120__), .dout(new_new_n1716__));
  and1  g0738(.dina(new_new_n1716__), .dinb(new_new_n1714__), .dout(new_new_n1717__));
  or1   g0739(.dina(new_new_n1715__), .dinb(new_new_n1713__), .dout(new_new_n1718__));
  and1  g0740(.dina(new_new_n1055__), .dinb(new_new_n1025__), .dout(new_new_n1719__));
  or1   g0741(.dina(new_new_n1056__), .dinb(new_new_n1026__), .dout(new_new_n1720__));
  and1  g0742(.dina(new_new_n3121__), .dinb(new_new_n3122__), .dout(new_new_n1721__));
  or1   g0743(.dina(new_new_n3123__), .dinb(new_new_n3124__), .dout(new_new_n1722__));
  and1  g0744(.dina(new_new_n3123__), .dinb(new_new_n3124__), .dout(new_new_n1723__));
  or1   g0745(.dina(new_new_n3121__), .dinb(new_new_n3122__), .dout(new_new_n1724__));
  and1  g0746(.dina(new_new_n1724__), .dinb(new_new_n1722__), .dout(new_new_n1725__));
  or1   g0747(.dina(new_new_n1723__), .dinb(new_new_n1721__), .dout(new_new_n1726__));
  and1  g0748(.dina(new_new_n1726__), .dinb(new_new_n993__), .dout(new_new_n1727__));
  or1   g0749(.dina(new_new_n1725__), .dinb(new_new_n994__), .dout(new_new_n1728__));
  and1  g0750(.dina(new_new_n3125__), .dinb(new_new_n3126__), .dout(new_new_n1729__));
  or1   g0751(.dina(new_new_n3127__), .dinb(new_new_n3128__), .dout(new_new_n1730__));
  and1  g0752(.dina(new_new_n3127__), .dinb(new_new_n3128__), .dout(new_new_n1731__));
  or1   g0753(.dina(new_new_n3125__), .dinb(new_new_n3126__), .dout(new_new_n1732__));
  and1  g0754(.dina(new_new_n1732__), .dinb(new_new_n1730__), .dout(new_new_n1733__));
  or1   g0755(.dina(new_new_n1731__), .dinb(new_new_n1729__), .dout(new_new_n1734__));
  and1  g0756(.dina(new_new_n1733__), .dinb(new_new_n1727__), .dout(new_new_n1735__));
  and1  g0757(.dina(new_new_n1734__), .dinb(new_new_n1728__), .dout(new_new_n1736__));
  or1   g0758(.dina(new_new_n1736__), .dinb(new_new_n1735__), .dout(new_new_n1737__));
  and1  g0759(.dina(new_new_n3092__), .dinb(new_new_n1017__), .dout(new_new_n1738__));
  and1  g0760(.dina(new_new_n1738__), .dinb(new_new_n1737__), .dout(new_new_n1739__));
  and1  g0761(.dina(new_new_n1635__), .dinb(new_new_n3109__), .dout(new_new_n1740__));
  and1  g0762(.dina(new_new_n1740__), .dinb(new_new_n1012__), .dout(new_new_n1741__));
  and1  g0763(.dina(new_new_n1016__), .dinb(new_new_n3063__), .dout(new_new_n1742__));
  or1   g0764(.dina(new_new_n1742__), .dinb(new_new_n3074__), .dout(new_new_n1743__));
  or1   g0765(.dina(new_new_n904__), .dinb(new_new_n900__), .dout(new_new_n1744__));
  and1  g0766(.dina(new_new_n1744__), .dinb(new_new_n1018__), .dout(new_new_n1745__));
  and1  g0767(.dina(new_new_n1745__), .dinb(new_new_n1743__), .dout(new_new_n1746__));
  or1   g0768(.dina(new_new_n1746__), .dinb(new_new_n1741__), .dout(new_new_n1747__));
  or1   g0769(.dina(new_new_n1747__), .dinb(new_new_n1739__), .dout(new_new_n1748__));
  and1  g0770(.dina(new_new_n1336__), .dinb(new_new_n1331__), .dout(new_new_n1749__));
  or1   g0771(.dina(new_new_n1335__), .dinb(new_new_n1332__), .dout(new_new_n1750__));
  and1  g0772(.dina(new_new_n1359__), .dinb(new_new_n1320__), .dout(new_new_n1751__));
  or1   g0773(.dina(new_new_n1360__), .dinb(new_new_n1319__), .dout(new_new_n1752__));
  and1  g0774(.dina(new_new_n1752__), .dinb(new_new_n1750__), .dout(new_new_n1753__));
  or1   g0775(.dina(new_new_n1751__), .dinb(new_new_n1749__), .dout(new_new_n1754__));
  and1  g0776(.dina(new_new_n1343__), .dinb(new_new_n3118__), .dout(new_new_n1755__));
  or1   g0777(.dina(new_new_n1344__), .dinb(new_new_n3129__), .dout(new_new_n1756__));
  and1  g0778(.dina(new_new_n1348__), .dinb(new_new_n1322__), .dout(new_new_n1757__));
  or1   g0779(.dina(new_new_n1347__), .dinb(new_new_n1321__), .dout(new_new_n1758__));
  and1  g0780(.dina(new_new_n1757__), .dinb(new_new_n1756__), .dout(new_new_n1759__));
  or1   g0781(.dina(new_new_n1758__), .dinb(new_new_n1755__), .dout(new_new_n1760__));
  and1  g0782(.dina(new_new_n1353__), .dinb(new_new_n3117__), .dout(new_new_n1761__));
  or1   g0783(.dina(new_new_n1354__), .dinb(new_new_n3129__), .dout(new_new_n1762__));
  and1  g0784(.dina(new_new_n1352__), .dinb(new_new_n1324__), .dout(new_new_n1763__));
  or1   g0785(.dina(new_new_n1351__), .dinb(new_new_n1323__), .dout(new_new_n1764__));
  and1  g0786(.dina(new_new_n1763__), .dinb(new_new_n1762__), .dout(new_new_n1765__));
  or1   g0787(.dina(new_new_n1764__), .dinb(new_new_n1761__), .dout(new_new_n1766__));
  and1  g0788(.dina(new_new_n1333__), .dinb(new_new_n1306__), .dout(new_new_n1767__));
  or1   g0789(.dina(new_new_n1334__), .dinb(new_new_n1305__), .dout(new_new_n1768__));
  and1  g0790(.dina(new_new_n1349__), .dinb(new_new_n1318__), .dout(new_new_n1769__));
  or1   g0791(.dina(new_new_n1350__), .dinb(new_new_n1317__), .dout(new_new_n1770__));
  and1  g0792(.dina(new_new_n1770__), .dinb(new_new_n1768__), .dout(new_new_n1771__));
  or1   g0793(.dina(new_new_n1769__), .dinb(new_new_n1767__), .dout(new_new_n1772__));
  and1  g0794(.dina(new_new_n3130__), .dinb(new_new_n3131__), .dout(new_new_n1773__));
  or1   g0795(.dina(new_new_n3133__), .dinb(new_new_n3135__), .dout(new_new_n1774__));
  and1  g0796(.dina(new_new_n3136__), .dinb(new_new_n3137__), .dout(new_new_n1775__));
  or1   g0797(.dina(new_new_n3139__), .dinb(new_new_n3141__), .dout(new_new_n1776__));
  and1  g0798(.dina(new_new_n3142__), .dinb(new_new_n3143__), .dout(new_new_n1777__));
  or1   g0799(.dina(new_new_n3145__), .dinb(new_new_n3147__), .dout(new_new_n1778__));
  or1   g0800(.dina(new_new_n3148__), .dinb(new_new_n3149__), .dout(new_new_n1779__));
  or1   g0801(.dina(new_new_n1779__), .dinb(new_new_n3150__), .dout(new_new_n1780__));
  or1   g0802(.dina(new_new_n1780__), .dinb(new_new_n3152__), .dout(new_new_n1781__));
  and1  g0803(.dina(new_new_n997__), .dinb(new_new_n3153__), .dout(new_new_n1782__));
  or1   g0804(.dina(new_new_n998__), .dinb(new_new_n946__), .dout(new_new_n1783__));
  or1   g0805(.dina(new_new_n3154__), .dinb(new_new_n3152__), .dout(new_new_n1784__));
  and1  g0806(.dina(new_new_n1784__), .dinb(new_new_n3153__), .dout(new_new_n1785__));
  and1  g0807(.dina(new_new_n1785__), .dinb(new_new_n3155__), .dout(new_new_n1786__));
  and1  g0808(.dina(new_new_n3145__), .dinb(new_new_n3147__), .dout(new_new_n1787__));
  or1   g0809(.dina(new_new_n3142__), .dinb(new_new_n3143__), .dout(new_new_n1788__));
  and1  g0810(.dina(new_new_n1788__), .dinb(new_new_n3148__), .dout(new_new_n1789__));
  or1   g0811(.dina(new_new_n1787__), .dinb(new_new_n1777__), .dout(new_new_n1790__));
  and1  g0812(.dina(new_new_n3139__), .dinb(new_new_n3141__), .dout(new_new_n1791__));
  or1   g0813(.dina(new_new_n3136__), .dinb(new_new_n3137__), .dout(new_new_n1792__));
  and1  g0814(.dina(new_new_n1792__), .dinb(new_new_n3149__), .dout(new_new_n1793__));
  or1   g0815(.dina(new_new_n1791__), .dinb(new_new_n1775__), .dout(new_new_n1794__));
  and1  g0816(.dina(new_new_n3156__), .dinb(new_new_n3157__), .dout(new_new_n1795__));
  or1   g0817(.dina(new_new_n3158__), .dinb(new_new_n3159__), .dout(new_new_n1796__));
  and1  g0818(.dina(new_new_n3158__), .dinb(new_new_n3159__), .dout(new_new_n1797__));
  or1   g0819(.dina(new_new_n3156__), .dinb(new_new_n3157__), .dout(new_new_n1798__));
  and1  g0820(.dina(new_new_n1798__), .dinb(new_new_n1796__), .dout(new_new_n1799__));
  or1   g0821(.dina(new_new_n1797__), .dinb(new_new_n1795__), .dout(new_new_n1800__));
  and1  g0822(.dina(new_new_n3133__), .dinb(new_new_n3135__), .dout(new_new_n1801__));
  or1   g0823(.dina(new_new_n3130__), .dinb(new_new_n3131__), .dout(new_new_n1802__));
  and1  g0824(.dina(new_new_n1802__), .dinb(new_new_n3150__), .dout(new_new_n1803__));
  or1   g0825(.dina(new_new_n1801__), .dinb(new_new_n1773__), .dout(new_new_n1804__));
  and1  g0826(.dina(new_new_n1364__), .dinb(new_new_n3151__), .dout(new_new_n1805__));
  or1   g0827(.dina(new_new_n1363__), .dinb(new_new_n1362__), .dout(new_new_n1806__));
  and1  g0828(.dina(new_new_n3161__), .dinb(new_new_n3163__), .dout(new_new_n1807__));
  or1   g0829(.dina(new_new_n3165__), .dinb(new_new_n3167__), .dout(new_new_n1808__));
  and1  g0830(.dina(new_new_n3165__), .dinb(new_new_n3167__), .dout(new_new_n1809__));
  or1   g0831(.dina(new_new_n3161__), .dinb(new_new_n3163__), .dout(new_new_n1810__));
  and1  g0832(.dina(new_new_n1810__), .dinb(new_new_n1808__), .dout(new_new_n1811__));
  or1   g0833(.dina(new_new_n1809__), .dinb(new_new_n1807__), .dout(new_new_n1812__));
  and1  g0834(.dina(new_new_n1812__), .dinb(new_new_n3154__), .dout(new_new_n1813__));
  or1   g0835(.dina(new_new_n1811__), .dinb(new_new_n1782__), .dout(new_new_n1814__));
  and1  g0836(.dina(new_new_n3168__), .dinb(new_new_n3170__), .dout(new_new_n1815__));
  or1   g0837(.dina(new_new_n3172__), .dinb(new_new_n3174__), .dout(new_new_n1816__));
  and1  g0838(.dina(new_new_n3172__), .dinb(new_new_n3174__), .dout(new_new_n1817__));
  or1   g0839(.dina(new_new_n3168__), .dinb(new_new_n3170__), .dout(new_new_n1818__));
  and1  g0840(.dina(new_new_n1818__), .dinb(new_new_n1816__), .dout(new_new_n1819__));
  or1   g0841(.dina(new_new_n1817__), .dinb(new_new_n1815__), .dout(new_new_n1820__));
  and1  g0842(.dina(new_new_n1820__), .dinb(new_new_n3176__), .dout(new_new_n1821__));
  and1  g0843(.dina(new_new_n1819__), .dinb(new_new_n3177__), .dout(new_new_n1822__));
  or1   g0844(.dina(new_new_n1822__), .dinb(new_new_n1821__), .dout(new_new_n1823__));
  and1  g0845(.dina(new_new_n3162__), .dinb(new_new_n3175__), .dout(new_new_n1824__));
  or1   g0846(.dina(new_new_n3166__), .dinb(new_new_n3171__), .dout(new_new_n1825__));
  and1  g0847(.dina(new_new_n3166__), .dinb(new_new_n3171__), .dout(new_new_n1826__));
  or1   g0848(.dina(new_new_n3162__), .dinb(new_new_n3175__), .dout(new_new_n1827__));
  and1  g0849(.dina(new_new_n1827__), .dinb(new_new_n1825__), .dout(new_new_n1828__));
  or1   g0850(.dina(new_new_n1826__), .dinb(new_new_n1824__), .dout(new_new_n1829__));
  or1   g0851(.dina(new_new_n1828__), .dinb(new_new_n3177__), .dout(new_new_n1830__));
  or1   g0852(.dina(new_new_n1829__), .dinb(new_new_n3176__), .dout(new_new_n1831__));
  and1  g0853(.dina(new_new_n1831__), .dinb(new_new_n1830__), .dout(new_new_n1832__));
  or1   g0854(.dina(new_new_n1110__), .dinb(new_new_n3179__), .dout(new_new_n1833__));
  or1   g0855(.dina(new_new_n1068__), .dinb(new_new_n3181__), .dout(new_new_n1834__));
  and1  g0856(.dina(new_new_n1433__), .dinb(new_new_n3183__), .dout(new_new_n1835__));
  or1   g0857(.dina(new_new_n1434__), .dinb(new_new_n3184__), .dout(new_new_n1836__));
  and1  g0858(.dina(new_new_n1472__), .dinb(new_new_n1428__), .dout(new_new_n1837__));
  or1   g0859(.dina(new_new_n1471__), .dinb(new_new_n1427__), .dout(new_new_n1838__));
  and1  g0860(.dina(new_new_n1476__), .dinb(new_new_n1443__), .dout(new_new_n1839__));
  or1   g0861(.dina(new_new_n3185__), .dinb(new_new_n1444__), .dout(new_new_n1840__));
  and1  g0862(.dina(new_new_n3186__), .dinb(new_new_n1057__), .dout(new_new_n1841__));
  or1   g0863(.dina(new_new_n3188__), .dinb(new_new_n1058__), .dout(new_new_n1842__));
  and1  g0864(.dina(new_new_n1464__), .dinb(new_new_n1421__), .dout(new_new_n1843__));
  and1  g0865(.dina(new_new_n1463__), .dinb(new_new_n1422__), .dout(new_new_n1844__));
  or1   g0866(.dina(new_new_n1844__), .dinb(new_new_n1843__), .dout(new_new_n1845__));
  and1  g0867(.dina(new_new_n1404__), .dinb(new_new_n3189__), .dout(new_new_n1846__));
  or1   g0868(.dina(new_new_n3190__), .dinb(new_new_n3191__), .dout(new_new_n1847__));
  and1  g0869(.dina(new_new_n1847__), .dinb(new_new_n1030__), .dout(new_new_n1848__));
  or1   g0870(.dina(new_new_n1846__), .dinb(new_new_n3192__), .dout(new_new_n1849__));
  and1  g0871(.dina(new_new_n3193__), .dinb(new_new_n3195__), .dout(new_new_n1850__));
  or1   g0872(.dina(new_new_n3198__), .dinb(new_new_n3202__), .dout(new_new_n1851__));
  and1  g0873(.dina(new_new_n3204__), .dinb(new_new_n3205__), .dout(new_new_n1852__));
  or1   g0874(.dina(new_new_n3206__), .dinb(new_new_n3207__), .dout(new_new_n1853__));
  and1  g0875(.dina(new_new_n1518__), .dinb(new_new_n1516__), .dout(new_new_n1854__));
  or1   g0876(.dina(new_new_n1517__), .dinb(new_new_n1515__), .dout(new_new_n1855__));
  and1  g0877(.dina(new_new_n1854__), .dinb(new_new_n3211__), .dout(new_new_n1856__));
  or1   g0878(.dina(new_new_n1855__), .dinb(new_new_n3220__), .dout(new_new_n1857__));
  and1  g0879(.dina(new_new_n3228__), .dinb(new_new_n3220__), .dout(new_new_n1858__));
  or1   g0880(.dina(new_new_n1853__), .dinb(new_new_n3211__), .dout(new_new_n1859__));
  and1  g0881(.dina(new_new_n1859__), .dinb(new_new_n1857__), .dout(new_new_n1860__));
  or1   g0882(.dina(new_new_n1858__), .dinb(new_new_n1856__), .dout(new_new_n1861__));
  and1  g0883(.dina(new_new_n1537__), .dinb(new_new_n3230__), .dout(new_new_n1862__));
  or1   g0884(.dina(new_new_n1538__), .dinb(new_new_n3231__), .dout(new_new_n1863__));
  and1  g0885(.dina(new_new_n3221__), .dinb(new_new_n1479__), .dout(new_new_n1864__));
  or1   g0886(.dina(new_new_n3212__), .dinb(new_new_n1480__), .dout(new_new_n1865__));
  and1  g0887(.dina(new_new_n3232__), .dinb(new_new_n3234__), .dout(new_new_n1866__));
  or1   g0888(.dina(new_new_n3235__), .dinb(new_new_n3236__), .dout(new_new_n1867__));
  and1  g0889(.dina(new_new_n3235__), .dinb(new_new_n3236__), .dout(new_new_n1868__));
  or1   g0890(.dina(new_new_n3232__), .dinb(new_new_n3234__), .dout(new_new_n1869__));
  and1  g0891(.dina(new_new_n1869__), .dinb(new_new_n1867__), .dout(new_new_n1870__));
  or1   g0892(.dina(new_new_n1868__), .dinb(new_new_n1866__), .dout(new_new_n1871__));
  and1  g0893(.dina(new_new_n1539__), .dinb(new_new_n3238__), .dout(new_new_n1872__));
  or1   g0894(.dina(new_new_n1540__), .dinb(new_new_n3239__), .dout(new_new_n1873__));
  and1  g0895(.dina(new_new_n3221__), .dinb(new_new_n1485__), .dout(new_new_n1874__));
  or1   g0896(.dina(new_new_n3212__), .dinb(new_new_n1486__), .dout(new_new_n1875__));
  and1  g0897(.dina(new_new_n3240__), .dinb(new_new_n3242__), .dout(new_new_n1876__));
  or1   g0898(.dina(new_new_n3243__), .dinb(new_new_n3244__), .dout(new_new_n1877__));
  and1  g0899(.dina(new_new_n3243__), .dinb(new_new_n3244__), .dout(new_new_n1878__));
  or1   g0900(.dina(new_new_n3240__), .dinb(new_new_n3242__), .dout(new_new_n1879__));
  and1  g0901(.dina(new_new_n1879__), .dinb(new_new_n1877__), .dout(new_new_n1880__));
  or1   g0902(.dina(new_new_n1878__), .dinb(new_new_n1876__), .dout(new_new_n1881__));
  and1  g0903(.dina(new_new_n1225__), .dinb(new_new_n3247__), .dout(new_new_n1882__));
  or1   g0904(.dina(new_new_n1226__), .dinb(new_new_n3250__), .dout(new_new_n1883__));
  and1  g0905(.dina(new_new_n1227__), .dinb(new_new_n3247__), .dout(new_new_n1884__));
  or1   g0906(.dina(new_new_n1228__), .dinb(new_new_n3250__), .dout(new_new_n1885__));
  or1   g0907(.dina(new_new_n3253__), .dinb(new_new_n3256__), .dout(new_new_n1886__));
  or1   g0908(.dina(new_new_n1886__), .dinb(new_new_n3258__), .dout(new_new_n1887__));
  or1   g0909(.dina(new_new_n3253__), .dinb(new_new_n3260__), .dout(new_new_n1888__));
  or1   g0910(.dina(new_new_n1888__), .dinb(new_new_n3258__), .dout(new_new_n1889__));
  and1  g0911(.dina(new_new_n3204__), .dinb(new_new_n1489__), .dout(new_new_n1890__));
  or1   g0912(.dina(new_new_n3206__), .dinb(new_new_n3261__), .dout(new_new_n1891__));
  and1  g0913(.dina(new_new_n1495__), .dinb(new_new_n3262__), .dout(new_new_n1892__));
  or1   g0914(.dina(new_new_n1496__), .dinb(new_new_n1374__), .dout(new_new_n1893__));
  and1  g0915(.dina(new_new_n3263__), .dinb(new_new_n3264__), .dout(new_new_n1894__));
  or1   g0916(.dina(new_new_n1376__), .dinb(new_new_n1296__), .dout(new_new_n1895__));
  and1  g0917(.dina(new_new_n1895__), .dinb(new_new_n1294__), .dout(new_new_n1896__));
  or1   g0918(.dina(new_new_n1894__), .dinb(new_new_n1293__), .dout(new_new_n1897__));
  and1  g0919(.dina(new_new_n1896__), .dinb(new_new_n1893__), .dout(new_new_n1898__));
  or1   g0920(.dina(new_new_n1897__), .dinb(new_new_n1892__), .dout(new_new_n1899__));
  and1  g0921(.dina(new_new_n1898__), .dinb(new_new_n1891__), .dout(new_new_n1900__));
  or1   g0922(.dina(new_new_n1899__), .dinb(new_new_n1890__), .dout(new_new_n1901__));
  and1  g0923(.dina(new_new_n3266__), .dinb(new_new_n3268__), .dout(new_new_n1902__));
  or1   g0924(.dina(new_new_n1871__), .dinb(new_new_n1861__), .dout(new_new_n1903__));
  or1   g0925(.dina(new_new_n3269__), .dinb(new_new_n3271__), .dout(new_new_n1904__));
  and1  g0926(.dina(new_new_n3272__), .dinb(new_new_n3213__), .dout(new_new_n1905__));
  or1   g0927(.dina(new_new_n1900__), .dinb(new_new_n3223__), .dout(new_new_n1906__));
  and1  g0928(.dina(new_new_n3260__), .dinb(new_new_n3246__), .dout(new_new_n1907__));
  or1   g0929(.dina(new_new_n3256__), .dinb(new_new_n3249__), .dout(new_new_n1908__));
  and1  g0930(.dina(new_new_n3273__), .dinb(new_new_n3274__), .dout(new_new_n1909__));
  or1   g0931(.dina(new_new_n3275__), .dinb(new_new_n3259__), .dout(new_new_n1910__));
  and1  g0932(.dina(new_new_n3276__), .dinb(new_new_n3278__), .dout(new_new_n1911__));
  or1   g0933(.dina(new_new_n3280__), .dinb(new_new_n3254__), .dout(new_new_n1912__));
  and1  g0934(.dina(new_new_n3275__), .dinb(new_new_n3274__), .dout(new_new_n1913__));
  or1   g0935(.dina(new_new_n3273__), .dinb(new_new_n3259__), .dout(new_new_n1914__));
  and1  g0936(.dina(new_new_n3281__), .dinb(new_new_n3254__), .dout(new_new_n1915__));
  or1   g0937(.dina(new_new_n3282__), .dinb(new_new_n3278__), .dout(new_new_n1916__));
  and1  g0938(.dina(new_new_n3276__), .dinb(new_new_n3255__), .dout(new_new_n1917__));
  or1   g0939(.dina(new_new_n3280__), .dinb(new_new_n3279__), .dout(new_new_n1918__));
  and1  g0940(.dina(new_new_n3281__), .dinb(new_new_n3279__), .dout(new_new_n1919__));
  or1   g0941(.dina(new_new_n3282__), .dinb(new_new_n3255__), .dout(new_new_n1920__));
  and1  g0942(.dina(new_new_n1448__), .dinb(new_new_n3283__), .dout(new_new_n1921__));
  or1   g0943(.dina(new_new_n1447__), .dinb(new_new_n3284__), .dout(new_new_n1922__));
  and1  g0944(.dina(new_new_n1484__), .dinb(new_new_n1481__), .dout(new_new_n1923__));
  or1   g0945(.dina(new_new_n1483__), .dinb(new_new_n1482__), .dout(new_new_n1924__));
  and1  g0946(.dina(new_new_n3285__), .dinb(new_new_n3287__), .dout(new_new_n1925__));
  or1   g0947(.dina(new_new_n1430__), .dinb(new_new_n3290__), .dout(new_new_n1926__));
  and1  g0948(.dina(new_new_n1925__), .dinb(new_new_n1840__), .dout(new_new_n1927__));
  or1   g0949(.dina(new_new_n1926__), .dinb(new_new_n3292__), .dout(new_new_n1928__));
  and1  g0950(.dina(new_new_n3293__), .dinb(new_new_n3295__), .dout(new_new_n1929__));
  or1   g0951(.dina(new_new_n3296__), .dinb(new_new_n3297__), .dout(new_new_n1930__));
  and1  g0952(.dina(new_new_n3298__), .dinb(new_new_n1921__), .dout(new_new_n1931__));
  and1  g0953(.dina(new_new_n1929__), .dinb(new_new_n3300__), .dout(new_new_n1932__));
  or1   g0954(.dina(new_new_n1932__), .dinb(new_new_n1931__), .dout(new_new_n1933__));
  and1  g0955(.dina(new_new_n1933__), .dinb(new_new_n3202__), .dout(new_new_n1934__));
  or1   g0956(.dina(new_new_n3303__), .dinb(new_new_n1033__), .dout(new_new_n1935__));
  or1   g0957(.dina(new_new_n3308__), .dinb(new_new_n1254__), .dout(new_new_n1936__));
  and1  g0958(.dina(new_new_n1106__), .dinb(new_new_n3310__), .dout(new_new_n1937__));
  or1   g0959(.dina(new_new_n1105__), .dinb(new_new_n1032__), .dout(new_new_n1938__));
  and1  g0960(.dina(new_new_n1938__), .dinb(new_new_n3311__), .dout(new_new_n1939__));
  or1   g0961(.dina(new_new_n1937__), .dinb(new_new_n1064__), .dout(new_new_n1940__));
  or1   g0962(.dina(new_new_n1469__), .dinb(new_new_n1458__), .dout(new_new_n1941__));
  or1   g0963(.dina(new_new_n1492__), .dinb(new_new_n1456__), .dout(new_new_n1942__));
  and1  g0964(.dina(new_new_n1942__), .dinb(new_new_n1941__), .dout(new_new_n1943__));
  or1   g0965(.dina(new_new_n1943__), .dinb(new_new_n3314__), .dout(new_new_n1944__));
  and1  g0966(.dina(new_new_n1944__), .dinb(new_new_n3320__), .dout(new_new_n1945__));
  and1  g0967(.dina(new_new_n1945__), .dinb(new_new_n1936__), .dout(new_new_n1946__));
  and1  g0968(.dina(new_new_n3300__), .dinb(new_new_n3198__), .dout(new_new_n1947__));
  or1   g0969(.dina(new_new_n1947__), .dinb(new_new_n1946__), .dout(new_new_n1948__));
  or1   g0970(.dina(new_new_n1948__), .dinb(new_new_n1934__), .dout(new_new_n1949__));
  and1  g0971(.dina(new_new_n1442__), .dinb(new_new_n1439__), .dout(new_new_n1950__));
  or1   g0972(.dina(new_new_n1441__), .dinb(new_new_n1440__), .dout(new_new_n1951__));
  or1   g0973(.dina(new_new_n3325__), .dinb(new_new_n3308__), .dout(new_new_n1952__));
  or1   g0974(.dina(new_new_n1487__), .dinb(new_new_n1431__), .dout(new_new_n1953__));
  or1   g0975(.dina(new_new_n1467__), .dinb(new_new_n1414__), .dout(new_new_n1954__));
  or1   g0976(.dina(new_new_n1954__), .dinb(new_new_n1953__), .dout(new_new_n1955__));
  or1   g0977(.dina(new_new_n1462__), .dinb(new_new_n1410__), .dout(new_new_n1956__));
  or1   g0978(.dina(new_new_n1466__), .dinb(new_new_n1460__), .dout(new_new_n1957__));
  or1   g0979(.dina(new_new_n1957__), .dinb(new_new_n1956__), .dout(new_new_n1958__));
  and1  g0980(.dina(new_new_n1958__), .dinb(new_new_n1955__), .dout(new_new_n1959__));
  or1   g0981(.dina(new_new_n1959__), .dinb(new_new_n3314__), .dout(new_new_n1960__));
  and1  g0982(.dina(new_new_n1960__), .dinb(new_new_n3320__), .dout(new_new_n1961__));
  and1  g0983(.dina(new_new_n1961__), .dinb(new_new_n1952__), .dout(new_new_n1962__));
  and1  g0984(.dina(new_new_n3325__), .dinb(new_new_n3327__), .dout(new_new_n1963__));
  or1   g0985(.dina(new_new_n3328__), .dinb(new_new_n3329__), .dout(new_new_n1964__));
  and1  g0986(.dina(new_new_n3328__), .dinb(new_new_n3329__), .dout(new_new_n1965__));
  or1   g0987(.dina(new_new_n3324__), .dinb(new_new_n3327__), .dout(new_new_n1966__));
  and1  g0988(.dina(new_new_n1966__), .dinb(new_new_n1964__), .dout(new_new_n1967__));
  or1   g0989(.dina(new_new_n1965__), .dinb(new_new_n1963__), .dout(new_new_n1968__));
  and1  g0990(.dina(new_new_n1968__), .dinb(new_new_n3283__), .dout(new_new_n1969__));
  and1  g0991(.dina(new_new_n1967__), .dinb(new_new_n3284__), .dout(new_new_n1970__));
  or1   g0992(.dina(new_new_n1970__), .dinb(new_new_n1969__), .dout(new_new_n1971__));
  and1  g0993(.dina(new_new_n3295__), .dinb(new_new_n3299__), .dout(new_new_n1972__));
  or1   g0994(.dina(new_new_n1972__), .dinb(new_new_n3293__), .dout(new_new_n1973__));
  and1  g0995(.dina(new_new_n1973__), .dinb(new_new_n3203__), .dout(new_new_n1974__));
  or1   g0996(.dina(new_new_n1974__), .dinb(new_new_n3199__), .dout(new_new_n1975__));
  and1  g0997(.dina(new_new_n1975__), .dinb(new_new_n1971__), .dout(new_new_n1976__));
  or1   g0998(.dina(new_new_n1976__), .dinb(new_new_n1962__), .dout(new_new_n1977__));
  or1   g0999(.dina(new_new_n3332__), .dinb(new_new_n3335__), .dout(new_new_n1978__));
  and1  g1000(.dina(new_new_n3337__), .dinb(new_new_n1259__), .dout(new_new_n1979__));
  or1   g1001(.dina(new_new_n3338__), .dinb(new_new_n3339__), .dout(new_new_n1980__));
  and1  g1002(.dina(new_new_n1532__), .dinb(new_new_n1512__), .dout(new_new_n1981__));
  or1   g1003(.dina(new_new_n1531__), .dinb(new_new_n1511__), .dout(new_new_n1982__));
  and1  g1004(.dina(new_new_n3341__), .dinb(new_new_n1980__), .dout(new_new_n1983__));
  or1   g1005(.dina(new_new_n3343__), .dinb(new_new_n1979__), .dout(new_new_n1984__));
  and1  g1006(.dina(new_new_n3337__), .dinb(new_new_n3344__), .dout(new_new_n1985__));
  or1   g1007(.dina(new_new_n3338__), .dinb(new_new_n3345__), .dout(new_new_n1986__));
  and1  g1008(.dina(new_new_n1985__), .dinb(new_new_n3343__), .dout(new_new_n1987__));
  or1   g1009(.dina(new_new_n1986__), .dinb(new_new_n3341__), .dout(new_new_n1988__));
  and1  g1010(.dina(new_new_n3346__), .dinb(new_new_n1984__), .dout(new_new_n1989__));
  or1   g1011(.dina(new_new_n3347__), .dinb(new_new_n1983__), .dout(new_new_n1990__));
  and1  g1012(.dina(new_new_n3342__), .dinb(new_new_n1477__), .dout(new_new_n1991__));
  or1   g1013(.dina(new_new_n3340__), .dinb(new_new_n3349__), .dout(new_new_n1992__));
  and1  g1014(.dina(new_new_n3350__), .dinb(new_new_n3352__), .dout(new_new_n1993__));
  or1   g1015(.dina(new_new_n3353__), .dinb(new_new_n3354__), .dout(new_new_n1994__));
  and1  g1016(.dina(new_new_n3353__), .dinb(new_new_n3354__), .dout(new_new_n1995__));
  or1   g1017(.dina(new_new_n3350__), .dinb(new_new_n3352__), .dout(new_new_n1996__));
  and1  g1018(.dina(new_new_n1996__), .dinb(new_new_n1994__), .dout(new_new_n1997__));
  or1   g1019(.dina(new_new_n1995__), .dinb(new_new_n1993__), .dout(new_new_n1998__));
  or1   g1020(.dina(new_new_n3335__), .dinb(new_new_n3356__), .dout(new_new_n1999__));
  and1  g1021(.dina(new_new_n3358__), .dinb(new_new_n1564__), .dout(new_new_n2000__));
  or1   g1022(.dina(new_new_n3360__), .dinb(new_new_n3361__), .dout(new_new_n2001__));
  or1   g1023(.dina(new_new_n3362__), .dinb(new_new_n3363__), .dout(new_new_n2002__));
  and1  g1024(.dina(new_new_n3365__), .dinb(new_new_n3366__), .dout(new_new_n2003__));
  or1   g1025(.dina(new_new_n3368__), .dinb(new_new_n3369__), .dout(new_new_n2004__));
  or1   g1026(.dina(new_new_n3370__), .dinb(new_new_n1174__), .dout(new_new_n2005__));
  and1  g1027(.dina(new_new_n3372__), .dinb(new_new_n3374__), .dout(new_new_n2006__));
  or1   g1028(.dina(new_new_n3375__), .dinb(new_new_n3378__), .dout(new_new_n2007__));
  or1   g1029(.dina(new_new_n3381__), .dinb(new_new_n3383__), .dout(new_new_n2008__));
  and1  g1030(.dina(new_new_n3384__), .dinb(new_new_n3266__), .dout(new_new_n2009__));
  or1   g1031(.dina(new_new_n3385__), .dinb(new_new_n3332__), .dout(new_new_n2010__));
  and1  g1032(.dina(new_new_n3386__), .dinb(new_new_n1572__), .dout(new_new_n2011__));
  or1   g1033(.dina(new_new_n1601__), .dinb(new_new_n1571__), .dout(new_new_n2012__));
  and1  g1034(.dina(new_new_n3388__), .dinb(new_new_n3392__), .dout(new_new_n2013__));
  or1   g1035(.dina(new_new_n3395__), .dinb(new_new_n3398__), .dout(new_new_n2014__));
  and1  g1036(.dina(new_new_n3401__), .dinb(new_new_n3398__), .dout(new_new_n2015__));
  or1   g1037(.dina(new_new_n3405__), .dinb(new_new_n3392__), .dout(new_new_n2016__));
  and1  g1038(.dina(new_new_n2016__), .dinb(new_new_n2014__), .dout(new_new_n2017__));
  or1   g1039(.dina(new_new_n2015__), .dinb(new_new_n2013__), .dout(new_new_n2018__));
  and1  g1040(.dina(new_new_n3410__), .dinb(new_new_n3413__), .dout(new_new_n2019__));
  or1   g1041(.dina(new_new_n3331__), .dinb(new_new_n3416__), .dout(new_new_n2020__));
  and1  g1042(.dina(new_new_n1586__), .dinb(new_new_n1578__), .dout(new_new_n2021__));
  or1   g1043(.dina(new_new_n1585__), .dinb(new_new_n1577__), .dout(new_new_n2022__));
  and1  g1044(.dina(new_new_n2021__), .dinb(new_new_n2020__), .dout(new_new_n2023__));
  or1   g1045(.dina(new_new_n2022__), .dinb(new_new_n2019__), .dout(new_new_n2024__));
  and1  g1046(.dina(new_new_n2024__), .dinb(new_new_n3420__), .dout(new_new_n2025__));
  or1   g1047(.dina(new_new_n2023__), .dinb(new_new_n3427__), .dout(new_new_n2026__));
  and1  g1048(.dina(new_new_n2026__), .dinb(new_new_n2018__), .dout(new_new_n2027__));
  or1   g1049(.dina(new_new_n2025__), .dinb(new_new_n2017__), .dout(new_new_n2028__));
  and1  g1050(.dina(new_new_n3388__), .dinb(new_new_n3430__), .dout(new_new_n2029__));
  or1   g1051(.dina(new_new_n3395__), .dinb(new_new_n3433__), .dout(new_new_n2030__));
  and1  g1052(.dina(new_new_n3401__), .dinb(new_new_n3433__), .dout(new_new_n2031__));
  or1   g1053(.dina(new_new_n3405__), .dinb(new_new_n3430__), .dout(new_new_n2032__));
  and1  g1054(.dina(new_new_n2032__), .dinb(new_new_n2030__), .dout(new_new_n2033__));
  or1   g1055(.dina(new_new_n2031__), .dinb(new_new_n2029__), .dout(new_new_n2034__));
  and1  g1056(.dina(new_new_n3437__), .dinb(new_new_n3440__), .dout(new_new_n2035__));
  or1   g1057(.dina(new_new_n3442__), .dinb(new_new_n1575__), .dout(new_new_n2036__));
  and1  g1058(.dina(new_new_n1588__), .dinb(new_new_n1580__), .dout(new_new_n2037__));
  or1   g1059(.dina(new_new_n1587__), .dinb(new_new_n1579__), .dout(new_new_n2038__));
  and1  g1060(.dina(new_new_n2037__), .dinb(new_new_n2036__), .dout(new_new_n2039__));
  or1   g1061(.dina(new_new_n2038__), .dinb(new_new_n2035__), .dout(new_new_n2040__));
  and1  g1062(.dina(new_new_n2040__), .dinb(new_new_n3420__), .dout(new_new_n2041__));
  or1   g1063(.dina(new_new_n2039__), .dinb(new_new_n3427__), .dout(new_new_n2042__));
  and1  g1064(.dina(new_new_n2042__), .dinb(new_new_n2034__), .dout(new_new_n2043__));
  or1   g1065(.dina(new_new_n2041__), .dinb(new_new_n2033__), .dout(new_new_n2044__));
  or1   g1066(.dina(new_new_n3410__), .dinb(new_new_n3444__), .dout(new_new_n2045__));
  and1  g1067(.dina(new_new_n2045__), .dinb(new_new_n3446__), .dout(new_new_n2046__));
  or1   g1068(.dina(new_new_n3447__), .dinb(new_new_n3449__), .dout(new_new_n2047__));
  and1  g1069(.dina(new_new_n1615__), .dinb(new_new_n3453__), .dout(new_new_n2048__));
  or1   g1070(.dina(new_new_n1616__), .dinb(new_new_n3459__), .dout(new_new_n2049__));
  and1  g1071(.dina(new_new_n1498__), .dinb(new_new_n1384__), .dout(new_new_n2050__));
  or1   g1072(.dina(new_new_n3463__), .dinb(new_new_n3464__), .dout(new_new_n2051__));
  and1  g1073(.dina(new_new_n2051__), .dinb(new_new_n1298__), .dout(new_new_n2052__));
  or1   g1074(.dina(new_new_n2050__), .dinb(new_new_n3449__), .dout(new_new_n2053__));
  and1  g1075(.dina(new_new_n3466__), .dinb(new_new_n3468__), .dout(new_new_n2054__));
  or1   g1076(.dina(new_new_n3470__), .dinb(new_new_n3472__), .dout(new_new_n2055__));
  and1  g1077(.dina(new_new_n3419__), .dinb(new_new_n3475__), .dout(new_new_n2056__));
  or1   g1078(.dina(new_new_n3426__), .dinb(new_new_n3477__), .dout(new_new_n2057__));
  and1  g1079(.dina(new_new_n3478__), .dinb(new_new_n3402__), .dout(new_new_n2058__));
  or1   g1080(.dina(new_new_n3480__), .dinb(new_new_n3406__), .dout(new_new_n2059__));
  and1  g1081(.dina(new_new_n3481__), .dinb(new_new_n3483__), .dout(new_new_n2060__));
  or1   g1082(.dina(new_new_n2058__), .dinb(new_new_n3485__), .dout(new_new_n2061__));
  and1  g1083(.dina(new_new_n3413__), .dinb(new_new_n3399__), .dout(new_new_n2062__));
  or1   g1084(.dina(new_new_n3416__), .dinb(new_new_n3391__), .dout(new_new_n2063__));
  and1  g1085(.dina(new_new_n3487__), .dinb(new_new_n3489__), .dout(new_new_n2064__));
  or1   g1086(.dina(new_new_n3491__), .dinb(new_new_n3493__), .dout(new_new_n2065__));
  and1  g1087(.dina(new_new_n2065__), .dinb(new_new_n2063__), .dout(new_new_n2066__));
  or1   g1088(.dina(new_new_n2064__), .dinb(new_new_n2062__), .dout(new_new_n2067__));
  and1  g1089(.dina(new_new_n2067__), .dinb(new_new_n3421__), .dout(new_new_n2068__));
  or1   g1090(.dina(new_new_n2066__), .dinb(new_new_n3428__), .dout(new_new_n2069__));
  and1  g1091(.dina(new_new_n3396__), .dinb(new_new_n3485__), .dout(new_new_n2070__));
  or1   g1092(.dina(new_new_n3389__), .dinb(new_new_n3483__), .dout(new_new_n2071__));
  and1  g1093(.dina(new_new_n2071__), .dinb(new_new_n2069__), .dout(new_new_n2072__));
  or1   g1094(.dina(new_new_n2070__), .dinb(new_new_n2068__), .dout(new_new_n2073__));
  and1  g1095(.dina(new_new_n2072__), .dinb(new_new_n2061__), .dout(new_new_n2074__));
  or1   g1096(.dina(new_new_n2073__), .dinb(new_new_n2060__), .dout(new_new_n2075__));
  and1  g1097(.dina(new_new_n3468__), .dinb(new_new_n1452__), .dout(new_new_n2076__));
  or1   g1098(.dina(new_new_n3472__), .dinb(new_new_n1451__), .dout(new_new_n2077__));
  and1  g1099(.dina(new_new_n1608__), .dinb(new_new_n1596__), .dout(new_new_n2078__));
  or1   g1100(.dina(new_new_n1607__), .dinb(new_new_n1595__), .dout(new_new_n2079__));
  and1  g1101(.dina(new_new_n2079__), .dinb(new_new_n3453__), .dout(new_new_n2080__));
  or1   g1102(.dina(new_new_n2078__), .dinb(new_new_n3459__), .dout(new_new_n2081__));
  and1  g1103(.dina(new_new_n2081__), .dinb(new_new_n2077__), .dout(new_new_n2082__));
  or1   g1104(.dina(new_new_n2080__), .dinb(new_new_n2076__), .dout(new_new_n2083__));
  or1   g1105(.dina(new_new_n3494__), .dinb(new_new_n3496__), .dout(new_new_n2084__));
  or1   g1106(.dina(new_new_n2084__), .dinb(new_new_n2027__), .dout(new_new_n2085__));
  and1  g1107(.dina(new_new_n3467__), .dinb(new_new_n3499__), .dout(new_new_n2086__));
  or1   g1108(.dina(new_new_n3471__), .dinb(new_new_n3501__), .dout(new_new_n2087__));
  and1  g1109(.dina(new_new_n1606__), .dinb(new_new_n1594__), .dout(new_new_n2088__));
  or1   g1110(.dina(new_new_n1605__), .dinb(new_new_n1593__), .dout(new_new_n2089__));
  and1  g1111(.dina(new_new_n2089__), .dinb(new_new_n3454__), .dout(new_new_n2090__));
  or1   g1112(.dina(new_new_n2088__), .dinb(new_new_n3460__), .dout(new_new_n2091__));
  and1  g1113(.dina(new_new_n2091__), .dinb(new_new_n3503__), .dout(new_new_n2092__));
  or1   g1114(.dina(new_new_n2090__), .dinb(new_new_n3505__), .dout(new_new_n2093__));
  or1   g1115(.dina(new_new_n3506__), .dinb(new_new_n3496__), .dout(new_new_n2094__));
  or1   g1116(.dina(new_new_n2094__), .dinb(new_new_n2043__), .dout(new_new_n2095__));
  or1   g1117(.dina(new_new_n3309__), .dinb(new_new_n1194__), .dout(new_new_n2096__));
  or1   g1118(.dina(new_new_n3309__), .dinb(new_new_n3507__), .dout(new_new_n2097__));
  and1  g1119(.dina(new_new_n3508__), .dinb(new_new_n3510__), .dout(new_new_n2098__));
  or1   g1120(.dina(new_new_n3190__), .dinb(new_new_n3303__), .dout(new_new_n2099__));
  or1   g1121(.dina(new_new_n3512__), .dinb(new_new_n3514__), .dout(new_new_n2100__));
  or1   g1122(.dina(new_new_n3375__), .dinb(new_new_n3516__), .dout(new_new_n2101__));
  or1   g1123(.dina(new_new_n3518__), .dinb(new_new_n3378__), .dout(new_new_n2102__));
  and1  g1124(.dina(new_new_n3296__), .dinb(new_new_n3297__), .dout(new_new_n2103__));
  and1  g1125(.dina(new_new_n3514__), .dinb(new_new_n3287__), .dout(new_new_n2104__));
  or1   g1126(.dina(new_new_n3519__), .dinb(new_new_n3290__), .dout(new_new_n2105__));
  and1  g1127(.dina(new_new_n3184__), .dinb(new_new_n1337__), .dout(new_new_n2106__));
  or1   g1128(.dina(new_new_n3183__), .dinb(new_new_n1338__), .dout(new_new_n2107__));
  and1  g1129(.dina(new_new_n2107__), .dinb(new_new_n3520__), .dout(new_new_n2108__));
  or1   g1130(.dina(new_new_n2106__), .dinb(new_new_n3521__), .dout(new_new_n2109__));
  and1  g1131(.dina(new_new_n3522__), .dinb(new_new_n3523__), .dout(new_new_n2110__));
  or1   g1132(.dina(new_new_n3524__), .dinb(new_new_n3526__), .dout(new_new_n2111__));
  and1  g1133(.dina(new_new_n3524__), .dinb(new_new_n3526__), .dout(new_new_n2112__));
  or1   g1134(.dina(new_new_n3522__), .dinb(new_new_n3523__), .dout(new_new_n2113__));
  and1  g1135(.dina(new_new_n2113__), .dinb(new_new_n2111__), .dout(new_new_n2114__));
  or1   g1136(.dina(new_new_n2112__), .dinb(new_new_n2110__), .dout(new_new_n2115__));
  and1  g1137(.dina(new_new_n3527__), .dinb(new_new_n3528__), .dout(new_new_n2116__));
  or1   g1138(.dina(new_new_n3529__), .dinb(new_new_n3530__), .dout(new_new_n2117__));
  and1  g1139(.dina(new_new_n3529__), .dinb(new_new_n3530__), .dout(new_new_n2118__));
  or1   g1140(.dina(new_new_n3527__), .dinb(new_new_n3528__), .dout(new_new_n2119__));
  and1  g1141(.dina(new_new_n2119__), .dinb(new_new_n2117__), .dout(new_new_n2120__));
  or1   g1142(.dina(new_new_n2118__), .dinb(new_new_n2116__), .dout(new_new_n2121__));
  and1  g1143(.dina(new_new_n3520__), .dinb(new_new_n1426__), .dout(new_new_n2122__));
  or1   g1144(.dina(new_new_n3521__), .dinb(new_new_n1425__), .dout(new_new_n2123__));
  and1  g1145(.dina(new_new_n3531__), .dinb(new_new_n3532__), .dout(new_new_n2124__));
  or1   g1146(.dina(new_new_n3533__), .dinb(new_new_n3535__), .dout(new_new_n2125__));
  and1  g1147(.dina(new_new_n3536__), .dinb(new_new_n3538__), .dout(new_new_n2126__));
  or1   g1148(.dina(new_new_n3540__), .dinb(new_new_n3543__), .dout(new_new_n2127__));
  and1  g1149(.dina(new_new_n3540__), .dinb(new_new_n3543__), .dout(new_new_n2128__));
  or1   g1150(.dina(new_new_n3536__), .dinb(new_new_n3538__), .dout(new_new_n2129__));
  and1  g1151(.dina(new_new_n2129__), .dinb(new_new_n2127__), .dout(new_new_n2130__));
  or1   g1152(.dina(new_new_n2128__), .dinb(new_new_n2126__), .dout(new_new_n2131__));
  or1   g1153(.dina(new_new_n3545__), .dinb(new_new_n3546__), .dout(new_new_n2132__));
  and1  g1154(.dina(new_new_n2132__), .dinb(new_new_n3548__), .dout(new_new_n2133__));
  or1   g1155(.dina(new_new_n2133__), .dinb(new_new_n3195__), .dout(new_new_n2134__));
  and1  g1156(.dina(new_new_n2134__), .dinb(new_new_n3193__), .dout(new_new_n2135__));
  and1  g1157(.dina(new_new_n3551__), .dinb(new_new_n3199__), .dout(new_new_n2136__));
  and1  g1158(.dina(new_new_n3552__), .dinb(new_new_n3200__), .dout(new_new_n2137__));
  and1  g1159(.dina(new_new_n3519__), .dinb(new_new_n3291__), .dout(new_new_n2138__));
  or1   g1160(.dina(new_new_n2138__), .dinb(new_new_n3525__), .dout(new_new_n2139__));
  and1  g1161(.dina(new_new_n3186__), .dinb(new_new_n3304__), .dout(new_new_n2140__));
  or1   g1162(.dina(new_new_n3188__), .dinb(new_new_n3555__), .dout(new_new_n2141__));
  or1   g1163(.dina(new_new_n2140__), .dinb(new_new_n3560__), .dout(new_new_n2142__));
  and1  g1164(.dina(new_new_n3562__), .dinb(new_new_n3191__), .dout(new_new_n2143__));
  and1  g1165(.dina(new_new_n3563__), .dinb(new_new_n3189__), .dout(new_new_n2144__));
  or1   g1166(.dina(new_new_n2141__), .dinb(new_new_n3564__), .dout(new_new_n2145__));
  or1   g1167(.dina(new_new_n2145__), .dinb(new_new_n2144__), .dout(new_new_n2146__));
  or1   g1168(.dina(new_new_n2146__), .dinb(new_new_n2143__), .dout(new_new_n2147__));
  and1  g1169(.dina(new_new_n2147__), .dinb(new_new_n2142__), .dout(new_new_n2148__));
  or1   g1170(.dina(new_new_n2148__), .dinb(new_new_n3565__), .dout(new_new_n2149__));
  or1   g1171(.dina(new_new_n3568__), .dinb(new_new_n988__), .dout(new_new_n2150__));
  or1   g1172(.dina(new_new_n1400__), .dinb(new_new_n3571__), .dout(new_new_n2151__));
  or1   g1173(.dina(new_new_n1304__), .dinb(new_new_n3574__), .dout(new_new_n2152__));
  and1  g1174(.dina(new_new_n2152__), .dinb(new_new_n2151__), .dout(new_new_n2153__));
  and1  g1175(.dina(new_new_n2153__), .dinb(new_new_n2150__), .dout(new_new_n2154__));
  or1   g1176(.dina(new_new_n3574__), .dinb(new_new_n1052__), .dout(new_new_n2155__));
  or1   g1177(.dina(new_new_n1302__), .dinb(new_new_n3568__), .dout(new_new_n2156__));
  and1  g1178(.dina(new_new_n2156__), .dinb(new_new_n2155__), .dout(new_new_n2157__));
  or1   g1179(.dina(new_new_n3577__), .dinb(new_new_n3578__), .dout(new_new_n2158__));
  and1  g1180(.dina(new_new_n2158__), .dinb(new_new_n3555__), .dout(new_new_n2159__));
  or1   g1181(.dina(new_new_n1402__), .dinb(new_new_n3580__), .dout(new_new_n2160__));
  or1   g1182(.dina(new_new_n3583__), .dinb(new_new_n3584__), .dout(new_new_n2161__));
  and1  g1183(.dina(new_new_n2161__), .dinb(new_new_n2160__), .dout(new_new_n2162__));
  and1  g1184(.dina(new_new_n2162__), .dinb(new_new_n2159__), .dout(new_new_n2163__));
  and1  g1185(.dina(new_new_n2163__), .dinb(new_new_n3585__), .dout(new_new_n2164__));
  and1  g1186(.dina(new_new_n2164__), .dinb(new_new_n2154__), .dout(new_new_n2165__));
  or1   g1187(.dina(new_new_n3571__), .dinb(new_new_n3587__), .dout(new_new_n2166__));
  and1  g1188(.dina(new_new_n2166__), .dinb(new_new_n1267__), .dout(new_new_n2167__));
  or1   g1189(.dina(new_new_n3583__), .dinb(new_new_n3588__), .dout(new_new_n2168__));
  and1  g1190(.dina(new_new_n3589__), .dinb(new_new_n1263__), .dout(new_new_n2169__));
  and1  g1191(.dina(new_new_n2169__), .dinb(new_new_n2167__), .dout(new_new_n2170__));
  or1   g1192(.dina(new_new_n1417__), .dinb(new_new_n3567__), .dout(new_new_n2171__));
  and1  g1193(.dina(new_new_n2171__), .dinb(new_new_n3304__), .dout(new_new_n2172__));
  or1   g1194(.dina(new_new_n3580__), .dinb(new_new_n3179__), .dout(new_new_n2173__));
  and1  g1195(.dina(new_new_n2173__), .dinb(new_new_n1261__), .dout(new_new_n2174__));
  and1  g1196(.dina(new_new_n2174__), .dinb(new_new_n2172__), .dout(new_new_n2175__));
  and1  g1197(.dina(new_new_n2175__), .dinb(new_new_n2170__), .dout(new_new_n2176__));
  or1   g1198(.dina(new_new_n2176__), .dinb(new_new_n3315__), .dout(new_new_n2177__));
  or1   g1199(.dina(new_new_n2177__), .dinb(new_new_n2165__), .dout(new_new_n2178__));
  and1  g1200(.dina(new_new_n2178__), .dinb(new_new_n2149__), .dout(new_new_n2179__));
  or1   g1201(.dina(new_new_n2179__), .dinb(new_new_n3590__), .dout(new_new_n2180__));
  or1   g1202(.dina(new_new_n3569__), .dinb(new_new_n3591__), .dout(new_new_n2181__));
  or1   g1203(.dina(new_new_n3575__), .dinb(new_new_n3592__), .dout(new_new_n2182__));
  or1   g1204(.dina(new_new_n3581__), .dinb(new_new_n3578__), .dout(new_new_n2183__));
  and1  g1205(.dina(new_new_n2183__), .dinb(new_new_n2182__), .dout(new_new_n2184__));
  and1  g1206(.dina(new_new_n2184__), .dinb(new_new_n2181__), .dout(new_new_n2185__));
  and1  g1207(.dina(new_new_n3589__), .dinb(new_new_n3556__), .dout(new_new_n2186__));
  or1   g1208(.dina(new_new_n3577__), .dinb(new_new_n3593__), .dout(new_new_n2187__));
  or1   g1209(.dina(new_new_n3572__), .dinb(new_new_n3584__), .dout(new_new_n2188__));
  and1  g1210(.dina(new_new_n2188__), .dinb(new_new_n2187__), .dout(new_new_n2189__));
  and1  g1211(.dina(new_new_n2189__), .dinb(new_new_n2186__), .dout(new_new_n2190__));
  and1  g1212(.dina(new_new_n2190__), .dinb(new_new_n3585__), .dout(new_new_n2191__));
  and1  g1213(.dina(new_new_n2191__), .dinb(new_new_n2185__), .dout(new_new_n2192__));
  or1   g1214(.dina(new_new_n3582__), .dinb(new_new_n3587__), .dout(new_new_n2193__));
  or1   g1215(.dina(new_new_n3581__), .dinb(new_new_n1202__), .dout(new_new_n2194__));
  or1   g1216(.dina(new_new_n3572__), .dinb(new_new_n1204__), .dout(new_new_n2195__));
  and1  g1217(.dina(new_new_n2195__), .dinb(new_new_n2194__), .dout(new_new_n2196__));
  and1  g1218(.dina(new_new_n2196__), .dinb(new_new_n2193__), .dout(new_new_n2197__));
  or1   g1219(.dina(new_new_n1272__), .dinb(new_new_n3569__), .dout(new_new_n2198__));
  and1  g1220(.dina(new_new_n2198__), .dinb(new_new_n3306__), .dout(new_new_n2199__));
  or1   g1221(.dina(new_new_n3576__), .dinb(new_new_n3180__), .dout(new_new_n2200__));
  or1   g1222(.dina(new_new_n1415__), .dinb(new_new_n3575__), .dout(new_new_n2201__));
  and1  g1223(.dina(new_new_n2201__), .dinb(new_new_n2200__), .dout(new_new_n2202__));
  and1  g1224(.dina(new_new_n2202__), .dinb(new_new_n2199__), .dout(new_new_n2203__));
  and1  g1225(.dina(new_new_n2203__), .dinb(new_new_n2197__), .dout(new_new_n2204__));
  or1   g1226(.dina(new_new_n2204__), .dinb(new_new_n2192__), .dout(new_new_n2205__));
  and1  g1227(.dina(new_new_n2205__), .dinb(new_new_n3565__), .dout(new_new_n2206__));
  or1   g1228(.dina(new_new_n2206__), .dinb(new_new_n3590__), .dout(new_new_n2207__));
  and1  g1229(.dina(new_new_n3596__), .dinb(new_new_n3598__), .dout(new_new_n2208__));
  and1  g1230(.dina(new_new_n1301__), .dinb(new_new_n3601__), .dout(new_new_n2209__));
  or1   g1231(.dina(new_new_n3605__), .dinb(new_new_n3607__), .dout(new_new_n2210__));
  and1  g1232(.dina(new_new_n2210__), .dinb(new_new_n3612__), .dout(new_new_n2211__));
  or1   g1233(.dina(new_new_n2211__), .dinb(new_new_n2209__), .dout(new_new_n2212__));
  or1   g1234(.dina(new_new_n2212__), .dinb(new_new_n2208__), .dout(new_new_n2213__));
  or1   g1235(.dina(new_new_n3618__), .dinb(new_new_n3619__), .dout(new_new_n2214__));
  and1  g1236(.dina(new_new_n2214__), .dinb(new_new_n3622__), .dout(new_new_n2215__));
  or1   g1237(.dina(new_new_n2215__), .dinb(new_new_n3306__), .dout(new_new_n2216__));
  and1  g1238(.dina(new_new_n3627__), .dinb(new_new_n3560__), .dout(new_new_n2217__));
  and1  g1239(.dina(new_new_n3633__), .dinb(new_new_n3637__), .dout(new_new_n2218__));
  or1   g1240(.dina(new_new_n2218__), .dinb(new_new_n2217__), .dout(new_new_n2219__));
  or1   g1241(.dina(new_new_n2219__), .dinb(new_new_n2216__), .dout(new_new_n2220__));
  or1   g1242(.dina(new_new_n2220__), .dinb(new_new_n2213__), .dout(new_new_n2221__));
  and1  g1243(.dina(new_new_n3633__), .dinb(new_new_n3639__), .dout(new_new_n2222__));
  and1  g1244(.dina(new_new_n3601__), .dinb(new_new_n1203__), .dout(new_new_n2223__));
  and1  g1245(.dina(new_new_n1418__), .dinb(new_new_n3622__), .dout(new_new_n2224__));
  or1   g1246(.dina(new_new_n2224__), .dinb(new_new_n2223__), .dout(new_new_n2225__));
  or1   g1247(.dina(new_new_n2225__), .dinb(new_new_n2222__), .dout(new_new_n2226__));
  and1  g1248(.dina(new_new_n3612__), .dinb(new_new_n1236__), .dout(new_new_n2227__));
  or1   g1249(.dina(new_new_n2227__), .dinb(new_new_n3556__), .dout(new_new_n2228__));
  and1  g1250(.dina(new_new_n3627__), .dinb(new_new_n1104__), .dout(new_new_n2229__));
  or1   g1251(.dina(new_new_n2229__), .dinb(new_new_n1313__), .dout(new_new_n2230__));
  or1   g1252(.dina(new_new_n2230__), .dinb(new_new_n2228__), .dout(new_new_n2231__));
  or1   g1253(.dina(new_new_n2231__), .dinb(new_new_n2226__), .dout(new_new_n2232__));
  and1  g1254(.dina(new_new_n2232__), .dinb(new_new_n2221__), .dout(new_new_n2233__));
  or1   g1255(.dina(new_new_n2233__), .dinb(new_new_n3315__), .dout(new_new_n2234__));
  and1  g1256(.dina(new_new_n2234__), .dinb(new_new_n3321__), .dout(new_new_n2235__));
  and1  g1257(.dina(new_new_n3611__), .dinb(new_new_n3598__), .dout(new_new_n2236__));
  and1  g1258(.dina(new_new_n3634__), .dinb(new_new_n3607__), .dout(new_new_n2237__));
  or1   g1259(.dina(new_new_n2237__), .dinb(new_new_n2236__), .dout(new_new_n2238__));
  and1  g1260(.dina(new_new_n3602__), .dinb(new_new_n3618__), .dout(new_new_n2239__));
  or1   g1261(.dina(new_new_n1084__), .dinb(new_new_n3561__), .dout(new_new_n2240__));
  and1  g1262(.dina(new_new_n2240__), .dinb(new_new_n3623__), .dout(new_new_n2241__));
  or1   g1263(.dina(new_new_n2241__), .dinb(new_new_n2239__), .dout(new_new_n2242__));
  or1   g1264(.dina(new_new_n2242__), .dinb(new_new_n2238__), .dout(new_new_n2243__));
  and1  g1265(.dina(new_new_n3613__), .dinb(new_new_n3637__), .dout(new_new_n2244__));
  or1   g1266(.dina(new_new_n2244__), .dinb(new_new_n3305__), .dout(new_new_n2245__));
  and1  g1267(.dina(new_new_n3596__), .dinb(new_new_n3181__), .dout(new_new_n2246__));
  and1  g1268(.dina(new_new_n3628__), .dinb(new_new_n3619__), .dout(new_new_n2247__));
  or1   g1269(.dina(new_new_n2247__), .dinb(new_new_n3640__), .dout(new_new_n2248__));
  or1   g1270(.dina(new_new_n2248__), .dinb(new_new_n3641__), .dout(new_new_n2249__));
  or1   g1271(.dina(new_new_n2249__), .dinb(new_new_n2243__), .dout(new_new_n2250__));
  or1   g1272(.dina(new_new_n1231__), .dinb(new_new_n3639__), .dout(new_new_n2251__));
  and1  g1273(.dina(new_new_n2251__), .dinb(new_new_n3613__), .dout(new_new_n2252__));
  and1  g1274(.dina(new_new_n3628__), .dinb(new_new_n3643__), .dout(new_new_n2253__));
  and1  g1275(.dina(new_new_n3644__), .dinb(new_new_n3623__), .dout(new_new_n2254__));
  or1   g1276(.dina(new_new_n2254__), .dinb(new_new_n2253__), .dout(new_new_n2255__));
  or1   g1277(.dina(new_new_n2255__), .dinb(new_new_n2252__), .dout(new_new_n2256__));
  and1  g1278(.dina(new_new_n3595__), .dinb(new_new_n3645__), .dout(new_new_n2257__));
  and1  g1279(.dina(new_new_n3634__), .dinb(new_new_n1201__), .dout(new_new_n2258__));
  or1   g1280(.dina(new_new_n2258__), .dinb(new_new_n2257__), .dout(new_new_n2259__));
  and1  g1281(.dina(new_new_n1233__), .dinb(new_new_n3602__), .dout(new_new_n2260__));
  or1   g1282(.dina(new_new_n2260__), .dinb(new_new_n3558__), .dout(new_new_n2261__));
  or1   g1283(.dina(new_new_n2261__), .dinb(new_new_n2259__), .dout(new_new_n2262__));
  or1   g1284(.dina(new_new_n2262__), .dinb(new_new_n2256__), .dout(new_new_n2263__));
  and1  g1285(.dina(new_new_n2263__), .dinb(new_new_n2250__), .dout(new_new_n2264__));
  or1   g1286(.dina(new_new_n2264__), .dinb(new_new_n3317__), .dout(new_new_n2265__));
  and1  g1287(.dina(new_new_n2265__), .dinb(new_new_n3321__), .dout(new_new_n2266__));
  and1  g1288(.dina(new_new_n3646__), .dinb(new_new_n1115__), .dout(new_new_n2267__));
  or1   g1289(.dina(new_new_n3647__), .dinb(new_new_n1116__), .dout(new_new_n2268__));
  and1  g1290(.dina(new_new_n3648__), .dinb(new_new_n3649__), .dout(new_new_n2269__));
  or1   g1291(.dina(new_new_n3650__), .dinb(new_new_n3651__), .dout(new_new_n2270__));
  and1  g1292(.dina(new_new_n3650__), .dinb(new_new_n3651__), .dout(new_new_n2271__));
  or1   g1293(.dina(new_new_n3648__), .dinb(new_new_n3649__), .dout(new_new_n2272__));
  and1  g1294(.dina(new_new_n2272__), .dinb(new_new_n2270__), .dout(new_new_n2273__));
  or1   g1295(.dina(new_new_n2271__), .dinb(new_new_n2269__), .dout(new_new_n2274__));
  or1   g1296(.dina(new_new_n3653__), .dinb(new_new_n3512__), .dout(new_new_n2275__));
  or1   g1297(.dina(new_new_n3223__), .dinb(new_new_n3261__), .dout(new_new_n2276__));
  or1   g1298(.dina(new_new_n3654__), .dinb(new_new_n3475__), .dout(new_new_n2277__));
  and1  g1299(.dina(new_new_n1530__), .dinb(new_new_n1510__), .dout(new_new_n2278__));
  or1   g1300(.dina(new_new_n1529__), .dinb(new_new_n1509__), .dout(new_new_n2279__));
  and1  g1301(.dina(new_new_n1514__), .dinb(new_new_n1286__), .dout(new_new_n2280__));
  or1   g1302(.dina(new_new_n1513__), .dinb(new_new_n1285__), .dout(new_new_n2281__));
  or1   g1303(.dina(new_new_n3655__), .dinb(new_new_n3339__), .dout(new_new_n2282__));
  and1  g1304(.dina(new_new_n2282__), .dinb(new_new_n3657__), .dout(new_new_n2283__));
  and1  g1305(.dina(new_new_n2279__), .dinb(new_new_n3344__), .dout(new_new_n2284__));
  or1   g1306(.dina(new_new_n3657__), .dinb(new_new_n3345__), .dout(new_new_n2285__));
  and1  g1307(.dina(new_new_n2284__), .dinb(new_new_n2280__), .dout(new_new_n2286__));
  or1   g1308(.dina(new_new_n2285__), .dinb(new_new_n3655__), .dout(new_new_n2287__));
  or1   g1309(.dina(new_new_n2286__), .dinb(new_new_n2283__), .dout(new_new_n2288__));
  or1   g1310(.dina(new_new_n3659__), .dinb(new_new_n3351__), .dout(new_new_n2289__));
  or1   g1311(.dina(new_new_n3661__), .dinb(new_new_n3241__), .dout(new_new_n2290__));
  or1   g1312(.dina(new_new_n3662__), .dinb(new_new_n3233__), .dout(new_new_n2291__));
  or1   g1313(.dina(new_new_n3551__), .dinb(new_new_n3664__), .dout(new_new_n2292__));
  and1  g1314(.dina(new_new_n3550__), .dinb(new_new_n3664__), .dout(new_new_n2293__));
  or1   g1315(.dina(new_new_n3546__), .dinb(new_new_n3548__), .dout(new_new_n2294__));
  and1  g1316(.dina(new_new_n3665__), .dinb(new_new_n2292__), .dout(new_new_n2295__));
  or1   g1317(.dina(new_new_n3666__), .dinb(new_new_n3668__), .dout(new_new_n2296__));
  or1   g1318(.dina(new_new_n3513__), .dinb(new_new_n3182__), .dout(new_new_n2297__));
  and1  g1319(.dina(new_new_n3669__), .dinb(new_new_n3604__), .dout(new_new_n2298__));
  and1  g1320(.dina(new_new_n3597__), .dinb(new_new_n3608__), .dout(new_new_n2299__));
  or1   g1321(.dina(new_new_n2299__), .dinb(new_new_n2298__), .dout(new_new_n2300__));
  and1  g1322(.dina(new_new_n1408__), .dinb(new_new_n3624__), .dout(new_new_n2301__));
  and1  g1323(.dina(new_new_n3605__), .dinb(new_new_n3636__), .dout(new_new_n2302__));
  or1   g1324(.dina(new_new_n2302__), .dinb(new_new_n2301__), .dout(new_new_n2303__));
  or1   g1325(.dina(new_new_n2303__), .dinb(new_new_n2300__), .dout(new_new_n2304__));
  and1  g1326(.dina(new_new_n3630__), .dinb(new_new_n3617__), .dout(new_new_n2305__));
  and1  g1327(.dina(new_new_n1401__), .dinb(new_new_n3615__), .dout(new_new_n2306__));
  or1   g1328(.dina(new_new_n2306__), .dinb(new_new_n2305__), .dout(new_new_n2307__));
  or1   g1329(.dina(new_new_n2307__), .dinb(new_new_n3641__), .dout(new_new_n2308__));
  or1   g1330(.dina(new_new_n2308__), .dinb(new_new_n2304__), .dout(new_new_n2309__));
  and1  g1331(.dina(new_new_n3604__), .dinb(new_new_n3643__), .dout(new_new_n2310__));
  and1  g1332(.dina(new_new_n1416__), .dinb(new_new_n3615__), .dout(new_new_n2311__));
  or1   g1333(.dina(new_new_n2311__), .dinb(new_new_n2310__), .dout(new_new_n2312__));
  or1   g1334(.dina(new_new_n2312__), .dinb(new_new_n1316__), .dout(new_new_n2313__));
  and1  g1335(.dina(new_new_n3636__), .dinb(new_new_n3645__), .dout(new_new_n2314__));
  or1   g1336(.dina(new_new_n2314__), .dinb(new_new_n3640__), .dout(new_new_n2315__));
  or1   g1337(.dina(new_new_n1356__), .dinb(new_new_n3558__), .dout(new_new_n2316__));
  or1   g1338(.dina(new_new_n2316__), .dinb(new_new_n2315__), .dout(new_new_n2317__));
  or1   g1339(.dina(new_new_n2317__), .dinb(new_new_n2313__), .dout(new_new_n2318__));
  and1  g1340(.dina(new_new_n2318__), .dinb(new_new_n2309__), .dout(new_new_n2319__));
  or1   g1341(.dina(new_new_n2319__), .dinb(new_new_n3317__), .dout(new_new_n2320__));
  and1  g1342(.dina(new_new_n2320__), .dinb(new_new_n3323__), .dout(new_new_n2321__));
  and1  g1343(.dina(new_new_n2321__), .dinb(new_new_n2297__), .dout(new_new_n2322__));
  and1  g1344(.dina(new_new_n3294__), .dinb(new_new_n3200__), .dout(new_new_n2323__));
  and1  g1345(.dina(new_new_n3298__), .dinb(new_new_n3203__), .dout(new_new_n2324__));
  or1   g1346(.dina(new_new_n2324__), .dinb(new_new_n2323__), .dout(new_new_n2325__));
  or1   g1347(.dina(new_new_n3542__), .dinb(new_new_n3513__), .dout(new_new_n2326__));
  and1  g1348(.dina(new_new_n3630__), .dinb(new_new_n1082__), .dout(new_new_n2327__));
  and1  g1349(.dina(new_new_n3603__), .dinb(new_new_n3638__), .dout(new_new_n2328__));
  and1  g1350(.dina(new_new_n3635__), .dinb(new_new_n3642__), .dout(new_new_n2329__));
  or1   g1351(.dina(new_new_n2329__), .dinb(new_new_n2328__), .dout(new_new_n2330__));
  or1   g1352(.dina(new_new_n2330__), .dinb(new_new_n2327__), .dout(new_new_n2331__));
  and1  g1353(.dina(new_new_n3644__), .dinb(new_new_n3616__), .dout(new_new_n2332__));
  or1   g1354(.dina(new_new_n2332__), .dinb(new_new_n3557__), .dout(new_new_n2333__));
  and1  g1355(.dina(new_new_n1406__), .dinb(new_new_n3624__), .dout(new_new_n2334__));
  or1   g1356(.dina(new_new_n2334__), .dinb(new_new_n1269__), .dout(new_new_n2335__));
  or1   g1357(.dina(new_new_n2335__), .dinb(new_new_n2333__), .dout(new_new_n2336__));
  or1   g1358(.dina(new_new_n2336__), .dinb(new_new_n2331__), .dout(new_new_n2337__));
  and1  g1359(.dina(new_new_n3629__), .dinb(new_new_n3608__), .dout(new_new_n2338__));
  and1  g1360(.dina(new_new_n3669__), .dinb(new_new_n3616__), .dout(new_new_n2339__));
  and1  g1361(.dina(new_new_n3597__), .dinb(new_new_n3561__), .dout(new_new_n2340__));
  or1   g1362(.dina(new_new_n2340__), .dinb(new_new_n2339__), .dout(new_new_n2341__));
  or1   g1363(.dina(new_new_n2341__), .dinb(new_new_n2338__), .dout(new_new_n2342__));
  or1   g1364(.dina(new_new_n1435__), .dinb(new_new_n1265__), .dout(new_new_n2343__));
  or1   g1365(.dina(new_new_n1437__), .dinb(new_new_n1411__), .dout(new_new_n2344__));
  or1   g1366(.dina(new_new_n2344__), .dinb(new_new_n2343__), .dout(new_new_n2345__));
  or1   g1367(.dina(new_new_n2345__), .dinb(new_new_n1310__), .dout(new_new_n2346__));
  or1   g1368(.dina(new_new_n2346__), .dinb(new_new_n2342__), .dout(new_new_n2347__));
  and1  g1369(.dina(new_new_n2347__), .dinb(new_new_n2337__), .dout(new_new_n2348__));
  or1   g1370(.dina(new_new_n2348__), .dinb(new_new_n3316__), .dout(new_new_n2349__));
  and1  g1371(.dina(new_new_n2349__), .dinb(new_new_n3323__), .dout(new_new_n2350__));
  and1  g1372(.dina(new_new_n2350__), .dinb(new_new_n2326__), .dout(new_new_n2351__));
  and1  g1373(.dina(new_new_n3665__), .dinb(new_new_n3545__), .dout(new_new_n2352__));
  and1  g1374(.dina(new_new_n2293__), .dinb(new_new_n3552__), .dout(new_new_n2353__));
  or1   g1375(.dina(new_new_n2353__), .dinb(new_new_n2352__), .dout(new_new_n2354__));
  and1  g1376(.dina(new_new_n3671__), .dinb(new_new_n3672__), .dout(new_new_n2355__));
  or1   g1377(.dina(new_new_n2355__), .dinb(new_new_n3368__), .dout(new_new_n2356__));
  and1  g1378(.dina(new_new_n3288__), .dinb(new_new_n1190__), .dout(new_new_n2357__));
  or1   g1379(.dina(new_new_n3291__), .dinb(new_new_n1189__), .dout(new_new_n2358__));
  and1  g1380(.dina(new_new_n3549__), .dinb(new_new_n3507__), .dout(new_new_n2359__));
  or1   g1381(.dina(new_new_n3663__), .dinb(new_new_n1191__), .dout(new_new_n2360__));
  and1  g1382(.dina(new_new_n2360__), .dinb(new_new_n1274__), .dout(new_new_n2361__));
  or1   g1383(.dina(new_new_n2359__), .dinb(new_new_n1273__), .dout(new_new_n2362__));
  and1  g1384(.dina(new_new_n2361__), .dinb(new_new_n2357__), .dout(new_new_n2363__));
  and1  g1385(.dina(new_new_n2362__), .dinb(new_new_n2358__), .dout(new_new_n2364__));
  or1   g1386(.dina(new_new_n2364__), .dinb(new_new_n2363__), .dout(new_new_n2365__));
  and1  g1387(.dina(new_new_n3544__), .dinb(new_new_n3535__), .dout(new_new_n2366__));
  or1   g1388(.dina(new_new_n3539__), .dinb(new_new_n3532__), .dout(new_new_n2367__));
  and1  g1389(.dina(new_new_n3647__), .dinb(new_new_n1127__), .dout(new_new_n2368__));
  or1   g1390(.dina(new_new_n3646__), .dinb(new_new_n1128__), .dout(new_new_n2369__));
  and1  g1391(.dina(new_new_n3531__), .dinb(new_new_n3544__), .dout(new_new_n2370__));
  or1   g1392(.dina(new_new_n3533__), .dinb(new_new_n3539__), .dout(new_new_n2371__));
  and1  g1393(.dina(new_new_n2371__), .dinb(new_new_n2369__), .dout(new_new_n2372__));
  or1   g1394(.dina(new_new_n2370__), .dinb(new_new_n2368__), .dout(new_new_n2373__));
  and1  g1395(.dina(new_new_n3673__), .dinb(new_new_n3653__), .dout(new_new_n2374__));
  or1   g1396(.dina(new_new_n3674__), .dinb(new_new_n3675__), .dout(new_new_n2375__));
  and1  g1397(.dina(new_new_n3674__), .dinb(new_new_n3675__), .dout(new_new_n2376__));
  or1   g1398(.dina(new_new_n3673__), .dinb(new_new_n3652__), .dout(new_new_n2377__));
  and1  g1399(.dina(new_new_n2377__), .dinb(new_new_n2375__), .dout(new_new_n2378__));
  or1   g1400(.dina(new_new_n2376__), .dinb(new_new_n2374__), .dout(new_new_n2379__));
  and1  g1401(.dina(new_new_n2379__), .dinb(new_new_n2367__), .dout(new_new_n2380__));
  and1  g1402(.dina(new_new_n2378__), .dinb(new_new_n2366__), .dout(new_new_n2381__));
  or1   g1403(.dina(new_new_n2381__), .dinb(new_new_n2380__), .dout(new_new_n2382__));
  or1   g1404(.dina(new_new_n3677__), .dinb(new_new_n3679__), .dout(new_new_n2383__));
  and1  g1405(.dina(new_new_n3677__), .dinb(new_new_n3679__), .dout(new_new_n2384__));
  and1  g1406(.dina(new_new_n3224__), .dinb(new_new_n1291__), .dout(new_new_n2385__));
  or1   g1407(.dina(new_new_n3213__), .dinb(new_new_n1292__), .dout(new_new_n2386__));
  and1  g1408(.dina(new_new_n2386__), .dinb(new_new_n1494__), .dout(new_new_n2387__));
  and1  g1409(.dina(new_new_n2385__), .dinb(new_new_n1493__), .dout(new_new_n2388__));
  or1   g1410(.dina(new_new_n2388__), .dinb(new_new_n2387__), .dout(new_new_n2389__));
  and1  g1411(.dina(new_new_n3224__), .dinb(new_new_n1371__), .dout(new_new_n2390__));
  or1   g1412(.dina(new_new_n3215__), .dinb(new_new_n1372__), .dout(new_new_n2391__));
  and1  g1413(.dina(new_new_n2391__), .dinb(new_new_n3207__), .dout(new_new_n2392__));
  and1  g1414(.dina(new_new_n2390__), .dinb(new_new_n3205__), .dout(new_new_n2393__));
  or1   g1415(.dina(new_new_n2393__), .dinb(new_new_n2392__), .dout(new_new_n2394__));
  and1  g1416(.dina(new_new_n3414__), .dinb(new_new_n3434__), .dout(new_new_n2395__));
  or1   g1417(.dina(new_new_n3415__), .dinb(new_new_n3431__), .dout(new_new_n2396__));
  and1  g1418(.dina(new_new_n3487__), .dinb(new_new_n3680__), .dout(new_new_n2397__));
  or1   g1419(.dina(new_new_n3491__), .dinb(new_new_n1398__), .dout(new_new_n2398__));
  and1  g1420(.dina(new_new_n2398__), .dinb(new_new_n2396__), .dout(new_new_n2399__));
  or1   g1421(.dina(new_new_n2397__), .dinb(new_new_n2395__), .dout(new_new_n2400__));
  and1  g1422(.dina(new_new_n2400__), .dinb(new_new_n3421__), .dout(new_new_n2401__));
  or1   g1423(.dina(new_new_n2399__), .dinb(new_new_n3428__), .dout(new_new_n2402__));
  and1  g1424(.dina(new_new_n3402__), .dinb(new_new_n3493__), .dout(new_new_n2403__));
  or1   g1425(.dina(new_new_n3406__), .dinb(new_new_n3489__), .dout(new_new_n2404__));
  and1  g1426(.dina(new_new_n3478__), .dinb(new_new_n3490__), .dout(new_new_n2405__));
  or1   g1427(.dina(new_new_n3480__), .dinb(new_new_n3492__), .dout(new_new_n2406__));
  and1  g1428(.dina(new_new_n2405__), .dinb(new_new_n3389__), .dout(new_new_n2407__));
  or1   g1429(.dina(new_new_n2406__), .dinb(new_new_n3396__), .dout(new_new_n2408__));
  and1  g1430(.dina(new_new_n2408__), .dinb(new_new_n2404__), .dout(new_new_n2409__));
  or1   g1431(.dina(new_new_n2407__), .dinb(new_new_n2403__), .dout(new_new_n2410__));
  and1  g1432(.dina(new_new_n2410__), .dinb(new_new_n2402__), .dout(new_new_n2411__));
  or1   g1433(.dina(new_new_n2409__), .dinb(new_new_n2401__), .dout(new_new_n2412__));
  and1  g1434(.dina(new_new_n3681__), .dinb(new_new_n3501__), .dout(new_new_n2413__));
  or1   g1435(.dina(new_new_n1548__), .dinb(new_new_n3499__), .dout(new_new_n2414__));
  and1  g1436(.dina(new_new_n1604__), .dinb(new_new_n1590__), .dout(new_new_n2415__));
  or1   g1437(.dina(new_new_n1603__), .dinb(new_new_n1589__), .dout(new_new_n2416__));
  and1  g1438(.dina(new_new_n2415__), .dinb(new_new_n2414__), .dout(new_new_n2417__));
  or1   g1439(.dina(new_new_n2416__), .dinb(new_new_n2413__), .dout(new_new_n2418__));
  and1  g1440(.dina(new_new_n2418__), .dinb(new_new_n3454__), .dout(new_new_n2419__));
  or1   g1441(.dina(new_new_n2417__), .dinb(new_new_n3460__), .dout(new_new_n2420__));
  and1  g1442(.dina(new_new_n2420__), .dinb(new_new_n3503__), .dout(new_new_n2421__));
  or1   g1443(.dina(new_new_n2419__), .dinb(new_new_n3505__), .dout(new_new_n2422__));
  or1   g1444(.dina(new_new_n3682__), .dinb(new_new_n3497__), .dout(new_new_n2423__));
  or1   g1445(.dina(new_new_n2423__), .dinb(new_new_n2074__), .dout(new_new_n2424__));
  and1  g1446(.dina(new_new_n3683__), .dinb(new_new_n3686__), .dout(new_new_n2425__));
  or1   g1447(.dina(new_new_n2425__), .dinb(new_new_n3690__), .dout(new_new_n2426__));
  and1  g1448(.dina(new_new_n2426__), .dinb(new_new_n3691__), .dout(new_new_n2427__));
  and1  g1449(.dina(new_new_n3692__), .dinb(new_new_n3686__), .dout(new_new_n2428__));
  or1   g1450(.dina(new_new_n2428__), .dinb(new_new_n3693__), .dout(new_new_n2429__));
  and1  g1451(.dina(new_new_n2429__), .dinb(new_new_n3694__), .dout(new_new_n2430__));
  or1   g1452(.dina(new_new_n3695__), .dinb(new_new_n3248__), .dout(new_new_n2431__));
  and1  g1453(.dina(new_new_n3696__), .dinb(new_new_n3697__), .dout(new_new_n2432__));
  and1  g1454(.dina(new_new_n3698__), .dinb(new_new_n970__), .dout(new_new_n2433__));
  and1  g1455(.dina(new_new_n3701__), .dinb(new_new_n3704__), .dout(new_new_n2434__));
  and1  g1456(.dina(new_new_n3372__), .dinb(new_new_n3705__), .dout(new_new_n2435__));
  and1  g1457(.dina(new_new_n3708__), .dinb(new_new_n3712__), .dout(new_new_n2436__));
  or1   g1458(.dina(new_new_n2436__), .dinb(new_new_n1180__), .dout(new_new_n2437__));
  and1  g1459(.dina(new_new_n1288__), .dinb(new_new_n3516__), .dout(new_new_n2438__));
  and1  g1460(.dina(new_new_n1290__), .dinb(new_new_n3377__), .dout(new_new_n2439__));
  and1  g1461(.dina(new_new_n3671__), .dinb(new_new_n938__), .dout(new_new_n2440__));
  or1   g1462(.dina(new_new_n1222__), .dinb(new_new_n3269__), .dout(new_new_n2441__));
  and1  g1463(.dina(new_new_n2441__), .dinb(new_new_n1255__), .dout(new_new_n2442__));
  and1  g1464(.dina(new_new_n3226__), .dinb(new_new_n1279__), .dout(new_new_n2443__));
  and1  g1465(.dina(new_new_n3215__), .dinb(new_new_n3262__), .dout(new_new_n2444__));
  and1  g1466(.dina(new_new_n3216__), .dinb(new_new_n3231__), .dout(new_new_n2445__));
  or1   g1467(.dina(new_new_n3226__), .dinb(new_new_n3230__), .dout(new_new_n2446__));
  or1   g1468(.dina(new_new_n3714__), .dinb(new_new_n3715__), .dout(new_new_n2447__));
  and1  g1469(.dina(new_new_n3717__), .dinb(new_new_n3268__), .dout(new_new_n2448__));
  and1  g1470(.dina(new_new_n3701__), .dinb(new_new_n3718__), .dout(new_new_n2449__));
  or1   g1471(.dina(new_new_n3719__), .dinb(new_new_n3720__), .dout(new_new_n2450__));
  and1  g1472(.dina(new_new_n3702__), .dinb(new_new_n3721__), .dout(new_new_n2451__));
  and1  g1473(.dina(new_new_n3708__), .dinb(new_new_n3722__), .dout(new_new_n2452__));
  or1   g1474(.dina(new_new_n3656__), .dinb(new_new_n3349__), .dout(new_new_n2453__));
  and1  g1475(.dina(new_new_n3723__), .dinb(new_new_n3659__), .dout(new_new_n2454__));
  or1   g1476(.dina(new_new_n3723__), .dinb(new_new_n3660__), .dout(new_new_n2455__));
  and1  g1477(.dina(new_new_n3717__), .dinb(new_new_n3384__), .dout(new_new_n2456__));
  and1  g1478(.dina(new_new_n3724__), .dinb(new_new_n3725__), .dout(new_new_n2457__));
  or1   g1479(.dina(new_new_n1903__), .dinb(new_new_n3720__), .dout(new_new_n2458__));
  or1   g1480(.dina(new_new_n2458__), .dinb(new_new_n3668__), .dout(new_new_n2459__));
  and1  g1481(.dina(new_new_n3216__), .dinb(new_new_n3239__), .dout(new_new_n2460__));
  or1   g1482(.dina(new_new_n3227__), .dinb(new_new_n3238__), .dout(new_new_n2461__));
  and1  g1483(.dina(new_new_n2446__), .dinb(new_new_n3727__), .dout(new_new_n2462__));
  or1   g1484(.dina(new_new_n3714__), .dinb(new_new_n3667__), .dout(new_new_n2463__));
  and1  g1485(.dina(new_new_n2463__), .dinb(new_new_n2461__), .dout(new_new_n2464__));
  or1   g1486(.dina(new_new_n2462__), .dinb(new_new_n3728__), .dout(new_new_n2465__));
  and1  g1487(.dina(new_new_n2464__), .dinb(new_new_n3730__), .dout(new_new_n2466__));
  and1  g1488(.dina(new_new_n2465__), .dinb(new_new_n3666__), .dout(new_new_n2467__));
  or1   g1489(.dina(new_new_n2467__), .dinb(new_new_n2466__), .dout(new_new_n2468__));
  or1   g1490(.dina(new_new_n3731__), .dinb(new_new_n3733__), .dout(new_new_n2469__));
  and1  g1491(.dina(new_new_n3731__), .dinb(new_new_n3733__), .dout(new_new_n2470__));
  or1   g1492(.dina(new_new_n3734__), .dinb(new_new_n3736__), .dout(new_new_n2471__));
  or1   g1493(.dina(new_new_n3737__), .dinb(new_new_n3736__), .dout(new_new_n2472__));
  and1  g1494(.dina(new_new_n3738__), .dinb(new_new_n3739__), .dout(new_new_n2473__));
  and1  g1495(.dina(new_new_n2473__), .dinb(new_new_n3740__), .dout(new_new_n2474__));
  and1  g1496(.dina(new_new_n3365__), .dinb(new_new_n3742__), .dout(new_new_n2475__));
  and1  g1497(.dina(new_new_n3373__), .dinb(new_new_n3743__), .dout(new_new_n2476__));
  or1   g1498(.dina(new_new_n2476__), .dinb(new_new_n2475__), .dout(new_new_n2477__));
  or1   g1499(.dina(new_new_n3745__), .dinb(new_new_n3718__), .dout(new_new_n2478__));
  and1  g1500(.dina(new_new_n2478__), .dinb(new_new_n3747__), .dout(new_new_n2479__));
  or1   g1501(.dina(new_new_n2479__), .dinb(new_new_n3510__), .dout(new_new_n2480__));
  or1   g1502(.dina(new_new_n2480__), .dinb(new_new_n2477__), .dout(new_new_n2481__));
  and1  g1503(.dina(new_new_n3749__), .dinb(new_new_n1150__), .dout(new_new_n2482__));
  and1  g1504(.dina(new_new_n2482__), .dinb(new_new_n3750__), .dout(new_new_n2483__));
  and1  g1505(.dina(new_new_n3709__), .dinb(new_new_n1158__), .dout(new_new_n2484__));
  or1   g1506(.dina(new_new_n3752__), .dinb(new_new_n3366__), .dout(new_new_n2485__));
  and1  g1507(.dina(new_new_n2485__), .dinb(new_new_n3747__), .dout(new_new_n2486__));
  or1   g1508(.dina(new_new_n2486__), .dinb(new_new_n2484__), .dout(new_new_n2487__));
  or1   g1509(.dina(new_new_n3379__), .dinb(new_new_n3517__), .dout(new_new_n2488__));
  or1   g1510(.dina(new_new_n1198__), .dinb(new_new_n3374__), .dout(new_new_n2489__));
  and1  g1511(.dina(new_new_n2489__), .dinb(new_new_n2488__), .dout(new_new_n2490__));
  and1  g1512(.dina(new_new_n3753__), .dinb(new_new_n3754__), .dout(new_new_n2491__));
  or1   g1513(.dina(new_new_n3271__), .dinb(new_new_n917__), .dout(new_new_n2492__));
  and1  g1514(.dina(new_new_n2492__), .dinb(new_new_n3748__), .dout(new_new_n2493__));
  and1  g1515(.dina(new_new_n3756__), .dinb(new_new_n3742__), .dout(new_new_n2494__));
  or1   g1516(.dina(new_new_n2494__), .dinb(new_new_n2493__), .dout(new_new_n2495__));
  and1  g1517(.dina(new_new_n3756__), .dinb(new_new_n3381__), .dout(new_new_n2496__));
  and1  g1518(.dina(new_new_n3702__), .dinb(new_new_n3712__), .dout(new_new_n2497__));
  and1  g1519(.dina(new_new_n3709__), .dinb(new_new_n3383__), .dout(new_new_n2498__));
  or1   g1520(.dina(new_new_n2498__), .dinb(new_new_n2497__), .dout(new_new_n2499__));
  or1   g1521(.dina(new_new_n2499__), .dinb(new_new_n2496__), .dout(new_new_n2500__));
  and1  g1522(.dina(new_new_n3728__), .dinb(new_new_n3730__), .dout(new_new_n2501__));
  and1  g1523(.dina(new_new_n3347__), .dinb(new_new_n3348__), .dout(new_new_n2502__));
  or1   g1524(.dina(new_new_n2502__), .dinb(new_new_n2501__), .dout(new_new_n2503__));
  and1  g1525(.dina(new_new_n3757__), .dinb(new_new_n3758__), .dout(new_new_n2504__));
  or1   g1526(.dina(new_new_n3662__), .dinb(new_new_n3229__), .dout(new_new_n2505__));
  or1   g1527(.dina(new_new_n3661__), .dinb(new_new_n3237__), .dout(new_new_n2506__));
  or1   g1528(.dina(new_new_n3660__), .dinb(new_new_n3346__), .dout(new_new_n2507__));
  and1  g1529(.dina(new_new_n2507__), .dinb(new_new_n2287__), .dout(new_new_n2508__));
  and1  g1530(.dina(new_new_n2508__), .dinb(new_new_n2506__), .dout(new_new_n2509__));
  and1  g1531(.dina(new_new_n2509__), .dinb(new_new_n2505__), .dout(new_new_n2510__));
  or1   g1532(.dina(new_new_n3759__), .dinb(new_new_n944__), .dout(new_new_n2511__));
  and1  g1533(.dina(new_new_n3414__), .dinb(new_new_n3444__), .dout(new_new_n2512__));
  and1  g1534(.dina(new_new_n3761__), .dinb(new_new_n3399__), .dout(new_new_n2513__));
  or1   g1535(.dina(new_new_n2513__), .dinb(new_new_n2512__), .dout(new_new_n2514__));
  and1  g1536(.dina(new_new_n2514__), .dinb(new_new_n3423__), .dout(new_new_n2515__));
  or1   g1537(.dina(new_new_n3437__), .dinb(new_new_n3408__), .dout(new_new_n2516__));
  or1   g1538(.dina(new_new_n3479__), .dinb(new_new_n3442__), .dout(new_new_n2517__));
  or1   g1539(.dina(new_new_n3477__), .dinb(new_new_n3450__), .dout(new_new_n2518__));
  and1  g1540(.dina(new_new_n2518__), .dinb(new_new_n3386__), .dout(new_new_n2519__));
  or1   g1541(.dina(new_new_n3763__), .dinb(new_new_n2517__), .dout(new_new_n2520__));
  and1  g1542(.dina(new_new_n2520__), .dinb(new_new_n2516__), .dout(new_new_n2521__));
  or1   g1543(.dina(new_new_n2521__), .dinb(new_new_n2515__), .dout(new_new_n2522__));
  or1   g1544(.dina(new_new_n3713__), .dinb(new_new_n3765__), .dout(new_new_n2523__));
  or1   g1545(.dina(new_new_n2457__), .dinb(new_new_n3727__), .dout(new_new_n2524__));
  and1  g1546(.dina(new_new_n2524__), .dinb(new_new_n3732__), .dout(new_new_n2525__));
  or1   g1547(.dina(new_new_n3766__), .dinb(new_new_n3767__), .dout(new_new_n2526__));
  and1  g1548(.dina(new_new_n3766__), .dinb(new_new_n3767__), .dout(new_new_n2527__));
  and1  g1549(.dina(new_new_n3481__), .dinb(new_new_n3411__), .dout(new_new_n2528__));
  and1  g1550(.dina(new_new_n3440__), .dinb(new_new_n3356__), .dout(new_new_n2529__));
  and1  g1551(.dina(new_new_n3436__), .dinb(new_new_n3486__), .dout(new_new_n2530__));
  or1   g1552(.dina(new_new_n2530__), .dinb(new_new_n2529__), .dout(new_new_n2531__));
  and1  g1553(.dina(new_new_n2531__), .dinb(new_new_n3423__), .dout(new_new_n2532__));
  and1  g1554(.dina(new_new_n3763__), .dinb(new_new_n3333__), .dout(new_new_n2533__));
  or1   g1555(.dina(new_new_n2533__), .dinb(new_new_n2532__), .dout(new_new_n2534__));
  or1   g1556(.dina(new_new_n2534__), .dinb(new_new_n2528__), .dout(new_new_n2535__));
  and1  g1557(.dina(new_new_n3364__), .dinb(new_new_n3745__), .dout(new_new_n2536__));
  and1  g1558(.dina(new_new_n3768__), .dinb(new_new_n3373__), .dout(new_new_n2537__));
  or1   g1559(.dina(new_new_n2537__), .dinb(new_new_n2536__), .dout(new_new_n2538__));
  and1  g1560(.dina(new_new_n3769__), .dinb(new_new_n3500__), .dout(new_new_n2539__));
  or1   g1561(.dina(new_new_n1600__), .dinb(new_new_n3498__), .dout(new_new_n2540__));
  and1  g1562(.dina(new_new_n1584__), .dinb(new_new_n1581__), .dout(new_new_n2541__));
  or1   g1563(.dina(new_new_n1583__), .dinb(new_new_n1582__), .dout(new_new_n2542__));
  and1  g1564(.dina(new_new_n3771__), .dinb(new_new_n3772__), .dout(new_new_n2543__));
  or1   g1565(.dina(new_new_n3774__), .dinb(new_new_n1500__), .dout(new_new_n2544__));
  and1  g1566(.dina(new_new_n2544__), .dinb(new_new_n2542__), .dout(new_new_n2545__));
  or1   g1567(.dina(new_new_n2543__), .dinb(new_new_n2541__), .dout(new_new_n2546__));
  and1  g1568(.dina(new_new_n2545__), .dinb(new_new_n2540__), .dout(new_new_n2547__));
  or1   g1569(.dina(new_new_n2546__), .dinb(new_new_n2539__), .dout(new_new_n2548__));
  and1  g1570(.dina(new_new_n2548__), .dinb(new_new_n3456__), .dout(new_new_n2549__));
  or1   g1571(.dina(new_new_n2547__), .dinb(new_new_n3462__), .dout(new_new_n2550__));
  and1  g1572(.dina(new_new_n2550__), .dinb(new_new_n3502__), .dout(new_new_n2551__));
  or1   g1573(.dina(new_new_n2549__), .dinb(new_new_n3504__), .dout(new_new_n2552__));
  or1   g1574(.dina(new_new_n3775__), .dinb(new_new_n3497__), .dout(new_new_n2553__));
  or1   g1575(.dina(new_new_n2553__), .dinb(new_new_n2411__), .dout(new_new_n2554__));
  and1  g1576(.dina(new_new_n3748__), .dinb(new_new_n1156__), .dout(new_new_n2555__));
  or1   g1577(.dina(new_new_n2555__), .dinb(new_new_n3776__), .dout(new_new_n2556__));
  and1  g1578(.dina(new_new_n3703__), .dinb(new_new_n3752__), .dout(new_new_n2557__));
  and1  g1579(.dina(new_new_n3710__), .dinb(new_new_n3704__), .dout(new_new_n2558__));
  or1   g1580(.dina(new_new_n2558__), .dinb(new_new_n2557__), .dout(new_new_n2559__));
  or1   g1581(.dina(new_new_n2559__), .dinb(new_new_n3777__), .dout(new_new_n2560__));
  or1   g1582(.dina(new_new_n2560__), .dinb(new_new_n2556__), .dout(new_new_n2561__));
  and1  g1583(.dina(new_new_n3778__), .dinb(new_new_n3687__), .dout(new_new_n2562__));
  or1   g1584(.dina(new_new_n2562__), .dinb(new_new_n3779__), .dout(new_new_n2563__));
  and1  g1585(.dina(new_new_n2563__), .dinb(new_new_n3780__), .dout(new_new_n2564__));
  and1  g1586(.dina(new_new_n3781__), .dinb(new_new_n3782__), .dout(new_new_n2565__));
  or1   g1587(.dina(new_new_n891__), .dinb(new_new_n3786__), .dout(new_new_n2566__));
  or1   g1588(.dina(new_new_n3793__), .dinb(new_new_n3795__), .dout(new_new_n2567__));
  or1   g1589(.dina(new_new_n3797__), .dinb(new_new_n3793__), .dout(new_new_n2568__));
  and1  g1590(.dina(new_new_n3441__), .dinb(new_new_n3798__), .dout(new_new_n2569__));
  and1  g1591(.dina(new_new_n3445__), .dinb(new_new_n3761__), .dout(new_new_n2570__));
  and1  g1592(.dina(new_new_n3799__), .dinb(new_new_n3474__), .dout(new_new_n2571__));
  or1   g1593(.dina(new_new_n2571__), .dinb(new_new_n2570__), .dout(new_new_n2572__));
  or1   g1594(.dina(new_new_n2572__), .dinb(new_new_n2569__), .dout(new_new_n2573__));
  and1  g1595(.dina(new_new_n2573__), .dinb(new_new_n3424__), .dout(new_new_n2574__));
  and1  g1596(.dina(new_new_n3441__), .dinb(new_new_n3800__), .dout(new_new_n2575__));
  and1  g1597(.dina(new_new_n3411__), .dinb(new_new_n3760__), .dout(new_new_n2576__));
  and1  g1598(.dina(new_new_n3801__), .dinb(new_new_n3476__), .dout(new_new_n2577__));
  or1   g1599(.dina(new_new_n2577__), .dinb(new_new_n2576__), .dout(new_new_n2578__));
  or1   g1600(.dina(new_new_n2578__), .dinb(new_new_n2575__), .dout(new_new_n2579__));
  and1  g1601(.dina(new_new_n2579__), .dinb(new_new_n3424__), .dout(new_new_n2580__));
  and1  g1602(.dina(new_new_n3470__), .dinb(new_new_n3803__), .dout(new_new_n2581__));
  or1   g1603(.dina(new_new_n3438__), .dinb(new_new_n3806__), .dout(new_new_n2582__));
  or1   g1604(.dina(new_new_n3809__), .dinb(new_new_n3811__), .dout(new_new_n2583__));
  and1  g1605(.dina(new_new_n2583__), .dinb(new_new_n2582__), .dout(new_new_n2584__));
  and1  g1606(.dina(new_new_n3771__), .dinb(new_new_n947__), .dout(new_new_n2585__));
  or1   g1607(.dina(new_new_n2585__), .dinb(new_new_n2584__), .dout(new_new_n2586__));
  or1   g1608(.dina(new_new_n2586__), .dinb(new_new_n2581__), .dout(new_new_n2587__));
  and1  g1609(.dina(new_new_n2587__), .dinb(new_new_n3456__), .dout(new_new_n2588__));
  or1   g1610(.dina(new_new_n3812__), .dinb(new_new_n3778__), .dout(new_new_n2589__));
  or1   g1611(.dina(new_new_n3692__), .dinb(new_new_n3683__), .dout(new_new_n2590__));
  or1   g1612(.dina(new_new_n2590__), .dinb(new_new_n2589__), .dout(new_new_n2591__));
  and1  g1613(.dina(new_new_n2591__), .dinb(new_new_n3360__), .dout(new_new_n2592__));
  or1   g1614(.dina(new_new_n3775__), .dinb(new_new_n3682__), .dout(new_new_n2593__));
  or1   g1615(.dina(new_new_n3506__), .dinb(new_new_n3494__), .dout(new_new_n2594__));
  or1   g1616(.dina(new_new_n2594__), .dinb(new_new_n2593__), .dout(new_new_n2595__));
  and1  g1617(.dina(new_new_n2595__), .dinb(new_new_n3358__), .dout(new_new_n2596__));
  and1  g1618(.dina(new_new_n3469__), .dinb(new_new_n3813__), .dout(new_new_n2597__));
  or1   g1619(.dina(new_new_n3393__), .dinb(new_new_n3806__), .dout(new_new_n2598__));
  or1   g1620(.dina(new_new_n3803__), .dinb(new_new_n3809__), .dout(new_new_n2599__));
  and1  g1621(.dina(new_new_n2599__), .dinb(new_new_n2598__), .dout(new_new_n2600__));
  and1  g1622(.dina(new_new_n3770__), .dinb(new_new_n3811__), .dout(new_new_n2601__));
  or1   g1623(.dina(new_new_n2601__), .dinb(new_new_n2600__), .dout(new_new_n2602__));
  or1   g1624(.dina(new_new_n2602__), .dinb(new_new_n2597__), .dout(new_new_n2603__));
  and1  g1625(.dina(new_new_n2603__), .dinb(new_new_n3455__), .dout(new_new_n2604__));
  or1   g1626(.dina(new_new_n2604__), .dinb(new_new_n3814__), .dout(new_new_n2605__));
  or1   g1627(.dina(new_new_n3817__), .dinb(new_new_n3821__), .dout(new_new_n2606__));
  or1   g1628(.dina(new_new_n3823__), .dinb(new_new_n3824__), .dout(new_new_n2607__));
  and1  g1629(.dina(new_new_n3826__), .dinb(new_new_n3786__), .dout(new_new_n2608__));
  or1   g1630(.dina(new_new_n3764__), .dinb(new_new_n1560__), .dout(new_new_n2609__));
  or1   g1631(.dina(new_new_n3357__), .dinb(new_new_n3408__), .dout(new_new_n2610__));
  and1  g1632(.dina(new_new_n2610__), .dinb(new_new_n2609__), .dout(new_new_n2611__));
  or1   g1633(.dina(new_new_n3764__), .dinb(new_new_n3445__), .dout(new_new_n2612__));
  or1   g1634(.dina(new_new_n3336__), .dinb(new_new_n3407__), .dout(new_new_n2613__));
  and1  g1635(.dina(new_new_n2613__), .dinb(new_new_n2612__), .dout(new_new_n2614__));
  or1   g1636(.dina(new_new_n3466__), .dinb(new_new_n1394__), .dout(new_new_n2615__));
  and1  g1637(.dina(new_new_n3482__), .dinb(new_new_n3810__), .dout(new_new_n2616__));
  and1  g1638(.dina(new_new_n3827__), .dinb(new_new_n3805__), .dout(new_new_n2617__));
  or1   g1639(.dina(new_new_n2617__), .dinb(new_new_n2616__), .dout(new_new_n2618__));
  or1   g1640(.dina(new_new_n3828__), .dinb(new_new_n3774__), .dout(new_new_n2619__));
  and1  g1641(.dina(new_new_n2619__), .dinb(new_new_n2618__), .dout(new_new_n2620__));
  and1  g1642(.dina(new_new_n2620__), .dinb(new_new_n2615__), .dout(new_new_n2621__));
  or1   g1643(.dina(new_new_n2621__), .dinb(new_new_n3462__), .dout(new_new_n2622__));
  and1  g1644(.dina(new_new_n2622__), .dinb(new_new_n3829__), .dout(new_new_n2623__));
  and1  g1645(.dina(new_new_n3830__), .dinb(new_new_n3832__), .dout(new_new_n2624__));
  and1  g1646(.dina(new_new_n2624__), .dinb(new_new_n3834__), .dout(new_new_n2625__));
  or1   g1647(.dina(new_new_n3465__), .dinb(new_new_n3827__), .dout(new_new_n2626__));
  and1  g1648(.dina(new_new_n3434__), .dinb(new_new_n3810__), .dout(new_new_n2627__));
  and1  g1649(.dina(new_new_n3828__), .dinb(new_new_n3807__), .dout(new_new_n2628__));
  or1   g1650(.dina(new_new_n2628__), .dinb(new_new_n2627__), .dout(new_new_n2629__));
  or1   g1651(.dina(new_new_n1598__), .dinb(new_new_n3773__), .dout(new_new_n2630__));
  and1  g1652(.dina(new_new_n2630__), .dinb(new_new_n2629__), .dout(new_new_n2631__));
  and1  g1653(.dina(new_new_n2631__), .dinb(new_new_n2626__), .dout(new_new_n2632__));
  or1   g1654(.dina(new_new_n2632__), .dinb(new_new_n3461__), .dout(new_new_n2633__));
  and1  g1655(.dina(new_new_n2633__), .dinb(new_new_n3829__), .dout(new_new_n2634__));
  and1  g1656(.dina(new_new_n3835__), .dinb(new_new_n3832__), .dout(new_new_n2635__));
  and1  g1657(.dina(new_new_n2635__), .dinb(new_new_n3837__), .dout(new_new_n2636__));
  and1  g1658(.dina(new_new_n3830__), .dinb(new_new_n3687__), .dout(new_new_n2637__));
  or1   g1659(.dina(new_new_n2637__), .dinb(new_new_n3834__), .dout(new_new_n2638__));
  and1  g1660(.dina(new_new_n3835__), .dinb(new_new_n3689__), .dout(new_new_n2639__));
  or1   g1661(.dina(new_new_n2639__), .dinb(new_new_n3837__), .dout(new_new_n2640__));
  or1   g1662(.dina(new_new_n3734__), .dinb(new_new_n3839__), .dout(new_new_n2641__));
  or1   g1663(.dina(new_new_n3824__), .dinb(new_new_n3839__), .dout(new_new_n2642__));
  or1   g1664(.dina(new_new_n2642__), .dinb(new_new_n3817__), .dout(new_new_n2643__));
  and1  g1665(.dina(new_new_n2643__), .dinb(new_new_n3840__), .dout(new_new_n2644__));
  or1   g1666(.dina(new_new_n3842__), .dinb(new_new_n3826__), .dout(new_new_n2645__));
  or1   g1667(.dina(new_new_n3843__), .dinb(new_new_n996__), .dout(new_new_n2646__));
  and1  g1668(.dina(new_new_n3812__), .dinb(new_new_n3689__), .dout(new_new_n2647__));
  or1   g1669(.dina(new_new_n2647__), .dinb(new_new_n3844__), .dout(new_new_n2648__));
  and1  g1670(.dina(new_new_n2648__), .dinb(new_new_n3845__), .dout(new_new_n2649__));
  and1  g1671(.dina(new_new_n3846__), .dinb(new_new_n3847__), .dout(new_new_n2650__));
  or1   g1672(.dina(new_new_n3848__), .dinb(new_new_n818__), .dout(new_new_n2651__));
  and1  g1673(.dina(new_new_n2651__), .dinb(new_new_n3849__), .dout(new_new_n2652__));
  and1  g1674(.dina(new_new_n3787__), .dinb(new_new_n3838__), .dout(new_new_n2653__));
  or1   g1675(.dina(new_new_n3787__), .dinb(new_new_n3821__), .dout(new_new_n2654__));
  or1   g1676(.dina(new_new_n3850__), .dinb(new_new_n3797__), .dout(new_new_n2655__));
  and1  g1677(.dina(new_new_n2655__), .dinb(new_new_n3820__), .dout(new_new_n2656__));
  and1  g1678(.dina(new_new_n3851__), .dinb(new_new_n3822__), .dout(new_new_n2657__));
  or1   g1679(.dina(new_new_n3852__), .dinb(new_new_n3788__), .dout(new_new_n2658__));
  and1  g1680(.dina(new_new_n866__), .dinb(new_new_n3788__), .dout(new_new_n2659__));
  or1   g1681(.dina(new_new_n3854__), .dinb(new_new_n3794__), .dout(new_new_n2660__));
  or1   g1682(.dina(new_new_n3854__), .dinb(new_new_n3848__), .dout(new_new_n2661__));
  or1   g1683(.dina(new_new_n3857__), .dinb(new_new_n3859__), .dout(new_new_n2662__));
  or1   g1684(.dina(new_new_n3840__), .dinb(new_new_n3860__), .dout(new_new_n2663__));
  and1  g1685(.dina(new_new_n3861__), .dinb(new_new_n3863__), .dout(new_new_n2664__));
  or1   g1686(.dina(new_new_n3857__), .dinb(new_new_n858__), .dout(new_new_n2665__));
  and1  g1687(.dina(new_new_n3864__), .dinb(new_new_n3865__), .dout(new_new_n2666__));
  or1   g1688(.dina(new_new_n3866__), .dinb(new_new_n3790__), .dout(new_new_n2667__));
  or1   g1689(.dina(new_new_n3863__), .dinb(new_new_n3816__), .dout(new_new_n2668__));
  and1  g1690(.dina(new_new_n2668__), .dinb(new_new_n2667__), .dout(new_new_n2669__));
  and1  g1691(.dina(new_new_n872__), .dinb(new_new_n3818__), .dout(new_new_n2670__));
  and1  g1692(.dina(new_new_n3859__), .dinb(new_new_n3790__), .dout(new_new_n2671__));
  or1   g1693(.dina(new_new_n2671__), .dinb(new_new_n2670__), .dout(new_new_n2672__));
  or1   g1694(.dina(new_new_n3858__), .dinb(new_new_n860__), .dout(new_new_n2673__));
  and1  g1695(.dina(new_new_n2673__), .dinb(new_new_n2672__), .dout(new_new_n2674__));
  and1  g1696(.dina(new_new_n3867__), .dinb(new_new_n3791__), .dout(new_new_n2675__));
  and1  g1697(.dina(new_new_n3868__), .dinb(new_new_n3818__), .dout(new_new_n2676__));
  or1   g1698(.dina(new_new_n2676__), .dinb(new_new_n2675__), .dout(new_new_n2677__));
  and1  g1699(.dina(new_new_n3842__), .dinb(new_new_n3869__), .dout(new_new_n2678__));
  or1   g1700(.dina(new_new_n2678__), .dinb(new_new_n2677__), .dout(new_new_n2679__));
  buf1  g1701(.din(new_new_n1617__), .dout(G3519));
  buf1  g1702(.din(new_new_n1090__), .dout(G3520));
  buf1  g1703(.din(new_new_n1642__), .dout(G3521));
  buf1  g1704(.din(new_new_n1681__), .dout(G3522));
  buf1  g1705(.din(new_new_n1700__), .dout(G3523));
  buf1  g1706(.din(new_new_n1701__), .dout(G3524));
  buf1  g1707(.din(new_new_n1703__), .dout(G3525));
  buf1  g1708(.din(new_new_n1095__), .dout(G3526));
  buf1  g1709(.din(new_new_n1706__), .dout(G3527));
  buf1  g1710(.din(new_new_n3146__), .dout(G3528));
  buf1  g1711(.din(new_new_n3134__), .dout(G3529));
  buf1  g1712(.din(new_new_n1748__), .dout(G3530));
  buf1  g1713(.din(new_new_n3140__), .dout(G3531));
  buf1  g1714(.din(new_new_n3144__), .dout(G3532));
  buf1  g1715(.din(new_new_n3138__), .dout(G3533));
  buf1  g1716(.din(new_new_n1247__), .dout(G3534));
  buf1  g1717(.din(new_new_n1249__), .dout(G3535));
  buf1  g1718(.din(new_new_n3132__), .dout(G3536));
  buf1  g1719(.din(new_new_n3155__), .dout(G3537));
  not1  g1720(.din(new_new_n1786__), .dout(G3538));
  buf1  g1721(.din(new_new_n1823__), .dout(G3539));
  buf1  g1722(.din(new_new_n1832__), .dout(G3540));
  buf1  g1723(.din(new_new_n3192__), .dout(n6268));
  buf1  g1724(.din(new_new_n3310__), .dout(n6271));
  buf1  g1725(.din(new_new_n3180__), .dout(n6274));
  buf1  g1726(.din(new_new_n3586__), .dout(n6277));
  buf1  g1727(.din(new_new_n1081__), .dout(n6280));
  buf1  g1728(.din(new_new_n1083__), .dout(n6283));
  buf1  g1729(.din(new_new_n3592__), .dout(n6286));
  buf1  g1730(.din(new_new_n3588__), .dout(n6289));
  buf1  g1731(.din(new_new_n3593__), .dout(n6292));
  buf1  g1732(.din(new_new_n3591__), .dout(n6295));
  buf1  g1733(.din(new_new_n823__), .dout(n6298));
  buf1  g1734(.din(new_new_n915__), .dout(n6301));
  buf1  g1735(.din(new_new_n825__), .dout(n6304));
  buf1  g1736(.din(new_new_n919__), .dout(n6307));
  buf1  g1737(.din(new_new_n827__), .dout(n6310));
  buf1  g1738(.din(new_new_n923__), .dout(n6313));
  buf1  g1739(.din(new_new_n829__), .dout(n6316));
  buf1  g1740(.din(new_new_n927__), .dout(n6319));
  buf1  g1741(.din(new_new_n831__), .dout(n6322));
  buf1  g1742(.din(new_new_n931__), .dout(n6325));
  buf1  g1743(.din(new_new_n833__), .dout(n6328));
  buf1  g1744(.din(new_new_n935__), .dout(n6331));
  buf1  g1745(.din(new_new_n835__), .dout(n6334));
  buf1  g1746(.din(new_new_n837__), .dout(n6337));
  buf1  g1747(.din(new_new_n847__), .dout(n6340));
  buf1  g1748(.din(new_new_n1129__), .dout(n6343));
  buf1  g1749(.din(new_new_n849__), .dout(n6346));
  buf1  g1750(.din(new_new_n851__), .dout(n6349));
  buf1  g1751(.din(new_new_n1091__), .dout(n6352));
  buf1  g1752(.din(new_new_n1085__), .dout(n6355));
  buf1  g1753(.din(new_new_n1069__), .dout(n6358));
  buf1  g1754(.din(new_new_n1047__), .dout(n6361));
  buf1  g1755(.din(new_new_n1049__), .dout(n6364));
  buf1  g1756(.din(new_new_n1059__), .dout(n6367));
  buf1  g1757(.din(new_new_n1071__), .dout(n6370));
  buf1  g1758(.din(new_new_n1093__), .dout(n6373));
  buf1  g1759(.din(new_new_n877__), .dout(n6376));
  buf1  g1760(.din(new_new_n967__), .dout(n6379));
  buf1  g1761(.din(new_new_n879__), .dout(n6382));
  buf1  g1762(.din(new_new_n971__), .dout(n6385));
  buf1  g1763(.din(new_new_n881__), .dout(n6388));
  buf1  g1764(.din(new_new_n975__), .dout(n6391));
  buf1  g1765(.din(new_new_n883__), .dout(n6394));
  buf1  g1766(.din(new_new_n979__), .dout(n6397));
  buf1  g1767(.din(new_new_n885__), .dout(n6400));
  buf1  g1768(.din(new_new_n983__), .dout(n6403));
  buf1  g1769(.din(new_new_n985__), .dout(n6406));
  buf1  g1770(.din(new_new_n887__), .dout(n6409));
  buf1  g1771(.din(new_new_n989__), .dout(n6412));
  buf1  g1772(.din(new_new_n3288__), .dout(n6415));
  buf1  g1773(.din(new_new_n889__), .dout(n6418));
  buf1  g1774(.din(new_new_n1137__), .dout(n6421));
  buf1  g1775(.din(new_new_n893__), .dout(n6424));
  buf1  g1776(.din(new_new_n999__), .dout(n6427));
  buf1  g1777(.din(new_new_n1001__), .dout(n6430));
  buf1  g1778(.din(new_new_n1003__), .dout(n6433));
  buf1  g1779(.din(new_new_n3311__), .dout(n6436));
  buf1  g1780(.din(new_new_n1065__), .dout(n6439));
  buf1  g1781(.din(new_new_n1079__), .dout(n6442));
  buf1  g1782(.din(new_new_n1113__), .dout(n6445));
  buf1  g1783(.din(new_new_n1117__), .dout(n6448));
  buf1  g1784(.din(new_new_n1123__), .dout(n6451));
  buf1  g1785(.din(new_new_n3187__), .dout(n6454));
  buf1  g1786(.din(new_new_n1145__), .dout(n6457));
  buf1  g1787(.din(new_new_n1215__), .dout(n6460));
  buf1  g1788(.din(new_new_n1217__), .dout(n6463));
  buf1  g1789(.din(new_new_n3549__), .dout(n6466));
  buf1  g1790(.din(new_new_n1141__), .dout(n6469));
  buf1  g1791(.din(new_new_n3248__), .dout(n6472));
  buf1  g1792(.din(new_new_n3695__), .dout(n6475));
  buf1  g1793(.din(new_new_n3509__), .dout(n6478));
  buf1  g1794(.din(new_new_n1151__), .dout(n6481));
  buf1  g1795(.din(new_new_n3697__), .dout(n6484));
  buf1  g1796(.din(new_new_n3672__), .dout(n6487));
  buf1  g1797(.din(new_new_n3369__), .dout(n6490));
  buf1  g1798(.din(new_new_n3698__), .dout(n6493));
  buf1  g1799(.din(new_new_n1161__), .dout(n6496));
  buf1  g1800(.din(new_new_n1163__), .dout(n6499));
  buf1  g1801(.din(new_new_n3751__), .dout(n6502));
  buf1  g1802(.din(new_new_n1341__), .dout(n6505));
  buf1  g1803(.din(new_new_n1345__), .dout(n6508));
  buf1  g1804(.din(new_new_n3749__), .dout(n6511));
  buf1  g1805(.din(new_new_n1171__), .dout(n6514));
  buf1  g1806(.din(new_new_n1173__), .dout(n6517));
  buf1  g1807(.din(new_new_n1167__), .dout(n6520));
  buf1  g1808(.din(new_new_n1175__), .dout(n6523));
  buf1  g1809(.din(new_new_n1177__), .dout(n6526));
  buf1  g1810(.din(new_new_n1181__), .dout(n6529));
  buf1  g1811(.din(new_new_n1183__), .dout(n6532));
  buf1  g1812(.din(new_new_n3705__), .dout(n6535));
  buf1  g1813(.din(new_new_n3285__), .dout(n6538));
  buf1  g1814(.din(new_new_n3185__), .dout(n6541));
  buf1  g1815(.din(new_new_n1187__), .dout(n6544));
  buf1  g1816(.din(new_new_n3517__), .dout(n6547));
  buf1  g1817(.din(new_new_n3379__), .dout(n6550));
  buf1  g1818(.din(new_new_n1199__), .dout(n6553));
  not1  g1819(.din(new_new_n3563__), .dout(n6556));
  not1  g1820(.din(new_new_n3564__), .dout(n6559));
  buf1  g1821(.din(new_new_n1207__), .dout(n6562));
  buf1  g1822(.din(new_new_n1209__), .dout(n6565));
  buf1  g1823(.din(new_new_n3534__), .dout(n6568));
  buf1  g1824(.din(new_new_n3326__), .dout(n6571));
  buf1  g1825(.din(new_new_n3292__), .dout(n6574));
  buf1  g1826(.din(new_new_n3696__), .dout(n6577));
  buf1  g1827(.din(new_new_n3670__), .dout(n6580));
  buf1  g1828(.din(new_new_n1223__), .dout(n6583));
  buf1  g1829(.din(new_new_n3194__), .dout(n6586));
  buf1  g1830(.din(new_new_n1251__), .dout(n6589));
  buf1  g1831(.din(new_new_n3562__), .dout(n6592));
  buf1  g1832(.din(new_new_n1275__), .dout(n6595));
  buf1  g1833(.din(new_new_n1277__), .dout(n6598));
  buf1  g1834(.din(new_new_n1281__), .dout(n6601));
  buf1  g1835(.din(new_new_n3741__), .dout(n6604));
  buf1  g1836(.din(new_new_n3380__), .dout(n6607));
  buf1  g1837(.din(new_new_n1283__), .dout(n6610));
  buf1  g1838(.din(new_new_n3322__), .dout(n6613));
  buf1  g1839(.din(new_new_n3264__), .dout(n6616));
  buf1  g1840(.din(new_new_n1369__), .dout(n6619));
  buf1  g1841(.din(new_new_n1339__), .dout(n6622));
  buf1  g1842(.din(new_new_n3263__), .dout(n6625));
  buf1  g1843(.din(new_new_n1377__), .dout(n6628));
  buf1  g1844(.din(new_new_n1453__), .dout(n6631));
  buf1  g1845(.din(new_new_n3227__), .dout(n6634));
  buf1  g1846(.din(new_new_n3450__), .dout(n6637));
  buf1  g1847(.din(new_new_n3476__), .dout(n6640));
  buf1  g1848(.din(new_new_n3228__), .dout(n6643));
  buf1  g1849(.din(new_new_n3447__), .dout(n6646));
  buf1  g1850(.din(new_new_n3807__), .dout(n6649));
  buf1  g1851(.din(new_new_n3464__), .dout(n6652));
  buf1  g1852(.din(new_new_n3393__), .dout(n6655));
  buf1  g1853(.din(new_new_n3431__), .dout(n6658));
  buf1  g1854(.din(new_new_n3484__), .dout(n6661));
  buf1  g1855(.din(new_new_n3490__), .dout(n6664));
  buf1  g1856(.din(new_new_n1393__), .dout(n6667));
  buf1  g1857(.din(new_new_n1395__), .dout(n6670));
  buf1  g1858(.din(new_new_n3680__), .dout(n6673));
  buf1  g1859(.din(new_new_n1449__), .dout(n6676));
  buf1  g1860(.din(new_new_n3463__), .dout(n6679));
  buf1  g1861(.din(new_new_n3772__), .dout(n6682));
  buf1  g1862(.din(new_new_n1501__), .dout(n6685));
  buf1  g1863(.din(new_new_n1505__), .dout(n6688));
  buf1  g1864(.din(new_new_n1507__), .dout(n6691));
  buf1  g1865(.din(new_new_n1527__), .dout(n6694));
  buf1  g1866(.din(new_new_n1545__), .dout(n6697));
  buf1  g1867(.din(new_new_n3681__), .dout(n6700));
  buf1  g1868(.din(new_new_n1549__), .dout(n6703));
  buf1  g1869(.din(new_new_n1557__), .dout(n6706));
  buf1  g1870(.din(new_new_n3267__), .dout(n6709));
  buf1  g1871(.din(new_new_n3265__), .dout(n6712));
  buf1  g1872(.din(new_new_n3726__), .dout(n6715));
  buf1  g1873(.din(new_new_n3333__), .dout(n6718));
  buf1  g1874(.din(new_new_n3438__), .dout(n6721));
  buf1  g1875(.din(new_new_n3813__), .dout(n6724));
  buf1  g1876(.din(new_new_n3270__), .dout(n6727));
  buf1  g1877(.din(new_new_n3744__), .dout(n6730));
  buf1  g1878(.din(new_new_n3725__), .dout(n6733));
  buf1  g1879(.din(new_new_n3802__), .dout(n6736));
  buf1  g1880(.din(new_new_n3769__), .dout(n6739));
  not1  g1881(.din(new_new_n3703__), .dout(n6742));
  buf1  g1882(.din(new_new_n3710__), .dout(n6745));
  buf1  g1883(.din(new_new_n3272__), .dout(n6748));
  buf1  g1884(.din(new_new_n3724__), .dout(n6751));
  buf1  g1885(.din(new_new_n3357__), .dout(n6754));
  buf1  g1886(.din(new_new_n3336__), .dout(n6757));
  buf1  g1887(.din(new_new_n3361__), .dout(n6760));
  buf1  g1888(.din(new_new_n3359__), .dout(n6763));
  buf1  g1889(.din(new_new_n3363__), .dout(n6766));
  buf1  g1890(.din(new_new_n3362__), .dout(n6769));
  buf1  g1891(.din(new_new_n3711__), .dout(n6772));
  buf1  g1892(.din(new_new_n3382__), .dout(n6775));
  not1  g1893(.din(new_new_n3743__), .dout(n6778));
  buf1  g1894(.din(new_new_n1905__), .dout(n6781));
  buf1  g1895(.din(new_new_n3755__), .dout(n6784));
  buf1  g1896(.din(new_new_n3367__), .dout(n6787));
  buf1  g1897(.din(new_new_n3370__), .dout(n6790));
  buf1  g1898(.din(new_new_n3518__), .dout(n6793));
  buf1  g1899(.din(new_new_n3678__), .dout(n6796));
  buf1  g1900(.din(new_new_n3676__), .dout(n6799));
  buf1  g1901(.din(new_new_n3446__), .dout(n6802));
  buf1  g1902(.din(new_new_n3729__), .dout(n6805));
  buf1  g1903(.din(new_new_n3385__), .dout(n6808));
  buf1  g1904(.din(new_new_n3831__), .dout(n6811));
  buf1  g1905(.din(new_new_n3688__), .dout(n6814));
  not1  g1906(.din(new_new_n3777__), .dout(n6817));
  buf1  g1907(.din(new_new_n3508__), .dout(n6820));
  not1  g1908(.din(new_new_n3739__), .dout(n6823));
  not1  g1909(.din(new_new_n3776__), .dout(n6826));
  not1  g1910(.din(new_new_n3738__), .dout(n6829));
  buf1  g1911(.din(new_new_n3768__), .dout(n6832));
  buf1  g1912(.din(new_new_n3765__), .dout(n6835));
  buf1  g1913(.din(new_new_n3799__), .dout(n6838));
  buf1  g1914(.din(new_new_n3690__), .dout(n6841));
  buf1  g1915(.din(new_new_n3693__), .dout(n6844));
  buf1  g1916(.din(new_new_n3801__), .dout(n6847));
  buf1  g1917(.din(new_new_n3654__), .dout(n6850));
  buf1  g1918(.din(new_new_n3814__), .dout(n6853));
  buf1  g1919(.din(new_new_n3798__), .dout(n6856));
  buf1  g1920(.din(new_new_n3800__), .dout(n6859));
  buf1  g1921(.din(new_new_n3779__), .dout(n6862));
  not1  g1922(.din(new_new_n3691__), .dout(n6865));
  not1  g1923(.din(new_new_n3694__), .dout(n6868));
  buf1  g1924(.din(new_new_n3735__), .dout(n6871));
  buf1  g1925(.din(new_new_n3822__), .dout(n6874));
  buf1  g1926(.din(new_new_n3722__), .dout(n6877));
  buf1  g1927(.din(new_new_n3721__), .dout(n6880));
  not1  g1928(.din(new_new_n2096__), .dout(n6883));
  not1  g1929(.din(new_new_n2097__), .dout(n6886));
  buf1  g1930(.din(new_new_n3740__), .dout(n6889));
  not1  g1931(.din(new_new_n2100__), .dout(n6892));
  not1  g1932(.din(new_new_n3750__), .dout(n6895));
  buf1  g1933(.din(new_new_n3754__), .dout(n6898));
  buf1  g1934(.din(new_new_n2103__), .dout(n6901));
  buf1  g1935(.din(new_new_n2135__), .dout(n6904));
  buf1  g1936(.din(new_new_n2136__), .dout(n6907));
  buf1  g1937(.din(new_new_n2137__), .dout(n6910));
  buf1  g1938(.din(new_new_n2139__), .dout(n6913));
  not1  g1939(.din(new_new_n2180__), .dout(n6916));
  not1  g1940(.din(new_new_n2207__), .dout(n6919));
  buf1  g1941(.din(new_new_n2235__), .dout(n6922));
  buf1  g1942(.din(new_new_n2266__), .dout(n6925));
  not1  g1943(.din(new_new_n2275__), .dout(n6928));
  not1  g1944(.din(new_new_n3758__), .dout(n6931));
  buf1  g1945(.din(new_new_n3759__), .dout(n6934));
  not1  g1946(.din(new_new_n3716__), .dout(n6937));
  buf1  g1947(.din(new_new_n2295__), .dout(n6940));
  not1  g1948(.din(new_new_n3715__), .dout(n6943));
  buf1  g1949(.din(new_new_n2322__), .dout(n6946));
  buf1  g1950(.din(new_new_n2325__), .dout(n6949));
  buf1  g1951(.din(new_new_n2351__), .dout(n6952));
  buf1  g1952(.din(new_new_n2354__), .dout(n6955));
  buf1  g1953(.din(new_new_n3753__), .dout(n6958));
  buf1  g1954(.din(new_new_n2365__), .dout(n6961));
  buf1  g1955(.din(new_new_n2382__), .dout(n6964));
  buf1  g1956(.din(new_new_n2383__), .dout(n6967));
  buf1  g1957(.din(new_new_n2384__), .dout(n6970));
  not1  g1958(.din(new_new_n3757__), .dout(n6973));
  not1  g1959(.din(new_new_n3719__), .dout(n6976));
  buf1  g1960(.din(new_new_n943__), .dout(n6979));
  buf1  g1961(.din(new_new_n3844__), .dout(n6982));
  not1  g1962(.din(new_new_n3780__), .dout(n6985));
  buf1  g1963(.din(new_new_n3782__), .dout(n6988));
  buf1  g1964(.din(new_new_n3781__), .dout(n6991));
  buf1  g1965(.din(new_new_n797__), .dout(n6994));
  buf1  g1966(.din(new_new_n3791__), .dout(n6997));
  buf1  g1967(.din(new_new_n3737__), .dout(n7000));
  buf1  g1968(.din(new_new_n3795__), .dout(n7003));
  buf1  g1969(.din(new_new_n3794__), .dout(n7006));
  buf1  g1970(.din(new_new_n3796__), .dout(n7009));
  buf1  g1971(.din(new_new_n3868__), .dout(n7012));
  buf1  g1972(.din(new_new_n3867__), .dout(n7015));
  buf1  g1973(.din(new_new_n3869__), .dout(n7018));
  buf1  g1974(.din(new_new_n871__), .dout(n7021));
  buf1  g1975(.din(new_new_n977__), .dout(n7024));
  buf1  g1976(.din(new_new_n981__), .dout(n7027));
  buf1  g1977(.din(new_new_n2431__), .dout(n7030));
  buf1  g1978(.din(new_new_n2432__), .dout(n7033));
  buf1  g1979(.din(new_new_n2433__), .dout(n7036));
  not1  g1980(.din(new_new_n2434__), .dout(n7039));
  buf1  g1981(.din(new_new_n2435__), .dout(n7042));
  not1  g1982(.din(new_new_n2437__), .dout(n7045));
  buf1  g1983(.din(new_new_n2438__), .dout(n7048));
  buf1  g1984(.din(new_new_n2439__), .dout(n7051));
  buf1  g1985(.din(new_new_n2440__), .dout(n7054));
  buf1  g1986(.din(new_new_n2442__), .dout(n7057));
  buf1  g1987(.din(new_new_n2443__), .dout(n7060));
  buf1  g1988(.din(new_new_n2444__), .dout(n7063));
  not1  g1989(.din(new_new_n2447__), .dout(n7066));
  buf1  g1990(.din(new_new_n2448__), .dout(n7069));
  buf1  g1991(.din(new_new_n2449__), .dout(n7072));
  not1  g1992(.din(new_new_n2450__), .dout(n7075));
  buf1  g1993(.din(new_new_n2451__), .dout(n7078));
  buf1  g1994(.din(new_new_n2452__), .dout(n7081));
  not1  g1995(.din(new_new_n2454__), .dout(n7084));
  not1  g1996(.din(new_new_n2455__), .dout(n7087));
  not1  g1997(.din(new_new_n2456__), .dout(n7090));
  not1  g1998(.din(new_new_n2469__), .dout(n7093));
  buf1  g1999(.din(new_new_n2470__), .dout(n7096));
  not1  g2000(.din(new_new_n3823__), .dout(n7099));
  buf1  g2001(.din(new_new_n3841__), .dout(n7102));
  buf1  g2002(.din(new_new_n995__), .dout(n7105));
  buf1  g2003(.din(new_new_n2474__), .dout(n7108));
  not1  g2004(.din(new_new_n2481__), .dout(n7111));
  buf1  g2005(.din(new_new_n2483__), .dout(n7114));
  not1  g2006(.din(new_new_n2487__), .dout(n7117));
  buf1  g2007(.din(new_new_n2490__), .dout(n7120));
  buf1  g2008(.din(new_new_n2491__), .dout(n7123));
  buf1  g2009(.din(new_new_n2495__), .dout(n7126));
  buf1  g2010(.din(new_new_n2500__), .dout(n7129));
  buf1  g2011(.din(new_new_n2503__), .dout(n7132));
  not1  g2012(.din(new_new_n2504__), .dout(n7135));
  not1  g2013(.din(new_new_n2510__), .dout(n7138));
  not1  g2014(.din(new_new_n3843__), .dout(n7141));
  buf1  g2015(.din(new_new_n3833__), .dout(n7144));
  buf1  g2016(.din(new_new_n2526__), .dout(n7147));
  buf1  g2017(.din(new_new_n2527__), .dout(n7150));
  buf1  g2018(.din(new_new_n3836__), .dout(n7153));
  buf1  g2019(.din(new_new_n2538__), .dout(n7156));
  not1  g2020(.din(new_new_n3845__), .dout(n7159));
  not1  g2021(.din(new_new_n2561__), .dout(n7162));
  buf1  g2022(.din(new_new_n3847__), .dout(n7165));
  buf1  g2023(.din(new_new_n3846__), .dout(n7168));
  buf1  g2024(.din(new_new_n3825__), .dout(n7171));
  buf1  g2025(.din(new_new_n3862__), .dout(n7174));
  buf1  g2026(.din(new_new_n3866__), .dout(n7177));
  buf1  g2027(.din(new_new_n3858__), .dout(n7180));
  buf1  g2028(.din(new_new_n3850__), .dout(n7183));
  buf1  g2029(.din(new_new_n3849__), .dout(n7186));
  buf1  g2030(.din(new_new_n2574__), .dout(n7189));
  buf1  g2031(.din(new_new_n2580__), .dout(n7192));
  buf1  g2032(.din(new_new_n2588__), .dout(n7195));
  buf1  g2033(.din(new_new_n2592__), .dout(n7198));
  buf1  g2034(.din(new_new_n2596__), .dout(n7201));
  buf1  g2035(.din(new_new_n2605__), .dout(n7204));
  not1  g2036(.din(new_new_n3855__), .dout(n7207));
  buf1  g2037(.din(n7207), .dout(n7210));
  not1  g2038(.din(new_new_n3865__), .dout(n7213));
  buf1  g2039(.din(new_new_n3860__), .dout(n7216));
  buf1  g2040(.din(new_new_n2611__), .dout(n7219));
  buf1  g2041(.din(new_new_n2614__), .dout(n7222));
  buf1  g2042(.din(new_new_n2625__), .dout(n7225));
  buf1  g2043(.din(new_new_n2636__), .dout(n7228));
  buf1  g2044(.din(new_new_n2638__), .dout(n7231));
  buf1  g2045(.din(new_new_n2640__), .dout(n7234));
  not1  g2046(.din(new_new_n3864__), .dout(n7237));
  buf1  g2047(.din(new_new_n3861__), .dout(n7240));
  buf1  g2048(.din(new_new_n857__), .dout(n7243));
  buf1  g2049(.din(new_new_n865__), .dout(n7246));
  buf1  g2050(.din(new_new_n3852__), .dout(n7249));
  not1  g2051(.din(new_new_n2646__), .dout(n7252));
  buf1  g2052(.din(new_new_n2649__), .dout(n7255));
  buf1  g2053(.din(new_new_n2650__), .dout(n7258));
  buf1  g2054(.din(new_new_n3851__), .dout(n7261));
  buf1  g2055(.din(new_new_n807__), .dout(n7264));
  buf1  g2056(.din(new_new_n809__), .dout(n7267));
  buf1  g2057(.din(new_new_n839__), .dout(n7270));
  buf1  g2058(.din(new_new_n841__), .dout(n7273));
  buf1  g2059(.din(new_new_n843__), .dout(n7276));
  buf1  g2060(.din(new_new_n845__), .dout(n7279));
  buf1  g2061(.din(new_new_n2653__), .dout(n7282));
  buf1  g2062(.din(new_new_n3870__), .dout(n7285));
  buf1  g2063(.din(n7285), .dout(n7288));
  buf1  g2064(.din(new_new_n2656__), .dout(n7291));
  buf1  g2065(.din(new_new_n2657__), .dout(n7294));
  buf1  g2066(.din(new_new_n2658__), .dout(n7297));
  buf1  g2067(.din(new_new_n2659__), .dout(n7300));
  not1  g2068(.din(new_new_n2660__), .dout(n7303));
  not1  g2069(.din(new_new_n2661__), .dout(n7306));
  not1  g2070(.din(new_new_n2662__), .dout(n7309));
  not1  g2071(.din(new_new_n2663__), .dout(n7312));
  buf1  g2072(.din(new_new_n2664__), .dout(n7315));
  not1  g2073(.din(new_new_n2665__), .dout(n7318));
  buf1  g2074(.din(new_new_n853__), .dout(n7321));
  buf1  g2075(.din(new_new_n867__), .dout(n7324));
  not1  g2076(.din(new_new_n2666__), .dout(n7327));
  buf1  g2077(.din(new_new_n2669__), .dout(n7330));
  not1  g2078(.din(new_new_n2674__), .dout(n7333));
  buf1  g2079(.din(new_new_n2679__), .dout(n7336));
  buf1  g2080(.din(new_new_n811__), .dout(n7339));
  buf1  g2081(.din(new_new_n813__), .dout(n7342));
  buf1  g2082(.din(new_new_n855__), .dout(n7345));
  buf1  g2083(.din(new_new_n869__), .dout(n7348));
  buf1  g2084(.din(new_new_n906__), .dout(new_new_n3063__));
  buf1  g2085(.din(new_new_n898__), .dout(new_new_n3064__));
  buf1  g2086(.din(new_new_n896__), .dout(new_new_n3065__));
  buf1  g2087(.din(new_new_n960__), .dout(new_new_n3066__));
  buf1  g2088(.din(new_new_n3066__), .dout(new_new_n3067__));
  buf1  g2089(.din(new_new_n3066__), .dout(new_new_n3068__));
  buf1  g2090(.din(new_new_n907__), .dout(new_new_n3069__));
  buf1  g2091(.din(new_new_n956__), .dout(new_new_n3070__));
  buf1  g2092(.din(new_new_n3070__), .dout(new_new_n3071__));
  buf1  g2093(.din(new_new_n952__), .dout(new_new_n3072__));
  buf1  g2094(.din(new_new_n3072__), .dout(new_new_n3073__));
  buf1  g2095(.din(new_new_n899__), .dout(new_new_n3074__));
  buf1  g2096(.din(new_new_n958__), .dout(new_new_n3075__));
  buf1  g2097(.din(new_new_n3075__), .dout(new_new_n3076__));
  buf1  g2098(.din(new_new_n966__), .dout(new_new_n3077__));
  buf1  g2099(.din(new_new_n3077__), .dout(new_new_n3078__));
  buf1  g2100(.din(new_new_n913__), .dout(new_new_n3079__));
  buf1  g2101(.din(new_new_n3079__), .dout(new_new_n3080__));
  buf1  g2102(.din(new_new_n954__), .dout(new_new_n3081__));
  buf1  g2103(.din(new_new_n3081__), .dout(new_new_n3082__));
  buf1  g2104(.din(new_new_n962__), .dout(new_new_n3083__));
  buf1  g2105(.din(new_new_n3083__), .dout(new_new_n3084__));
  buf1  g2106(.din(new_new_n3083__), .dout(new_new_n3085__));
  buf1  g2107(.din(new_new_n909__), .dout(new_new_n3086__));
  buf1  g2108(.din(new_new_n964__), .dout(new_new_n3087__));
  buf1  g2109(.din(new_new_n3087__), .dout(new_new_n3088__));
  buf1  g2110(.din(new_new_n3087__), .dout(new_new_n3089__));
  buf1  g2111(.din(new_new_n911__), .dout(new_new_n3090__));
  buf1  g2112(.din(new_new_n3090__), .dout(new_new_n3091__));
  buf1  g2113(.din(new_new_n1636__), .dout(new_new_n3092__));
  buf1  g2114(.din(new_new_n963__), .dout(new_new_n3093__));
  buf1  g2115(.din(new_new_n965__), .dout(new_new_n3094__));
  buf1  g2116(.din(new_new_n959__), .dout(new_new_n3095__));
  buf1  g2117(.din(new_new_n961__), .dout(new_new_n3096__));
  buf1  g2118(.din(new_new_n1653__), .dout(new_new_n3097__));
  buf1  g2119(.din(new_new_n1648__), .dout(new_new_n3098__));
  buf1  g2120(.din(new_new_n1654__), .dout(new_new_n3099__));
  buf1  g2121(.din(new_new_n1647__), .dout(new_new_n3100__));
  buf1  g2122(.din(new_new_n955__), .dout(new_new_n3101__));
  buf1  g2123(.din(new_new_n957__), .dout(new_new_n3102__));
  buf1  g2124(.din(new_new_n951__), .dout(new_new_n3103__));
  buf1  g2125(.din(new_new_n953__), .dout(new_new_n3104__));
  buf1  g2126(.din(new_new_n1672__), .dout(new_new_n3105__));
  buf1  g2127(.din(new_new_n1665__), .dout(new_new_n3106__));
  buf1  g2128(.din(new_new_n1671__), .dout(new_new_n3107__));
  buf1  g2129(.din(new_new_n1666__), .dout(new_new_n3108__));
  buf1  g2130(.din(new_new_n914__), .dout(new_new_n3109__));
  buf1  g2131(.din(new_new_n3109__), .dout(new_new_n3110__));
  buf1  g2132(.din(new_new_n912__), .dout(new_new_n3111__));
  buf1  g2133(.din(new_new_n1690__), .dout(new_new_n3112__));
  buf1  g2134(.din(new_new_n1684__), .dout(new_new_n3113__));
  buf1  g2135(.din(new_new_n1691__), .dout(new_new_n3114__));
  buf1  g2136(.din(new_new_n1685__), .dout(new_new_n3115__));
  buf1  g2137(.din(new_new_n1053__), .dout(new_new_n3116__));
  buf1  g2138(.din(new_new_n1108__), .dout(new_new_n3117__));
  buf1  g2139(.din(new_new_n3117__), .dout(new_new_n3118__));
  buf1  g2140(.din(new_new_n1126__), .dout(new_new_n3119__));
  buf1  g2141(.din(new_new_n1125__), .dout(new_new_n3120__));
  buf1  g2142(.din(new_new_n1720__), .dout(new_new_n3121__));
  buf1  g2143(.din(new_new_n1075__), .dout(new_new_n3122__));
  buf1  g2144(.din(new_new_n1719__), .dout(new_new_n3123__));
  buf1  g2145(.din(new_new_n1076__), .dout(new_new_n3124__));
  buf1  g2146(.din(new_new_n1099__), .dout(new_new_n3125__));
  buf1  g2147(.din(new_new_n1097__), .dout(new_new_n3126__));
  buf1  g2148(.din(new_new_n1100__), .dout(new_new_n3127__));
  buf1  g2149(.din(new_new_n1098__), .dout(new_new_n3128__));
  buf1  g2150(.din(new_new_n1107__), .dout(new_new_n3129__));
  buf1  g2151(.din(new_new_n1771__), .dout(new_new_n3130__));
  buf1  g2152(.din(new_new_n1717__), .dout(new_new_n3131__));
  buf1  g2153(.din(new_new_n1772__), .dout(new_new_n3132__));
  buf1  g2154(.din(new_new_n3132__), .dout(new_new_n3133__));
  buf1  g2155(.din(new_new_n1718__), .dout(new_new_n3134__));
  buf1  g2156(.din(new_new_n3134__), .dout(new_new_n3135__));
  buf1  g2157(.din(new_new_n1765__), .dout(new_new_n3136__));
  buf1  g2158(.din(new_new_n1753__), .dout(new_new_n3137__));
  buf1  g2159(.din(new_new_n1766__), .dout(new_new_n3138__));
  buf1  g2160(.din(new_new_n3138__), .dout(new_new_n3139__));
  buf1  g2161(.din(new_new_n1754__), .dout(new_new_n3140__));
  buf1  g2162(.din(new_new_n3140__), .dout(new_new_n3141__));
  buf1  g2163(.din(new_new_n1759__), .dout(new_new_n3142__));
  buf1  g2164(.din(new_new_n1711__), .dout(new_new_n3143__));
  buf1  g2165(.din(new_new_n1760__), .dout(new_new_n3144__));
  buf1  g2166(.din(new_new_n3144__), .dout(new_new_n3145__));
  buf1  g2167(.din(new_new_n1712__), .dout(new_new_n3146__));
  buf1  g2168(.din(new_new_n3146__), .dout(new_new_n3147__));
  buf1  g2169(.din(new_new_n1778__), .dout(new_new_n3148__));
  buf1  g2170(.din(new_new_n1776__), .dout(new_new_n3149__));
  buf1  g2171(.din(new_new_n1774__), .dout(new_new_n3150__));
  buf1  g2172(.din(new_new_n1361__), .dout(new_new_n3151__));
  buf1  g2173(.din(new_new_n3151__), .dout(new_new_n3152__));
  buf1  g2174(.din(new_new_n945__), .dout(new_new_n3153__));
  buf1  g2175(.din(new_new_n1783__), .dout(new_new_n3154__));
  buf1  g2176(.din(new_new_n1781__), .dout(new_new_n3155__));
  buf1  g2177(.din(new_new_n1794__), .dout(new_new_n3156__));
  buf1  g2178(.din(new_new_n1789__), .dout(new_new_n3157__));
  buf1  g2179(.din(new_new_n1793__), .dout(new_new_n3158__));
  buf1  g2180(.din(new_new_n1790__), .dout(new_new_n3159__));
  buf1  g2181(.din(new_new_n1806__), .dout(new_new_n3160__));
  buf1  g2182(.din(new_new_n3160__), .dout(new_new_n3161__));
  buf1  g2183(.din(new_new_n3160__), .dout(new_new_n3162__));
  buf1  g2184(.din(new_new_n1005__), .dout(new_new_n3163__));
  buf1  g2185(.din(new_new_n1805__), .dout(new_new_n3164__));
  buf1  g2186(.din(new_new_n3164__), .dout(new_new_n3165__));
  buf1  g2187(.din(new_new_n3164__), .dout(new_new_n3166__));
  buf1  g2188(.din(new_new_n1006__), .dout(new_new_n3167__));
  buf1  g2189(.din(new_new_n1813__), .dout(new_new_n3168__));
  buf1  g2190(.din(new_new_n1803__), .dout(new_new_n3169__));
  buf1  g2191(.din(new_new_n3169__), .dout(new_new_n3170__));
  buf1  g2192(.din(new_new_n3169__), .dout(new_new_n3171__));
  buf1  g2193(.din(new_new_n1814__), .dout(new_new_n3172__));
  buf1  g2194(.din(new_new_n1804__), .dout(new_new_n3173__));
  buf1  g2195(.din(new_new_n3173__), .dout(new_new_n3174__));
  buf1  g2196(.din(new_new_n3173__), .dout(new_new_n3175__));
  buf1  g2197(.din(new_new_n1800__), .dout(new_new_n3176__));
  buf1  g2198(.din(new_new_n1799__), .dout(new_new_n3177__));
  buf1  g2199(.din(new_new_n1101__), .dout(new_new_n3178__));
  buf1  g2200(.din(new_new_n3178__), .dout(new_new_n3179__));
  buf1  g2201(.din(new_new_n3178__), .dout(new_new_n3180__));
  buf1  g2202(.din(new_new_n1040__), .dout(new_new_n3181__));
  buf1  g2203(.din(new_new_n1366__), .dout(new_new_n3182__));
  buf1  g2204(.din(new_new_n3182__), .dout(new_new_n3183__));
  buf1  g2205(.din(new_new_n1365__), .dout(new_new_n3184__));
  buf1  g2206(.din(new_new_n1475__), .dout(new_new_n3185__));
  buf1  g2207(.din(new_new_n1132__), .dout(new_new_n3186__));
  buf1  g2208(.din(new_new_n1131__), .dout(new_new_n3187__));
  buf1  g2209(.din(new_new_n3187__), .dout(new_new_n3188__));
  buf1  g2210(.din(new_new_n1037__), .dout(new_new_n3189__));
  buf1  g2211(.din(new_new_n1403__), .dout(new_new_n3190__));
  buf1  g2212(.din(new_new_n1038__), .dout(new_new_n3191__));
  buf1  g2213(.din(new_new_n1029__), .dout(new_new_n3192__));
  buf1  g2214(.din(new_new_n1848__), .dout(new_new_n3193__));
  buf1  g2215(.din(new_new_n1841__), .dout(new_new_n3194__));
  buf1  g2216(.din(new_new_n3194__), .dout(new_new_n3195__));
  buf1  g2217(.din(new_new_n1849__), .dout(new_new_n3196__));
  buf1  g2218(.din(new_new_n3196__), .dout(new_new_n3197__));
  buf1  g2219(.din(new_new_n3197__), .dout(new_new_n3198__));
  buf1  g2220(.din(new_new_n3197__), .dout(new_new_n3199__));
  buf1  g2221(.din(new_new_n3196__), .dout(new_new_n3200__));
  buf1  g2222(.din(new_new_n1842__), .dout(new_new_n3201__));
  buf1  g2223(.din(new_new_n3201__), .dout(new_new_n3202__));
  buf1  g2224(.din(new_new_n3201__), .dout(new_new_n3203__));
  buf1  g2225(.din(new_new_n1555__), .dout(new_new_n3204__));
  buf1  g2226(.din(new_new_n1553__), .dout(new_new_n3205__));
  buf1  g2227(.din(new_new_n1556__), .dout(new_new_n3206__));
  buf1  g2228(.din(new_new_n1554__), .dout(new_new_n3207__));
  buf1  g2229(.din(new_new_n1552__), .dout(new_new_n3208__));
  buf1  g2230(.din(new_new_n3208__), .dout(new_new_n3209__));
  buf1  g2231(.din(new_new_n3209__), .dout(new_new_n3210__));
  buf1  g2232(.din(new_new_n3210__), .dout(new_new_n3211__));
  buf1  g2233(.din(new_new_n3210__), .dout(new_new_n3212__));
  buf1  g2234(.din(new_new_n3209__), .dout(new_new_n3213__));
  buf1  g2235(.din(new_new_n3208__), .dout(new_new_n3214__));
  buf1  g2236(.din(new_new_n3214__), .dout(new_new_n3215__));
  buf1  g2237(.din(new_new_n3214__), .dout(new_new_n3216__));
  buf1  g2238(.din(new_new_n1551__), .dout(new_new_n3217__));
  buf1  g2239(.din(new_new_n3217__), .dout(new_new_n3218__));
  buf1  g2240(.din(new_new_n3218__), .dout(new_new_n3219__));
  buf1  g2241(.din(new_new_n3219__), .dout(new_new_n3220__));
  buf1  g2242(.din(new_new_n3219__), .dout(new_new_n3221__));
  buf1  g2243(.din(new_new_n3218__), .dout(new_new_n3222__));
  buf1  g2244(.din(new_new_n3222__), .dout(new_new_n3223__));
  buf1  g2245(.din(new_new_n3222__), .dout(new_new_n3224__));
  buf1  g2246(.din(new_new_n3217__), .dout(new_new_n3225__));
  buf1  g2247(.din(new_new_n3225__), .dout(new_new_n3226__));
  buf1  g2248(.din(new_new_n3225__), .dout(new_new_n3227__));
  buf1  g2249(.din(new_new_n1852__), .dout(new_new_n3228__));
  buf1  g2250(.din(new_new_n1534__), .dout(new_new_n3229__));
  buf1  g2251(.din(new_new_n3229__), .dout(new_new_n3230__));
  buf1  g2252(.din(new_new_n1533__), .dout(new_new_n3231__));
  buf1  g2253(.din(new_new_n1865__), .dout(new_new_n3232__));
  buf1  g2254(.din(new_new_n1863__), .dout(new_new_n3233__));
  buf1  g2255(.din(new_new_n3233__), .dout(new_new_n3234__));
  buf1  g2256(.din(new_new_n1864__), .dout(new_new_n3235__));
  buf1  g2257(.din(new_new_n1862__), .dout(new_new_n3236__));
  buf1  g2258(.din(new_new_n1536__), .dout(new_new_n3237__));
  buf1  g2259(.din(new_new_n3237__), .dout(new_new_n3238__));
  buf1  g2260(.din(new_new_n1535__), .dout(new_new_n3239__));
  buf1  g2261(.din(new_new_n1875__), .dout(new_new_n3240__));
  buf1  g2262(.din(new_new_n1873__), .dout(new_new_n3241__));
  buf1  g2263(.din(new_new_n3241__), .dout(new_new_n3242__));
  buf1  g2264(.din(new_new_n1874__), .dout(new_new_n3243__));
  buf1  g2265(.din(new_new_n1872__), .dout(new_new_n3244__));
  buf1  g2266(.din(new_new_n1143__), .dout(new_new_n3245__));
  buf1  g2267(.din(new_new_n3245__), .dout(new_new_n3246__));
  buf1  g2268(.din(new_new_n3246__), .dout(new_new_n3247__));
  buf1  g2269(.din(new_new_n3245__), .dout(new_new_n3248__));
  buf1  g2270(.din(new_new_n1144__), .dout(new_new_n3249__));
  buf1  g2271(.din(new_new_n3249__), .dout(new_new_n3250__));
  buf1  g2272(.din(new_new_n1884__), .dout(new_new_n3251__));
  buf1  g2273(.din(new_new_n3251__), .dout(new_new_n3252__));
  buf1  g2274(.din(new_new_n3252__), .dout(new_new_n3253__));
  buf1  g2275(.din(new_new_n3252__), .dout(new_new_n3254__));
  buf1  g2276(.din(new_new_n3251__), .dout(new_new_n3255__));
  buf1  g2277(.din(new_new_n1230__), .dout(new_new_n3256__));
  buf1  g2278(.din(new_new_n1882__), .dout(new_new_n3257__));
  buf1  g2279(.din(new_new_n3257__), .dout(new_new_n3258__));
  buf1  g2280(.din(new_new_n3257__), .dout(new_new_n3259__));
  buf1  g2281(.din(new_new_n1229__), .dout(new_new_n3260__));
  buf1  g2282(.din(new_new_n1490__), .dout(new_new_n3261__));
  buf1  g2283(.din(new_new_n1373__), .dout(new_new_n3262__));
  buf1  g2284(.din(new_new_n1375__), .dout(new_new_n3263__));
  buf1  g2285(.din(new_new_n1295__), .dout(new_new_n3264__));
  buf1  g2286(.din(new_new_n1870__), .dout(new_new_n3265__));
  buf1  g2287(.din(new_new_n3265__), .dout(new_new_n3266__));
  buf1  g2288(.din(new_new_n1860__), .dout(new_new_n3267__));
  buf1  g2289(.din(new_new_n3267__), .dout(new_new_n3268__));
  buf1  g2290(.din(new_new_n1220__), .dout(new_new_n3269__));
  buf1  g2291(.din(new_new_n933__), .dout(new_new_n3270__));
  buf1  g2292(.din(new_new_n3270__), .dout(new_new_n3271__));
  buf1  g2293(.din(new_new_n1901__), .dout(new_new_n3272__));
  buf1  g2294(.din(new_new_n1908__), .dout(new_new_n3273__));
  buf1  g2295(.din(new_new_n1883__), .dout(new_new_n3274__));
  buf1  g2296(.din(new_new_n1907__), .dout(new_new_n3275__));
  buf1  g2297(.din(new_new_n1909__), .dout(new_new_n3276__));
  buf1  g2298(.din(new_new_n1885__), .dout(new_new_n3277__));
  buf1  g2299(.din(new_new_n3277__), .dout(new_new_n3278__));
  buf1  g2300(.din(new_new_n3277__), .dout(new_new_n3279__));
  buf1  g2301(.din(new_new_n1910__), .dout(new_new_n3280__));
  buf1  g2302(.din(new_new_n1913__), .dout(new_new_n3281__));
  buf1  g2303(.din(new_new_n1914__), .dout(new_new_n3282__));
  buf1  g2304(.din(new_new_n1446__), .dout(new_new_n3283__));
  buf1  g2305(.din(new_new_n1445__), .dout(new_new_n3284__));
  buf1  g2306(.din(new_new_n1429__), .dout(new_new_n3285__));
  buf1  g2307(.din(new_new_n1205__), .dout(new_new_n3286__));
  buf1  g2308(.din(new_new_n3286__), .dout(new_new_n3287__));
  buf1  g2309(.din(new_new_n3286__), .dout(new_new_n3288__));
  buf1  g2310(.din(new_new_n1206__), .dout(new_new_n3289__));
  buf1  g2311(.din(new_new_n3289__), .dout(new_new_n3290__));
  buf1  g2312(.din(new_new_n3289__), .dout(new_new_n3291__));
  buf1  g2313(.din(new_new_n1839__), .dout(new_new_n3292__));
  buf1  g2314(.din(new_new_n1928__), .dout(new_new_n3293__));
  buf1  g2315(.din(new_new_n1924__), .dout(new_new_n3294__));
  buf1  g2316(.din(new_new_n3294__), .dout(new_new_n3295__));
  buf1  g2317(.din(new_new_n1927__), .dout(new_new_n3296__));
  buf1  g2318(.din(new_new_n1923__), .dout(new_new_n3297__));
  buf1  g2319(.din(new_new_n1930__), .dout(new_new_n3298__));
  buf1  g2320(.din(new_new_n1922__), .dout(new_new_n3299__));
  buf1  g2321(.din(new_new_n3299__), .dout(new_new_n3300__));
  buf1  g2322(.din(new_new_n1036__), .dout(new_new_n3301__));
  buf1  g2323(.din(new_new_n3301__), .dout(new_new_n3302__));
  buf1  g2324(.din(new_new_n3302__), .dout(new_new_n3303__));
  buf1  g2325(.din(new_new_n3302__), .dout(new_new_n3304__));
  buf1  g2326(.din(new_new_n3301__), .dout(new_new_n3305__));
  buf1  g2327(.din(new_new_n3305__), .dout(new_new_n3306__));
  buf1  g2328(.din(new_new_n1935__), .dout(new_new_n3307__));
  buf1  g2329(.din(new_new_n3307__), .dout(new_new_n3308__));
  buf1  g2330(.din(new_new_n3307__), .dout(new_new_n3309__));
  buf1  g2331(.din(new_new_n1031__), .dout(new_new_n3310__));
  buf1  g2332(.din(new_new_n1063__), .dout(new_new_n3311__));
  buf1  g2333(.din(new_new_n1939__), .dout(new_new_n3312__));
  buf1  g2334(.din(new_new_n3312__), .dout(new_new_n3313__));
  buf1  g2335(.din(new_new_n3313__), .dout(new_new_n3314__));
  buf1  g2336(.din(new_new_n3313__), .dout(new_new_n3315__));
  buf1  g2337(.din(new_new_n3312__), .dout(new_new_n3316__));
  buf1  g2338(.din(new_new_n3316__), .dout(new_new_n3317__));
  buf1  g2339(.din(new_new_n1850__), .dout(new_new_n3318__));
  buf1  g2340(.din(new_new_n3318__), .dout(new_new_n3319__));
  buf1  g2341(.din(new_new_n3319__), .dout(new_new_n3320__));
  buf1  g2342(.din(new_new_n3319__), .dout(new_new_n3321__));
  buf1  g2343(.din(new_new_n3318__), .dout(new_new_n3322__));
  buf1  g2344(.din(new_new_n3322__), .dout(new_new_n3323__));
  buf1  g2345(.din(new_new_n1951__), .dout(new_new_n3324__));
  buf1  g2346(.din(new_new_n3324__), .dout(new_new_n3325__));
  buf1  g2347(.din(new_new_n1838__), .dout(new_new_n3326__));
  buf1  g2348(.din(new_new_n3326__), .dout(new_new_n3327__));
  buf1  g2349(.din(new_new_n1950__), .dout(new_new_n3328__));
  buf1  g2350(.din(new_new_n1837__), .dout(new_new_n3329__));
  buf1  g2351(.din(new_new_n1609__), .dout(new_new_n3330__));
  buf1  g2352(.din(new_new_n3330__), .dout(new_new_n3331__));
  buf1  g2353(.din(new_new_n3331__), .dout(new_new_n3332__));
  buf1  g2354(.din(new_new_n3330__), .dout(new_new_n3333__));
  buf1  g2355(.din(new_new_n1561__), .dout(new_new_n3334__));
  buf1  g2356(.din(new_new_n3334__), .dout(new_new_n3335__));
  buf1  g2357(.din(new_new_n3334__), .dout(new_new_n3336__));
  buf1  g2358(.din(new_new_n1520__), .dout(new_new_n3337__));
  buf1  g2359(.din(new_new_n1519__), .dout(new_new_n3338__));
  buf1  g2360(.din(new_new_n1260__), .dout(new_new_n3339__));
  buf1  g2361(.din(new_new_n1981__), .dout(new_new_n3340__));
  buf1  g2362(.din(new_new_n3340__), .dout(new_new_n3341__));
  buf1  g2363(.din(new_new_n1982__), .dout(new_new_n3342__));
  buf1  g2364(.din(new_new_n3342__), .dout(new_new_n3343__));
  buf1  g2365(.din(new_new_n1257__), .dout(new_new_n3344__));
  buf1  g2366(.din(new_new_n1258__), .dout(new_new_n3345__));
  buf1  g2367(.din(new_new_n1988__), .dout(new_new_n3346__));
  buf1  g2368(.din(new_new_n1987__), .dout(new_new_n3347__));
  buf1  g2369(.din(new_new_n1478__), .dout(new_new_n3348__));
  buf1  g2370(.din(new_new_n3348__), .dout(new_new_n3349__));
  buf1  g2371(.din(new_new_n1992__), .dout(new_new_n3350__));
  buf1  g2372(.din(new_new_n1990__), .dout(new_new_n3351__));
  buf1  g2373(.din(new_new_n3351__), .dout(new_new_n3352__));
  buf1  g2374(.din(new_new_n1991__), .dout(new_new_n3353__));
  buf1  g2375(.din(new_new_n1989__), .dout(new_new_n3354__));
  buf1  g2376(.din(new_new_n1559__), .dout(new_new_n3355__));
  buf1  g2377(.din(new_new_n3355__), .dout(new_new_n3356__));
  buf1  g2378(.din(new_new_n3355__), .dout(new_new_n3357__));
  buf1  g2379(.din(new_new_n1566__), .dout(new_new_n3358__));
  buf1  g2380(.din(new_new_n1565__), .dout(new_new_n3359__));
  buf1  g2381(.din(new_new_n3359__), .dout(new_new_n3360__));
  buf1  g2382(.din(new_new_n1563__), .dout(new_new_n3361__));
  buf1  g2383(.din(new_new_n1569__), .dout(new_new_n3362__));
  buf1  g2384(.din(new_new_n1567__), .dout(new_new_n3363__));
  buf1  g2385(.din(new_new_n1920__), .dout(new_new_n3364__));
  buf1  g2386(.din(new_new_n3364__), .dout(new_new_n3365__));
  buf1  g2387(.din(new_new_n1154__), .dout(new_new_n3366__));
  buf1  g2388(.din(new_new_n1915__), .dout(new_new_n3367__));
  buf1  g2389(.din(new_new_n3367__), .dout(new_new_n3368__));
  buf1  g2390(.din(new_new_n1157__), .dout(new_new_n3369__));
  buf1  g2391(.din(new_new_n1917__), .dout(new_new_n3370__));
  buf1  g2392(.din(new_new_n1916__), .dout(new_new_n3371__));
  buf1  g2393(.din(new_new_n3371__), .dout(new_new_n3372__));
  buf1  g2394(.din(new_new_n3371__), .dout(new_new_n3373__));
  buf1  g2395(.din(new_new_n1196__), .dout(new_new_n3374__));
  buf1  g2396(.din(new_new_n1911__), .dout(new_new_n3375__));
  buf1  g2397(.din(new_new_n1197__), .dout(new_new_n3376__));
  buf1  g2398(.din(new_new_n3376__), .dout(new_new_n3377__));
  buf1  g2399(.din(new_new_n3377__), .dout(new_new_n3378__));
  buf1  g2400(.din(new_new_n3376__), .dout(new_new_n3379__));
  buf1  g2401(.din(new_new_n1289__), .dout(new_new_n3380__));
  buf1  g2402(.din(new_new_n3380__), .dout(new_new_n3381__));
  buf1  g2403(.din(new_new_n929__), .dout(new_new_n3382__));
  buf1  g2404(.din(new_new_n3382__), .dout(new_new_n3383__));
  buf1  g2405(.din(new_new_n1906__), .dout(new_new_n3384__));
  buf1  g2406(.din(new_new_n1999__), .dout(new_new_n3385__));
  buf1  g2407(.din(new_new_n1602__), .dout(new_new_n3386__));
  buf1  g2408(.din(new_new_n2012__), .dout(new_new_n3387__));
  buf1  g2409(.din(new_new_n3387__), .dout(new_new_n3388__));
  buf1  g2410(.din(new_new_n3387__), .dout(new_new_n3389__));
  buf1  g2411(.din(new_new_n1385__), .dout(new_new_n3390__));
  buf1  g2412(.din(new_new_n3390__), .dout(new_new_n3391__));
  buf1  g2413(.din(new_new_n3391__), .dout(new_new_n3392__));
  buf1  g2414(.din(new_new_n3390__), .dout(new_new_n3393__));
  buf1  g2415(.din(new_new_n2011__), .dout(new_new_n3394__));
  buf1  g2416(.din(new_new_n3394__), .dout(new_new_n3395__));
  buf1  g2417(.din(new_new_n3394__), .dout(new_new_n3396__));
  buf1  g2418(.din(new_new_n1386__), .dout(new_new_n3397__));
  buf1  g2419(.din(new_new_n3397__), .dout(new_new_n3398__));
  buf1  g2420(.din(new_new_n3397__), .dout(new_new_n3399__));
  buf1  g2421(.din(new_new_n1526__), .dout(new_new_n3400__));
  buf1  g2422(.din(new_new_n3400__), .dout(new_new_n3401__));
  buf1  g2423(.din(new_new_n3400__), .dout(new_new_n3402__));
  buf1  g2424(.din(new_new_n1525__), .dout(new_new_n3403__));
  buf1  g2425(.din(new_new_n3403__), .dout(new_new_n3404__));
  buf1  g2426(.din(new_new_n3404__), .dout(new_new_n3405__));
  buf1  g2427(.din(new_new_n3404__), .dout(new_new_n3406__));
  buf1  g2428(.din(new_new_n3403__), .dout(new_new_n3407__));
  buf1  g2429(.din(new_new_n3407__), .dout(new_new_n3408__));
  buf1  g2430(.din(new_new_n1610__), .dout(new_new_n3409__));
  buf1  g2431(.din(new_new_n3409__), .dout(new_new_n3410__));
  buf1  g2432(.din(new_new_n3409__), .dout(new_new_n3411__));
  buf1  g2433(.din(new_new_n1574__), .dout(new_new_n3412__));
  buf1  g2434(.din(new_new_n3412__), .dout(new_new_n3413__));
  buf1  g2435(.din(new_new_n3412__), .dout(new_new_n3414__));
  buf1  g2436(.din(new_new_n1573__), .dout(new_new_n3415__));
  buf1  g2437(.din(new_new_n3415__), .dout(new_new_n3416__));
  buf1  g2438(.din(new_new_n1541__), .dout(new_new_n3417__));
  buf1  g2439(.din(new_new_n3417__), .dout(new_new_n3418__));
  buf1  g2440(.din(new_new_n3418__), .dout(new_new_n3419__));
  buf1  g2441(.din(new_new_n3419__), .dout(new_new_n3420__));
  buf1  g2442(.din(new_new_n3418__), .dout(new_new_n3421__));
  buf1  g2443(.din(new_new_n3417__), .dout(new_new_n3422__));
  buf1  g2444(.din(new_new_n3422__), .dout(new_new_n3423__));
  buf1  g2445(.din(new_new_n3422__), .dout(new_new_n3424__));
  buf1  g2446(.din(new_new_n1542__), .dout(new_new_n3425__));
  buf1  g2447(.din(new_new_n3425__), .dout(new_new_n3426__));
  buf1  g2448(.din(new_new_n3426__), .dout(new_new_n3427__));
  buf1  g2449(.din(new_new_n3425__), .dout(new_new_n3428__));
  buf1  g2450(.din(new_new_n1387__), .dout(new_new_n3429__));
  buf1  g2451(.din(new_new_n3429__), .dout(new_new_n3430__));
  buf1  g2452(.din(new_new_n3429__), .dout(new_new_n3431__));
  buf1  g2453(.din(new_new_n1388__), .dout(new_new_n3432__));
  buf1  g2454(.din(new_new_n3432__), .dout(new_new_n3433__));
  buf1  g2455(.din(new_new_n3432__), .dout(new_new_n3434__));
  buf1  g2456(.din(new_new_n1611__), .dout(new_new_n3435__));
  buf1  g2457(.din(new_new_n3435__), .dout(new_new_n3436__));
  buf1  g2458(.din(new_new_n3436__), .dout(new_new_n3437__));
  buf1  g2459(.din(new_new_n3435__), .dout(new_new_n3438__));
  buf1  g2460(.din(new_new_n1576__), .dout(new_new_n3439__));
  buf1  g2461(.din(new_new_n3439__), .dout(new_new_n3440__));
  buf1  g2462(.din(new_new_n3439__), .dout(new_new_n3441__));
  buf1  g2463(.din(new_new_n1612__), .dout(new_new_n3442__));
  buf1  g2464(.din(new_new_n1562__), .dout(new_new_n3443__));
  buf1  g2465(.din(new_new_n3443__), .dout(new_new_n3444__));
  buf1  g2466(.din(new_new_n3443__), .dout(new_new_n3445__));
  buf1  g2467(.din(new_new_n1978__), .dout(new_new_n3446__));
  buf1  g2468(.din(new_new_n1379__), .dout(new_new_n3447__));
  buf1  g2469(.din(new_new_n1297__), .dout(new_new_n3448__));
  buf1  g2470(.din(new_new_n3448__), .dout(new_new_n3449__));
  buf1  g2471(.din(new_new_n3448__), .dout(new_new_n3450__));
  buf1  g2472(.din(new_new_n1592__), .dout(new_new_n3451__));
  buf1  g2473(.din(new_new_n3451__), .dout(new_new_n3452__));
  buf1  g2474(.din(new_new_n3452__), .dout(new_new_n3453__));
  buf1  g2475(.din(new_new_n3452__), .dout(new_new_n3454__));
  buf1  g2476(.din(new_new_n3451__), .dout(new_new_n3455__));
  buf1  g2477(.din(new_new_n3455__), .dout(new_new_n3456__));
  buf1  g2478(.din(new_new_n1591__), .dout(new_new_n3457__));
  buf1  g2479(.din(new_new_n3457__), .dout(new_new_n3458__));
  buf1  g2480(.din(new_new_n3458__), .dout(new_new_n3459__));
  buf1  g2481(.din(new_new_n3458__), .dout(new_new_n3460__));
  buf1  g2482(.din(new_new_n3457__), .dout(new_new_n3461__));
  buf1  g2483(.din(new_new_n3461__), .dout(new_new_n3462__));
  buf1  g2484(.din(new_new_n1497__), .dout(new_new_n3463__));
  buf1  g2485(.din(new_new_n1383__), .dout(new_new_n3464__));
  buf1  g2486(.din(new_new_n2052__), .dout(new_new_n3465__));
  buf1  g2487(.din(new_new_n3465__), .dout(new_new_n3466__));
  buf1  g2488(.din(new_new_n2048__), .dout(new_new_n3467__));
  buf1  g2489(.din(new_new_n3467__), .dout(new_new_n3468__));
  buf1  g2490(.din(new_new_n2053__), .dout(new_new_n3469__));
  buf1  g2491(.din(new_new_n3469__), .dout(new_new_n3470__));
  buf1  g2492(.din(new_new_n2049__), .dout(new_new_n3471__));
  buf1  g2493(.din(new_new_n3471__), .dout(new_new_n3472__));
  buf1  g2494(.din(new_new_n1299__), .dout(new_new_n3473__));
  buf1  g2495(.din(new_new_n3473__), .dout(new_new_n3474__));
  buf1  g2496(.din(new_new_n3474__), .dout(new_new_n3475__));
  buf1  g2497(.din(new_new_n3473__), .dout(new_new_n3476__));
  buf1  g2498(.din(new_new_n1300__), .dout(new_new_n3477__));
  buf1  g2499(.din(new_new_n2057__), .dout(new_new_n3478__));
  buf1  g2500(.din(new_new_n2056__), .dout(new_new_n3479__));
  buf1  g2501(.din(new_new_n3479__), .dout(new_new_n3480__));
  buf1  g2502(.din(new_new_n2059__), .dout(new_new_n3481__));
  buf1  g2503(.din(new_new_n1390__), .dout(new_new_n3482__));
  buf1  g2504(.din(new_new_n3482__), .dout(new_new_n3483__));
  buf1  g2505(.din(new_new_n1389__), .dout(new_new_n3484__));
  buf1  g2506(.din(new_new_n3484__), .dout(new_new_n3485__));
  buf1  g2507(.din(new_new_n1523__), .dout(new_new_n3486__));
  buf1  g2508(.din(new_new_n3486__), .dout(new_new_n3487__));
  buf1  g2509(.din(new_new_n1391__), .dout(new_new_n3488__));
  buf1  g2510(.din(new_new_n3488__), .dout(new_new_n3489__));
  buf1  g2511(.din(new_new_n3488__), .dout(new_new_n3490__));
  buf1  g2512(.din(new_new_n1524__), .dout(new_new_n3491__));
  buf1  g2513(.din(new_new_n1392__), .dout(new_new_n3492__));
  buf1  g2514(.din(new_new_n3492__), .dout(new_new_n3493__));
  buf1  g2515(.din(new_new_n2083__), .dout(new_new_n3494__));
  buf1  g2516(.din(new_new_n2000__), .dout(new_new_n3495__));
  buf1  g2517(.din(new_new_n3495__), .dout(new_new_n3496__));
  buf1  g2518(.din(new_new_n3495__), .dout(new_new_n3497__));
  buf1  g2519(.din(new_new_n1544__), .dout(new_new_n3498__));
  buf1  g2520(.din(new_new_n3498__), .dout(new_new_n3499__));
  buf1  g2521(.din(new_new_n1543__), .dout(new_new_n3500__));
  buf1  g2522(.din(new_new_n3500__), .dout(new_new_n3501__));
  buf1  g2523(.din(new_new_n2087__), .dout(new_new_n3502__));
  buf1  g2524(.din(new_new_n3502__), .dout(new_new_n3503__));
  buf1  g2525(.din(new_new_n2086__), .dout(new_new_n3504__));
  buf1  g2526(.din(new_new_n3504__), .dout(new_new_n3505__));
  buf1  g2527(.din(new_new_n2093__), .dout(new_new_n3506__));
  buf1  g2528(.din(new_new_n1192__), .dout(new_new_n3507__));
  buf1  g2529(.din(new_new_n2004__), .dout(new_new_n3508__));
  buf1  g2530(.din(new_new_n1149__), .dout(new_new_n3509__));
  buf1  g2531(.din(new_new_n3509__), .dout(new_new_n3510__));
  buf1  g2532(.din(new_new_n2099__), .dout(new_new_n3511__));
  buf1  g2533(.din(new_new_n3511__), .dout(new_new_n3512__));
  buf1  g2534(.din(new_new_n3511__), .dout(new_new_n3513__));
  buf1  g2535(.din(new_new_n1368__), .dout(new_new_n3514__));
  buf1  g2536(.din(new_new_n1195__), .dout(new_new_n3515__));
  buf1  g2537(.din(new_new_n3515__), .dout(new_new_n3516__));
  buf1  g2538(.din(new_new_n3515__), .dout(new_new_n3517__));
  buf1  g2539(.din(new_new_n1919__), .dout(new_new_n3518__));
  buf1  g2540(.din(new_new_n1367__), .dout(new_new_n3519__));
  buf1  g2541(.din(new_new_n1473__), .dout(new_new_n3520__));
  buf1  g2542(.din(new_new_n1474__), .dout(new_new_n3521__));
  buf1  g2543(.din(new_new_n2109__), .dout(new_new_n3522__));
  buf1  g2544(.din(new_new_n2105__), .dout(new_new_n3523__));
  buf1  g2545(.din(new_new_n2108__), .dout(new_new_n3524__));
  buf1  g2546(.din(new_new_n2104__), .dout(new_new_n3525__));
  buf1  g2547(.din(new_new_n3525__), .dout(new_new_n3526__));
  buf1  g2548(.din(new_new_n1424__), .dout(new_new_n3527__));
  buf1  g2549(.din(new_new_n1136__), .dout(new_new_n3528__));
  buf1  g2550(.din(new_new_n1423__), .dout(new_new_n3529__));
  buf1  g2551(.din(new_new_n1135__), .dout(new_new_n3530__));
  buf1  g2552(.din(new_new_n2123__), .dout(new_new_n3531__));
  buf1  g2553(.din(new_new_n1836__), .dout(new_new_n3532__));
  buf1  g2554(.din(new_new_n2122__), .dout(new_new_n3533__));
  buf1  g2555(.din(new_new_n1835__), .dout(new_new_n3534__));
  buf1  g2556(.din(new_new_n3534__), .dout(new_new_n3535__));
  buf1  g2557(.din(new_new_n2124__), .dout(new_new_n3536__));
  buf1  g2558(.din(new_new_n2120__), .dout(new_new_n3537__));
  buf1  g2559(.din(new_new_n3537__), .dout(new_new_n3538__));
  buf1  g2560(.din(new_new_n3537__), .dout(new_new_n3539__));
  buf1  g2561(.din(new_new_n2125__), .dout(new_new_n3540__));
  buf1  g2562(.din(new_new_n2121__), .dout(new_new_n3541__));
  buf1  g2563(.din(new_new_n3541__), .dout(new_new_n3542__));
  buf1  g2564(.din(new_new_n3542__), .dout(new_new_n3543__));
  buf1  g2565(.din(new_new_n3541__), .dout(new_new_n3544__));
  buf1  g2566(.din(new_new_n2130__), .dout(new_new_n3545__));
  buf1  g2567(.din(new_new_n2114__), .dout(new_new_n3546__));
  buf1  g2568(.din(new_new_n1237__), .dout(new_new_n3547__));
  buf1  g2569(.din(new_new_n3547__), .dout(new_new_n3548__));
  buf1  g2570(.din(new_new_n3547__), .dout(new_new_n3549__));
  buf1  g2571(.din(new_new_n2115__), .dout(new_new_n3550__));
  buf1  g2572(.din(new_new_n3550__), .dout(new_new_n3551__));
  buf1  g2573(.din(new_new_n2131__), .dout(new_new_n3552__));
  buf1  g2574(.din(new_new_n1035__), .dout(new_new_n3553__));
  buf1  g2575(.din(new_new_n3553__), .dout(new_new_n3554__));
  buf1  g2576(.din(new_new_n3554__), .dout(new_new_n3555__));
  buf1  g2577(.din(new_new_n3554__), .dout(new_new_n3556__));
  buf1  g2578(.din(new_new_n3553__), .dout(new_new_n3557__));
  buf1  g2579(.din(new_new_n3557__), .dout(new_new_n3558__));
  buf1  g2580(.din(new_new_n1046__), .dout(new_new_n3559__));
  buf1  g2581(.din(new_new_n3559__), .dout(new_new_n3560__));
  buf1  g2582(.din(new_new_n3559__), .dout(new_new_n3561__));
  buf1  g2583(.din(new_new_n1845__), .dout(new_new_n3562__));
  buf1  g2584(.din(new_new_n1833__), .dout(new_new_n3563__));
  buf1  g2585(.din(new_new_n1834__), .dout(new_new_n3564__));
  buf1  g2586(.din(new_new_n1940__), .dout(new_new_n3565__));
  buf1  g2587(.din(new_new_n1243__), .dout(new_new_n3566__));
  buf1  g2588(.din(new_new_n3566__), .dout(new_new_n3567__));
  buf1  g2589(.din(new_new_n3567__), .dout(new_new_n3568__));
  buf1  g2590(.din(new_new_n3566__), .dout(new_new_n3569__));
  buf1  g2591(.din(new_new_n1214__), .dout(new_new_n3570__));
  buf1  g2592(.din(new_new_n3570__), .dout(new_new_n3571__));
  buf1  g2593(.din(new_new_n3570__), .dout(new_new_n3572__));
  buf1  g2594(.din(new_new_n1241__), .dout(new_new_n3573__));
  buf1  g2595(.din(new_new_n3573__), .dout(new_new_n3574__));
  buf1  g2596(.din(new_new_n3573__), .dout(new_new_n3575__));
  buf1  g2597(.din(new_new_n1245__), .dout(new_new_n3576__));
  buf1  g2598(.din(new_new_n3576__), .dout(new_new_n3577__));
  buf1  g2599(.din(new_new_n1074__), .dout(new_new_n3578__));
  buf1  g2600(.din(new_new_n1211__), .dout(new_new_n3579__));
  buf1  g2601(.din(new_new_n3579__), .dout(new_new_n3580__));
  buf1  g2602(.din(new_new_n3579__), .dout(new_new_n3581__));
  buf1  g2603(.din(new_new_n1240__), .dout(new_new_n3582__));
  buf1  g2604(.din(new_new_n3582__), .dout(new_new_n3583__));
  buf1  g2605(.din(new_new_n1062__), .dout(new_new_n3584__));
  buf1  g2606(.din(new_new_n2157__), .dout(new_new_n3585__));
  buf1  g2607(.din(new_new_n1103__), .dout(new_new_n3586__));
  buf1  g2608(.din(new_new_n3586__), .dout(new_new_n3587__));
  buf1  g2609(.din(new_new_n1041__), .dout(new_new_n3588__));
  buf1  g2610(.din(new_new_n2168__), .dout(new_new_n3589__));
  buf1  g2611(.din(new_new_n1851__), .dout(new_new_n3590__));
  buf1  g2612(.din(new_new_n1045__), .dout(new_new_n3591__));
  buf1  g2613(.din(new_new_n1039__), .dout(new_new_n3592__));
  buf1  g2614(.din(new_new_n1043__), .dout(new_new_n3593__));
  buf1  g2615(.din(new_new_n1239__), .dout(new_new_n3594__));
  buf1  g2616(.din(new_new_n3594__), .dout(new_new_n3595__));
  buf1  g2617(.din(new_new_n3595__), .dout(new_new_n3596__));
  buf1  g2618(.din(new_new_n3594__), .dout(new_new_n3597__));
  buf1  g2619(.din(new_new_n1044__), .dout(new_new_n3598__));
  buf1  g2620(.din(new_new_n1212__), .dout(new_new_n3599__));
  buf1  g2621(.din(new_new_n3599__), .dout(new_new_n3600__));
  buf1  g2622(.din(new_new_n3600__), .dout(new_new_n3601__));
  buf1  g2623(.din(new_new_n3600__), .dout(new_new_n3602__));
  buf1  g2624(.din(new_new_n3599__), .dout(new_new_n3603__));
  buf1  g2625(.din(new_new_n3603__), .dout(new_new_n3604__));
  buf1  g2626(.din(new_new_n1303__), .dout(new_new_n3605__));
  buf1  g2627(.din(new_new_n1051__), .dout(new_new_n3606__));
  buf1  g2628(.din(new_new_n3606__), .dout(new_new_n3607__));
  buf1  g2629(.din(new_new_n3606__), .dout(new_new_n3608__));
  buf1  g2630(.din(new_new_n1244__), .dout(new_new_n3609__));
  buf1  g2631(.din(new_new_n3609__), .dout(new_new_n3610__));
  buf1  g2632(.din(new_new_n3610__), .dout(new_new_n3611__));
  buf1  g2633(.din(new_new_n3611__), .dout(new_new_n3612__));
  buf1  g2634(.din(new_new_n3610__), .dout(new_new_n3613__));
  buf1  g2635(.din(new_new_n3609__), .dout(new_new_n3614__));
  buf1  g2636(.din(new_new_n3614__), .dout(new_new_n3615__));
  buf1  g2637(.din(new_new_n3614__), .dout(new_new_n3616__));
  buf1  g2638(.din(new_new_n1061__), .dout(new_new_n3617__));
  buf1  g2639(.din(new_new_n3617__), .dout(new_new_n3618__));
  buf1  g2640(.din(new_new_n1042__), .dout(new_new_n3619__));
  buf1  g2641(.din(new_new_n1242__), .dout(new_new_n3620__));
  buf1  g2642(.din(new_new_n3620__), .dout(new_new_n3621__));
  buf1  g2643(.din(new_new_n3621__), .dout(new_new_n3622__));
  buf1  g2644(.din(new_new_n3621__), .dout(new_new_n3623__));
  buf1  g2645(.din(new_new_n3620__), .dout(new_new_n3624__));
  buf1  g2646(.din(new_new_n1246__), .dout(new_new_n3625__));
  buf1  g2647(.din(new_new_n3625__), .dout(new_new_n3626__));
  buf1  g2648(.din(new_new_n3626__), .dout(new_new_n3627__));
  buf1  g2649(.din(new_new_n3626__), .dout(new_new_n3628__));
  buf1  g2650(.din(new_new_n3625__), .dout(new_new_n3629__));
  buf1  g2651(.din(new_new_n3629__), .dout(new_new_n3630__));
  buf1  g2652(.din(new_new_n1213__), .dout(new_new_n3631__));
  buf1  g2653(.din(new_new_n3631__), .dout(new_new_n3632__));
  buf1  g2654(.din(new_new_n3632__), .dout(new_new_n3633__));
  buf1  g2655(.din(new_new_n3632__), .dout(new_new_n3634__));
  buf1  g2656(.din(new_new_n3631__), .dout(new_new_n3635__));
  buf1  g2657(.din(new_new_n3635__), .dout(new_new_n3636__));
  buf1  g2658(.din(new_new_n1073__), .dout(new_new_n3637__));
  buf1  g2659(.din(new_new_n1119__), .dout(new_new_n3638__));
  buf1  g2660(.din(new_new_n3638__), .dout(new_new_n3639__));
  buf1  g2661(.din(new_new_n2246__), .dout(new_new_n3640__));
  buf1  g2662(.din(new_new_n2245__), .dout(new_new_n3641__));
  buf1  g2663(.din(new_new_n1121__), .dout(new_new_n3642__));
  buf1  g2664(.din(new_new_n3642__), .dout(new_new_n3643__));
  buf1  g2665(.din(new_new_n1420__), .dout(new_new_n3644__));
  buf1  g2666(.din(new_new_n1102__), .dout(new_new_n3645__));
  buf1  g2667(.din(new_new_n1139__), .dout(new_new_n3646__));
  buf1  g2668(.din(new_new_n1140__), .dout(new_new_n3647__));
  buf1  g2669(.din(new_new_n2268__), .dout(new_new_n3648__));
  buf1  g2670(.din(new_new_n1134__), .dout(new_new_n3649__));
  buf1  g2671(.din(new_new_n2267__), .dout(new_new_n3650__));
  buf1  g2672(.din(new_new_n1133__), .dout(new_new_n3651__));
  buf1  g2673(.din(new_new_n2274__), .dout(new_new_n3652__));
  buf1  g2674(.din(new_new_n3652__), .dout(new_new_n3653__));
  buf1  g2675(.din(new_new_n2047__), .dout(new_new_n3654__));
  buf1  g2676(.din(new_new_n2281__), .dout(new_new_n3655__));
  buf1  g2677(.din(new_new_n2278__), .dout(new_new_n3656__));
  buf1  g2678(.din(new_new_n3656__), .dout(new_new_n3657__));
  buf1  g2679(.din(new_new_n2288__), .dout(new_new_n3658__));
  buf1  g2680(.din(new_new_n3658__), .dout(new_new_n3659__));
  buf1  g2681(.din(new_new_n3658__), .dout(new_new_n3660__));
  buf1  g2682(.din(new_new_n2289__), .dout(new_new_n3661__));
  buf1  g2683(.din(new_new_n2290__), .dout(new_new_n3662__));
  buf1  g2684(.din(new_new_n1238__), .dout(new_new_n3663__));
  buf1  g2685(.din(new_new_n3663__), .dout(new_new_n3664__));
  buf1  g2686(.din(new_new_n2294__), .dout(new_new_n3665__));
  buf1  g2687(.din(new_new_n1998__), .dout(new_new_n3666__));
  buf1  g2688(.din(new_new_n1881__), .dout(new_new_n3667__));
  buf1  g2689(.din(new_new_n3667__), .dout(new_new_n3668__));
  buf1  g2690(.din(new_new_n1399__), .dout(new_new_n3669__));
  buf1  g2691(.din(new_new_n1221__), .dout(new_new_n3670__));
  buf1  g2692(.din(new_new_n3670__), .dout(new_new_n3671__));
  buf1  g2693(.din(new_new_n1155__), .dout(new_new_n3672__));
  buf1  g2694(.din(new_new_n2372__), .dout(new_new_n3673__));
  buf1  g2695(.din(new_new_n2373__), .dout(new_new_n3674__));
  buf1  g2696(.din(new_new_n2273__), .dout(new_new_n3675__));
  buf1  g2697(.din(new_new_n1977__), .dout(new_new_n3676__));
  buf1  g2698(.din(new_new_n3676__), .dout(new_new_n3677__));
  buf1  g2699(.din(new_new_n1949__), .dout(new_new_n3678__));
  buf1  g2700(.din(new_new_n3678__), .dout(new_new_n3679__));
  buf1  g2701(.din(new_new_n1397__), .dout(new_new_n3680__));
  buf1  g2702(.din(new_new_n1547__), .dout(new_new_n3681__));
  buf1  g2703(.din(new_new_n2422__), .dout(new_new_n3682__));
  buf1  g2704(.din(new_new_n2082__), .dout(new_new_n3683__));
  buf1  g2705(.din(new_new_n2002__), .dout(new_new_n3684__));
  buf1  g2706(.din(new_new_n3684__), .dout(new_new_n3685__));
  buf1  g2707(.din(new_new_n3685__), .dout(new_new_n3686__));
  buf1  g2708(.din(new_new_n3685__), .dout(new_new_n3687__));
  buf1  g2709(.din(new_new_n3684__), .dout(new_new_n3688__));
  buf1  g2710(.din(new_new_n3688__), .dout(new_new_n3689__));
  buf1  g2711(.din(new_new_n2028__), .dout(new_new_n3690__));
  buf1  g2712(.din(new_new_n2085__), .dout(new_new_n3691__));
  buf1  g2713(.din(new_new_n2092__), .dout(new_new_n3692__));
  buf1  g2714(.din(new_new_n2044__), .dout(new_new_n3693__));
  buf1  g2715(.din(new_new_n2095__), .dout(new_new_n3694__));
  buf1  g2716(.din(new_new_n1147__), .dout(new_new_n3695__));
  buf1  g2717(.din(new_new_n1219__), .dout(new_new_n3696__));
  buf1  g2718(.din(new_new_n1153__), .dout(new_new_n3697__));
  buf1  g2719(.din(new_new_n1159__), .dout(new_new_n3698__));
  buf1  g2720(.din(new_new_n1887__), .dout(new_new_n3699__));
  buf1  g2721(.din(new_new_n3699__), .dout(new_new_n3700__));
  buf1  g2722(.din(new_new_n3700__), .dout(new_new_n3701__));
  buf1  g2723(.din(new_new_n3700__), .dout(new_new_n3702__));
  buf1  g2724(.din(new_new_n3699__), .dout(new_new_n3703__));
  buf1  g2725(.din(new_new_n1160__), .dout(new_new_n3704__));
  buf1  g2726(.din(new_new_n1185__), .dout(new_new_n3705__));
  buf1  g2727(.din(new_new_n1889__), .dout(new_new_n3706__));
  buf1  g2728(.din(new_new_n3706__), .dout(new_new_n3707__));
  buf1  g2729(.din(new_new_n3707__), .dout(new_new_n3708__));
  buf1  g2730(.din(new_new_n3707__), .dout(new_new_n3709__));
  buf1  g2731(.din(new_new_n3706__), .dout(new_new_n3710__));
  buf1  g2732(.din(new_new_n925__), .dout(new_new_n3711__));
  buf1  g2733(.din(new_new_n3711__), .dout(new_new_n3712__));
  buf1  g2734(.din(new_new_n2445__), .dout(new_new_n3713__));
  buf1  g2735(.din(new_new_n3713__), .dout(new_new_n3714__));
  buf1  g2736(.din(new_new_n2296__), .dout(new_new_n3715__));
  buf1  g2737(.din(new_new_n2291__), .dout(new_new_n3716__));
  buf1  g2738(.din(new_new_n3716__), .dout(new_new_n3717__));
  buf1  g2739(.din(new_new_n921__), .dout(new_new_n3718__));
  buf1  g2740(.din(new_new_n2394__), .dout(new_new_n3719__));
  buf1  g2741(.din(new_new_n992__), .dout(new_new_n3720__));
  buf1  g2742(.din(new_new_n973__), .dout(new_new_n3721__));
  buf1  g2743(.din(new_new_n969__), .dout(new_new_n3722__));
  buf1  g2744(.din(new_new_n2453__), .dout(new_new_n3723__));
  buf1  g2745(.din(new_new_n1902__), .dout(new_new_n3724__));
  buf1  g2746(.din(new_new_n991__), .dout(new_new_n3725__));
  buf1  g2747(.din(new_new_n1880__), .dout(new_new_n3726__));
  buf1  g2748(.din(new_new_n3726__), .dout(new_new_n3727__));
  buf1  g2749(.din(new_new_n2460__), .dout(new_new_n3728__));
  buf1  g2750(.din(new_new_n1997__), .dout(new_new_n3729__));
  buf1  g2751(.din(new_new_n3729__), .dout(new_new_n3730__));
  buf1  g2752(.din(new_new_n2468__), .dout(new_new_n3731__));
  buf1  g2753(.din(new_new_n2459__), .dout(new_new_n3732__));
  buf1  g2754(.din(new_new_n3732__), .dout(new_new_n3733__));
  buf1  g2755(.din(new_new_n798__), .dout(new_new_n3734__));
  buf1  g2756(.din(new_new_n795__), .dout(new_new_n3735__));
  buf1  g2757(.din(new_new_n3735__), .dout(new_new_n3736__));
  buf1  g2758(.din(new_new_n805__), .dout(new_new_n3737__));
  buf1  g2759(.din(new_new_n2007__), .dout(new_new_n3738__));
  buf1  g2760(.din(new_new_n2005__), .dout(new_new_n3739__));
  buf1  g2761(.din(new_new_n2098__), .dout(new_new_n3740__));
  buf1  g2762(.din(new_new_n1287__), .dout(new_new_n3741__));
  buf1  g2763(.din(new_new_n3741__), .dout(new_new_n3742__));
  buf1  g2764(.din(new_new_n1904__), .dout(new_new_n3743__));
  buf1  g2765(.din(new_new_n937__), .dout(new_new_n3744__));
  buf1  g2766(.din(new_new_n3744__), .dout(new_new_n3745__));
  buf1  g2767(.din(new_new_n1918__), .dout(new_new_n3746__));
  buf1  g2768(.din(new_new_n3746__), .dout(new_new_n3747__));
  buf1  g2769(.din(new_new_n3746__), .dout(new_new_n3748__));
  buf1  g2770(.din(new_new_n1169__), .dout(new_new_n3749__));
  buf1  g2771(.din(new_new_n2101__), .dout(new_new_n3750__));
  buf1  g2772(.din(new_new_n1165__), .dout(new_new_n3751__));
  buf1  g2773(.din(new_new_n3751__), .dout(new_new_n3752__));
  buf1  g2774(.din(new_new_n2356__), .dout(new_new_n3753__));
  buf1  g2775(.din(new_new_n2102__), .dout(new_new_n3754__));
  buf1  g2776(.din(new_new_n1912__), .dout(new_new_n3755__));
  buf1  g2777(.din(new_new_n3755__), .dout(new_new_n3756__));
  buf1  g2778(.din(new_new_n2389__), .dout(new_new_n3757__));
  buf1  g2779(.din(new_new_n2276__), .dout(new_new_n3758__));
  buf1  g2780(.din(new_new_n2277__), .dout(new_new_n3759__));
  buf1  g2781(.din(new_new_n1521__), .dout(new_new_n3760__));
  buf1  g2782(.din(new_new_n3760__), .dout(new_new_n3761__));
  buf1  g2783(.din(new_new_n2519__), .dout(new_new_n3762__));
  buf1  g2784(.din(new_new_n3762__), .dout(new_new_n3763__));
  buf1  g2785(.din(new_new_n3762__), .dout(new_new_n3764__));
  buf1  g2786(.din(new_new_n2009__), .dout(new_new_n3765__));
  buf1  g2787(.din(new_new_n2525__), .dout(new_new_n3766__));
  buf1  g2788(.din(new_new_n2523__), .dout(new_new_n3767__));
  buf1  g2789(.din(new_new_n2008__), .dout(new_new_n3768__));
  buf1  g2790(.din(new_new_n1599__), .dout(new_new_n3769__));
  buf1  g2791(.din(new_new_n1504__), .dout(new_new_n3770__));
  buf1  g2792(.din(new_new_n3770__), .dout(new_new_n3771__));
  buf1  g2793(.din(new_new_n1499__), .dout(new_new_n3772__));
  buf1  g2794(.din(new_new_n1503__), .dout(new_new_n3773__));
  buf1  g2795(.din(new_new_n3773__), .dout(new_new_n3774__));
  buf1  g2796(.din(new_new_n2552__), .dout(new_new_n3775__));
  buf1  g2797(.din(new_new_n2006__), .dout(new_new_n3776__));
  buf1  g2798(.din(new_new_n2003__), .dout(new_new_n3777__));
  buf1  g2799(.din(new_new_n2421__), .dout(new_new_n3778__));
  buf1  g2800(.din(new_new_n2075__), .dout(new_new_n3779__));
  buf1  g2801(.din(new_new_n2424__), .dout(new_new_n3780__));
  buf1  g2802(.din(new_new_n2430__), .dout(new_new_n3781__));
  buf1  g2803(.din(new_new_n2427__), .dout(new_new_n3782__));
  buf1  g2804(.din(new_new_n801__), .dout(new_new_n3783__));
  buf1  g2805(.din(new_new_n3783__), .dout(new_new_n3784__));
  buf1  g2806(.din(new_new_n3784__), .dout(new_new_n3785__));
  buf1  g2807(.din(new_new_n3785__), .dout(new_new_n3786__));
  buf1  g2808(.din(new_new_n3785__), .dout(new_new_n3787__));
  buf1  g2809(.din(new_new_n3784__), .dout(new_new_n3788__));
  buf1  g2810(.din(new_new_n3783__), .dout(new_new_n3789__));
  buf1  g2811(.din(new_new_n3789__), .dout(new_new_n3790__));
  buf1  g2812(.din(new_new_n3789__), .dout(new_new_n3791__));
  buf1  g2813(.din(new_new_n817__), .dout(new_new_n3792__));
  buf1  g2814(.din(new_new_n3792__), .dout(new_new_n3793__));
  buf1  g2815(.din(new_new_n3792__), .dout(new_new_n3794__));
  buf1  g2816(.din(new_new_n815__), .dout(new_new_n3795__));
  buf1  g2817(.din(new_new_n819__), .dout(new_new_n3796__));
  buf1  g2818(.din(new_new_n3796__), .dout(new_new_n3797__));
  buf1  g2819(.din(new_new_n939__), .dout(new_new_n3798__));
  buf1  g2820(.din(new_new_n2010__), .dout(new_new_n3799__));
  buf1  g2821(.din(new_new_n941__), .dout(new_new_n3800__));
  buf1  g2822(.din(new_new_n2046__), .dout(new_new_n3801__));
  buf1  g2823(.din(new_new_n1597__), .dout(new_new_n3802__));
  buf1  g2824(.din(new_new_n3802__), .dout(new_new_n3803__));
  buf1  g2825(.din(new_new_n1381__), .dout(new_new_n3804__));
  buf1  g2826(.din(new_new_n3804__), .dout(new_new_n3805__));
  buf1  g2827(.din(new_new_n3805__), .dout(new_new_n3806__));
  buf1  g2828(.din(new_new_n3804__), .dout(new_new_n3807__));
  buf1  g2829(.din(new_new_n1382__), .dout(new_new_n3808__));
  buf1  g2830(.din(new_new_n3808__), .dout(new_new_n3809__));
  buf1  g2831(.din(new_new_n3808__), .dout(new_new_n3810__));
  buf1  g2832(.din(new_new_n949__), .dout(new_new_n3811__));
  buf1  g2833(.din(new_new_n2551__), .dout(new_new_n3812__));
  buf1  g2834(.din(new_new_n1613__), .dout(new_new_n3813__));
  buf1  g2835(.din(new_new_n2054__), .dout(new_new_n3814__));
  buf1  g2836(.din(new_new_n802__), .dout(new_new_n3815__));
  buf1  g2837(.din(new_new_n3815__), .dout(new_new_n3816__));
  buf1  g2838(.din(new_new_n3816__), .dout(new_new_n3817__));
  buf1  g2839(.din(new_new_n3815__), .dout(new_new_n3818__));
  buf1  g2840(.din(new_new_n799__), .dout(new_new_n3819__));
  buf1  g2841(.din(new_new_n3819__), .dout(new_new_n3820__));
  buf1  g2842(.din(new_new_n3820__), .dout(new_new_n3821__));
  buf1  g2843(.din(new_new_n3819__), .dout(new_new_n3822__));
  buf1  g2844(.din(new_new_n2471__), .dout(new_new_n3823__));
  buf1  g2845(.din(new_new_n800__), .dout(new_new_n3824__));
  buf1  g2846(.din(new_new_n803__), .dout(new_new_n3825__));
  buf1  g2847(.din(new_new_n3825__), .dout(new_new_n3826__));
  buf1  g2848(.din(new_new_n1546__), .dout(new_new_n3827__));
  buf1  g2849(.din(new_new_n1614__), .dout(new_new_n3828__));
  buf1  g2850(.din(new_new_n2055__), .dout(new_new_n3829__));
  buf1  g2851(.din(new_new_n2623__), .dout(new_new_n3830__));
  buf1  g2852(.din(new_new_n2001__), .dout(new_new_n3831__));
  buf1  g2853(.din(new_new_n3831__), .dout(new_new_n3832__));
  buf1  g2854(.din(new_new_n2522__), .dout(new_new_n3833__));
  buf1  g2855(.din(new_new_n3833__), .dout(new_new_n3834__));
  buf1  g2856(.din(new_new_n2634__), .dout(new_new_n3835__));
  buf1  g2857(.din(new_new_n2535__), .dout(new_new_n3836__));
  buf1  g2858(.din(new_new_n3836__), .dout(new_new_n3837__));
  buf1  g2859(.din(new_new_n796__), .dout(new_new_n3838__));
  buf1  g2860(.din(new_new_n3838__), .dout(new_new_n3839__));
  buf1  g2861(.din(new_new_n2641__), .dout(new_new_n3840__));
  buf1  g2862(.din(new_new_n2472__), .dout(new_new_n3841__));
  buf1  g2863(.din(new_new_n3841__), .dout(new_new_n3842__));
  buf1  g2864(.din(new_new_n2511__), .dout(new_new_n3843__));
  buf1  g2865(.din(new_new_n2412__), .dout(new_new_n3844__));
  buf1  g2866(.din(new_new_n2554__), .dout(new_new_n3845__));
  buf1  g2867(.din(new_new_n2565__), .dout(new_new_n3846__));
  buf1  g2868(.din(new_new_n2564__), .dout(new_new_n3847__));
  buf1  g2869(.din(new_new_n820__), .dout(new_new_n3848__));
  buf1  g2870(.din(new_new_n2568__), .dout(new_new_n3849__));
  buf1  g2871(.din(new_new_n2567__), .dout(new_new_n3850__));
  buf1  g2872(.din(new_new_n2652__), .dout(new_new_n3851__));
  buf1  g2873(.din(new_new_n875__), .dout(new_new_n3852__));
  buf1  g2874(.din(new_new_n2606__), .dout(new_new_n3853__));
  buf1  g2875(.din(new_new_n3853__), .dout(new_new_n3854__));
  buf1  g2876(.din(new_new_n3853__), .dout(new_new_n3855__));
  buf1  g2877(.din(new_new_n2566__), .dout(new_new_n3856__));
  buf1  g2878(.din(new_new_n3856__), .dout(new_new_n3857__));
  buf1  g2879(.din(new_new_n3856__), .dout(new_new_n3858__));
  buf1  g2880(.din(new_new_n862__), .dout(new_new_n3859__));
  buf1  g2881(.din(new_new_n2608__), .dout(new_new_n3860__));
  buf1  g2882(.din(new_new_n2645__), .dout(new_new_n3861__));
  buf1  g2883(.din(new_new_n863__), .dout(new_new_n3862__));
  buf1  g2884(.din(new_new_n3862__), .dout(new_new_n3863__));
  buf1  g2885(.din(new_new_n2644__), .dout(new_new_n3864__));
  buf1  g2886(.din(new_new_n2607__), .dout(new_new_n3865__));
  buf1  g2887(.din(new_new_n873__), .dout(new_new_n3866__));
  buf1  g2888(.din(new_new_n859__), .dout(new_new_n3867__));
  buf1  g2889(.din(new_new_n821__), .dout(new_new_n3868__));
  buf1  g2890(.din(new_new_n861__), .dout(new_new_n3869__));
  buf1  g2891(.din(new_new_n2654__), .dout(new_new_n3870__));
  always @ (posedge clock) begin
    n1752_lo <= n6268;
    n1776_lo <= n6271;
    n1824_lo <= n6274;
    n1836_lo <= n6277;
    n1848_lo <= n6280;
    n1860_lo <= n6283;
    n1872_lo <= n6286;
    n1884_lo <= n6289;
    n1896_lo <= n6292;
    n1908_lo <= n6295;
    n1911_lo <= n6298;
    n1914_lo <= n6301;
    n1923_lo <= n6304;
    n1926_lo <= n6307;
    n1935_lo <= n6310;
    n1938_lo <= n6313;
    n1947_lo <= n6316;
    n1950_lo <= n6319;
    n1959_lo <= n6322;
    n1962_lo <= n6325;
    n1971_lo <= n6328;
    n1974_lo <= n6331;
    n1983_lo <= n6334;
    n1995_lo <= n6337;
    n2055_lo <= n6340;
    n2064_lo <= n6343;
    n2067_lo <= n6346;
    n2079_lo <= n6349;
    n2100_lo <= n6352;
    n2112_lo <= n6355;
    n2124_lo <= n6358;
    n2136_lo <= n6361;
    n2148_lo <= n6364;
    n2160_lo <= n6367;
    n2172_lo <= n6370;
    n2184_lo <= n6373;
    n2235_lo <= n6376;
    n2238_lo <= n6379;
    n2247_lo <= n6382;
    n2250_lo <= n6385;
    n2259_lo <= n6388;
    n2262_lo <= n6391;
    n2271_lo <= n6394;
    n2274_lo <= n6397;
    n2283_lo <= n6400;
    n2286_lo <= n6403;
    n2289_lo <= n6406;
    n2295_lo <= n6409;
    n2298_lo <= n6412;
    n2304_lo <= n6415;
    n2307_lo <= n6418;
    n2316_lo <= n6421;
    n2331_lo <= n6424;
    n2334_lo <= n6427;
    n2337_lo <= n6430;
    n2340_lo <= n6433;
    n2071_o2 <= n6436;
    n2080_o2 <= n6439;
    n2137_o2 <= n6442;
    n2368_o2 <= n6445;
    n2383_o2 <= n6448;
    n2405_o2 <= n6451;
    n2471_o2 <= n6454;
    n2617_o2 <= n6457;
    n2765_o2 <= n6460;
    n2775_o2 <= n6463;
    n2829_o2 <= n6466;
    n2579_o2 <= n6469;
    n2580_o2 <= n6472;
    n2618_o2 <= n6475;
    n2619_o2 <= n6478;
    n2620_o2 <= n6481;
    n2621_o2 <= n6484;
    n2622_o2 <= n6487;
    n2623_o2 <= n6490;
    n2624_o2 <= n6493;
    n2625_o2 <= n6496;
    n2626_o2 <= n6499;
    n2627_o2 <= n6502;
    n3029_o2 <= n6505;
    n3035_o2 <= n6508;
    n2643_o2 <= n6511;
    n2644_o2 <= n6514;
    n2645_o2 <= n6517;
    n327_inv <= n6520;
    n2658_o2 <= n6523;
    n2659_o2 <= n6526;
    n2674_o2 <= n6529;
    n2675_o2 <= n6532;
    n2676_o2 <= n6535;
    n3119_o2 <= n6538;
    n3153_o2 <= n6541;
    n351_inv <= n6544;
    n2729_o2 <= n6547;
    n2730_o2 <= n6550;
    n2731_o2 <= n6553;
    n698_o2 <= n6556;
    n366_inv <= n6559;
    n2757_o2 <= n6562;
    n2758_o2 <= n6565;
    n1000_o2 <= n6568;
    n1160_o2 <= n6571;
    n1153_o2 <= n6574;
    n2793_o2 <= n6577;
    n2794_o2 <= n6580;
    n2795_o2 <= n6583;
    n1001_o2 <= n6586;
    n2859_o2 <= n6589;
    n744_o2 <= n6592;
    n402_inv <= n6595;
    n2926_o2 <= n6598;
    n408_inv <= n6601;
    n2966_o2 <= n6604;
    n2967_o2 <= n6607;
    n2947_o2 <= n6610;
    n1010_o2 <= n6613;
    n2976_o2 <= n6616;
    n3069_o2 <= n6619;
    n3028_o2 <= n6622;
    n3081_o2 <= n6625;
    n3082_o2 <= n6628;
    n3142_o2 <= n6631;
    n3214_o2 <= n6634;
    n2992_o2 <= n6637;
    n2993_o2 <= n6640;
    n870_o2 <= n6643;
    n3086_o2 <= n6646;
    n3087_o2 <= n6649;
    n3088_o2 <= n6652;
    n3089_o2 <= n6655;
    n3090_o2 <= n6658;
    n3091_o2 <= n6661;
    n3092_o2 <= n6664;
    n3093_o2 <= n6667;
    n3094_o2 <= n6670;
    n3095_o2 <= n6673;
    n483_inv <= n6676;
    n3170_o2 <= n6679;
    n3171_o2 <= n6682;
    n3172_o2 <= n6685;
    n3179_o2 <= n6688;
    n498_inv <= n6691;
    n3193_o2 <= n6694;
    n3211_o2 <= n6697;
    n3212_o2 <= n6700;
    n3213_o2 <= n6703;
    n513_inv <= n6706;
    n1125_o2 <= n6709;
    n1081_o2 <= n6712;
    n1139_o2 <= n6715;
    n3245_o2 <= n6718;
    n3246_o2 <= n6721;
    n3247_o2 <= n6724;
    lo074_buf_o2 <= n6727;
    lo078_buf_o2 <= n6730;
    lo186_buf_o2 <= n6733;
    lo118_buf_o2 <= n6736;
    lo146_buf_o2 <= n6739;
    n1038_o2 <= n6742;
    n1044_o2 <= n6745;
    n555_inv <= n6748;
    n558_inv <= n6751;
    lo026_buf_o2 <= n6754;
    lo030_buf_o2 <= n6757;
    lo090_buf_o2 <= n6760;
    lo094_buf_o2 <= n6763;
    lo098_buf_o2 <= n6766;
    lo102_buf_o2 <= n6769;
    lo066_buf_o2 <= n6772;
    lo070_buf_o2 <= n6775;
    n1202_o2 <= n6778;
    n1003_o2 <= n6781;
    n1031_o2 <= n6784;
    n1034_o2 <= n6787;
    n1040_o2 <= n6790;
    n1046_o2 <= n6793;
    n1380_o2 <= n6796;
    n1425_o2 <= n6799;
    n697_o2 <= n6802;
    n1143_o2 <= n6805;
    n673_o2 <= n6808;
    n789_o2 <= n6811;
    n786_o2 <= n6814;
    n1047_o2 <= n6817;
    n1036_o2 <= n6820;
    n1307_o2 <= n6823;
    n1035_o2 <= n6826;
    n1297_o2 <= n6829;
    n1099_o2 <= n6832;
    n1128_o2 <= n6835;
    n645_inv <= n6838;
    n826_o2 <= n6841;
    n853_o2 <= n6844;
    n654_inv <= n6847;
    n700_o2 <= n6850;
    n884_o2 <= n6853;
    lo082_buf_o2 <= n6856;
    lo086_buf_o2 <= n6859;
    n801_o2 <= n6862;
    n840_o2 <= n6865;
    n675_inv <= n6868;
    lo002_buf_o2 <= n6871;
    lo010_buf_o2 <= n6874;
    lo166_buf_o2 <= n6877;
    lo170_buf_o2 <= n6880;
    n1426_o2 <= n6883;
    n1082_o2 <= n6886;
    n1310_o2 <= n6889;
    n1015_o2 <= n6892;
    n1206_o2 <= n6895;
    n1262_o2 <= n6898;
    n1456_o2 <= n6901;
    n1244_o2 <= n6904;
    n1280_o2 <= n6907;
    n1290_o2 <= n6910;
    n1012_o2 <= n6913;
    n1074_o2 <= n6916;
    n1112_o2 <= n6919;
    n1212_o2 <= n6922;
    n1454_o2 <= n6925;
    n1182_o2 <= n6928;
    n1220_o2 <= n6931;
    n701_o2 <= n6934;
    n744_inv <= n6937;
    n1282_o2 <= n6940;
    n1144_o2 <= n6943;
    n1278_o2 <= n6946;
    n1459_o2 <= n6949;
    n1324_o2 <= n6952;
    n1288_o2 <= n6955;
    n1271_o2 <= n6958;
    n1132_o2 <= n6961;
    n1231_o2 <= n6964;
    n1462_o2 <= n6967;
    n1482_o2 <= n6970;
    n994_o2 <= n6973;
    n998_o2 <= n6976;
    lo106_buf_o2 <= n6979;
    n769_o2 <= n6982;
    n814_o2 <= n6985;
    n841_o2 <= n6988;
    n867_o2 <= n6991;
    lo006_buf_o2 <= n6994;
    lo014_buf_o2 <= n6997;
    lo022_buf_o2 <= n7000;
    lo042_buf_o2 <= n7003;
    lo046_buf_o2 <= n7006;
    lo050_buf_o2 <= n7009;
    lo054_buf_o2 <= n7012;
    lo130_buf_o2 <= n7015;
    lo134_buf_o2 <= n7018;
    lo154_buf_o2 <= n7021;
    lo174_buf_o2 <= n7024;
    lo178_buf_o2 <= n7027;
    n1007_o2 <= n7030;
    n1294_o2 <= n7033;
    n1084_o2 <= n7036;
    n1399_o2 <= n7039;
    n1311_o2 <= n7042;
    n1392_o2 <= n7045;
    n1102_o2 <= n7048;
    n1041_o2 <= n7051;
    n1298_o2 <= n7054;
    n738_o2 <= n7057;
    n1214_o2 <= n7060;
    n1222_o2 <= n7063;
    n1155_o2 <= n7066;
    n1147_o2 <= n7069;
    n1393_o2 <= n7072;
    n999_o2 <= n7075;
    n1306_o2 <= n7078;
    n1312_o2 <= n7081;
    n1382_o2 <= n7084;
    n1383_o2 <= n7087;
    n1152_o2 <= n7090;
    n1334_o2 <= n7093;
    n1335_o2 <= n7096;
    n906_inv <= n7099;
    n773_o2 <= n7102;
    lo190_buf_o2 <= n7105;
    n1368_o2 <= n7108;
    n1362_o2 <= n7111;
    n1406_o2 <= n7114;
    n1403_o2 <= n7117;
    n741_o2 <= n7120;
    n1407_o2 <= n7123;
    n1395_o2 <= n7126;
    n1359_o2 <= n7129;
    n1159_o2 <= n7132;
    n1221_o2 <= n7135;
    n945_inv <= n7138;
    n989_o2 <= n7141;
    n881_o2 <= n7144;
    n1340_o2 <= n7147;
    n1341_o2 <= n7150;
    n906_o2 <= n7153;
    n1388_o2 <= n7156;
    n791_o2 <= n7159;
    n1372_o2 <= n7162;
    n815_o2 <= n7165;
    n868_o2 <= n7168;
    lo018_buf_o2 <= n7171;
    lo138_buf_o2 <= n7174;
    lo158_buf_o2 <= n7177;
    n780_o2 <= n7180;
    n728_o2 <= n7183;
    n993_inv <= n7186;
    n929_o2 <= n7189;
    n955_o2 <= n7192;
    n938_o2 <= n7195;
    n1117_o2 <= n7198;
    n1121_o2 <= n7201;
    n965_o2 <= n7204;
    n752_o2 <= n7207;
    n753_o2 <= n7210;
    n760_o2 <= n7213;
    n770_o2 <= n7216;
    n923_o2 <= n7219;
    n947_o2 <= n7222;
    n897_o2 <= n7225;
    n919_o2 <= n7228;
    n895_o2 <= n7231;
    n917_o2 <= n7234;
    n751_o2 <= n7237;
    n774_o2 <= n7240;
    lo126_buf_o2 <= n7243;
    lo142_buf_o2 <= n7246;
    lo162_buf_o2 <= n7249;
    n1059_inv <= n7252;
    n792_o2 <= n7255;
    n869_o2 <= n7258;
    n1068_inv <= n7261;
    lo024_buf_o2 <= n7264;
    lo028_buf_o2 <= n7267;
    lo088_buf_o2 <= n7270;
    lo092_buf_o2 <= n7273;
    lo096_buf_o2 <= n7276;
    lo100_buf_o2 <= n7279;
    n763_o2 <= n7282;
    n754_o2 <= n7285;
    n755_o2 <= n7288;
    n822_o2 <= n7291;
    n849_o2 <= n7294;
    n777_o2 <= n7297;
    n778_o2 <= n7300;
    n820_o2 <= n7303;
    n846_o2 <= n7306;
    n806_o2 <= n7309;
    n771_o2 <= n7312;
    n854_o2 <= n7315;
    n828_o2 <= n7318;
    lo117_buf_o2 <= n7321;
    lo145_buf_o2 <= n7324;
    n762_o2 <= n7327;
    n805_o2 <= n7330;
    n859_o2 <= n7333;
    n833_o2 <= n7336;
    lo034_buf_o2 <= n7339;
    lo038_buf_o2 <= n7342;
    lo122_buf_o2 <= n7345;
    lo150_buf_o2 <= n7348;
  end
  initial begin
    n1752_lo <= 1'b0;
    n1776_lo <= 1'b0;
    n1824_lo <= 1'b0;
    n1836_lo <= 1'b0;
    n1848_lo <= 1'b0;
    n1860_lo <= 1'b0;
    n1872_lo <= 1'b0;
    n1884_lo <= 1'b0;
    n1896_lo <= 1'b0;
    n1908_lo <= 1'b0;
    n1911_lo <= 1'b0;
    n1914_lo <= 1'b0;
    n1923_lo <= 1'b0;
    n1926_lo <= 1'b0;
    n1935_lo <= 1'b0;
    n1938_lo <= 1'b0;
    n1947_lo <= 1'b0;
    n1950_lo <= 1'b0;
    n1959_lo <= 1'b0;
    n1962_lo <= 1'b0;
    n1971_lo <= 1'b0;
    n1974_lo <= 1'b0;
    n1983_lo <= 1'b0;
    n1995_lo <= 1'b0;
    n2055_lo <= 1'b0;
    n2064_lo <= 1'b0;
    n2067_lo <= 1'b0;
    n2079_lo <= 1'b0;
    n2100_lo <= 1'b0;
    n2112_lo <= 1'b0;
    n2124_lo <= 1'b0;
    n2136_lo <= 1'b0;
    n2148_lo <= 1'b0;
    n2160_lo <= 1'b0;
    n2172_lo <= 1'b0;
    n2184_lo <= 1'b0;
    n2235_lo <= 1'b0;
    n2238_lo <= 1'b0;
    n2247_lo <= 1'b0;
    n2250_lo <= 1'b0;
    n2259_lo <= 1'b0;
    n2262_lo <= 1'b0;
    n2271_lo <= 1'b0;
    n2274_lo <= 1'b0;
    n2283_lo <= 1'b0;
    n2286_lo <= 1'b0;
    n2289_lo <= 1'b0;
    n2295_lo <= 1'b0;
    n2298_lo <= 1'b0;
    n2304_lo <= 1'b0;
    n2307_lo <= 1'b0;
    n2316_lo <= 1'b0;
    n2331_lo <= 1'b0;
    n2334_lo <= 1'b0;
    n2337_lo <= 1'b0;
    n2340_lo <= 1'b0;
    n2071_o2 <= 1'b0;
    n2080_o2 <= 1'b0;
    n2137_o2 <= 1'b0;
    n2368_o2 <= 1'b0;
    n2383_o2 <= 1'b0;
    n2405_o2 <= 1'b0;
    n2471_o2 <= 1'b0;
    n2617_o2 <= 1'b0;
    n2765_o2 <= 1'b0;
    n2775_o2 <= 1'b0;
    n2829_o2 <= 1'b0;
    n2579_o2 <= 1'b0;
    n2580_o2 <= 1'b0;
    n2618_o2 <= 1'b0;
    n2619_o2 <= 1'b0;
    n2620_o2 <= 1'b0;
    n2621_o2 <= 1'b0;
    n2622_o2 <= 1'b0;
    n2623_o2 <= 1'b0;
    n2624_o2 <= 1'b0;
    n2625_o2 <= 1'b0;
    n2626_o2 <= 1'b0;
    n2627_o2 <= 1'b0;
    n3029_o2 <= 1'b0;
    n3035_o2 <= 1'b0;
    n2643_o2 <= 1'b0;
    n2644_o2 <= 1'b0;
    n2645_o2 <= 1'b0;
    n327_inv <= 1'b0;
    n2658_o2 <= 1'b0;
    n2659_o2 <= 1'b0;
    n2674_o2 <= 1'b0;
    n2675_o2 <= 1'b0;
    n2676_o2 <= 1'b0;
    n3119_o2 <= 1'b0;
    n3153_o2 <= 1'b0;
    n351_inv <= 1'b0;
    n2729_o2 <= 1'b0;
    n2730_o2 <= 1'b0;
    n2731_o2 <= 1'b0;
    n698_o2 <= 1'b0;
    n366_inv <= 1'b0;
    n2757_o2 <= 1'b0;
    n2758_o2 <= 1'b0;
    n1000_o2 <= 1'b0;
    n1160_o2 <= 1'b0;
    n1153_o2 <= 1'b0;
    n2793_o2 <= 1'b0;
    n2794_o2 <= 1'b0;
    n2795_o2 <= 1'b0;
    n1001_o2 <= 1'b0;
    n2859_o2 <= 1'b0;
    n744_o2 <= 1'b0;
    n402_inv <= 1'b0;
    n2926_o2 <= 1'b0;
    n408_inv <= 1'b0;
    n2966_o2 <= 1'b0;
    n2967_o2 <= 1'b0;
    n2947_o2 <= 1'b0;
    n1010_o2 <= 1'b0;
    n2976_o2 <= 1'b0;
    n3069_o2 <= 1'b0;
    n3028_o2 <= 1'b0;
    n3081_o2 <= 1'b0;
    n3082_o2 <= 1'b0;
    n3142_o2 <= 1'b0;
    n3214_o2 <= 1'b0;
    n2992_o2 <= 1'b0;
    n2993_o2 <= 1'b0;
    n870_o2 <= 1'b0;
    n3086_o2 <= 1'b0;
    n3087_o2 <= 1'b0;
    n3088_o2 <= 1'b0;
    n3089_o2 <= 1'b0;
    n3090_o2 <= 1'b0;
    n3091_o2 <= 1'b0;
    n3092_o2 <= 1'b0;
    n3093_o2 <= 1'b0;
    n3094_o2 <= 1'b0;
    n3095_o2 <= 1'b0;
    n483_inv <= 1'b0;
    n3170_o2 <= 1'b0;
    n3171_o2 <= 1'b0;
    n3172_o2 <= 1'b0;
    n3179_o2 <= 1'b0;
    n498_inv <= 1'b0;
    n3193_o2 <= 1'b0;
    n3211_o2 <= 1'b0;
    n3212_o2 <= 1'b0;
    n3213_o2 <= 1'b0;
    n513_inv <= 1'b0;
    n1125_o2 <= 1'b0;
    n1081_o2 <= 1'b0;
    n1139_o2 <= 1'b0;
    n3245_o2 <= 1'b0;
    n3246_o2 <= 1'b0;
    n3247_o2 <= 1'b0;
    lo074_buf_o2 <= 1'b0;
    lo078_buf_o2 <= 1'b0;
    lo186_buf_o2 <= 1'b0;
    lo118_buf_o2 <= 1'b0;
    lo146_buf_o2 <= 1'b0;
    n1038_o2 <= 1'b0;
    n1044_o2 <= 1'b0;
    n555_inv <= 1'b0;
    n558_inv <= 1'b0;
    lo026_buf_o2 <= 1'b0;
    lo030_buf_o2 <= 1'b0;
    lo090_buf_o2 <= 1'b0;
    lo094_buf_o2 <= 1'b0;
    lo098_buf_o2 <= 1'b0;
    lo102_buf_o2 <= 1'b0;
    lo066_buf_o2 <= 1'b0;
    lo070_buf_o2 <= 1'b0;
    n1202_o2 <= 1'b0;
    n1003_o2 <= 1'b0;
    n1031_o2 <= 1'b0;
    n1034_o2 <= 1'b0;
    n1040_o2 <= 1'b0;
    n1046_o2 <= 1'b0;
    n1380_o2 <= 1'b0;
    n1425_o2 <= 1'b0;
    n697_o2 <= 1'b0;
    n1143_o2 <= 1'b0;
    n673_o2 <= 1'b0;
    n789_o2 <= 1'b0;
    n786_o2 <= 1'b0;
    n1047_o2 <= 1'b0;
    n1036_o2 <= 1'b0;
    n1307_o2 <= 1'b0;
    n1035_o2 <= 1'b0;
    n1297_o2 <= 1'b0;
    n1099_o2 <= 1'b0;
    n1128_o2 <= 1'b0;
    n645_inv <= 1'b0;
    n826_o2 <= 1'b0;
    n853_o2 <= 1'b0;
    n654_inv <= 1'b0;
    n700_o2 <= 1'b0;
    n884_o2 <= 1'b0;
    lo082_buf_o2 <= 1'b0;
    lo086_buf_o2 <= 1'b0;
    n801_o2 <= 1'b0;
    n840_o2 <= 1'b0;
    n675_inv <= 1'b0;
    lo002_buf_o2 <= 1'b0;
    lo010_buf_o2 <= 1'b0;
    lo166_buf_o2 <= 1'b0;
    lo170_buf_o2 <= 1'b0;
    n1426_o2 <= 1'b0;
    n1082_o2 <= 1'b0;
    n1310_o2 <= 1'b0;
    n1015_o2 <= 1'b0;
    n1206_o2 <= 1'b0;
    n1262_o2 <= 1'b0;
    n1456_o2 <= 1'b0;
    n1244_o2 <= 1'b0;
    n1280_o2 <= 1'b0;
    n1290_o2 <= 1'b0;
    n1012_o2 <= 1'b0;
    n1074_o2 <= 1'b0;
    n1112_o2 <= 1'b0;
    n1212_o2 <= 1'b0;
    n1454_o2 <= 1'b0;
    n1182_o2 <= 1'b0;
    n1220_o2 <= 1'b0;
    n701_o2 <= 1'b0;
    n744_inv <= 1'b0;
    n1282_o2 <= 1'b0;
    n1144_o2 <= 1'b0;
    n1278_o2 <= 1'b0;
    n1459_o2 <= 1'b0;
    n1324_o2 <= 1'b0;
    n1288_o2 <= 1'b0;
    n1271_o2 <= 1'b0;
    n1132_o2 <= 1'b0;
    n1231_o2 <= 1'b0;
    n1462_o2 <= 1'b0;
    n1482_o2 <= 1'b0;
    n994_o2 <= 1'b0;
    n998_o2 <= 1'b0;
    lo106_buf_o2 <= 1'b0;
    n769_o2 <= 1'b0;
    n814_o2 <= 1'b0;
    n841_o2 <= 1'b0;
    n867_o2 <= 1'b0;
    lo006_buf_o2 <= 1'b0;
    lo014_buf_o2 <= 1'b0;
    lo022_buf_o2 <= 1'b0;
    lo042_buf_o2 <= 1'b0;
    lo046_buf_o2 <= 1'b0;
    lo050_buf_o2 <= 1'b0;
    lo054_buf_o2 <= 1'b0;
    lo130_buf_o2 <= 1'b0;
    lo134_buf_o2 <= 1'b0;
    lo154_buf_o2 <= 1'b0;
    lo174_buf_o2 <= 1'b0;
    lo178_buf_o2 <= 1'b0;
    n1007_o2 <= 1'b0;
    n1294_o2 <= 1'b0;
    n1084_o2 <= 1'b0;
    n1399_o2 <= 1'b0;
    n1311_o2 <= 1'b0;
    n1392_o2 <= 1'b0;
    n1102_o2 <= 1'b0;
    n1041_o2 <= 1'b0;
    n1298_o2 <= 1'b0;
    n738_o2 <= 1'b0;
    n1214_o2 <= 1'b0;
    n1222_o2 <= 1'b0;
    n1155_o2 <= 1'b0;
    n1147_o2 <= 1'b0;
    n1393_o2 <= 1'b0;
    n999_o2 <= 1'b0;
    n1306_o2 <= 1'b0;
    n1312_o2 <= 1'b0;
    n1382_o2 <= 1'b0;
    n1383_o2 <= 1'b0;
    n1152_o2 <= 1'b0;
    n1334_o2 <= 1'b0;
    n1335_o2 <= 1'b0;
    n906_inv <= 1'b0;
    n773_o2 <= 1'b0;
    lo190_buf_o2 <= 1'b0;
    n1368_o2 <= 1'b0;
    n1362_o2 <= 1'b0;
    n1406_o2 <= 1'b0;
    n1403_o2 <= 1'b0;
    n741_o2 <= 1'b0;
    n1407_o2 <= 1'b0;
    n1395_o2 <= 1'b0;
    n1359_o2 <= 1'b0;
    n1159_o2 <= 1'b0;
    n1221_o2 <= 1'b0;
    n945_inv <= 1'b0;
    n989_o2 <= 1'b0;
    n881_o2 <= 1'b0;
    n1340_o2 <= 1'b0;
    n1341_o2 <= 1'b0;
    n906_o2 <= 1'b0;
    n1388_o2 <= 1'b0;
    n791_o2 <= 1'b0;
    n1372_o2 <= 1'b0;
    n815_o2 <= 1'b0;
    n868_o2 <= 1'b0;
    lo018_buf_o2 <= 1'b0;
    lo138_buf_o2 <= 1'b0;
    lo158_buf_o2 <= 1'b0;
    n780_o2 <= 1'b0;
    n728_o2 <= 1'b0;
    n993_inv <= 1'b0;
    n929_o2 <= 1'b0;
    n955_o2 <= 1'b0;
    n938_o2 <= 1'b0;
    n1117_o2 <= 1'b0;
    n1121_o2 <= 1'b0;
    n965_o2 <= 1'b0;
    n752_o2 <= 1'b0;
    n753_o2 <= 1'b0;
    n760_o2 <= 1'b0;
    n770_o2 <= 1'b0;
    n923_o2 <= 1'b0;
    n947_o2 <= 1'b0;
    n897_o2 <= 1'b0;
    n919_o2 <= 1'b0;
    n895_o2 <= 1'b0;
    n917_o2 <= 1'b0;
    n751_o2 <= 1'b0;
    n774_o2 <= 1'b0;
    lo126_buf_o2 <= 1'b0;
    lo142_buf_o2 <= 1'b0;
    lo162_buf_o2 <= 1'b0;
    n1059_inv <= 1'b0;
    n792_o2 <= 1'b0;
    n869_o2 <= 1'b0;
    n1068_inv <= 1'b0;
    lo024_buf_o2 <= 1'b0;
    lo028_buf_o2 <= 1'b0;
    lo088_buf_o2 <= 1'b0;
    lo092_buf_o2 <= 1'b0;
    lo096_buf_o2 <= 1'b0;
    lo100_buf_o2 <= 1'b0;
    n763_o2 <= 1'b0;
    n754_o2 <= 1'b0;
    n755_o2 <= 1'b0;
    n822_o2 <= 1'b0;
    n849_o2 <= 1'b0;
    n777_o2 <= 1'b0;
    n778_o2 <= 1'b0;
    n820_o2 <= 1'b0;
    n846_o2 <= 1'b0;
    n806_o2 <= 1'b0;
    n771_o2 <= 1'b0;
    n854_o2 <= 1'b0;
    n828_o2 <= 1'b0;
    lo117_buf_o2 <= 1'b0;
    lo145_buf_o2 <= 1'b0;
    n762_o2 <= 1'b0;
    n805_o2 <= 1'b0;
    n859_o2 <= 1'b0;
    n833_o2 <= 1'b0;
    lo034_buf_o2 <= 1'b0;
    lo038_buf_o2 <= 1'b0;
    lo122_buf_o2 <= 1'b0;
    lo150_buf_o2 <= 1'b0;
  end
endmodule


