
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G1884,
  G1885,
  G1886,
  G1887,
  G1888,
  G1889,
  G1890,
  G1891,
  G1892,
  G1893,
  G1894,
  G1895,
  G1896,
  G1897,
  G1898,
  G1899,
  G1900,
  G1901,
  G1902,
  G1903,
  G1904,
  G1905,
  G1906,
  G1907,
  G1908
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;
  output G1884;output G1885;output G1886;output G1887;output G1888;output G1889;output G1890;output G1891;output G1892;output G1893;output G1894;output G1895;output G1896;output G1897;output G1898;output G1899;output G1900;output G1901;output G1902;output G1903;output G1904;output G1905;output G1906;output G1907;output G1908;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire g34_p;
  wire g34_n;
  wire g35_p;
  wire g35_n;
  wire g36_p;
  wire g36_n;
  wire g37_p;
  wire g37_n;
  wire g38_p;
  wire g38_n;
  wire g39_p;
  wire g39_n;
  wire g40_p;
  wire g40_n;
  wire g41_p;
  wire g41_n;
  wire g42_p;
  wire g42_n;
  wire g43_p;
  wire g43_n;
  wire g44_p;
  wire g44_n;
  wire g45_p;
  wire g45_n;
  wire g46_p;
  wire g46_n;
  wire g47_p;
  wire g47_n;
  wire g48_p;
  wire g48_n;
  wire g49_p;
  wire g49_n;
  wire g50_p;
  wire g50_n;
  wire g51_p;
  wire g51_n;
  wire g52_p;
  wire g52_n;
  wire g53_p;
  wire g53_n;
  wire g54_p;
  wire g54_n;
  wire g55_p;
  wire g55_n;
  wire g56_p;
  wire g56_n;
  wire g57_p;
  wire g57_n;
  wire g58_p;
  wire g58_n;
  wire g59_p;
  wire g59_n;
  wire g60_p;
  wire g60_n;
  wire g61_p;
  wire g61_n;
  wire g62_p;
  wire g62_n;
  wire g63_p;
  wire g63_n;
  wire g64_p;
  wire g64_n;
  wire g65_p;
  wire g65_n;
  wire g66_p;
  wire g66_n;
  wire g67_p;
  wire g67_n;
  wire g68_p;
  wire g68_n;
  wire g69_p;
  wire g69_n;
  wire g70_p;
  wire g70_n;
  wire g71_p;
  wire g71_n;
  wire g72_p;
  wire g72_n;
  wire g73_p;
  wire g73_n;
  wire g74_p;
  wire g74_n;
  wire g75_p;
  wire g75_n;
  wire g76_p;
  wire g76_n;
  wire g77_p;
  wire g77_n;
  wire g78_p;
  wire g78_n;
  wire g79_p;
  wire g79_n;
  wire g80_p;
  wire g80_n;
  wire g81_p;
  wire g81_n;
  wire g82_p;
  wire g82_n;
  wire g83_p;
  wire g83_n;
  wire g84_p;
  wire g84_n;
  wire g85_p;
  wire g85_n;
  wire g86_p;
  wire g86_n;
  wire g87_p;
  wire g87_n;
  wire g88_p;
  wire g88_n;
  wire g89_p;
  wire g89_n;
  wire g90_p;
  wire g90_n;
  wire g91_p;
  wire g91_n;
  wire g92_p;
  wire g92_n;
  wire g93_p;
  wire g93_n;
  wire g94_p;
  wire g94_n;
  wire g95_p;
  wire g95_n;
  wire g96_p;
  wire g96_n;
  wire g97_p;
  wire g97_n;
  wire g98_p;
  wire g98_n;
  wire g99_p;
  wire g99_n;
  wire g100_p;
  wire g100_n;
  wire g101_p;
  wire g101_n;
  wire g102_p;
  wire g102_n;
  wire g103_p;
  wire g103_n;
  wire g104_p;
  wire g104_n;
  wire g105_p;
  wire g105_n;
  wire g106_p;
  wire g106_n;
  wire g107_p;
  wire g107_n;
  wire g108_p;
  wire g108_n;
  wire g109_p;
  wire g109_n;
  wire g110_p;
  wire g110_n;
  wire g111_p;
  wire g111_n;
  wire g112_p;
  wire g112_n;
  wire g113_p;
  wire g113_n;
  wire g114_p;
  wire g114_n;
  wire g115_p;
  wire g115_n;
  wire g116_p;
  wire g116_n;
  wire g117_p;
  wire g117_n;
  wire g118_p;
  wire g118_n;
  wire g119_p;
  wire g119_n;
  wire g120_p;
  wire g120_n;
  wire g121_p;
  wire g121_n;
  wire g122_p;
  wire g122_n;
  wire g123_p;
  wire g123_n;
  wire g124_p;
  wire g124_n;
  wire g125_p;
  wire g125_n;
  wire g126_p;
  wire g126_n;
  wire g127_p;
  wire g127_n;
  wire g128_p;
  wire g128_n;
  wire g129_p;
  wire g129_n;
  wire g130_p;
  wire g130_n;
  wire g131_p;
  wire g131_n;
  wire g132_p;
  wire g132_n;
  wire g133_p;
  wire g133_n;
  wire g134_p;
  wire g134_n;
  wire g135_p;
  wire g135_n;
  wire g136_p;
  wire g136_n;
  wire g137_p;
  wire g137_n;
  wire g138_p;
  wire g138_n;
  wire g139_p;
  wire g139_n;
  wire g140_p;
  wire g140_n;
  wire g141_p;
  wire g141_n;
  wire g142_p;
  wire g142_n;
  wire g143_p;
  wire g143_n;
  wire g144_p;
  wire g144_n;
  wire g145_p;
  wire g145_n;
  wire g146_p;
  wire g146_n;
  wire g147_p;
  wire g147_n;
  wire g148_p;
  wire g148_n;
  wire g149_p;
  wire g149_n;
  wire g150_p;
  wire g150_n;
  wire g151_p;
  wire g151_n;
  wire g152_p;
  wire g152_n;
  wire g153_p;
  wire g153_n;
  wire g154_p;
  wire g154_n;
  wire g155_p;
  wire g155_n;
  wire g156_p;
  wire g156_n;
  wire g157_p;
  wire g157_n;
  wire g158_p;
  wire g158_n;
  wire g159_p;
  wire g159_n;
  wire g160_p;
  wire g160_n;
  wire g161_p;
  wire g161_n;
  wire g162_p;
  wire g162_n;
  wire g163_p;
  wire g163_n;
  wire g164_p;
  wire g164_n;
  wire g165_p;
  wire g165_n;
  wire g166_p;
  wire g166_n;
  wire g167_p;
  wire g167_n;
  wire g168_p;
  wire g168_n;
  wire g169_p;
  wire g169_n;
  wire g170_p;
  wire g170_n;
  wire g171_p;
  wire g171_n;
  wire g172_p;
  wire g172_n;
  wire g173_p;
  wire g173_n;
  wire g174_p;
  wire g174_n;
  wire g175_p;
  wire g175_n;
  wire g176_p;
  wire g176_n;
  wire g177_p;
  wire g177_n;
  wire g178_p;
  wire g178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire G33_n_spl_;
  wire G33_n_spl_0;
  wire G33_n_spl_00;
  wire G33_n_spl_000;
  wire G33_n_spl_001;
  wire G33_n_spl_01;
  wire G33_n_spl_010;
  wire G33_n_spl_011;
  wire G33_n_spl_1;
  wire G33_n_spl_10;
  wire G33_n_spl_11;
  wire G29_n_spl_;
  wire G33_p_spl_;
  wire G33_p_spl_0;
  wire G33_p_spl_00;
  wire G33_p_spl_000;
  wire G33_p_spl_001;
  wire G33_p_spl_01;
  wire G33_p_spl_010;
  wire G33_p_spl_1;
  wire G33_p_spl_10;
  wire G33_p_spl_11;
  wire G29_p_spl_;
  wire G24_p_spl_;
  wire G24_p_spl_0;
  wire G24_p_spl_1;
  wire G23_n_spl_;
  wire G23_n_spl_0;
  wire G23_n_spl_1;
  wire G24_n_spl_;
  wire G24_n_spl_0;
  wire G24_n_spl_1;
  wire G23_p_spl_;
  wire G23_p_spl_0;
  wire G23_p_spl_1;
  wire g35_n_spl_;
  wire G31_n_spl_;
  wire G31_n_spl_0;
  wire G31_n_spl_00;
  wire G31_n_spl_000;
  wire G31_n_spl_001;
  wire G31_n_spl_01;
  wire G31_n_spl_010;
  wire G31_n_spl_011;
  wire G31_n_spl_1;
  wire G31_n_spl_10;
  wire G31_n_spl_11;
  wire g35_p_spl_;
  wire G31_p_spl_;
  wire G31_p_spl_0;
  wire G31_p_spl_00;
  wire G31_p_spl_000;
  wire G31_p_spl_001;
  wire G31_p_spl_01;
  wire G31_p_spl_010;
  wire G31_p_spl_011;
  wire G31_p_spl_1;
  wire G31_p_spl_10;
  wire G31_p_spl_100;
  wire G31_p_spl_101;
  wire G31_p_spl_11;
  wire G31_p_spl_110;
  wire g36_p_spl_;
  wire g34_p_spl_;
  wire g36_n_spl_;
  wire g34_n_spl_;
  wire G32_n_spl_;
  wire g38_p_spl_;
  wire g38_p_spl_0;
  wire g38_p_spl_00;
  wire g38_p_spl_01;
  wire g38_p_spl_1;
  wire g38_p_spl_10;
  wire g39_n_spl_;
  wire g39_p_spl_;
  wire g41_n_spl_;
  wire G20_p_spl_;
  wire g41_p_spl_;
  wire G20_n_spl_;
  wire G22_p_spl_;
  wire G22_n_spl_;
  wire G14_n_spl_;
  wire G14_n_spl_0;
  wire G14_n_spl_00;
  wire G14_n_spl_1;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_00;
  wire G4_p_spl_01;
  wire G4_p_spl_1;
  wire G4_p_spl_10;
  wire G14_p_spl_;
  wire G14_p_spl_0;
  wire G14_p_spl_00;
  wire G14_p_spl_1;
  wire G4_n_spl_;
  wire G4_n_spl_0;
  wire G4_n_spl_00;
  wire G4_n_spl_01;
  wire G4_n_spl_1;
  wire G4_n_spl_10;
  wire g46_p_spl_;
  wire g43_p_spl_;
  wire g46_n_spl_;
  wire g43_n_spl_;
  wire G13_n_spl_;
  wire G13_n_spl_0;
  wire G13_n_spl_00;
  wire G13_n_spl_1;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire G12_p_spl_00;
  wire G12_p_spl_1;
  wire G13_p_spl_;
  wire G13_p_spl_0;
  wire G13_p_spl_00;
  wire G13_p_spl_1;
  wire G12_n_spl_;
  wire G12_n_spl_0;
  wire G12_n_spl_00;
  wire G12_n_spl_1;
  wire g52_p_spl_;
  wire G11_p_spl_;
  wire G11_p_spl_0;
  wire G11_p_spl_00;
  wire G11_p_spl_1;
  wire g52_n_spl_;
  wire G11_n_spl_;
  wire G11_n_spl_0;
  wire G11_n_spl_00;
  wire G11_n_spl_1;
  wire G15_n_spl_;
  wire G15_n_spl_0;
  wire G15_n_spl_00;
  wire G15_n_spl_1;
  wire G10_n_spl_;
  wire G10_n_spl_0;
  wire G10_n_spl_00;
  wire G10_n_spl_1;
  wire G15_p_spl_;
  wire G15_p_spl_0;
  wire G15_p_spl_00;
  wire G15_p_spl_1;
  wire G10_p_spl_;
  wire G10_p_spl_0;
  wire G10_p_spl_00;
  wire G10_p_spl_1;
  wire g58_n_spl_;
  wire g58_n_spl_0;
  wire g58_n_spl_1;
  wire G16_p_spl_;
  wire G16_p_spl_0;
  wire G16_p_spl_00;
  wire G16_p_spl_1;
  wire g58_p_spl_;
  wire g58_p_spl_0;
  wire g58_p_spl_1;
  wire G16_n_spl_;
  wire G16_n_spl_0;
  wire G16_n_spl_00;
  wire G16_n_spl_1;
  wire g61_p_spl_;
  wire g61_p_spl_0;
  wire g61_p_spl_1;
  wire g55_n_spl_;
  wire g61_n_spl_;
  wire g61_n_spl_0;
  wire g61_n_spl_1;
  wire g55_p_spl_;
  wire G3_n_spl_;
  wire G3_n_spl_0;
  wire G3_n_spl_00;
  wire G3_n_spl_1;
  wire G2_p_spl_;
  wire G2_p_spl_0;
  wire G2_p_spl_00;
  wire G2_p_spl_1;
  wire G3_p_spl_;
  wire G3_p_spl_0;
  wire G3_p_spl_00;
  wire G3_p_spl_1;
  wire G2_n_spl_;
  wire G2_n_spl_0;
  wire G2_n_spl_00;
  wire G2_n_spl_1;
  wire g67_p_spl_;
  wire G1_p_spl_;
  wire G1_p_spl_0;
  wire G1_p_spl_00;
  wire G1_p_spl_1;
  wire g67_n_spl_;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire G1_n_spl_00;
  wire G1_n_spl_1;
  wire g70_n_spl_;
  wire g70_n_spl_0;
  wire g70_n_spl_1;
  wire g64_n_spl_;
  wire g64_n_spl_0;
  wire g64_n_spl_00;
  wire g64_n_spl_01;
  wire g64_n_spl_1;
  wire g70_p_spl_;
  wire g70_p_spl_0;
  wire g70_p_spl_1;
  wire g64_p_spl_;
  wire g64_p_spl_0;
  wire g64_p_spl_00;
  wire g64_p_spl_01;
  wire g64_p_spl_1;
  wire g73_n_spl_;
  wire g49_n_spl_;
  wire g73_p_spl_;
  wire g49_p_spl_;
  wire g76_n_spl_;
  wire g76_p_spl_;
  wire g77_p_spl_;
  wire G25_n_spl_;
  wire G25_n_spl_0;
  wire g77_n_spl_;
  wire G25_p_spl_;
  wire G25_p_spl_0;
  wire g80_n_spl_;
  wire g80_n_spl_0;
  wire g42_p_spl_;
  wire g42_p_spl_0;
  wire g80_p_spl_;
  wire g42_n_spl_;
  wire G18_p_spl_;
  wire G18_n_spl_;
  wire g83_n_spl_;
  wire g83_p_spl_;
  wire g86_n_spl_;
  wire g86_p_spl_;
  wire G9_p_spl_;
  wire G9_p_spl_0;
  wire G9_p_spl_00;
  wire G9_p_spl_1;
  wire G9_n_spl_;
  wire G9_n_spl_0;
  wire G9_n_spl_00;
  wire G9_n_spl_1;
  wire g92_n_spl_;
  wire g92_n_spl_0;
  wire g92_n_spl_1;
  wire g92_p_spl_;
  wire g92_p_spl_0;
  wire g92_p_spl_1;
  wire g95_p_spl_;
  wire g95_p_spl_0;
  wire g95_p_spl_1;
  wire g89_p_spl_;
  wire g95_n_spl_;
  wire g95_n_spl_0;
  wire g95_n_spl_1;
  wire g89_n_spl_;
  wire G8_n_spl_;
  wire G8_n_spl_0;
  wire G8_n_spl_00;
  wire G8_n_spl_01;
  wire G8_n_spl_1;
  wire G8_n_spl_10;
  wire G5_n_spl_;
  wire G5_n_spl_0;
  wire G5_n_spl_00;
  wire G5_n_spl_1;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire G8_p_spl_00;
  wire G8_p_spl_01;
  wire G8_p_spl_1;
  wire G8_p_spl_10;
  wire G5_p_spl_;
  wire G5_p_spl_0;
  wire G5_p_spl_00;
  wire G5_p_spl_1;
  wire g101_p_spl_;
  wire g101_n_spl_;
  wire g104_p_spl_;
  wire g98_n_spl_;
  wire g104_n_spl_;
  wire g98_p_spl_;
  wire g107_n_spl_;
  wire g108_p_spl_;
  wire G27_n_spl_;
  wire G27_n_spl_0;
  wire g108_n_spl_;
  wire G27_p_spl_;
  wire G6_n_spl_;
  wire G6_n_spl_0;
  wire G6_n_spl_00;
  wire G6_n_spl_1;
  wire G6_p_spl_;
  wire G6_p_spl_0;
  wire G6_p_spl_00;
  wire G6_p_spl_1;
  wire g112_p_spl_;
  wire g112_n_spl_;
  wire g118_n_spl_;
  wire g115_n_spl_;
  wire g118_p_spl_;
  wire g115_p_spl_;
  wire G19_p_spl_;
  wire G19_n_spl_;
  wire g123_n_spl_;
  wire g121_n_spl_;
  wire g123_p_spl_;
  wire g121_p_spl_;
  wire g126_n_spl_;
  wire g127_p_spl_;
  wire G28_n_spl_;
  wire G28_n_spl_0;
  wire g127_n_spl_;
  wire G28_p_spl_;
  wire G7_n_spl_;
  wire G7_n_spl_0;
  wire G7_n_spl_00;
  wire G7_n_spl_1;
  wire G7_p_spl_;
  wire G7_p_spl_0;
  wire G7_p_spl_00;
  wire G7_p_spl_1;
  wire g133_p_spl_;
  wire g133_n_spl_;
  wire g136_n_spl_;
  wire g136_p_spl_;
  wire g141_p_spl_;
  wire g141_n_spl_;
  wire g144_n_spl_;
  wire g139_n_spl_;
  wire g144_p_spl_;
  wire g139_p_spl_;
  wire g147_n_spl_;
  wire g149_n_spl_;
  wire g149_n_spl_0;
  wire g148_p_spl_;
  wire g149_p_spl_;
  wire g148_n_spl_;
  wire G17_p_spl_;
  wire G17_n_spl_;
  wire g156_p_spl_;
  wire g156_n_spl_;
  wire g162_p_spl_;
  wire g162_n_spl_;
  wire g165_n_spl_;
  wire g165_n_spl_0;
  wire g165_n_spl_1;
  wire g165_p_spl_;
  wire g165_p_spl_0;
  wire g165_p_spl_1;
  wire g168_p_spl_;
  wire g159_p_spl_;
  wire g168_n_spl_;
  wire g159_n_spl_;
  wire g171_n_spl_;
  wire g171_p_spl_;
  wire g172_n_spl_;
  wire G26_p_spl_;
  wire G26_p_spl_0;
  wire g172_p_spl_;
  wire G26_n_spl_;
  wire G26_n_spl_0;
  wire g179_n_spl_;
  wire g179_p_spl_;
  wire G21_p_spl_;
  wire G21_n_spl_;
  wire g184_p_spl_;
  wire g181_p_spl_;
  wire g184_n_spl_;
  wire g181_n_spl_;
  wire g193_n_spl_;
  wire g190_p_spl_;
  wire g193_p_spl_;
  wire g190_n_spl_;
  wire g196_n_spl_;
  wire g196_n_spl_0;
  wire g187_p_spl_;
  wire g196_p_spl_;
  wire g196_p_spl_0;
  wire g187_n_spl_;
  wire g199_p_spl_;
  wire g199_n_spl_;
  wire g201_n_spl_;
  wire g201_n_spl_0;
  wire g200_p_spl_;
  wire g201_p_spl_;
  wire g201_p_spl_0;
  wire g200_n_spl_;
  wire g204_n_spl_;
  wire g204_n_spl_0;
  wire g180_p_spl_;
  wire g180_p_spl_0;
  wire g204_p_spl_;
  wire g180_n_spl_;
  wire g178_p_spl_;
  wire g178_n_spl_;
  wire g178_n_spl_0;
  wire g206_p_spl_;
  wire g81_n_spl_;
  wire g206_n_spl_;
  wire g81_p_spl_;
  wire g207_p_spl_;
  wire g40_n_spl_;
  wire g207_n_spl_;
  wire g40_p_spl_;
  wire g208_n_spl_;
  wire g208_n_spl_0;
  wire g208_n_spl_00;
  wire g208_n_spl_01;
  wire g208_n_spl_1;
  wire g208_n_spl_10;
  wire g208_p_spl_;
  wire g208_p_spl_0;
  wire g208_p_spl_00;
  wire g208_p_spl_01;
  wire g208_p_spl_1;
  wire g208_p_spl_10;
  wire G30_n_spl_;
  wire G30_p_spl_;
  wire g221_p_spl_;
  wire g221_n_spl_;
  wire g223_n_spl_;
  wire g223_n_spl_0;
  wire g223_p_spl_;
  wire g223_p_spl_0;
  wire g224_n_spl_;
  wire g224_n_spl_0;
  wire g224_n_spl_00;
  wire g224_n_spl_01;
  wire g224_n_spl_1;
  wire g224_p_spl_;
  wire g224_p_spl_0;
  wire g224_p_spl_00;
  wire g224_p_spl_01;
  wire g224_p_spl_1;
  wire g235_p_spl_;
  wire g235_n_spl_;
  wire g236_n_spl_;
  wire g236_n_spl_0;
  wire g236_n_spl_1;
  wire g236_p_spl_;
  wire g236_p_spl_0;
  wire g236_p_spl_1;
  wire g256_n_spl_;
  wire g256_n_spl_0;
  wire g256_n_spl_1;
  wire g256_p_spl_;
  wire g256_p_spl_0;
  wire g256_p_spl_1;
  wire g269_p_spl_;
  wire g269_p_spl_0;
  wire g269_p_spl_00;
  wire g269_p_spl_01;
  wire g269_p_spl_1;
  wire g269_p_spl_10;
  wire g269_n_spl_;
  wire g269_n_spl_0;
  wire g303_n_spl_;
  wire g303_p_spl_;
  wire g315_n_spl_;
  wire g315_p_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  and

  (
    g34_p,
    G33_n_spl_000,
    G29_n_spl_
  );


  or

  (
    g34_n,
    G33_p_spl_000,
    G29_p_spl_
  );


  and

  (
    g35_p,
    G24_p_spl_0,
    G23_n_spl_0
  );


  or

  (
    g35_n,
    G24_n_spl_0,
    G23_p_spl_0
  );


  and

  (
    g36_p,
    g35_n_spl_,
    G31_n_spl_000
  );


  or

  (
    g36_n,
    g35_p_spl_,
    G31_p_spl_000
  );


  and

  (
    g37_p,
    g36_p_spl_,
    g34_p_spl_
  );


  or

  (
    g37_n,
    g36_n_spl_,
    g34_n_spl_
  );


  and

  (
    g38_p,
    G33_n_spl_000,
    G32_n_spl_
  );


  or

  (
    g38_n,
    G33_p_spl_000,
    G32_p
  );


  and

  (
    g39_p,
    g38_p_spl_00,
    g35_n_spl_
  );


  or

  (
    g39_n,
    g38_n,
    g35_p_spl_
  );


  and

  (
    g40_p,
    g39_n_spl_,
    g37_n
  );


  or

  (
    g40_n,
    g39_p_spl_,
    g37_p
  );


  and

  (
    g41_p,
    G31_n_spl_000,
    G23_n_spl_0
  );


  or

  (
    g41_n,
    G31_p_spl_000,
    G23_p_spl_0
  );


  and

  (
    g42_p,
    g41_n_spl_,
    G20_p_spl_
  );


  or

  (
    g42_n,
    g41_p_spl_,
    G20_n_spl_
  );


  and

  (
    g43_p,
    G33_n_spl_001,
    G22_p_spl_
  );


  or

  (
    g43_n,
    G33_p_spl_001,
    G22_n_spl_
  );


  and

  (
    g44_p,
    G14_n_spl_00,
    G4_p_spl_00
  );


  or

  (
    g44_n,
    G14_p_spl_00,
    G4_n_spl_00
  );


  and

  (
    g45_p,
    G14_p_spl_00,
    G4_n_spl_00
  );


  or

  (
    g45_n,
    G14_n_spl_00,
    G4_p_spl_00
  );


  and

  (
    g46_p,
    g45_n,
    g44_n
  );


  or

  (
    g46_n,
    g45_p,
    g44_p
  );


  and

  (
    g47_p,
    g46_p_spl_,
    g43_p_spl_
  );


  or

  (
    g47_n,
    g46_n_spl_,
    g43_n_spl_
  );


  and

  (
    g48_p,
    g46_n_spl_,
    g43_n_spl_
  );


  or

  (
    g48_n,
    g46_p_spl_,
    g43_p_spl_
  );


  and

  (
    g49_p,
    g48_n,
    g47_n
  );


  or

  (
    g49_n,
    g48_p,
    g47_p
  );


  and

  (
    g50_p,
    G13_n_spl_00,
    G12_p_spl_00
  );


  or

  (
    g50_n,
    G13_p_spl_00,
    G12_n_spl_00
  );


  and

  (
    g51_p,
    G13_p_spl_00,
    G12_n_spl_00
  );


  or

  (
    g51_n,
    G13_n_spl_00,
    G12_p_spl_00
  );


  and

  (
    g52_p,
    g51_n,
    g50_n
  );


  or

  (
    g52_n,
    g51_p,
    g50_p
  );


  and

  (
    g53_p,
    g52_p_spl_,
    G11_p_spl_00
  );


  or

  (
    g53_n,
    g52_n_spl_,
    G11_n_spl_00
  );


  and

  (
    g54_p,
    g52_n_spl_,
    G11_n_spl_00
  );


  or

  (
    g54_n,
    g52_p_spl_,
    G11_p_spl_00
  );


  and

  (
    g55_p,
    g54_n,
    g53_n
  );


  or

  (
    g55_n,
    g54_p,
    g53_p
  );


  and

  (
    g56_p,
    G15_n_spl_00,
    G10_n_spl_00
  );


  or

  (
    g56_n,
    G15_p_spl_00,
    G10_p_spl_00
  );


  and

  (
    g57_p,
    G15_p_spl_00,
    G10_p_spl_00
  );


  or

  (
    g57_n,
    G15_n_spl_00,
    G10_n_spl_00
  );


  and

  (
    g58_p,
    g57_n,
    g56_n
  );


  or

  (
    g58_n,
    g57_p,
    g56_p
  );


  and

  (
    g59_p,
    g58_n_spl_0,
    G16_p_spl_00
  );


  or

  (
    g59_n,
    g58_p_spl_0,
    G16_n_spl_00
  );


  and

  (
    g60_p,
    g58_p_spl_0,
    G16_n_spl_00
  );


  or

  (
    g60_n,
    g58_n_spl_0,
    G16_p_spl_00
  );


  and

  (
    g61_p,
    g60_n,
    g59_n
  );


  or

  (
    g61_n,
    g60_p,
    g59_p
  );


  and

  (
    g62_p,
    g61_p_spl_0,
    g55_n_spl_
  );


  or

  (
    g62_n,
    g61_n_spl_0,
    g55_p_spl_
  );


  and

  (
    g63_p,
    g61_n_spl_0,
    g55_p_spl_
  );


  or

  (
    g63_n,
    g61_p_spl_0,
    g55_n_spl_
  );


  and

  (
    g64_p,
    g63_n,
    g62_n
  );


  or

  (
    g64_n,
    g63_p,
    g62_p
  );


  and

  (
    g65_p,
    G3_n_spl_00,
    G2_p_spl_00
  );


  or

  (
    g65_n,
    G3_p_spl_00,
    G2_n_spl_00
  );


  and

  (
    g66_p,
    G3_p_spl_00,
    G2_n_spl_00
  );


  or

  (
    g66_n,
    G3_n_spl_00,
    G2_p_spl_00
  );


  and

  (
    g67_p,
    g66_n,
    g65_n
  );


  or

  (
    g67_n,
    g66_p,
    g65_p
  );


  and

  (
    g68_p,
    g67_p_spl_,
    G1_p_spl_00
  );


  or

  (
    g68_n,
    g67_n_spl_,
    G1_n_spl_00
  );


  and

  (
    g69_p,
    g67_n_spl_,
    G1_n_spl_00
  );


  or

  (
    g69_n,
    g67_p_spl_,
    G1_p_spl_00
  );


  and

  (
    g70_p,
    g69_n,
    g68_n
  );


  or

  (
    g70_n,
    g69_p,
    g68_p
  );


  and

  (
    g71_p,
    g70_n_spl_0,
    g64_n_spl_00
  );


  or

  (
    g71_n,
    g70_p_spl_0,
    g64_p_spl_00
  );


  and

  (
    g72_p,
    g70_p_spl_0,
    g64_p_spl_00
  );


  or

  (
    g72_n,
    g70_n_spl_0,
    g64_n_spl_00
  );


  and

  (
    g73_p,
    g72_n,
    g71_n
  );


  or

  (
    g73_n,
    g72_p,
    g71_p
  );


  and

  (
    g74_p,
    g73_n_spl_,
    g49_n_spl_
  );


  or

  (
    g74_n,
    g73_p_spl_,
    g49_p_spl_
  );


  and

  (
    g75_p,
    g73_p_spl_,
    g49_p_spl_
  );


  or

  (
    g75_n,
    g73_n_spl_,
    g49_n_spl_
  );


  and

  (
    g76_p,
    g75_n,
    g74_n
  );


  or

  (
    g76_n,
    g75_p,
    g74_p
  );


  and

  (
    g77_p,
    g76_n_spl_,
    G31_n_spl_001
  );


  or

  (
    g77_n,
    g76_p_spl_,
    G31_p_spl_001
  );


  and

  (
    g78_p,
    g77_p_spl_,
    G25_n_spl_0
  );


  or

  (
    g78_n,
    g77_n_spl_,
    G25_p_spl_0
  );


  and

  (
    g79_p,
    g77_n_spl_,
    G25_p_spl_0
  );


  or

  (
    g79_n,
    g77_p_spl_,
    G25_n_spl_0
  );


  and

  (
    g80_p,
    g79_n,
    g78_n
  );


  or

  (
    g80_n,
    g79_p,
    g78_p
  );


  and

  (
    g81_p,
    g80_n_spl_0,
    g42_p_spl_0
  );


  or

  (
    g81_n,
    g80_p_spl_,
    g42_n_spl_
  );


  and

  (
    g82_p,
    G33_n_spl_001,
    G18_p_spl_
  );


  or

  (
    g82_n,
    G33_p_spl_001,
    G18_n_spl_
  );


  and

  (
    g83_p,
    g82_p,
    G24_n_spl_0
  );


  or

  (
    g83_n,
    g82_n,
    G24_p_spl_0
  );


  and

  (
    g84_p,
    g83_n_spl_,
    G15_p_spl_0
  );


  or

  (
    g84_n,
    g83_p_spl_,
    G15_n_spl_0
  );


  and

  (
    g85_p,
    g83_p_spl_,
    G15_n_spl_1
  );


  or

  (
    g85_n,
    g83_n_spl_,
    G15_p_spl_1
  );


  and

  (
    g86_p,
    g85_n,
    g84_n
  );


  or

  (
    g86_n,
    g85_p,
    g84_p
  );


  and

  (
    g87_p,
    g86_n_spl_,
    G11_n_spl_0
  );


  or

  (
    g87_n,
    g86_p_spl_,
    G11_p_spl_0
  );


  and

  (
    g88_p,
    g86_p_spl_,
    G11_p_spl_1
  );


  or

  (
    g88_n,
    g86_n_spl_,
    G11_n_spl_1
  );


  and

  (
    g89_p,
    g88_n,
    g87_n
  );


  or

  (
    g89_n,
    g88_p,
    g87_p
  );


  and

  (
    g90_p,
    G14_n_spl_0,
    G9_p_spl_00
  );


  or

  (
    g90_n,
    G14_p_spl_0,
    G9_n_spl_00
  );


  and

  (
    g91_p,
    G14_p_spl_1,
    G9_n_spl_00
  );


  or

  (
    g91_n,
    G14_n_spl_1,
    G9_p_spl_00
  );


  and

  (
    g92_p,
    g91_n,
    g90_n
  );


  or

  (
    g92_n,
    g91_p,
    g90_p
  );


  and

  (
    g93_p,
    g92_n_spl_0,
    G16_p_spl_0
  );


  or

  (
    g93_n,
    g92_p_spl_0,
    G16_n_spl_0
  );


  and

  (
    g94_p,
    g92_p_spl_0,
    G16_n_spl_1
  );


  or

  (
    g94_n,
    g92_n_spl_0,
    G16_p_spl_1
  );


  and

  (
    g95_p,
    g94_n,
    g93_n
  );


  or

  (
    g95_n,
    g94_p,
    g93_p
  );


  and

  (
    g96_p,
    g95_p_spl_0,
    g89_p_spl_
  );


  or

  (
    g96_n,
    g95_n_spl_0,
    g89_n_spl_
  );


  and

  (
    g97_p,
    g95_n_spl_0,
    g89_n_spl_
  );


  or

  (
    g97_n,
    g95_p_spl_0,
    g89_p_spl_
  );


  and

  (
    g98_p,
    g97_n,
    g96_n
  );


  or

  (
    g98_n,
    g97_p,
    g96_p
  );


  and

  (
    g99_p,
    G8_n_spl_00,
    G5_n_spl_00
  );


  or

  (
    g99_n,
    G8_p_spl_00,
    G5_p_spl_00
  );


  and

  (
    g100_p,
    G8_p_spl_00,
    G5_p_spl_00
  );


  or

  (
    g100_n,
    G8_n_spl_00,
    G5_n_spl_00
  );


  and

  (
    g101_p,
    g100_n,
    g99_n
  );


  or

  (
    g101_n,
    g100_p,
    g99_p
  );


  and

  (
    g102_p,
    g101_p_spl_,
    G2_n_spl_0
  );


  or

  (
    g102_n,
    g101_n_spl_,
    G2_p_spl_0
  );


  and

  (
    g103_p,
    g101_n_spl_,
    G2_p_spl_1
  );


  or

  (
    g103_n,
    g101_p_spl_,
    G2_n_spl_1
  );


  and

  (
    g104_p,
    g103_n,
    g102_n
  );


  or

  (
    g104_n,
    g103_p,
    g102_p
  );


  and

  (
    g105_p,
    g104_p_spl_,
    g98_n_spl_
  );


  or

  (
    g105_n,
    g104_n_spl_,
    g98_p_spl_
  );


  and

  (
    g106_p,
    g104_n_spl_,
    g98_p_spl_
  );


  or

  (
    g106_n,
    g104_p_spl_,
    g98_n_spl_
  );


  and

  (
    g107_p,
    g106_n,
    g105_n
  );


  or

  (
    g107_n,
    g106_p,
    g105_p
  );


  and

  (
    g108_p,
    g107_n_spl_,
    G31_n_spl_001
  );


  or

  (
    g108_n,
    g107_p,
    G31_p_spl_001
  );


  and

  (
    g109_p,
    g108_p_spl_,
    G27_n_spl_0
  );


  or

  (
    g109_n,
    g108_n_spl_,
    G27_p_spl_
  );


  and

  (
    g110_p,
    G8_n_spl_01,
    G6_n_spl_00
  );


  or

  (
    g110_n,
    G8_p_spl_01,
    G6_p_spl_00
  );


  and

  (
    g111_p,
    G8_p_spl_01,
    G6_p_spl_00
  );


  or

  (
    g111_n,
    G8_n_spl_01,
    G6_n_spl_00
  );


  and

  (
    g112_p,
    g111_n,
    g110_n
  );


  or

  (
    g112_n,
    g111_p,
    g110_p
  );


  and

  (
    g113_p,
    g112_p_spl_,
    G3_n_spl_0
  );


  or

  (
    g113_n,
    g112_n_spl_,
    G3_p_spl_0
  );


  and

  (
    g114_p,
    g112_n_spl_,
    G3_p_spl_1
  );


  or

  (
    g114_n,
    g112_p_spl_,
    G3_n_spl_1
  );


  and

  (
    g115_p,
    g114_n,
    g113_n
  );


  or

  (
    g115_n,
    g114_p,
    g113_p
  );


  and

  (
    g116_p,
    g58_n_spl_1,
    G12_n_spl_0
  );


  or

  (
    g116_n,
    g58_p_spl_1,
    G12_p_spl_0
  );


  and

  (
    g117_p,
    g58_p_spl_1,
    G12_p_spl_1
  );


  or

  (
    g117_n,
    g58_n_spl_1,
    G12_n_spl_1
  );


  and

  (
    g118_p,
    g117_n,
    g116_n
  );


  or

  (
    g118_n,
    g117_p,
    g116_p
  );


  and

  (
    g119_p,
    g118_n_spl_,
    g115_n_spl_
  );


  or

  (
    g119_n,
    g118_p_spl_,
    g115_p_spl_
  );


  and

  (
    g120_p,
    g118_p_spl_,
    g115_p_spl_
  );


  or

  (
    g120_n,
    g118_n_spl_,
    g115_n_spl_
  );


  and

  (
    g121_p,
    g120_n,
    g119_n
  );


  or

  (
    g121_n,
    g120_p,
    g119_p
  );


  and

  (
    g122_p,
    G33_n_spl_010,
    G19_p_spl_
  );


  or

  (
    g122_n,
    G33_p_spl_010,
    G19_n_spl_
  );


  and

  (
    g123_p,
    g122_p,
    G23_n_spl_1
  );


  or

  (
    g123_n,
    g122_n,
    G23_p_spl_1
  );


  and

  (
    g124_p,
    g123_n_spl_,
    g121_n_spl_
  );


  or

  (
    g124_n,
    g123_p_spl_,
    g121_p_spl_
  );


  and

  (
    g125_p,
    g123_p_spl_,
    g121_p_spl_
  );


  or

  (
    g125_n,
    g123_n_spl_,
    g121_n_spl_
  );


  and

  (
    g126_p,
    g125_n,
    g124_n
  );


  or

  (
    g126_n,
    g125_p,
    g124_p
  );


  and

  (
    g127_p,
    g126_n_spl_,
    G31_n_spl_010
  );


  or

  (
    g127_n,
    g126_p,
    G31_p_spl_010
  );


  and

  (
    g128_p,
    g127_p_spl_,
    G28_n_spl_0
  );


  or

  (
    g128_n,
    g127_n_spl_,
    G28_p_spl_
  );


  and

  (
    g129_p,
    g127_n_spl_,
    G28_p_spl_
  );


  or

  (
    g129_n,
    g127_p_spl_,
    G28_n_spl_0
  );


  and

  (
    g130_p,
    g129_n,
    g128_n
  );


  or

  (
    g130_n,
    g129_p,
    g128_p
  );


  and

  (
    g131_p,
    G10_n_spl_0,
    G7_n_spl_00
  );


  or

  (
    g131_n,
    G10_p_spl_0,
    G7_p_spl_00
  );


  and

  (
    g132_p,
    G10_p_spl_1,
    G7_p_spl_00
  );


  or

  (
    g132_n,
    G10_n_spl_1,
    G7_n_spl_00
  );


  and

  (
    g133_p,
    g132_n,
    g131_n
  );


  or

  (
    g133_n,
    g132_p,
    g131_p
  );


  and

  (
    g134_p,
    g133_p_spl_,
    G4_n_spl_01
  );


  or

  (
    g134_n,
    g133_n_spl_,
    G4_p_spl_01
  );


  and

  (
    g135_p,
    g133_n_spl_,
    G4_p_spl_01
  );


  or

  (
    g135_n,
    g133_p_spl_,
    G4_n_spl_01
  );


  and

  (
    g136_p,
    g135_n,
    g134_n
  );


  or

  (
    g136_n,
    g135_p,
    g134_p
  );


  and

  (
    g137_p,
    g136_n_spl_,
    g95_n_spl_1
  );


  or

  (
    g137_n,
    g136_p_spl_,
    g95_p_spl_1
  );


  and

  (
    g138_p,
    g136_p_spl_,
    g95_p_spl_1
  );


  or

  (
    g138_n,
    g136_n_spl_,
    g95_n_spl_1
  );


  and

  (
    g139_p,
    g138_n,
    g137_n
  );


  or

  (
    g139_n,
    g138_p,
    g137_p
  );


  and

  (
    g140_p,
    G33_n_spl_010,
    G20_p_spl_
  );


  or

  (
    g140_n,
    G33_p_spl_010,
    G20_n_spl_
  );


  and

  (
    g141_p,
    g140_p,
    G23_n_spl_1
  );


  or

  (
    g141_n,
    g140_n,
    G23_p_spl_1
  );


  and

  (
    g142_p,
    g141_p_spl_,
    G13_n_spl_0
  );


  or

  (
    g142_n,
    g141_n_spl_,
    G13_p_spl_0
  );


  and

  (
    g143_p,
    g141_n_spl_,
    G13_p_spl_1
  );


  or

  (
    g143_n,
    g141_p_spl_,
    G13_n_spl_1
  );


  and

  (
    g144_p,
    g143_n,
    g142_n
  );


  or

  (
    g144_n,
    g143_p,
    g142_p
  );


  and

  (
    g145_p,
    g144_n_spl_,
    g139_n_spl_
  );


  or

  (
    g145_n,
    g144_p_spl_,
    g139_p_spl_
  );


  and

  (
    g146_p,
    g144_p_spl_,
    g139_p_spl_
  );


  or

  (
    g146_n,
    g144_n_spl_,
    g139_n_spl_
  );


  and

  (
    g147_p,
    g146_n,
    g145_n
  );


  or

  (
    g147_n,
    g146_p,
    g145_p
  );


  and

  (
    g148_p,
    g147_n_spl_,
    G31_n_spl_010
  );


  or

  (
    g148_n,
    g147_p,
    G31_p_spl_010
  );


  and

  (
    g149_p,
    g41_n_spl_,
    G19_p_spl_
  );


  or

  (
    g149_n,
    g41_p_spl_,
    G19_n_spl_
  );


  and

  (
    g150_p,
    g149_n_spl_0,
    g148_p_spl_
  );


  or

  (
    g150_n,
    g149_p_spl_,
    g148_n_spl_
  );


  and

  (
    g151_p,
    g149_p_spl_,
    g148_n_spl_
  );


  or

  (
    g151_n,
    g149_n_spl_0,
    g148_p_spl_
  );


  and

  (
    g152_p,
    g151_n,
    g150_n
  );


  or

  (
    g152_n,
    g151_p,
    g150_p
  );


  and

  (
    g153_p,
    g152_p,
    g130_p
  );


  or

  (
    g153_n,
    g152_n,
    g130_n
  );


  and

  (
    g154_p,
    g153_p,
    g109_n
  );


  or

  (
    g154_n,
    g153_n,
    g109_p
  );


  and

  (
    g155_p,
    G33_n_spl_011,
    G17_p_spl_
  );


  or

  (
    g155_n,
    G33_p_spl_01,
    G17_n_spl_
  );


  and

  (
    g156_p,
    g155_p,
    G24_n_spl_1
  );


  or

  (
    g156_n,
    g155_n,
    G24_p_spl_1
  );


  and

  (
    g157_p,
    g156_p_spl_,
    G1_p_spl_0
  );


  or

  (
    g157_n,
    g156_n_spl_,
    G1_n_spl_0
  );


  and

  (
    g158_p,
    g156_n_spl_,
    G1_n_spl_1
  );


  or

  (
    g158_n,
    g156_p_spl_,
    G1_p_spl_1
  );


  and

  (
    g159_p,
    g158_n,
    g157_n
  );


  or

  (
    g159_n,
    g158_p,
    g157_p
  );


  and

  (
    g160_p,
    G7_n_spl_0,
    G6_p_spl_0
  );


  or

  (
    g160_n,
    G7_p_spl_0,
    G6_n_spl_0
  );


  and

  (
    g161_p,
    G7_p_spl_1,
    G6_n_spl_1
  );


  or

  (
    g161_n,
    G7_n_spl_1,
    G6_p_spl_1
  );


  and

  (
    g162_p,
    g161_n,
    g160_n
  );


  or

  (
    g162_n,
    g161_p,
    g160_p
  );


  and

  (
    g163_p,
    g162_p_spl_,
    G5_p_spl_0
  );


  or

  (
    g163_n,
    g162_n_spl_,
    G5_n_spl_0
  );


  and

  (
    g164_p,
    g162_n_spl_,
    G5_n_spl_1
  );


  or

  (
    g164_n,
    g162_p_spl_,
    G5_p_spl_1
  );


  and

  (
    g165_p,
    g164_n,
    g163_n
  );


  or

  (
    g165_n,
    g164_p,
    g163_p
  );


  and

  (
    g166_p,
    g165_n_spl_0,
    g64_n_spl_01
  );


  or

  (
    g166_n,
    g165_p_spl_0,
    g64_p_spl_01
  );


  and

  (
    g167_p,
    g165_p_spl_0,
    g64_p_spl_01
  );


  or

  (
    g167_n,
    g165_n_spl_0,
    g64_n_spl_01
  );


  and

  (
    g168_p,
    g167_n,
    g166_n
  );


  or

  (
    g168_n,
    g167_p,
    g166_p
  );


  and

  (
    g169_p,
    g168_p_spl_,
    g159_p_spl_
  );


  or

  (
    g169_n,
    g168_n_spl_,
    g159_n_spl_
  );


  and

  (
    g170_p,
    g168_n_spl_,
    g159_n_spl_
  );


  or

  (
    g170_n,
    g168_p_spl_,
    g159_p_spl_
  );


  and

  (
    g171_p,
    g170_n,
    g169_n
  );


  or

  (
    g171_n,
    g170_p,
    g169_p
  );


  and

  (
    g172_p,
    g171_n_spl_,
    G31_n_spl_011
  );


  or

  (
    g172_n,
    g171_p_spl_,
    G31_p_spl_011
  );


  and

  (
    g173_p,
    g172_n_spl_,
    G26_p_spl_0
  );


  or

  (
    g173_n,
    g172_p_spl_,
    G26_n_spl_0
  );


  and

  (
    g174_p,
    g108_n_spl_,
    G27_p_spl_
  );


  or

  (
    g174_n,
    g108_p_spl_,
    G27_n_spl_0
  );


  and

  (
    g175_p,
    g172_p_spl_,
    G26_n_spl_0
  );


  or

  (
    g175_n,
    g172_n_spl_,
    G26_p_spl_0
  );


  and

  (
    g176_p,
    g175_n,
    g174_n
  );


  or

  (
    g176_n,
    g175_p,
    g174_p
  );


  and

  (
    g177_p,
    g176_p,
    g173_n
  );


  or

  (
    g177_n,
    g176_n,
    g173_p
  );


  and

  (
    g178_p,
    g177_p,
    g154_p
  );


  or

  (
    g178_n,
    g177_n,
    g154_n
  );


  and

  (
    g179_p,
    G31_n_spl_011,
    G24_n_spl_1
  );


  or

  (
    g179_n,
    G31_p_spl_011,
    G24_p_spl_1
  );


  and

  (
    g180_p,
    g179_n_spl_,
    G18_p_spl_
  );


  or

  (
    g180_n,
    g179_p_spl_,
    G18_n_spl_
  );


  and

  (
    g181_p,
    G33_n_spl_011,
    G21_p_spl_
  );


  or

  (
    g181_n,
    G33_p_spl_10,
    G21_n_spl_
  );


  and

  (
    g182_p,
    g61_n_spl_1,
    G9_p_spl_0
  );


  or

  (
    g182_n,
    g61_p_spl_1,
    G9_n_spl_0
  );


  and

  (
    g183_p,
    g61_p_spl_1,
    G9_n_spl_1
  );


  or

  (
    g183_n,
    g61_n_spl_1,
    G9_p_spl_1
  );


  and

  (
    g184_p,
    g183_n,
    g182_n
  );


  or

  (
    g184_n,
    g183_p,
    g182_p
  );


  and

  (
    g185_p,
    g184_p_spl_,
    g181_p_spl_
  );


  or

  (
    g185_n,
    g184_n_spl_,
    g181_n_spl_
  );


  and

  (
    g186_p,
    g184_n_spl_,
    g181_n_spl_
  );


  or

  (
    g186_n,
    g184_p_spl_,
    g181_p_spl_
  );


  and

  (
    g187_p,
    g186_n,
    g185_n
  );


  or

  (
    g187_n,
    g186_p,
    g185_p
  );


  and

  (
    g188_p,
    g165_p_spl_1,
    g70_n_spl_1
  );


  or

  (
    g188_n,
    g165_n_spl_1,
    g70_p_spl_1
  );


  and

  (
    g189_p,
    g165_n_spl_1,
    g70_p_spl_1
  );


  or

  (
    g189_n,
    g165_p_spl_1,
    g70_n_spl_1
  );


  and

  (
    g190_p,
    g189_n,
    g188_n
  );


  or

  (
    g190_n,
    g189_p,
    g188_p
  );


  and

  (
    g191_p,
    G8_n_spl_10,
    G4_n_spl_10
  );


  or

  (
    g191_n,
    G8_p_spl_10,
    G4_p_spl_10
  );


  and

  (
    g192_p,
    G8_p_spl_10,
    G4_p_spl_10
  );


  or

  (
    g192_n,
    G8_n_spl_10,
    G4_n_spl_10
  );


  and

  (
    g193_p,
    g192_n,
    g191_n
  );


  or

  (
    g193_n,
    g192_p,
    g191_p
  );


  and

  (
    g194_p,
    g193_n_spl_,
    g190_p_spl_
  );


  or

  (
    g194_n,
    g193_p_spl_,
    g190_n_spl_
  );


  and

  (
    g195_p,
    g193_p_spl_,
    g190_n_spl_
  );


  or

  (
    g195_n,
    g193_n_spl_,
    g190_p_spl_
  );


  and

  (
    g196_p,
    g195_n,
    g194_n
  );


  or

  (
    g196_n,
    g195_p,
    g194_p
  );


  and

  (
    g197_p,
    g196_n_spl_0,
    g187_p_spl_
  );


  or

  (
    g197_n,
    g196_p_spl_0,
    g187_n_spl_
  );


  and

  (
    g198_p,
    g196_p_spl_0,
    g187_n_spl_
  );


  or

  (
    g198_n,
    g196_n_spl_0,
    g187_p_spl_
  );


  and

  (
    g199_p,
    g198_n,
    g197_n
  );


  or

  (
    g199_n,
    g198_p,
    g197_p
  );


  and

  (
    g200_p,
    g199_p_spl_,
    G31_n_spl_10
  );


  or

  (
    g200_n,
    g199_n_spl_,
    G31_p_spl_100
  );


  and

  (
    g201_p,
    g179_n_spl_,
    G17_p_spl_
  );


  or

  (
    g201_n,
    g179_p_spl_,
    G17_n_spl_
  );


  and

  (
    g202_p,
    g201_n_spl_0,
    g200_p_spl_
  );


  or

  (
    g202_n,
    g201_p_spl_0,
    g200_n_spl_
  );


  and

  (
    g203_p,
    g201_p_spl_0,
    g200_n_spl_
  );


  or

  (
    g203_n,
    g201_n_spl_0,
    g200_p_spl_
  );


  and

  (
    g204_p,
    g203_n,
    g202_n
  );


  or

  (
    g204_n,
    g203_p,
    g202_p
  );


  and

  (
    g205_p,
    g204_n_spl_0,
    g180_p_spl_0
  );


  or

  (
    g205_n,
    g204_p_spl_,
    g180_n_spl_
  );


  and

  (
    g206_p,
    g205_n,
    g178_p_spl_
  );


  or

  (
    g206_n,
    g205_p,
    g178_n_spl_0
  );


  and

  (
    g207_p,
    g206_p_spl_,
    g81_n_spl_
  );


  or

  (
    g207_n,
    g206_n_spl_,
    g81_p_spl_
  );


  and

  (
    g208_p,
    g207_p_spl_,
    g40_n_spl_
  );


  or

  (
    g208_n,
    g207_n_spl_,
    g40_p_spl_
  );


  and

  (
    g209_p,
    g208_n_spl_00,
    G1_p_spl_1
  );


  and

  (
    g210_p,
    g208_p_spl_00,
    G1_n_spl_1
  );


  or

  (
    g211_n,
    g210_p,
    g209_p
  );


  and

  (
    g212_p,
    g208_n_spl_00,
    G2_p_spl_1
  );


  and

  (
    g213_p,
    g208_p_spl_00,
    G2_n_spl_1
  );


  or

  (
    g214_n,
    g213_p,
    g212_p
  );


  and

  (
    g215_p,
    g208_n_spl_01,
    G3_p_spl_1
  );


  and

  (
    g216_p,
    g208_p_spl_01,
    G3_n_spl_1
  );


  or

  (
    g217_n,
    g216_p,
    g215_p
  );


  and

  (
    g218_p,
    g208_n_spl_01,
    G4_p_spl_1
  );


  and

  (
    g219_p,
    g208_p_spl_01,
    G4_n_spl_1
  );


  or

  (
    g220_n,
    g219_p,
    g218_p
  );


  and

  (
    g221_p,
    G33_n_spl_10,
    G30_n_spl_
  );


  or

  (
    g221_n,
    G33_p_spl_10,
    G30_p_spl_
  );


  and

  (
    g222_p,
    g221_p_spl_,
    g36_p_spl_
  );


  or

  (
    g222_n,
    g221_n_spl_,
    g36_n_spl_
  );


  and

  (
    g223_p,
    g222_n,
    g39_n_spl_
  );


  or

  (
    g223_n,
    g222_p,
    g39_p_spl_
  );


  and

  (
    g224_p,
    g223_n_spl_0,
    g207_p_spl_
  );


  or

  (
    g224_n,
    g223_p_spl_0,
    g207_n_spl_
  );


  and

  (
    g225_p,
    g224_n_spl_00,
    G10_p_spl_1
  );


  and

  (
    g226_p,
    g224_p_spl_00,
    G10_n_spl_1
  );


  or

  (
    g227_n,
    g226_p,
    g225_p
  );


  and

  (
    g228_p,
    g224_n_spl_00,
    G15_p_spl_1
  );


  and

  (
    g229_p,
    g224_p_spl_00,
    G15_n_spl_1
  );


  or

  (
    g230_n,
    g229_p,
    g228_p
  );


  and

  (
    g231_p,
    g224_n_spl_01,
    G16_p_spl_1
  );


  and

  (
    g232_p,
    g224_p_spl_01,
    G16_n_spl_1
  );


  or

  (
    g233_n,
    g232_p,
    g231_p
  );


  and

  (
    g234_p,
    g80_p_spl_,
    g42_p_spl_0
  );


  or

  (
    g234_n,
    g80_n_spl_0,
    g42_n_spl_
  );


  and

  (
    g235_p,
    g234_p,
    g206_p_spl_
  );


  or

  (
    g235_n,
    g234_n,
    g206_n_spl_
  );


  and

  (
    g236_p,
    g235_p_spl_,
    g40_n_spl_
  );


  or

  (
    g236_n,
    g235_n_spl_,
    g40_p_spl_
  );


  and

  (
    g237_p,
    g236_n_spl_0,
    G5_p_spl_1
  );


  and

  (
    g238_p,
    g236_p_spl_0,
    G5_n_spl_1
  );


  or

  (
    g239_n,
    g238_p,
    g237_p
  );


  and

  (
    g240_p,
    g236_n_spl_0,
    G6_p_spl_1
  );


  and

  (
    g241_p,
    g236_p_spl_0,
    G6_n_spl_1
  );


  or

  (
    g242_n,
    g241_p,
    g240_p
  );


  and

  (
    g243_p,
    g236_n_spl_1,
    G7_p_spl_1
  );


  and

  (
    g244_p,
    g236_p_spl_1,
    G7_n_spl_1
  );


  or

  (
    g245_n,
    g244_p,
    g243_p
  );


  and

  (
    g246_p,
    g236_n_spl_1,
    G8_p_spl_1
  );


  and

  (
    g247_p,
    g236_p_spl_1,
    G8_n_spl_1
  );


  or

  (
    g248_n,
    g247_p,
    g246_p
  );


  and

  (
    g249_p,
    g235_p_spl_,
    g223_n_spl_0
  );


  or

  (
    g249_n,
    g235_n_spl_,
    g223_p_spl_0
  );


  or

  (
    g250_n,
    g249_n,
    G9_n_spl_1
  );


  or

  (
    g251_n,
    g249_p,
    G9_p_spl_1
  );


  and

  (
    g252_p,
    g251_n,
    g250_n
  );


  and

  (
    g253_p,
    g180_p_spl_0,
    g178_p_spl_
  );


  or

  (
    g253_n,
    g180_n_spl_,
    g178_n_spl_0
  );


  and

  (
    g254_p,
    g223_n_spl_,
    g81_n_spl_
  );


  or

  (
    g254_n,
    g223_p_spl_,
    g81_p_spl_
  );


  and

  (
    g255_p,
    g254_p,
    g204_p_spl_
  );


  or

  (
    g255_n,
    g254_n,
    g204_n_spl_0
  );


  and

  (
    g256_p,
    g255_p,
    g253_p
  );


  or

  (
    g256_n,
    g255_n,
    g253_n
  );


  and

  (
    g257_p,
    g256_n_spl_0,
    G11_p_spl_1
  );


  and

  (
    g258_p,
    g256_p_spl_0,
    G11_n_spl_1
  );


  or

  (
    g259_n,
    g258_p,
    g257_p
  );


  and

  (
    g260_p,
    g256_n_spl_0,
    G12_p_spl_1
  );


  and

  (
    g261_p,
    g256_p_spl_0,
    G12_n_spl_1
  );


  or

  (
    g262_n,
    g261_p,
    g260_p
  );


  and

  (
    g263_p,
    g256_n_spl_1,
    G13_p_spl_1
  );


  and

  (
    g264_p,
    g256_p_spl_1,
    G13_n_spl_1
  );


  or

  (
    g265_n,
    g264_p,
    g263_p
  );


  and

  (
    g266_p,
    g256_n_spl_1,
    G14_p_spl_1
  );


  and

  (
    g267_p,
    g256_p_spl_1,
    G14_n_spl_1
  );


  or

  (
    g268_n,
    g267_p,
    g266_p
  );


  and

  (
    g269_p,
    g224_n_spl_01,
    g208_n_spl_10
  );


  or

  (
    g269_n,
    g224_p_spl_01,
    g208_p_spl_10
  );


  or

  (
    g270_n,
    g269_p_spl_00,
    G32_n_spl_
  );


  or

  (
    g271_n,
    g204_n_spl_,
    g80_n_spl_
  );


  or

  (
    g272_n,
    g180_p_spl_,
    g42_p_spl_
  );


  or

  (
    g273_n,
    g272_n,
    g178_n_spl_
  );


  or

  (
    g274_n,
    g273_n,
    g271_n
  );


  and

  (
    g275_p,
    g274_n,
    g270_n
  );


  and

  (
    g276_p,
    g275_p,
    G33_n_spl_10
  );


  and

  (
    g277_p,
    g201_p_spl_,
    G31_n_spl_10
  );


  or

  (
    g277_n,
    g201_n_spl_,
    G31_p_spl_100
  );


  and

  (
    g278_p,
    g277_p,
    g269_n_spl_0
  );


  or

  (
    g278_n,
    g277_n,
    g269_p_spl_00
  );


  or

  (
    g279_n,
    g278_p,
    g199_n_spl_
  );


  or

  (
    g280_n,
    g278_n,
    g199_p_spl_
  );


  and

  (
    g281_p,
    g280_n,
    g279_n
  );


  or

  (
    g282_n,
    g281_p,
    g38_p_spl_00
  );


  and

  (
    g283_p,
    G31_n_spl_11,
    G25_p_spl_
  );


  or

  (
    g283_n,
    G31_p_spl_101,
    G25_n_spl_
  );


  and

  (
    g284_p,
    g283_p,
    g269_n_spl_0
  );


  or

  (
    g284_n,
    g283_n,
    g269_p_spl_01
  );


  or

  (
    g285_n,
    g284_p,
    g76_p_spl_
  );


  or

  (
    g286_n,
    g284_n,
    g76_n_spl_
  );


  and

  (
    g287_p,
    g286_n,
    g285_n
  );


  or

  (
    g288_n,
    g287_p,
    g38_p_spl_01
  );


  or

  (
    g289_n,
    G31_p_spl_101,
    G27_n_spl_
  );


  or

  (
    g290_n,
    g289_n,
    g269_p_spl_01
  );


  and

  (
    g291_p,
    g290_n,
    g107_n_spl_
  );


  or

  (
    g292_n,
    g291_p,
    g38_p_spl_01
  );


  or

  (
    g293_n,
    G31_p_spl_110,
    G28_n_spl_
  );


  or

  (
    g294_n,
    g293_n,
    g269_p_spl_10
  );


  and

  (
    g295_p,
    g294_n,
    g126_n_spl_
  );


  or

  (
    g296_n,
    g295_p,
    g38_p_spl_10
  );


  or

  (
    g297_n,
    g149_n_spl_,
    G31_p_spl_110
  );


  or

  (
    g298_n,
    g297_n,
    g269_p_spl_10
  );


  and

  (
    g299_p,
    g298_n,
    g147_n_spl_
  );


  or

  (
    g300_n,
    g299_p,
    g38_p_spl_10
  );


  and

  (
    g301_p,
    G29_p_spl_,
    G21_p_spl_
  );


  or

  (
    g301_n,
    G29_n_spl_,
    G21_n_spl_
  );


  and

  (
    g302_p,
    g301_n,
    G33_n_spl_11
  );


  or

  (
    g302_n,
    g301_p,
    G33_p_spl_11
  );


  and

  (
    g303_p,
    g196_p_spl_,
    g34_n_spl_
  );


  or

  (
    g303_n,
    g196_n_spl_,
    g34_p_spl_
  );


  and

  (
    g304_p,
    g303_n_spl_,
    g208_n_spl_10
  );


  or

  (
    g304_n,
    g303_p_spl_,
    g208_p_spl_10
  );


  and

  (
    g305_p,
    g303_p_spl_,
    g208_p_spl_1
  );


  or

  (
    g305_n,
    g303_n_spl_,
    g208_n_spl_1
  );


  and

  (
    g306_p,
    g305_n,
    g304_n
  );


  or

  (
    g306_n,
    g305_p,
    g304_p
  );


  or

  (
    g307_n,
    g306_n,
    g302_p
  );


  or

  (
    g308_n,
    g306_p,
    g302_n
  );


  and

  (
    g309_p,
    g308_n,
    g307_n
  );


  and

  (
    g310_p,
    G30_p_spl_,
    G22_p_spl_
  );


  or

  (
    g310_n,
    G30_n_spl_,
    G22_n_spl_
  );


  and

  (
    g311_p,
    g310_n,
    G33_n_spl_11
  );


  or

  (
    g311_n,
    g310_p,
    G33_p_spl_11
  );


  and

  (
    g312_p,
    g92_n_spl_1,
    g64_p_spl_1
  );


  or

  (
    g312_n,
    g92_p_spl_1,
    g64_n_spl_1
  );


  and

  (
    g313_p,
    g92_p_spl_1,
    g64_n_spl_1
  );


  or

  (
    g313_n,
    g92_n_spl_1,
    g64_p_spl_1
  );


  and

  (
    g314_p,
    g313_n,
    g312_n
  );


  or

  (
    g314_n,
    g313_p,
    g312_p
  );


  and

  (
    g315_p,
    g314_n,
    g221_n_spl_
  );


  or

  (
    g315_n,
    g314_p,
    g221_p_spl_
  );


  and

  (
    g316_p,
    g315_n_spl_,
    g224_n_spl_1
  );


  or

  (
    g316_n,
    g315_p_spl_,
    g224_p_spl_1
  );


  and

  (
    g317_p,
    g315_p_spl_,
    g224_p_spl_1
  );


  or

  (
    g317_n,
    g315_n_spl_,
    g224_n_spl_1
  );


  and

  (
    g318_p,
    g317_n,
    g316_n
  );


  or

  (
    g318_n,
    g317_p,
    g316_p
  );


  or

  (
    g319_n,
    g318_n,
    g311_p
  );


  or

  (
    g320_n,
    g318_p,
    g311_n
  );


  and

  (
    g321_p,
    g320_n,
    g319_n
  );


  and

  (
    g322_p,
    G31_n_spl_11,
    G26_p_spl_
  );


  or

  (
    g322_n,
    G31_p_spl_11,
    G26_n_spl_
  );


  and

  (
    g323_p,
    g322_p,
    g269_n_spl_
  );


  or

  (
    g323_n,
    g322_n,
    g269_p_spl_1
  );


  or

  (
    g324_n,
    g323_p,
    g171_p_spl_
  );


  or

  (
    g325_n,
    g323_n,
    g171_n_spl_
  );


  and

  (
    g326_p,
    g325_n,
    g324_n
  );


  or

  (
    g327_n,
    g326_p,
    g38_p_spl_1
  );


  not

  (
    G1884,
    g211_n
  );


  not

  (
    G1885,
    g214_n
  );


  not

  (
    G1886,
    g217_n
  );


  not

  (
    G1887,
    g220_n
  );


  not

  (
    G1888,
    g227_n
  );


  not

  (
    G1889,
    g230_n
  );


  not

  (
    G1890,
    g233_n
  );


  not

  (
    G1891,
    g239_n
  );


  not

  (
    G1892,
    g242_n
  );


  not

  (
    G1893,
    g245_n
  );


  not

  (
    G1894,
    g248_n
  );


  not

  (
    G1895,
    g252_p
  );


  not

  (
    G1896,
    g259_n
  );


  not

  (
    G1897,
    g262_n
  );


  not

  (
    G1898,
    g265_n
  );


  not

  (
    G1899,
    g268_n
  );


  not

  (
    G1900,
    g276_p
  );


  not

  (
    G1901,
    g282_n
  );


  not

  (
    G1902,
    g288_n
  );


  not

  (
    G1903,
    g292_n
  );


  not

  (
    G1904,
    g296_n
  );


  not

  (
    G1905,
    g300_n
  );


  not

  (
    G1906,
    g309_p
  );


  not

  (
    G1907,
    g321_p
  );


  not

  (
    G1908,
    g327_n
  );


  buf

  (
    G33_n_spl_,
    G33_n
  );


  buf

  (
    G33_n_spl_0,
    G33_n_spl_
  );


  buf

  (
    G33_n_spl_00,
    G33_n_spl_0
  );


  buf

  (
    G33_n_spl_000,
    G33_n_spl_00
  );


  buf

  (
    G33_n_spl_001,
    G33_n_spl_00
  );


  buf

  (
    G33_n_spl_01,
    G33_n_spl_0
  );


  buf

  (
    G33_n_spl_010,
    G33_n_spl_01
  );


  buf

  (
    G33_n_spl_011,
    G33_n_spl_01
  );


  buf

  (
    G33_n_spl_1,
    G33_n_spl_
  );


  buf

  (
    G33_n_spl_10,
    G33_n_spl_1
  );


  buf

  (
    G33_n_spl_11,
    G33_n_spl_1
  );


  buf

  (
    G29_n_spl_,
    G29_n
  );


  buf

  (
    G33_p_spl_,
    G33_p
  );


  buf

  (
    G33_p_spl_0,
    G33_p_spl_
  );


  buf

  (
    G33_p_spl_00,
    G33_p_spl_0
  );


  buf

  (
    G33_p_spl_000,
    G33_p_spl_00
  );


  buf

  (
    G33_p_spl_001,
    G33_p_spl_00
  );


  buf

  (
    G33_p_spl_01,
    G33_p_spl_0
  );


  buf

  (
    G33_p_spl_010,
    G33_p_spl_01
  );


  buf

  (
    G33_p_spl_1,
    G33_p_spl_
  );


  buf

  (
    G33_p_spl_10,
    G33_p_spl_1
  );


  buf

  (
    G33_p_spl_11,
    G33_p_spl_1
  );


  buf

  (
    G29_p_spl_,
    G29_p
  );


  buf

  (
    G24_p_spl_,
    G24_p
  );


  buf

  (
    G24_p_spl_0,
    G24_p_spl_
  );


  buf

  (
    G24_p_spl_1,
    G24_p_spl_
  );


  buf

  (
    G23_n_spl_,
    G23_n
  );


  buf

  (
    G23_n_spl_0,
    G23_n_spl_
  );


  buf

  (
    G23_n_spl_1,
    G23_n_spl_
  );


  buf

  (
    G24_n_spl_,
    G24_n
  );


  buf

  (
    G24_n_spl_0,
    G24_n_spl_
  );


  buf

  (
    G24_n_spl_1,
    G24_n_spl_
  );


  buf

  (
    G23_p_spl_,
    G23_p
  );


  buf

  (
    G23_p_spl_0,
    G23_p_spl_
  );


  buf

  (
    G23_p_spl_1,
    G23_p_spl_
  );


  buf

  (
    g35_n_spl_,
    g35_n
  );


  buf

  (
    G31_n_spl_,
    G31_n
  );


  buf

  (
    G31_n_spl_0,
    G31_n_spl_
  );


  buf

  (
    G31_n_spl_00,
    G31_n_spl_0
  );


  buf

  (
    G31_n_spl_000,
    G31_n_spl_00
  );


  buf

  (
    G31_n_spl_001,
    G31_n_spl_00
  );


  buf

  (
    G31_n_spl_01,
    G31_n_spl_0
  );


  buf

  (
    G31_n_spl_010,
    G31_n_spl_01
  );


  buf

  (
    G31_n_spl_011,
    G31_n_spl_01
  );


  buf

  (
    G31_n_spl_1,
    G31_n_spl_
  );


  buf

  (
    G31_n_spl_10,
    G31_n_spl_1
  );


  buf

  (
    G31_n_spl_11,
    G31_n_spl_1
  );


  buf

  (
    g35_p_spl_,
    g35_p
  );


  buf

  (
    G31_p_spl_,
    G31_p
  );


  buf

  (
    G31_p_spl_0,
    G31_p_spl_
  );


  buf

  (
    G31_p_spl_00,
    G31_p_spl_0
  );


  buf

  (
    G31_p_spl_000,
    G31_p_spl_00
  );


  buf

  (
    G31_p_spl_001,
    G31_p_spl_00
  );


  buf

  (
    G31_p_spl_01,
    G31_p_spl_0
  );


  buf

  (
    G31_p_spl_010,
    G31_p_spl_01
  );


  buf

  (
    G31_p_spl_011,
    G31_p_spl_01
  );


  buf

  (
    G31_p_spl_1,
    G31_p_spl_
  );


  buf

  (
    G31_p_spl_10,
    G31_p_spl_1
  );


  buf

  (
    G31_p_spl_100,
    G31_p_spl_10
  );


  buf

  (
    G31_p_spl_101,
    G31_p_spl_10
  );


  buf

  (
    G31_p_spl_11,
    G31_p_spl_1
  );


  buf

  (
    G31_p_spl_110,
    G31_p_spl_11
  );


  buf

  (
    g36_p_spl_,
    g36_p
  );


  buf

  (
    g34_p_spl_,
    g34_p
  );


  buf

  (
    g36_n_spl_,
    g36_n
  );


  buf

  (
    g34_n_spl_,
    g34_n
  );


  buf

  (
    G32_n_spl_,
    G32_n
  );


  buf

  (
    g38_p_spl_,
    g38_p
  );


  buf

  (
    g38_p_spl_0,
    g38_p_spl_
  );


  buf

  (
    g38_p_spl_00,
    g38_p_spl_0
  );


  buf

  (
    g38_p_spl_01,
    g38_p_spl_0
  );


  buf

  (
    g38_p_spl_1,
    g38_p_spl_
  );


  buf

  (
    g38_p_spl_10,
    g38_p_spl_1
  );


  buf

  (
    g39_n_spl_,
    g39_n
  );


  buf

  (
    g39_p_spl_,
    g39_p
  );


  buf

  (
    g41_n_spl_,
    g41_n
  );


  buf

  (
    G20_p_spl_,
    G20_p
  );


  buf

  (
    g41_p_spl_,
    g41_p
  );


  buf

  (
    G20_n_spl_,
    G20_n
  );


  buf

  (
    G22_p_spl_,
    G22_p
  );


  buf

  (
    G22_n_spl_,
    G22_n
  );


  buf

  (
    G14_n_spl_,
    G14_n
  );


  buf

  (
    G14_n_spl_0,
    G14_n_spl_
  );


  buf

  (
    G14_n_spl_00,
    G14_n_spl_0
  );


  buf

  (
    G14_n_spl_1,
    G14_n_spl_
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_00,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_01,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_10,
    G4_p_spl_1
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G14_p_spl_0,
    G14_p_spl_
  );


  buf

  (
    G14_p_spl_00,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_1,
    G14_p_spl_
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    G4_n_spl_0,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_00,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_01,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_1,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_10,
    G4_n_spl_1
  );


  buf

  (
    g46_p_spl_,
    g46_p
  );


  buf

  (
    g43_p_spl_,
    g43_p
  );


  buf

  (
    g46_n_spl_,
    g46_n
  );


  buf

  (
    g43_n_spl_,
    g43_n
  );


  buf

  (
    G13_n_spl_,
    G13_n
  );


  buf

  (
    G13_n_spl_0,
    G13_n_spl_
  );


  buf

  (
    G13_n_spl_00,
    G13_n_spl_0
  );


  buf

  (
    G13_n_spl_1,
    G13_n_spl_
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_00,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_1,
    G12_p_spl_
  );


  buf

  (
    G13_p_spl_,
    G13_p
  );


  buf

  (
    G13_p_spl_0,
    G13_p_spl_
  );


  buf

  (
    G13_p_spl_00,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_1,
    G13_p_spl_
  );


  buf

  (
    G12_n_spl_,
    G12_n
  );


  buf

  (
    G12_n_spl_0,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_00,
    G12_n_spl_0
  );


  buf

  (
    G12_n_spl_1,
    G12_n_spl_
  );


  buf

  (
    g52_p_spl_,
    g52_p
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    G11_p_spl_0,
    G11_p_spl_
  );


  buf

  (
    G11_p_spl_00,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_1,
    G11_p_spl_
  );


  buf

  (
    g52_n_spl_,
    g52_n
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    G11_n_spl_0,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_00,
    G11_n_spl_0
  );


  buf

  (
    G11_n_spl_1,
    G11_n_spl_
  );


  buf

  (
    G15_n_spl_,
    G15_n
  );


  buf

  (
    G15_n_spl_0,
    G15_n_spl_
  );


  buf

  (
    G15_n_spl_00,
    G15_n_spl_0
  );


  buf

  (
    G15_n_spl_1,
    G15_n_spl_
  );


  buf

  (
    G10_n_spl_,
    G10_n
  );


  buf

  (
    G10_n_spl_0,
    G10_n_spl_
  );


  buf

  (
    G10_n_spl_00,
    G10_n_spl_0
  );


  buf

  (
    G10_n_spl_1,
    G10_n_spl_
  );


  buf

  (
    G15_p_spl_,
    G15_p
  );


  buf

  (
    G15_p_spl_0,
    G15_p_spl_
  );


  buf

  (
    G15_p_spl_00,
    G15_p_spl_0
  );


  buf

  (
    G15_p_spl_1,
    G15_p_spl_
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


  buf

  (
    G10_p_spl_0,
    G10_p_spl_
  );


  buf

  (
    G10_p_spl_00,
    G10_p_spl_0
  );


  buf

  (
    G10_p_spl_1,
    G10_p_spl_
  );


  buf

  (
    g58_n_spl_,
    g58_n
  );


  buf

  (
    g58_n_spl_0,
    g58_n_spl_
  );


  buf

  (
    g58_n_spl_1,
    g58_n_spl_
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    G16_p_spl_0,
    G16_p_spl_
  );


  buf

  (
    G16_p_spl_00,
    G16_p_spl_0
  );


  buf

  (
    G16_p_spl_1,
    G16_p_spl_
  );


  buf

  (
    g58_p_spl_,
    g58_p
  );


  buf

  (
    g58_p_spl_0,
    g58_p_spl_
  );


  buf

  (
    g58_p_spl_1,
    g58_p_spl_
  );


  buf

  (
    G16_n_spl_,
    G16_n
  );


  buf

  (
    G16_n_spl_0,
    G16_n_spl_
  );


  buf

  (
    G16_n_spl_00,
    G16_n_spl_0
  );


  buf

  (
    G16_n_spl_1,
    G16_n_spl_
  );


  buf

  (
    g61_p_spl_,
    g61_p
  );


  buf

  (
    g61_p_spl_0,
    g61_p_spl_
  );


  buf

  (
    g61_p_spl_1,
    g61_p_spl_
  );


  buf

  (
    g55_n_spl_,
    g55_n
  );


  buf

  (
    g61_n_spl_,
    g61_n
  );


  buf

  (
    g61_n_spl_0,
    g61_n_spl_
  );


  buf

  (
    g61_n_spl_1,
    g61_n_spl_
  );


  buf

  (
    g55_p_spl_,
    g55_p
  );


  buf

  (
    G3_n_spl_,
    G3_n
  );


  buf

  (
    G3_n_spl_0,
    G3_n_spl_
  );


  buf

  (
    G3_n_spl_00,
    G3_n_spl_0
  );


  buf

  (
    G3_n_spl_1,
    G3_n_spl_
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G2_p_spl_0,
    G2_p_spl_
  );


  buf

  (
    G2_p_spl_00,
    G2_p_spl_0
  );


  buf

  (
    G2_p_spl_1,
    G2_p_spl_
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G3_p_spl_0,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_00,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_1,
    G3_p_spl_
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G2_n_spl_0,
    G2_n_spl_
  );


  buf

  (
    G2_n_spl_00,
    G2_n_spl_0
  );


  buf

  (
    G2_n_spl_1,
    G2_n_spl_
  );


  buf

  (
    g67_p_spl_,
    g67_p
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G1_p_spl_0,
    G1_p_spl_
  );


  buf

  (
    G1_p_spl_00,
    G1_p_spl_0
  );


  buf

  (
    G1_p_spl_1,
    G1_p_spl_
  );


  buf

  (
    g67_n_spl_,
    g67_n
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    G1_n_spl_00,
    G1_n_spl_0
  );


  buf

  (
    G1_n_spl_1,
    G1_n_spl_
  );


  buf

  (
    g70_n_spl_,
    g70_n
  );


  buf

  (
    g70_n_spl_0,
    g70_n_spl_
  );


  buf

  (
    g70_n_spl_1,
    g70_n_spl_
  );


  buf

  (
    g64_n_spl_,
    g64_n
  );


  buf

  (
    g64_n_spl_0,
    g64_n_spl_
  );


  buf

  (
    g64_n_spl_00,
    g64_n_spl_0
  );


  buf

  (
    g64_n_spl_01,
    g64_n_spl_0
  );


  buf

  (
    g64_n_spl_1,
    g64_n_spl_
  );


  buf

  (
    g70_p_spl_,
    g70_p
  );


  buf

  (
    g70_p_spl_0,
    g70_p_spl_
  );


  buf

  (
    g70_p_spl_1,
    g70_p_spl_
  );


  buf

  (
    g64_p_spl_,
    g64_p
  );


  buf

  (
    g64_p_spl_0,
    g64_p_spl_
  );


  buf

  (
    g64_p_spl_00,
    g64_p_spl_0
  );


  buf

  (
    g64_p_spl_01,
    g64_p_spl_0
  );


  buf

  (
    g64_p_spl_1,
    g64_p_spl_
  );


  buf

  (
    g73_n_spl_,
    g73_n
  );


  buf

  (
    g49_n_spl_,
    g49_n
  );


  buf

  (
    g73_p_spl_,
    g73_p
  );


  buf

  (
    g49_p_spl_,
    g49_p
  );


  buf

  (
    g76_n_spl_,
    g76_n
  );


  buf

  (
    g76_p_spl_,
    g76_p
  );


  buf

  (
    g77_p_spl_,
    g77_p
  );


  buf

  (
    G25_n_spl_,
    G25_n
  );


  buf

  (
    G25_n_spl_0,
    G25_n_spl_
  );


  buf

  (
    g77_n_spl_,
    g77_n
  );


  buf

  (
    G25_p_spl_,
    G25_p
  );


  buf

  (
    G25_p_spl_0,
    G25_p_spl_
  );


  buf

  (
    g80_n_spl_,
    g80_n
  );


  buf

  (
    g80_n_spl_0,
    g80_n_spl_
  );


  buf

  (
    g42_p_spl_,
    g42_p
  );


  buf

  (
    g42_p_spl_0,
    g42_p_spl_
  );


  buf

  (
    g80_p_spl_,
    g80_p
  );


  buf

  (
    g42_n_spl_,
    g42_n
  );


  buf

  (
    G18_p_spl_,
    G18_p
  );


  buf

  (
    G18_n_spl_,
    G18_n
  );


  buf

  (
    g83_n_spl_,
    g83_n
  );


  buf

  (
    g83_p_spl_,
    g83_p
  );


  buf

  (
    g86_n_spl_,
    g86_n
  );


  buf

  (
    g86_p_spl_,
    g86_p
  );


  buf

  (
    G9_p_spl_,
    G9_p
  );


  buf

  (
    G9_p_spl_0,
    G9_p_spl_
  );


  buf

  (
    G9_p_spl_00,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_1,
    G9_p_spl_
  );


  buf

  (
    G9_n_spl_,
    G9_n
  );


  buf

  (
    G9_n_spl_0,
    G9_n_spl_
  );


  buf

  (
    G9_n_spl_00,
    G9_n_spl_0
  );


  buf

  (
    G9_n_spl_1,
    G9_n_spl_
  );


  buf

  (
    g92_n_spl_,
    g92_n
  );


  buf

  (
    g92_n_spl_0,
    g92_n_spl_
  );


  buf

  (
    g92_n_spl_1,
    g92_n_spl_
  );


  buf

  (
    g92_p_spl_,
    g92_p
  );


  buf

  (
    g92_p_spl_0,
    g92_p_spl_
  );


  buf

  (
    g92_p_spl_1,
    g92_p_spl_
  );


  buf

  (
    g95_p_spl_,
    g95_p
  );


  buf

  (
    g95_p_spl_0,
    g95_p_spl_
  );


  buf

  (
    g95_p_spl_1,
    g95_p_spl_
  );


  buf

  (
    g89_p_spl_,
    g89_p
  );


  buf

  (
    g95_n_spl_,
    g95_n
  );


  buf

  (
    g95_n_spl_0,
    g95_n_spl_
  );


  buf

  (
    g95_n_spl_1,
    g95_n_spl_
  );


  buf

  (
    g89_n_spl_,
    g89_n
  );


  buf

  (
    G8_n_spl_,
    G8_n
  );


  buf

  (
    G8_n_spl_0,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_00,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_01,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_1,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_10,
    G8_n_spl_1
  );


  buf

  (
    G5_n_spl_,
    G5_n
  );


  buf

  (
    G5_n_spl_0,
    G5_n_spl_
  );


  buf

  (
    G5_n_spl_00,
    G5_n_spl_0
  );


  buf

  (
    G5_n_spl_1,
    G5_n_spl_
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_00,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_01,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_1,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_10,
    G8_p_spl_1
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G5_p_spl_0,
    G5_p_spl_
  );


  buf

  (
    G5_p_spl_00,
    G5_p_spl_0
  );


  buf

  (
    G5_p_spl_1,
    G5_p_spl_
  );


  buf

  (
    g101_p_spl_,
    g101_p
  );


  buf

  (
    g101_n_spl_,
    g101_n
  );


  buf

  (
    g104_p_spl_,
    g104_p
  );


  buf

  (
    g98_n_spl_,
    g98_n
  );


  buf

  (
    g104_n_spl_,
    g104_n
  );


  buf

  (
    g98_p_spl_,
    g98_p
  );


  buf

  (
    g107_n_spl_,
    g107_n
  );


  buf

  (
    g108_p_spl_,
    g108_p
  );


  buf

  (
    G27_n_spl_,
    G27_n
  );


  buf

  (
    G27_n_spl_0,
    G27_n_spl_
  );


  buf

  (
    g108_n_spl_,
    g108_n
  );


  buf

  (
    G27_p_spl_,
    G27_p
  );


  buf

  (
    G6_n_spl_,
    G6_n
  );


  buf

  (
    G6_n_spl_0,
    G6_n_spl_
  );


  buf

  (
    G6_n_spl_00,
    G6_n_spl_0
  );


  buf

  (
    G6_n_spl_1,
    G6_n_spl_
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G6_p_spl_0,
    G6_p_spl_
  );


  buf

  (
    G6_p_spl_00,
    G6_p_spl_0
  );


  buf

  (
    G6_p_spl_1,
    G6_p_spl_
  );


  buf

  (
    g112_p_spl_,
    g112_p
  );


  buf

  (
    g112_n_spl_,
    g112_n
  );


  buf

  (
    g118_n_spl_,
    g118_n
  );


  buf

  (
    g115_n_spl_,
    g115_n
  );


  buf

  (
    g118_p_spl_,
    g118_p
  );


  buf

  (
    g115_p_spl_,
    g115_p
  );


  buf

  (
    G19_p_spl_,
    G19_p
  );


  buf

  (
    G19_n_spl_,
    G19_n
  );


  buf

  (
    g123_n_spl_,
    g123_n
  );


  buf

  (
    g121_n_spl_,
    g121_n
  );


  buf

  (
    g123_p_spl_,
    g123_p
  );


  buf

  (
    g121_p_spl_,
    g121_p
  );


  buf

  (
    g126_n_spl_,
    g126_n
  );


  buf

  (
    g127_p_spl_,
    g127_p
  );


  buf

  (
    G28_n_spl_,
    G28_n
  );


  buf

  (
    G28_n_spl_0,
    G28_n_spl_
  );


  buf

  (
    g127_n_spl_,
    g127_n
  );


  buf

  (
    G28_p_spl_,
    G28_p
  );


  buf

  (
    G7_n_spl_,
    G7_n
  );


  buf

  (
    G7_n_spl_0,
    G7_n_spl_
  );


  buf

  (
    G7_n_spl_00,
    G7_n_spl_0
  );


  buf

  (
    G7_n_spl_1,
    G7_n_spl_
  );


  buf

  (
    G7_p_spl_,
    G7_p
  );


  buf

  (
    G7_p_spl_0,
    G7_p_spl_
  );


  buf

  (
    G7_p_spl_00,
    G7_p_spl_0
  );


  buf

  (
    G7_p_spl_1,
    G7_p_spl_
  );


  buf

  (
    g133_p_spl_,
    g133_p
  );


  buf

  (
    g133_n_spl_,
    g133_n
  );


  buf

  (
    g136_n_spl_,
    g136_n
  );


  buf

  (
    g136_p_spl_,
    g136_p
  );


  buf

  (
    g141_p_spl_,
    g141_p
  );


  buf

  (
    g141_n_spl_,
    g141_n
  );


  buf

  (
    g144_n_spl_,
    g144_n
  );


  buf

  (
    g139_n_spl_,
    g139_n
  );


  buf

  (
    g144_p_spl_,
    g144_p
  );


  buf

  (
    g139_p_spl_,
    g139_p
  );


  buf

  (
    g147_n_spl_,
    g147_n
  );


  buf

  (
    g149_n_spl_,
    g149_n
  );


  buf

  (
    g149_n_spl_0,
    g149_n_spl_
  );


  buf

  (
    g148_p_spl_,
    g148_p
  );


  buf

  (
    g149_p_spl_,
    g149_p
  );


  buf

  (
    g148_n_spl_,
    g148_n
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    G17_n_spl_,
    G17_n
  );


  buf

  (
    g156_p_spl_,
    g156_p
  );


  buf

  (
    g156_n_spl_,
    g156_n
  );


  buf

  (
    g162_p_spl_,
    g162_p
  );


  buf

  (
    g162_n_spl_,
    g162_n
  );


  buf

  (
    g165_n_spl_,
    g165_n
  );


  buf

  (
    g165_n_spl_0,
    g165_n_spl_
  );


  buf

  (
    g165_n_spl_1,
    g165_n_spl_
  );


  buf

  (
    g165_p_spl_,
    g165_p
  );


  buf

  (
    g165_p_spl_0,
    g165_p_spl_
  );


  buf

  (
    g165_p_spl_1,
    g165_p_spl_
  );


  buf

  (
    g168_p_spl_,
    g168_p
  );


  buf

  (
    g159_p_spl_,
    g159_p
  );


  buf

  (
    g168_n_spl_,
    g168_n
  );


  buf

  (
    g159_n_spl_,
    g159_n
  );


  buf

  (
    g171_n_spl_,
    g171_n
  );


  buf

  (
    g171_p_spl_,
    g171_p
  );


  buf

  (
    g172_n_spl_,
    g172_n
  );


  buf

  (
    G26_p_spl_,
    G26_p
  );


  buf

  (
    G26_p_spl_0,
    G26_p_spl_
  );


  buf

  (
    g172_p_spl_,
    g172_p
  );


  buf

  (
    G26_n_spl_,
    G26_n
  );


  buf

  (
    G26_n_spl_0,
    G26_n_spl_
  );


  buf

  (
    g179_n_spl_,
    g179_n
  );


  buf

  (
    g179_p_spl_,
    g179_p
  );


  buf

  (
    G21_p_spl_,
    G21_p
  );


  buf

  (
    G21_n_spl_,
    G21_n
  );


  buf

  (
    g184_p_spl_,
    g184_p
  );


  buf

  (
    g181_p_spl_,
    g181_p
  );


  buf

  (
    g184_n_spl_,
    g184_n
  );


  buf

  (
    g181_n_spl_,
    g181_n
  );


  buf

  (
    g193_n_spl_,
    g193_n
  );


  buf

  (
    g190_p_spl_,
    g190_p
  );


  buf

  (
    g193_p_spl_,
    g193_p
  );


  buf

  (
    g190_n_spl_,
    g190_n
  );


  buf

  (
    g196_n_spl_,
    g196_n
  );


  buf

  (
    g196_n_spl_0,
    g196_n_spl_
  );


  buf

  (
    g187_p_spl_,
    g187_p
  );


  buf

  (
    g196_p_spl_,
    g196_p
  );


  buf

  (
    g196_p_spl_0,
    g196_p_spl_
  );


  buf

  (
    g187_n_spl_,
    g187_n
  );


  buf

  (
    g199_p_spl_,
    g199_p
  );


  buf

  (
    g199_n_spl_,
    g199_n
  );


  buf

  (
    g201_n_spl_,
    g201_n
  );


  buf

  (
    g201_n_spl_0,
    g201_n_spl_
  );


  buf

  (
    g200_p_spl_,
    g200_p
  );


  buf

  (
    g201_p_spl_,
    g201_p
  );


  buf

  (
    g201_p_spl_0,
    g201_p_spl_
  );


  buf

  (
    g200_n_spl_,
    g200_n
  );


  buf

  (
    g204_n_spl_,
    g204_n
  );


  buf

  (
    g204_n_spl_0,
    g204_n_spl_
  );


  buf

  (
    g180_p_spl_,
    g180_p
  );


  buf

  (
    g180_p_spl_0,
    g180_p_spl_
  );


  buf

  (
    g204_p_spl_,
    g204_p
  );


  buf

  (
    g180_n_spl_,
    g180_n
  );


  buf

  (
    g178_p_spl_,
    g178_p
  );


  buf

  (
    g178_n_spl_,
    g178_n
  );


  buf

  (
    g178_n_spl_0,
    g178_n_spl_
  );


  buf

  (
    g206_p_spl_,
    g206_p
  );


  buf

  (
    g81_n_spl_,
    g81_n
  );


  buf

  (
    g206_n_spl_,
    g206_n
  );


  buf

  (
    g81_p_spl_,
    g81_p
  );


  buf

  (
    g207_p_spl_,
    g207_p
  );


  buf

  (
    g40_n_spl_,
    g40_n
  );


  buf

  (
    g207_n_spl_,
    g207_n
  );


  buf

  (
    g40_p_spl_,
    g40_p
  );


  buf

  (
    g208_n_spl_,
    g208_n
  );


  buf

  (
    g208_n_spl_0,
    g208_n_spl_
  );


  buf

  (
    g208_n_spl_00,
    g208_n_spl_0
  );


  buf

  (
    g208_n_spl_01,
    g208_n_spl_0
  );


  buf

  (
    g208_n_spl_1,
    g208_n_spl_
  );


  buf

  (
    g208_n_spl_10,
    g208_n_spl_1
  );


  buf

  (
    g208_p_spl_,
    g208_p
  );


  buf

  (
    g208_p_spl_0,
    g208_p_spl_
  );


  buf

  (
    g208_p_spl_00,
    g208_p_spl_0
  );


  buf

  (
    g208_p_spl_01,
    g208_p_spl_0
  );


  buf

  (
    g208_p_spl_1,
    g208_p_spl_
  );


  buf

  (
    g208_p_spl_10,
    g208_p_spl_1
  );


  buf

  (
    G30_n_spl_,
    G30_n
  );


  buf

  (
    G30_p_spl_,
    G30_p
  );


  buf

  (
    g221_p_spl_,
    g221_p
  );


  buf

  (
    g221_n_spl_,
    g221_n
  );


  buf

  (
    g223_n_spl_,
    g223_n
  );


  buf

  (
    g223_n_spl_0,
    g223_n_spl_
  );


  buf

  (
    g223_p_spl_,
    g223_p
  );


  buf

  (
    g223_p_spl_0,
    g223_p_spl_
  );


  buf

  (
    g224_n_spl_,
    g224_n
  );


  buf

  (
    g224_n_spl_0,
    g224_n_spl_
  );


  buf

  (
    g224_n_spl_00,
    g224_n_spl_0
  );


  buf

  (
    g224_n_spl_01,
    g224_n_spl_0
  );


  buf

  (
    g224_n_spl_1,
    g224_n_spl_
  );


  buf

  (
    g224_p_spl_,
    g224_p
  );


  buf

  (
    g224_p_spl_0,
    g224_p_spl_
  );


  buf

  (
    g224_p_spl_00,
    g224_p_spl_0
  );


  buf

  (
    g224_p_spl_01,
    g224_p_spl_0
  );


  buf

  (
    g224_p_spl_1,
    g224_p_spl_
  );


  buf

  (
    g235_p_spl_,
    g235_p
  );


  buf

  (
    g235_n_spl_,
    g235_n
  );


  buf

  (
    g236_n_spl_,
    g236_n
  );


  buf

  (
    g236_n_spl_0,
    g236_n_spl_
  );


  buf

  (
    g236_n_spl_1,
    g236_n_spl_
  );


  buf

  (
    g236_p_spl_,
    g236_p
  );


  buf

  (
    g236_p_spl_0,
    g236_p_spl_
  );


  buf

  (
    g236_p_spl_1,
    g236_p_spl_
  );


  buf

  (
    g256_n_spl_,
    g256_n
  );


  buf

  (
    g256_n_spl_0,
    g256_n_spl_
  );


  buf

  (
    g256_n_spl_1,
    g256_n_spl_
  );


  buf

  (
    g256_p_spl_,
    g256_p
  );


  buf

  (
    g256_p_spl_0,
    g256_p_spl_
  );


  buf

  (
    g256_p_spl_1,
    g256_p_spl_
  );


  buf

  (
    g269_p_spl_,
    g269_p
  );


  buf

  (
    g269_p_spl_0,
    g269_p_spl_
  );


  buf

  (
    g269_p_spl_00,
    g269_p_spl_0
  );


  buf

  (
    g269_p_spl_01,
    g269_p_spl_0
  );


  buf

  (
    g269_p_spl_1,
    g269_p_spl_
  );


  buf

  (
    g269_p_spl_10,
    g269_p_spl_1
  );


  buf

  (
    g269_n_spl_,
    g269_n
  );


  buf

  (
    g269_n_spl_0,
    g269_n_spl_
  );


  buf

  (
    g303_n_spl_,
    g303_n
  );


  buf

  (
    g303_p_spl_,
    g303_p
  );


  buf

  (
    g315_n_spl_,
    g315_n
  );


  buf

  (
    g315_p_spl_,
    g315_p
  );


endmodule
