// Benchmark "mymod" written by ABC on Sun Oct 29 19:31:56 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50,
    G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528,
    G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538,
    G3539, G3540  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50;
  output G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528,
    G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538,
    G3539, G3540;
  reg n1836_lo, n1872_lo, n1884_lo, n1911_lo, n1914_lo, n1917_lo, n1923_lo,
    n1926_lo, n1929_lo, n1935_lo, n1938_lo, n1947_lo, n1950_lo, n1959_lo,
    n1962_lo, n1971_lo, n1974_lo, n1983_lo, n1995_lo, n2007_lo, n2019_lo,
    n2031_lo, n2043_lo, n2055_lo, n2064_lo, n2067_lo, n2100_lo, n2112_lo,
    n2124_lo, n2136_lo, n2148_lo, n2160_lo, n2163_lo, n2172_lo, n2175_lo,
    n2184_lo, n2223_lo, n2235_lo, n2238_lo, n2247_lo, n2250_lo, n2259_lo,
    n2262_lo, n2271_lo, n2274_lo, n2283_lo, n2286_lo, n2295_lo, n2298_lo,
    n2304_lo, n2307_lo, n2331_lo, n2334_lo, n2337_lo, n2340_lo, n3241_o2,
    n3242_o2, n3610_o2, n3980_o2, n3968_o2, n4298_o2, n4371_o2, n4413_o2,
    n4418_o2, n4628_o2, n4629_o2, n4633_o2, n4634_o2, n4732_o2, n4733_o2,
    n4884_o2, n4886_o2, n4890_o2, n5011_o2, n5012_o2, n5013_o2, n5014_o2,
    n5015_o2, n5021_o2, n5016_o2, n5026_o2, n4377_o2, n4378_o2, n4389_o2,
    n327_inv, n330_inv, n4398_o2, n4401_o2, n5117_o2, n5115_o2, n5122_o2,
    n5121_o2, n5119_o2, n5116_o2, n5123_o2, n5156_o2, n5167_o2, n4454_o2,
    n4455_o2, n4456_o2, n4505_o2, G742_o2, G727_o2, n4567_o2, n4568_o2,
    n4569_o2, n4571_o2, n4572_o2, n399_inv, n4539_o2, n4651_o2, n4652_o2,
    n4653_o2, G1514_o2, G1823_o2, n4783_o2, n4787_o2, n426_inv, n429_inv,
    n4816_o2, n435_inv, G572_o2, n4919_o2, n4920_o2, n4921_o2, G1048_o2,
    n5041_o2, n5094_o2, n5278_o2, n5301_o2, G2610_o2, G3174_o2, G3146_o2,
    G3217_o2, G3220_o2, G2839_o2, G3251_o2, G3042_o2, G3045_o2, G3262_o2,
    G2845_o2, G2929_o2, G2848_o2, G2851_o2, G3291_o2, G3254_o2, G2666_o2,
    n5099_o2, n5100_o2, n5101_o2, G2558_o2, n5266_o2, n5267_o2, G2759_o2,
    n537_inv, n540_inv, n543_inv, n5292_o2, n5293_o2, n5294_o2, n5295_o2,
    G618_o2, G621_o2, G384_o2, G377_o2, n570_inv, G3171_o2, G2552_o2,
    G3272_o2, G2015_o2, G3294_o2, G3281_o2, G3320_o2, G3275_o2, G3140_o2,
    G2836_o2, G2926_o2, G2842_o2, G3302_o2, G3288_o2, G3143_o2, G3100_o2,
    G2512_o2, n5325_o2, n5326_o2, n5327_o2, n1857_lo_buf_o2,
    n2097_lo_buf_o2, G2669_o2, n642_inv, G568_o2, n648_inv, G565_o2,
    G559_o2, n1821_lo_buf_o2, n1905_lo_buf_o2, n2133_lo_buf_o2,
    n2145_lo_buf_o2, n2157_lo_buf_o2, n2205_lo_buf_o2, n2217_lo_buf_o2,
    G447_o2, G434_o2, G422_o2, G461_o2, G3312_o2, G3332_o2, G3195_o2,
    G2607_o2, n702_inv, G1005_o2, G1008_o2, n2001_lo_buf_o2,
    n2169_lo_buf_o2, n2229_lo_buf_o2, n2301_lo_buf_o2, n723_inv, G2947_o2,
    n2013_lo_buf_o2, n2025_lo_buf_o2, n2037_lo_buf_o2, n2049_lo_buf_o2,
    n2181_lo_buf_o2, n744_inv, n747_inv, n750_inv, n753_inv, G3350_o2,
    G3360_o2, G3373_o2, G3237_o2, G2773_o2, G1733_o2, G1738_o2, G1751_o2,
    G2216_o2, G2219_o2, n786_inv, n789_inv, G787_o2, G2823_o2, G2796_o2,
    G875_o2, G2208_o2, G2211_o2, n1989_lo_buf_o2, n2061_lo_buf_o2,
    n2313_lo_buf_o2, G2232_o2, G1725_o2, G1764_o2, G2356_o2, G2359_o2,
    G1180_o2, G1756_o2, G2441_o2, G2887_o2, G2991_o2, n849_inv, n852_inv,
    n855_inv, n858_inv, n861_inv, G2805_o2, G2906_o2, G2833_o2, n873_inv,
    G3353_o2, G3367_o2, G3346_o2, G3340_o2, G3376_o2, G3359_o2, G3240_o2,
    G3344_o2, G2880_o2, G2939_o2, G2248_o2, G2251_o2, G2021_o2, G3383_o2,
    G3399_o2, G3404_o2, G3265_o2, G2866_o2, G2999_o2, G736_o2, G739_o2,
    G1200_o2, G1203_o2, G3027_o2, G1463_o2, G1460_o2, G3012_o2, G1574_o2,
    G1646_o2, G1592_o2, G1664_o2, G1547_o2, G1619_o2, G1556_o2, G1628_o2,
    G1583_o2, G1655_o2, G1529_o2, G1601_o2, G1538_o2, G1610_o2, G1565_o2,
    G1637_o2, G2437_o2, n1008_inv, n1785_lo_buf_o2, n1845_lo_buf_o2,
    n1893_lo_buf_o2, n1941_lo_buf_o2, n1953_lo_buf_o2, n1965_lo_buf_o2,
    n1977_lo_buf_o2, n2241_lo_buf_o2, n2253_lo_buf_o2, n2265_lo_buf_o2,
    n2277_lo_buf_o2, n2289_lo_buf_o2, G519_o2, n1050_inv, n1053_inv,
    n1056_inv, G1318_o2, n1062_inv, G593_o2, n1068_inv, n1071_inv,
    n1074_inv, G2284_o2, G2580_o2, G2302_o2, G2598_o2, G2497_o2, G2651_o2,
    G2296_o2, G2308_o2, G2592_o2, G2604_o2, G2902_o2, G2975_o2, G2962_o2,
    G3069_o2, G2018_o2, G1176_o2, G1189_o2, G3066_o2, G3137_o2, G3038_o2,
    G3117_o2, G2384_o2, G2472_o2, G772_o2, G935_o2, G2923_o2, G2971_o2,
    G2980_o2, G3039_o2, G2388_o2, G2287_o2, G3024_o2, G2916_o2, n1176_inv,
    G3035_o2, G3107_o2, G1023_o2, G1024_o2, G1311_o2, G1312_o2, G3063_o2,
    G1520_o2, G1519_o2, G3078_o2, G2038_o2, G1848_o2, G1864_o2, G1872_o2,
    G1880_o2, G1888_o2, G1912_o2, G1928_o2, G1936_o2, G1944_o2, G1952_o2,
    G1850_o2, G1866_o2, G1874_o2, G1882_o2, G1890_o2, G1914_o2, G1930_o2,
    G1938_o2, G1946_o2, G1954_o2, G1845_o2, G1861_o2, G1869_o2, G1877_o2,
    G1885_o2, G1909_o2, G1925_o2, G1933_o2, G1941_o2, G1949_o2, G1846_o2,
    G1862_o2, G1870_o2, G1878_o2, G1886_o2, G1910_o2, G1926_o2, G1934_o2,
    G1942_o2, G1950_o2, G1849_o2, G1865_o2, G1873_o2, G1881_o2, G1889_o2,
    G1913_o2, G1929_o2, G1937_o2, G1945_o2, G1953_o2, G1843_o2, G1859_o2,
    G1867_o2, G1875_o2, G1883_o2, G1907_o2, G1923_o2, G1931_o2, G1939_o2,
    G1947_o2, G1844_o2, G1860_o2, G1868_o2, G1876_o2, G1884_o2, G1908_o2,
    G1924_o2, G1932_o2, G1940_o2, G1948_o2, G1847_o2, G1863_o2, G1871_o2,
    G1879_o2, G1887_o2, G1911_o2, G1927_o2, G1935_o2, G1943_o2, G1951_o2,
    G2444_o2, G2451_o2, G2502_o2, G2507_o2, n1464_inv, G2583_o2,
    n1797_lo_buf_o2, n1833_lo_buf_o2, n1881_lo_buf_o2, n1479_inv,
    n1482_inv, n1485_inv, G615_o2, G2254_o2, G2255_o2, G2027_o2, G2393_o2,
    G527_o2, G594_o2, G1689_o2, G1693_o2, G2281_o2, G2014_o2, G2459_o2,
    G2561_o2, G2533_o2, n1749_lo_buf_o2, n1761_lo_buf_o2, n1773_lo_buf_o2,
    n1809_lo_buf_o2, G1955_o2, G1958_o2, G2562_o2, G2398_o2, n1554_inv,
    n1557_inv, G2577_o2, G2627_o2, G654_o2, G660_o2, G831_o2, G919_o2,
    G925_o2, n1815_lo_buf_o2, n1899_lo_buf_o2, n2079_lo_buf_o2,
    n2127_lo_buf_o2, n2139_lo_buf_o2, n2151_lo_buf_o2, n2187_lo_buf_o2,
    n2199_lo_buf_o2, n2211_lo_buf_o2, G533_o2, n1854_lo_buf_o2,
    n2094_lo_buf_o2, G667_o2, G874_o2, G851_o2, G1127_o2, n1869_lo_buf_o2,
    n2109_lo_buf_o2, n2121_lo_buf_o2, G477_o2, G491_o2, G501_o2, G786_o2,
    G791_o2, G1126_o2, G1052_o2, G1054_o2;
  wire new_new_n1131__, new_new_n1133__, new_new_n1135__, new_new_n1136__,
    new_new_n1137__, new_new_n1139__, new_new_n1141__, new_new_n1143__,
    new_new_n1145__, new_new_n1147__, new_new_n1149__, new_new_n1151__,
    new_new_n1153__, new_new_n1155__, new_new_n1157__, new_new_n1159__,
    new_new_n1161__, new_new_n1163__, new_new_n1165__, new_new_n1167__,
    new_new_n1169__, new_new_n1171__, new_new_n1173__, new_new_n1175__,
    new_new_n1177__, new_new_n1179__, new_new_n1181__, new_new_n1183__,
    new_new_n1185__, new_new_n1187__, new_new_n1189__, new_new_n1191__,
    new_new_n1193__, new_new_n1195__, new_new_n1197__, new_new_n1199__,
    new_new_n1201__, new_new_n1203__, new_new_n1205__, new_new_n1207__,
    new_new_n1209__, new_new_n1211__, new_new_n1213__, new_new_n1215__,
    new_new_n1217__, new_new_n1219__, new_new_n1221__, new_new_n1223__,
    new_new_n1225__, new_new_n1227__, new_new_n1229__, new_new_n1231__,
    new_new_n1232__, new_new_n1234__, new_new_n1235__, new_new_n1236__,
    new_new_n1237__, new_new_n1239__, new_new_n1242__, new_new_n1243__,
    new_new_n1245__, new_new_n1248__, new_new_n1249__, new_new_n1251__,
    new_new_n1253__, new_new_n1255__, new_new_n1257__, new_new_n1259__,
    new_new_n1261__, new_new_n1263__, new_new_n1265__, new_new_n1267__,
    new_new_n1268__, new_new_n1269__, new_new_n1270__, new_new_n1271__,
    new_new_n1272__, new_new_n1273__, new_new_n1274__, new_new_n1275__,
    new_new_n1276__, new_new_n1277__, new_new_n1278__, new_new_n1279__,
    new_new_n1281__, new_new_n1284__, new_new_n1286__, new_new_n1288__,
    new_new_n1290__, new_new_n1292__, new_new_n1294__, new_new_n1295__,
    new_new_n1296__, new_new_n1298__, new_new_n1299__, new_new_n1302__,
    new_new_n1303__, new_new_n1305__, new_new_n1307__, new_new_n1309__,
    new_new_n1311__, new_new_n1313__, new_new_n1315__, new_new_n1317__,
    new_new_n1319__, new_new_n1321__, new_new_n1323__, new_new_n1325__,
    new_new_n1327__, new_new_n1328__, new_new_n1329__, new_new_n1330__,
    new_new_n1331__, new_new_n1332__, new_new_n1333__, new_new_n1335__,
    new_new_n1337__, new_new_n1339__, new_new_n1340__, new_new_n1341__,
    new_new_n1342__, new_new_n1343__, new_new_n1344__, new_new_n1346__,
    new_new_n1348__, new_new_n1350__, new_new_n1351__, new_new_n1353__,
    new_new_n1356__, new_new_n1357__, new_new_n1359__, new_new_n1362__,
    new_new_n1363__, new_new_n1364__, new_new_n1365__, new_new_n1366__,
    new_new_n1367__, new_new_n1368__, new_new_n1369__, new_new_n1370__,
    new_new_n1372__, new_new_n1374__, new_new_n1375__, new_new_n1377__,
    new_new_n1378__, new_new_n1379__, new_new_n1380__, new_new_n1381__,
    new_new_n1382__, new_new_n1383__, new_new_n1385__, new_new_n1386__,
    new_new_n1387__, new_new_n1389__, new_new_n1392__, new_new_n1393__,
    new_new_n1395__, new_new_n1397__, new_new_n1398__, new_new_n1399__,
    new_new_n1401__, new_new_n1403__, new_new_n1404__, new_new_n1405__,
    new_new_n1406__, new_new_n1407__, new_new_n1409__, new_new_n1411__,
    new_new_n1413__, new_new_n1415__, new_new_n1417__, new_new_n1419__,
    new_new_n1420__, new_new_n1421__, new_new_n1422__, new_new_n1423__,
    new_new_n1424__, new_new_n1425__, new_new_n1427__, new_new_n1429__,
    new_new_n1431__, new_new_n1433__, new_new_n1434__, new_new_n1436__,
    new_new_n1437__, new_new_n1439__, new_new_n1441__, new_new_n1443__,
    new_new_n1444__, new_new_n1445__, new_new_n1446__, new_new_n1447__,
    new_new_n1449__, new_new_n1450__, new_new_n1451__, new_new_n1452__,
    new_new_n1453__, new_new_n1455__, new_new_n1456__, new_new_n1457__,
    new_new_n1458__, new_new_n1459__, new_new_n1460__, new_new_n1461__,
    new_new_n1462__, new_new_n1463__, new_new_n1465__, new_new_n1467__,
    new_new_n1468__, new_new_n1469__, new_new_n1470__, new_new_n1471__,
    new_new_n1473__, new_new_n1474__, new_new_n1475__, new_new_n1476__,
    new_new_n1477__, new_new_n1479__, new_new_n1481__, new_new_n1482__,
    new_new_n1483__, new_new_n1484__, new_new_n1485__, new_new_n1486__,
    new_new_n1487__, new_new_n1488__, new_new_n1489__, new_new_n1490__,
    new_new_n1491__, new_new_n1493__, new_new_n1495__, new_new_n1497__,
    new_new_n1499__, new_new_n1501__, new_new_n1503__, new_new_n1505__,
    new_new_n1508__, new_new_n1509__, new_new_n1511__, new_new_n1513__,
    new_new_n1515__, new_new_n1517__, new_new_n1519__, new_new_n1521__,
    new_new_n1523__, new_new_n1524__, new_new_n1525__, new_new_n1527__,
    new_new_n1528__, new_new_n1529__, new_new_n1530__, new_new_n1531__,
    new_new_n1533__, new_new_n1534__, new_new_n1535__, new_new_n1536__,
    new_new_n1537__, new_new_n1538__, new_new_n1539__, new_new_n1541__,
    new_new_n1543__, new_new_n1545__, new_new_n1547__, new_new_n1549__,
    new_new_n1550__, new_new_n1551__, new_new_n1553__, new_new_n1554__,
    new_new_n1555__, new_new_n1556__, new_new_n1558__, new_new_n1560__,
    new_new_n1561__, new_new_n1562__, new_new_n1563__, new_new_n1565__,
    new_new_n1567__, new_new_n1569__, new_new_n1570__, new_new_n1571__,
    new_new_n1573__, new_new_n1575__, new_new_n1577__, new_new_n1579__,
    new_new_n1581__, new_new_n1583__, new_new_n1585__, new_new_n1587__,
    new_new_n1589__, new_new_n1591__, new_new_n1594__, new_new_n1595__,
    new_new_n1596__, new_new_n1597__, new_new_n1598__, new_new_n1599__,
    new_new_n1600__, new_new_n1601__, new_new_n1602__, new_new_n1603__,
    new_new_n1604__, new_new_n1605__, new_new_n1606__, new_new_n1607__,
    new_new_n1608__, new_new_n1609__, new_new_n1611__, new_new_n1613__,
    new_new_n1615__, new_new_n1617__, new_new_n1619__, new_new_n1620__,
    new_new_n1621__, new_new_n1622__, new_new_n1623__, new_new_n1624__,
    new_new_n1625__, new_new_n1626__, new_new_n1627__, new_new_n1628__,
    new_new_n1629__, new_new_n1631__, new_new_n1633__, new_new_n1634__,
    new_new_n1635__, new_new_n1638__, new_new_n1639__, new_new_n1641__,
    new_new_n1643__, new_new_n1645__, new_new_n1647__, new_new_n1649__,
    new_new_n1651__, new_new_n1653__, new_new_n1655__, new_new_n1657__,
    new_new_n1658__, new_new_n1659__, new_new_n1661__, new_new_n1662__,
    new_new_n1663__, new_new_n1665__, new_new_n1667__, new_new_n1668__,
    new_new_n1669__, new_new_n1670__, new_new_n1671__, new_new_n1672__,
    new_new_n1673__, new_new_n1674__, new_new_n1675__, new_new_n1676__,
    new_new_n1677__, new_new_n1679__, new_new_n1681__, new_new_n1683__,
    new_new_n1685__, new_new_n1686__, new_new_n1687__, new_new_n1688__,
    new_new_n1689__, new_new_n1690__, new_new_n1691__, new_new_n1692__,
    new_new_n1693__, new_new_n1694__, new_new_n1695__, new_new_n1696__,
    new_new_n1697__, new_new_n1698__, new_new_n1699__, new_new_n1700__,
    new_new_n1701__, new_new_n1702__, new_new_n1703__, new_new_n1704__,
    new_new_n1705__, new_new_n1707__, new_new_n1709__, new_new_n1711__,
    new_new_n1713__, new_new_n1715__, new_new_n1716__, new_new_n1717__,
    new_new_n1718__, new_new_n1719__, new_new_n1720__, new_new_n1721__,
    new_new_n1723__, new_new_n1724__, new_new_n1725__, new_new_n1726__,
    new_new_n1727__, new_new_n1728__, new_new_n1729__, new_new_n1730__,
    new_new_n1731__, new_new_n1732__, new_new_n1733__, new_new_n1734__,
    new_new_n1735__, new_new_n1736__, new_new_n1737__, new_new_n1738__,
    new_new_n1739__, new_new_n1740__, new_new_n1742__, new_new_n1743__,
    new_new_n1744__, new_new_n1745__, new_new_n1746__, new_new_n1747__,
    new_new_n1748__, new_new_n1749__, new_new_n1750__, new_new_n1751__,
    new_new_n1752__, new_new_n1753__, new_new_n1754__, new_new_n1755__,
    new_new_n1756__, new_new_n1757__, new_new_n1759__, new_new_n1761__,
    new_new_n1763__, new_new_n1765__, new_new_n1766__, new_new_n1767__,
    new_new_n1768__, new_new_n1769__, new_new_n1770__, new_new_n1771__,
    new_new_n1772__, new_new_n1773__, new_new_n1774__, new_new_n1775__,
    new_new_n1776__, new_new_n1777__, new_new_n1778__, new_new_n1779__,
    new_new_n1780__, new_new_n1781__, new_new_n1782__, new_new_n1783__,
    new_new_n1784__, new_new_n1785__, new_new_n1786__, new_new_n1787__,
    new_new_n1788__, new_new_n1789__, new_new_n1791__, new_new_n1792__,
    new_new_n1793__, new_new_n1794__, new_new_n1795__, new_new_n1796__,
    new_new_n1797__, new_new_n1798__, new_new_n1799__, new_new_n1800__,
    new_new_n1801__, new_new_n1802__, new_new_n1804__, new_new_n1805__,
    new_new_n1807__, new_new_n1809__, new_new_n1811__, new_new_n1812__,
    new_new_n1814__, new_new_n1816__, new_new_n1817__, new_new_n1818__,
    new_new_n1819__, new_new_n1821__, new_new_n1823__, new_new_n1825__,
    new_new_n1828__, new_new_n1830__, new_new_n1831__, new_new_n1833__,
    new_new_n1836__, new_new_n1838__, new_new_n1839__, new_new_n1841__,
    new_new_n1843__, new_new_n1845__, new_new_n1847__, new_new_n1849__,
    new_new_n1851__, new_new_n1852__, new_new_n1853__, new_new_n1855__,
    new_new_n1856__, new_new_n1857__, new_new_n1858__, new_new_n1859__,
    new_new_n1860__, new_new_n1862__, new_new_n1864__, new_new_n1866__,
    new_new_n1867__, new_new_n1868__, new_new_n1869__, new_new_n1870__,
    new_new_n1871__, new_new_n1872__, new_new_n1873__, new_new_n1874__,
    new_new_n1875__, new_new_n1876__, new_new_n1877__, new_new_n1879__,
    new_new_n1880__, new_new_n1881__, new_new_n1882__, new_new_n1883__,
    new_new_n1884__, new_new_n1885__, new_new_n1886__, new_new_n1888__,
    new_new_n1889__, new_new_n1890__, new_new_n1891__, new_new_n1892__,
    new_new_n1893__, new_new_n1894__, new_new_n1895__, new_new_n1896__,
    new_new_n1897__, new_new_n1898__, new_new_n1899__, new_new_n1900__,
    new_new_n1901__, new_new_n1902__, new_new_n1903__, new_new_n1904__,
    new_new_n1905__, new_new_n1906__, new_new_n1907__, new_new_n1908__,
    new_new_n1909__, new_new_n1910__, new_new_n1911__, new_new_n1912__,
    new_new_n1913__, new_new_n1914__, new_new_n1915__, new_new_n1916__,
    new_new_n1917__, new_new_n1918__, new_new_n1919__, new_new_n1920__,
    new_new_n1921__, new_new_n1922__, new_new_n1923__, new_new_n1924__,
    new_new_n1925__, new_new_n1926__, new_new_n1927__, new_new_n1929__,
    new_new_n1930__, new_new_n1931__, new_new_n1932__, new_new_n1933__,
    new_new_n1934__, new_new_n1935__, new_new_n1936__, new_new_n1937__,
    new_new_n1938__, new_new_n1939__, new_new_n1940__, new_new_n1941__,
    new_new_n1942__, new_new_n1943__, new_new_n1944__, new_new_n1945__,
    new_new_n1946__, new_new_n1947__, new_new_n1949__, new_new_n1950__,
    new_new_n1951__, new_new_n1952__, new_new_n1953__, new_new_n1954__,
    new_new_n1955__, new_new_n1956__, new_new_n1957__, new_new_n1958__,
    new_new_n1959__, new_new_n1960__, new_new_n1961__, new_new_n1962__,
    new_new_n1963__, new_new_n1964__, new_new_n1965__, new_new_n1966__,
    new_new_n1967__, new_new_n1968__, new_new_n1969__, new_new_n1970__,
    new_new_n1971__, new_new_n1974__, new_new_n1976__, new_new_n1978__,
    new_new_n1979__, new_new_n1980__, new_new_n1981__, new_new_n1983__,
    new_new_n1985__, new_new_n1986__, new_new_n1987__, new_new_n1989__,
    new_new_n1991__, new_new_n1994__, new_new_n1995__, new_new_n1998__,
    new_new_n1999__, new_new_n2001__, new_new_n2004__, new_new_n2005__,
    new_new_n2008__, new_new_n2009__, new_new_n2011__, new_new_n2014__,
    new_new_n2015__, new_new_n2018__, new_new_n2019__, new_new_n2021__,
    new_new_n2024__, new_new_n2025__, new_new_n2028__, new_new_n2030__,
    new_new_n2032__, new_new_n2033__, new_new_n2036__, new_new_n2037__,
    new_new_n2040__, new_new_n2042__, new_new_n2043__, new_new_n2046__,
    new_new_n2047__, new_new_n2049__, new_new_n2051__, new_new_n2054__,
    new_new_n2055__, new_new_n2058__, new_new_n2059__, new_new_n2061__,
    new_new_n2064__, new_new_n2065__, new_new_n2068__, new_new_n2070__,
    new_new_n2072__, new_new_n2073__, new_new_n2076__, new_new_n2077__,
    new_new_n2080__, new_new_n2082__, new_new_n2083__, new_new_n2086__,
    new_new_n2087__, new_new_n2089__, new_new_n2091__, new_new_n2094__,
    new_new_n2095__, new_new_n2098__, new_new_n2099__, new_new_n2101__,
    new_new_n2104__, new_new_n2105__, new_new_n2108__, new_new_n2109__,
    new_new_n2111__, new_new_n2114__, new_new_n2115__, new_new_n2118__,
    new_new_n2119__, new_new_n2121__, new_new_n2124__, new_new_n2125__,
    new_new_n2128__, new_new_n2129__, new_new_n2131__, new_new_n2134__,
    new_new_n2135__, new_new_n2138__, new_new_n2139__, new_new_n2141__,
    new_new_n2144__, new_new_n2145__, new_new_n2148__, new_new_n2149__,
    new_new_n2150__, new_new_n2151__, new_new_n2152__, new_new_n2153__,
    new_new_n2154__, new_new_n2155__, new_new_n2156__, new_new_n2157__,
    new_new_n2159__, new_new_n2160__, new_new_n2161__, new_new_n2162__,
    new_new_n2163__, new_new_n2164__, new_new_n2165__, new_new_n2166__,
    new_new_n2167__, new_new_n2169__, new_new_n2171__, new_new_n2173__,
    new_new_n2174__, new_new_n2175__, new_new_n2176__, new_new_n2177__,
    new_new_n2178__, new_new_n2179__, new_new_n2180__, new_new_n2181__,
    new_new_n2182__, new_new_n2183__, new_new_n2184__, new_new_n2185__,
    new_new_n2186__, new_new_n2187__, new_new_n2188__, new_new_n2189__,
    new_new_n2190__, new_new_n2191__, new_new_n2192__, new_new_n2193__,
    new_new_n2194__, new_new_n2195__, new_new_n2196__, new_new_n2197__,
    new_new_n2198__, new_new_n2199__, new_new_n2200__, new_new_n2201__,
    new_new_n2202__, new_new_n2203__, new_new_n2204__, new_new_n2205__,
    new_new_n2206__, new_new_n2207__, new_new_n2208__, new_new_n2209__,
    new_new_n2210__, new_new_n2211__, new_new_n2212__, new_new_n2213__,
    new_new_n2214__, new_new_n2215__, new_new_n2216__, new_new_n2217__,
    new_new_n2218__, new_new_n2219__, new_new_n2220__, new_new_n2221__,
    new_new_n2222__, new_new_n2223__, new_new_n2224__, new_new_n2225__,
    new_new_n2226__, new_new_n2227__, new_new_n2228__, new_new_n2229__,
    new_new_n2230__, new_new_n2231__, new_new_n2232__, new_new_n2233__,
    new_new_n2234__, new_new_n2235__, new_new_n2236__, new_new_n2237__,
    new_new_n2238__, new_new_n2239__, new_new_n2240__, new_new_n2241__,
    new_new_n2242__, new_new_n2243__, new_new_n2244__, new_new_n2245__,
    new_new_n2246__, new_new_n2247__, new_new_n2248__, new_new_n2249__,
    new_new_n2250__, new_new_n2251__, new_new_n2252__, new_new_n2253__,
    new_new_n2254__, new_new_n2255__, new_new_n2256__, new_new_n2257__,
    new_new_n2258__, new_new_n2259__, new_new_n2260__, new_new_n2261__,
    new_new_n2262__, new_new_n2263__, new_new_n2264__, new_new_n2265__,
    new_new_n2266__, new_new_n2267__, new_new_n2268__, new_new_n2269__,
    new_new_n2270__, new_new_n2271__, new_new_n2272__, new_new_n2273__,
    new_new_n2274__, new_new_n2275__, new_new_n2276__, new_new_n2277__,
    new_new_n2278__, new_new_n2279__, new_new_n2280__, new_new_n2281__,
    new_new_n2282__, new_new_n2283__, new_new_n2284__, new_new_n2285__,
    new_new_n2286__, new_new_n2287__, new_new_n2288__, new_new_n2289__,
    new_new_n2290__, new_new_n2291__, new_new_n2292__, new_new_n2293__,
    new_new_n2294__, new_new_n2295__, new_new_n2296__, new_new_n2297__,
    new_new_n2298__, new_new_n2299__, new_new_n2300__, new_new_n2301__,
    new_new_n2302__, new_new_n2303__, new_new_n2304__, new_new_n2305__,
    new_new_n2306__, new_new_n2307__, new_new_n2308__, new_new_n2309__,
    new_new_n2310__, new_new_n2311__, new_new_n2312__, new_new_n2313__,
    new_new_n2314__, new_new_n2315__, new_new_n2316__, new_new_n2317__,
    new_new_n2318__, new_new_n2319__, new_new_n2320__, new_new_n2321__,
    new_new_n2322__, new_new_n2323__, new_new_n2324__, new_new_n2325__,
    new_new_n2326__, new_new_n2327__, new_new_n2328__, new_new_n2329__,
    new_new_n2330__, new_new_n2331__, new_new_n2332__, new_new_n2333__,
    new_new_n2334__, new_new_n2335__, new_new_n2336__, new_new_n2337__,
    new_new_n2338__, new_new_n2339__, new_new_n2340__, new_new_n2341__,
    new_new_n2342__, new_new_n2343__, new_new_n2344__, new_new_n2345__,
    new_new_n2346__, new_new_n2347__, new_new_n2348__, new_new_n2349__,
    new_new_n2350__, new_new_n2351__, new_new_n2352__, new_new_n2353__,
    new_new_n2354__, new_new_n2355__, new_new_n2356__, new_new_n2357__,
    new_new_n2358__, new_new_n2359__, new_new_n2360__, new_new_n2361__,
    new_new_n2362__, new_new_n2363__, new_new_n2364__, new_new_n2365__,
    new_new_n2366__, new_new_n2367__, new_new_n2368__, new_new_n2369__,
    new_new_n2370__, new_new_n2371__, new_new_n2372__, new_new_n2373__,
    new_new_n2374__, new_new_n2375__, new_new_n2376__, new_new_n2377__,
    new_new_n2378__, new_new_n2379__, new_new_n2380__, new_new_n2381__,
    new_new_n2382__, new_new_n2383__, new_new_n2384__, new_new_n2385__,
    new_new_n2386__, new_new_n2387__, new_new_n2388__, new_new_n2389__,
    new_new_n2390__, new_new_n2391__, new_new_n2392__, new_new_n2393__,
    new_new_n2394__, new_new_n2395__, new_new_n2396__, new_new_n2397__,
    new_new_n2398__, new_new_n2399__, new_new_n2400__, new_new_n2401__,
    new_new_n2402__, new_new_n2403__, new_new_n2404__, new_new_n2405__,
    new_new_n2406__, new_new_n2407__, new_new_n2408__, new_new_n2409__,
    new_new_n2410__, new_new_n2411__, new_new_n2412__, new_new_n2413__,
    new_new_n2414__, new_new_n2415__, new_new_n2416__, new_new_n2417__,
    new_new_n2418__, new_new_n2419__, new_new_n2420__, new_new_n2421__,
    new_new_n2422__, new_new_n2423__, new_new_n2424__, new_new_n2425__,
    new_new_n2426__, new_new_n2427__, new_new_n2428__, new_new_n2429__,
    new_new_n2430__, new_new_n2431__, new_new_n2432__, new_new_n2433__,
    new_new_n2434__, new_new_n2435__, new_new_n2436__, new_new_n2437__,
    new_new_n2438__, new_new_n2439__, new_new_n2440__, new_new_n2441__,
    new_new_n2442__, new_new_n2443__, new_new_n2444__, new_new_n2445__,
    new_new_n2446__, new_new_n2447__, new_new_n2448__, new_new_n2449__,
    new_new_n2450__, new_new_n2451__, new_new_n2452__, new_new_n2453__,
    new_new_n2454__, new_new_n2455__, new_new_n2456__, new_new_n2457__,
    new_new_n2458__, new_new_n2459__, new_new_n2460__, new_new_n2461__,
    new_new_n2462__, new_new_n2463__, new_new_n2464__, new_new_n2465__,
    new_new_n2466__, new_new_n2467__, new_new_n2468__, new_new_n2469__,
    new_new_n2470__, new_new_n2471__, new_new_n2472__, new_new_n2473__,
    new_new_n2474__, new_new_n2475__, new_new_n2476__, new_new_n2477__,
    new_new_n2478__, new_new_n2479__, new_new_n2480__, new_new_n2481__,
    new_new_n2482__, new_new_n2483__, new_new_n2484__, new_new_n2485__,
    new_new_n2486__, new_new_n2487__, new_new_n2488__, new_new_n2489__,
    new_new_n2490__, new_new_n2491__, new_new_n2492__, new_new_n2493__,
    new_new_n2494__, new_new_n2495__, new_new_n2496__, new_new_n2497__,
    new_new_n2498__, new_new_n2499__, new_new_n2500__, new_new_n2501__,
    new_new_n2502__, new_new_n2503__, new_new_n2504__, new_new_n2505__,
    new_new_n2506__, new_new_n2507__, new_new_n2508__, new_new_n2509__,
    new_new_n2510__, new_new_n2511__, new_new_n2512__, new_new_n2513__,
    new_new_n2514__, new_new_n2515__, new_new_n2516__, new_new_n2517__,
    new_new_n2518__, new_new_n2519__, new_new_n2520__, new_new_n2521__,
    new_new_n2522__, new_new_n2523__, new_new_n2524__, new_new_n2525__,
    new_new_n2526__, new_new_n2527__, new_new_n2528__, new_new_n2529__,
    new_new_n2530__, new_new_n2531__, new_new_n2532__, new_new_n2533__,
    new_new_n2534__, new_new_n2535__, new_new_n2536__, new_new_n2537__,
    new_new_n2538__, new_new_n2539__, new_new_n2540__, new_new_n2541__,
    new_new_n2542__, new_new_n2543__, new_new_n2544__, new_new_n2545__,
    new_new_n2546__, new_new_n2547__, new_new_n2548__, new_new_n2549__,
    new_new_n2550__, new_new_n2551__, new_new_n2552__, new_new_n2553__,
    new_new_n2554__, new_new_n2555__, new_new_n2556__, new_new_n2557__,
    new_new_n2558__, new_new_n2559__, new_new_n2560__, new_new_n2561__,
    new_new_n2562__, new_new_n2563__, new_new_n2564__, new_new_n2565__,
    new_new_n2566__, new_new_n2567__, new_new_n2568__, new_new_n2569__,
    new_new_n2570__, new_new_n2571__, new_new_n2572__, new_new_n2573__,
    new_new_n2574__, new_new_n2575__, new_new_n2576__, new_new_n2577__,
    new_new_n2578__, new_new_n2579__, new_new_n2580__, new_new_n2581__,
    new_new_n2582__, new_new_n2583__, new_new_n2584__, new_new_n2585__,
    new_new_n2586__, new_new_n2587__, new_new_n2588__, new_new_n2589__,
    new_new_n2590__, new_new_n2591__, new_new_n2592__, new_new_n2593__,
    new_new_n2594__, new_new_n2595__, new_new_n2596__, new_new_n2597__,
    new_new_n2598__, new_new_n2599__, new_new_n2600__, new_new_n2601__,
    new_new_n2602__, new_new_n2603__, new_new_n2604__, new_new_n2605__,
    new_new_n2606__, new_new_n2607__, new_new_n2608__, new_new_n2609__,
    new_new_n2610__, new_new_n2611__, new_new_n2612__, new_new_n2613__,
    new_new_n2614__, new_new_n2615__, new_new_n2616__, new_new_n2617__,
    new_new_n2618__, new_new_n2619__, new_new_n2620__, new_new_n2621__,
    new_new_n2622__, new_new_n2623__, new_new_n2624__, new_new_n2625__,
    new_new_n2626__, new_new_n2627__, new_new_n2628__, new_new_n2629__,
    new_new_n2630__, new_new_n2631__, new_new_n2632__, new_new_n2633__,
    new_new_n2634__, new_new_n2635__, new_new_n2636__, new_new_n2637__,
    new_new_n2638__, new_new_n2639__, new_new_n2640__, new_new_n2641__,
    new_new_n2642__, new_new_n2643__, new_new_n2644__, new_new_n2645__,
    new_new_n2646__, new_new_n2647__, new_new_n2648__, new_new_n2649__,
    new_new_n2650__, new_new_n2651__, new_new_n2652__, new_new_n2653__,
    new_new_n2654__, new_new_n2655__, new_new_n2656__, new_new_n2657__,
    new_new_n2658__, new_new_n2659__, new_new_n2660__, new_new_n2661__,
    new_new_n2662__, new_new_n2663__, new_new_n2664__, new_new_n2665__,
    new_new_n2666__, new_new_n2667__, new_new_n2668__, new_new_n2669__,
    new_new_n2670__, new_new_n2671__, new_new_n2672__, new_new_n2673__,
    new_new_n2674__, new_new_n2675__, new_new_n2676__, new_new_n2677__,
    new_new_n2678__, new_new_n2679__, new_new_n2680__, new_new_n2681__,
    new_new_n2682__, new_new_n2683__, new_new_n2684__, new_new_n2685__,
    new_new_n2686__, new_new_n2687__, new_new_n2688__, new_new_n2689__,
    new_new_n2690__, new_new_n2691__, new_new_n2692__, new_new_n2693__,
    new_new_n2694__, new_new_n2695__, new_new_n2696__, new_new_n2697__,
    new_new_n2698__, new_new_n2699__, new_new_n2700__, new_new_n2701__,
    new_new_n2702__, new_new_n2703__, new_new_n2704__, new_new_n2705__,
    new_new_n2706__, new_new_n2707__, new_new_n2708__, new_new_n2709__,
    new_new_n2710__, new_new_n2711__, new_new_n2712__, new_new_n2713__,
    new_new_n2714__, new_new_n2715__, new_new_n2716__, new_new_n2717__,
    new_new_n2718__, new_new_n2719__, new_new_n2720__, new_new_n2721__,
    new_new_n2722__, new_new_n2723__, new_new_n2724__, new_new_n2725__,
    new_new_n2726__, new_new_n2727__, new_new_n2728__, new_new_n2729__,
    new_new_n2730__, new_new_n2731__, new_new_n2732__, new_new_n2733__,
    new_new_n2734__, new_new_n2735__, new_new_n2736__, new_new_n2737__,
    new_new_n2738__, new_new_n2739__, new_new_n2740__, new_new_n2741__,
    new_new_n2742__, new_new_n2743__, new_new_n2744__, new_new_n2745__,
    new_new_n2746__, new_new_n2747__, new_new_n2748__, new_new_n2749__,
    new_new_n2750__, new_new_n2751__, new_new_n2752__, new_new_n2753__,
    new_new_n2754__, new_new_n2755__, new_new_n2756__, new_new_n2757__,
    new_new_n2758__, new_new_n2759__, new_new_n2760__, new_new_n2761__,
    new_new_n2762__, new_new_n2763__, new_new_n2764__, new_new_n2765__,
    new_new_n2766__, new_new_n2767__, new_new_n2768__, new_new_n2769__,
    new_new_n2770__, new_new_n2771__, new_new_n2772__, new_new_n2773__,
    new_new_n2774__, new_new_n2775__, new_new_n2776__, new_new_n2777__,
    new_new_n2778__, new_new_n2779__, new_new_n2780__, new_new_n2781__,
    new_new_n2782__, new_new_n2783__, new_new_n2784__, new_new_n2785__,
    new_new_n2786__, new_new_n2787__, new_new_n2788__, new_new_n2789__,
    new_new_n2790__, new_new_n2791__, new_new_n2792__, new_new_n2793__,
    new_new_n2794__, new_new_n2795__, new_new_n2796__, new_new_n2797__,
    new_new_n2798__, new_new_n2799__, new_new_n2800__, new_new_n2801__,
    new_new_n2802__, new_new_n2803__, new_new_n2804__, new_new_n2805__,
    new_new_n2806__, new_new_n2807__, new_new_n2808__, new_new_n2809__,
    new_new_n2810__, new_new_n2811__, new_new_n2812__, new_new_n2813__,
    new_new_n2814__, new_new_n2815__, new_new_n2816__, new_new_n2817__,
    new_new_n2818__, new_new_n2819__, new_new_n2820__, new_new_n2821__,
    new_new_n2822__, new_new_n2823__, new_new_n2824__, new_new_n2825__,
    new_new_n2826__, new_new_n2827__, new_new_n2828__, new_new_n2829__,
    new_new_n2830__, new_new_n2831__, new_new_n2832__, new_new_n2833__,
    new_new_n2834__, new_new_n2835__, new_new_n2836__, new_new_n2837__,
    new_new_n2838__, new_new_n2839__, new_new_n2840__, new_new_n2841__,
    new_new_n2842__, new_new_n2843__, new_new_n2844__, new_new_n2845__,
    new_new_n2846__, new_new_n2847__, new_new_n2848__, new_new_n2849__,
    new_new_n2850__, new_new_n2851__, new_new_n2852__, new_new_n2853__,
    new_new_n2854__, new_new_n2855__, new_new_n2856__, new_new_n2857__,
    new_new_n2858__, new_new_n2859__, new_new_n2860__, new_new_n2861__,
    new_new_n2862__, new_new_n2863__, new_new_n2864__, new_new_n2865__,
    new_new_n2866__, new_new_n2867__, new_new_n2868__, new_new_n2869__,
    new_new_n2870__, new_new_n2871__, new_new_n2872__, new_new_n2873__,
    new_new_n2874__, new_new_n2875__, new_new_n2876__, new_new_n2877__,
    new_new_n2878__, new_new_n2879__, new_new_n2880__, new_new_n2881__,
    new_new_n2882__, new_new_n2883__, new_new_n2884__, new_new_n2885__,
    new_new_n2886__, new_new_n2887__, new_new_n2888__, new_new_n2889__,
    new_new_n2890__, new_new_n2891__, new_new_n2892__, new_new_n2893__,
    new_new_n2894__, new_new_n2895__, new_new_n2896__, new_new_n2897__,
    new_new_n2898__, new_new_n2899__, new_new_n2900__, new_new_n2901__,
    new_new_n2902__, new_new_n2903__, new_new_n2904__, new_new_n2905__,
    new_new_n2906__, new_new_n2907__, new_new_n2908__, new_new_n2909__,
    new_new_n2910__, new_new_n2911__, new_new_n2912__, new_new_n2913__,
    new_new_n2914__, new_new_n2915__, new_new_n2916__, new_new_n2917__,
    new_new_n2918__, new_new_n2919__, new_new_n2920__, new_new_n2921__,
    new_new_n2922__, new_new_n2923__, new_new_n2924__, new_new_n2925__,
    new_new_n2926__, new_new_n2927__, new_new_n2928__, new_new_n2929__,
    new_new_n2930__, new_new_n2931__, new_new_n2932__, new_new_n2933__,
    new_new_n2934__, new_new_n2935__, new_new_n2936__, new_new_n2937__,
    new_new_n2938__, new_new_n2939__, new_new_n2940__, new_new_n2941__,
    new_new_n2942__, new_new_n2943__, new_new_n2944__, new_new_n2945__,
    new_new_n2946__, new_new_n2947__, new_new_n2948__, new_new_n2949__,
    new_new_n2950__, new_new_n2951__, new_new_n2952__, new_new_n2953__,
    new_new_n2954__, new_new_n2955__, new_new_n2956__, new_new_n2957__,
    new_new_n2958__, new_new_n2959__, new_new_n2960__, new_new_n2961__,
    new_new_n2962__, new_new_n2963__, new_new_n2964__, new_new_n2965__,
    new_new_n2966__, new_new_n2967__, new_new_n2968__, new_new_n2969__,
    new_new_n2970__, new_new_n2971__, new_new_n2972__, new_new_n2973__,
    new_new_n2974__, new_new_n2975__, new_new_n2976__, new_new_n2977__,
    new_new_n2978__, new_new_n2979__, new_new_n2980__, new_new_n2981__,
    new_new_n2982__, new_new_n2983__, new_new_n2984__, new_new_n2985__,
    new_new_n2986__, new_new_n2987__, new_new_n2988__, new_new_n2989__,
    new_new_n2990__, new_new_n2991__, new_new_n2992__, new_new_n2993__,
    new_new_n2994__, new_new_n2995__, new_new_n2996__, new_new_n2997__,
    new_new_n2998__, new_new_n2999__, new_new_n3000__, new_new_n3001__,
    new_new_n3002__, new_new_n3003__, new_new_n3004__, new_new_n3005__,
    new_new_n3006__, new_new_n3007__, new_new_n3008__, new_new_n3009__,
    new_new_n3010__, new_new_n3011__, new_new_n3012__, new_new_n3013__,
    new_new_n3014__, new_new_n3015__, new_new_n3016__, new_new_n3017__,
    new_new_n3018__, new_new_n3019__, new_new_n3020__, new_new_n3021__,
    new_new_n3022__, new_new_n3023__, new_new_n3024__, new_new_n3025__,
    new_new_n3026__, new_new_n3027__, new_new_n3028__, new_new_n3029__,
    new_new_n3030__, new_new_n3031__, new_new_n3032__, new_new_n3033__,
    new_new_n3034__, new_new_n3035__, new_new_n3036__, new_new_n3037__,
    new_new_n3038__, new_new_n3039__, new_new_n3040__, new_new_n3041__,
    new_new_n3042__, new_new_n3043__, new_new_n3044__, new_new_n3045__,
    new_new_n3046__, new_new_n3047__, new_new_n3048__, new_new_n3049__,
    new_new_n3050__, new_new_n3051__, new_new_n3052__, new_new_n3053__,
    new_new_n3054__, new_new_n3055__, new_new_n3056__, new_new_n3057__,
    new_new_n3058__, new_new_n3059__, new_new_n3060__, new_new_n3061__,
    new_new_n3062__, new_new_n3063__, new_new_n3064__, new_new_n3065__,
    new_new_n3066__, new_new_n3067__, new_new_n3068__, new_new_n3069__,
    new_new_n3070__, new_new_n3071__, new_new_n3072__, new_new_n3073__,
    new_new_n3074__, new_new_n3075__, new_new_n3076__, new_new_n3077__,
    new_new_n3078__, new_new_n3079__, new_new_n3080__, new_new_n3081__,
    new_new_n3082__, new_new_n3083__, new_new_n3084__, new_new_n3085__,
    new_new_n3086__, new_new_n3087__, new_new_n3088__, new_new_n3089__,
    new_new_n3090__, new_new_n3091__, new_new_n3092__, new_new_n3093__,
    new_new_n3094__, new_new_n3095__, new_new_n3096__, new_new_n3097__,
    new_new_n3098__, new_new_n3099__, new_new_n3100__, new_new_n3101__,
    new_new_n3102__, new_new_n3103__, new_new_n3104__, new_new_n3105__,
    new_new_n3106__, new_new_n3107__, new_new_n3108__, new_new_n3109__,
    new_new_n3110__, new_new_n3111__, new_new_n3112__, new_new_n3113__,
    new_new_n3114__, new_new_n3115__, new_new_n3116__, new_new_n3117__,
    new_new_n3118__, new_new_n3119__, new_new_n3120__, new_new_n3121__,
    new_new_n3122__, new_new_n3123__, new_new_n3124__, new_new_n3125__,
    new_new_n3126__, new_new_n3127__, new_new_n3128__, new_new_n3129__,
    new_new_n3130__, new_new_n3131__, new_new_n3132__, new_new_n3133__,
    new_new_n3134__, new_new_n3135__, new_new_n3136__, new_new_n3137__,
    new_new_n3138__, new_new_n3139__, new_new_n3140__, new_new_n3141__,
    new_new_n3142__, new_new_n3143__, new_new_n3144__, new_new_n3145__,
    new_new_n3146__, new_new_n3147__, new_new_n3148__, new_new_n3149__,
    new_new_n3150__, new_new_n3151__, new_new_n3152__, new_new_n3153__,
    new_new_n3154__, new_new_n3155__, new_new_n3156__, new_new_n3157__,
    new_new_n3158__, new_new_n3159__, new_new_n3160__, new_new_n3161__,
    new_new_n3162__, new_new_n3163__, new_new_n3164__, new_new_n3165__,
    new_new_n3166__, new_new_n3167__, new_new_n3168__, new_new_n3169__,
    new_new_n3170__, new_new_n3171__, new_new_n3172__, new_new_n3173__,
    new_new_n3174__, new_new_n3175__, new_new_n3176__, new_new_n3177__,
    new_new_n3178__, new_new_n3179__, new_new_n3180__, new_new_n3181__,
    new_new_n3182__, new_new_n3183__, new_new_n3184__, new_new_n3185__,
    new_new_n3186__, new_new_n3187__, new_new_n3188__, new_new_n3189__,
    new_new_n3190__, new_new_n3191__, new_new_n3192__, new_new_n3193__,
    new_new_n3194__, new_new_n3195__, new_new_n3196__, new_new_n3197__,
    new_new_n3198__, new_new_n3199__, new_new_n3200__, new_new_n3201__,
    new_new_n3202__, new_new_n3203__, new_new_n3204__, new_new_n3205__,
    new_new_n3206__, new_new_n3207__, new_new_n3208__, new_new_n3209__,
    new_new_n3210__, new_new_n3211__, new_new_n3212__, new_new_n3213__,
    new_new_n3214__, new_new_n3215__, new_new_n3216__, new_new_n3217__,
    new_new_n3218__, new_new_n3219__, new_new_n3220__, new_new_n3221__,
    new_new_n3222__, new_new_n3223__, new_new_n3224__, new_new_n3225__,
    new_new_n3226__, new_new_n3227__, new_new_n3228__, new_new_n3229__,
    new_new_n3230__, new_new_n3231__, new_new_n3232__, new_new_n3233__,
    new_new_n3234__, new_new_n3235__, new_new_n3236__, new_new_n3237__,
    new_new_n3238__, new_new_n3239__, new_new_n3240__, new_new_n3241__,
    new_new_n3242__, new_new_n3243__, new_new_n3244__, new_new_n3245__,
    new_new_n3246__, new_new_n3247__, new_new_n3248__, new_new_n3249__,
    new_new_n3250__, new_new_n3251__, new_new_n3252__, new_new_n3253__,
    new_new_n3254__, new_new_n3255__, new_new_n3256__, new_new_n3257__,
    new_new_n3258__, new_new_n3259__, new_new_n3260__, new_new_n3261__,
    new_new_n3262__, new_new_n3263__, new_new_n3264__, new_new_n3265__,
    new_new_n3266__, new_new_n3267__, new_new_n3268__, new_new_n3269__,
    new_new_n3270__, new_new_n3271__, new_new_n3272__, new_new_n3273__,
    new_new_n3274__, new_new_n3275__, new_new_n3276__, new_new_n3277__,
    new_new_n3278__, new_new_n3279__, new_new_n3280__, new_new_n3281__,
    new_new_n3282__, new_new_n3283__, new_new_n3284__, new_new_n3285__,
    new_new_n3286__, new_new_n3287__, new_new_n3288__, new_new_n3289__,
    new_new_n3290__, new_new_n3291__, new_new_n3292__, new_new_n3293__,
    new_new_n3294__, new_new_n3295__, new_new_n3296__, new_new_n3297__,
    new_new_n3298__, new_new_n3299__, new_new_n3300__, new_new_n3301__,
    new_new_n3302__, new_new_n3303__, new_new_n3304__, new_new_n3305__,
    new_new_n3306__, new_new_n3307__, new_new_n3308__, new_new_n3309__,
    new_new_n3310__, new_new_n3311__, new_new_n3312__, new_new_n3313__,
    new_new_n3314__, new_new_n3315__, new_new_n3316__, new_new_n3317__,
    new_new_n3318__, new_new_n3319__, new_new_n3320__, new_new_n3321__,
    new_new_n3322__, new_new_n3323__, new_new_n3324__, new_new_n3325__,
    new_new_n3326__, new_new_n3327__, new_new_n3328__, new_new_n3329__,
    new_new_n3330__, new_new_n3331__, new_new_n3332__, new_new_n3333__,
    new_new_n3334__, new_new_n3335__, new_new_n3336__, new_new_n3337__,
    new_new_n3338__, new_new_n3339__, new_new_n3340__, new_new_n3341__,
    new_new_n3342__, new_new_n3343__, new_new_n3344__, new_new_n3345__,
    new_new_n3346__, new_new_n3347__, new_new_n3348__, new_new_n3349__,
    new_new_n3350__, new_new_n3351__, new_new_n3352__, new_new_n3353__,
    new_new_n3354__, new_new_n3355__, new_new_n3356__, new_new_n3357__,
    new_new_n3358__, new_new_n3359__, new_new_n3360__, new_new_n3361__,
    new_new_n3362__, new_new_n3363__, new_new_n3364__, new_new_n3365__,
    new_new_n3366__, new_new_n3367__, new_new_n3368__, new_new_n3369__,
    new_new_n3370__, new_new_n3371__, new_new_n3372__, new_new_n3373__,
    new_new_n3374__, new_new_n3375__, new_new_n3376__, new_new_n3377__,
    new_new_n3378__, new_new_n3379__, new_new_n3380__, new_new_n3381__,
    new_new_n3382__, new_new_n3383__, new_new_n3384__, new_new_n3385__,
    new_new_n3386__, new_new_n3387__, new_new_n3388__, new_new_n3389__,
    new_new_n3390__, new_new_n3391__, new_new_n3392__, new_new_n3393__,
    new_new_n3394__, new_new_n3395__, new_new_n3396__, new_new_n3397__,
    new_new_n3398__, new_new_n3399__, new_new_n3400__, new_new_n3401__,
    new_new_n3402__, new_new_n3403__, new_new_n3404__, new_new_n3405__,
    new_new_n3406__, new_new_n3407__, new_new_n3408__, new_new_n3409__,
    new_new_n3410__, new_new_n3411__, new_new_n3412__, new_new_n3413__,
    new_new_n3414__, new_new_n3415__, new_new_n3416__, new_new_n3417__,
    new_new_n3418__, new_new_n3419__, new_new_n3420__, new_new_n3421__,
    new_new_n3422__, new_new_n3423__, new_new_n3424__, new_new_n3425__,
    new_new_n3426__, new_new_n3427__, new_new_n3428__, new_new_n3429__,
    new_new_n3430__, new_new_n3431__, new_new_n3432__, new_new_n3433__,
    new_new_n3434__, new_new_n3435__, new_new_n3436__, new_new_n3437__,
    new_new_n3438__, new_new_n3439__, new_new_n3440__, new_new_n3441__,
    new_new_n3442__, new_new_n3443__, new_new_n3444__, new_new_n3445__,
    new_new_n3446__, new_new_n3447__, new_new_n3448__, new_new_n3449__,
    new_new_n3450__, new_new_n3451__, new_new_n3452__, new_new_n3453__,
    new_new_n3454__, new_new_n3455__, new_new_n3456__, new_new_n3457__,
    new_new_n3458__, new_new_n3459__, new_new_n3460__, new_new_n3461__,
    new_new_n3462__, new_new_n3463__, new_new_n3464__, new_new_n3465__,
    new_new_n3466__, new_new_n3467__, new_new_n3468__, new_new_n3469__,
    new_new_n3470__, new_new_n3471__, new_new_n3472__, new_new_n3473__,
    new_new_n3474__, new_new_n3475__, new_new_n3476__, new_new_n3477__,
    new_new_n3478__, new_new_n3479__, new_new_n3480__, new_new_n3481__,
    new_new_n3482__, new_new_n3483__, new_new_n3484__, new_new_n3485__,
    new_new_n3486__, new_new_n3487__, new_new_n3488__, new_new_n3489__,
    new_new_n3490__, new_new_n3491__, new_new_n3492__, new_new_n3493__,
    new_new_n3494__, new_new_n3495__, new_new_n3496__, new_new_n3497__,
    new_new_n3498__, new_new_n3499__, new_new_n3500__, new_new_n3501__,
    new_new_n3502__, new_new_n3503__, new_new_n3504__, new_new_n3505__,
    new_new_n3506__, new_new_n3507__, new_new_n3508__, new_new_n3509__,
    new_new_n3510__, new_new_n3511__, new_new_n3512__, new_new_n3513__,
    new_new_n3514__, new_new_n3515__, new_new_n3516__, new_new_n3517__,
    new_new_n3518__, new_new_n3519__, new_new_n3520__, new_new_n3521__,
    new_new_n3522__, new_new_n3523__, new_new_n3524__, new_new_n3525__,
    new_new_n3526__, new_new_n3527__, new_new_n3528__, new_new_n3529__,
    new_new_n3530__, new_new_n3531__, new_new_n3532__, new_new_n3533__,
    new_new_n3534__, new_new_n3535__, new_new_n3536__, new_new_n3537__,
    new_new_n3538__, new_new_n3539__, new_new_n3540__, new_new_n3541__,
    new_new_n3542__, new_new_n3543__, new_new_n3544__, new_new_n3545__,
    new_new_n3546__, new_new_n3547__, new_new_n3548__, new_new_n3549__,
    new_new_n3550__, new_new_n3551__, new_new_n3552__, new_new_n3553__,
    new_new_n3554__, new_new_n3555__, new_new_n3556__, new_new_n3557__,
    new_new_n3558__, new_new_n3559__, new_new_n3560__, new_new_n3561__,
    new_new_n3562__, new_new_n3563__, new_new_n3564__, new_new_n3565__,
    new_new_n3566__, new_new_n3567__, new_new_n3568__, new_new_n3569__,
    new_new_n3570__, new_new_n3571__, new_new_n3572__, new_new_n3573__,
    new_new_n3574__, new_new_n3575__, new_new_n3576__, new_new_n3577__,
    new_new_n3578__, new_new_n3579__, new_new_n3580__, new_new_n3581__,
    new_new_n3582__, new_new_n3583__, new_new_n3584__, new_new_n3585__,
    new_new_n3586__, new_new_n3587__, new_new_n3588__, new_new_n3589__,
    new_new_n3590__, new_new_n3591__, new_new_n3592__, new_new_n3593__,
    new_new_n3594__, new_new_n3595__, new_new_n3596__, new_new_n3597__,
    new_new_n3598__, new_new_n3599__, new_new_n3600__, new_new_n3601__,
    new_new_n3602__, new_new_n3603__, new_new_n3604__, new_new_n3605__,
    new_new_n3606__, new_new_n3607__, new_new_n3608__, new_new_n3609__,
    new_new_n3610__, new_new_n3611__, new_new_n3612__, new_new_n3613__,
    new_new_n3614__, new_new_n3615__, new_new_n3616__, new_new_n3617__,
    new_new_n3618__, new_new_n3619__, new_new_n3620__, new_new_n3621__,
    new_new_n3622__, new_new_n3623__, new_new_n3624__, new_new_n3625__,
    new_new_n3626__, new_new_n3627__, new_new_n3628__, new_new_n3629__,
    new_new_n3630__, new_new_n3631__, new_new_n3632__, new_new_n3633__,
    new_new_n3634__, new_new_n3635__, new_new_n3636__, new_new_n3637__,
    new_new_n3638__, new_new_n3639__, new_new_n3640__, new_new_n3641__,
    new_new_n3642__, new_new_n3643__, new_new_n3644__, new_new_n3645__,
    new_new_n3646__, new_new_n3647__, new_new_n3648__, new_new_n3649__,
    new_new_n3650__, new_new_n3651__, new_new_n3652__, new_new_n3653__,
    new_new_n3654__, new_new_n3655__, new_new_n3656__, new_new_n3657__,
    new_new_n3658__, new_new_n3659__, new_new_n3660__, new_new_n3661__,
    new_new_n3662__, new_new_n3663__, new_new_n3664__, new_new_n3665__,
    new_new_n3666__, new_new_n3667__, new_new_n3668__, new_new_n3669__,
    new_new_n3670__, new_new_n3671__, new_new_n3672__, new_new_n3673__,
    new_new_n3674__, new_new_n3675__, new_new_n3676__, new_new_n3677__,
    new_new_n3678__, new_new_n3679__, new_new_n3680__, new_new_n3681__,
    new_new_n3682__, new_new_n3683__, new_new_n3684__, new_new_n3685__,
    new_new_n3686__, new_new_n3687__, new_new_n3688__, new_new_n3689__,
    new_new_n3690__, new_new_n3691__, new_new_n3692__, new_new_n3693__,
    new_new_n3694__, new_new_n3695__, new_new_n3696__, new_new_n3697__,
    new_new_n3698__, new_new_n3699__, new_new_n3700__, new_new_n3701__,
    new_new_n3702__, new_new_n3703__, new_new_n3704__, new_new_n3705__,
    new_new_n3706__, new_new_n3707__, new_new_n3708__, new_new_n3709__,
    new_new_n3710__, new_new_n3711__, new_new_n3712__, new_new_n3713__,
    new_new_n3714__, new_new_n3715__, new_new_n3716__, new_new_n3717__,
    new_new_n3718__, new_new_n3719__, new_new_n3720__, new_new_n3721__,
    new_new_n3722__, new_new_n3723__, new_new_n3724__, new_new_n3725__,
    new_new_n3726__, new_new_n3727__, new_new_n3728__, new_new_n3729__,
    new_new_n3730__, new_new_n3731__, new_new_n3732__, new_new_n3733__,
    new_new_n3734__, new_new_n3735__, new_new_n3736__, new_new_n3737__,
    new_new_n3738__, new_new_n3739__, new_new_n3740__, new_new_n3741__,
    new_new_n3742__, new_new_n3743__, new_new_n3744__, new_new_n3745__,
    new_new_n3746__, new_new_n3747__, new_new_n3748__, new_new_n3749__,
    new_new_n3750__, new_new_n3751__, new_new_n3752__, new_new_n3753__,
    new_new_n3754__, new_new_n3755__, new_new_n3756__, new_new_n3757__,
    new_new_n3758__, new_new_n3759__, new_new_n3760__, new_new_n3761__,
    new_new_n3762__, new_new_n3763__, new_new_n3764__, new_new_n3765__,
    new_new_n3766__, new_new_n3767__, new_new_n3768__, new_new_n3769__,
    new_new_n3770__, new_new_n3771__, new_new_n3772__, new_new_n3773__,
    new_new_n3774__, new_new_n3775__, new_new_n3776__, new_new_n3777__,
    new_new_n3778__, new_new_n3779__, new_new_n3780__, new_new_n3781__,
    new_new_n3782__, new_new_n3783__, new_new_n3784__, new_new_n3785__,
    new_new_n3786__, new_new_n3787__, new_new_n3788__, new_new_n3789__,
    new_new_n3790__, new_new_n3791__, new_new_n3792__, new_new_n3793__,
    new_new_n3794__, new_new_n3795__, new_new_n3796__, new_new_n3797__,
    new_new_n3798__, new_new_n3799__, new_new_n3800__, new_new_n3801__,
    new_new_n3802__, new_new_n3803__, new_new_n3804__, new_new_n3805__,
    new_new_n3806__, new_new_n3807__, new_new_n3808__, new_new_n3809__,
    new_new_n3810__, new_new_n3811__, new_new_n4363__, new_new_n4364__,
    new_new_n4365__, new_new_n4366__, new_new_n4367__, new_new_n4368__,
    new_new_n4369__, new_new_n4370__, new_new_n4371__, new_new_n4372__,
    new_new_n4373__, new_new_n4374__, new_new_n4375__, new_new_n4376__,
    new_new_n4377__, new_new_n4378__, new_new_n4379__, new_new_n4380__,
    new_new_n4381__, new_new_n4382__, new_new_n4383__, new_new_n4384__,
    new_new_n4385__, new_new_n4386__, new_new_n4387__, new_new_n4388__,
    new_new_n4389__, new_new_n4390__, new_new_n4391__, new_new_n4392__,
    new_new_n4393__, new_new_n4394__, new_new_n4395__, new_new_n4396__,
    new_new_n4397__, new_new_n4398__, new_new_n4399__, new_new_n4400__,
    new_new_n4401__, new_new_n4402__, new_new_n4403__, new_new_n4404__,
    new_new_n4405__, new_new_n4406__, new_new_n4407__, new_new_n4408__,
    new_new_n4409__, new_new_n4410__, new_new_n4411__, new_new_n4412__,
    new_new_n4413__, new_new_n4414__, new_new_n4415__, new_new_n4416__,
    new_new_n4417__, new_new_n4418__, new_new_n4419__, new_new_n4420__,
    new_new_n4421__, new_new_n4422__, new_new_n4423__, new_new_n4424__,
    new_new_n4425__, new_new_n4426__, new_new_n4427__, new_new_n4428__,
    new_new_n4429__, new_new_n4430__, new_new_n4431__, new_new_n4432__,
    new_new_n4433__, new_new_n4434__, new_new_n4435__, new_new_n4436__,
    new_new_n4437__, new_new_n4438__, new_new_n4439__, new_new_n4440__,
    new_new_n4441__, new_new_n4442__, new_new_n4443__, new_new_n4444__,
    new_new_n4445__, new_new_n4446__, new_new_n4447__, new_new_n4448__,
    new_new_n4449__, new_new_n4450__, new_new_n4451__, new_new_n4452__,
    new_new_n4453__, new_new_n4454__, new_new_n4455__, new_new_n4456__,
    new_new_n4457__, new_new_n4458__, new_new_n4459__, new_new_n4460__,
    new_new_n4461__, new_new_n4462__, new_new_n4463__, new_new_n4464__,
    new_new_n4465__, new_new_n4466__, new_new_n4467__, new_new_n4468__,
    new_new_n4469__, new_new_n4470__, new_new_n4471__, new_new_n4472__,
    new_new_n4473__, new_new_n4474__, new_new_n4475__, new_new_n4476__,
    new_new_n4477__, new_new_n4478__, new_new_n4479__, new_new_n4480__,
    new_new_n4481__, new_new_n4482__, new_new_n4483__, new_new_n4484__,
    new_new_n4485__, new_new_n4486__, new_new_n4487__, new_new_n4488__,
    new_new_n4489__, new_new_n4490__, new_new_n4491__, new_new_n4492__,
    new_new_n4493__, new_new_n4494__, new_new_n4495__, new_new_n4496__,
    new_new_n4497__, new_new_n4498__, new_new_n4499__, new_new_n4500__,
    new_new_n4501__, new_new_n4502__, new_new_n4503__, new_new_n4504__,
    new_new_n4505__, new_new_n4506__, new_new_n4507__, new_new_n4508__,
    new_new_n4509__, new_new_n4510__, new_new_n4511__, new_new_n4512__,
    new_new_n4513__, new_new_n4514__, new_new_n4515__, new_new_n4516__,
    new_new_n4517__, new_new_n4518__, new_new_n4519__, new_new_n4520__,
    new_new_n4521__, new_new_n4522__, new_new_n4523__, new_new_n4524__,
    new_new_n4525__, new_new_n4526__, new_new_n4527__, new_new_n4528__,
    new_new_n4529__, new_new_n4530__, new_new_n4531__, new_new_n4532__,
    new_new_n4533__, new_new_n4534__, new_new_n4535__, new_new_n4536__,
    new_new_n4537__, new_new_n4538__, new_new_n4539__, new_new_n4540__,
    new_new_n4541__, new_new_n4542__, new_new_n4543__, new_new_n4544__,
    new_new_n4545__, new_new_n4546__, new_new_n4547__, new_new_n4548__,
    new_new_n4549__, new_new_n4550__, new_new_n4551__, new_new_n4552__,
    new_new_n4553__, new_new_n4554__, new_new_n4555__, new_new_n4556__,
    new_new_n4557__, new_new_n4558__, new_new_n4559__, new_new_n4560__,
    new_new_n4561__, new_new_n4562__, new_new_n4563__, new_new_n4564__,
    new_new_n4565__, new_new_n4566__, new_new_n4567__, new_new_n4568__,
    new_new_n4569__, new_new_n4570__, new_new_n4571__, new_new_n4572__,
    new_new_n4573__, new_new_n4574__, new_new_n4575__, new_new_n4576__,
    new_new_n4577__, new_new_n4578__, new_new_n4579__, new_new_n4580__,
    new_new_n4581__, new_new_n4582__, new_new_n4583__, new_new_n4584__,
    new_new_n4585__, new_new_n4586__, new_new_n4587__, new_new_n4588__,
    new_new_n4589__, new_new_n4590__, new_new_n4591__, new_new_n4592__,
    new_new_n4593__, new_new_n4594__, new_new_n4595__, new_new_n4596__,
    new_new_n4597__, new_new_n4598__, new_new_n4599__, new_new_n4600__,
    new_new_n4601__, new_new_n4602__, new_new_n4603__, new_new_n4604__,
    new_new_n4605__, new_new_n4606__, new_new_n4607__, new_new_n4608__,
    new_new_n4609__, new_new_n4610__, new_new_n4611__, new_new_n4612__,
    new_new_n4613__, new_new_n4614__, new_new_n4615__, new_new_n4616__,
    new_new_n4617__, new_new_n4618__, new_new_n4619__, new_new_n4620__,
    new_new_n4621__, new_new_n4622__, new_new_n4623__, new_new_n4624__,
    new_new_n4625__, new_new_n4626__, new_new_n4627__, new_new_n4628__,
    new_new_n4629__, new_new_n4630__, new_new_n4631__, new_new_n4632__,
    new_new_n4633__, new_new_n4634__, new_new_n4635__, new_new_n4636__,
    new_new_n4637__, new_new_n4638__, new_new_n4639__, new_new_n4640__,
    new_new_n4641__, new_new_n4642__, new_new_n4643__, new_new_n4644__,
    new_new_n4645__, new_new_n4646__, new_new_n4647__, new_new_n4648__,
    new_new_n4649__, new_new_n4650__, new_new_n4651__, new_new_n4652__,
    new_new_n4653__, new_new_n4654__, new_new_n4655__, new_new_n4656__,
    new_new_n4657__, new_new_n4658__, new_new_n4659__, new_new_n4660__,
    new_new_n4661__, new_new_n4662__, new_new_n4663__, new_new_n4664__,
    new_new_n4665__, new_new_n4666__, new_new_n4667__, new_new_n4668__,
    new_new_n4669__, new_new_n4670__, new_new_n4671__, new_new_n4672__,
    new_new_n4673__, new_new_n4674__, new_new_n4675__, new_new_n4676__,
    new_new_n4677__, new_new_n4678__, new_new_n4679__, new_new_n4680__,
    new_new_n4681__, new_new_n4682__, new_new_n4683__, new_new_n4684__,
    new_new_n4685__, new_new_n4686__, new_new_n4687__, new_new_n4688__,
    new_new_n4689__, new_new_n4690__, new_new_n4691__, new_new_n4692__,
    new_new_n4693__, new_new_n4694__, new_new_n4695__, new_new_n4696__,
    new_new_n4697__, new_new_n4698__, new_new_n4699__, new_new_n4700__,
    new_new_n4701__, new_new_n4702__, new_new_n4703__, new_new_n4704__,
    new_new_n4705__, new_new_n4706__, new_new_n4707__, new_new_n4708__,
    new_new_n4709__, new_new_n4710__, new_new_n4711__, new_new_n4712__,
    new_new_n4713__, new_new_n4714__, new_new_n4715__, new_new_n4716__,
    new_new_n4717__, new_new_n4718__, new_new_n4719__, new_new_n4720__,
    new_new_n4721__, new_new_n4722__, new_new_n4723__, new_new_n4724__,
    new_new_n4725__, new_new_n4726__, new_new_n4727__, new_new_n4728__,
    new_new_n4729__, new_new_n4730__, new_new_n4731__, new_new_n4732__,
    new_new_n4733__, new_new_n4734__, new_new_n4735__, new_new_n4736__,
    new_new_n4737__, new_new_n4738__, new_new_n4739__, new_new_n4740__,
    new_new_n4741__, new_new_n4742__, new_new_n4743__, new_new_n4744__,
    new_new_n4745__, new_new_n4746__, new_new_n4747__, new_new_n4748__,
    new_new_n4749__, new_new_n4750__, new_new_n4751__, new_new_n4752__,
    new_new_n4753__, new_new_n4754__, new_new_n4755__, new_new_n4756__,
    new_new_n4757__, new_new_n4758__, new_new_n4759__, new_new_n4760__,
    new_new_n4761__, new_new_n4762__, new_new_n4763__, new_new_n4764__,
    new_new_n4765__, new_new_n4766__, new_new_n4767__, new_new_n4768__,
    new_new_n4769__, new_new_n4770__, new_new_n4771__, new_new_n4772__,
    new_new_n4773__, new_new_n4774__, new_new_n4775__, new_new_n4776__,
    new_new_n4777__, new_new_n4778__, new_new_n4779__, new_new_n4780__,
    new_new_n4781__, new_new_n4782__, new_new_n4783__, new_new_n4784__,
    new_new_n4785__, new_new_n4786__, new_new_n4787__, new_new_n4788__,
    new_new_n4789__, new_new_n4790__, new_new_n4791__, new_new_n4792__,
    new_new_n4793__, new_new_n4794__, new_new_n4795__, new_new_n4796__,
    new_new_n4797__, new_new_n4798__, new_new_n4799__, new_new_n4800__,
    new_new_n4801__, new_new_n4802__, new_new_n4803__, new_new_n4804__,
    new_new_n4805__, new_new_n4806__, new_new_n4807__, new_new_n4808__,
    new_new_n4809__, new_new_n4810__, new_new_n4811__, new_new_n4812__,
    new_new_n4813__, new_new_n4814__, new_new_n4815__, new_new_n4816__,
    new_new_n4817__, new_new_n4818__, new_new_n4819__, new_new_n4820__,
    new_new_n4821__, new_new_n4822__, new_new_n4823__, new_new_n4824__,
    new_new_n4825__, new_new_n4826__, new_new_n4827__, new_new_n4828__,
    new_new_n4829__, new_new_n4830__, new_new_n4831__, new_new_n4832__,
    new_new_n4833__, new_new_n4834__, new_new_n4835__, new_new_n4836__,
    new_new_n4837__, new_new_n4838__, new_new_n4839__, new_new_n4840__,
    new_new_n4841__, new_new_n4842__, new_new_n4843__, new_new_n4844__,
    new_new_n4845__, new_new_n4846__, new_new_n4847__, new_new_n4848__,
    new_new_n4849__, new_new_n4850__, new_new_n4851__, new_new_n4852__,
    new_new_n4853__, new_new_n4854__, new_new_n4855__, new_new_n4856__,
    new_new_n4857__, new_new_n4858__, new_new_n4859__, new_new_n4860__,
    new_new_n4861__, new_new_n4862__, new_new_n4863__, new_new_n4864__,
    new_new_n4865__, new_new_n4866__, new_new_n4867__, new_new_n4868__,
    new_new_n4869__, new_new_n4870__, new_new_n4871__, new_new_n4872__,
    new_new_n4873__, new_new_n4874__, new_new_n4875__, new_new_n4876__,
    new_new_n4877__, new_new_n4878__, new_new_n4879__, new_new_n4880__,
    new_new_n4881__, new_new_n4882__, new_new_n4883__, new_new_n4884__,
    new_new_n4885__, new_new_n4886__, new_new_n4887__, new_new_n4888__,
    new_new_n4889__, new_new_n4890__, new_new_n4891__, new_new_n4892__,
    new_new_n4893__, new_new_n4894__, new_new_n4895__, new_new_n4896__,
    new_new_n4897__, new_new_n4898__, new_new_n4899__, new_new_n4900__,
    new_new_n4901__, new_new_n4902__, new_new_n4903__, new_new_n4904__,
    new_new_n4905__, new_new_n4906__, new_new_n4907__, new_new_n4908__,
    new_new_n4909__, new_new_n4910__, new_new_n4911__, new_new_n4912__,
    new_new_n4913__, new_new_n4914__, new_new_n4915__, new_new_n4916__,
    new_new_n4917__, new_new_n4918__, new_new_n4919__, new_new_n4920__,
    new_new_n4921__, new_new_n4922__, new_new_n4923__, new_new_n4924__,
    new_new_n4925__, new_new_n4926__, new_new_n4927__, new_new_n4928__,
    new_new_n4929__, new_new_n4930__, new_new_n4931__, new_new_n4932__,
    new_new_n4933__, new_new_n4934__, new_new_n4935__, new_new_n4936__,
    new_new_n4937__, new_new_n4938__, new_new_n4939__, new_new_n4940__,
    new_new_n4941__, new_new_n4942__, new_new_n4943__, new_new_n4944__,
    new_new_n4945__, new_new_n4946__, new_new_n4947__, new_new_n4948__,
    new_new_n4949__, new_new_n4950__, new_new_n4951__, new_new_n4952__,
    new_new_n4953__, new_new_n4954__, new_new_n4955__, new_new_n4956__,
    new_new_n4957__, new_new_n4958__, new_new_n4959__, new_new_n4960__,
    new_new_n4961__, new_new_n4962__, new_new_n4963__, new_new_n4964__,
    new_new_n4965__, new_new_n4966__, new_new_n4967__, new_new_n4968__,
    new_new_n4969__, new_new_n4970__, new_new_n4971__, new_new_n4972__,
    new_new_n4973__, new_new_n4974__, new_new_n4975__, new_new_n4976__,
    new_new_n4977__, new_new_n4978__, new_new_n4979__, new_new_n4980__,
    new_new_n4981__, new_new_n4982__, new_new_n4983__, new_new_n4984__,
    new_new_n4985__, new_new_n4986__, new_new_n4987__, new_new_n4988__,
    new_new_n4989__, new_new_n4990__, new_new_n4991__, new_new_n4992__,
    new_new_n4993__, new_new_n4994__, new_new_n4995__, new_new_n4996__,
    new_new_n4997__, new_new_n4998__, new_new_n4999__, new_new_n5000__,
    new_new_n5001__, new_new_n5002__, new_new_n5003__, new_new_n5004__,
    new_new_n5005__, new_new_n5006__, new_new_n5007__, new_new_n5008__,
    new_new_n5009__, new_new_n5010__, new_new_n5011__, new_new_n5012__,
    new_new_n5013__, new_new_n5014__, new_new_n5015__, new_new_n5016__,
    new_new_n5017__, new_new_n5018__, new_new_n5019__, new_new_n5020__,
    new_new_n5021__, new_new_n5022__, new_new_n5023__, new_new_n5024__,
    new_new_n5025__, new_new_n5026__, new_new_n5027__, new_new_n5028__,
    new_new_n5029__, new_new_n5030__, new_new_n5031__, new_new_n5032__,
    new_new_n5033__, new_new_n5034__, new_new_n5035__, new_new_n5036__,
    new_new_n5037__, new_new_n5038__, new_new_n5039__, new_new_n5040__,
    new_new_n5041__, new_new_n5042__, new_new_n5043__, new_new_n5044__,
    new_new_n5045__, new_new_n5046__, new_new_n5047__, new_new_n5048__,
    new_new_n5049__, new_new_n5050__, new_new_n5051__, new_new_n5052__,
    new_new_n5053__, new_new_n5054__, new_new_n5055__, new_new_n5056__,
    new_new_n5057__, new_new_n5058__, new_new_n5059__, new_new_n5060__,
    new_new_n5061__, new_new_n5062__, new_new_n5063__, new_new_n5064__,
    new_new_n5065__, new_new_n5066__, new_new_n5067__, new_new_n5068__,
    new_new_n5069__, new_new_n5070__, new_new_n5071__, new_new_n5072__,
    new_new_n5073__, new_new_n5074__, new_new_n5075__, new_new_n5076__,
    new_new_n5077__, new_new_n5078__, new_new_n5079__, new_new_n5080__,
    new_new_n5081__, new_new_n5082__, new_new_n5083__, new_new_n5084__,
    new_new_n5085__, new_new_n5086__, new_new_n5087__, new_new_n5088__,
    new_new_n5089__, new_new_n5090__, new_new_n5091__, new_new_n5092__,
    new_new_n5093__, new_new_n5094__, new_new_n5095__, new_new_n5096__,
    new_new_n5097__, new_new_n5098__, new_new_n5099__, new_new_n5100__,
    new_new_n5101__, new_new_n5102__, new_new_n5103__, new_new_n5104__,
    new_new_n5105__, new_new_n5106__, new_new_n5107__, new_new_n5108__,
    new_new_n5109__, new_new_n5110__, new_new_n5111__, new_new_n5112__,
    new_new_n5113__, new_new_n5114__, new_new_n5115__, new_new_n5116__,
    new_new_n5117__, new_new_n5118__, new_new_n5119__, new_new_n5120__,
    new_new_n5121__, new_new_n5122__, new_new_n5123__, new_new_n5124__,
    new_new_n5125__, new_new_n5126__, new_new_n5127__, new_new_n5128__,
    new_new_n5129__, new_new_n5130__, new_new_n5131__, new_new_n5132__,
    new_new_n5133__, new_new_n5134__, new_new_n5135__, new_new_n5136__,
    new_new_n5137__, new_new_n5138__, new_new_n5139__, new_new_n5140__,
    new_new_n5141__, new_new_n5142__, new_new_n5143__, new_new_n5144__,
    new_new_n5145__, new_new_n5146__, new_new_n5147__, new_new_n5148__,
    new_new_n5149__, new_new_n5150__, new_new_n5151__, new_new_n5152__,
    new_new_n5153__, new_new_n5154__, new_new_n5155__, new_new_n5156__,
    new_new_n5157__, new_new_n5158__, new_new_n5159__, new_new_n5160__,
    new_new_n5161__, new_new_n5162__, new_new_n5163__, new_new_n5164__,
    new_new_n5165__, new_new_n5166__, new_new_n5167__, new_new_n5168__,
    new_new_n5169__, new_new_n5170__, new_new_n5171__, new_new_n5172__,
    new_new_n5173__, new_new_n5174__, new_new_n5175__, new_new_n5176__,
    new_new_n5177__, new_new_n5178__, new_new_n5179__, new_new_n5180__,
    new_new_n5181__, new_new_n5182__, new_new_n5183__, new_new_n5184__,
    new_new_n5185__, new_new_n5186__, new_new_n5187__, new_new_n5188__,
    new_new_n5189__, new_new_n5190__, new_new_n5191__, new_new_n5192__,
    new_new_n5193__, new_new_n5194__, new_new_n5195__, new_new_n5196__,
    new_new_n5197__, new_new_n5198__, new_new_n5199__, new_new_n5200__,
    new_new_n5201__, new_new_n5202__, new_new_n5203__, new_new_n5204__,
    new_new_n5205__, new_new_n5206__, new_new_n5207__, new_new_n5208__,
    new_new_n5209__, new_new_n5210__, new_new_n5211__, new_new_n5212__,
    new_new_n5213__, new_new_n5214__, new_new_n5215__, new_new_n5216__,
    new_new_n5217__, new_new_n5218__, new_new_n5219__, new_new_n5220__,
    new_new_n5221__, new_new_n5222__, new_new_n5223__, new_new_n5224__,
    new_new_n5225__, new_new_n5226__, new_new_n5227__, new_new_n5228__,
    new_new_n5229__, new_new_n5230__, new_new_n5231__, new_new_n5232__,
    new_new_n5233__, new_new_n5234__, new_new_n5235__, new_new_n5236__,
    new_new_n5237__, new_new_n5238__, new_new_n5239__, new_new_n5240__,
    new_new_n5241__, new_new_n5242__, new_new_n5243__, new_new_n5244__,
    new_new_n5245__, new_new_n5246__, new_new_n5247__, new_new_n5248__,
    new_new_n5249__, new_new_n5250__, new_new_n5251__, new_new_n5252__,
    new_new_n5253__, new_new_n5254__, new_new_n5255__, new_new_n5256__,
    new_new_n5257__, new_new_n5258__, new_new_n5259__, new_new_n5260__,
    new_new_n5261__, new_new_n5262__, new_new_n5263__, new_new_n5264__,
    new_new_n5265__, new_new_n5266__, new_new_n5267__, new_new_n5268__,
    new_new_n5269__, new_new_n5270__, new_new_n5271__, new_new_n5272__,
    new_new_n5273__, new_new_n5274__, new_new_n5275__, new_new_n5276__,
    new_new_n5277__, new_new_n5278__, new_new_n5279__, new_new_n5280__,
    new_new_n5281__, new_new_n5282__, new_new_n5283__, new_new_n5284__,
    new_new_n5285__, new_new_n5286__, new_new_n5287__, new_new_n5288__,
    new_new_n5289__, new_new_n5290__, new_new_n5291__, new_new_n5292__,
    new_new_n5293__, new_new_n5294__, new_new_n5295__, new_new_n5296__,
    new_new_n5297__, new_new_n5298__, new_new_n5299__, new_new_n5300__,
    new_new_n5301__, new_new_n5302__, new_new_n5303__, new_new_n5304__,
    new_new_n5305__, new_new_n5306__, new_new_n5307__, new_new_n5308__,
    new_new_n5309__, new_new_n5310__, new_new_n5311__, new_new_n5312__,
    new_new_n5313__, new_new_n5314__, new_new_n5315__, new_new_n5316__,
    new_new_n5317__, new_new_n5318__, new_new_n5319__, new_new_n5320__,
    new_new_n5321__, new_new_n5322__, new_new_n5323__, new_new_n5324__,
    new_new_n5325__, new_new_n5326__, new_new_n5327__, new_new_n5328__,
    new_new_n5329__, new_new_n5330__, new_new_n5331__, new_new_n5332__,
    new_new_n5333__, new_new_n5334__, new_new_n5335__, new_new_n5336__,
    new_new_n5337__, new_new_n5338__, new_new_n5339__, new_new_n5340__,
    new_new_n5341__, new_new_n5342__, new_new_n5343__, new_new_n5344__,
    new_new_n5345__, new_new_n5346__, new_new_n5347__, new_new_n5348__,
    new_new_n5349__, new_new_n5350__, new_new_n5351__, new_new_n5352__,
    new_new_n5353__, new_new_n5354__, new_new_n5355__, new_new_n5356__,
    new_new_n5357__, new_new_n5358__, new_new_n5359__, new_new_n5360__,
    new_new_n5361__, new_new_n5362__, new_new_n5363__, new_new_n5364__,
    new_new_n5365__, new_new_n5366__, new_new_n5367__, new_new_n5368__,
    new_new_n5369__, new_new_n5370__, new_new_n5371__, new_new_n5372__,
    new_new_n5373__, new_new_n5374__, new_new_n5375__, new_new_n5376__,
    new_new_n5377__, new_new_n5378__, new_new_n5379__, new_new_n5380__,
    new_new_n5381__, new_new_n5382__, new_new_n5383__, new_new_n5384__,
    new_new_n5385__, new_new_n5386__, new_new_n5387__, new_new_n5388__,
    new_new_n5389__, new_new_n5390__, new_new_n5391__, new_new_n5392__,
    new_new_n5393__, new_new_n5394__, new_new_n5395__, new_new_n5396__,
    new_new_n5397__, new_new_n5398__, new_new_n5399__, new_new_n5400__,
    new_new_n5401__, new_new_n5402__, new_new_n5403__, new_new_n5404__,
    new_new_n5405__, new_new_n5406__, new_new_n5407__, new_new_n5408__,
    new_new_n5409__, new_new_n5410__, new_new_n5411__, new_new_n5412__,
    new_new_n5413__, new_new_n5414__, new_new_n5415__, new_new_n5416__,
    new_new_n5417__, new_new_n5418__, new_new_n5419__, new_new_n5420__,
    new_new_n5421__, new_new_n5422__, new_new_n5423__, new_new_n5424__,
    new_new_n5425__, new_new_n5426__, new_new_n5427__, new_new_n5428__,
    new_new_n5429__, new_new_n5430__, new_new_n5431__, new_new_n5432__,
    new_new_n5433__, new_new_n5434__, new_new_n5435__, new_new_n5436__,
    new_new_n5437__, new_new_n5438__, new_new_n5439__, new_new_n5440__,
    new_new_n5441__, new_new_n5442__, new_new_n5443__, new_new_n5444__,
    new_new_n5445__, new_new_n5446__, new_new_n5447__, new_new_n5448__,
    new_new_n5449__, new_new_n5450__, new_new_n5451__, new_new_n5452__,
    new_new_n5453__, new_new_n5454__, new_new_n5455__, new_new_n5456__,
    new_new_n5457__, new_new_n5458__, new_new_n5459__, new_new_n5460__,
    new_new_n5461__, new_new_n5462__, new_new_n5463__, new_new_n5464__,
    new_new_n5465__, new_new_n5466__, new_new_n5467__, new_new_n5468__,
    new_new_n5469__, new_new_n5470__, new_new_n5471__, new_new_n5472__,
    new_new_n5473__, new_new_n5474__, new_new_n5475__, new_new_n5476__,
    new_new_n5477__, new_new_n5478__, new_new_n5479__, new_new_n5480__,
    new_new_n5481__, new_new_n5482__, new_new_n5483__, new_new_n5484__,
    new_new_n5485__, new_new_n5486__, new_new_n5487__, new_new_n5488__,
    new_new_n5489__, new_new_n5490__, new_new_n5491__, new_new_n5492__,
    new_new_n5493__, new_new_n5494__, new_new_n5495__, new_new_n5496__,
    new_new_n5497__, new_new_n5498__, new_new_n5499__, new_new_n5500__,
    new_new_n5501__, new_new_n5502__, new_new_n5503__, new_new_n5504__,
    new_new_n5505__, new_new_n5506__, new_new_n5507__, new_new_n5508__,
    new_new_n5509__, new_new_n5510__, new_new_n5511__, new_new_n5512__,
    new_new_n5513__, new_new_n5514__, new_new_n5515__, new_new_n5516__,
    new_new_n5517__, new_new_n5518__, new_new_n5519__, new_new_n5520__,
    new_new_n5521__, new_new_n5522__, new_new_n5523__, new_new_n5524__,
    new_new_n5525__, new_new_n5526__, new_new_n5527__, new_new_n5528__,
    new_new_n5529__, new_new_n5530__, new_new_n5531__, new_new_n5532__,
    new_new_n5533__, new_new_n5534__, new_new_n5535__, new_new_n5536__,
    new_new_n5537__, new_new_n5538__, new_new_n5539__, new_new_n5540__,
    new_new_n5541__, new_new_n5542__, new_new_n5543__, new_new_n5544__,
    new_new_n5545__, new_new_n5546__, new_new_n5547__, new_new_n5548__,
    new_new_n5549__, new_new_n5550__, new_new_n5551__, new_new_n5552__,
    new_new_n5553__, new_new_n5554__, new_new_n5555__, new_new_n5556__,
    new_new_n5557__, new_new_n5558__, new_new_n5559__, new_new_n5560__,
    new_new_n5561__, new_new_n5562__, new_new_n5563__, new_new_n5564__,
    new_new_n5565__, new_new_n5566__, new_new_n5567__, new_new_n5568__,
    new_new_n5569__, new_new_n5570__, new_new_n5571__, new_new_n5572__,
    new_new_n5573__, new_new_n5574__, new_new_n5575__, new_new_n5576__,
    new_new_n5577__, new_new_n5578__, new_new_n5579__, new_new_n5580__,
    new_new_n5581__, new_new_n5582__, new_new_n5583__, new_new_n5584__,
    new_new_n5585__, new_new_n5586__, new_new_n5587__, new_new_n5588__,
    new_new_n5589__, new_new_n5590__, new_new_n5591__, new_new_n5592__,
    new_new_n5593__, new_new_n5594__, new_new_n5595__, new_new_n5596__,
    new_new_n5597__, new_new_n5598__, new_new_n5599__, new_new_n5600__,
    new_new_n5601__, new_new_n5602__, new_new_n5603__, new_new_n5604__,
    new_new_n5605__, new_new_n5606__, new_new_n5607__, new_new_n5608__,
    new_new_n5609__, n8948, n8951, n8954, n8957, n8960, n8963, n8966,
    n8969, n8972, n8975, n8978, n8981, n8984, n8987, n8990, n8993, n8996,
    n8999, n9002, n9005, n9008, n9011, n9014, n9017, n9020, n9023, n9026,
    n9029, n9032, n9035, n9038, n9041, n9044, n9047, n9050, n9053, n9056,
    n9059, n9062, n9065, n9068, n9071, n9074, n9077, n9080, n9083, n9086,
    n9089, n9092, n9095, n9098, n9101, n9104, n9107, n9110, n9113, n9116,
    n9119, n9122, n9125, n9128, n9131, n9134, n9137, n9140, n9143, n9146,
    n9149, n9152, n9155, n9158, n9161, n9164, n9167, n9170, n9173, n9176,
    n9179, n9182, n9185, n9188, n9191, n9194, n9197, n9200, n9203, n9206,
    n9209, n9212, n9215, n9218, n9221, n9224, n9227, n9230, n9233, n9236,
    n9239, n9242, n9245, n9248, n9251, n9254, n9257, n9260, n9263, n9266,
    n9269, n9272, n9275, n9278, n9281, n9284, n9287, n9290, n9293, n9296,
    n9299, n9302, n9305, n9308, n9311, n9314, n9317, n9320, n9323, n9326,
    n9329, n9332, n9335, n9338, n9341, n9344, n9347, n9350, n9353, n9356,
    n9359, n9362, n9365, n9368, n9371, n9374, n9377, n9380, n9383, n9386,
    n9389, n9392, n9395, n9398, n9401, n9404, n9407, n9410, n9413, n9416,
    n9419, n9422, n9425, n9428, n9431, n9434, n9437, n9440, n9443, n9446,
    n9449, n9452, n9455, n9458, n9461, n9464, n9467, n9470, n9473, n9476,
    n9479, n9482, n9485, n9488, n9491, n9494, n9497, n9500, n9503, n9506,
    n9509, n9512, n9515, n9518, n9521, n9524, n9527, n9530, n9533, n9536,
    n9539, n9542, n9545, n9548, n9551, n9554, n9557, n9560, n9563, n9566,
    n9569, n9572, n9575, n9578, n9581, n9584, n9587, n9590, n9593, n9596,
    n9599, n9602, n9605, n9608, n9611, n9614, n9617, n9620, n9623, n9626,
    n9629, n9632, n9635, n9638, n9641, n9644, n9647, n9650, n9653, n9656,
    n9659, n9662, n9665, n9668, n9671, n9674, n9677, n9680, n9683, n9686,
    n9689, n9692, n9695, n9698, n9701, n9704, n9707, n9710, n9713, n9716,
    n9719, n9722, n9725, n9728, n9731, n9734, n9737, n9740, n9743, n9746,
    n9749, n9752, n9755, n9758, n9761, n9764, n9767, n9770, n9773, n9776,
    n9779, n9782, n9785, n9788, n9791, n9794, n9797, n9800, n9803, n9806,
    n9809, n9812, n9815, n9818, n9821, n9824, n9827, n9830, n9833, n9836,
    n9839, n9842, n9845, n9848, n9851, n9854, n9857, n9860, n9863, n9866,
    n9869, n9872, n9875, n9878, n9881, n9884, n9887, n9890, n9893, n9896,
    n9899, n9902, n9905, n9908, n9911, n9914, n9917, n9920, n9923, n9926,
    n9929, n9932, n9935, n9938, n9941, n9944, n9947, n9950, n9953, n9956,
    n9959, n9962, n9965, n9968, n9971, n9974, n9977, n9980, n9983, n9986,
    n9989, n9992, n9995, n9998, n10001, n10004, n10007, n10010, n10013,
    n10016, n10019, n10022, n10025, n10028, n10031, n10034, n10037, n10040,
    n10043, n10046, n10049, n10052, n10055, n10058, n10061, n10064, n10067,
    n10070, n10073, n10076, n10079, n10082, n10085, n10088, n10091, n10094,
    n10097, n10100, n10103, n10106, n10109, n10112, n10115, n10118, n10121,
    n10124, n10127, n10130, n10133, n10136, n10139, n10142, n10145, n10148,
    n10151, n10154, n10157, n10160, n10163, n10166, n10169, n10172, n10175,
    n10178, n10181, n10184, n10187, n10190, n10193, n10196, n10199, n10202,
    n10205, n10208, n10211, n10214, n10217, n10220, n10223, n10226, n10229,
    n10232, n10235, n10238, n10241, n10244, n10247, n10250, n10253, n10256,
    n10259, n10262, n10265, n10268, n10271, n10274, n10277, n10280, n10283,
    n10286, n10289, n10292, n10295, n10298, n10301, n10304, n10307, n10310,
    n10313, n10316, n10319, n10322, n10325, n10328, n10331, n10334, n10337,
    n10340, n10343, n10346, n10349, n10352, n10355, n10358, n10361, n10364,
    n10367, n10370, n10373, n10376, n10379, n10382, n10385, n10388, n10391,
    n10394, n10397, n10400, n10403, n10406, n10409, n10412, n10415, n10418,
    n10421, n10424, n10427, n10430, n10433, n10436, n10439, n10442, n10445,
    n10448, n10451, n10454, n10457, n10460, n10463, n10466, n10469, n10472,
    n10475, n10478, n10481, n10484, n10487, n10490, n10493, n10496, n10499,
    n10502, n10505, n10508, n10511, n10514, n10517, n10520, n10523, n10526,
    n10529, n10532;
  buf1  g0000(.din(G1), .dout(new_new_n1131__));
  buf1  g0001(.din(G2), .dout(new_new_n1133__));
  buf1  g0002(.din(G3), .dout(new_new_n1135__));
  not1  g0003(.din(G3), .dout(new_new_n1136__));
  buf1  g0004(.din(G4), .dout(new_new_n1137__));
  buf1  g0005(.din(G5), .dout(new_new_n1139__));
  buf1  g0006(.din(G6), .dout(new_new_n1141__));
  buf1  g0007(.din(G7), .dout(new_new_n1143__));
  buf1  g0008(.din(G8), .dout(new_new_n1145__));
  buf1  g0009(.din(G9), .dout(new_new_n1147__));
  buf1  g0010(.din(G10), .dout(new_new_n1149__));
  buf1  g0011(.din(G11), .dout(new_new_n1151__));
  buf1  g0012(.din(G12), .dout(new_new_n1153__));
  buf1  g0013(.din(G13), .dout(new_new_n1155__));
  buf1  g0014(.din(G14), .dout(new_new_n1157__));
  buf1  g0015(.din(G15), .dout(new_new_n1159__));
  buf1  g0016(.din(G16), .dout(new_new_n1161__));
  buf1  g0017(.din(G17), .dout(new_new_n1163__));
  buf1  g0018(.din(G18), .dout(new_new_n1165__));
  buf1  g0019(.din(G19), .dout(new_new_n1167__));
  buf1  g0020(.din(G20), .dout(new_new_n1169__));
  buf1  g0021(.din(G21), .dout(new_new_n1171__));
  buf1  g0022(.din(G22), .dout(new_new_n1173__));
  buf1  g0023(.din(G23), .dout(new_new_n1175__));
  buf1  g0024(.din(G24), .dout(new_new_n1177__));
  buf1  g0025(.din(G25), .dout(new_new_n1179__));
  buf1  g0026(.din(G26), .dout(new_new_n1181__));
  buf1  g0027(.din(G27), .dout(new_new_n1183__));
  buf1  g0028(.din(G28), .dout(new_new_n1185__));
  buf1  g0029(.din(G29), .dout(new_new_n1187__));
  buf1  g0030(.din(G30), .dout(new_new_n1189__));
  buf1  g0031(.din(G31), .dout(new_new_n1191__));
  buf1  g0032(.din(G32), .dout(new_new_n1193__));
  buf1  g0033(.din(G33), .dout(new_new_n1195__));
  buf1  g0034(.din(G34), .dout(new_new_n1197__));
  buf1  g0035(.din(G35), .dout(new_new_n1199__));
  buf1  g0036(.din(G36), .dout(new_new_n1201__));
  buf1  g0037(.din(G37), .dout(new_new_n1203__));
  buf1  g0038(.din(G38), .dout(new_new_n1205__));
  buf1  g0039(.din(G39), .dout(new_new_n1207__));
  buf1  g0040(.din(G40), .dout(new_new_n1209__));
  buf1  g0041(.din(G41), .dout(new_new_n1211__));
  buf1  g0042(.din(G42), .dout(new_new_n1213__));
  buf1  g0043(.din(G43), .dout(new_new_n1215__));
  buf1  g0044(.din(G44), .dout(new_new_n1217__));
  buf1  g0045(.din(G45), .dout(new_new_n1219__));
  buf1  g0046(.din(G46), .dout(new_new_n1221__));
  buf1  g0047(.din(G47), .dout(new_new_n1223__));
  buf1  g0048(.din(G48), .dout(new_new_n1225__));
  buf1  g0049(.din(G49), .dout(new_new_n1227__));
  buf1  g0050(.din(G50), .dout(new_new_n1229__));
  buf1  g0051(.din(n1836_lo), .dout(new_new_n1231__));
  not1  g0052(.din(n1836_lo), .dout(new_new_n1232__));
  not1  g0053(.din(n1872_lo), .dout(new_new_n1234__));
  buf1  g0054(.din(n1884_lo), .dout(new_new_n1235__));
  not1  g0055(.din(n1884_lo), .dout(new_new_n1236__));
  buf1  g0056(.din(n1911_lo), .dout(new_new_n1237__));
  buf1  g0057(.din(n1914_lo), .dout(new_new_n1239__));
  not1  g0058(.din(n1917_lo), .dout(new_new_n1242__));
  buf1  g0059(.din(n1923_lo), .dout(new_new_n1243__));
  buf1  g0060(.din(n1926_lo), .dout(new_new_n1245__));
  not1  g0061(.din(n1929_lo), .dout(new_new_n1248__));
  buf1  g0062(.din(n1935_lo), .dout(new_new_n1249__));
  buf1  g0063(.din(n1938_lo), .dout(new_new_n1251__));
  buf1  g0064(.din(n1947_lo), .dout(new_new_n1253__));
  buf1  g0065(.din(n1950_lo), .dout(new_new_n1255__));
  buf1  g0066(.din(n1959_lo), .dout(new_new_n1257__));
  buf1  g0067(.din(n1962_lo), .dout(new_new_n1259__));
  buf1  g0068(.din(n1971_lo), .dout(new_new_n1261__));
  buf1  g0069(.din(n1974_lo), .dout(new_new_n1263__));
  buf1  g0070(.din(n1983_lo), .dout(new_new_n1265__));
  buf1  g0071(.din(n1995_lo), .dout(new_new_n1267__));
  not1  g0072(.din(n1995_lo), .dout(new_new_n1268__));
  buf1  g0073(.din(n2007_lo), .dout(new_new_n1269__));
  not1  g0074(.din(n2007_lo), .dout(new_new_n1270__));
  buf1  g0075(.din(n2019_lo), .dout(new_new_n1271__));
  not1  g0076(.din(n2019_lo), .dout(new_new_n1272__));
  buf1  g0077(.din(n2031_lo), .dout(new_new_n1273__));
  not1  g0078(.din(n2031_lo), .dout(new_new_n1274__));
  buf1  g0079(.din(n2043_lo), .dout(new_new_n1275__));
  not1  g0080(.din(n2043_lo), .dout(new_new_n1276__));
  buf1  g0081(.din(n2055_lo), .dout(new_new_n1277__));
  not1  g0082(.din(n2055_lo), .dout(new_new_n1278__));
  buf1  g0083(.din(n2064_lo), .dout(new_new_n1279__));
  buf1  g0084(.din(n2067_lo), .dout(new_new_n1281__));
  not1  g0085(.din(n2100_lo), .dout(new_new_n1284__));
  not1  g0086(.din(n2112_lo), .dout(new_new_n1286__));
  not1  g0087(.din(n2124_lo), .dout(new_new_n1288__));
  not1  g0088(.din(n2136_lo), .dout(new_new_n1290__));
  not1  g0089(.din(n2148_lo), .dout(new_new_n1292__));
  not1  g0090(.din(n2160_lo), .dout(new_new_n1294__));
  buf1  g0091(.din(n2163_lo), .dout(new_new_n1295__));
  not1  g0092(.din(n2163_lo), .dout(new_new_n1296__));
  not1  g0093(.din(n2172_lo), .dout(new_new_n1298__));
  buf1  g0094(.din(n2175_lo), .dout(new_new_n1299__));
  not1  g0095(.din(n2184_lo), .dout(new_new_n1302__));
  buf1  g0096(.din(n2223_lo), .dout(new_new_n1303__));
  buf1  g0097(.din(n2235_lo), .dout(new_new_n1305__));
  buf1  g0098(.din(n2238_lo), .dout(new_new_n1307__));
  buf1  g0099(.din(n2247_lo), .dout(new_new_n1309__));
  buf1  g0100(.din(n2250_lo), .dout(new_new_n1311__));
  buf1  g0101(.din(n2259_lo), .dout(new_new_n1313__));
  buf1  g0102(.din(n2262_lo), .dout(new_new_n1315__));
  buf1  g0103(.din(n2271_lo), .dout(new_new_n1317__));
  buf1  g0104(.din(n2274_lo), .dout(new_new_n1319__));
  buf1  g0105(.din(n2283_lo), .dout(new_new_n1321__));
  buf1  g0106(.din(n2286_lo), .dout(new_new_n1323__));
  buf1  g0107(.din(n2295_lo), .dout(new_new_n1325__));
  buf1  g0108(.din(n2298_lo), .dout(new_new_n1327__));
  not1  g0109(.din(n2298_lo), .dout(new_new_n1328__));
  buf1  g0110(.din(n2304_lo), .dout(new_new_n1329__));
  not1  g0111(.din(n2304_lo), .dout(new_new_n1330__));
  buf1  g0112(.din(n2307_lo), .dout(new_new_n1331__));
  not1  g0113(.din(n2307_lo), .dout(new_new_n1332__));
  buf1  g0114(.din(n2331_lo), .dout(new_new_n1333__));
  buf1  g0115(.din(n2334_lo), .dout(new_new_n1335__));
  buf1  g0116(.din(n2337_lo), .dout(new_new_n1337__));
  buf1  g0117(.din(n2340_lo), .dout(new_new_n1339__));
  not1  g0118(.din(n2340_lo), .dout(new_new_n1340__));
  buf1  g0119(.din(n3241_o2), .dout(new_new_n1341__));
  not1  g0120(.din(n3241_o2), .dout(new_new_n1342__));
  buf1  g0121(.din(n3242_o2), .dout(new_new_n1343__));
  not1  g0122(.din(n3242_o2), .dout(new_new_n1344__));
  not1  g0123(.din(n3610_o2), .dout(new_new_n1346__));
  not1  g0124(.din(n3980_o2), .dout(new_new_n1348__));
  not1  g0125(.din(n3968_o2), .dout(new_new_n1350__));
  buf1  g0126(.din(n4298_o2), .dout(new_new_n1351__));
  buf1  g0127(.din(n4371_o2), .dout(new_new_n1353__));
  not1  g0128(.din(n4413_o2), .dout(new_new_n1356__));
  buf1  g0129(.din(n4418_o2), .dout(new_new_n1357__));
  buf1  g0130(.din(n4628_o2), .dout(new_new_n1359__));
  not1  g0131(.din(n4629_o2), .dout(new_new_n1362__));
  buf1  g0132(.din(n4633_o2), .dout(new_new_n1363__));
  not1  g0133(.din(n4633_o2), .dout(new_new_n1364__));
  buf1  g0134(.din(n4634_o2), .dout(new_new_n1365__));
  not1  g0135(.din(n4634_o2), .dout(new_new_n1366__));
  buf1  g0136(.din(n4732_o2), .dout(new_new_n1367__));
  not1  g0137(.din(n4732_o2), .dout(new_new_n1368__));
  buf1  g0138(.din(n4733_o2), .dout(new_new_n1369__));
  not1  g0139(.din(n4733_o2), .dout(new_new_n1370__));
  not1  g0140(.din(n4884_o2), .dout(new_new_n1372__));
  not1  g0141(.din(n4886_o2), .dout(new_new_n1374__));
  buf1  g0142(.din(n4890_o2), .dout(new_new_n1375__));
  buf1  g0143(.din(n5011_o2), .dout(new_new_n1377__));
  not1  g0144(.din(n5011_o2), .dout(new_new_n1378__));
  buf1  g0145(.din(n5012_o2), .dout(new_new_n1379__));
  not1  g0146(.din(n5012_o2), .dout(new_new_n1380__));
  buf1  g0147(.din(n5013_o2), .dout(new_new_n1381__));
  not1  g0148(.din(n5013_o2), .dout(new_new_n1382__));
  buf1  g0149(.din(n5014_o2), .dout(new_new_n1383__));
  buf1  g0150(.din(n5015_o2), .dout(new_new_n1385__));
  not1  g0151(.din(n5015_o2), .dout(new_new_n1386__));
  buf1  g0152(.din(n5021_o2), .dout(new_new_n1387__));
  buf1  g0153(.din(n5016_o2), .dout(new_new_n1389__));
  not1  g0154(.din(n5026_o2), .dout(new_new_n1392__));
  buf1  g0155(.din(n4377_o2), .dout(new_new_n1393__));
  buf1  g0156(.din(n4378_o2), .dout(new_new_n1395__));
  buf1  g0157(.din(n4389_o2), .dout(new_new_n1397__));
  not1  g0158(.din(n4389_o2), .dout(new_new_n1398__));
  buf1  g0159(.din(n327_inv), .dout(new_new_n1399__));
  buf1  g0160(.din(n330_inv), .dout(new_new_n1401__));
  buf1  g0161(.din(n4398_o2), .dout(new_new_n1403__));
  not1  g0162(.din(n4398_o2), .dout(new_new_n1404__));
  buf1  g0163(.din(n4401_o2), .dout(new_new_n1405__));
  not1  g0164(.din(n4401_o2), .dout(new_new_n1406__));
  buf1  g0165(.din(n5117_o2), .dout(new_new_n1407__));
  buf1  g0166(.din(n5115_o2), .dout(new_new_n1409__));
  buf1  g0167(.din(n5122_o2), .dout(new_new_n1411__));
  buf1  g0168(.din(n5121_o2), .dout(new_new_n1413__));
  buf1  g0169(.din(n5119_o2), .dout(new_new_n1415__));
  buf1  g0170(.din(n5116_o2), .dout(new_new_n1417__));
  buf1  g0171(.din(n5123_o2), .dout(new_new_n1419__));
  not1  g0172(.din(n5123_o2), .dout(new_new_n1420__));
  buf1  g0173(.din(n5156_o2), .dout(new_new_n1421__));
  not1  g0174(.din(n5156_o2), .dout(new_new_n1422__));
  buf1  g0175(.din(n5167_o2), .dout(new_new_n1423__));
  not1  g0176(.din(n5167_o2), .dout(new_new_n1424__));
  buf1  g0177(.din(n4454_o2), .dout(new_new_n1425__));
  buf1  g0178(.din(n4455_o2), .dout(new_new_n1427__));
  buf1  g0179(.din(n4456_o2), .dout(new_new_n1429__));
  buf1  g0180(.din(n4505_o2), .dout(new_new_n1431__));
  buf1  g0181(.din(G742_o2), .dout(new_new_n1433__));
  not1  g0182(.din(G742_o2), .dout(new_new_n1434__));
  not1  g0183(.din(G727_o2), .dout(new_new_n1436__));
  buf1  g0184(.din(n4567_o2), .dout(new_new_n1437__));
  buf1  g0185(.din(n4568_o2), .dout(new_new_n1439__));
  buf1  g0186(.din(n4569_o2), .dout(new_new_n1441__));
  buf1  g0187(.din(n4571_o2), .dout(new_new_n1443__));
  not1  g0188(.din(n4571_o2), .dout(new_new_n1444__));
  buf1  g0189(.din(n4572_o2), .dout(new_new_n1445__));
  not1  g0190(.din(n4572_o2), .dout(new_new_n1446__));
  buf1  g0191(.din(n399_inv), .dout(new_new_n1447__));
  buf1  g0192(.din(n4539_o2), .dout(new_new_n1449__));
  not1  g0193(.din(n4539_o2), .dout(new_new_n1450__));
  buf1  g0194(.din(n4651_o2), .dout(new_new_n1451__));
  not1  g0195(.din(n4651_o2), .dout(new_new_n1452__));
  buf1  g0196(.din(n4652_o2), .dout(new_new_n1453__));
  buf1  g0197(.din(n4653_o2), .dout(new_new_n1455__));
  not1  g0198(.din(n4653_o2), .dout(new_new_n1456__));
  buf1  g0199(.din(G1514_o2), .dout(new_new_n1457__));
  not1  g0200(.din(G1514_o2), .dout(new_new_n1458__));
  buf1  g0201(.din(G1823_o2), .dout(new_new_n1459__));
  not1  g0202(.din(G1823_o2), .dout(new_new_n1460__));
  buf1  g0203(.din(n4783_o2), .dout(new_new_n1461__));
  not1  g0204(.din(n4783_o2), .dout(new_new_n1462__));
  buf1  g0205(.din(n4787_o2), .dout(new_new_n1463__));
  buf1  g0206(.din(n426_inv), .dout(new_new_n1465__));
  buf1  g0207(.din(n429_inv), .dout(new_new_n1467__));
  not1  g0208(.din(n429_inv), .dout(new_new_n1468__));
  buf1  g0209(.din(n4816_o2), .dout(new_new_n1469__));
  not1  g0210(.din(n4816_o2), .dout(new_new_n1470__));
  buf1  g0211(.din(n435_inv), .dout(new_new_n1471__));
  buf1  g0212(.din(G572_o2), .dout(new_new_n1473__));
  not1  g0213(.din(G572_o2), .dout(new_new_n1474__));
  buf1  g0214(.din(n4919_o2), .dout(new_new_n1475__));
  not1  g0215(.din(n4919_o2), .dout(new_new_n1476__));
  buf1  g0216(.din(n4920_o2), .dout(new_new_n1477__));
  buf1  g0217(.din(n4921_o2), .dout(new_new_n1479__));
  buf1  g0218(.din(G1048_o2), .dout(new_new_n1481__));
  not1  g0219(.din(G1048_o2), .dout(new_new_n1482__));
  buf1  g0220(.din(n5041_o2), .dout(new_new_n1483__));
  not1  g0221(.din(n5041_o2), .dout(new_new_n1484__));
  buf1  g0222(.din(n5094_o2), .dout(new_new_n1485__));
  not1  g0223(.din(n5094_o2), .dout(new_new_n1486__));
  buf1  g0224(.din(n5278_o2), .dout(new_new_n1487__));
  not1  g0225(.din(n5278_o2), .dout(new_new_n1488__));
  buf1  g0226(.din(n5301_o2), .dout(new_new_n1489__));
  not1  g0227(.din(n5301_o2), .dout(new_new_n1490__));
  buf1  g0228(.din(G2610_o2), .dout(new_new_n1491__));
  buf1  g0229(.din(G3174_o2), .dout(new_new_n1493__));
  buf1  g0230(.din(G3146_o2), .dout(new_new_n1495__));
  buf1  g0231(.din(G3217_o2), .dout(new_new_n1497__));
  buf1  g0232(.din(G3220_o2), .dout(new_new_n1499__));
  buf1  g0233(.din(G2839_o2), .dout(new_new_n1501__));
  buf1  g0234(.din(G3251_o2), .dout(new_new_n1503__));
  buf1  g0235(.din(G3042_o2), .dout(new_new_n1505__));
  not1  g0236(.din(G3045_o2), .dout(new_new_n1508__));
  buf1  g0237(.din(G3262_o2), .dout(new_new_n1509__));
  buf1  g0238(.din(G2845_o2), .dout(new_new_n1511__));
  buf1  g0239(.din(G2929_o2), .dout(new_new_n1513__));
  buf1  g0240(.din(G2848_o2), .dout(new_new_n1515__));
  buf1  g0241(.din(G2851_o2), .dout(new_new_n1517__));
  buf1  g0242(.din(G3291_o2), .dout(new_new_n1519__));
  buf1  g0243(.din(G3254_o2), .dout(new_new_n1521__));
  buf1  g0244(.din(G2666_o2), .dout(new_new_n1523__));
  not1  g0245(.din(G2666_o2), .dout(new_new_n1524__));
  buf1  g0246(.din(n5099_o2), .dout(new_new_n1525__));
  buf1  g0247(.din(n5100_o2), .dout(new_new_n1527__));
  not1  g0248(.din(n5100_o2), .dout(new_new_n1528__));
  buf1  g0249(.din(n5101_o2), .dout(new_new_n1529__));
  not1  g0250(.din(n5101_o2), .dout(new_new_n1530__));
  buf1  g0251(.din(G2558_o2), .dout(new_new_n1531__));
  buf1  g0252(.din(n5266_o2), .dout(new_new_n1533__));
  not1  g0253(.din(n5266_o2), .dout(new_new_n1534__));
  buf1  g0254(.din(n5267_o2), .dout(new_new_n1535__));
  not1  g0255(.din(n5267_o2), .dout(new_new_n1536__));
  buf1  g0256(.din(G2759_o2), .dout(new_new_n1537__));
  not1  g0257(.din(G2759_o2), .dout(new_new_n1538__));
  buf1  g0258(.din(n537_inv), .dout(new_new_n1539__));
  buf1  g0259(.din(n540_inv), .dout(new_new_n1541__));
  buf1  g0260(.din(n543_inv), .dout(new_new_n1543__));
  buf1  g0261(.din(n5292_o2), .dout(new_new_n1545__));
  buf1  g0262(.din(n5293_o2), .dout(new_new_n1547__));
  buf1  g0263(.din(n5294_o2), .dout(new_new_n1549__));
  not1  g0264(.din(n5294_o2), .dout(new_new_n1550__));
  buf1  g0265(.din(n5295_o2), .dout(new_new_n1551__));
  buf1  g0266(.din(G618_o2), .dout(new_new_n1553__));
  not1  g0267(.din(G618_o2), .dout(new_new_n1554__));
  buf1  g0268(.din(G621_o2), .dout(new_new_n1555__));
  not1  g0269(.din(G621_o2), .dout(new_new_n1556__));
  not1  g0270(.din(G384_o2), .dout(new_new_n1558__));
  not1  g0271(.din(G377_o2), .dout(new_new_n1560__));
  buf1  g0272(.din(n570_inv), .dout(new_new_n1561__));
  not1  g0273(.din(n570_inv), .dout(new_new_n1562__));
  buf1  g0274(.din(G3171_o2), .dout(new_new_n1563__));
  buf1  g0275(.din(G2552_o2), .dout(new_new_n1565__));
  buf1  g0276(.din(G3272_o2), .dout(new_new_n1567__));
  buf1  g0277(.din(G2015_o2), .dout(new_new_n1569__));
  not1  g0278(.din(G2015_o2), .dout(new_new_n1570__));
  buf1  g0279(.din(G3294_o2), .dout(new_new_n1571__));
  buf1  g0280(.din(G3281_o2), .dout(new_new_n1573__));
  buf1  g0281(.din(G3320_o2), .dout(new_new_n1575__));
  buf1  g0282(.din(G3275_o2), .dout(new_new_n1577__));
  buf1  g0283(.din(G3140_o2), .dout(new_new_n1579__));
  buf1  g0284(.din(G2836_o2), .dout(new_new_n1581__));
  buf1  g0285(.din(G2926_o2), .dout(new_new_n1583__));
  buf1  g0286(.din(G2842_o2), .dout(new_new_n1585__));
  buf1  g0287(.din(G3302_o2), .dout(new_new_n1587__));
  buf1  g0288(.din(G3288_o2), .dout(new_new_n1589__));
  buf1  g0289(.din(G3143_o2), .dout(new_new_n1591__));
  not1  g0290(.din(G3100_o2), .dout(new_new_n1594__));
  buf1  g0291(.din(G2512_o2), .dout(new_new_n1595__));
  not1  g0292(.din(G2512_o2), .dout(new_new_n1596__));
  buf1  g0293(.din(n5325_o2), .dout(new_new_n1597__));
  not1  g0294(.din(n5325_o2), .dout(new_new_n1598__));
  buf1  g0295(.din(n5326_o2), .dout(new_new_n1599__));
  not1  g0296(.din(n5326_o2), .dout(new_new_n1600__));
  buf1  g0297(.din(n5327_o2), .dout(new_new_n1601__));
  not1  g0298(.din(n5327_o2), .dout(new_new_n1602__));
  buf1  g0299(.din(n1857_lo_buf_o2), .dout(new_new_n1603__));
  not1  g0300(.din(n1857_lo_buf_o2), .dout(new_new_n1604__));
  buf1  g0301(.din(n2097_lo_buf_o2), .dout(new_new_n1605__));
  not1  g0302(.din(n2097_lo_buf_o2), .dout(new_new_n1606__));
  buf1  g0303(.din(G2669_o2), .dout(new_new_n1607__));
  not1  g0304(.din(G2669_o2), .dout(new_new_n1608__));
  buf1  g0305(.din(n642_inv), .dout(new_new_n1609__));
  buf1  g0306(.din(G568_o2), .dout(new_new_n1611__));
  buf1  g0307(.din(n648_inv), .dout(new_new_n1613__));
  buf1  g0308(.din(G565_o2), .dout(new_new_n1615__));
  buf1  g0309(.din(G559_o2), .dout(new_new_n1617__));
  buf1  g0310(.din(n1821_lo_buf_o2), .dout(new_new_n1619__));
  not1  g0311(.din(n1821_lo_buf_o2), .dout(new_new_n1620__));
  buf1  g0312(.din(n1905_lo_buf_o2), .dout(new_new_n1621__));
  not1  g0313(.din(n1905_lo_buf_o2), .dout(new_new_n1622__));
  buf1  g0314(.din(n2133_lo_buf_o2), .dout(new_new_n1623__));
  not1  g0315(.din(n2133_lo_buf_o2), .dout(new_new_n1624__));
  buf1  g0316(.din(n2145_lo_buf_o2), .dout(new_new_n1625__));
  not1  g0317(.din(n2145_lo_buf_o2), .dout(new_new_n1626__));
  buf1  g0318(.din(n2157_lo_buf_o2), .dout(new_new_n1627__));
  not1  g0319(.din(n2157_lo_buf_o2), .dout(new_new_n1628__));
  buf1  g0320(.din(n2205_lo_buf_o2), .dout(new_new_n1629__));
  buf1  g0321(.din(n2217_lo_buf_o2), .dout(new_new_n1631__));
  buf1  g0322(.din(G447_o2), .dout(new_new_n1633__));
  not1  g0323(.din(G447_o2), .dout(new_new_n1634__));
  buf1  g0324(.din(G434_o2), .dout(new_new_n1635__));
  not1  g0325(.din(G422_o2), .dout(new_new_n1638__));
  buf1  g0326(.din(G461_o2), .dout(new_new_n1639__));
  buf1  g0327(.din(G3312_o2), .dout(new_new_n1641__));
  buf1  g0328(.din(G3332_o2), .dout(new_new_n1643__));
  buf1  g0329(.din(G3195_o2), .dout(new_new_n1645__));
  buf1  g0330(.din(G2607_o2), .dout(new_new_n1647__));
  buf1  g0331(.din(n702_inv), .dout(new_new_n1649__));
  buf1  g0332(.din(G1005_o2), .dout(new_new_n1651__));
  buf1  g0333(.din(G1008_o2), .dout(new_new_n1653__));
  buf1  g0334(.din(n2001_lo_buf_o2), .dout(new_new_n1655__));
  buf1  g0335(.din(n2169_lo_buf_o2), .dout(new_new_n1657__));
  not1  g0336(.din(n2169_lo_buf_o2), .dout(new_new_n1658__));
  buf1  g0337(.din(n2229_lo_buf_o2), .dout(new_new_n1659__));
  buf1  g0338(.din(n2301_lo_buf_o2), .dout(new_new_n1661__));
  not1  g0339(.din(n2301_lo_buf_o2), .dout(new_new_n1662__));
  buf1  g0340(.din(n723_inv), .dout(new_new_n1663__));
  buf1  g0341(.din(G2947_o2), .dout(new_new_n1665__));
  buf1  g0342(.din(n2013_lo_buf_o2), .dout(new_new_n1667__));
  not1  g0343(.din(n2013_lo_buf_o2), .dout(new_new_n1668__));
  buf1  g0344(.din(n2025_lo_buf_o2), .dout(new_new_n1669__));
  not1  g0345(.din(n2025_lo_buf_o2), .dout(new_new_n1670__));
  buf1  g0346(.din(n2037_lo_buf_o2), .dout(new_new_n1671__));
  not1  g0347(.din(n2037_lo_buf_o2), .dout(new_new_n1672__));
  buf1  g0348(.din(n2049_lo_buf_o2), .dout(new_new_n1673__));
  not1  g0349(.din(n2049_lo_buf_o2), .dout(new_new_n1674__));
  buf1  g0350(.din(n2181_lo_buf_o2), .dout(new_new_n1675__));
  not1  g0351(.din(n2181_lo_buf_o2), .dout(new_new_n1676__));
  buf1  g0352(.din(n744_inv), .dout(new_new_n1677__));
  buf1  g0353(.din(n747_inv), .dout(new_new_n1679__));
  buf1  g0354(.din(n750_inv), .dout(new_new_n1681__));
  buf1  g0355(.din(n753_inv), .dout(new_new_n1683__));
  buf1  g0356(.din(G3350_o2), .dout(new_new_n1685__));
  not1  g0357(.din(G3350_o2), .dout(new_new_n1686__));
  buf1  g0358(.din(G3360_o2), .dout(new_new_n1687__));
  not1  g0359(.din(G3360_o2), .dout(new_new_n1688__));
  buf1  g0360(.din(G3373_o2), .dout(new_new_n1689__));
  not1  g0361(.din(G3373_o2), .dout(new_new_n1690__));
  buf1  g0362(.din(G3237_o2), .dout(new_new_n1691__));
  not1  g0363(.din(G3237_o2), .dout(new_new_n1692__));
  buf1  g0364(.din(G2773_o2), .dout(new_new_n1693__));
  not1  g0365(.din(G2773_o2), .dout(new_new_n1694__));
  buf1  g0366(.din(G1733_o2), .dout(new_new_n1695__));
  not1  g0367(.din(G1733_o2), .dout(new_new_n1696__));
  buf1  g0368(.din(G1738_o2), .dout(new_new_n1697__));
  not1  g0369(.din(G1738_o2), .dout(new_new_n1698__));
  buf1  g0370(.din(G1751_o2), .dout(new_new_n1699__));
  not1  g0371(.din(G1751_o2), .dout(new_new_n1700__));
  buf1  g0372(.din(G2216_o2), .dout(new_new_n1701__));
  not1  g0373(.din(G2216_o2), .dout(new_new_n1702__));
  buf1  g0374(.din(G2219_o2), .dout(new_new_n1703__));
  not1  g0375(.din(G2219_o2), .dout(new_new_n1704__));
  buf1  g0376(.din(n786_inv), .dout(new_new_n1705__));
  buf1  g0377(.din(n789_inv), .dout(new_new_n1707__));
  buf1  g0378(.din(G787_o2), .dout(new_new_n1709__));
  buf1  g0379(.din(G2823_o2), .dout(new_new_n1711__));
  buf1  g0380(.din(G2796_o2), .dout(new_new_n1713__));
  buf1  g0381(.din(G875_o2), .dout(new_new_n1715__));
  not1  g0382(.din(G875_o2), .dout(new_new_n1716__));
  buf1  g0383(.din(G2208_o2), .dout(new_new_n1717__));
  not1  g0384(.din(G2208_o2), .dout(new_new_n1718__));
  buf1  g0385(.din(G2211_o2), .dout(new_new_n1719__));
  not1  g0386(.din(G2211_o2), .dout(new_new_n1720__));
  buf1  g0387(.din(n1989_lo_buf_o2), .dout(new_new_n1721__));
  buf1  g0388(.din(n2061_lo_buf_o2), .dout(new_new_n1723__));
  not1  g0389(.din(n2061_lo_buf_o2), .dout(new_new_n1724__));
  buf1  g0390(.din(n2313_lo_buf_o2), .dout(new_new_n1725__));
  not1  g0391(.din(n2313_lo_buf_o2), .dout(new_new_n1726__));
  buf1  g0392(.din(G2232_o2), .dout(new_new_n1727__));
  not1  g0393(.din(G2232_o2), .dout(new_new_n1728__));
  buf1  g0394(.din(G1725_o2), .dout(new_new_n1729__));
  not1  g0395(.din(G1725_o2), .dout(new_new_n1730__));
  buf1  g0396(.din(G1764_o2), .dout(new_new_n1731__));
  not1  g0397(.din(G1764_o2), .dout(new_new_n1732__));
  buf1  g0398(.din(G2356_o2), .dout(new_new_n1733__));
  not1  g0399(.din(G2356_o2), .dout(new_new_n1734__));
  buf1  g0400(.din(G2359_o2), .dout(new_new_n1735__));
  not1  g0401(.din(G2359_o2), .dout(new_new_n1736__));
  buf1  g0402(.din(G1180_o2), .dout(new_new_n1737__));
  not1  g0403(.din(G1180_o2), .dout(new_new_n1738__));
  buf1  g0404(.din(G1756_o2), .dout(new_new_n1739__));
  not1  g0405(.din(G1756_o2), .dout(new_new_n1740__));
  not1  g0406(.din(G2441_o2), .dout(new_new_n1742__));
  buf1  g0407(.din(G2887_o2), .dout(new_new_n1743__));
  not1  g0408(.din(G2887_o2), .dout(new_new_n1744__));
  buf1  g0409(.din(G2991_o2), .dout(new_new_n1745__));
  not1  g0410(.din(G2991_o2), .dout(new_new_n1746__));
  buf1  g0411(.din(n849_inv), .dout(new_new_n1747__));
  not1  g0412(.din(n849_inv), .dout(new_new_n1748__));
  buf1  g0413(.din(n852_inv), .dout(new_new_n1749__));
  not1  g0414(.din(n852_inv), .dout(new_new_n1750__));
  buf1  g0415(.din(n855_inv), .dout(new_new_n1751__));
  not1  g0416(.din(n855_inv), .dout(new_new_n1752__));
  buf1  g0417(.din(n858_inv), .dout(new_new_n1753__));
  not1  g0418(.din(n858_inv), .dout(new_new_n1754__));
  buf1  g0419(.din(n861_inv), .dout(new_new_n1755__));
  not1  g0420(.din(n861_inv), .dout(new_new_n1756__));
  buf1  g0421(.din(G2805_o2), .dout(new_new_n1757__));
  buf1  g0422(.din(G2906_o2), .dout(new_new_n1759__));
  buf1  g0423(.din(G2833_o2), .dout(new_new_n1761__));
  buf1  g0424(.din(n873_inv), .dout(new_new_n1763__));
  buf1  g0425(.din(G3353_o2), .dout(new_new_n1765__));
  not1  g0426(.din(G3353_o2), .dout(new_new_n1766__));
  buf1  g0427(.din(G3367_o2), .dout(new_new_n1767__));
  not1  g0428(.din(G3367_o2), .dout(new_new_n1768__));
  buf1  g0429(.din(G3346_o2), .dout(new_new_n1769__));
  not1  g0430(.din(G3346_o2), .dout(new_new_n1770__));
  buf1  g0431(.din(G3340_o2), .dout(new_new_n1771__));
  not1  g0432(.din(G3340_o2), .dout(new_new_n1772__));
  buf1  g0433(.din(G3376_o2), .dout(new_new_n1773__));
  not1  g0434(.din(G3376_o2), .dout(new_new_n1774__));
  buf1  g0435(.din(G3359_o2), .dout(new_new_n1775__));
  not1  g0436(.din(G3359_o2), .dout(new_new_n1776__));
  buf1  g0437(.din(G3240_o2), .dout(new_new_n1777__));
  not1  g0438(.din(G3240_o2), .dout(new_new_n1778__));
  buf1  g0439(.din(G3344_o2), .dout(new_new_n1779__));
  not1  g0440(.din(G3344_o2), .dout(new_new_n1780__));
  buf1  g0441(.din(G2880_o2), .dout(new_new_n1781__));
  not1  g0442(.din(G2880_o2), .dout(new_new_n1782__));
  buf1  g0443(.din(G2939_o2), .dout(new_new_n1783__));
  not1  g0444(.din(G2939_o2), .dout(new_new_n1784__));
  buf1  g0445(.din(G2248_o2), .dout(new_new_n1785__));
  not1  g0446(.din(G2248_o2), .dout(new_new_n1786__));
  buf1  g0447(.din(G2251_o2), .dout(new_new_n1787__));
  not1  g0448(.din(G2251_o2), .dout(new_new_n1788__));
  buf1  g0449(.din(G2021_o2), .dout(new_new_n1789__));
  buf1  g0450(.din(G3383_o2), .dout(new_new_n1791__));
  not1  g0451(.din(G3383_o2), .dout(new_new_n1792__));
  buf1  g0452(.din(G3399_o2), .dout(new_new_n1793__));
  not1  g0453(.din(G3399_o2), .dout(new_new_n1794__));
  buf1  g0454(.din(G3404_o2), .dout(new_new_n1795__));
  not1  g0455(.din(G3404_o2), .dout(new_new_n1796__));
  buf1  g0456(.din(G3265_o2), .dout(new_new_n1797__));
  not1  g0457(.din(G3265_o2), .dout(new_new_n1798__));
  buf1  g0458(.din(G2866_o2), .dout(new_new_n1799__));
  not1  g0459(.din(G2866_o2), .dout(new_new_n1800__));
  buf1  g0460(.din(G2999_o2), .dout(new_new_n1801__));
  not1  g0461(.din(G2999_o2), .dout(new_new_n1802__));
  not1  g0462(.din(G736_o2), .dout(new_new_n1804__));
  buf1  g0463(.din(G739_o2), .dout(new_new_n1805__));
  buf1  g0464(.din(G1200_o2), .dout(new_new_n1807__));
  buf1  g0465(.din(G1203_o2), .dout(new_new_n1809__));
  buf1  g0466(.din(G3027_o2), .dout(new_new_n1811__));
  not1  g0467(.din(G3027_o2), .dout(new_new_n1812__));
  not1  g0468(.din(G1463_o2), .dout(new_new_n1814__));
  not1  g0469(.din(G1460_o2), .dout(new_new_n1816__));
  buf1  g0470(.din(G3012_o2), .dout(new_new_n1817__));
  not1  g0471(.din(G3012_o2), .dout(new_new_n1818__));
  buf1  g0472(.din(G1574_o2), .dout(new_new_n1819__));
  buf1  g0473(.din(G1646_o2), .dout(new_new_n1821__));
  buf1  g0474(.din(G1592_o2), .dout(new_new_n1823__));
  buf1  g0475(.din(G1664_o2), .dout(new_new_n1825__));
  not1  g0476(.din(G1547_o2), .dout(new_new_n1828__));
  not1  g0477(.din(G1619_o2), .dout(new_new_n1830__));
  buf1  g0478(.din(G1556_o2), .dout(new_new_n1831__));
  buf1  g0479(.din(G1628_o2), .dout(new_new_n1833__));
  not1  g0480(.din(G1583_o2), .dout(new_new_n1836__));
  not1  g0481(.din(G1655_o2), .dout(new_new_n1838__));
  buf1  g0482(.din(G1529_o2), .dout(new_new_n1839__));
  buf1  g0483(.din(G1601_o2), .dout(new_new_n1841__));
  buf1  g0484(.din(G1538_o2), .dout(new_new_n1843__));
  buf1  g0485(.din(G1610_o2), .dout(new_new_n1845__));
  buf1  g0486(.din(G1565_o2), .dout(new_new_n1847__));
  buf1  g0487(.din(G1637_o2), .dout(new_new_n1849__));
  buf1  g0488(.din(G2437_o2), .dout(new_new_n1851__));
  not1  g0489(.din(G2437_o2), .dout(new_new_n1852__));
  buf1  g0490(.din(n1008_inv), .dout(new_new_n1853__));
  buf1  g0491(.din(n1785_lo_buf_o2), .dout(new_new_n1855__));
  not1  g0492(.din(n1785_lo_buf_o2), .dout(new_new_n1856__));
  buf1  g0493(.din(n1845_lo_buf_o2), .dout(new_new_n1857__));
  not1  g0494(.din(n1845_lo_buf_o2), .dout(new_new_n1858__));
  buf1  g0495(.din(n1893_lo_buf_o2), .dout(new_new_n1859__));
  not1  g0496(.din(n1893_lo_buf_o2), .dout(new_new_n1860__));
  not1  g0497(.din(n1941_lo_buf_o2), .dout(new_new_n1862__));
  not1  g0498(.din(n1953_lo_buf_o2), .dout(new_new_n1864__));
  not1  g0499(.din(n1965_lo_buf_o2), .dout(new_new_n1866__));
  buf1  g0500(.din(n1977_lo_buf_o2), .dout(new_new_n1867__));
  not1  g0501(.din(n1977_lo_buf_o2), .dout(new_new_n1868__));
  buf1  g0502(.din(n2241_lo_buf_o2), .dout(new_new_n1869__));
  not1  g0503(.din(n2241_lo_buf_o2), .dout(new_new_n1870__));
  buf1  g0504(.din(n2253_lo_buf_o2), .dout(new_new_n1871__));
  not1  g0505(.din(n2253_lo_buf_o2), .dout(new_new_n1872__));
  buf1  g0506(.din(n2265_lo_buf_o2), .dout(new_new_n1873__));
  not1  g0507(.din(n2265_lo_buf_o2), .dout(new_new_n1874__));
  buf1  g0508(.din(n2277_lo_buf_o2), .dout(new_new_n1875__));
  not1  g0509(.din(n2277_lo_buf_o2), .dout(new_new_n1876__));
  buf1  g0510(.din(n2289_lo_buf_o2), .dout(new_new_n1877__));
  buf1  g0511(.din(G519_o2), .dout(new_new_n1879__));
  not1  g0512(.din(G519_o2), .dout(new_new_n1880__));
  buf1  g0513(.din(n1050_inv), .dout(new_new_n1881__));
  not1  g0514(.din(n1050_inv), .dout(new_new_n1882__));
  buf1  g0515(.din(n1053_inv), .dout(new_new_n1883__));
  not1  g0516(.din(n1053_inv), .dout(new_new_n1884__));
  buf1  g0517(.din(n1056_inv), .dout(new_new_n1885__));
  not1  g0518(.din(n1056_inv), .dout(new_new_n1886__));
  not1  g0519(.din(G1318_o2), .dout(new_new_n1888__));
  buf1  g0520(.din(n1062_inv), .dout(new_new_n1889__));
  not1  g0521(.din(n1062_inv), .dout(new_new_n1890__));
  buf1  g0522(.din(G593_o2), .dout(new_new_n1891__));
  not1  g0523(.din(G593_o2), .dout(new_new_n1892__));
  buf1  g0524(.din(n1068_inv), .dout(new_new_n1893__));
  not1  g0525(.din(n1068_inv), .dout(new_new_n1894__));
  buf1  g0526(.din(n1071_inv), .dout(new_new_n1895__));
  not1  g0527(.din(n1071_inv), .dout(new_new_n1896__));
  buf1  g0528(.din(n1074_inv), .dout(new_new_n1897__));
  not1  g0529(.din(n1074_inv), .dout(new_new_n1898__));
  buf1  g0530(.din(G2284_o2), .dout(new_new_n1899__));
  not1  g0531(.din(G2284_o2), .dout(new_new_n1900__));
  buf1  g0532(.din(G2580_o2), .dout(new_new_n1901__));
  not1  g0533(.din(G2580_o2), .dout(new_new_n1902__));
  buf1  g0534(.din(G2302_o2), .dout(new_new_n1903__));
  not1  g0535(.din(G2302_o2), .dout(new_new_n1904__));
  buf1  g0536(.din(G2598_o2), .dout(new_new_n1905__));
  not1  g0537(.din(G2598_o2), .dout(new_new_n1906__));
  buf1  g0538(.din(G2497_o2), .dout(new_new_n1907__));
  not1  g0539(.din(G2497_o2), .dout(new_new_n1908__));
  buf1  g0540(.din(G2651_o2), .dout(new_new_n1909__));
  not1  g0541(.din(G2651_o2), .dout(new_new_n1910__));
  buf1  g0542(.din(G2296_o2), .dout(new_new_n1911__));
  not1  g0543(.din(G2296_o2), .dout(new_new_n1912__));
  buf1  g0544(.din(G2308_o2), .dout(new_new_n1913__));
  not1  g0545(.din(G2308_o2), .dout(new_new_n1914__));
  buf1  g0546(.din(G2592_o2), .dout(new_new_n1915__));
  not1  g0547(.din(G2592_o2), .dout(new_new_n1916__));
  buf1  g0548(.din(G2604_o2), .dout(new_new_n1917__));
  not1  g0549(.din(G2604_o2), .dout(new_new_n1918__));
  buf1  g0550(.din(G2902_o2), .dout(new_new_n1919__));
  not1  g0551(.din(G2902_o2), .dout(new_new_n1920__));
  buf1  g0552(.din(G2975_o2), .dout(new_new_n1921__));
  not1  g0553(.din(G2975_o2), .dout(new_new_n1922__));
  buf1  g0554(.din(G2962_o2), .dout(new_new_n1923__));
  not1  g0555(.din(G2962_o2), .dout(new_new_n1924__));
  buf1  g0556(.din(G3069_o2), .dout(new_new_n1925__));
  not1  g0557(.din(G3069_o2), .dout(new_new_n1926__));
  buf1  g0558(.din(G2018_o2), .dout(new_new_n1927__));
  buf1  g0559(.din(G1176_o2), .dout(new_new_n1929__));
  not1  g0560(.din(G1176_o2), .dout(new_new_n1930__));
  buf1  g0561(.din(G1189_o2), .dout(new_new_n1931__));
  not1  g0562(.din(G1189_o2), .dout(new_new_n1932__));
  buf1  g0563(.din(G3066_o2), .dout(new_new_n1933__));
  not1  g0564(.din(G3066_o2), .dout(new_new_n1934__));
  buf1  g0565(.din(G3137_o2), .dout(new_new_n1935__));
  not1  g0566(.din(G3137_o2), .dout(new_new_n1936__));
  buf1  g0567(.din(G3038_o2), .dout(new_new_n1937__));
  not1  g0568(.din(G3038_o2), .dout(new_new_n1938__));
  buf1  g0569(.din(G3117_o2), .dout(new_new_n1939__));
  not1  g0570(.din(G3117_o2), .dout(new_new_n1940__));
  buf1  g0571(.din(G2384_o2), .dout(new_new_n1941__));
  not1  g0572(.din(G2384_o2), .dout(new_new_n1942__));
  buf1  g0573(.din(G2472_o2), .dout(new_new_n1943__));
  not1  g0574(.din(G2472_o2), .dout(new_new_n1944__));
  buf1  g0575(.din(G772_o2), .dout(new_new_n1945__));
  not1  g0576(.din(G772_o2), .dout(new_new_n1946__));
  buf1  g0577(.din(G935_o2), .dout(new_new_n1947__));
  buf1  g0578(.din(G2923_o2), .dout(new_new_n1949__));
  not1  g0579(.din(G2923_o2), .dout(new_new_n1950__));
  buf1  g0580(.din(G2971_o2), .dout(new_new_n1951__));
  not1  g0581(.din(G2971_o2), .dout(new_new_n1952__));
  buf1  g0582(.din(G2980_o2), .dout(new_new_n1953__));
  not1  g0583(.din(G2980_o2), .dout(new_new_n1954__));
  buf1  g0584(.din(G3039_o2), .dout(new_new_n1955__));
  not1  g0585(.din(G3039_o2), .dout(new_new_n1956__));
  buf1  g0586(.din(G2388_o2), .dout(new_new_n1957__));
  not1  g0587(.din(G2388_o2), .dout(new_new_n1958__));
  buf1  g0588(.din(G2287_o2), .dout(new_new_n1959__));
  not1  g0589(.din(G2287_o2), .dout(new_new_n1960__));
  buf1  g0590(.din(G3024_o2), .dout(new_new_n1961__));
  not1  g0591(.din(G3024_o2), .dout(new_new_n1962__));
  buf1  g0592(.din(G2916_o2), .dout(new_new_n1963__));
  not1  g0593(.din(G2916_o2), .dout(new_new_n1964__));
  buf1  g0594(.din(n1176_inv), .dout(new_new_n1965__));
  not1  g0595(.din(n1176_inv), .dout(new_new_n1966__));
  buf1  g0596(.din(G3035_o2), .dout(new_new_n1967__));
  not1  g0597(.din(G3035_o2), .dout(new_new_n1968__));
  buf1  g0598(.din(G3107_o2), .dout(new_new_n1969__));
  not1  g0599(.din(G3107_o2), .dout(new_new_n1970__));
  buf1  g0600(.din(G1023_o2), .dout(new_new_n1971__));
  not1  g0601(.din(G1024_o2), .dout(new_new_n1974__));
  not1  g0602(.din(G1311_o2), .dout(new_new_n1976__));
  not1  g0603(.din(G1312_o2), .dout(new_new_n1978__));
  buf1  g0604(.din(G3063_o2), .dout(new_new_n1979__));
  not1  g0605(.din(G3063_o2), .dout(new_new_n1980__));
  buf1  g0606(.din(G1520_o2), .dout(new_new_n1981__));
  buf1  g0607(.din(G1519_o2), .dout(new_new_n1983__));
  buf1  g0608(.din(G3078_o2), .dout(new_new_n1985__));
  not1  g0609(.din(G3078_o2), .dout(new_new_n1986__));
  buf1  g0610(.din(G2038_o2), .dout(new_new_n1987__));
  buf1  g0611(.din(G1848_o2), .dout(new_new_n1989__));
  buf1  g0612(.din(G1864_o2), .dout(new_new_n1991__));
  not1  g0613(.din(G1872_o2), .dout(new_new_n1994__));
  buf1  g0614(.din(G1880_o2), .dout(new_new_n1995__));
  not1  g0615(.din(G1888_o2), .dout(new_new_n1998__));
  buf1  g0616(.din(G1912_o2), .dout(new_new_n1999__));
  buf1  g0617(.din(G1928_o2), .dout(new_new_n2001__));
  not1  g0618(.din(G1936_o2), .dout(new_new_n2004__));
  buf1  g0619(.din(G1944_o2), .dout(new_new_n2005__));
  not1  g0620(.din(G1952_o2), .dout(new_new_n2008__));
  buf1  g0621(.din(G1850_o2), .dout(new_new_n2009__));
  buf1  g0622(.din(G1866_o2), .dout(new_new_n2011__));
  not1  g0623(.din(G1874_o2), .dout(new_new_n2014__));
  buf1  g0624(.din(G1882_o2), .dout(new_new_n2015__));
  not1  g0625(.din(G1890_o2), .dout(new_new_n2018__));
  buf1  g0626(.din(G1914_o2), .dout(new_new_n2019__));
  buf1  g0627(.din(G1930_o2), .dout(new_new_n2021__));
  not1  g0628(.din(G1938_o2), .dout(new_new_n2024__));
  buf1  g0629(.din(G1946_o2), .dout(new_new_n2025__));
  not1  g0630(.din(G1954_o2), .dout(new_new_n2028__));
  not1  g0631(.din(G1845_o2), .dout(new_new_n2030__));
  not1  g0632(.din(G1861_o2), .dout(new_new_n2032__));
  buf1  g0633(.din(G1869_o2), .dout(new_new_n2033__));
  not1  g0634(.din(G1877_o2), .dout(new_new_n2036__));
  buf1  g0635(.din(G1885_o2), .dout(new_new_n2037__));
  not1  g0636(.din(G1909_o2), .dout(new_new_n2040__));
  not1  g0637(.din(G1925_o2), .dout(new_new_n2042__));
  buf1  g0638(.din(G1933_o2), .dout(new_new_n2043__));
  not1  g0639(.din(G1941_o2), .dout(new_new_n2046__));
  buf1  g0640(.din(G1949_o2), .dout(new_new_n2047__));
  buf1  g0641(.din(G1846_o2), .dout(new_new_n2049__));
  buf1  g0642(.din(G1862_o2), .dout(new_new_n2051__));
  not1  g0643(.din(G1870_o2), .dout(new_new_n2054__));
  buf1  g0644(.din(G1878_o2), .dout(new_new_n2055__));
  not1  g0645(.din(G1886_o2), .dout(new_new_n2058__));
  buf1  g0646(.din(G1910_o2), .dout(new_new_n2059__));
  buf1  g0647(.din(G1926_o2), .dout(new_new_n2061__));
  not1  g0648(.din(G1934_o2), .dout(new_new_n2064__));
  buf1  g0649(.din(G1942_o2), .dout(new_new_n2065__));
  not1  g0650(.din(G1950_o2), .dout(new_new_n2068__));
  not1  g0651(.din(G1849_o2), .dout(new_new_n2070__));
  not1  g0652(.din(G1865_o2), .dout(new_new_n2072__));
  buf1  g0653(.din(G1873_o2), .dout(new_new_n2073__));
  not1  g0654(.din(G1881_o2), .dout(new_new_n2076__));
  buf1  g0655(.din(G1889_o2), .dout(new_new_n2077__));
  not1  g0656(.din(G1913_o2), .dout(new_new_n2080__));
  not1  g0657(.din(G1929_o2), .dout(new_new_n2082__));
  buf1  g0658(.din(G1937_o2), .dout(new_new_n2083__));
  not1  g0659(.din(G1945_o2), .dout(new_new_n2086__));
  buf1  g0660(.din(G1953_o2), .dout(new_new_n2087__));
  buf1  g0661(.din(G1843_o2), .dout(new_new_n2089__));
  buf1  g0662(.din(G1859_o2), .dout(new_new_n2091__));
  not1  g0663(.din(G1867_o2), .dout(new_new_n2094__));
  buf1  g0664(.din(G1875_o2), .dout(new_new_n2095__));
  not1  g0665(.din(G1883_o2), .dout(new_new_n2098__));
  buf1  g0666(.din(G1907_o2), .dout(new_new_n2099__));
  buf1  g0667(.din(G1923_o2), .dout(new_new_n2101__));
  not1  g0668(.din(G1931_o2), .dout(new_new_n2104__));
  buf1  g0669(.din(G1939_o2), .dout(new_new_n2105__));
  not1  g0670(.din(G1947_o2), .dout(new_new_n2108__));
  buf1  g0671(.din(G1844_o2), .dout(new_new_n2109__));
  buf1  g0672(.din(G1860_o2), .dout(new_new_n2111__));
  not1  g0673(.din(G1868_o2), .dout(new_new_n2114__));
  buf1  g0674(.din(G1876_o2), .dout(new_new_n2115__));
  not1  g0675(.din(G1884_o2), .dout(new_new_n2118__));
  buf1  g0676(.din(G1908_o2), .dout(new_new_n2119__));
  buf1  g0677(.din(G1924_o2), .dout(new_new_n2121__));
  not1  g0678(.din(G1932_o2), .dout(new_new_n2124__));
  buf1  g0679(.din(G1940_o2), .dout(new_new_n2125__));
  not1  g0680(.din(G1948_o2), .dout(new_new_n2128__));
  buf1  g0681(.din(G1847_o2), .dout(new_new_n2129__));
  buf1  g0682(.din(G1863_o2), .dout(new_new_n2131__));
  not1  g0683(.din(G1871_o2), .dout(new_new_n2134__));
  buf1  g0684(.din(G1879_o2), .dout(new_new_n2135__));
  not1  g0685(.din(G1887_o2), .dout(new_new_n2138__));
  buf1  g0686(.din(G1911_o2), .dout(new_new_n2139__));
  buf1  g0687(.din(G1927_o2), .dout(new_new_n2141__));
  not1  g0688(.din(G1935_o2), .dout(new_new_n2144__));
  buf1  g0689(.din(G1943_o2), .dout(new_new_n2145__));
  not1  g0690(.din(G1951_o2), .dout(new_new_n2148__));
  buf1  g0691(.din(G2444_o2), .dout(new_new_n2149__));
  not1  g0692(.din(G2444_o2), .dout(new_new_n2150__));
  buf1  g0693(.din(G2451_o2), .dout(new_new_n2151__));
  not1  g0694(.din(G2451_o2), .dout(new_new_n2152__));
  buf1  g0695(.din(G2502_o2), .dout(new_new_n2153__));
  not1  g0696(.din(G2502_o2), .dout(new_new_n2154__));
  buf1  g0697(.din(G2507_o2), .dout(new_new_n2155__));
  not1  g0698(.din(G2507_o2), .dout(new_new_n2156__));
  buf1  g0699(.din(n1464_inv), .dout(new_new_n2157__));
  buf1  g0700(.din(G2583_o2), .dout(new_new_n2159__));
  not1  g0701(.din(G2583_o2), .dout(new_new_n2160__));
  buf1  g0702(.din(n1797_lo_buf_o2), .dout(new_new_n2161__));
  not1  g0703(.din(n1797_lo_buf_o2), .dout(new_new_n2162__));
  buf1  g0704(.din(n1833_lo_buf_o2), .dout(new_new_n2163__));
  not1  g0705(.din(n1833_lo_buf_o2), .dout(new_new_n2164__));
  buf1  g0706(.din(n1881_lo_buf_o2), .dout(new_new_n2165__));
  not1  g0707(.din(n1881_lo_buf_o2), .dout(new_new_n2166__));
  buf1  g0708(.din(n1479_inv), .dout(new_new_n2167__));
  buf1  g0709(.din(n1482_inv), .dout(new_new_n2169__));
  buf1  g0710(.din(n1485_inv), .dout(new_new_n2171__));
  buf1  g0711(.din(G615_o2), .dout(new_new_n2173__));
  not1  g0712(.din(G615_o2), .dout(new_new_n2174__));
  buf1  g0713(.din(G2254_o2), .dout(new_new_n2175__));
  not1  g0714(.din(G2254_o2), .dout(new_new_n2176__));
  buf1  g0715(.din(G2255_o2), .dout(new_new_n2177__));
  not1  g0716(.din(G2255_o2), .dout(new_new_n2178__));
  buf1  g0717(.din(G2027_o2), .dout(new_new_n2179__));
  not1  g0718(.din(G2027_o2), .dout(new_new_n2180__));
  buf1  g0719(.din(G2393_o2), .dout(new_new_n2181__));
  not1  g0720(.din(G2393_o2), .dout(new_new_n2182__));
  buf1  g0721(.din(G527_o2), .dout(new_new_n2183__));
  not1  g0722(.din(G527_o2), .dout(new_new_n2184__));
  buf1  g0723(.din(G594_o2), .dout(new_new_n2185__));
  not1  g0724(.din(G594_o2), .dout(new_new_n2186__));
  buf1  g0725(.din(G1689_o2), .dout(new_new_n2187__));
  not1  g0726(.din(G1689_o2), .dout(new_new_n2188__));
  buf1  g0727(.din(G1693_o2), .dout(new_new_n2189__));
  not1  g0728(.din(G1693_o2), .dout(new_new_n2190__));
  buf1  g0729(.din(G2281_o2), .dout(new_new_n2191__));
  not1  g0730(.din(G2281_o2), .dout(new_new_n2192__));
  buf1  g0731(.din(G2014_o2), .dout(new_new_n2193__));
  not1  g0732(.din(G2014_o2), .dout(new_new_n2194__));
  buf1  g0733(.din(G2459_o2), .dout(new_new_n2195__));
  not1  g0734(.din(G2459_o2), .dout(new_new_n2196__));
  buf1  g0735(.din(G2561_o2), .dout(new_new_n2197__));
  not1  g0736(.din(G2561_o2), .dout(new_new_n2198__));
  buf1  g0737(.din(G2533_o2), .dout(new_new_n2199__));
  not1  g0738(.din(G2533_o2), .dout(new_new_n2200__));
  buf1  g0739(.din(n1749_lo_buf_o2), .dout(new_new_n2201__));
  not1  g0740(.din(n1749_lo_buf_o2), .dout(new_new_n2202__));
  buf1  g0741(.din(n1761_lo_buf_o2), .dout(new_new_n2203__));
  not1  g0742(.din(n1761_lo_buf_o2), .dout(new_new_n2204__));
  buf1  g0743(.din(n1773_lo_buf_o2), .dout(new_new_n2205__));
  not1  g0744(.din(n1773_lo_buf_o2), .dout(new_new_n2206__));
  buf1  g0745(.din(n1809_lo_buf_o2), .dout(new_new_n2207__));
  not1  g0746(.din(n1809_lo_buf_o2), .dout(new_new_n2208__));
  buf1  g0747(.din(G1955_o2), .dout(new_new_n2209__));
  not1  g0748(.din(G1955_o2), .dout(new_new_n2210__));
  buf1  g0749(.din(G1958_o2), .dout(new_new_n2211__));
  not1  g0750(.din(G1958_o2), .dout(new_new_n2212__));
  buf1  g0751(.din(G2562_o2), .dout(new_new_n2213__));
  not1  g0752(.din(G2562_o2), .dout(new_new_n2214__));
  buf1  g0753(.din(G2398_o2), .dout(new_new_n2215__));
  not1  g0754(.din(G2398_o2), .dout(new_new_n2216__));
  buf1  g0755(.din(n1554_inv), .dout(new_new_n2217__));
  not1  g0756(.din(n1554_inv), .dout(new_new_n2218__));
  buf1  g0757(.din(n1557_inv), .dout(new_new_n2219__));
  not1  g0758(.din(n1557_inv), .dout(new_new_n2220__));
  buf1  g0759(.din(G2577_o2), .dout(new_new_n2221__));
  not1  g0760(.din(G2577_o2), .dout(new_new_n2222__));
  buf1  g0761(.din(G2627_o2), .dout(new_new_n2223__));
  not1  g0762(.din(G2627_o2), .dout(new_new_n2224__));
  buf1  g0763(.din(G654_o2), .dout(new_new_n2225__));
  not1  g0764(.din(G654_o2), .dout(new_new_n2226__));
  buf1  g0765(.din(G660_o2), .dout(new_new_n2227__));
  not1  g0766(.din(G660_o2), .dout(new_new_n2228__));
  buf1  g0767(.din(G831_o2), .dout(new_new_n2229__));
  not1  g0768(.din(G831_o2), .dout(new_new_n2230__));
  buf1  g0769(.din(G919_o2), .dout(new_new_n2231__));
  not1  g0770(.din(G919_o2), .dout(new_new_n2232__));
  buf1  g0771(.din(G925_o2), .dout(new_new_n2233__));
  not1  g0772(.din(G925_o2), .dout(new_new_n2234__));
  buf1  g0773(.din(n1815_lo_buf_o2), .dout(new_new_n2235__));
  not1  g0774(.din(n1815_lo_buf_o2), .dout(new_new_n2236__));
  buf1  g0775(.din(n1899_lo_buf_o2), .dout(new_new_n2237__));
  not1  g0776(.din(n1899_lo_buf_o2), .dout(new_new_n2238__));
  buf1  g0777(.din(n2079_lo_buf_o2), .dout(new_new_n2239__));
  not1  g0778(.din(n2079_lo_buf_o2), .dout(new_new_n2240__));
  buf1  g0779(.din(n2127_lo_buf_o2), .dout(new_new_n2241__));
  not1  g0780(.din(n2127_lo_buf_o2), .dout(new_new_n2242__));
  buf1  g0781(.din(n2139_lo_buf_o2), .dout(new_new_n2243__));
  not1  g0782(.din(n2139_lo_buf_o2), .dout(new_new_n2244__));
  buf1  g0783(.din(n2151_lo_buf_o2), .dout(new_new_n2245__));
  not1  g0784(.din(n2151_lo_buf_o2), .dout(new_new_n2246__));
  buf1  g0785(.din(n2187_lo_buf_o2), .dout(new_new_n2247__));
  not1  g0786(.din(n2187_lo_buf_o2), .dout(new_new_n2248__));
  buf1  g0787(.din(n2199_lo_buf_o2), .dout(new_new_n2249__));
  not1  g0788(.din(n2199_lo_buf_o2), .dout(new_new_n2250__));
  buf1  g0789(.din(n2211_lo_buf_o2), .dout(new_new_n2251__));
  not1  g0790(.din(n2211_lo_buf_o2), .dout(new_new_n2252__));
  buf1  g0791(.din(G533_o2), .dout(new_new_n2253__));
  not1  g0792(.din(G533_o2), .dout(new_new_n2254__));
  buf1  g0793(.din(n1854_lo_buf_o2), .dout(new_new_n2255__));
  not1  g0794(.din(n1854_lo_buf_o2), .dout(new_new_n2256__));
  buf1  g0795(.din(n2094_lo_buf_o2), .dout(new_new_n2257__));
  not1  g0796(.din(n2094_lo_buf_o2), .dout(new_new_n2258__));
  buf1  g0797(.din(G667_o2), .dout(new_new_n2259__));
  not1  g0798(.din(G667_o2), .dout(new_new_n2260__));
  buf1  g0799(.din(G874_o2), .dout(new_new_n2261__));
  not1  g0800(.din(G874_o2), .dout(new_new_n2262__));
  buf1  g0801(.din(G851_o2), .dout(new_new_n2263__));
  not1  g0802(.din(G851_o2), .dout(new_new_n2264__));
  buf1  g0803(.din(G1127_o2), .dout(new_new_n2265__));
  not1  g0804(.din(G1127_o2), .dout(new_new_n2266__));
  buf1  g0805(.din(n1869_lo_buf_o2), .dout(new_new_n2267__));
  not1  g0806(.din(n1869_lo_buf_o2), .dout(new_new_n2268__));
  buf1  g0807(.din(n2109_lo_buf_o2), .dout(new_new_n2269__));
  not1  g0808(.din(n2109_lo_buf_o2), .dout(new_new_n2270__));
  buf1  g0809(.din(n2121_lo_buf_o2), .dout(new_new_n2271__));
  not1  g0810(.din(n2121_lo_buf_o2), .dout(new_new_n2272__));
  buf1  g0811(.din(G477_o2), .dout(new_new_n2273__));
  not1  g0812(.din(G477_o2), .dout(new_new_n2274__));
  buf1  g0813(.din(G491_o2), .dout(new_new_n2275__));
  not1  g0814(.din(G491_o2), .dout(new_new_n2276__));
  buf1  g0815(.din(G501_o2), .dout(new_new_n2277__));
  not1  g0816(.din(G501_o2), .dout(new_new_n2278__));
  buf1  g0817(.din(G786_o2), .dout(new_new_n2279__));
  not1  g0818(.din(G786_o2), .dout(new_new_n2280__));
  buf1  g0819(.din(G791_o2), .dout(new_new_n2281__));
  not1  g0820(.din(G791_o2), .dout(new_new_n2282__));
  buf1  g0821(.din(G1126_o2), .dout(new_new_n2283__));
  not1  g0822(.din(G1126_o2), .dout(new_new_n2284__));
  buf1  g0823(.din(G1052_o2), .dout(new_new_n2285__));
  not1  g0824(.din(G1052_o2), .dout(new_new_n2286__));
  buf1  g0825(.din(G1054_o2), .dout(new_new_n2287__));
  not1  g0826(.din(G1054_o2), .dout(new_new_n2288__));
  and1  g0827(.dina(new_new_n1350__), .dinb(new_new_n1348__), .dout(new_new_n2289__));
  and1  g0828(.dina(new_new_n2289__), .dinb(new_new_n1346__), .dout(new_new_n2290__));
  and1  g0829(.dina(new_new_n2290__), .dinb(new_new_n1356__), .dout(new_new_n2291__));
  or1   g0830(.dina(new_new_n1436__), .dinb(new_new_n1234__), .dout(new_new_n2292__));
  and1  g0831(.dina(new_new_n1433__), .dinb(new_new_n4363__), .dout(new_new_n2293__));
  or1   g0832(.dina(new_new_n1434__), .dinb(new_new_n4364__), .dout(new_new_n2294__));
  and1  g0833(.dina(new_new_n2293__), .dinb(new_new_n4365__), .dout(new_new_n2295__));
  or1   g0834(.dina(new_new_n2294__), .dinb(new_new_n4366__), .dout(new_new_n2296__));
  or1   g0835(.dina(new_new_n4367__), .dinb(new_new_n1422__), .dout(new_new_n2297__));
  and1  g0836(.dina(new_new_n4368__), .dinb(new_new_n4369__), .dout(new_new_n2298__));
  or1   g0837(.dina(new_new_n2298__), .dinb(new_new_n4370__), .dout(new_new_n2299__));
  and1  g0838(.dina(new_new_n1380__), .dinb(new_new_n4363__), .dout(new_new_n2300__));
  or1   g0839(.dina(new_new_n1379__), .dinb(new_new_n4364__), .dout(new_new_n2301__));
  and1  g0840(.dina(new_new_n4371__), .dinb(new_new_n4365__), .dout(new_new_n2302__));
  or1   g0841(.dina(new_new_n4372__), .dinb(new_new_n4366__), .dout(new_new_n2303__));
  or1   g0842(.dina(new_new_n2303__), .dinb(new_new_n2299__), .dout(new_new_n2304__));
  or1   g0843(.dina(new_new_n1383__), .dinb(new_new_n1284__), .dout(new_new_n2305__));
  or1   g0844(.dina(new_new_n1407__), .dinb(new_new_n1286__), .dout(new_new_n2306__));
  or1   g0845(.dina(new_new_n1409__), .dinb(new_new_n1288__), .dout(new_new_n2307__));
  or1   g0846(.dina(new_new_n1411__), .dinb(new_new_n1290__), .dout(new_new_n2308__));
  and1  g0847(.dina(new_new_n2306__), .dinb(new_new_n2305__), .dout(new_new_n2309__));
  and1  g0848(.dina(new_new_n2309__), .dinb(new_new_n2307__), .dout(new_new_n2310__));
  and1  g0849(.dina(new_new_n2310__), .dinb(new_new_n2308__), .dout(new_new_n2311__));
  or1   g0850(.dina(new_new_n1413__), .dinb(new_new_n4370__), .dout(new_new_n2312__));
  or1   g0851(.dina(new_new_n1415__), .dinb(new_new_n4369__), .dout(new_new_n2313__));
  or1   g0852(.dina(new_new_n1417__), .dinb(new_new_n4368__), .dout(new_new_n2314__));
  or1   g0853(.dina(new_new_n1419__), .dinb(new_new_n1302__), .dout(new_new_n2315__));
  and1  g0854(.dina(new_new_n2313__), .dinb(new_new_n2312__), .dout(new_new_n2316__));
  and1  g0855(.dina(new_new_n2316__), .dinb(new_new_n2314__), .dout(new_new_n2317__));
  and1  g0856(.dina(new_new_n2317__), .dinb(new_new_n2315__), .dout(new_new_n2318__));
  and1  g0857(.dina(new_new_n2318__), .dinb(new_new_n2311__), .dout(new_new_n2319__));
  or1   g0858(.dina(new_new_n2302__), .dinb(new_new_n4373__), .dout(new_new_n2320__));
  or1   g0859(.dina(new_new_n2320__), .dinb(new_new_n2319__), .dout(new_new_n2321__));
  and1  g0860(.dina(new_new_n2304__), .dinb(new_new_n2297__), .dout(new_new_n2322__));
  and1  g0861(.dina(new_new_n2322__), .dinb(new_new_n2321__), .dout(new_new_n2323__));
  and1  g0862(.dina(new_new_n4374__), .dinb(new_new_n4375__), .dout(new_new_n2324__));
  or1   g0863(.dina(new_new_n4376__), .dinb(new_new_n4377__), .dout(new_new_n2325__));
  and1  g0864(.dina(new_new_n4376__), .dinb(new_new_n4377__), .dout(new_new_n2326__));
  or1   g0865(.dina(new_new_n4374__), .dinb(new_new_n4375__), .dout(new_new_n2327__));
  and1  g0866(.dina(new_new_n2327__), .dinb(new_new_n2325__), .dout(new_new_n2328__));
  or1   g0867(.dina(new_new_n2326__), .dinb(new_new_n2324__), .dout(new_new_n2329__));
  or1   g0868(.dina(new_new_n2328__), .dinb(new_new_n1458__), .dout(new_new_n2330__));
  or1   g0869(.dina(new_new_n2329__), .dinb(new_new_n1457__), .dout(new_new_n2331__));
  and1  g0870(.dina(new_new_n2331__), .dinb(new_new_n2330__), .dout(new_new_n2332__));
  and1  g0871(.dina(new_new_n1459__), .dinb(new_new_n1424__), .dout(new_new_n2333__));
  and1  g0872(.dina(new_new_n1460__), .dinb(new_new_n1423__), .dout(new_new_n2334__));
  or1   g0873(.dina(new_new_n2334__), .dinb(new_new_n2333__), .dout(new_new_n2335__));
  and1  g0874(.dina(new_new_n4378__), .dinb(new_new_n1353__), .dout(new_new_n2336__));
  and1  g0875(.dina(new_new_n4378__), .dinb(new_new_n1351__), .dout(new_new_n2337__));
  or1   g0876(.dina(new_new_n2337__), .dinb(new_new_n1359__), .dout(new_new_n2338__));
  and1  g0877(.dina(new_new_n1375__), .dinb(new_new_n4379__), .dout(new_new_n2339__));
  and1  g0878(.dina(new_new_n2339__), .dinb(new_new_n1362__), .dout(new_new_n2340__));
  and1  g0879(.dina(new_new_n1482__), .dinb(new_new_n1421__), .dout(new_new_n2341__));
  or1   g0880(.dina(new_new_n1389__), .dinb(new_new_n1387__), .dout(new_new_n2342__));
  and1  g0881(.dina(new_new_n2342__), .dinb(new_new_n1474__), .dout(new_new_n2343__));
  and1  g0882(.dina(new_new_n1481__), .dinb(new_new_n1473__), .dout(new_new_n2344__));
  and1  g0883(.dina(new_new_n2344__), .dinb(new_new_n1392__), .dout(new_new_n2345__));
  or1   g0884(.dina(new_new_n2343__), .dinb(new_new_n2341__), .dout(new_new_n2346__));
  or1   g0885(.dina(new_new_n2346__), .dinb(new_new_n2345__), .dout(new_new_n2347__));
  or1   g0886(.dina(new_new_n1508__), .dinb(new_new_n1505__), .dout(new_new_n2348__));
  or1   g0887(.dina(new_new_n2348__), .dinb(new_new_n1517__), .dout(new_new_n2349__));
  and1  g0888(.dina(new_new_n4380__), .dinb(new_new_n1594__), .dout(new_new_n2350__));
  or1   g0889(.dina(new_new_n1591__), .dinb(new_new_n1579__), .dout(new_new_n2351__));
  or1   g0890(.dina(new_new_n2351__), .dinb(new_new_n1585__), .dout(new_new_n2352__));
  and1  g0891(.dina(new_new_n4381__), .dinb(new_new_n1645__), .dout(new_new_n2353__));
  and1  g0892(.dina(new_new_n1341__), .dinb(new_new_n1231__), .dout(new_new_n2354__));
  and1  g0893(.dina(new_new_n1342__), .dinb(new_new_n1232__), .dout(new_new_n2355__));
  or1   g0894(.dina(new_new_n2355__), .dinb(new_new_n2354__), .dout(new_new_n2356__));
  and1  g0895(.dina(new_new_n2356__), .dinb(new_new_n1374__), .dout(new_new_n2357__));
  and1  g0896(.dina(new_new_n2357__), .dinb(new_new_n1386__), .dout(new_new_n2358__));
  and1  g0897(.dina(new_new_n1385__), .dinb(new_new_n1372__), .dout(new_new_n2359__));
  or1   g0898(.dina(new_new_n2359__), .dinb(new_new_n2358__), .dout(new_new_n2360__));
  and1  g0899(.dina(new_new_n2360__), .dinb(new_new_n4371__), .dout(new_new_n2361__));
  and1  g0900(.dina(new_new_n1343__), .dinb(new_new_n1235__), .dout(new_new_n2362__));
  and1  g0901(.dina(new_new_n1344__), .dinb(new_new_n1236__), .dout(new_new_n2363__));
  or1   g0902(.dina(new_new_n2363__), .dinb(new_new_n2362__), .dout(new_new_n2364__));
  and1  g0903(.dina(new_new_n2364__), .dinb(new_new_n1420__), .dout(new_new_n2365__));
  and1  g0904(.dina(new_new_n2365__), .dinb(new_new_n4373__), .dout(new_new_n2366__));
  and1  g0905(.dina(new_new_n4382__), .dinb(new_new_n4383__), .dout(new_new_n2367__));
  or1   g0906(.dina(new_new_n4384__), .dinb(new_new_n4385__), .dout(new_new_n2368__));
  and1  g0907(.dina(new_new_n4384__), .dinb(new_new_n4385__), .dout(new_new_n2369__));
  or1   g0908(.dina(new_new_n4382__), .dinb(new_new_n4383__), .dout(new_new_n2370__));
  and1  g0909(.dina(new_new_n2370__), .dinb(new_new_n2368__), .dout(new_new_n2371__));
  or1   g0910(.dina(new_new_n2369__), .dinb(new_new_n2367__), .dout(new_new_n2372__));
  and1  g0911(.dina(new_new_n2372__), .dinb(new_new_n4379__), .dout(new_new_n2373__));
  or1   g0912(.dina(new_new_n2371__), .dinb(new_new_n1330__), .dout(new_new_n2374__));
  and1  g0913(.dina(new_new_n4386__), .dinb(new_new_n4387__), .dout(new_new_n2375__));
  or1   g0914(.dina(new_new_n4388__), .dinb(new_new_n4389__), .dout(new_new_n2376__));
  and1  g0915(.dina(new_new_n4388__), .dinb(new_new_n4389__), .dout(new_new_n2377__));
  or1   g0916(.dina(new_new_n4386__), .dinb(new_new_n4387__), .dout(new_new_n2378__));
  and1  g0917(.dina(new_new_n2378__), .dinb(new_new_n2376__), .dout(new_new_n2379__));
  or1   g0918(.dina(new_new_n2377__), .dinb(new_new_n2375__), .dout(new_new_n2380__));
  and1  g0919(.dina(new_new_n2379__), .dinb(new_new_n2373__), .dout(new_new_n2381__));
  and1  g0920(.dina(new_new_n2380__), .dinb(new_new_n2374__), .dout(new_new_n2382__));
  or1   g0921(.dina(new_new_n2382__), .dinb(new_new_n2381__), .dout(new_new_n2383__));
  and1  g0922(.dina(new_new_n4372__), .dinb(new_new_n4367__), .dout(new_new_n2384__));
  and1  g0923(.dina(new_new_n2384__), .dinb(new_new_n2383__), .dout(new_new_n2385__));
  or1   g0924(.dina(new_new_n2366__), .dinb(new_new_n2361__), .dout(new_new_n2386__));
  or1   g0925(.dina(new_new_n2386__), .dinb(new_new_n2385__), .dout(new_new_n2387__));
  or1   g0926(.dina(new_new_n1503__), .dinb(new_new_n1499__), .dout(new_new_n2388__));
  or1   g0927(.dina(new_new_n2388__), .dinb(new_new_n1511__), .dout(new_new_n2389__));
  and1  g0928(.dina(new_new_n4390__), .dinb(new_new_n1577__), .dout(new_new_n2390__));
  or1   g0929(.dina(new_new_n1521__), .dinb(new_new_n1495__), .dout(new_new_n2391__));
  or1   g0930(.dina(new_new_n2391__), .dinb(new_new_n1515__), .dout(new_new_n2392__));
  and1  g0931(.dina(new_new_n4391__), .dinb(new_new_n1573__), .dout(new_new_n2393__));
  or1   g0932(.dina(new_new_n1509__), .dinb(new_new_n1493__), .dout(new_new_n2394__));
  or1   g0933(.dina(new_new_n2394__), .dinb(new_new_n1513__), .dout(new_new_n2395__));
  and1  g0934(.dina(new_new_n4392__), .dinb(new_new_n1571__), .dout(new_new_n2396__));
  or1   g0935(.dina(new_new_n1519__), .dinb(new_new_n1497__), .dout(new_new_n2397__));
  or1   g0936(.dina(new_new_n2397__), .dinb(new_new_n1501__), .dout(new_new_n2398__));
  and1  g0937(.dina(new_new_n4393__), .dinb(new_new_n1575__), .dout(new_new_n2399__));
  or1   g0938(.dina(new_new_n4391__), .dinb(new_new_n4380__), .dout(new_new_n2400__));
  or1   g0939(.dina(new_new_n2400__), .dinb(new_new_n4392__), .dout(new_new_n2401__));
  or1   g0940(.dina(new_new_n2401__), .dinb(new_new_n4390__), .dout(new_new_n2402__));
  or1   g0941(.dina(new_new_n1589__), .dinb(new_new_n1563__), .dout(new_new_n2403__));
  or1   g0942(.dina(new_new_n2403__), .dinb(new_new_n1583__), .dout(new_new_n2404__));
  or1   g0943(.dina(new_new_n1587__), .dinb(new_new_n1567__), .dout(new_new_n2405__));
  or1   g0944(.dina(new_new_n2405__), .dinb(new_new_n1581__), .dout(new_new_n2406__));
  or1   g0945(.dina(new_new_n4393__), .dinb(new_new_n4381__), .dout(new_new_n2407__));
  or1   g0946(.dina(new_new_n2407__), .dinb(new_new_n4394__), .dout(new_new_n2408__));
  or1   g0947(.dina(new_new_n2408__), .dinb(new_new_n4395__), .dout(new_new_n2409__));
  or1   g0948(.dina(new_new_n2409__), .dinb(new_new_n2402__), .dout(new_new_n2410__));
  and1  g0949(.dina(new_new_n1555__), .dinb(new_new_n1553__), .dout(new_new_n2411__));
  or1   g0950(.dina(new_new_n1556__), .dinb(new_new_n1554__), .dout(new_new_n2412__));
  or1   g0951(.dina(new_new_n4395__), .dinb(new_new_n4394__), .dout(new_new_n2413__));
  or1   g0952(.dina(new_new_n2413__), .dinb(new_new_n4396__), .dout(new_new_n2414__));
  and1  g0953(.dina(new_new_n2414__), .dinb(new_new_n4397__), .dout(new_new_n2415__));
  and1  g0954(.dina(new_new_n2415__), .dinb(new_new_n1279__), .dout(new_new_n2416__));
  and1  g0955(.dina(new_new_n1776__), .dinb(new_new_n1770__), .dout(new_new_n2417__));
  or1   g0956(.dina(new_new_n1775__), .dinb(new_new_n1769__), .dout(new_new_n2418__));
  and1  g0957(.dina(new_new_n1780__), .dinb(new_new_n1771__), .dout(new_new_n2419__));
  or1   g0958(.dina(new_new_n1779__), .dinb(new_new_n1772__), .dout(new_new_n2420__));
  and1  g0959(.dina(new_new_n4398__), .dinb(new_new_n4399__), .dout(new_new_n2421__));
  or1   g0960(.dina(new_new_n4400__), .dinb(new_new_n4401__), .dout(new_new_n2422__));
  and1  g0961(.dina(new_new_n4400__), .dinb(new_new_n4401__), .dout(new_new_n2423__));
  or1   g0962(.dina(new_new_n4398__), .dinb(new_new_n4399__), .dout(new_new_n2424__));
  and1  g0963(.dina(new_new_n2424__), .dinb(new_new_n2422__), .dout(new_new_n2425__));
  or1   g0964(.dina(new_new_n2423__), .dinb(new_new_n2421__), .dout(new_new_n2426__));
  and1  g0965(.dina(new_new_n1797__), .dinb(new_new_n1689__), .dout(new_new_n2427__));
  or1   g0966(.dina(new_new_n1798__), .dinb(new_new_n1690__), .dout(new_new_n2428__));
  and1  g0967(.dina(new_new_n1796__), .dinb(new_new_n1692__), .dout(new_new_n2429__));
  or1   g0968(.dina(new_new_n1795__), .dinb(new_new_n1691__), .dout(new_new_n2430__));
  and1  g0969(.dina(new_new_n2430__), .dinb(new_new_n2428__), .dout(new_new_n2431__));
  or1   g0970(.dina(new_new_n2429__), .dinb(new_new_n2427__), .dout(new_new_n2432__));
  and1  g0971(.dina(new_new_n4402__), .dinb(new_new_n4403__), .dout(new_new_n2433__));
  or1   g0972(.dina(new_new_n4404__), .dinb(new_new_n4405__), .dout(new_new_n2434__));
  and1  g0973(.dina(new_new_n4404__), .dinb(new_new_n4405__), .dout(new_new_n2435__));
  or1   g0974(.dina(new_new_n4402__), .dinb(new_new_n4403__), .dout(new_new_n2436__));
  and1  g0975(.dina(new_new_n2436__), .dinb(new_new_n2434__), .dout(new_new_n2437__));
  or1   g0976(.dina(new_new_n2435__), .dinb(new_new_n2433__), .dout(new_new_n2438__));
  and1  g0977(.dina(new_new_n4396__), .dinb(new_new_n1339__), .dout(new_new_n2439__));
  or1   g0978(.dina(new_new_n2411__), .dinb(new_new_n1340__), .dout(new_new_n2440__));
  and1  g0979(.dina(new_new_n4406__), .dinb(new_new_n4408__), .dout(new_new_n2441__));
  or1   g0980(.dina(new_new_n4410__), .dinb(new_new_n4412__), .dout(new_new_n2442__));
  and1  g0981(.dina(new_new_n2441__), .dinb(new_new_n4415__), .dout(new_new_n2443__));
  or1   g0982(.dina(new_new_n2442__), .dinb(new_new_n4418__), .dout(new_new_n2444__));
  and1  g0983(.dina(new_new_n4420__), .dinb(new_new_n4421__), .dout(new_new_n2445__));
  or1   g0984(.dina(new_new_n4422__), .dinb(new_new_n4423__), .dout(new_new_n2446__));
  and1  g0985(.dina(new_new_n4422__), .dinb(new_new_n4423__), .dout(new_new_n2447__));
  or1   g0986(.dina(new_new_n4420__), .dinb(new_new_n4421__), .dout(new_new_n2448__));
  and1  g0987(.dina(new_new_n2448__), .dinb(new_new_n2446__), .dout(new_new_n2449__));
  or1   g0988(.dina(new_new_n2447__), .dinb(new_new_n2445__), .dout(new_new_n2450__));
  and1  g0989(.dina(new_new_n4424__), .dinb(new_new_n4408__), .dout(new_new_n2451__));
  or1   g0990(.dina(new_new_n4425__), .dinb(new_new_n4412__), .dout(new_new_n2452__));
  and1  g0991(.dina(new_new_n2451__), .dinb(new_new_n4418__), .dout(new_new_n2453__));
  or1   g0992(.dina(new_new_n2452__), .dinb(new_new_n4415__), .dout(new_new_n2454__));
  and1  g0993(.dina(new_new_n4426__), .dinb(new_new_n4427__), .dout(new_new_n2455__));
  or1   g0994(.dina(new_new_n4428__), .dinb(new_new_n4429__), .dout(new_new_n2456__));
  and1  g0995(.dina(new_new_n4428__), .dinb(new_new_n4429__), .dout(new_new_n2457__));
  or1   g0996(.dina(new_new_n4426__), .dinb(new_new_n4427__), .dout(new_new_n2458__));
  and1  g0997(.dina(new_new_n2458__), .dinb(new_new_n2456__), .dout(new_new_n2459__));
  or1   g0998(.dina(new_new_n2457__), .dinb(new_new_n2455__), .dout(new_new_n2460__));
  and1  g0999(.dina(new_new_n4430__), .dinb(new_new_n4406__), .dout(new_new_n2461__));
  or1   g1000(.dina(new_new_n4431__), .dinb(new_new_n4410__), .dout(new_new_n2462__));
  and1  g1001(.dina(new_new_n2461__), .dinb(new_new_n4419__), .dout(new_new_n2463__));
  or1   g1002(.dina(new_new_n2462__), .dinb(new_new_n4416__), .dout(new_new_n2464__));
  and1  g1003(.dina(new_new_n4430__), .dinb(new_new_n4424__), .dout(new_new_n2465__));
  or1   g1004(.dina(new_new_n4431__), .dinb(new_new_n4425__), .dout(new_new_n2466__));
  and1  g1005(.dina(new_new_n2465__), .dinb(new_new_n4416__), .dout(new_new_n2467__));
  or1   g1006(.dina(new_new_n2466__), .dinb(new_new_n4419__), .dout(new_new_n2468__));
  and1  g1007(.dina(new_new_n2454__), .dinb(new_new_n2444__), .dout(new_new_n2469__));
  or1   g1008(.dina(new_new_n2453__), .dinb(new_new_n2443__), .dout(new_new_n2470__));
  and1  g1009(.dina(new_new_n2469__), .dinb(new_new_n2464__), .dout(new_new_n2471__));
  or1   g1010(.dina(new_new_n2470__), .dinb(new_new_n2463__), .dout(new_new_n2472__));
  and1  g1011(.dina(new_new_n2471__), .dinb(new_new_n2468__), .dout(new_new_n2473__));
  or1   g1012(.dina(new_new_n2472__), .dinb(new_new_n2467__), .dout(new_new_n2474__));
  and1  g1013(.dina(new_new_n2474__), .dinb(new_new_n4432__), .dout(new_new_n2475__));
  and1  g1014(.dina(new_new_n2473__), .dinb(new_new_n4433__), .dout(new_new_n2476__));
  or1   g1015(.dina(new_new_n2476__), .dinb(new_new_n2475__), .dout(new_new_n2477__));
  and1  g1016(.dina(new_new_n4434__), .dinb(new_new_n4435__), .dout(new_new_n2478__));
  or1   g1017(.dina(new_new_n4436__), .dinb(new_new_n4437__), .dout(new_new_n2479__));
  and1  g1018(.dina(new_new_n4436__), .dinb(new_new_n4437__), .dout(new_new_n2480__));
  or1   g1019(.dina(new_new_n4434__), .dinb(new_new_n4435__), .dout(new_new_n2481__));
  and1  g1020(.dina(new_new_n2481__), .dinb(new_new_n2479__), .dout(new_new_n2482__));
  or1   g1021(.dina(new_new_n2480__), .dinb(new_new_n2478__), .dout(new_new_n2483__));
  and1  g1022(.dina(new_new_n4438__), .dinb(new_new_n4409__), .dout(new_new_n2484__));
  or1   g1023(.dina(new_new_n4439__), .dinb(new_new_n4413__), .dout(new_new_n2485__));
  and1  g1024(.dina(new_new_n4439__), .dinb(new_new_n4413__), .dout(new_new_n2486__));
  or1   g1025(.dina(new_new_n4438__), .dinb(new_new_n4409__), .dout(new_new_n2487__));
  and1  g1026(.dina(new_new_n2487__), .dinb(new_new_n2485__), .dout(new_new_n2488__));
  or1   g1027(.dina(new_new_n2486__), .dinb(new_new_n2484__), .dout(new_new_n2489__));
  or1   g1028(.dina(new_new_n2489__), .dinb(new_new_n4433__), .dout(new_new_n2490__));
  or1   g1029(.dina(new_new_n2488__), .dinb(new_new_n4432__), .dout(new_new_n2491__));
  and1  g1030(.dina(new_new_n2491__), .dinb(new_new_n2490__), .dout(new_new_n2492__));
  or1   g1031(.dina(new_new_n4440__), .dinb(new_new_n1633__), .dout(new_new_n2493__));
  and1  g1032(.dina(new_new_n1976__), .dinb(new_new_n1809__), .dout(new_new_n2494__));
  and1  g1033(.dina(new_new_n1978__), .dinb(new_new_n1807__), .dout(new_new_n2495__));
  or1   g1034(.dina(new_new_n2495__), .dinb(new_new_n2494__), .dout(new_new_n2496__));
  or1   g1035(.dina(new_new_n1983__), .dinb(new_new_n1814__), .dout(new_new_n2497__));
  or1   g1036(.dina(new_new_n1981__), .dinb(new_new_n1816__), .dout(new_new_n2498__));
  and1  g1037(.dina(new_new_n2498__), .dinb(new_new_n2497__), .dout(new_new_n2499__));
  and1  g1038(.dina(new_new_n4442__), .dinb(new_new_n4443__), .dout(new_new_n2500__));
  or1   g1039(.dina(new_new_n4445__), .dinb(new_new_n4448__), .dout(new_new_n2501__));
  and1  g1040(.dina(new_new_n2500__), .dinb(new_new_n1752__), .dout(new_new_n2502__));
  or1   g1041(.dina(new_new_n2501__), .dinb(new_new_n4449__), .dout(new_new_n2503__));
  and1  g1042(.dina(new_new_n2502__), .dinb(new_new_n4451__), .dout(new_new_n2504__));
  or1   g1043(.dina(new_new_n2503__), .dinb(new_new_n4453__), .dout(new_new_n2505__));
  and1  g1044(.dina(new_new_n2200__), .dinb(new_new_n2196__), .dout(new_new_n2506__));
  or1   g1045(.dina(new_new_n2199__), .dinb(new_new_n2195__), .dout(new_new_n2507__));
  and1  g1046(.dina(new_new_n2506__), .dinb(new_new_n2198__), .dout(new_new_n2508__));
  or1   g1047(.dina(new_new_n2507__), .dinb(new_new_n2197__), .dout(new_new_n2509__));
  and1  g1048(.dina(new_new_n2508__), .dinb(new_new_n2214__), .dout(new_new_n2510__));
  or1   g1049(.dina(new_new_n2509__), .dinb(new_new_n2213__), .dout(new_new_n2511__));
  and1  g1050(.dina(new_new_n1980__), .dinb(new_new_n1783__), .dout(new_new_n2512__));
  or1   g1051(.dina(new_new_n1979__), .dinb(new_new_n1784__), .dout(new_new_n2513__));
  and1  g1052(.dina(new_new_n1954__), .dinb(new_new_n1811__), .dout(new_new_n2514__));
  or1   g1053(.dina(new_new_n1953__), .dinb(new_new_n1812__), .dout(new_new_n2515__));
  and1  g1054(.dina(new_new_n2515__), .dinb(new_new_n2513__), .dout(new_new_n2516__));
  or1   g1055(.dina(new_new_n2514__), .dinb(new_new_n2512__), .dout(new_new_n2517__));
  and1  g1056(.dina(new_new_n4454__), .dinb(new_new_n4455__), .dout(new_new_n2518__));
  or1   g1057(.dina(new_new_n4456__), .dinb(new_new_n4458__), .dout(new_new_n2519__));
  and1  g1058(.dina(new_new_n2518__), .dinb(new_new_n1405__), .dout(new_new_n2520__));
  or1   g1059(.dina(new_new_n2519__), .dinb(new_new_n1406__), .dout(new_new_n2521__));
  and1  g1060(.dina(new_new_n2521__), .dinb(new_new_n1404__), .dout(new_new_n2522__));
  or1   g1061(.dina(new_new_n2520__), .dinb(new_new_n4459__), .dout(new_new_n2523__));
  and1  g1062(.dina(new_new_n4461__), .dinb(new_new_n4462__), .dout(new_new_n2524__));
  and1  g1063(.dina(new_new_n1968__), .dinb(new_new_n1800__), .dout(new_new_n2525__));
  or1   g1064(.dina(new_new_n1967__), .dinb(new_new_n1799__), .dout(new_new_n2526__));
  and1  g1065(.dina(new_new_n1963__), .dinb(new_new_n1801__), .dout(new_new_n2527__));
  or1   g1066(.dina(new_new_n1964__), .dinb(new_new_n1802__), .dout(new_new_n2528__));
  and1  g1067(.dina(new_new_n2528__), .dinb(new_new_n2526__), .dout(new_new_n2529__));
  or1   g1068(.dina(new_new_n2527__), .dinb(new_new_n2525__), .dout(new_new_n2530__));
  or1   g1069(.dina(new_new_n4464__), .dinb(new_new_n4467__), .dout(new_new_n2531__));
  and1  g1070(.dina(new_new_n4471__), .dinb(new_new_n4472__), .dout(new_new_n2532__));
  or1   g1071(.dina(new_new_n4473__), .dinb(new_new_n4474__), .dout(new_new_n2533__));
  and1  g1072(.dina(new_new_n4473__), .dinb(new_new_n4474__), .dout(new_new_n2534__));
  or1   g1073(.dina(new_new_n4471__), .dinb(new_new_n4472__), .dout(new_new_n2535__));
  and1  g1074(.dina(new_new_n2535__), .dinb(new_new_n2533__), .dout(new_new_n2536__));
  or1   g1075(.dina(new_new_n2534__), .dinb(new_new_n2532__), .dout(new_new_n2537__));
  or1   g1076(.dina(new_new_n4476__), .dinb(new_new_n4467__), .dout(new_new_n2538__));
  or1   g1077(.dina(new_new_n1818__), .dinb(new_new_n1781__), .dout(new_new_n2539__));
  or1   g1078(.dina(new_new_n1817__), .dinb(new_new_n1782__), .dout(new_new_n2540__));
  and1  g1079(.dina(new_new_n2540__), .dinb(new_new_n2539__), .dout(new_new_n2541__));
  or1   g1080(.dina(new_new_n4477__), .dinb(new_new_n4468__), .dout(new_new_n2542__));
  or1   g1081(.dina(new_new_n2089__), .dinb(new_new_n4479__), .dout(new_new_n2543__));
  or1   g1082(.dina(new_new_n2109__), .dinb(new_new_n4482__), .dout(new_new_n2544__));
  or1   g1083(.dina(new_new_n2030__), .dinb(new_new_n4487__), .dout(new_new_n2545__));
  or1   g1084(.dina(new_new_n2049__), .dinb(new_new_n4492__), .dout(new_new_n2546__));
  or1   g1085(.dina(new_new_n2129__), .dinb(new_new_n4497__), .dout(new_new_n2547__));
  or1   g1086(.dina(new_new_n1989__), .dinb(new_new_n4502__), .dout(new_new_n2548__));
  or1   g1087(.dina(new_new_n2070__), .dinb(new_new_n4506__), .dout(new_new_n2549__));
  or1   g1088(.dina(new_new_n2009__), .dinb(new_new_n4509__), .dout(new_new_n2550__));
  and1  g1089(.dina(new_new_n2544__), .dinb(new_new_n2543__), .dout(new_new_n2551__));
  and1  g1090(.dina(new_new_n2551__), .dinb(new_new_n2545__), .dout(new_new_n2552__));
  and1  g1091(.dina(new_new_n2552__), .dinb(new_new_n2546__), .dout(new_new_n2553__));
  and1  g1092(.dina(new_new_n2553__), .dinb(new_new_n2547__), .dout(new_new_n2554__));
  and1  g1093(.dina(new_new_n2554__), .dinb(new_new_n2548__), .dout(new_new_n2555__));
  and1  g1094(.dina(new_new_n2555__), .dinb(new_new_n2549__), .dout(new_new_n2556__));
  and1  g1095(.dina(new_new_n2556__), .dinb(new_new_n2550__), .dout(new_new_n2557__));
  and1  g1096(.dina(new_new_n2557__), .dinb(new_new_n4514__), .dout(new_new_n2558__));
  or1   g1097(.dina(new_new_n2099__), .dinb(new_new_n4520__), .dout(new_new_n2559__));
  or1   g1098(.dina(new_new_n2119__), .dinb(new_new_n4524__), .dout(new_new_n2560__));
  or1   g1099(.dina(new_new_n2040__), .dinb(new_new_n4529__), .dout(new_new_n2561__));
  or1   g1100(.dina(new_new_n2059__), .dinb(new_new_n4534__), .dout(new_new_n2562__));
  or1   g1101(.dina(new_new_n2139__), .dinb(new_new_n4540__), .dout(new_new_n2563__));
  or1   g1102(.dina(new_new_n1999__), .dinb(new_new_n4545__), .dout(new_new_n2564__));
  or1   g1103(.dina(new_new_n2080__), .dinb(new_new_n4551__), .dout(new_new_n2565__));
  or1   g1104(.dina(new_new_n2019__), .dinb(new_new_n4556__), .dout(new_new_n2566__));
  and1  g1105(.dina(new_new_n2560__), .dinb(new_new_n2559__), .dout(new_new_n2567__));
  and1  g1106(.dina(new_new_n2567__), .dinb(new_new_n2561__), .dout(new_new_n2568__));
  and1  g1107(.dina(new_new_n2568__), .dinb(new_new_n2562__), .dout(new_new_n2569__));
  and1  g1108(.dina(new_new_n2569__), .dinb(new_new_n2563__), .dout(new_new_n2570__));
  and1  g1109(.dina(new_new_n2570__), .dinb(new_new_n2564__), .dout(new_new_n2571__));
  and1  g1110(.dina(new_new_n2571__), .dinb(new_new_n2565__), .dout(new_new_n2572__));
  and1  g1111(.dina(new_new_n2572__), .dinb(new_new_n2566__), .dout(new_new_n2573__));
  and1  g1112(.dina(new_new_n2573__), .dinb(new_new_n4561__), .dout(new_new_n2574__));
  or1   g1113(.dina(new_new_n2574__), .dinb(new_new_n2558__), .dout(new_new_n2575__));
  and1  g1114(.dina(new_new_n1891__), .dinb(new_new_n1462__), .dout(new_new_n2576__));
  or1   g1115(.dina(new_new_n1892__), .dinb(new_new_n1461__), .dout(new_new_n2577__));
  and1  g1116(.dina(new_new_n4443__), .dinb(new_new_n4458__), .dout(new_new_n2578__));
  or1   g1117(.dina(new_new_n4448__), .dinb(new_new_n4455__), .dout(new_new_n2579__));
  and1  g1118(.dina(new_new_n2578__), .dinb(new_new_n2577__), .dout(new_new_n2580__));
  or1   g1119(.dina(new_new_n2579__), .dinb(new_new_n2576__), .dout(new_new_n2581__));
  and1  g1120(.dina(new_new_n4568__), .dinb(new_new_n2575__), .dout(new_new_n2582__));
  or1   g1121(.dina(new_new_n1901__), .dinb(new_new_n1899__), .dout(new_new_n2583__));
  or1   g1122(.dina(new_new_n1902__), .dinb(new_new_n1900__), .dout(new_new_n2584__));
  and1  g1123(.dina(new_new_n2584__), .dinb(new_new_n2583__), .dout(new_new_n2585__));
  and1  g1124(.dina(new_new_n4442__), .dinb(new_new_n4573__), .dout(new_new_n2586__));
  or1   g1125(.dina(new_new_n4445__), .dinb(new_new_n4576__), .dout(new_new_n2587__));
  and1  g1126(.dina(new_new_n4579__), .dinb(new_new_n2585__), .dout(new_new_n2588__));
  and1  g1127(.dina(new_new_n2587__), .dinb(new_new_n4582__), .dout(new_new_n2589__));
  and1  g1128(.dina(new_new_n4585__), .dinb(new_new_n1558__), .dout(new_new_n2590__));
  or1   g1129(.dina(new_new_n2588__), .dinb(new_new_n2582__), .dout(new_new_n2591__));
  or1   g1130(.dina(new_new_n2591__), .dinb(new_new_n2590__), .dout(new_new_n2592__));
  and1  g1131(.dina(new_new_n4468__), .dinb(new_new_n4589__), .dout(new_new_n2593__));
  or1   g1132(.dina(new_new_n4461__), .dinb(new_new_n4595__), .dout(new_new_n2594__));
  or1   g1133(.dina(new_new_n4598__), .dinb(new_new_n2592__), .dout(new_new_n2595__));
  or1   g1134(.dina(new_new_n1986__), .dinb(new_new_n1951__), .dout(new_new_n2596__));
  or1   g1135(.dina(new_new_n1985__), .dinb(new_new_n1952__), .dout(new_new_n2597__));
  and1  g1136(.dina(new_new_n2597__), .dinb(new_new_n2596__), .dout(new_new_n2598__));
  or1   g1137(.dina(new_new_n2598__), .dinb(new_new_n4602__), .dout(new_new_n2599__));
  or1   g1138(.dina(new_new_n4464__), .dinb(new_new_n4603__), .dout(new_new_n2600__));
  or1   g1139(.dina(new_new_n2600__), .dinb(new_new_n4477__), .dout(new_new_n2601__));
  or1   g1140(.dina(new_new_n2601__), .dinb(new_new_n4605__), .dout(new_new_n2602__));
  and1  g1141(.dina(new_new_n2602__), .dinb(new_new_n2599__), .dout(new_new_n2603__));
  or1   g1142(.dina(new_new_n2603__), .dinb(new_new_n4589__), .dout(new_new_n2604__));
  and1  g1143(.dina(new_new_n1693__), .dinb(new_new_n4607__), .dout(new_new_n2605__));
  and1  g1144(.dina(new_new_n1694__), .dinb(new_new_n4608__), .dout(new_new_n2606__));
  or1   g1145(.dina(new_new_n2606__), .dinb(new_new_n2605__), .dout(new_new_n2607__));
  and1  g1146(.dina(new_new_n4609__), .dinb(new_new_n4460__), .dout(new_new_n2608__));
  and1  g1147(.dina(new_new_n4609__), .dinb(new_new_n4595__), .dout(new_new_n2609__));
  and1  g1148(.dina(new_new_n2530__), .dinb(new_new_n4605__), .dout(new_new_n2610__));
  or1   g1149(.dina(new_new_n4463__), .dinb(new_new_n4602__), .dout(new_new_n2611__));
  and1  g1150(.dina(new_new_n2610__), .dinb(new_new_n4462__), .dout(new_new_n2612__));
  and1  g1151(.dina(new_new_n2611__), .dinb(new_new_n4603__), .dout(new_new_n2613__));
  or1   g1152(.dina(new_new_n2613__), .dinb(new_new_n2612__), .dout(new_new_n2614__));
  and1  g1153(.dina(new_new_n2614__), .dinb(new_new_n4594__), .dout(new_new_n2615__));
  or1   g1154(.dina(new_new_n2091__), .dinb(new_new_n4506__), .dout(new_new_n2616__));
  or1   g1155(.dina(new_new_n2111__), .dinb(new_new_n4524__), .dout(new_new_n2617__));
  or1   g1156(.dina(new_new_n2032__), .dinb(new_new_n4612__), .dout(new_new_n2618__));
  or1   g1157(.dina(new_new_n2051__), .dinb(new_new_n4482__), .dout(new_new_n2619__));
  or1   g1158(.dina(new_new_n2131__), .dinb(new_new_n4487__), .dout(new_new_n2620__));
  or1   g1159(.dina(new_new_n1991__), .dinb(new_new_n4492__), .dout(new_new_n2621__));
  or1   g1160(.dina(new_new_n2072__), .dinb(new_new_n4497__), .dout(new_new_n2622__));
  or1   g1161(.dina(new_new_n2011__), .dinb(new_new_n4502__), .dout(new_new_n2623__));
  and1  g1162(.dina(new_new_n2617__), .dinb(new_new_n2616__), .dout(new_new_n2624__));
  and1  g1163(.dina(new_new_n2624__), .dinb(new_new_n2618__), .dout(new_new_n2625__));
  and1  g1164(.dina(new_new_n2625__), .dinb(new_new_n2619__), .dout(new_new_n2626__));
  and1  g1165(.dina(new_new_n2626__), .dinb(new_new_n2620__), .dout(new_new_n2627__));
  and1  g1166(.dina(new_new_n2627__), .dinb(new_new_n2621__), .dout(new_new_n2628__));
  and1  g1167(.dina(new_new_n2628__), .dinb(new_new_n2622__), .dout(new_new_n2629__));
  and1  g1168(.dina(new_new_n2629__), .dinb(new_new_n2623__), .dout(new_new_n2630__));
  and1  g1169(.dina(new_new_n2630__), .dinb(new_new_n4514__), .dout(new_new_n2631__));
  or1   g1170(.dina(new_new_n2101__), .dinb(new_new_n4615__), .dout(new_new_n2632__));
  or1   g1171(.dina(new_new_n2121__), .dinb(new_new_n4534__), .dout(new_new_n2633__));
  or1   g1172(.dina(new_new_n2042__), .dinb(new_new_n4540__), .dout(new_new_n2634__));
  or1   g1173(.dina(new_new_n2061__), .dinb(new_new_n4545__), .dout(new_new_n2635__));
  or1   g1174(.dina(new_new_n2141__), .dinb(new_new_n4551__), .dout(new_new_n2636__));
  or1   g1175(.dina(new_new_n2001__), .dinb(new_new_n4556__), .dout(new_new_n2637__));
  or1   g1176(.dina(new_new_n2082__), .dinb(new_new_n4520__), .dout(new_new_n2638__));
  or1   g1177(.dina(new_new_n2021__), .dinb(new_new_n4617__), .dout(new_new_n2639__));
  and1  g1178(.dina(new_new_n2633__), .dinb(new_new_n2632__), .dout(new_new_n2640__));
  and1  g1179(.dina(new_new_n2640__), .dinb(new_new_n2634__), .dout(new_new_n2641__));
  and1  g1180(.dina(new_new_n2641__), .dinb(new_new_n2635__), .dout(new_new_n2642__));
  and1  g1181(.dina(new_new_n2642__), .dinb(new_new_n2636__), .dout(new_new_n2643__));
  and1  g1182(.dina(new_new_n2643__), .dinb(new_new_n2637__), .dout(new_new_n2644__));
  and1  g1183(.dina(new_new_n2644__), .dinb(new_new_n2638__), .dout(new_new_n2645__));
  and1  g1184(.dina(new_new_n2645__), .dinb(new_new_n2639__), .dout(new_new_n2646__));
  and1  g1185(.dina(new_new_n2646__), .dinb(new_new_n4561__), .dout(new_new_n2647__));
  or1   g1186(.dina(new_new_n2647__), .dinb(new_new_n2631__), .dout(new_new_n2648__));
  and1  g1187(.dina(new_new_n2648__), .dinb(new_new_n4568__), .dout(new_new_n2649__));
  or1   g1188(.dina(new_new_n1915__), .dinb(new_new_n1911__), .dout(new_new_n2650__));
  or1   g1189(.dina(new_new_n1916__), .dinb(new_new_n1912__), .dout(new_new_n2651__));
  and1  g1190(.dina(new_new_n2651__), .dinb(new_new_n2650__), .dout(new_new_n2652__));
  and1  g1191(.dina(new_new_n4441__), .dinb(new_new_n4454__), .dout(new_new_n2653__));
  or1   g1192(.dina(new_new_n4446__), .dinb(new_new_n4456__), .dout(new_new_n2654__));
  and1  g1193(.dina(new_new_n2653__), .dinb(new_new_n4573__), .dout(new_new_n2655__));
  or1   g1194(.dina(new_new_n2654__), .dinb(new_new_n4576__), .dout(new_new_n2656__));
  and1  g1195(.dina(new_new_n4619__), .dinb(new_new_n2652__), .dout(new_new_n2657__));
  and1  g1196(.dina(new_new_n4620__), .dinb(new_new_n4513__), .dout(new_new_n2658__));
  or1   g1197(.dina(new_new_n4621__), .dinb(new_new_n4560__), .dout(new_new_n2659__));
  and1  g1198(.dina(new_new_n4623__), .dinb(new_new_n4624__), .dout(new_new_n2660__));
  and1  g1199(.dina(new_new_n4620__), .dinb(new_new_n4577__), .dout(new_new_n2661__));
  or1   g1200(.dina(new_new_n4621__), .dinb(new_new_n4574__), .dout(new_new_n2662__));
  and1  g1201(.dina(new_new_n4626__), .dinb(new_new_n4628__), .dout(new_new_n2663__));
  or1   g1202(.dina(new_new_n4630__), .dinb(new_new_n4623__), .dout(new_new_n2664__));
  and1  g1203(.dina(new_new_n4631__), .dinb(new_new_n1638__), .dout(new_new_n2665__));
  or1   g1204(.dina(new_new_n4630__), .dinb(new_new_n2660__), .dout(new_new_n2666__));
  or1   g1205(.dina(new_new_n2666__), .dinb(new_new_n2665__), .dout(new_new_n2667__));
  and1  g1206(.dina(new_new_n4633__), .dinb(new_new_n4582__), .dout(new_new_n2668__));
  or1   g1207(.dina(new_new_n4619__), .dinb(new_new_n4569__), .dout(new_new_n2669__));
  and1  g1208(.dina(new_new_n4634__), .dinb(new_new_n2667__), .dout(new_new_n2670__));
  or1   g1209(.dina(new_new_n2657__), .dinb(new_new_n2649__), .dout(new_new_n2671__));
  or1   g1210(.dina(new_new_n2671__), .dinb(new_new_n2670__), .dout(new_new_n2672__));
  or1   g1211(.dina(new_new_n2672__), .dinb(new_new_n4598__), .dout(new_new_n2673__));
  and1  g1212(.dina(new_new_n2094__), .dinb(new_new_n1867__), .dout(new_new_n2674__));
  and1  g1213(.dina(new_new_n2114__), .dinb(new_new_n4635__), .dout(new_new_n2675__));
  and1  g1214(.dina(new_new_n2033__), .dinb(new_new_n4636__), .dout(new_new_n2676__));
  and1  g1215(.dina(new_new_n2054__), .dinb(new_new_n4637__), .dout(new_new_n2677__));
  and1  g1216(.dina(new_new_n2134__), .dinb(new_new_n4638__), .dout(new_new_n2678__));
  and1  g1217(.dina(new_new_n1994__), .dinb(new_new_n4639__), .dout(new_new_n2679__));
  and1  g1218(.dina(new_new_n2073__), .dinb(new_new_n4640__), .dout(new_new_n2680__));
  and1  g1219(.dina(new_new_n2014__), .dinb(new_new_n1475__), .dout(new_new_n2681__));
  or1   g1220(.dina(new_new_n2675__), .dinb(new_new_n2674__), .dout(new_new_n2682__));
  or1   g1221(.dina(new_new_n2682__), .dinb(new_new_n2676__), .dout(new_new_n2683__));
  or1   g1222(.dina(new_new_n2683__), .dinb(new_new_n2677__), .dout(new_new_n2684__));
  or1   g1223(.dina(new_new_n2684__), .dinb(new_new_n2678__), .dout(new_new_n2685__));
  or1   g1224(.dina(new_new_n2685__), .dinb(new_new_n2679__), .dout(new_new_n2686__));
  or1   g1225(.dina(new_new_n2686__), .dinb(new_new_n2680__), .dout(new_new_n2687__));
  or1   g1226(.dina(new_new_n2687__), .dinb(new_new_n2681__), .dout(new_new_n2688__));
  or1   g1227(.dina(new_new_n2688__), .dinb(new_new_n4562__), .dout(new_new_n2689__));
  and1  g1228(.dina(new_new_n2104__), .dinb(new_new_n4641__), .dout(new_new_n2690__));
  and1  g1229(.dina(new_new_n2124__), .dinb(new_new_n4642__), .dout(new_new_n2691__));
  and1  g1230(.dina(new_new_n2043__), .dinb(new_new_n1898__), .dout(new_new_n2692__));
  and1  g1231(.dina(new_new_n2064__), .dinb(new_new_n4643__), .dout(new_new_n2693__));
  and1  g1232(.dina(new_new_n2144__), .dinb(new_new_n4644__), .dout(new_new_n2694__));
  and1  g1233(.dina(new_new_n2004__), .dinb(new_new_n4645__), .dout(new_new_n2695__));
  and1  g1234(.dina(new_new_n2083__), .dinb(new_new_n4646__), .dout(new_new_n2696__));
  and1  g1235(.dina(new_new_n2024__), .dinb(new_new_n4647__), .dout(new_new_n2697__));
  or1   g1236(.dina(new_new_n2691__), .dinb(new_new_n2690__), .dout(new_new_n2698__));
  or1   g1237(.dina(new_new_n2698__), .dinb(new_new_n2692__), .dout(new_new_n2699__));
  or1   g1238(.dina(new_new_n2699__), .dinb(new_new_n2693__), .dout(new_new_n2700__));
  or1   g1239(.dina(new_new_n2700__), .dinb(new_new_n2694__), .dout(new_new_n2701__));
  or1   g1240(.dina(new_new_n2701__), .dinb(new_new_n2695__), .dout(new_new_n2702__));
  or1   g1241(.dina(new_new_n2702__), .dinb(new_new_n2696__), .dout(new_new_n2703__));
  or1   g1242(.dina(new_new_n2703__), .dinb(new_new_n2697__), .dout(new_new_n2704__));
  or1   g1243(.dina(new_new_n2704__), .dinb(new_new_n4515__), .dout(new_new_n2705__));
  and1  g1244(.dina(new_new_n2705__), .dinb(new_new_n2689__), .dout(new_new_n2706__));
  or1   g1245(.dina(new_new_n2706__), .dinb(new_new_n4583__), .dout(new_new_n2707__));
  and1  g1246(.dina(new_new_n1910__), .dinb(new_new_n1908__), .dout(new_new_n2708__));
  and1  g1247(.dina(new_new_n1909__), .dinb(new_new_n1907__), .dout(new_new_n2709__));
  or1   g1248(.dina(new_new_n2709__), .dinb(new_new_n2708__), .dout(new_new_n2710__));
  or1   g1249(.dina(new_new_n2710__), .dinb(new_new_n4633__), .dout(new_new_n2711__));
  or1   g1250(.dina(new_new_n4628__), .dinb(new_new_n4648__), .dout(new_new_n2712__));
  or1   g1251(.dina(new_new_n4649__), .dinb(new_new_n4440__), .dout(new_new_n2713__));
  and1  g1252(.dina(new_new_n2712__), .dinb(new_new_n4626__), .dout(new_new_n2714__));
  and1  g1253(.dina(new_new_n2714__), .dinb(new_new_n2713__), .dout(new_new_n2715__));
  or1   g1254(.dina(new_new_n2715__), .dinb(new_new_n4650__), .dout(new_new_n2716__));
  and1  g1255(.dina(new_new_n2711__), .dinb(new_new_n2707__), .dout(new_new_n2717__));
  and1  g1256(.dina(new_new_n2717__), .dinb(new_new_n2716__), .dout(new_new_n2718__));
  and1  g1257(.dina(new_new_n2718__), .dinb(new_new_n4651__), .dout(new_new_n2719__));
  or1   g1258(.dina(new_new_n2095__), .dinb(new_new_n4498__), .dout(new_new_n2720__));
  or1   g1259(.dina(new_new_n2115__), .dinb(new_new_n4535__), .dout(new_new_n2721__));
  or1   g1260(.dina(new_new_n2036__), .dinb(new_new_n4529__), .dout(new_new_n2722__));
  or1   g1261(.dina(new_new_n2055__), .dinb(new_new_n4525__), .dout(new_new_n2723__));
  or1   g1262(.dina(new_new_n2135__), .dinb(new_new_n4612__), .dout(new_new_n2724__));
  or1   g1263(.dina(new_new_n1995__), .dinb(new_new_n4483__), .dout(new_new_n2725__));
  or1   g1264(.dina(new_new_n2076__), .dinb(new_new_n4488__), .dout(new_new_n2726__));
  or1   g1265(.dina(new_new_n2015__), .dinb(new_new_n4493__), .dout(new_new_n2727__));
  and1  g1266(.dina(new_new_n2721__), .dinb(new_new_n2720__), .dout(new_new_n2728__));
  and1  g1267(.dina(new_new_n2728__), .dinb(new_new_n2722__), .dout(new_new_n2729__));
  and1  g1268(.dina(new_new_n2729__), .dinb(new_new_n2723__), .dout(new_new_n2730__));
  and1  g1269(.dina(new_new_n2730__), .dinb(new_new_n2724__), .dout(new_new_n2731__));
  and1  g1270(.dina(new_new_n2731__), .dinb(new_new_n2725__), .dout(new_new_n2732__));
  and1  g1271(.dina(new_new_n2732__), .dinb(new_new_n2726__), .dout(new_new_n2733__));
  and1  g1272(.dina(new_new_n2733__), .dinb(new_new_n2727__), .dout(new_new_n2734__));
  and1  g1273(.dina(new_new_n2734__), .dinb(new_new_n4515__), .dout(new_new_n2735__));
  or1   g1274(.dina(new_new_n2105__), .dinb(new_new_n1876__), .dout(new_new_n2736__));
  or1   g1275(.dina(new_new_n2125__), .dinb(new_new_n4546__), .dout(new_new_n2737__));
  or1   g1276(.dina(new_new_n2046__), .dinb(new_new_n4552__), .dout(new_new_n2738__));
  or1   g1277(.dina(new_new_n2065__), .dinb(new_new_n4555__), .dout(new_new_n2739__));
  or1   g1278(.dina(new_new_n2145__), .dinb(new_new_n4521__), .dout(new_new_n2740__));
  or1   g1279(.dina(new_new_n2005__), .dinb(new_new_n4617__), .dout(new_new_n2741__));
  or1   g1280(.dina(new_new_n2086__), .dinb(new_new_n4615__), .dout(new_new_n2742__));
  or1   g1281(.dina(new_new_n2025__), .dinb(new_new_n1874__), .dout(new_new_n2743__));
  and1  g1282(.dina(new_new_n2737__), .dinb(new_new_n2736__), .dout(new_new_n2744__));
  and1  g1283(.dina(new_new_n2744__), .dinb(new_new_n2738__), .dout(new_new_n2745__));
  and1  g1284(.dina(new_new_n2745__), .dinb(new_new_n2739__), .dout(new_new_n2746__));
  and1  g1285(.dina(new_new_n2746__), .dinb(new_new_n2740__), .dout(new_new_n2747__));
  and1  g1286(.dina(new_new_n2747__), .dinb(new_new_n2741__), .dout(new_new_n2748__));
  and1  g1287(.dina(new_new_n2748__), .dinb(new_new_n2742__), .dout(new_new_n2749__));
  and1  g1288(.dina(new_new_n2749__), .dinb(new_new_n2743__), .dout(new_new_n2750__));
  and1  g1289(.dina(new_new_n2750__), .dinb(new_new_n4562__), .dout(new_new_n2751__));
  or1   g1290(.dina(new_new_n2751__), .dinb(new_new_n2735__), .dout(new_new_n2752__));
  and1  g1291(.dina(new_new_n2752__), .dinb(new_new_n4569__), .dout(new_new_n2753__));
  or1   g1292(.dina(new_new_n1905__), .dinb(new_new_n1903__), .dout(new_new_n2754__));
  or1   g1293(.dina(new_new_n1906__), .dinb(new_new_n1904__), .dout(new_new_n2755__));
  and1  g1294(.dina(new_new_n2755__), .dinb(new_new_n2754__), .dout(new_new_n2756__));
  and1  g1295(.dina(new_new_n2756__), .dinb(new_new_n4618__), .dout(new_new_n2757__));
  or1   g1296(.dina(new_new_n1987__), .dinb(new_new_n1971__), .dout(new_new_n2758__));
  or1   g1297(.dina(new_new_n1888__), .dinb(new_new_n1804__), .dout(new_new_n2759__));
  and1  g1298(.dina(new_new_n2759__), .dinb(new_new_n2758__), .dout(new_new_n2760__));
  and1  g1299(.dina(new_new_n2760__), .dinb(new_new_n4622__), .dout(new_new_n2761__));
  or1   g1300(.dina(new_new_n1709__), .dinb(new_new_n4652__), .dout(new_new_n2762__));
  and1  g1301(.dina(new_new_n2762__), .dinb(new_new_n4629__), .dout(new_new_n2763__));
  and1  g1302(.dina(new_new_n4631__), .dinb(new_new_n1634__), .dout(new_new_n2764__));
  or1   g1303(.dina(new_new_n2763__), .dinb(new_new_n2761__), .dout(new_new_n2765__));
  or1   g1304(.dina(new_new_n2765__), .dinb(new_new_n2764__), .dout(new_new_n2766__));
  and1  g1305(.dina(new_new_n2766__), .dinb(new_new_n4634__), .dout(new_new_n2767__));
  or1   g1306(.dina(new_new_n2757__), .dinb(new_new_n2753__), .dout(new_new_n2768__));
  or1   g1307(.dina(new_new_n2768__), .dinb(new_new_n2767__), .dout(new_new_n2769__));
  or1   g1308(.dina(new_new_n2769__), .dinb(new_new_n4599__), .dout(new_new_n2770__));
  and1  g1309(.dina(new_new_n2098__), .dinb(new_new_n4640__), .dout(new_new_n2771__));
  and1  g1310(.dina(new_new_n2118__), .dinb(new_new_n4642__), .dout(new_new_n2772__));
  and1  g1311(.dina(new_new_n2037__), .dinb(new_new_n1890__), .dout(new_new_n2773__));
  and1  g1312(.dina(new_new_n2058__), .dinb(new_new_n4635__), .dout(new_new_n2774__));
  and1  g1313(.dina(new_new_n2138__), .dinb(new_new_n4636__), .dout(new_new_n2775__));
  and1  g1314(.dina(new_new_n1998__), .dinb(new_new_n4637__), .dout(new_new_n2776__));
  and1  g1315(.dina(new_new_n2077__), .dinb(new_new_n4638__), .dout(new_new_n2777__));
  and1  g1316(.dina(new_new_n2018__), .dinb(new_new_n4639__), .dout(new_new_n2778__));
  or1   g1317(.dina(new_new_n2772__), .dinb(new_new_n2771__), .dout(new_new_n2779__));
  or1   g1318(.dina(new_new_n2779__), .dinb(new_new_n2773__), .dout(new_new_n2780__));
  or1   g1319(.dina(new_new_n2780__), .dinb(new_new_n2774__), .dout(new_new_n2781__));
  or1   g1320(.dina(new_new_n2781__), .dinb(new_new_n2775__), .dout(new_new_n2782__));
  or1   g1321(.dina(new_new_n2782__), .dinb(new_new_n2776__), .dout(new_new_n2783__));
  or1   g1322(.dina(new_new_n2783__), .dinb(new_new_n2777__), .dout(new_new_n2784__));
  or1   g1323(.dina(new_new_n2784__), .dinb(new_new_n2778__), .dout(new_new_n2785__));
  or1   g1324(.dina(new_new_n2785__), .dinb(new_new_n4564__), .dout(new_new_n2786__));
  and1  g1325(.dina(new_new_n2108__), .dinb(new_new_n1877__), .dout(new_new_n2787__));
  and1  g1326(.dina(new_new_n2128__), .dinb(new_new_n4643__), .dout(new_new_n2788__));
  and1  g1327(.dina(new_new_n2047__), .dinb(new_new_n4644__), .dout(new_new_n2789__));
  and1  g1328(.dina(new_new_n2068__), .dinb(new_new_n4645__), .dout(new_new_n2790__));
  and1  g1329(.dina(new_new_n2148__), .dinb(new_new_n4646__), .dout(new_new_n2791__));
  and1  g1330(.dina(new_new_n2008__), .dinb(new_new_n4647__), .dout(new_new_n2792__));
  and1  g1331(.dina(new_new_n2087__), .dinb(new_new_n4641__), .dout(new_new_n2793__));
  and1  g1332(.dina(new_new_n2028__), .dinb(new_new_n1875__), .dout(new_new_n2794__));
  or1   g1333(.dina(new_new_n2788__), .dinb(new_new_n2787__), .dout(new_new_n2795__));
  or1   g1334(.dina(new_new_n2795__), .dinb(new_new_n2789__), .dout(new_new_n2796__));
  or1   g1335(.dina(new_new_n2796__), .dinb(new_new_n2790__), .dout(new_new_n2797__));
  or1   g1336(.dina(new_new_n2797__), .dinb(new_new_n2791__), .dout(new_new_n2798__));
  or1   g1337(.dina(new_new_n2798__), .dinb(new_new_n2792__), .dout(new_new_n2799__));
  or1   g1338(.dina(new_new_n2799__), .dinb(new_new_n2793__), .dout(new_new_n2800__));
  or1   g1339(.dina(new_new_n2800__), .dinb(new_new_n2794__), .dout(new_new_n2801__));
  or1   g1340(.dina(new_new_n2801__), .dinb(new_new_n4517__), .dout(new_new_n2802__));
  and1  g1341(.dina(new_new_n2802__), .dinb(new_new_n2786__), .dout(new_new_n2803__));
  or1   g1342(.dina(new_new_n2803__), .dinb(new_new_n4583__), .dout(new_new_n2804__));
  and1  g1343(.dina(new_new_n1918__), .dinb(new_new_n1914__), .dout(new_new_n2805__));
  and1  g1344(.dina(new_new_n1917__), .dinb(new_new_n1913__), .dout(new_new_n2806__));
  or1   g1345(.dina(new_new_n2806__), .dinb(new_new_n2805__), .dout(new_new_n2807__));
  or1   g1346(.dina(new_new_n2807__), .dinb(new_new_n4632__), .dout(new_new_n2808__));
  and1  g1347(.dina(new_new_n1974__), .dinb(new_new_n1966__), .dout(new_new_n2809__));
  and1  g1348(.dina(new_new_n4653__), .dinb(new_new_n1805__), .dout(new_new_n2810__));
  or1   g1349(.dina(new_new_n2810__), .dinb(new_new_n2809__), .dout(new_new_n2811__));
  or1   g1350(.dina(new_new_n2811__), .dinb(new_new_n4627__), .dout(new_new_n2812__));
  and1  g1351(.dina(new_new_n4654__), .dinb(new_new_n4655__), .dout(new_new_n2813__));
  or1   g1352(.dina(new_new_n2813__), .dinb(new_new_n4625__), .dout(new_new_n2814__));
  or1   g1353(.dina(new_new_n4649__), .dinb(new_new_n4652__), .dout(new_new_n2815__));
  and1  g1354(.dina(new_new_n2814__), .dinb(new_new_n2812__), .dout(new_new_n2816__));
  and1  g1355(.dina(new_new_n2816__), .dinb(new_new_n2815__), .dout(new_new_n2817__));
  or1   g1356(.dina(new_new_n2817__), .dinb(new_new_n4650__), .dout(new_new_n2818__));
  and1  g1357(.dina(new_new_n2808__), .dinb(new_new_n2804__), .dout(new_new_n2819__));
  and1  g1358(.dina(new_new_n2819__), .dinb(new_new_n2818__), .dout(new_new_n2820__));
  and1  g1359(.dina(new_new_n2820__), .dinb(new_new_n4651__), .dout(new_new_n2821__));
  and1  g1360(.dina(new_new_n1940__), .dinb(new_new_n1935__), .dout(new_new_n2822__));
  or1   g1361(.dina(new_new_n1939__), .dinb(new_new_n1936__), .dout(new_new_n2823__));
  and1  g1362(.dina(new_new_n2823__), .dinb(new_new_n4657__), .dout(new_new_n2824__));
  and1  g1363(.dina(new_new_n2822__), .dinb(new_new_n4659__), .dout(new_new_n2825__));
  or1   g1364(.dina(new_new_n2825__), .dinb(new_new_n2824__), .dout(new_new_n2826__));
  or1   g1365(.dina(new_new_n2826__), .dinb(new_new_n4590__), .dout(new_new_n2827__));
  and1  g1366(.dina(new_new_n1938__), .dinb(new_new_n1933__), .dout(new_new_n2828__));
  or1   g1367(.dina(new_new_n1937__), .dinb(new_new_n1934__), .dout(new_new_n2829__));
  and1  g1368(.dina(new_new_n2829__), .dinb(new_new_n4604__), .dout(new_new_n2830__));
  and1  g1369(.dina(new_new_n2828__), .dinb(new_new_n4601__), .dout(new_new_n2831__));
  or1   g1370(.dina(new_new_n2831__), .dinb(new_new_n2830__), .dout(new_new_n2832__));
  or1   g1371(.dina(new_new_n2832__), .dinb(new_new_n4590__), .dout(new_new_n2833__));
  and1  g1372(.dina(new_new_n4660__), .dinb(new_new_n1716__), .dout(new_new_n2834__));
  or1   g1373(.dina(new_new_n1724__), .dinb(new_new_n1715__), .dout(new_new_n2835__));
  and1  g1374(.dina(new_new_n4661__), .dinb(new_new_n4662__), .dout(new_new_n2836__));
  or1   g1375(.dina(new_new_n4663__), .dinb(new_new_n1726__), .dout(new_new_n2837__));
  and1  g1376(.dina(new_new_n4666__), .dinb(new_new_n4671__), .dout(new_new_n2838__));
  or1   g1377(.dina(new_new_n4674__), .dinb(new_new_n2510__), .dout(new_new_n2839__));
  and1  g1378(.dina(new_new_n1788__), .dinb(new_new_n1786__), .dout(new_new_n2840__));
  or1   g1379(.dina(new_new_n1787__), .dinb(new_new_n1785__), .dout(new_new_n2841__));
  and1  g1380(.dina(new_new_n2178__), .dinb(new_new_n2176__), .dout(new_new_n2842__));
  or1   g1381(.dina(new_new_n2177__), .dinb(new_new_n2175__), .dout(new_new_n2843__));
  and1  g1382(.dina(new_new_n2842__), .dinb(new_new_n2194__), .dout(new_new_n2844__));
  or1   g1383(.dina(new_new_n2843__), .dinb(new_new_n2193__), .dout(new_new_n2845__));
  and1  g1384(.dina(new_new_n2845__), .dinb(new_new_n2840__), .dout(new_new_n2846__));
  or1   g1385(.dina(new_new_n2844__), .dinb(new_new_n2841__), .dout(new_new_n2847__));
  and1  g1386(.dina(new_new_n4680__), .dinb(new_new_n4683__), .dout(new_new_n2848__));
  or1   g1387(.dina(new_new_n4686__), .dinb(new_new_n4688__), .dout(new_new_n2849__));
  and1  g1388(.dina(new_new_n2848__), .dinb(new_new_n2151__), .dout(new_new_n2850__));
  or1   g1389(.dina(new_new_n2849__), .dinb(new_new_n2152__), .dout(new_new_n2851__));
  and1  g1390(.dina(new_new_n2850__), .dinb(new_new_n4690__), .dout(new_new_n2852__));
  or1   g1391(.dina(new_new_n2851__), .dinb(new_new_n4693__), .dout(new_new_n2853__));
  and1  g1392(.dina(new_new_n2224__), .dinb(new_new_n1960__), .dout(new_new_n2854__));
  or1   g1393(.dina(new_new_n2223__), .dinb(new_new_n1959__), .dout(new_new_n2855__));
  and1  g1394(.dina(new_new_n2215__), .dinb(new_new_n2159__), .dout(new_new_n2856__));
  or1   g1395(.dina(new_new_n2216__), .dinb(new_new_n2160__), .dout(new_new_n2857__));
  and1  g1396(.dina(new_new_n2857__), .dinb(new_new_n2855__), .dout(new_new_n2858__));
  or1   g1397(.dina(new_new_n2856__), .dinb(new_new_n2854__), .dout(new_new_n2859__));
  and1  g1398(.dina(new_new_n4694__), .dinb(new_new_n4695__), .dout(new_new_n2860__));
  or1   g1399(.dina(new_new_n4696__), .dinb(new_new_n4697__), .dout(new_new_n2861__));
  and1  g1400(.dina(new_new_n4696__), .dinb(new_new_n4697__), .dout(new_new_n2862__));
  or1   g1401(.dina(new_new_n4694__), .dinb(new_new_n4695__), .dout(new_new_n2863__));
  and1  g1402(.dina(new_new_n2863__), .dinb(new_new_n2861__), .dout(new_new_n2864__));
  or1   g1403(.dina(new_new_n2862__), .dinb(new_new_n2860__), .dout(new_new_n2865__));
  or1   g1404(.dina(new_new_n4699__), .dinb(new_new_n4470__), .dout(new_new_n2866__));
  and1  g1405(.dina(new_new_n4701__), .dinb(new_new_n4702__), .dout(new_new_n2867__));
  or1   g1406(.dina(new_new_n4704__), .dinb(new_new_n1668__), .dout(new_new_n2868__));
  and1  g1407(.dina(new_new_n2867__), .dinb(new_new_n4705__), .dout(new_new_n2869__));
  or1   g1408(.dina(new_new_n2868__), .dinb(new_new_n4706__), .dout(new_new_n2870__));
  and1  g1409(.dina(new_new_n4701__), .dinb(new_new_n4707__), .dout(new_new_n2871__));
  or1   g1410(.dina(new_new_n4704__), .dinb(new_new_n4708__), .dout(new_new_n2872__));
  and1  g1411(.dina(new_new_n2871__), .dinb(new_new_n4709__), .dout(new_new_n2873__));
  or1   g1412(.dina(new_new_n2872__), .dinb(new_new_n4710__), .dout(new_new_n2874__));
  and1  g1413(.dina(new_new_n2874__), .dinb(new_new_n2870__), .dout(new_new_n2875__));
  or1   g1414(.dina(new_new_n2873__), .dinb(new_new_n2869__), .dout(new_new_n2876__));
  and1  g1415(.dina(new_new_n4712__), .dinb(new_new_n4713__), .dout(new_new_n2877__));
  or1   g1416(.dina(new_new_n4715__), .dinb(new_new_n4716__), .dout(new_new_n2878__));
  and1  g1417(.dina(new_new_n2877__), .dinb(new_new_n4709__), .dout(new_new_n2879__));
  or1   g1418(.dina(new_new_n2878__), .dinb(new_new_n4710__), .dout(new_new_n2880__));
  and1  g1419(.dina(new_new_n4712__), .dinb(new_new_n4717__), .dout(new_new_n2881__));
  or1   g1420(.dina(new_new_n4715__), .dinb(new_new_n4719__), .dout(new_new_n2882__));
  and1  g1421(.dina(new_new_n2881__), .dinb(new_new_n4705__), .dout(new_new_n2883__));
  or1   g1422(.dina(new_new_n2882__), .dinb(new_new_n4706__), .dout(new_new_n2884__));
  and1  g1423(.dina(new_new_n2884__), .dinb(new_new_n2880__), .dout(new_new_n2885__));
  or1   g1424(.dina(new_new_n2883__), .dinb(new_new_n2879__), .dout(new_new_n2886__));
  and1  g1425(.dina(new_new_n2885__), .dinb(new_new_n4711__), .dout(new_new_n2887__));
  or1   g1426(.dina(new_new_n2886__), .dinb(new_new_n4714__), .dout(new_new_n2888__));
  and1  g1427(.dina(new_new_n2888__), .dinb(new_new_n2875__), .dout(new_new_n2889__));
  or1   g1428(.dina(new_new_n2887__), .dinb(new_new_n4720__), .dout(new_new_n2890__));
  and1  g1429(.dina(new_new_n4723__), .dinb(new_new_n4726__), .dout(new_new_n2891__));
  or1   g1430(.dina(new_new_n4728__), .dinb(new_new_n2154__), .dout(new_new_n2892__));
  or1   g1431(.dina(new_new_n2892__), .dinb(new_new_n1852__), .dout(new_new_n2893__));
  or1   g1432(.dina(new_new_n2893__), .dinb(new_new_n1742__), .dout(new_new_n2894__));
  or1   g1433(.dina(new_new_n1970__), .dinb(new_new_n1921__), .dout(new_new_n2895__));
  or1   g1434(.dina(new_new_n1969__), .dinb(new_new_n1922__), .dout(new_new_n2896__));
  and1  g1435(.dina(new_new_n2896__), .dinb(new_new_n2895__), .dout(new_new_n2897__));
  or1   g1436(.dina(new_new_n4730__), .dinb(new_new_n4470__), .dout(new_new_n2898__));
  and1  g1437(.dina(new_new_n4700__), .dinb(new_new_n1929__), .dout(new_new_n2899__));
  or1   g1438(.dina(new_new_n4703__), .dinb(new_new_n1930__), .dout(new_new_n2900__));
  or1   g1439(.dina(new_new_n4731__), .dinb(new_new_n4732__), .dout(new_new_n2901__));
  or1   g1440(.dina(new_new_n2901__), .dinb(new_new_n4733__), .dout(new_new_n2902__));
  and1  g1441(.dina(new_new_n4734__), .dinb(new_new_n4735__), .dout(new_new_n2903__));
  and1  g1442(.dina(new_new_n2903__), .dinb(new_new_n4736__), .dout(new_new_n2904__));
  and1  g1443(.dina(new_new_n4737__), .dinb(new_new_n4738__), .dout(new_new_n2905__));
  and1  g1444(.dina(new_new_n2905__), .dinb(new_new_n4739__), .dout(new_new_n2906__));
  and1  g1445(.dina(new_new_n4740__), .dinb(new_new_n4741__), .dout(new_new_n2907__));
  and1  g1446(.dina(new_new_n2907__), .dinb(new_new_n4742__), .dout(new_new_n2908__));
  and1  g1447(.dina(new_new_n4607__), .dinb(new_new_n1608__), .dout(new_new_n2909__));
  or1   g1448(.dina(new_new_n4608__), .dinb(new_new_n1607__), .dout(new_new_n2910__));
  and1  g1449(.dina(new_new_n4743__), .dinb(new_new_n4744__), .dout(new_new_n2911__));
  or1   g1450(.dina(new_new_n4745__), .dinb(new_new_n4746__), .dout(new_new_n2912__));
  and1  g1451(.dina(new_new_n4745__), .dinb(new_new_n4746__), .dout(new_new_n2913__));
  or1   g1452(.dina(new_new_n4743__), .dinb(new_new_n4744__), .dout(new_new_n2914__));
  and1  g1453(.dina(new_new_n2914__), .dinb(new_new_n2912__), .dout(new_new_n2915__));
  or1   g1454(.dina(new_new_n2913__), .dinb(new_new_n2911__), .dout(new_new_n2916__));
  or1   g1455(.dina(new_new_n2916__), .dinb(new_new_n2910__), .dout(new_new_n2917__));
  or1   g1456(.dina(new_new_n2915__), .dinb(new_new_n2909__), .dout(new_new_n2918__));
  and1  g1457(.dina(new_new_n2918__), .dinb(new_new_n2917__), .dout(new_new_n2919__));
  or1   g1458(.dina(new_new_n4747__), .dinb(new_new_n4469__), .dout(new_new_n2920__));
  or1   g1459(.dina(new_new_n4749__), .dinb(new_new_n1242__), .dout(new_new_n2921__));
  or1   g1460(.dina(new_new_n4751__), .dinb(new_new_n4493__), .dout(new_new_n2922__));
  or1   g1461(.dina(new_new_n4753__), .dinb(new_new_n4498__), .dout(new_new_n2923__));
  or1   g1462(.dina(new_new_n4501__), .dinb(new_new_n4755__), .dout(new_new_n2924__));
  or1   g1463(.dina(new_new_n4505__), .dinb(new_new_n4757__), .dout(new_new_n2925__));
  or1   g1464(.dina(new_new_n4509__), .dinb(new_new_n4759__), .dout(new_new_n2926__));
  or1   g1465(.dina(new_new_n4479__), .dinb(new_new_n4761__), .dout(new_new_n2927__));
  or1   g1466(.dina(new_new_n4763__), .dinb(new_new_n4764__), .dout(new_new_n2928__));
  and1  g1467(.dina(new_new_n2922__), .dinb(new_new_n2921__), .dout(new_new_n2929__));
  and1  g1468(.dina(new_new_n2929__), .dinb(new_new_n2923__), .dout(new_new_n2930__));
  and1  g1469(.dina(new_new_n2930__), .dinb(new_new_n2924__), .dout(new_new_n2931__));
  and1  g1470(.dina(new_new_n2931__), .dinb(new_new_n2925__), .dout(new_new_n2932__));
  and1  g1471(.dina(new_new_n2932__), .dinb(new_new_n2926__), .dout(new_new_n2933__));
  and1  g1472(.dina(new_new_n2933__), .dinb(new_new_n2927__), .dout(new_new_n2934__));
  and1  g1473(.dina(new_new_n2934__), .dinb(new_new_n2928__), .dout(new_new_n2935__));
  and1  g1474(.dina(new_new_n4451__), .dinb(new_new_n4574__), .dout(new_new_n2936__));
  or1   g1475(.dina(new_new_n4453__), .dinb(new_new_n4577__), .dout(new_new_n2937__));
  and1  g1476(.dina(new_new_n2936__), .dinb(new_new_n2935__), .dout(new_new_n2938__));
  or1   g1477(.dina(new_new_n4766__), .dinb(new_new_n4552__), .dout(new_new_n2939__));
  or1   g1478(.dina(new_new_n4483__), .dinb(new_new_n4768__), .dout(new_new_n2940__));
  or1   g1479(.dina(new_new_n4613__), .dinb(new_new_n4770__), .dout(new_new_n2941__));
  or1   g1480(.dina(new_new_n4525__), .dinb(new_new_n4772__), .dout(new_new_n2942__));
  or1   g1481(.dina(new_new_n4530__), .dinb(new_new_n4774__), .dout(new_new_n2943__));
  or1   g1482(.dina(new_new_n4535__), .dinb(new_new_n4776__), .dout(new_new_n2944__));
  or1   g1483(.dina(new_new_n4541__), .dinb(new_new_n4778__), .dout(new_new_n2945__));
  or1   g1484(.dina(new_new_n4546__), .dinb(new_new_n4780__), .dout(new_new_n2946__));
  and1  g1485(.dina(new_new_n2940__), .dinb(new_new_n2939__), .dout(new_new_n2947__));
  and1  g1486(.dina(new_new_n2947__), .dinb(new_new_n2941__), .dout(new_new_n2948__));
  and1  g1487(.dina(new_new_n2948__), .dinb(new_new_n2942__), .dout(new_new_n2949__));
  and1  g1488(.dina(new_new_n2949__), .dinb(new_new_n2943__), .dout(new_new_n2950__));
  and1  g1489(.dina(new_new_n2950__), .dinb(new_new_n2944__), .dout(new_new_n2951__));
  and1  g1490(.dina(new_new_n2951__), .dinb(new_new_n2945__), .dout(new_new_n2952__));
  and1  g1491(.dina(new_new_n2952__), .dinb(new_new_n2946__), .dout(new_new_n2953__));
  and1  g1492(.dina(new_new_n4517__), .dinb(new_new_n4450__), .dout(new_new_n2954__));
  or1   g1493(.dina(new_new_n4564__), .dinb(new_new_n4452__), .dout(new_new_n2955__));
  and1  g1494(.dina(new_new_n2954__), .dinb(new_new_n2953__), .dout(new_new_n2956__));
  and1  g1495(.dina(new_new_n2955__), .dinb(new_new_n2937__), .dout(new_new_n2957__));
  and1  g1496(.dina(new_new_n2957__), .dinb(new_new_n4781__), .dout(new_new_n2958__));
  or1   g1497(.dina(new_new_n2956__), .dinb(new_new_n2938__), .dout(new_new_n2959__));
  or1   g1498(.dina(new_new_n2959__), .dinb(new_new_n2958__), .dout(new_new_n2960__));
  and1  g1499(.dina(new_new_n2960__), .dinb(new_new_n4571__), .dout(new_new_n2961__));
  or1   g1500(.dina(new_new_n1595__), .dinb(new_new_n1569__), .dout(new_new_n2962__));
  or1   g1501(.dina(new_new_n1596__), .dinb(new_new_n1570__), .dout(new_new_n2963__));
  and1  g1502(.dina(new_new_n2963__), .dinb(new_new_n2962__), .dout(new_new_n2964__));
  and1  g1503(.dina(new_new_n2964__), .dinb(new_new_n4579__), .dout(new_new_n2965__));
  and1  g1504(.dina(new_new_n4585__), .dinb(new_new_n4781__), .dout(new_new_n2966__));
  or1   g1505(.dina(new_new_n2965__), .dinb(new_new_n2961__), .dout(new_new_n2967__));
  or1   g1506(.dina(new_new_n2967__), .dinb(new_new_n2966__), .dout(new_new_n2968__));
  or1   g1507(.dina(new_new_n2968__), .dinb(new_new_n4599__), .dout(new_new_n2969__));
  or1   g1508(.dina(new_new_n4749__), .dinb(new_new_n4764__), .dout(new_new_n2970__));
  or1   g1509(.dina(new_new_n4751__), .dinb(new_new_n4488__), .dout(new_new_n2971__));
  or1   g1510(.dina(new_new_n4753__), .dinb(new_new_n4494__), .dout(new_new_n2972__));
  or1   g1511(.dina(new_new_n4755__), .dinb(new_new_n4499__), .dout(new_new_n2973__));
  or1   g1512(.dina(new_new_n4503__), .dinb(new_new_n4757__), .dout(new_new_n2974__));
  or1   g1513(.dina(new_new_n4507__), .dinb(new_new_n4759__), .dout(new_new_n2975__));
  or1   g1514(.dina(new_new_n4510__), .dinb(new_new_n4761__), .dout(new_new_n2976__));
  or1   g1515(.dina(new_new_n4478__), .dinb(new_new_n4763__), .dout(new_new_n2977__));
  and1  g1516(.dina(new_new_n2971__), .dinb(new_new_n2970__), .dout(new_new_n2978__));
  and1  g1517(.dina(new_new_n2978__), .dinb(new_new_n2972__), .dout(new_new_n2979__));
  and1  g1518(.dina(new_new_n2979__), .dinb(new_new_n2973__), .dout(new_new_n2980__));
  and1  g1519(.dina(new_new_n2980__), .dinb(new_new_n2974__), .dout(new_new_n2981__));
  and1  g1520(.dina(new_new_n2981__), .dinb(new_new_n2975__), .dout(new_new_n2982__));
  and1  g1521(.dina(new_new_n2982__), .dinb(new_new_n2976__), .dout(new_new_n2983__));
  and1  g1522(.dina(new_new_n2983__), .dinb(new_new_n2977__), .dout(new_new_n2984__));
  and1  g1523(.dina(new_new_n2984__), .dinb(new_new_n4518__), .dout(new_new_n2985__));
  or1   g1524(.dina(new_new_n4766__), .dinb(new_new_n4557__), .dout(new_new_n2986__));
  or1   g1525(.dina(new_new_n4613__), .dinb(new_new_n4768__), .dout(new_new_n2987__));
  or1   g1526(.dina(new_new_n4526__), .dinb(new_new_n4770__), .dout(new_new_n2988__));
  or1   g1527(.dina(new_new_n4530__), .dinb(new_new_n4772__), .dout(new_new_n2989__));
  or1   g1528(.dina(new_new_n4537__), .dinb(new_new_n4774__), .dout(new_new_n2990__));
  or1   g1529(.dina(new_new_n4541__), .dinb(new_new_n4776__), .dout(new_new_n2991__));
  or1   g1530(.dina(new_new_n4548__), .dinb(new_new_n4778__), .dout(new_new_n2992__));
  or1   g1531(.dina(new_new_n4780__), .dinb(new_new_n4553__), .dout(new_new_n2993__));
  and1  g1532(.dina(new_new_n2987__), .dinb(new_new_n2986__), .dout(new_new_n2994__));
  and1  g1533(.dina(new_new_n2994__), .dinb(new_new_n2988__), .dout(new_new_n2995__));
  and1  g1534(.dina(new_new_n2995__), .dinb(new_new_n2989__), .dout(new_new_n2996__));
  and1  g1535(.dina(new_new_n2996__), .dinb(new_new_n2990__), .dout(new_new_n2997__));
  and1  g1536(.dina(new_new_n2997__), .dinb(new_new_n2991__), .dout(new_new_n2998__));
  and1  g1537(.dina(new_new_n2998__), .dinb(new_new_n2992__), .dout(new_new_n2999__));
  and1  g1538(.dina(new_new_n2999__), .dinb(new_new_n2993__), .dout(new_new_n3000__));
  and1  g1539(.dina(new_new_n3000__), .dinb(new_new_n4565__), .dout(new_new_n3001__));
  or1   g1540(.dina(new_new_n3001__), .dinb(new_new_n2985__), .dout(new_new_n3002__));
  and1  g1541(.dina(new_new_n3002__), .dinb(new_new_n4571__), .dout(new_new_n3003__));
  or1   g1542(.dina(new_new_n1489__), .dinb(new_new_n1487__), .dout(new_new_n3004__));
  or1   g1543(.dina(new_new_n1490__), .dinb(new_new_n1488__), .dout(new_new_n3005__));
  and1  g1544(.dina(new_new_n3005__), .dinb(new_new_n3004__), .dout(new_new_n3006__));
  and1  g1545(.dina(new_new_n3006__), .dinb(new_new_n4580__), .dout(new_new_n3007__));
  and1  g1546(.dina(new_new_n4586__), .dinb(new_new_n1560__), .dout(new_new_n3008__));
  or1   g1547(.dina(new_new_n3007__), .dinb(new_new_n3003__), .dout(new_new_n3009__));
  or1   g1548(.dina(new_new_n3009__), .dinb(new_new_n3008__), .dout(new_new_n3010__));
  or1   g1549(.dina(new_new_n3010__), .dinb(new_new_n4600__), .dout(new_new_n3011__));
  or1   g1550(.dina(new_new_n4510__), .dinb(new_new_n4748__), .dout(new_new_n3012__));
  or1   g1551(.dina(new_new_n4614__), .dinb(new_new_n4750__), .dout(new_new_n3013__));
  or1   g1552(.dina(new_new_n4484__), .dinb(new_new_n4752__), .dout(new_new_n3014__));
  or1   g1553(.dina(new_new_n4754__), .dinb(new_new_n4489__), .dout(new_new_n3015__));
  or1   g1554(.dina(new_new_n4756__), .dinb(new_new_n4494__), .dout(new_new_n3016__));
  or1   g1555(.dina(new_new_n4758__), .dinb(new_new_n4499__), .dout(new_new_n3017__));
  or1   g1556(.dina(new_new_n4503__), .dinb(new_new_n4760__), .dout(new_new_n3018__));
  or1   g1557(.dina(new_new_n4507__), .dinb(new_new_n4762__), .dout(new_new_n3019__));
  and1  g1558(.dina(new_new_n3013__), .dinb(new_new_n3012__), .dout(new_new_n3020__));
  and1  g1559(.dina(new_new_n3020__), .dinb(new_new_n3014__), .dout(new_new_n3021__));
  and1  g1560(.dina(new_new_n3021__), .dinb(new_new_n3015__), .dout(new_new_n3022__));
  and1  g1561(.dina(new_new_n3022__), .dinb(new_new_n3016__), .dout(new_new_n3023__));
  and1  g1562(.dina(new_new_n3023__), .dinb(new_new_n3017__), .dout(new_new_n3024__));
  and1  g1563(.dina(new_new_n3024__), .dinb(new_new_n3018__), .dout(new_new_n3025__));
  and1  g1564(.dina(new_new_n3025__), .dinb(new_new_n3019__), .dout(new_new_n3026__));
  and1  g1565(.dina(new_new_n3026__), .dinb(new_new_n4518__), .dout(new_new_n3027__));
  or1   g1566(.dina(new_new_n4616__), .dinb(new_new_n4765__), .dout(new_new_n3028__));
  or1   g1567(.dina(new_new_n4531__), .dinb(new_new_n4767__), .dout(new_new_n3029__));
  or1   g1568(.dina(new_new_n4537__), .dinb(new_new_n4769__), .dout(new_new_n3030__));
  or1   g1569(.dina(new_new_n4542__), .dinb(new_new_n4771__), .dout(new_new_n3031__));
  or1   g1570(.dina(new_new_n4548__), .dinb(new_new_n4773__), .dout(new_new_n3032__));
  or1   g1571(.dina(new_new_n4775__), .dinb(new_new_n4553__), .dout(new_new_n3033__));
  or1   g1572(.dina(new_new_n4777__), .dinb(new_new_n4557__), .dout(new_new_n3034__));
  or1   g1573(.dina(new_new_n4779__), .dinb(new_new_n4521__), .dout(new_new_n3035__));
  and1  g1574(.dina(new_new_n3029__), .dinb(new_new_n3028__), .dout(new_new_n3036__));
  and1  g1575(.dina(new_new_n3036__), .dinb(new_new_n3030__), .dout(new_new_n3037__));
  and1  g1576(.dina(new_new_n3037__), .dinb(new_new_n3031__), .dout(new_new_n3038__));
  and1  g1577(.dina(new_new_n3038__), .dinb(new_new_n3032__), .dout(new_new_n3039__));
  and1  g1578(.dina(new_new_n3039__), .dinb(new_new_n3033__), .dout(new_new_n3040__));
  and1  g1579(.dina(new_new_n3040__), .dinb(new_new_n3034__), .dout(new_new_n3041__));
  and1  g1580(.dina(new_new_n3041__), .dinb(new_new_n3035__), .dout(new_new_n3042__));
  and1  g1581(.dina(new_new_n3042__), .dinb(new_new_n4565__), .dout(new_new_n3043__));
  or1   g1582(.dina(new_new_n3043__), .dinb(new_new_n3027__), .dout(new_new_n3044__));
  and1  g1583(.dina(new_new_n3044__), .dinb(new_new_n4570__), .dout(new_new_n3045__));
  or1   g1584(.dina(new_new_n1485__), .dinb(new_new_n1483__), .dout(new_new_n3046__));
  or1   g1585(.dina(new_new_n1486__), .dinb(new_new_n1484__), .dout(new_new_n3047__));
  and1  g1586(.dina(new_new_n3047__), .dinb(new_new_n3046__), .dout(new_new_n3048__));
  and1  g1587(.dina(new_new_n3048__), .dinb(new_new_n4580__), .dout(new_new_n3049__));
  and1  g1588(.dina(new_new_n4586__), .dinb(new_new_n1562__), .dout(new_new_n3050__));
  or1   g1589(.dina(new_new_n3049__), .dinb(new_new_n3045__), .dout(new_new_n3051__));
  or1   g1590(.dina(new_new_n3051__), .dinb(new_new_n3050__), .dout(new_new_n3052__));
  or1   g1591(.dina(new_new_n3052__), .dinb(new_new_n4600__), .dout(new_new_n3053__));
  or1   g1592(.dina(new_new_n4730__), .dinb(new_new_n4659__), .dout(new_new_n3054__));
  or1   g1593(.dina(new_new_n4699__), .dinb(new_new_n4476__), .dout(new_new_n3055__));
  or1   g1594(.dina(new_new_n3055__), .dinb(new_new_n4729__), .dout(new_new_n3056__));
  or1   g1595(.dina(new_new_n3056__), .dinb(new_new_n4657__), .dout(new_new_n3057__));
  and1  g1596(.dina(new_new_n3057__), .dinb(new_new_n3054__), .dout(new_new_n3058__));
  or1   g1597(.dina(new_new_n3058__), .dinb(new_new_n4592__), .dout(new_new_n3059__));
  and1  g1598(.dina(new_new_n2537__), .dinb(new_new_n4656__), .dout(new_new_n3060__));
  or1   g1599(.dina(new_new_n4475__), .dinb(new_new_n4658__), .dout(new_new_n3061__));
  or1   g1600(.dina(new_new_n3061__), .dinb(new_new_n4698__), .dout(new_new_n3062__));
  or1   g1601(.dina(new_new_n3060__), .dinb(new_new_n2865__), .dout(new_new_n3063__));
  and1  g1602(.dina(new_new_n3063__), .dinb(new_new_n3062__), .dout(new_new_n3064__));
  or1   g1603(.dina(new_new_n3064__), .dinb(new_new_n4592__), .dout(new_new_n3065__));
  or1   g1604(.dina(new_new_n4747__), .dinb(new_new_n4593__), .dout(new_new_n3066__));
  or1   g1605(.dina(new_new_n4782__), .dinb(new_new_n4783__), .dout(new_new_n3067__));
  or1   g1606(.dina(new_new_n3067__), .dinb(new_new_n4784__), .dout(new_new_n3068__));
  and1  g1607(.dina(new_new_n4785__), .dinb(new_new_n4786__), .dout(new_new_n3069__));
  or1   g1608(.dina(new_new_n4787__), .dinb(new_new_n4788__), .dout(new_new_n3070__));
  and1  g1609(.dina(new_new_n3069__), .dinb(new_new_n4789__), .dout(new_new_n3071__));
  or1   g1610(.dina(new_new_n3070__), .dinb(new_new_n4790__), .dout(new_new_n3072__));
  and1  g1611(.dina(new_new_n3071__), .dinb(new_new_n4791__), .dout(new_new_n3073__));
  or1   g1612(.dina(new_new_n3072__), .dinb(new_new_n4792__), .dout(new_new_n3074__));
  and1  g1613(.dina(new_new_n3073__), .dinb(new_new_n4793__), .dout(new_new_n3075__));
  or1   g1614(.dina(new_new_n3074__), .dinb(new_new_n4794__), .dout(new_new_n3076__));
  and1  g1615(.dina(new_new_n4787__), .dinb(new_new_n4788__), .dout(new_new_n3077__));
  or1   g1616(.dina(new_new_n4785__), .dinb(new_new_n4786__), .dout(new_new_n3078__));
  and1  g1617(.dina(new_new_n3077__), .dinb(new_new_n4790__), .dout(new_new_n3079__));
  or1   g1618(.dina(new_new_n3078__), .dinb(new_new_n4789__), .dout(new_new_n3080__));
  and1  g1619(.dina(new_new_n3079__), .dinb(new_new_n4792__), .dout(new_new_n3081__));
  or1   g1620(.dina(new_new_n3080__), .dinb(new_new_n4791__), .dout(new_new_n3082__));
  and1  g1621(.dina(new_new_n3081__), .dinb(new_new_n4794__), .dout(new_new_n3083__));
  or1   g1622(.dina(new_new_n3082__), .dinb(new_new_n4793__), .dout(new_new_n3084__));
  and1  g1623(.dina(new_new_n3084__), .dinb(new_new_n3076__), .dout(new_new_n3085__));
  or1   g1624(.dina(new_new_n3083__), .dinb(new_new_n3075__), .dout(new_new_n3086__));
  and1  g1625(.dina(new_new_n3086__), .dinb(new_new_n4666__), .dout(new_new_n3087__));
  or1   g1626(.dina(new_new_n3085__), .dinb(new_new_n4674__), .dout(new_new_n3088__));
  and1  g1627(.dina(new_new_n4795__), .dinb(new_new_n4675__), .dout(new_new_n3089__));
  or1   g1628(.dina(new_new_n2853__), .dinb(new_new_n4667__), .dout(new_new_n3090__));
  and1  g1629(.dina(new_new_n3090__), .dinb(new_new_n3088__), .dout(new_new_n3091__));
  or1   g1630(.dina(new_new_n3089__), .dinb(new_new_n3087__), .dout(new_new_n3092__));
  and1  g1631(.dina(new_new_n4796__), .dinb(new_new_n4797__), .dout(new_new_n3093__));
  and1  g1632(.dina(new_new_n3093__), .dinb(new_new_n4798__), .dout(new_new_n3094__));
  and1  g1633(.dina(new_new_n4799__), .dinb(new_new_n4800__), .dout(new_new_n3095__));
  and1  g1634(.dina(new_new_n3095__), .dinb(new_new_n4801__), .dout(new_new_n3096__));
  and1  g1635(.dina(new_new_n4802__), .dinb(new_new_n4803__), .dout(new_new_n3097__));
  and1  g1636(.dina(new_new_n3097__), .dinb(new_new_n4804__), .dout(new_new_n3098__));
  and1  g1637(.dina(new_new_n1736__), .dinb(new_new_n1734__), .dout(new_new_n3099__));
  or1   g1638(.dina(new_new_n1735__), .dinb(new_new_n1733__), .dout(new_new_n3100__));
  and1  g1639(.dina(new_new_n4805__), .dinb(new_new_n4723__), .dout(new_new_n3101__));
  and1  g1640(.dina(new_new_n1720__), .dinb(new_new_n1718__), .dout(new_new_n3102__));
  or1   g1641(.dina(new_new_n1719__), .dinb(new_new_n1717__), .dout(new_new_n3103__));
  and1  g1642(.dina(new_new_n4806__), .dinb(new_new_n2891__), .dout(new_new_n3104__));
  and1  g1643(.dina(new_new_n1704__), .dinb(new_new_n1702__), .dout(new_new_n3105__));
  or1   g1644(.dina(new_new_n1703__), .dinb(new_new_n1701__), .dout(new_new_n3106__));
  and1  g1645(.dina(new_new_n4807__), .dinb(new_new_n4726__), .dout(new_new_n3107__));
  and1  g1646(.dina(new_new_n3107__), .dinb(new_new_n1851__), .dout(new_new_n3108__));
  and1  g1647(.dina(new_new_n3108__), .dinb(new_new_n4724__), .dout(new_new_n3109__));
  or1   g1648(.dina(new_new_n3101__), .dinb(new_new_n4720__), .dout(new_new_n3110__));
  or1   g1649(.dina(new_new_n3110__), .dinb(new_new_n3104__), .dout(new_new_n3111__));
  or1   g1650(.dina(new_new_n3111__), .dinb(new_new_n3109__), .dout(new_new_n3112__));
  and1  g1651(.dina(new_new_n4667__), .dinb(new_new_n1941__), .dout(new_new_n3113__));
  or1   g1652(.dina(new_new_n4675__), .dinb(new_new_n1942__), .dout(new_new_n3114__));
  and1  g1653(.dina(new_new_n4808__), .dinb(new_new_n4809__), .dout(new_new_n3115__));
  or1   g1654(.dina(new_new_n4811__), .dinb(new_new_n4813__), .dout(new_new_n3116__));
  and1  g1655(.dina(new_new_n4811__), .dinb(new_new_n4813__), .dout(new_new_n3117__));
  or1   g1656(.dina(new_new_n4808__), .dinb(new_new_n4809__), .dout(new_new_n3118__));
  and1  g1657(.dina(new_new_n3118__), .dinb(new_new_n3116__), .dout(new_new_n3119__));
  or1   g1658(.dina(new_new_n3117__), .dinb(new_new_n3115__), .dout(new_new_n3120__));
  and1  g1659(.dina(new_new_n4669__), .dinb(new_new_n1957__), .dout(new_new_n3121__));
  or1   g1660(.dina(new_new_n4677__), .dinb(new_new_n1958__), .dout(new_new_n3122__));
  and1  g1661(.dina(new_new_n4814__), .dinb(new_new_n4815__), .dout(new_new_n3123__));
  or1   g1662(.dina(new_new_n4817__), .dinb(new_new_n4819__), .dout(new_new_n3124__));
  and1  g1663(.dina(new_new_n3124__), .dinb(new_new_n4821__), .dout(new_new_n3125__));
  or1   g1664(.dina(new_new_n4822__), .dinb(new_new_n4823__), .dout(new_new_n3126__));
  and1  g1665(.dina(new_new_n4825__), .dinb(new_new_n4826__), .dout(new_new_n3127__));
  or1   g1666(.dina(new_new_n4827__), .dinb(new_new_n4829__), .dout(new_new_n3128__));
  and1  g1667(.dina(new_new_n4827__), .dinb(new_new_n4829__), .dout(new_new_n3129__));
  or1   g1668(.dina(new_new_n4825__), .dinb(new_new_n4826__), .dout(new_new_n3130__));
  and1  g1669(.dina(new_new_n3130__), .dinb(new_new_n3128__), .dout(new_new_n3131__));
  or1   g1670(.dina(new_new_n3129__), .dinb(new_new_n3127__), .dout(new_new_n3132__));
  and1  g1671(.dina(new_new_n4830__), .dinb(new_new_n4832__), .dout(new_new_n3133__));
  or1   g1672(.dina(new_new_n4834__), .dinb(new_new_n4835__), .dout(new_new_n3134__));
  and1  g1673(.dina(new_new_n4834__), .dinb(new_new_n4835__), .dout(new_new_n3135__));
  or1   g1674(.dina(new_new_n4830__), .dinb(new_new_n4832__), .dout(new_new_n3136__));
  and1  g1675(.dina(new_new_n3136__), .dinb(new_new_n3134__), .dout(new_new_n3137__));
  or1   g1676(.dina(new_new_n3135__), .dinb(new_new_n3133__), .dout(new_new_n3138__));
  and1  g1677(.dina(new_new_n4837__), .dinb(new_new_n4840__), .dout(new_new_n3139__));
  or1   g1678(.dina(new_new_n3139__), .dinb(new_new_n4843__), .dout(new_new_n3140__));
  and1  g1679(.dina(new_new_n4805__), .dinb(new_new_n4663__), .dout(new_new_n3141__));
  or1   g1680(.dina(new_new_n3099__), .dinb(new_new_n4661__), .dout(new_new_n3142__));
  and1  g1681(.dina(new_new_n4844__), .dinb(new_new_n4845__), .dout(new_new_n3143__));
  or1   g1682(.dina(new_new_n4847__), .dinb(new_new_n4849__), .dout(new_new_n3144__));
  and1  g1683(.dina(new_new_n4847__), .dinb(new_new_n4849__), .dout(new_new_n3145__));
  or1   g1684(.dina(new_new_n4844__), .dinb(new_new_n4845__), .dout(new_new_n3146__));
  and1  g1685(.dina(new_new_n3146__), .dinb(new_new_n3144__), .dout(new_new_n3147__));
  or1   g1686(.dina(new_new_n3145__), .dinb(new_new_n3143__), .dout(new_new_n3148__));
  and1  g1687(.dina(new_new_n4806__), .dinb(new_new_n4669__), .dout(new_new_n3149__));
  or1   g1688(.dina(new_new_n3102__), .dinb(new_new_n4677__), .dout(new_new_n3150__));
  and1  g1689(.dina(new_new_n4850__), .dinb(new_new_n4852__), .dout(new_new_n3151__));
  or1   g1690(.dina(new_new_n4853__), .dinb(new_new_n4855__), .dout(new_new_n3152__));
  and1  g1691(.dina(new_new_n4857__), .dinb(new_new_n4858__), .dout(new_new_n3153__));
  or1   g1692(.dina(new_new_n4859__), .dinb(new_new_n4860__), .dout(new_new_n3154__));
  and1  g1693(.dina(new_new_n4859__), .dinb(new_new_n4860__), .dout(new_new_n3155__));
  or1   g1694(.dina(new_new_n4857__), .dinb(new_new_n4858__), .dout(new_new_n3156__));
  and1  g1695(.dina(new_new_n3156__), .dinb(new_new_n3154__), .dout(new_new_n3157__));
  or1   g1696(.dina(new_new_n3155__), .dinb(new_new_n3153__), .dout(new_new_n3158__));
  and1  g1697(.dina(new_new_n4807__), .dinb(new_new_n4670__), .dout(new_new_n3159__));
  or1   g1698(.dina(new_new_n3105__), .dinb(new_new_n4678__), .dout(new_new_n3160__));
  and1  g1699(.dina(new_new_n4862__), .dinb(new_new_n4852__), .dout(new_new_n3161__));
  or1   g1700(.dina(new_new_n4866__), .dinb(new_new_n4855__), .dout(new_new_n3162__));
  and1  g1701(.dina(new_new_n4869__), .dinb(new_new_n4871__), .dout(new_new_n3163__));
  or1   g1702(.dina(new_new_n4872__), .dinb(new_new_n4874__), .dout(new_new_n3164__));
  and1  g1703(.dina(new_new_n4869__), .dinb(new_new_n4876__), .dout(new_new_n3165__));
  or1   g1704(.dina(new_new_n4872__), .dinb(new_new_n4880__), .dout(new_new_n3166__));
  and1  g1705(.dina(new_new_n3165__), .dinb(new_new_n4840__), .dout(new_new_n3167__));
  or1   g1706(.dina(new_new_n3166__), .dinb(new_new_n4884__), .dout(new_new_n3168__));
  and1  g1707(.dina(new_new_n3152__), .dinb(new_new_n3142__), .dout(new_new_n3169__));
  or1   g1708(.dina(new_new_n3151__), .dinb(new_new_n3141__), .dout(new_new_n3170__));
  and1  g1709(.dina(new_new_n3169__), .dinb(new_new_n3164__), .dout(new_new_n3171__));
  or1   g1710(.dina(new_new_n3170__), .dinb(new_new_n3163__), .dout(new_new_n3172__));
  and1  g1711(.dina(new_new_n3171__), .dinb(new_new_n3168__), .dout(new_new_n3173__));
  or1   g1712(.dina(new_new_n3172__), .dinb(new_new_n3167__), .dout(new_new_n3174__));
  and1  g1713(.dina(new_new_n4886__), .dinb(new_new_n4888__), .dout(new_new_n3175__));
  or1   g1714(.dina(new_new_n4889__), .dinb(new_new_n4891__), .dout(new_new_n3176__));
  or1   g1715(.dina(new_new_n4889__), .dinb(new_new_n4893__), .dout(new_new_n3177__));
  and1  g1716(.dina(new_new_n4894__), .dinb(new_new_n1739__), .dout(new_new_n3178__));
  or1   g1717(.dina(new_new_n4895__), .dinb(new_new_n1740__), .dout(new_new_n3179__));
  and1  g1718(.dina(new_new_n4896__), .dinb(new_new_n4693__), .dout(new_new_n3180__));
  or1   g1719(.dina(new_new_n4898__), .dinb(new_new_n4690__), .dout(new_new_n3181__));
  and1  g1720(.dina(new_new_n4898__), .dinb(new_new_n4691__), .dout(new_new_n3182__));
  or1   g1721(.dina(new_new_n4896__), .dinb(new_new_n4692__), .dout(new_new_n3183__));
  and1  g1722(.dina(new_new_n3183__), .dinb(new_new_n3181__), .dout(new_new_n3184__));
  or1   g1723(.dina(new_new_n3182__), .dinb(new_new_n3180__), .dout(new_new_n3185__));
  and1  g1724(.dina(new_new_n4900__), .dinb(new_new_n4904__), .dout(new_new_n3186__));
  or1   g1725(.dina(new_new_n2204__), .dinb(new_new_n4911__), .dout(new_new_n3187__));
  and1  g1726(.dina(new_new_n4915__), .dinb(new_new_n2184__), .dout(new_new_n3188__));
  or1   g1727(.dina(new_new_n4917__), .dinb(new_new_n2183__), .dout(new_new_n3189__));
  and1  g1728(.dina(new_new_n4918__), .dinb(new_new_n4911__), .dout(new_new_n3190__));
  or1   g1729(.dina(new_new_n4920__), .dinb(new_new_n4904__), .dout(new_new_n3191__));
  and1  g1730(.dina(new_new_n4924__), .dinb(new_new_n4930__), .dout(new_new_n3192__));
  or1   g1731(.dina(new_new_n4934__), .dinb(new_new_n4939__), .dout(new_new_n3193__));
  and1  g1732(.dina(new_new_n3192__), .dinb(new_new_n4940__), .dout(new_new_n3194__));
  or1   g1733(.dina(new_new_n3193__), .dinb(new_new_n4941__), .dout(new_new_n3195__));
  and1  g1734(.dina(new_new_n4924__), .dinb(new_new_n4942__), .dout(new_new_n3196__));
  or1   g1735(.dina(new_new_n4934__), .dinb(new_new_n4943__), .dout(new_new_n3197__));
  and1  g1736(.dina(new_new_n4944__), .dinb(new_new_n4941__), .dout(new_new_n3198__));
  or1   g1737(.dina(new_new_n4945__), .dinb(new_new_n4940__), .dout(new_new_n3199__));
  and1  g1738(.dina(new_new_n4948__), .dinb(new_new_n4953__), .dout(new_new_n3200__));
  or1   g1739(.dina(new_new_n4960__), .dinb(new_new_n4964__), .dout(new_new_n3201__));
  and1  g1740(.dina(new_new_n4968__), .dinb(new_new_n4972__), .dout(new_new_n3202__));
  or1   g1741(.dina(new_new_n4978__), .dinb(new_new_n4981__), .dout(new_new_n3203__));
  and1  g1742(.dina(new_new_n4964__), .dinb(new_new_n4981__), .dout(new_new_n3204__));
  or1   g1743(.dina(new_new_n4953__), .dinb(new_new_n4972__), .dout(new_new_n3205__));
  and1  g1744(.dina(new_new_n4986__), .dinb(new_new_n4991__), .dout(new_new_n3206__));
  or1   g1745(.dina(new_new_n4995__), .dinb(new_new_n4998__), .dout(new_new_n3207__));
  and1  g1746(.dina(new_new_n3203__), .dinb(new_new_n3201__), .dout(new_new_n3208__));
  or1   g1747(.dina(new_new_n3202__), .dinb(new_new_n3200__), .dout(new_new_n3209__));
  and1  g1748(.dina(new_new_n3208__), .dinb(new_new_n3207__), .dout(new_new_n3210__));
  or1   g1749(.dina(new_new_n3209__), .dinb(new_new_n3206__), .dout(new_new_n3211__));
  and1  g1750(.dina(new_new_n3211__), .dinb(new_new_n4923__), .dout(new_new_n3212__));
  or1   g1751(.dina(new_new_n3210__), .dinb(new_new_n4935__), .dout(new_new_n3213__));
  and1  g1752(.dina(new_new_n3199__), .dinb(new_new_n3195__), .dout(new_new_n3214__));
  or1   g1753(.dina(new_new_n3198__), .dinb(new_new_n3194__), .dout(new_new_n3215__));
  and1  g1754(.dina(new_new_n3214__), .dinb(new_new_n3213__), .dout(new_new_n3216__));
  or1   g1755(.dina(new_new_n3215__), .dinb(new_new_n3212__), .dout(new_new_n3217__));
  and1  g1756(.dina(new_new_n4999__), .dinb(new_new_n4918__), .dout(new_new_n3218__));
  or1   g1757(.dina(new_new_n5000__), .dinb(new_new_n4920__), .dout(new_new_n3219__));
  and1  g1758(.dina(new_new_n3218__), .dinb(new_new_n2162__), .dout(new_new_n3220__));
  or1   g1759(.dina(new_new_n3219__), .dinb(new_new_n5001__), .dout(new_new_n3221__));
  and1  g1760(.dina(new_new_n4925__), .dinb(new_new_n5003__), .dout(new_new_n3222__));
  or1   g1761(.dina(new_new_n4935__), .dinb(new_new_n5005__), .dout(new_new_n3223__));
  and1  g1762(.dina(new_new_n3222__), .dinb(new_new_n5007__), .dout(new_new_n3224__));
  or1   g1763(.dina(new_new_n3223__), .dinb(new_new_n5010__), .dout(new_new_n3225__));
  and1  g1764(.dina(new_new_n5010__), .dinb(new_new_n4944__), .dout(new_new_n3226__));
  or1   g1765(.dina(new_new_n5007__), .dinb(new_new_n4945__), .dout(new_new_n3227__));
  and1  g1766(.dina(new_new_n5012__), .dinb(new_new_n4954__), .dout(new_new_n3228__));
  or1   g1767(.dina(new_new_n5013__), .dinb(new_new_n4965__), .dout(new_new_n3229__));
  and1  g1768(.dina(new_new_n4991__), .dinb(new_new_n4973__), .dout(new_new_n3230__));
  or1   g1769(.dina(new_new_n4998__), .dinb(new_new_n4982__), .dout(new_new_n3231__));
  and1  g1770(.dina(new_new_n4986__), .dinb(new_new_n4930__), .dout(new_new_n3232__));
  or1   g1771(.dina(new_new_n4995__), .dinb(new_new_n4939__), .dout(new_new_n3233__));
  and1  g1772(.dina(new_new_n3231__), .dinb(new_new_n3229__), .dout(new_new_n3234__));
  or1   g1773(.dina(new_new_n3230__), .dinb(new_new_n3228__), .dout(new_new_n3235__));
  and1  g1774(.dina(new_new_n3234__), .dinb(new_new_n3233__), .dout(new_new_n3236__));
  or1   g1775(.dina(new_new_n3235__), .dinb(new_new_n3232__), .dout(new_new_n3237__));
  and1  g1776(.dina(new_new_n3237__), .dinb(new_new_n4925__), .dout(new_new_n3238__));
  or1   g1777(.dina(new_new_n3236__), .dinb(new_new_n4937__), .dout(new_new_n3239__));
  and1  g1778(.dina(new_new_n5014__), .dinb(new_new_n3225__), .dout(new_new_n3240__));
  or1   g1779(.dina(new_new_n5016__), .dinb(new_new_n3224__), .dout(new_new_n3241__));
  and1  g1780(.dina(new_new_n3240__), .dinb(new_new_n3239__), .dout(new_new_n3242__));
  or1   g1781(.dina(new_new_n3241__), .dinb(new_new_n3238__), .dout(new_new_n3243__));
  and1  g1782(.dina(new_new_n4927__), .dinb(new_new_n5018__), .dout(new_new_n3244__));
  or1   g1783(.dina(new_new_n4937__), .dinb(new_new_n1296__), .dout(new_new_n3245__));
  and1  g1784(.dina(new_new_n3244__), .dinb(new_new_n5008__), .dout(new_new_n3246__));
  or1   g1785(.dina(new_new_n3245__), .dinb(new_new_n5009__), .dout(new_new_n3247__));
  and1  g1786(.dina(new_new_n5019__), .dinb(new_new_n4954__), .dout(new_new_n3248__));
  or1   g1787(.dina(new_new_n2252__), .dinb(new_new_n4965__), .dout(new_new_n3249__));
  and1  g1788(.dina(new_new_n4931__), .dinb(new_new_n4973__), .dout(new_new_n3250__));
  or1   g1789(.dina(new_new_n4938__), .dinb(new_new_n4982__), .dout(new_new_n3251__));
  and1  g1790(.dina(new_new_n4987__), .dinb(new_new_n5003__), .dout(new_new_n3252__));
  or1   g1791(.dina(new_new_n4994__), .dinb(new_new_n5005__), .dout(new_new_n3253__));
  and1  g1792(.dina(new_new_n3251__), .dinb(new_new_n3249__), .dout(new_new_n3254__));
  or1   g1793(.dina(new_new_n3250__), .dinb(new_new_n3248__), .dout(new_new_n3255__));
  and1  g1794(.dina(new_new_n3254__), .dinb(new_new_n3253__), .dout(new_new_n3256__));
  or1   g1795(.dina(new_new_n3255__), .dinb(new_new_n3252__), .dout(new_new_n3257__));
  and1  g1796(.dina(new_new_n3257__), .dinb(new_new_n4927__), .dout(new_new_n3258__));
  or1   g1797(.dina(new_new_n3256__), .dinb(new_new_n4936__), .dout(new_new_n3259__));
  and1  g1798(.dina(new_new_n3247__), .dinb(new_new_n5014__), .dout(new_new_n3260__));
  or1   g1799(.dina(new_new_n3246__), .dinb(new_new_n5016__), .dout(new_new_n3261__));
  and1  g1800(.dina(new_new_n3260__), .dinb(new_new_n3259__), .dout(new_new_n3262__));
  or1   g1801(.dina(new_new_n3261__), .dinb(new_new_n3258__), .dout(new_new_n3263__));
  and1  g1802(.dina(new_new_n5023__), .dinb(new_new_n5030__), .dout(new_new_n3264__));
  or1   g1803(.dina(new_new_n5036__), .dinb(new_new_n5043__), .dout(new_new_n3265__));
  and1  g1804(.dina(new_new_n5047__), .dinb(new_new_n5053__), .dout(new_new_n3266__));
  or1   g1805(.dina(new_new_n5060__), .dinb(new_new_n5067__), .dout(new_new_n3267__));
  and1  g1806(.dina(new_new_n5036__), .dinb(new_new_n5067__), .dout(new_new_n3268__));
  or1   g1807(.dina(new_new_n5023__), .dinb(new_new_n5053__), .dout(new_new_n3269__));
  and1  g1808(.dina(new_new_n5074__), .dinb(new_new_n5080__), .dout(new_new_n3270__));
  or1   g1809(.dina(new_new_n5084__), .dinb(new_new_n5090__), .dout(new_new_n3271__));
  and1  g1810(.dina(new_new_n3267__), .dinb(new_new_n3265__), .dout(new_new_n3272__));
  or1   g1811(.dina(new_new_n3266__), .dinb(new_new_n3264__), .dout(new_new_n3273__));
  and1  g1812(.dina(new_new_n3272__), .dinb(new_new_n3271__), .dout(new_new_n3274__));
  or1   g1813(.dina(new_new_n3273__), .dinb(new_new_n3270__), .dout(new_new_n3275__));
  and1  g1814(.dina(new_new_n5095__), .dinb(new_new_n4905__), .dout(new_new_n3276__));
  or1   g1815(.dina(new_new_n5097__), .dinb(new_new_n4912__), .dout(new_new_n3277__));
  and1  g1816(.dina(new_new_n3276__), .dinb(new_new_n5099__), .dout(new_new_n3278__));
  or1   g1817(.dina(new_new_n3277__), .dinb(new_new_n5100__), .dout(new_new_n3279__));
  and1  g1818(.dina(new_new_n3279__), .dinb(new_new_n4917__), .dout(new_new_n3280__));
  or1   g1819(.dina(new_new_n3278__), .dinb(new_new_n4915__), .dout(new_new_n3281__));
  and1  g1820(.dina(new_new_n5104__), .dinb(new_new_n3275__), .dout(new_new_n3282__));
  or1   g1821(.dina(new_new_n5111__), .dinb(new_new_n3274__), .dout(new_new_n3283__));
  and1  g1822(.dina(new_new_n2275__), .dinb(new_new_n4912__), .dout(new_new_n3284__));
  or1   g1823(.dina(new_new_n2276__), .dinb(new_new_n4905__), .dout(new_new_n3285__));
  and1  g1824(.dina(new_new_n5119__), .dinb(new_new_n5043__), .dout(new_new_n3286__));
  or1   g1825(.dina(new_new_n5126__), .dinb(new_new_n5030__), .dout(new_new_n3287__));
  and1  g1826(.dina(new_new_n5095__), .dinb(new_new_n4913__), .dout(new_new_n3288__));
  or1   g1827(.dina(new_new_n5097__), .dinb(new_new_n4907__), .dout(new_new_n3289__));
  and1  g1828(.dina(new_new_n5126__), .dinb(new_new_n5111__), .dout(new_new_n3290__));
  or1   g1829(.dina(new_new_n5119__), .dinb(new_new_n5104__), .dout(new_new_n3291__));
  and1  g1830(.dina(new_new_n5132__), .dinb(new_new_n5031__), .dout(new_new_n3292__));
  or1   g1831(.dina(new_new_n5135__), .dinb(new_new_n5042__), .dout(new_new_n3293__));
  and1  g1832(.dina(new_new_n3292__), .dinb(new_new_n5138__), .dout(new_new_n3294__));
  or1   g1833(.dina(new_new_n3293__), .dinb(new_new_n5145__), .dout(new_new_n3295__));
  and1  g1834(.dina(new_new_n3287__), .dinb(new_new_n3283__), .dout(new_new_n3296__));
  or1   g1835(.dina(new_new_n3286__), .dinb(new_new_n3282__), .dout(new_new_n3297__));
  and1  g1836(.dina(new_new_n3296__), .dinb(new_new_n3295__), .dout(new_new_n3298__));
  or1   g1837(.dina(new_new_n3297__), .dinb(new_new_n3294__), .dout(new_new_n3299__));
  and1  g1838(.dina(new_new_n4914__), .dinb(new_new_n2262__), .dout(new_new_n3300__));
  or1   g1839(.dina(new_new_n4916__), .dinb(new_new_n2261__), .dout(new_new_n3301__));
  and1  g1840(.dina(new_new_n4999__), .dinb(new_new_n2253__), .dout(new_new_n3302__));
  or1   g1841(.dina(new_new_n5000__), .dinb(new_new_n2254__), .dout(new_new_n3303__));
  and1  g1842(.dina(new_new_n5152__), .dinb(new_new_n4992__), .dout(new_new_n3304__));
  or1   g1843(.dina(new_new_n5159__), .dinb(new_new_n4997__), .dout(new_new_n3305__));
  and1  g1844(.dina(new_new_n3304__), .dinb(new_new_n5165__), .dout(new_new_n3306__));
  or1   g1845(.dina(new_new_n3305__), .dinb(new_new_n5168__), .dout(new_new_n3307__));
  and1  g1846(.dina(new_new_n5152__), .dinb(new_new_n4942__), .dout(new_new_n3308__));
  or1   g1847(.dina(new_new_n5159__), .dinb(new_new_n4943__), .dout(new_new_n3309__));
  and1  g1848(.dina(new_new_n3308__), .dinb(new_new_n5168__), .dout(new_new_n3310__));
  or1   g1849(.dina(new_new_n3309__), .dinb(new_new_n5165__), .dout(new_new_n3311__));
  and1  g1850(.dina(new_new_n2284__), .dinb(new_new_n5172__), .dout(new_new_n3312__));
  or1   g1851(.dina(new_new_n2283__), .dinb(new_new_n5179__), .dout(new_new_n3313__));
  and1  g1852(.dina(new_new_n5183__), .dinb(new_new_n2264__), .dout(new_new_n3314__));
  or1   g1853(.dina(new_new_n5186__), .dinb(new_new_n2263__), .dout(new_new_n3315__));
  and1  g1854(.dina(new_new_n4968__), .dinb(new_new_n2265__), .dout(new_new_n3316__));
  or1   g1855(.dina(new_new_n4978__), .dinb(new_new_n2266__), .dout(new_new_n3317__));
  and1  g1856(.dina(new_new_n3315__), .dinb(new_new_n3313__), .dout(new_new_n3318__));
  or1   g1857(.dina(new_new_n3314__), .dinb(new_new_n3312__), .dout(new_new_n3319__));
  and1  g1858(.dina(new_new_n3318__), .dinb(new_new_n3317__), .dout(new_new_n3320__));
  or1   g1859(.dina(new_new_n3319__), .dinb(new_new_n3316__), .dout(new_new_n3321__));
  and1  g1860(.dina(new_new_n3321__), .dinb(new_new_n5151__), .dout(new_new_n3322__));
  or1   g1861(.dina(new_new_n3320__), .dinb(new_new_n5160__), .dout(new_new_n3323__));
  and1  g1862(.dina(new_new_n5188__), .dinb(new_new_n3307__), .dout(new_new_n3324__));
  or1   g1863(.dina(new_new_n5190__), .dinb(new_new_n3306__), .dout(new_new_n3325__));
  and1  g1864(.dina(new_new_n3324__), .dinb(new_new_n3323__), .dout(new_new_n3326__));
  or1   g1865(.dina(new_new_n3325__), .dinb(new_new_n3322__), .dout(new_new_n3327__));
  or1   g1866(.dina(new_new_n5194__), .dinb(new_new_n5198__), .dout(new_new_n3328__));
  or1   g1867(.dina(new_new_n3328__), .dinb(new_new_n5201__), .dout(new_new_n3329__));
  or1   g1868(.dina(new_new_n5194__), .dinb(new_new_n5204__), .dout(new_new_n3330__));
  or1   g1869(.dina(new_new_n3330__), .dinb(new_new_n5201__), .dout(new_new_n3331__));
  or1   g1870(.dina(new_new_n1617__), .dinb(new_new_n1615__), .dout(new_new_n3332__));
  or1   g1871(.dina(new_new_n3332__), .dinb(new_new_n1611__), .dout(new_new_n3333__));
  or1   g1872(.dina(new_new_n3185__), .dinb(new_new_n4819__), .dout(new_new_n3334__));
  and1  g1873(.dina(new_new_n5208__), .dinb(new_new_n4837__), .dout(new_new_n3335__));
  or1   g1874(.dina(new_new_n4900__), .dinb(new_new_n4907__), .dout(new_new_n3336__));
  or1   g1875(.dina(new_new_n3336__), .dinb(new_new_n5094__), .dout(new_new_n3337__));
  and1  g1876(.dina(new_new_n5022__), .dinb(new_new_n5211__), .dout(new_new_n3338__));
  or1   g1877(.dina(new_new_n5037__), .dinb(new_new_n5215__), .dout(new_new_n3339__));
  and1  g1878(.dina(new_new_n5052__), .dinb(new_new_n5031__), .dout(new_new_n3340__));
  or1   g1879(.dina(new_new_n5068__), .dinb(new_new_n5044__), .dout(new_new_n3341__));
  and1  g1880(.dina(new_new_n5074__), .dinb(new_new_n5222__), .dout(new_new_n3342__));
  or1   g1881(.dina(new_new_n5084__), .dinb(new_new_n5224__), .dout(new_new_n3343__));
  and1  g1882(.dina(new_new_n3341__), .dinb(new_new_n3339__), .dout(new_new_n3344__));
  or1   g1883(.dina(new_new_n3340__), .dinb(new_new_n3338__), .dout(new_new_n3345__));
  and1  g1884(.dina(new_new_n3344__), .dinb(new_new_n3343__), .dout(new_new_n3346__));
  or1   g1885(.dina(new_new_n3345__), .dinb(new_new_n3342__), .dout(new_new_n3347__));
  and1  g1886(.dina(new_new_n3347__), .dinb(new_new_n5103__), .dout(new_new_n3348__));
  or1   g1887(.dina(new_new_n3346__), .dinb(new_new_n5112__), .dout(new_new_n3349__));
  and1  g1888(.dina(new_new_n5118__), .dinb(new_new_n5211__), .dout(new_new_n3350__));
  or1   g1889(.dina(new_new_n5127__), .dinb(new_new_n5215__), .dout(new_new_n3351__));
  and1  g1890(.dina(new_new_n5132__), .dinb(new_new_n5216__), .dout(new_new_n3352__));
  or1   g1891(.dina(new_new_n5135__), .dinb(new_new_n5210__), .dout(new_new_n3353__));
  and1  g1892(.dina(new_new_n3352__), .dinb(new_new_n5138__), .dout(new_new_n3354__));
  or1   g1893(.dina(new_new_n3353__), .dinb(new_new_n5145__), .dout(new_new_n3355__));
  and1  g1894(.dina(new_new_n3351__), .dinb(new_new_n3349__), .dout(new_new_n3356__));
  or1   g1895(.dina(new_new_n3350__), .dinb(new_new_n3348__), .dout(new_new_n3357__));
  and1  g1896(.dina(new_new_n3356__), .dinb(new_new_n3355__), .dout(new_new_n3358__));
  or1   g1897(.dina(new_new_n3357__), .dinb(new_new_n3354__), .dout(new_new_n3359__));
  and1  g1898(.dina(new_new_n5153__), .dinb(new_new_n4969__), .dout(new_new_n3360__));
  or1   g1899(.dina(new_new_n5160__), .dinb(new_new_n4977__), .dout(new_new_n3361__));
  and1  g1900(.dina(new_new_n3360__), .dinb(new_new_n5164__), .dout(new_new_n3362__));
  or1   g1901(.dina(new_new_n3361__), .dinb(new_new_n5169__), .dout(new_new_n3363__));
  and1  g1902(.dina(new_new_n4956__), .dinb(new_new_n5227__), .dout(new_new_n3364__));
  or1   g1903(.dina(new_new_n4966__), .dinb(new_new_n5234__), .dout(new_new_n3365__));
  and1  g1904(.dina(new_new_n5238__), .dinb(new_new_n4975__), .dout(new_new_n3366__));
  or1   g1905(.dina(new_new_n5240__), .dinb(new_new_n4983__), .dout(new_new_n3367__));
  and1  g1906(.dina(new_new_n4987__), .dinb(new_new_n5183__), .dout(new_new_n3368__));
  or1   g1907(.dina(new_new_n4996__), .dinb(new_new_n5186__), .dout(new_new_n3369__));
  and1  g1908(.dina(new_new_n3367__), .dinb(new_new_n3365__), .dout(new_new_n3370__));
  or1   g1909(.dina(new_new_n3366__), .dinb(new_new_n3364__), .dout(new_new_n3371__));
  and1  g1910(.dina(new_new_n3370__), .dinb(new_new_n3369__), .dout(new_new_n3372__));
  or1   g1911(.dina(new_new_n3371__), .dinb(new_new_n3368__), .dout(new_new_n3373__));
  and1  g1912(.dina(new_new_n3373__), .dinb(new_new_n5153__), .dout(new_new_n3374__));
  or1   g1913(.dina(new_new_n3372__), .dinb(new_new_n5162__), .dout(new_new_n3375__));
  and1  g1914(.dina(new_new_n3363__), .dinb(new_new_n5188__), .dout(new_new_n3376__));
  or1   g1915(.dina(new_new_n3362__), .dinb(new_new_n5190__), .dout(new_new_n3377__));
  and1  g1916(.dina(new_new_n3376__), .dinb(new_new_n3375__), .dout(new_new_n3378__));
  or1   g1917(.dina(new_new_n3377__), .dinb(new_new_n3374__), .dout(new_new_n3379__));
  or1   g1918(.dina(new_new_n5243__), .dinb(new_new_n5198__), .dout(new_new_n3380__));
  or1   g1919(.dina(new_new_n3380__), .dinb(new_new_n5245__), .dout(new_new_n3381__));
  or1   g1920(.dina(new_new_n5243__), .dinb(new_new_n5204__), .dout(new_new_n3382__));
  or1   g1921(.dina(new_new_n3382__), .dinb(new_new_n5245__), .dout(new_new_n3383__));
  and1  g1922(.dina(new_new_n2281__), .dinb(new_new_n2233__), .dout(new_new_n3384__));
  or1   g1923(.dina(new_new_n2282__), .dinb(new_new_n2234__), .dout(new_new_n3385__));
  and1  g1924(.dina(new_new_n2288__), .dinb(new_new_n2228__), .dout(new_new_n3386__));
  or1   g1925(.dina(new_new_n2287__), .dinb(new_new_n2227__), .dout(new_new_n3387__));
  and1  g1926(.dina(new_new_n3387__), .dinb(new_new_n3385__), .dout(new_new_n3388__));
  or1   g1927(.dina(new_new_n3386__), .dinb(new_new_n3384__), .dout(new_new_n3389__));
  and1  g1928(.dina(new_new_n3388__), .dinb(new_new_n5024__), .dout(new_new_n3390__));
  or1   g1929(.dina(new_new_n3389__), .dinb(new_new_n5037__), .dout(new_new_n3391__));
  and1  g1930(.dina(new_new_n5054__), .dinb(new_new_n5172__), .dout(new_new_n3392__));
  or1   g1931(.dina(new_new_n5068__), .dinb(new_new_n5179__), .dout(new_new_n3393__));
  and1  g1932(.dina(new_new_n5075__), .dinb(new_new_n5033__), .dout(new_new_n3394__));
  or1   g1933(.dina(new_new_n5085__), .dinb(new_new_n5044__), .dout(new_new_n3395__));
  and1  g1934(.dina(new_new_n3393__), .dinb(new_new_n3391__), .dout(new_new_n3396__));
  or1   g1935(.dina(new_new_n3392__), .dinb(new_new_n3390__), .dout(new_new_n3397__));
  and1  g1936(.dina(new_new_n3396__), .dinb(new_new_n3395__), .dout(new_new_n3398__));
  or1   g1937(.dina(new_new_n3397__), .dinb(new_new_n3394__), .dout(new_new_n3399__));
  and1  g1938(.dina(new_new_n3399__), .dinb(new_new_n5105__), .dout(new_new_n3400__));
  or1   g1939(.dina(new_new_n3398__), .dinb(new_new_n5112__), .dout(new_new_n3401__));
  and1  g1940(.dina(new_new_n5120__), .dinb(new_new_n5234__), .dout(new_new_n3402__));
  or1   g1941(.dina(new_new_n5127__), .dinb(new_new_n5227__), .dout(new_new_n3403__));
  and1  g1942(.dina(new_new_n4913__), .dinb(new_new_n5099__), .dout(new_new_n3404__));
  or1   g1943(.dina(new_new_n4908__), .dinb(new_new_n5100__), .dout(new_new_n3405__));
  and1  g1944(.dina(new_new_n5247__), .dinb(new_new_n5228__), .dout(new_new_n3406__));
  or1   g1945(.dina(new_new_n5250__), .dinb(new_new_n5235__), .dout(new_new_n3407__));
  and1  g1946(.dina(new_new_n3406__), .dinb(new_new_n5139__), .dout(new_new_n3408__));
  or1   g1947(.dina(new_new_n3407__), .dinb(new_new_n5146__), .dout(new_new_n3409__));
  and1  g1948(.dina(new_new_n3403__), .dinb(new_new_n3401__), .dout(new_new_n3410__));
  or1   g1949(.dina(new_new_n3402__), .dinb(new_new_n3400__), .dout(new_new_n3411__));
  and1  g1950(.dina(new_new_n3410__), .dinb(new_new_n3409__), .dout(new_new_n3412__));
  or1   g1951(.dina(new_new_n3411__), .dinb(new_new_n3408__), .dout(new_new_n3413__));
  and1  g1952(.dina(new_new_n5047__), .dinb(new_new_n5235__), .dout(new_new_n3414__));
  or1   g1953(.dina(new_new_n5060__), .dinb(new_new_n5228__), .dout(new_new_n3415__));
  and1  g1954(.dina(new_new_n3414__), .dinb(new_new_n5180__), .dout(new_new_n3416__));
  or1   g1955(.dina(new_new_n3415__), .dinb(new_new_n5173__), .dout(new_new_n3417__));
  and1  g1956(.dina(new_new_n3417__), .dinb(new_new_n5024__), .dout(new_new_n3418__));
  or1   g1957(.dina(new_new_n3416__), .dinb(new_new_n5039__), .dout(new_new_n3419__));
  and1  g1958(.dina(new_new_n5054__), .dinb(new_new_n5236__), .dout(new_new_n3420__));
  or1   g1959(.dina(new_new_n5070__), .dinb(new_new_n5230__), .dout(new_new_n3421__));
  and1  g1960(.dina(new_new_n5075__), .dinb(new_new_n5212__), .dout(new_new_n3422__));
  or1   g1961(.dina(new_new_n5085__), .dinb(new_new_n5216__), .dout(new_new_n3423__));
  and1  g1962(.dina(new_new_n3421__), .dinb(new_new_n3419__), .dout(new_new_n3424__));
  or1   g1963(.dina(new_new_n3420__), .dinb(new_new_n3418__), .dout(new_new_n3425__));
  and1  g1964(.dina(new_new_n3424__), .dinb(new_new_n3423__), .dout(new_new_n3426__));
  or1   g1965(.dina(new_new_n3425__), .dinb(new_new_n3422__), .dout(new_new_n3427__));
  and1  g1966(.dina(new_new_n3427__), .dinb(new_new_n5105__), .dout(new_new_n3428__));
  or1   g1967(.dina(new_new_n3426__), .dinb(new_new_n5114__), .dout(new_new_n3429__));
  and1  g1968(.dina(new_new_n5120__), .dinb(new_new_n5048__), .dout(new_new_n3430__));
  or1   g1969(.dina(new_new_n5129__), .dinb(new_new_n5061__), .dout(new_new_n3431__));
  and1  g1970(.dina(new_new_n5247__), .dinb(new_new_n5061__), .dout(new_new_n3432__));
  or1   g1971(.dina(new_new_n5250__), .dinb(new_new_n5048__), .dout(new_new_n3433__));
  and1  g1972(.dina(new_new_n3432__), .dinb(new_new_n5139__), .dout(new_new_n3434__));
  or1   g1973(.dina(new_new_n3433__), .dinb(new_new_n5146__), .dout(new_new_n3435__));
  and1  g1974(.dina(new_new_n3431__), .dinb(new_new_n3429__), .dout(new_new_n3436__));
  or1   g1975(.dina(new_new_n3430__), .dinb(new_new_n3428__), .dout(new_new_n3437__));
  and1  g1976(.dina(new_new_n3436__), .dinb(new_new_n3435__), .dout(new_new_n3438__));
  or1   g1977(.dina(new_new_n3437__), .dinb(new_new_n3434__), .dout(new_new_n3439__));
  and1  g1978(.dina(new_new_n4928__), .dinb(new_new_n5252__), .dout(new_new_n3440__));
  and1  g1979(.dina(new_new_n3440__), .dinb(new_new_n5008__), .dout(new_new_n3441__));
  and1  g1980(.dina(new_new_n4956__), .dinb(new_new_n5253__), .dout(new_new_n3442__));
  and1  g1981(.dina(new_new_n5004__), .dinb(new_new_n4975__), .dout(new_new_n3443__));
  and1  g1982(.dina(new_new_n4989__), .dinb(new_new_n5018__), .dout(new_new_n3444__));
  or1   g1983(.dina(new_new_n3443__), .dinb(new_new_n3442__), .dout(new_new_n3445__));
  or1   g1984(.dina(new_new_n3445__), .dinb(new_new_n3444__), .dout(new_new_n3446__));
  and1  g1985(.dina(new_new_n3446__), .dinb(new_new_n4928__), .dout(new_new_n3447__));
  or1   g1986(.dina(new_new_n3441__), .dinb(new_new_n5015__), .dout(new_new_n3448__));
  or1   g1987(.dina(new_new_n3448__), .dinb(new_new_n3447__), .dout(new_new_n3449__));
  and1  g1988(.dina(new_new_n2279__), .dinb(new_new_n2231__), .dout(new_new_n3450__));
  or1   g1989(.dina(new_new_n2280__), .dinb(new_new_n2232__), .dout(new_new_n3451__));
  and1  g1990(.dina(new_new_n2286__), .dinb(new_new_n2226__), .dout(new_new_n3452__));
  or1   g1991(.dina(new_new_n2285__), .dinb(new_new_n2225__), .dout(new_new_n3453__));
  and1  g1992(.dina(new_new_n3453__), .dinb(new_new_n3451__), .dout(new_new_n3454__));
  or1   g1993(.dina(new_new_n3452__), .dinb(new_new_n3450__), .dout(new_new_n3455__));
  and1  g1994(.dina(new_new_n3454__), .dinb(new_new_n5026__), .dout(new_new_n3456__));
  or1   g1995(.dina(new_new_n3455__), .dinb(new_new_n5039__), .dout(new_new_n3457__));
  and1  g1996(.dina(new_new_n5056__), .dinb(new_new_n5212__), .dout(new_new_n3458__));
  or1   g1997(.dina(new_new_n5070__), .dinb(new_new_n5218__), .dout(new_new_n3459__));
  and1  g1998(.dina(new_new_n5077__), .dinb(new_new_n5254__), .dout(new_new_n3460__));
  or1   g1999(.dina(new_new_n5087__), .dinb(new_new_n1268__), .dout(new_new_n3461__));
  and1  g2000(.dina(new_new_n3459__), .dinb(new_new_n3457__), .dout(new_new_n3462__));
  or1   g2001(.dina(new_new_n3458__), .dinb(new_new_n3456__), .dout(new_new_n3463__));
  and1  g2002(.dina(new_new_n3462__), .dinb(new_new_n3461__), .dout(new_new_n3464__));
  or1   g2003(.dina(new_new_n3463__), .dinb(new_new_n3460__), .dout(new_new_n3465__));
  and1  g2004(.dina(new_new_n3465__), .dinb(new_new_n5107__), .dout(new_new_n3466__));
  or1   g2005(.dina(new_new_n3464__), .dinb(new_new_n5114__), .dout(new_new_n3467__));
  and1  g2006(.dina(new_new_n5122__), .dinb(new_new_n5080__), .dout(new_new_n3468__));
  or1   g2007(.dina(new_new_n5129__), .dinb(new_new_n5090__), .dout(new_new_n3469__));
  and1  g2008(.dina(new_new_n5133__), .dinb(new_new_n5091__), .dout(new_new_n3470__));
  or1   g2009(.dina(new_new_n5134__), .dinb(new_new_n5081__), .dout(new_new_n3471__));
  and1  g2010(.dina(new_new_n3470__), .dinb(new_new_n5141__), .dout(new_new_n3472__));
  or1   g2011(.dina(new_new_n3471__), .dinb(new_new_n5148__), .dout(new_new_n3473__));
  and1  g2012(.dina(new_new_n3469__), .dinb(new_new_n3467__), .dout(new_new_n3474__));
  or1   g2013(.dina(new_new_n3468__), .dinb(new_new_n3466__), .dout(new_new_n3475__));
  and1  g2014(.dina(new_new_n3474__), .dinb(new_new_n3473__), .dout(new_new_n3476__));
  or1   g2015(.dina(new_new_n3475__), .dinb(new_new_n3472__), .dout(new_new_n3477__));
  and1  g2016(.dina(new_new_n5155__), .dinb(new_new_n5184__), .dout(new_new_n3478__));
  or1   g2017(.dina(new_new_n5162__), .dinb(new_new_n5185__), .dout(new_new_n3479__));
  and1  g2018(.dina(new_new_n3478__), .dinb(new_new_n5166__), .dout(new_new_n3480__));
  or1   g2019(.dina(new_new_n3479__), .dinb(new_new_n5169__), .dout(new_new_n3481__));
  and1  g2020(.dina(new_new_n5063__), .dinb(new_new_n4957__), .dout(new_new_n3482__));
  or1   g2021(.dina(new_new_n5049__), .dinb(new_new_n4966__), .dout(new_new_n3483__));
  and1  g2022(.dina(new_new_n5255__), .dinb(new_new_n4976__), .dout(new_new_n3484__));
  or1   g2023(.dina(new_new_n2240__), .dinb(new_new_n4983__), .dout(new_new_n3485__));
  and1  g2024(.dina(new_new_n4989__), .dinb(new_new_n5238__), .dout(new_new_n3486__));
  or1   g2025(.dina(new_new_n4996__), .dinb(new_new_n5240__), .dout(new_new_n3487__));
  and1  g2026(.dina(new_new_n3485__), .dinb(new_new_n3483__), .dout(new_new_n3488__));
  or1   g2027(.dina(new_new_n3484__), .dinb(new_new_n3482__), .dout(new_new_n3489__));
  and1  g2028(.dina(new_new_n3488__), .dinb(new_new_n3487__), .dout(new_new_n3490__));
  or1   g2029(.dina(new_new_n3489__), .dinb(new_new_n3486__), .dout(new_new_n3491__));
  and1  g2030(.dina(new_new_n3491__), .dinb(new_new_n5155__), .dout(new_new_n3492__));
  or1   g2031(.dina(new_new_n3490__), .dinb(new_new_n5161__), .dout(new_new_n3493__));
  and1  g2032(.dina(new_new_n3481__), .dinb(new_new_n5187__), .dout(new_new_n3494__));
  or1   g2033(.dina(new_new_n3480__), .dinb(new_new_n5191__), .dout(new_new_n3495__));
  and1  g2034(.dina(new_new_n3494__), .dinb(new_new_n3493__), .dout(new_new_n3496__));
  or1   g2035(.dina(new_new_n3495__), .dinb(new_new_n3492__), .dout(new_new_n3497__));
  or1   g2036(.dina(new_new_n5258__), .dinb(new_new_n5199__), .dout(new_new_n3498__));
  or1   g2037(.dina(new_new_n3498__), .dinb(new_new_n5260__), .dout(new_new_n3499__));
  or1   g2038(.dina(new_new_n5258__), .dinb(new_new_n5205__), .dout(new_new_n3500__));
  or1   g2039(.dina(new_new_n3500__), .dinb(new_new_n5260__), .dout(new_new_n3501__));
  or1   g2040(.dina(new_new_n5261__), .dinb(new_new_n1278__), .dout(new_new_n3502__));
  or1   g2041(.dina(new_new_n5263__), .dinb(new_new_n1332__), .dout(new_new_n3503__));
  and1  g2042(.dina(new_new_n5026__), .dinb(new_new_n4948__), .dout(new_new_n3504__));
  or1   g2043(.dina(new_new_n5040__), .dinb(new_new_n4960__), .dout(new_new_n3505__));
  and1  g2044(.dina(new_new_n5056__), .dinb(new_new_n5012__), .dout(new_new_n3506__));
  or1   g2045(.dina(new_new_n5071__), .dinb(new_new_n5013__), .dout(new_new_n3507__));
  and1  g2046(.dina(new_new_n5077__), .dinb(new_new_n5236__), .dout(new_new_n3508__));
  or1   g2047(.dina(new_new_n5087__), .dinb(new_new_n5230__), .dout(new_new_n3509__));
  and1  g2048(.dina(new_new_n3507__), .dinb(new_new_n3505__), .dout(new_new_n3510__));
  or1   g2049(.dina(new_new_n3506__), .dinb(new_new_n3504__), .dout(new_new_n3511__));
  and1  g2050(.dina(new_new_n3510__), .dinb(new_new_n3509__), .dout(new_new_n3512__));
  or1   g2051(.dina(new_new_n3511__), .dinb(new_new_n3508__), .dout(new_new_n3513__));
  and1  g2052(.dina(new_new_n3513__), .dinb(new_new_n5107__), .dout(new_new_n3514__));
  or1   g2053(.dina(new_new_n3512__), .dinb(new_new_n5115__), .dout(new_new_n3515__));
  and1  g2054(.dina(new_new_n5122__), .dinb(new_new_n4959__), .dout(new_new_n3516__));
  or1   g2055(.dina(new_new_n5130__), .dinb(new_new_n4949__), .dout(new_new_n3517__));
  and1  g2056(.dina(new_new_n5248__), .dinb(new_new_n4949__), .dout(new_new_n3518__));
  or1   g2057(.dina(new_new_n5251__), .dinb(new_new_n4961__), .dout(new_new_n3519__));
  and1  g2058(.dina(new_new_n3518__), .dinb(new_new_n5141__), .dout(new_new_n3520__));
  or1   g2059(.dina(new_new_n3519__), .dinb(new_new_n5148__), .dout(new_new_n3521__));
  and1  g2060(.dina(new_new_n3517__), .dinb(new_new_n3515__), .dout(new_new_n3522__));
  or1   g2061(.dina(new_new_n3516__), .dinb(new_new_n3514__), .dout(new_new_n3523__));
  and1  g2062(.dina(new_new_n3522__), .dinb(new_new_n3521__), .dout(new_new_n3524__));
  or1   g2063(.dina(new_new_n3523__), .dinb(new_new_n3520__), .dout(new_new_n3525__));
  and1  g2064(.dina(new_new_n5264__), .dinb(new_new_n5265__), .dout(new_new_n3526__));
  and1  g2065(.dina(new_new_n5193__), .dinb(new_new_n5267__), .dout(new_new_n3527__));
  and1  g2066(.dina(new_new_n3527__), .dinb(new_new_n5269__), .dout(new_new_n3528__));
  and1  g2067(.dina(new_new_n5195__), .dinb(new_new_n5271__), .dout(new_new_n3529__));
  and1  g2068(.dina(new_new_n3529__), .dinb(new_new_n5269__), .dout(new_new_n3530__));
  or1   g2069(.dina(new_new_n3530__), .dinb(new_new_n3528__), .dout(new_new_n3531__));
  or1   g2070(.dina(new_new_n3531__), .dinb(new_new_n3299__), .dout(new_new_n3532__));
  and1  g2071(.dina(new_new_n3532__), .dinb(new_new_n3526__), .dout(new_new_n3533__));
  or1   g2072(.dina(new_new_n4856__), .dinb(new_new_n5273__), .dout(new_new_n3534__));
  or1   g2073(.dina(new_new_n3534__), .dinb(new_new_n4866__), .dout(new_new_n3535__));
  or1   g2074(.dina(new_new_n3535__), .dinb(new_new_n4880__), .dout(new_new_n3536__));
  or1   g2075(.dina(new_new_n5208__), .dinb(new_new_n5276__), .dout(new_new_n3537__));
  or1   g2076(.dina(new_new_n3537__), .dinb(new_new_n4841__), .dout(new_new_n3538__));
  or1   g2077(.dina(new_new_n5280__), .dinb(new_new_n5282__), .dout(new_new_n3539__));
  or1   g2078(.dina(new_new_n5285__), .dinb(new_new_n5287__), .dout(new_new_n3540__));
  and1  g2079(.dina(new_new_n5289__), .dinb(new_new_n5291__), .dout(new_new_n3541__));
  and1  g2080(.dina(new_new_n5285__), .dinb(new_new_n5287__), .dout(new_new_n3542__));
  or1   g2081(.dina(new_new_n5289__), .dinb(new_new_n5291__), .dout(new_new_n3543__));
  and1  g2082(.dina(new_new_n4894__), .dinb(new_new_n1727__), .dout(new_new_n3544__));
  or1   g2083(.dina(new_new_n4895__), .dinb(new_new_n1728__), .dout(new_new_n3545__));
  and1  g2084(.dina(new_new_n5292__), .dinb(new_new_n4686__), .dout(new_new_n3546__));
  or1   g2085(.dina(new_new_n5294__), .dinb(new_new_n4680__), .dout(new_new_n3547__));
  and1  g2086(.dina(new_new_n5294__), .dinb(new_new_n4681__), .dout(new_new_n3548__));
  or1   g2087(.dina(new_new_n5292__), .dinb(new_new_n4685__), .dout(new_new_n3549__));
  and1  g2088(.dina(new_new_n3549__), .dinb(new_new_n3547__), .dout(new_new_n3550__));
  or1   g2089(.dina(new_new_n3548__), .dinb(new_new_n3546__), .dout(new_new_n3551__));
  or1   g2090(.dina(new_new_n5296__), .dinb(new_new_n5299__), .dout(new_new_n3552__));
  or1   g2091(.dina(new_new_n3552__), .dinb(new_new_n5276__), .dout(new_new_n3553__));
  or1   g2092(.dina(new_new_n5299__), .dinb(new_new_n5277__), .dout(new_new_n3554__));
  or1   g2093(.dina(new_new_n5300__), .dinb(new_new_n5199__), .dout(new_new_n3555__));
  or1   g2094(.dina(new_new_n3555__), .dinb(new_new_n5303__), .dout(new_new_n3556__));
  or1   g2095(.dina(new_new_n5300__), .dinb(new_new_n5205__), .dout(new_new_n3557__));
  or1   g2096(.dina(new_new_n3557__), .dinb(new_new_n5303__), .dout(new_new_n3558__));
  or1   g2097(.dina(new_new_n5307__), .dinb(new_new_n5195__), .dout(new_new_n3559__));
  or1   g2098(.dina(new_new_n5309__), .dinb(new_new_n5277__), .dout(new_new_n3560__));
  and1  g2099(.dina(new_new_n4817__), .dinb(new_new_n4820__), .dout(new_new_n3561__));
  or1   g2100(.dina(new_new_n3561__), .dinb(new_new_n4822__), .dout(new_new_n3562__));
  and1  g2101(.dina(new_new_n1628__), .dinb(new_new_n5310__), .dout(new_new_n3563__));
  and1  g2102(.dina(new_new_n5311__), .dinb(new_new_n1626__), .dout(new_new_n3564__));
  or1   g2103(.dina(new_new_n3564__), .dinb(new_new_n3563__), .dout(new_new_n3565__));
  and1  g2104(.dina(new_new_n1676__), .dinb(new_new_n5312__), .dout(new_new_n3566__));
  and1  g2105(.dina(new_new_n5313__), .dinb(new_new_n1658__), .dout(new_new_n3567__));
  or1   g2106(.dina(new_new_n3567__), .dinb(new_new_n3566__), .dout(new_new_n3568__));
  and1  g2107(.dina(new_new_n5296__), .dinb(new_new_n3126__), .dout(new_new_n3569__));
  and1  g2108(.dina(new_new_n5315__), .dinb(new_new_n5316__), .dout(new_new_n3570__));
  or1   g2109(.dina(new_new_n3570__), .dinb(new_new_n3569__), .dout(new_new_n3571__));
  and1  g2110(.dina(new_new_n5282__), .dinb(new_new_n1530__), .dout(new_new_n3572__));
  and1  g2111(.dina(new_new_n1622__), .dinb(new_new_n5318__), .dout(new_new_n3573__));
  or1   g2112(.dina(new_new_n3573__), .dinb(new_new_n3572__), .dout(new_new_n3574__));
  and1  g2113(.dina(new_new_n1598__), .dinb(new_new_n5320__), .dout(new_new_n3575__));
  and1  g2114(.dina(new_new_n5323__), .dinb(new_new_n1536__), .dout(new_new_n3576__));
  or1   g2115(.dina(new_new_n3576__), .dinb(new_new_n3575__), .dout(new_new_n3577__));
  and1  g2116(.dina(new_new_n1737__), .dinb(new_new_n1729__), .dout(new_new_n3578__));
  or1   g2117(.dina(new_new_n1738__), .dinb(new_new_n1730__), .dout(new_new_n3579__));
  and1  g2118(.dina(new_new_n5325__), .dinb(new_new_n4688__), .dout(new_new_n3580__));
  or1   g2119(.dina(new_new_n5327__), .dinb(new_new_n4683__), .dout(new_new_n3581__));
  and1  g2120(.dina(new_new_n5327__), .dinb(new_new_n4684__), .dout(new_new_n3582__));
  or1   g2121(.dina(new_new_n5325__), .dinb(new_new_n4687__), .dout(new_new_n3583__));
  and1  g2122(.dina(new_new_n3583__), .dinb(new_new_n3581__), .dout(new_new_n3584__));
  or1   g2123(.dina(new_new_n3582__), .dinb(new_new_n3580__), .dout(new_new_n3585__));
  and1  g2124(.dina(new_new_n4670__), .dinb(new_new_n1943__), .dout(new_new_n3586__));
  or1   g2125(.dina(new_new_n4678__), .dinb(new_new_n1944__), .dout(new_new_n3587__));
  and1  g2126(.dina(new_new_n5315__), .dinb(new_new_n4823__), .dout(new_new_n3588__));
  or1   g2127(.dina(new_new_n5297__), .dinb(new_new_n4821__), .dout(new_new_n3589__));
  and1  g2128(.dina(new_new_n5314__), .dinb(new_new_n4815__), .dout(new_new_n3590__));
  or1   g2129(.dina(new_new_n5297__), .dinb(new_new_n4820__), .dout(new_new_n3591__));
  and1  g2130(.dina(new_new_n3590__), .dinb(new_new_n4814__), .dout(new_new_n3592__));
  or1   g2131(.dina(new_new_n3591__), .dinb(new_new_n4816__), .dout(new_new_n3593__));
  and1  g2132(.dina(new_new_n3589__), .dinb(new_new_n3587__), .dout(new_new_n3594__));
  or1   g2133(.dina(new_new_n3588__), .dinb(new_new_n3586__), .dout(new_new_n3595__));
  and1  g2134(.dina(new_new_n3594__), .dinb(new_new_n3593__), .dout(new_new_n3596__));
  or1   g2135(.dina(new_new_n3595__), .dinb(new_new_n3592__), .dout(new_new_n3597__));
  and1  g2136(.dina(new_new_n3596__), .dinb(new_new_n3585__), .dout(new_new_n3598__));
  and1  g2137(.dina(new_new_n3597__), .dinb(new_new_n3584__), .dout(new_new_n3599__));
  or1   g2138(.dina(new_new_n3599__), .dinb(new_new_n3598__), .dout(new_new_n3600__));
  and1  g2139(.dina(new_new_n4713__), .dinb(new_new_n5330__), .dout(new_new_n3601__));
  or1   g2140(.dina(new_new_n4716__), .dinb(new_new_n5333__), .dout(new_new_n3602__));
  and1  g2141(.dina(new_new_n4707__), .dinb(new_new_n5330__), .dout(new_new_n3603__));
  or1   g2142(.dina(new_new_n4708__), .dinb(new_new_n5333__), .dout(new_new_n3604__));
  or1   g2143(.dina(new_new_n5335__), .dinb(new_new_n4719__), .dout(new_new_n3605__));
  or1   g2144(.dina(new_new_n5336__), .dinb(new_new_n5338__), .dout(new_new_n3606__));
  or1   g2145(.dina(new_new_n5336__), .dinb(new_new_n5341__), .dout(new_new_n3607__));
  or1   g2146(.dina(new_new_n4718__), .dinb(new_new_n5332__), .dout(new_new_n3608__));
  and1  g2147(.dina(new_new_n5343__), .dinb(new_new_n3604__), .dout(new_new_n3609__));
  and1  g2148(.dina(new_new_n5344__), .dinb(new_new_n5338__), .dout(new_new_n3610__));
  or1   g2149(.dina(new_new_n5343__), .dinb(new_new_n5335__), .dout(new_new_n3611__));
  or1   g2150(.dina(new_new_n5345__), .dinb(new_new_n5341__), .dout(new_new_n3612__));
  or1   g2151(.dina(new_new_n5334__), .dinb(new_new_n4717__), .dout(new_new_n3613__));
  or1   g2152(.dina(new_new_n5346__), .dinb(new_new_n5342__), .dout(new_new_n3614__));
  and1  g2153(.dina(new_new_n5344__), .dinb(new_new_n5342__), .dout(new_new_n3615__));
  or1   g2154(.dina(new_new_n5345__), .dinb(new_new_n5339__), .dout(new_new_n3616__));
  or1   g2155(.dina(new_new_n5346__), .dinb(new_new_n5339__), .dout(new_new_n3617__));
  and1  g2156(.dina(new_new_n5347__), .dinb(new_new_n5348__), .dout(new_new_n3618__));
  and1  g2157(.dina(new_new_n5242__), .dinb(new_new_n5267__), .dout(new_new_n3619__));
  and1  g2158(.dina(new_new_n3619__), .dinb(new_new_n5349__), .dout(new_new_n3620__));
  and1  g2159(.dina(new_new_n5244__), .dinb(new_new_n5271__), .dout(new_new_n3621__));
  and1  g2160(.dina(new_new_n3621__), .dinb(new_new_n5349__), .dout(new_new_n3622__));
  or1   g2161(.dina(new_new_n3622__), .dinb(new_new_n3620__), .dout(new_new_n3623__));
  or1   g2162(.dina(new_new_n3623__), .dinb(new_new_n3359__), .dout(new_new_n3624__));
  and1  g2163(.dina(new_new_n3624__), .dinb(new_new_n3618__), .dout(new_new_n3625__));
  and1  g2164(.dina(new_new_n5351__), .dinb(new_new_n5353__), .dout(new_new_n3626__));
  or1   g2165(.dina(new_new_n3626__), .dinb(new_new_n5354__), .dout(new_new_n3627__));
  or1   g2166(.dina(new_new_n3627__), .dinb(new_new_n5357__), .dout(new_new_n3628__));
  or1   g2167(.dina(new_new_n3628__), .dinb(new_new_n5360__), .dout(new_new_n3629__));
  or1   g2168(.dina(new_new_n5273__), .dinb(new_new_n4879__), .dout(new_new_n3630__));
  or1   g2169(.dina(new_new_n5361__), .dinb(new_new_n4867__), .dout(new_new_n3631__));
  or1   g2170(.dina(new_new_n3631__), .dinb(new_new_n5279__), .dout(new_new_n3632__));
  or1   g2171(.dina(new_new_n5362__), .dinb(new_new_n5279__), .dout(new_new_n3633__));
  or1   g2172(.dina(new_new_n5361__), .dinb(new_new_n5278__), .dout(new_new_n3634__));
  and1  g2173(.dina(new_new_n4876__), .dinb(new_new_n4841__), .dout(new_new_n3635__));
  or1   g2174(.dina(new_new_n4881__), .dinb(new_new_n4884__), .dout(new_new_n3636__));
  and1  g2175(.dina(new_new_n3636__), .dinb(new_new_n4871__), .dout(new_new_n3637__));
  or1   g2176(.dina(new_new_n3635__), .dinb(new_new_n4874__), .dout(new_new_n3638__));
  and1  g2177(.dina(new_new_n3637__), .dinb(new_new_n4867__), .dout(new_new_n3639__));
  and1  g2178(.dina(new_new_n3638__), .dinb(new_new_n4862__), .dout(new_new_n3640__));
  or1   g2179(.dina(new_new_n3640__), .dinb(new_new_n3639__), .dout(new_new_n3641__));
  or1   g2180(.dina(new_new_n5307__), .dinb(new_new_n5244__), .dout(new_new_n3642__));
  and1  g2181(.dina(new_new_n5364__), .dinb(new_new_n5367__), .dout(new_new_n3643__));
  and1  g2182(.dina(new_new_n5370__), .dinb(new_new_n5372__), .dout(new_new_n3644__));
  or1   g2183(.dina(new_new_n5364__), .dinb(new_new_n5367__), .dout(new_new_n3645__));
  or1   g2184(.dina(new_new_n5370__), .dinb(new_new_n5372__), .dout(new_new_n3646__));
  and1  g2185(.dina(new_new_n5027__), .dinb(new_new_n5180__), .dout(new_new_n3647__));
  or1   g2186(.dina(new_new_n5040__), .dinb(new_new_n5173__), .dout(new_new_n3648__));
  and1  g2187(.dina(new_new_n5057__), .dinb(new_new_n4950__), .dout(new_new_n3649__));
  or1   g2188(.dina(new_new_n5071__), .dinb(new_new_n4961__), .dout(new_new_n3650__));
  and1  g2189(.dina(new_new_n5078__), .dinb(new_new_n5049__), .dout(new_new_n3651__));
  or1   g2190(.dina(new_new_n5086__), .dinb(new_new_n5063__), .dout(new_new_n3652__));
  and1  g2191(.dina(new_new_n3650__), .dinb(new_new_n3648__), .dout(new_new_n3653__));
  or1   g2192(.dina(new_new_n3649__), .dinb(new_new_n3647__), .dout(new_new_n3654__));
  and1  g2193(.dina(new_new_n3653__), .dinb(new_new_n3652__), .dout(new_new_n3655__));
  or1   g2194(.dina(new_new_n3654__), .dinb(new_new_n3651__), .dout(new_new_n3656__));
  and1  g2195(.dina(new_new_n3656__), .dinb(new_new_n5108__), .dout(new_new_n3657__));
  or1   g2196(.dina(new_new_n3655__), .dinb(new_new_n5115__), .dout(new_new_n3658__));
  and1  g2197(.dina(new_new_n5123__), .dinb(new_new_n5181__), .dout(new_new_n3659__));
  or1   g2198(.dina(new_new_n5130__), .dinb(new_new_n5175__), .dout(new_new_n3660__));
  and1  g2199(.dina(new_new_n5248__), .dinb(new_new_n5175__), .dout(new_new_n3661__));
  or1   g2200(.dina(new_new_n5251__), .dinb(new_new_n5181__), .dout(new_new_n3662__));
  and1  g2201(.dina(new_new_n3661__), .dinb(new_new_n5142__), .dout(new_new_n3663__));
  or1   g2202(.dina(new_new_n3662__), .dinb(new_new_n5147__), .dout(new_new_n3664__));
  and1  g2203(.dina(new_new_n3660__), .dinb(new_new_n3658__), .dout(new_new_n3665__));
  or1   g2204(.dina(new_new_n3659__), .dinb(new_new_n3657__), .dout(new_new_n3666__));
  and1  g2205(.dina(new_new_n3665__), .dinb(new_new_n3664__), .dout(new_new_n3667__));
  or1   g2206(.dina(new_new_n3666__), .dinb(new_new_n3663__), .dout(new_new_n3668__));
  and1  g2207(.dina(new_new_n5374__), .dinb(new_new_n5377__), .dout(new_new_n3669__));
  or1   g2208(.dina(new_new_n5380__), .dinb(new_new_n5200__), .dout(new_new_n3670__));
  and1  g2209(.dina(new_new_n3669__), .dinb(new_new_n5382__), .dout(new_new_n3671__));
  or1   g2210(.dina(new_new_n3670__), .dinb(new_new_n5385__), .dout(new_new_n3672__));
  and1  g2211(.dina(new_new_n5374__), .dinb(new_new_n5389__), .dout(new_new_n3673__));
  or1   g2212(.dina(new_new_n5380__), .dinb(new_new_n5206__), .dout(new_new_n3674__));
  and1  g2213(.dina(new_new_n3673__), .dinb(new_new_n5382__), .dout(new_new_n3675__));
  or1   g2214(.dina(new_new_n3674__), .dinb(new_new_n5385__), .dout(new_new_n3676__));
  and1  g2215(.dina(new_new_n3676__), .dinb(new_new_n3672__), .dout(new_new_n3677__));
  or1   g2216(.dina(new_new_n3675__), .dinb(new_new_n3671__), .dout(new_new_n3678__));
  and1  g2217(.dina(new_new_n5393__), .dinb(new_new_n5377__), .dout(new_new_n3679__));
  or1   g2218(.dina(new_new_n5396__), .dinb(new_new_n5200__), .dout(new_new_n3680__));
  and1  g2219(.dina(new_new_n3679__), .dinb(new_new_n5397__), .dout(new_new_n3681__));
  or1   g2220(.dina(new_new_n3680__), .dinb(new_new_n5400__), .dout(new_new_n3682__));
  and1  g2221(.dina(new_new_n5393__), .dinb(new_new_n5389__), .dout(new_new_n3683__));
  or1   g2222(.dina(new_new_n5396__), .dinb(new_new_n5206__), .dout(new_new_n3684__));
  and1  g2223(.dina(new_new_n3683__), .dinb(new_new_n5397__), .dout(new_new_n3685__));
  or1   g2224(.dina(new_new_n3684__), .dinb(new_new_n5400__), .dout(new_new_n3686__));
  and1  g2225(.dina(new_new_n3686__), .dinb(new_new_n3682__), .dout(new_new_n3687__));
  or1   g2226(.dina(new_new_n3685__), .dinb(new_new_n3681__), .dout(new_new_n3688__));
  or1   g2227(.dina(new_new_n5402__), .dinb(new_new_n5404__), .dout(new_new_n3689__));
  or1   g2228(.dina(new_new_n3689__), .dinb(new_new_n5329__), .dout(new_new_n3690__));
  or1   g2229(.dina(new_new_n5407__), .dinb(new_new_n5412__), .dout(new_new_n3691__));
  and1  g2230(.dina(new_new_n3691__), .dinb(new_new_n5416__), .dout(new_new_n3692__));
  and1  g2231(.dina(new_new_n5417__), .dinb(new_new_n4842__), .dout(new_new_n3693__));
  and1  g2232(.dina(new_new_n5418__), .dinb(new_new_n5419__), .dout(new_new_n3694__));
  and1  g2233(.dina(new_new_n3694__), .dinb(new_new_n5420__), .dout(new_new_n3695__));
  and1  g2234(.dina(new_new_n5421__), .dinb(new_new_n5422__), .dout(new_new_n3696__));
  and1  g2235(.dina(new_new_n4870__), .dinb(new_new_n4863__), .dout(new_new_n3697__));
  or1   g2236(.dina(new_new_n4873__), .dinb(new_new_n4868__), .dout(new_new_n3698__));
  and1  g2237(.dina(new_new_n4863__), .dinb(new_new_n4877__), .dout(new_new_n3699__));
  or1   g2238(.dina(new_new_n4868__), .dinb(new_new_n4881__), .dout(new_new_n3700__));
  and1  g2239(.dina(new_new_n3699__), .dinb(new_new_n4842__), .dout(new_new_n3701__));
  or1   g2240(.dina(new_new_n3700__), .dinb(new_new_n4883__), .dout(new_new_n3702__));
  and1  g2241(.dina(new_new_n3698__), .dinb(new_new_n4853__), .dout(new_new_n3703__));
  or1   g2242(.dina(new_new_n3697__), .dinb(new_new_n4850__), .dout(new_new_n3704__));
  and1  g2243(.dina(new_new_n3703__), .dinb(new_new_n3702__), .dout(new_new_n3705__));
  or1   g2244(.dina(new_new_n3704__), .dinb(new_new_n3701__), .dout(new_new_n3706__));
  and1  g2245(.dina(new_new_n3705__), .dinb(new_new_n4851__), .dout(new_new_n3707__));
  and1  g2246(.dina(new_new_n3706__), .dinb(new_new_n4856__), .dout(new_new_n3708__));
  or1   g2247(.dina(new_new_n3708__), .dinb(new_new_n3707__), .dout(new_new_n3709__));
  and1  g2248(.dina(new_new_n5425__), .dinb(new_new_n5353__), .dout(new_new_n3710__));
  or1   g2249(.dina(new_new_n5351__), .dinb(new_new_n5412__), .dout(new_new_n3711__));
  and1  g2250(.dina(new_new_n5350__), .dinb(new_new_n5413__), .dout(new_new_n3712__));
  or1   g2251(.dina(new_new_n5425__), .dinb(new_new_n5352__), .dout(new_new_n3713__));
  and1  g2252(.dina(new_new_n3713__), .dinb(new_new_n3711__), .dout(new_new_n3714__));
  or1   g2253(.dina(new_new_n3712__), .dinb(new_new_n3710__), .dout(new_new_n3715__));
  and1  g2254(.dina(new_new_n5357__), .dinb(new_new_n5407__), .dout(new_new_n3716__));
  or1   g2255(.dina(new_new_n5416__), .dinb(new_new_n5360__), .dout(new_new_n3717__));
  and1  g2256(.dina(new_new_n5415__), .dinb(new_new_n5359__), .dout(new_new_n3718__));
  or1   g2257(.dina(new_new_n5356__), .dinb(new_new_n5408__), .dout(new_new_n3719__));
  and1  g2258(.dina(new_new_n3719__), .dinb(new_new_n3717__), .dout(new_new_n3720__));
  or1   g2259(.dina(new_new_n3718__), .dinb(new_new_n3716__), .dout(new_new_n3721__));
  or1   g2260(.dina(new_new_n3721__), .dinb(new_new_n3714__), .dout(new_new_n3722__));
  or1   g2261(.dina(new_new_n3720__), .dinb(new_new_n3715__), .dout(new_new_n3723__));
  and1  g2262(.dina(new_new_n3723__), .dinb(new_new_n3722__), .dout(new_new_n3724__));
  and1  g2263(.dina(new_new_n5427__), .dinb(new_new_n4728__), .dout(new_new_n3725__));
  or1   g2264(.dina(new_new_n5429__), .dinb(new_new_n4724__), .dout(new_new_n3726__));
  and1  g2265(.dina(new_new_n5429__), .dinb(new_new_n4725__), .dout(new_new_n3727__));
  or1   g2266(.dina(new_new_n5427__), .dinb(new_new_n4727__), .dout(new_new_n3728__));
  and1  g2267(.dina(new_new_n3728__), .dinb(new_new_n3726__), .dout(new_new_n3729__));
  or1   g2268(.dina(new_new_n3727__), .dinb(new_new_n3725__), .dout(new_new_n3730__));
  and1  g2269(.dina(new_new_n3730__), .dinb(new_new_n5430__), .dout(new_new_n3731__));
  and1  g2270(.dina(new_new_n3729__), .dinb(new_new_n3173__), .dout(new_new_n3732__));
  or1   g2271(.dina(new_new_n3732__), .dinb(new_new_n3731__), .dout(new_new_n3733__));
  and1  g2272(.dina(new_new_n3137__), .dinb(new_new_n5431__), .dout(new_new_n3734__));
  and1  g2273(.dina(new_new_n5432__), .dinb(new_new_n3131__), .dout(new_new_n3735__));
  or1   g2274(.dina(new_new_n3735__), .dinb(new_new_n3734__), .dout(new_new_n3736__));
  and1  g2275(.dina(new_new_n5435__), .dinb(new_new_n5378__), .dout(new_new_n3737__));
  and1  g2276(.dina(new_new_n3737__), .dinb(new_new_n5437__), .dout(new_new_n3738__));
  and1  g2277(.dina(new_new_n5435__), .dinb(new_new_n5388__), .dout(new_new_n3739__));
  and1  g2278(.dina(new_new_n3739__), .dinb(new_new_n5437__), .dout(new_new_n3740__));
  or1   g2279(.dina(new_new_n3740__), .dinb(new_new_n3738__), .dout(new_new_n3741__));
  or1   g2280(.dina(new_new_n5434__), .dinb(new_new_n5439__), .dout(new_new_n3742__));
  or1   g2281(.dina(new_new_n3742__), .dinb(new_new_n5442__), .dout(new_new_n3743__));
  or1   g2282(.dina(new_new_n5436__), .dinb(new_new_n5444__), .dout(new_new_n3744__));
  or1   g2283(.dina(new_new_n3744__), .dinb(new_new_n5442__), .dout(new_new_n3745__));
  and1  g2284(.dina(new_new_n3745__), .dinb(new_new_n3743__), .dout(new_new_n3746__));
  and1  g2285(.dina(new_new_n3746__), .dinb(new_new_n3438__), .dout(new_new_n3747__));
  or1   g2286(.dina(new_new_n3747__), .dinb(new_new_n5446__), .dout(new_new_n3748__));
  or1   g2287(.dina(new_new_n5375__), .dinb(new_new_n5439__), .dout(new_new_n3749__));
  or1   g2288(.dina(new_new_n3749__), .dinb(new_new_n5384__), .dout(new_new_n3750__));
  or1   g2289(.dina(new_new_n5375__), .dinb(new_new_n5444__), .dout(new_new_n3751__));
  or1   g2290(.dina(new_new_n3751__), .dinb(new_new_n5386__), .dout(new_new_n3752__));
  and1  g2291(.dina(new_new_n3752__), .dinb(new_new_n3750__), .dout(new_new_n3753__));
  and1  g2292(.dina(new_new_n3753__), .dinb(new_new_n5381__), .dout(new_new_n3754__));
  or1   g2293(.dina(new_new_n3754__), .dinb(new_new_n5447__), .dout(new_new_n3755__));
  and1  g2294(.dina(new_new_n5448__), .dinb(new_new_n5449__), .dout(new_new_n3756__));
  and1  g2295(.dina(new_new_n5257__), .dinb(new_new_n5268__), .dout(new_new_n3757__));
  and1  g2296(.dina(new_new_n3757__), .dinb(new_new_n5450__), .dout(new_new_n3758__));
  and1  g2297(.dina(new_new_n5259__), .dinb(new_new_n5272__), .dout(new_new_n3759__));
  and1  g2298(.dina(new_new_n3759__), .dinb(new_new_n5450__), .dout(new_new_n3760__));
  or1   g2299(.dina(new_new_n3760__), .dinb(new_new_n3758__), .dout(new_new_n3761__));
  or1   g2300(.dina(new_new_n3761__), .dinb(new_new_n3477__), .dout(new_new_n3762__));
  and1  g2301(.dina(new_new_n3762__), .dinb(new_new_n3756__), .dout(new_new_n3763__));
  or1   g2302(.dina(new_new_n5392__), .dinb(new_new_n5440__), .dout(new_new_n3764__));
  or1   g2303(.dina(new_new_n3764__), .dinb(new_new_n5399__), .dout(new_new_n3765__));
  or1   g2304(.dina(new_new_n5394__), .dinb(new_new_n5445__), .dout(new_new_n3766__));
  or1   g2305(.dina(new_new_n3766__), .dinb(new_new_n5401__), .dout(new_new_n3767__));
  and1  g2306(.dina(new_new_n3767__), .dinb(new_new_n3765__), .dout(new_new_n3768__));
  and1  g2307(.dina(new_new_n3768__), .dinb(new_new_n5395__), .dout(new_new_n3769__));
  or1   g2308(.dina(new_new_n3769__), .dinb(new_new_n5451__), .dout(new_new_n3770__));
  or1   g2309(.dina(new_new_n5453__), .dinb(new_new_n5440__), .dout(new_new_n3771__));
  or1   g2310(.dina(new_new_n3771__), .dinb(new_new_n5302__), .dout(new_new_n3772__));
  or1   g2311(.dina(new_new_n5453__), .dinb(new_new_n5445__), .dout(new_new_n3773__));
  or1   g2312(.dina(new_new_n3773__), .dinb(new_new_n5304__), .dout(new_new_n3774__));
  or1   g2313(.dina(new_new_n5381__), .dinb(new_new_n5306__), .dout(new_new_n3775__));
  or1   g2314(.dina(new_new_n5263__), .dinb(new_new_n5259__), .dout(new_new_n3776__));
  and1  g2315(.dina(new_new_n5456__), .dinb(new_new_n5459__), .dout(new_new_n3777__));
  or1   g2316(.dina(new_new_n1227__), .dinb(new_new_n5459__), .dout(new_new_n3778__));
  or1   g2317(.dina(new_new_n5222__), .dinb(new_new_n5091__), .dout(new_new_n3779__));
  or1   g2318(.dina(new_new_n3779__), .dinb(new_new_n5218__), .dout(new_new_n3780__));
  and1  g2319(.dina(new_new_n3780__), .dinb(new_new_n5027__), .dout(new_new_n3781__));
  and1  g2320(.dina(new_new_n5057__), .dinb(new_new_n5081__), .dout(new_new_n3782__));
  and1  g2321(.dina(new_new_n5078__), .dinb(new_new_n5464__), .dout(new_new_n3783__));
  or1   g2322(.dina(new_new_n3782__), .dinb(new_new_n3781__), .dout(new_new_n3784__));
  or1   g2323(.dina(new_new_n3784__), .dinb(new_new_n3783__), .dout(new_new_n3785__));
  and1  g2324(.dina(new_new_n3785__), .dinb(new_new_n5108__), .dout(new_new_n3786__));
  and1  g2325(.dina(new_new_n5123__), .dinb(new_new_n5224__), .dout(new_new_n3787__));
  and1  g2326(.dina(new_new_n5133__), .dinb(new_new_n5221__), .dout(new_new_n3788__));
  and1  g2327(.dina(new_new_n3788__), .dinb(new_new_n5142__), .dout(new_new_n3789__));
  or1   g2328(.dina(new_new_n3787__), .dinb(new_new_n3786__), .dout(new_new_n3790__));
  or1   g2329(.dina(new_new_n3790__), .dinb(new_new_n3789__), .dout(new_new_n3791__));
  or1   g2330(.dina(new_new_n5466__), .dinb(new_new_n5468__), .dout(new_new_n3792__));
  or1   g2331(.dina(new_new_n3792__), .dinb(new_new_n3677__), .dout(new_new_n3793__));
  or1   g2332(.dina(new_new_n5468__), .dinb(new_new_n3687__), .dout(new_new_n3794__));
  and1  g2333(.dina(new_new_n5156__), .dinb(new_new_n5239__), .dout(new_new_n3795__));
  and1  g2334(.dina(new_new_n3795__), .dinb(new_new_n5166__), .dout(new_new_n3796__));
  and1  g2335(.dina(new_new_n5033__), .dinb(new_new_n4957__), .dout(new_new_n3797__));
  and1  g2336(.dina(new_new_n4976__), .dinb(new_new_n1281__), .dout(new_new_n3798__));
  and1  g2337(.dina(new_new_n4988__), .dinb(new_new_n5255__), .dout(new_new_n3799__));
  or1   g2338(.dina(new_new_n3798__), .dinb(new_new_n3797__), .dout(new_new_n3800__));
  or1   g2339(.dina(new_new_n3800__), .dinb(new_new_n3799__), .dout(new_new_n3801__));
  and1  g2340(.dina(new_new_n3801__), .dinb(new_new_n5156__), .dout(new_new_n3802__));
  or1   g2341(.dina(new_new_n3796__), .dinb(new_new_n5191__), .dout(new_new_n3803__));
  or1   g2342(.dina(new_new_n3803__), .dinb(new_new_n3802__), .dout(new_new_n3804__));
  or1   g2343(.dina(new_new_n5466__), .dinb(new_new_n5470__), .dout(new_new_n3805__));
  or1   g2344(.dina(new_new_n3805__), .dinb(new_new_n5472__), .dout(new_new_n3806__));
  or1   g2345(.dina(new_new_n3806__), .dinb(new_new_n5469__), .dout(new_new_n3807__));
  or1   g2346(.dina(new_new_n5473__), .dinb(new_new_n5456__), .dout(new_new_n3808__));
  and1  g2347(.dina(new_new_n5460__), .dinb(new_new_n1136__), .dout(new_new_n3809__));
  and1  g2348(.dina(new_new_n5475__), .dinb(new_new_n5460__), .dout(new_new_n3810__));
  and1  g2349(.dina(new_new_n5477__), .dinb(new_new_n5478__), .dout(new_new_n3811__));
  buf1  g2350(.din(new_new_n2291__), .dout(G3519));
  buf1  g2351(.din(new_new_n2292__), .dout(G3520));
  buf1  g2352(.din(new_new_n2323__), .dout(G3521));
  buf1  g2353(.din(new_new_n2332__), .dout(G3522));
  buf1  g2354(.din(new_new_n2335__), .dout(G3523));
  buf1  g2355(.din(new_new_n2336__), .dout(G3524));
  buf1  g2356(.din(new_new_n2338__), .dout(G3525));
  buf1  g2357(.din(new_new_n2340__), .dout(G3526));
  buf1  g2358(.din(new_new_n2347__), .dout(G3527));
  buf1  g2359(.din(new_new_n2350__), .dout(G3528));
  buf1  g2360(.din(new_new_n2353__), .dout(G3529));
  buf1  g2361(.din(new_new_n2387__), .dout(G3530));
  buf1  g2362(.din(new_new_n2390__), .dout(G3531));
  buf1  g2363(.din(new_new_n2393__), .dout(G3532));
  buf1  g2364(.din(new_new_n2396__), .dout(G3533));
  buf1  g2365(.din(new_new_n1641__), .dout(G3534));
  buf1  g2366(.din(new_new_n1643__), .dout(G3535));
  buf1  g2367(.din(new_new_n2399__), .dout(G3536));
  buf1  g2368(.din(new_new_n4397__), .dout(G3537));
  not1  g2369(.din(new_new_n2416__), .dout(G3538));
  buf1  g2370(.din(new_new_n2477__), .dout(G3539));
  buf1  g2371(.din(new_new_n2492__), .dout(G3540));
  buf1  g2372(.din(new_new_n1393__), .dout(n8948));
  buf1  g2373(.din(new_new_n4655__), .dout(n8951));
  buf1  g2374(.din(new_new_n1395__), .dout(n8954));
  buf1  g2375(.din(new_new_n1159__), .dout(n8957));
  buf1  g2376(.din(new_new_n1237__), .dout(n8960));
  buf1  g2377(.din(new_new_n1239__), .dout(n8963));
  buf1  g2378(.din(new_new_n1161__), .dout(n8966));
  buf1  g2379(.din(new_new_n1243__), .dout(n8969));
  buf1  g2380(.din(new_new_n1245__), .dout(n8972));
  buf1  g2381(.din(new_new_n1163__), .dout(n8975));
  buf1  g2382(.din(new_new_n1249__), .dout(n8978));
  buf1  g2383(.din(new_new_n1165__), .dout(n8981));
  buf1  g2384(.din(new_new_n1253__), .dout(n8984));
  buf1  g2385(.din(new_new_n1167__), .dout(n8987));
  buf1  g2386(.din(new_new_n1257__), .dout(n8990));
  buf1  g2387(.din(new_new_n1169__), .dout(n8993));
  buf1  g2388(.din(new_new_n1261__), .dout(n8996));
  buf1  g2389(.din(new_new_n1171__), .dout(n8999));
  buf1  g2390(.din(new_new_n1173__), .dout(n9002));
  buf1  g2391(.din(new_new_n1175__), .dout(n9005));
  buf1  g2392(.din(new_new_n1177__), .dout(n9008));
  buf1  g2393(.din(new_new_n1179__), .dout(n9011));
  buf1  g2394(.din(new_new_n1181__), .dout(n9014));
  buf1  g2395(.din(new_new_n1183__), .dout(n9017));
  buf1  g2396(.din(new_new_n4888__), .dout(n9020));
  buf1  g2397(.din(new_new_n1185__), .dout(n9023));
  buf1  g2398(.din(new_new_n1431__), .dout(n9026));
  buf1  g2399(.din(new_new_n1427__), .dout(n9029));
  buf1  g2400(.din(new_new_n1429__), .dout(n9032));
  buf1  g2401(.din(new_new_n1437__), .dout(n9035));
  buf1  g2402(.din(new_new_n1439__), .dout(n9038));
  buf1  g2403(.din(new_new_n1441__), .dout(n9041));
  buf1  g2404(.din(new_new_n1201__), .dout(n9044));
  buf1  g2405(.din(new_new_n1453__), .dout(n9047));
  buf1  g2406(.din(new_new_n1203__), .dout(n9050));
  buf1  g2407(.din(new_new_n1463__), .dout(n9053));
  buf1  g2408(.din(new_new_n1211__), .dout(n9056));
  buf1  g2409(.din(new_new_n1213__), .dout(n9059));
  buf1  g2410(.din(new_new_n1305__), .dout(n9062));
  buf1  g2411(.din(new_new_n1215__), .dout(n9065));
  buf1  g2412(.din(new_new_n1309__), .dout(n9068));
  buf1  g2413(.din(new_new_n1217__), .dout(n9071));
  buf1  g2414(.din(new_new_n1313__), .dout(n9074));
  buf1  g2415(.din(new_new_n1219__), .dout(n9077));
  buf1  g2416(.din(new_new_n1317__), .dout(n9080));
  buf1  g2417(.din(new_new_n1221__), .dout(n9083));
  buf1  g2418(.din(new_new_n1321__), .dout(n9086));
  buf1  g2419(.din(new_new_n1223__), .dout(n9089));
  buf1  g2420(.din(new_new_n1325__), .dout(n9092));
  buf1  g2421(.din(new_new_n4606__), .dout(n9095));
  buf1  g2422(.din(new_new_n1225__), .dout(n9098));
  buf1  g2423(.din(new_new_n1229__), .dout(n9101));
  buf1  g2424(.din(new_new_n1333__), .dout(n9104));
  buf1  g2425(.din(new_new_n1335__), .dout(n9107));
  buf1  g2426(.din(new_new_n1337__), .dout(n9110));
  buf1  g2427(.din(new_new_n1399__), .dout(n9113));
  buf1  g2428(.din(new_new_n1401__), .dout(n9116));
  buf1  g2429(.din(new_new_n1447__), .dout(n9119));
  buf1  g2430(.din(new_new_n1471__), .dout(n9122));
  buf1  g2431(.din(new_new_n1465__), .dout(n9125));
  buf1  g2432(.din(new_new_n1491__), .dout(n9128));
  buf1  g2433(.din(new_new_n1531__), .dout(n9131));
  buf1  g2434(.din(new_new_n1561__), .dout(n9134));
  buf1  g2435(.din(new_new_n1565__), .dout(n9137));
  buf1  g2436(.din(new_new_n1647__), .dout(n9140));
  buf1  g2437(.din(new_new_n1649__), .dout(n9143));
  buf1  g2438(.din(new_new_n1651__), .dout(n9146));
  buf1  g2439(.din(new_new_n1653__), .dout(n9149));
  buf1  g2440(.din(new_new_n1663__), .dout(n9152));
  buf1  g2441(.din(new_new_n1665__), .dout(n9155));
  buf1  g2442(.din(new_new_n1705__), .dout(n9158));
  buf1  g2443(.din(new_new_n1707__), .dout(n9161));
  buf1  g2444(.din(new_new_n1711__), .dout(n9164));
  buf1  g2445(.din(new_new_n4447__), .dout(n9167));
  buf1  g2446(.din(new_new_n4446__), .dout(n9170));
  buf1  g2447(.din(new_new_n4449__), .dout(n9173));
  buf1  g2448(.din(new_new_n4489__), .dout(n9176));
  buf1  g2449(.din(new_new_n1755__), .dout(n9179));
  buf1  g2450(.din(new_new_n1761__), .dout(n9182));
  buf1  g2451(.din(new_new_n1757__), .dout(n9185));
  buf1  g2452(.din(new_new_n1763__), .dout(n9188));
  buf1  g2453(.din(new_new_n5408__), .dout(n9191));
  buf1  g2454(.din(new_new_n5320__), .dout(n9194));
  buf1  g2455(.din(new_new_n1539__), .dout(n9197));
  buf1  g2456(.din(new_new_n1541__), .dout(n9200));
  buf1  g2457(.din(new_new_n1543__), .dout(n9203));
  buf1  g2458(.din(new_new_n5404__), .dout(n9206));
  buf1  g2459(.din(new_new_n5481__), .dout(n9209));
  buf1  g2460(.din(new_new_n4484__), .dout(n9212));
  buf1  g2461(.din(new_new_n4614__), .dout(n9215));
  buf1  g2462(.din(new_new_n4526__), .dout(n9218));
  buf1  g2463(.din(new_new_n4531__), .dout(n9221));
  buf1  g2464(.din(new_new_n4536__), .dout(n9224));
  buf1  g2465(.din(new_new_n4542__), .dout(n9227));
  buf1  g2466(.din(new_new_n4547__), .dout(n9230));
  buf1  g2467(.din(new_new_n4653__), .dout(n9233));
  buf1  g2468(.din(new_new_n1965__), .dout(n9236));
  buf1  g2469(.din(new_new_n5323__), .dout(n9239));
  buf1  g2470(.din(new_new_n4828__), .dout(n9242));
  buf1  g2471(.din(new_new_n4831__), .dout(n9245));
  buf1  g2472(.din(new_new_n4824__), .dout(n9248));
  buf1  g2473(.din(new_new_n4457__), .dout(n9251));
  buf1  g2474(.din(new_new_n4654__), .dout(n9254));
  buf1  g2475(.din(new_new_n4833__), .dout(n9257));
  buf1  g2476(.din(new_new_n5310__), .dout(n9260));
  buf1  g2477(.din(new_new_n5311__), .dout(n9263));
  buf1  g2478(.din(new_new_n1629__), .dout(n9266));
  buf1  g2479(.din(new_new_n1631__), .dout(n9269));
  buf1  g2480(.din(new_new_n1609__), .dout(n9272));
  buf1  g2481(.din(new_new_n1613__), .dout(n9275));
  buf1  g2482(.din(new_new_n1655__), .dout(n9278));
  buf1  g2483(.din(new_new_n5312__), .dout(n9281));
  buf1  g2484(.din(new_new_n1659__), .dout(n9284));
  buf1  g2485(.din(new_new_n4624__), .dout(n9287));
  not1  g2486(.din(new_new_n4648__), .dout(n9290));
  buf1  g2487(.din(new_new_n4702__), .dout(n9293));
  buf1  g2488(.din(new_new_n5313__), .dout(n9296));
  buf1  g2489(.din(new_new_n1677__), .dout(n9299));
  buf1  g2490(.din(new_new_n1679__), .dout(n9302));
  buf1  g2491(.din(new_new_n1681__), .dout(n9305));
  buf1  g2492(.din(new_new_n1683__), .dout(n9308));
  buf1  g2493(.din(new_new_n4459__), .dout(n9311));
  buf1  g2494(.din(new_new_n1721__), .dout(n9314));
  buf1  g2495(.din(new_new_n4660__), .dout(n9317));
  buf1  g2496(.din(new_new_n4662__), .dout(n9320));
  buf1  g2497(.din(new_new_n4593__), .dout(n9323));
  buf1  g2498(.din(new_new_n1789__), .dout(n9326));
  buf1  g2499(.din(new_new_n1853__), .dout(n9329));
  buf1  g2500(.din(new_new_n4848__), .dout(n9332));
  buf1  g2501(.din(new_new_n4846__), .dout(n9335));
  buf1  g2502(.din(new_new_n4671__), .dout(n9338));
  buf1  g2503(.din(new_new_n4732__), .dout(n9341));
  not1  g2504(.din(new_new_n4735__), .dout(n9344));
  not1  g2505(.din(new_new_n4738__), .dout(n9347));
  not1  g2506(.din(new_new_n4741__), .dout(n9350));
  not1  g2507(.din(new_new_n4739__), .dout(n9353));
  not1  g2508(.din(new_new_n4740__), .dout(n9356));
  buf1  g2509(.din(new_new_n4783__), .dout(n9359));
  not1  g2510(.din(new_new_n4782__), .dout(n9362));
  buf1  g2511(.din(new_new_n4731__), .dout(n9365));
  not1  g2512(.din(new_new_n4742__), .dout(n9368));
  buf1  g2513(.din(new_new_n4733__), .dout(n9371));
  not1  g2514(.din(new_new_n4736__), .dout(n9374));
  buf1  g2515(.din(new_new_n4784__), .dout(n9377));
  not1  g2516(.din(new_new_n4737__), .dout(n9380));
  not1  g2517(.din(new_new_n4734__), .dout(n9383));
  buf1  g2518(.din(new_new_n4885__), .dout(n9386));
  buf1  g2519(.din(new_new_n5098__), .dout(n9389));
  buf1  g2520(.din(new_new_n5219__), .dout(n9392));
  buf1  g2521(.din(new_new_n5176__), .dout(n9395));
  buf1  g2522(.din(new_new_n4795__), .dout(n9398));
  buf1  g2523(.din(new_new_n5092__), .dout(n9401));
  buf1  g2524(.din(new_new_n5231__), .dout(n9404));
  buf1  g2525(.din(new_new_n4877__), .dout(n9407));
  buf1  g2526(.din(new_new_n2167__), .dout(n9410));
  buf1  g2527(.din(new_new_n2169__), .dout(n9413));
  buf1  g2528(.din(new_new_n2171__), .dout(n9416));
  buf1  g2529(.din(new_new_n4908__), .dout(n9419));
  buf1  g2530(.din(new_new_n4901__), .dout(n9422));
  buf1  g2531(.din(new_new_n5096__), .dout(n9425));
  buf1  g2532(.din(new_new_n4919__), .dout(n9428));
  buf1  g2533(.din(new_new_n4887__), .dout(n9431));
  buf1  g2534(.din(new_new_n4886__), .dout(n9434));
  buf1  g2535(.din(new_new_n5413__), .dout(n9437));
  buf1  g2536(.din(new_new_n5409__), .dout(n9440));
  buf1  g2537(.din(new_new_n5424__), .dout(n9443));
  not1  g2538(.din(new_new_n4797__), .dout(n9446));
  not1  g2539(.din(new_new_n4836__), .dout(n9449));
  not1  g2540(.din(new_new_n4800__), .dout(n9452));
  buf1  g2541(.din(new_new_n5428__), .dout(n9455));
  buf1  g2542(.din(new_new_n5286__), .dout(n9458));
  not1  g2543(.din(new_new_n5290__), .dout(n9461));
  not1  g2544(.din(new_new_n5484__), .dout(n9464));
  not1  g2545(.din(new_new_n5284__), .dout(n9467));
  not1  g2546(.din(new_new_n4803__), .dout(n9470));
  not1  g2547(.din(new_new_n4801__), .dout(n9473));
  not1  g2548(.din(new_new_n4798__), .dout(n9476));
  not1  g2549(.din(new_new_n4804__), .dout(n9479));
  not1  g2550(.din(new_new_n4799__), .dout(n9482));
  not1  g2551(.din(new_new_n4796__), .dout(n9485));
  not1  g2552(.din(new_new_n4802__), .dout(n9488));
  not1  g2553(.din(new_new_n5288__), .dout(n9491));
  buf1  g2554(.din(new_new_n4725__), .dout(n9494));
  buf1  g2555(.din(new_new_n5064__), .dout(n9497));
  buf1  g2556(.din(new_new_n5184__), .dout(n9500));
  buf1  g2557(.din(new_new_n4969__), .dout(n9503));
  buf1  g2558(.din(new_new_n5032__), .dout(n9506));
  buf1  g2559(.din(new_new_n5239__), .dout(n9509));
  buf1  g2560(.din(new_new_n5207__), .dout(n9512));
  buf1  g2561(.din(n9392), .dout(n9515));
  buf1  g2562(.din(n9395), .dout(n9518));
  buf1  g2563(.din(new_new_n5001__), .dout(n9521));
  buf1  g2564(.din(n9404), .dout(n9524));
  buf1  g2565(.din(n9497), .dout(n9527));
  buf1  g2566(.din(new_new_n5223__), .dout(n9530));
  buf1  g2567(.din(new_new_n4950__), .dout(n9533));
  buf1  g2568(.din(new_new_n4992__), .dout(n9536));
  buf1  g2569(.din(new_new_n4931__), .dout(n9539));
  buf1  g2570(.din(new_new_n5004__), .dout(n9542));
  buf1  g2571(.din(new_new_n5011__), .dout(n9545));
  buf1  g2572(.din(new_new_n5019__), .dout(n9548));
  buf1  g2573(.din(new_new_n5318__), .dout(n9551));
  buf1  g2574(.din(new_new_n5321__), .dout(n9554));
  buf1  g2575(.din(new_new_n5324__), .dout(n9557));
  buf1  g2576(.din(new_new_n5283__), .dout(n9560));
  not1  g2577(.din(new_new_n4891__), .dout(n9563));
  not1  g2578(.din(new_new_n4893__), .dout(n9566));
  not1  g2579(.din(new_new_n5487__), .dout(n9569));
  buf1  g2580(.din(new_new_n4843__), .dout(n9572));
  buf1  g2581(.din(new_new_n5316__), .dout(n9575));
  buf1  g2582(.din(new_new_n5431__), .dout(n9578));
  buf1  g2583(.din(new_new_n5432__), .dout(n9581));
  buf1  g2584(.din(new_new_n5254__), .dout(n9584));
  buf1  g2585(.din(new_new_n5017__), .dout(n9587));
  buf1  g2586(.din(new_new_n5253__), .dout(n9590));
  buf1  g2587(.din(new_new_n5419__), .dout(n9593));
  not1  g2588(.din(new_new_n5420__), .dout(n9596));
  buf1  g2589(.din(new_new_n5430__), .dout(n9599));
  buf1  g2590(.din(new_new_n5378__), .dout(n9602));
  buf1  g2591(.din(new_new_n5390__), .dout(n9605));
  buf1  g2592(.din(new_new_n5268__), .dout(n9608));
  buf1  g2593(.din(new_new_n5272__), .dout(n9611));
  buf1  g2594(.din(new_new_n5252__), .dout(n9614));
  buf1  g2595(.din(n9401), .dout(n9617));
  buf1  g2596(.din(n9422), .dout(n9620));
  buf1  g2597(.din(n9425), .dout(n9623));
  buf1  g2598(.din(n9530), .dout(n9626));
  not1  g2599(.din(new_new_n5489__), .dout(n9629));
  not1  g2600(.din(new_new_n5490__), .dout(n9632));
  buf1  g2601(.din(n9464), .dout(n9635));
  buf1  g2602(.din(n9569), .dout(n9638));
  buf1  g2603(.din(new_new_n5309__), .dout(n9641));
  buf1  g2604(.din(new_new_n5441__), .dout(n9644));
  buf1  g2605(.din(new_new_n5401__), .dout(n9647));
  buf1  g2606(.din(new_new_n5386__), .dout(n9650));
  not1  g2607(.din(new_new_n5265__), .dout(n9653));
  not1  g2608(.din(new_new_n5264__), .dout(n9656));
  buf1  g2609(.din(new_new_n5414__), .dout(n9659));
  buf1  g2610(.din(new_new_n5426__), .dout(n9662));
  buf1  g2611(.din(new_new_n5280__), .dout(n9665));
  not1  g2612(.din(new_new_n5298__), .dout(n9668));
  buf1  g2613(.din(new_new_n5418__), .dout(n9671));
  buf1  g2614(.din(new_new_n5261__), .dout(n9674));
  not1  g2615(.din(new_new_n5348__), .dout(n9677));
  not1  g2616(.din(new_new_n5347__), .dout(n9680));
  buf1  g2617(.din(new_new_n5464__), .dout(n9683));
  buf1  g2618(.din(new_new_n1277__), .dout(n9686));
  buf1  g2619(.din(new_new_n1331__), .dout(n9689));
  buf1  g2620(.din(new_new_n5394__), .dout(n9692));
  buf1  g2621(.din(new_new_n5436__), .dout(n9695));
  buf1  g2622(.din(new_new_n5304__), .dout(n9698));
  not1  g2623(.din(new_new_n5449__), .dout(n9701));
  not1  g2624(.din(new_new_n5448__), .dout(n9704));
  not1  g2625(.din(new_new_n5308__), .dout(n9707));
  buf1  g2626(.din(new_new_n5454__), .dout(n9710));
  buf1  g2627(.din(new_new_n5492__), .dout(n9713));
  buf1  g2628(.din(new_new_n1713__), .dout(n9716));
  buf1  g2629(.din(new_new_n1759__), .dout(n9719));
  buf1  g2630(.din(new_new_n5403__), .dout(n9722));
  buf1  g2631(.din(new_new_n5402__), .dout(n9725));
  buf1  g2632(.din(new_new_n5331__), .dout(n9728));
  buf1  g2633(.din(new_new_n5358__), .dout(n9731));
  buf1  g2634(.din(n9731), .dout(n9734));
  buf1  g2635(.din(n9386), .dout(n9737));
  not1  g2636(.din(new_new_n5362__), .dout(n9740));
  not1  g2637(.din(new_new_n5417__), .dout(n9743));
  buf1  g2638(.din(new_new_n5354__), .dout(n9746));
  not1  g2639(.din(new_new_n4890__), .dout(n9749));
  not1  g2640(.din(new_new_n4892__), .dout(n9752));
  not1  g2641(.din(new_new_n3540__), .dout(n9755));
  not1  g2642(.din(new_new_n3541__), .dout(n9758));
  not1  g2643(.din(new_new_n5485__), .dout(n9761));
  buf1  g2644(.din(new_new_n3542__), .dout(n9764));
  not1  g2645(.din(new_new_n5488__), .dout(n9767));
  not1  g2646(.din(new_new_n3543__), .dout(n9770));
  not1  g2647(.din(new_new_n5494__), .dout(n9773));
  not1  g2648(.din(new_new_n5495__), .dout(n9776));
  not1  g2649(.din(new_new_n5422__), .dout(n9779));
  not1  g2650(.din(new_new_n5421__), .dout(n9782));
  not1  g2651(.din(new_new_n5497__), .dout(n9785));
  buf1  g2652(.din(n9629), .dout(n9788));
  buf1  g2653(.din(n9632), .dout(n9791));
  buf1  g2654(.din(n9761), .dout(n9794));
  buf1  g2655(.din(n9767), .dout(n9797));
  not1  g2656(.din(new_new_n5368__), .dout(n9800));
  not1  g2657(.din(new_new_n5365__), .dout(n9803));
  buf1  g2658(.din(n9209), .dout(n9806));
  buf1  g2659(.din(new_new_n5480__), .dout(n9809));
  buf1  g2660(.din(new_new_n5498__), .dout(n9812));
  buf1  g2661(.din(new_new_n5499__), .dout(n9815));
  buf1  g2662(.din(new_new_n5500__), .dout(n9818));
  buf1  g2663(.din(new_new_n5501__), .dout(n9821));
  buf1  g2664(.din(new_new_n5502__), .dout(n9824));
  buf1  g2665(.din(new_new_n5503__), .dout(n9827));
  not1  g2666(.din(new_new_n5507__), .dout(n9830));
  buf1  g2667(.din(n9830), .dout(n9833));
  not1  g2668(.din(new_new_n5518__), .dout(n9836));
  buf1  g2669(.din(n9836), .dout(n9839));
  not1  g2670(.din(new_new_n5529__), .dout(n9842));
  buf1  g2671(.din(n9842), .dout(n9845));
  not1  g2672(.din(new_new_n5540__), .dout(n9848));
  buf1  g2673(.din(n9848), .dout(n9851));
  buf1  g2674(.din(new_new_n5551__), .dout(n9854));
  buf1  g2675(.din(n9854), .dout(n9857));
  buf1  g2676(.din(new_new_n5562__), .dout(n9860));
  buf1  g2677(.din(n9860), .dout(n9863));
  not1  g2678(.din(new_new_n5573__), .dout(n9866));
  buf1  g2679(.din(n9866), .dout(n9869));
  not1  g2680(.din(new_new_n5584__), .dout(n9872));
  buf1  g2681(.din(n9872), .dout(n9875));
  buf1  g2682(.din(new_new_n5593__), .dout(n9878));
  buf1  g2683(.din(n9713), .dout(n9881));
  buf1  g2684(.din(new_new_n5462__), .dout(n9884));
  buf1  g2685(.din(new_new_n5595__), .dout(n9887));
  buf1  g2686(.din(new_new_n5598__), .dout(n9890));
  buf1  g2687(.din(new_new_n1251__), .dout(n9893));
  buf1  g2688(.din(new_new_n1255__), .dout(n9896));
  buf1  g2689(.din(new_new_n1259__), .dout(n9899));
  buf1  g2690(.din(new_new_n1263__), .dout(n9902));
  buf1  g2691(.din(new_new_n1307__), .dout(n9905));
  buf1  g2692(.din(new_new_n1311__), .dout(n9908));
  buf1  g2693(.din(new_new_n1315__), .dout(n9911));
  buf1  g2694(.din(new_new_n1319__), .dout(n9914));
  buf1  g2695(.din(new_new_n1323__), .dout(n9917));
  buf1  g2696(.din(new_new_n1525__), .dout(n9920));
  buf1  g2697(.din(n9659), .dout(n9923));
  buf1  g2698(.din(new_new_n5317__), .dout(n9926));
  buf1  g2699(.din(n9440), .dout(n9929));
  not1  g2700(.din(new_new_n3629__), .dout(n9932));
  buf1  g2701(.din(n9554), .dout(n9935));
  buf1  g2702(.din(n9728), .dout(n9938));
  buf1  g2703(.din(n9557), .dout(n9941));
  buf1  g2704(.din(n9662), .dout(n9944));
  buf1  g2705(.din(n9560), .dout(n9947));
  buf1  g2706(.din(new_new_n1927__), .dout(n9950));
  buf1  g2707(.din(new_new_n2157__), .dout(n9953));
  buf1  g2708(.din(new_new_n4812__), .dout(n9956));
  buf1  g2709(.din(new_new_n4810__), .dout(n9959));
  buf1  g2710(.din(new_new_n5293__), .dout(n9962));
  buf1  g2711(.din(new_new_n4681__), .dout(n9965));
  buf1  g2712(.din(new_new_n5326__), .dout(n9968));
  buf1  g2713(.din(new_new_n4897__), .dout(n9971));
  buf1  g2714(.din(new_new_n4684__), .dout(n9974));
  buf1  g2715(.din(new_new_n4691__), .dout(n9977));
  not1  g2716(.din(new_new_n3632__), .dout(n9980));
  not1  g2717(.din(new_new_n3633__), .dout(n9983));
  not1  g2718(.din(new_new_n5371__), .dout(n9986));
  not1  g2719(.din(new_new_n5369__), .dout(n9989));
  not1  g2720(.din(new_new_n5600__), .dout(n9992));
  not1  g2721(.din(new_new_n5262__), .dout(n9995));
  buf1  g2722(.din(n9707), .dout(n9998));
  not1  g2723(.din(new_new_n3643__), .dout(n10001));
  not1  g2724(.din(new_new_n3644__), .dout(n10004));
  not1  g2725(.din(new_new_n3645__), .dout(n10007));
  not1  g2726(.din(new_new_n3646__), .dout(n10010));
  buf1  g2727(.din(new_new_n5447__), .dout(n10013));
  buf1  g2728(.din(new_new_n5451__), .dout(n10016));
  buf1  g2729(.din(new_new_n3690__), .dout(n10019));
  buf1  g2730(.din(new_new_n3692__), .dout(n10022));
  not1  g2731(.din(new_new_n3693__), .dout(n10025));
  buf1  g2732(.din(n9773), .dout(n10028));
  buf1  g2733(.din(n9776), .dout(n10031));
  buf1  g2734(.din(new_new_n3695__), .dout(n10034));
  not1  g2735(.din(new_new_n5470__), .dout(n10037));
  buf1  g2736(.din(n9785), .dout(n10040));
  buf1  g2737(.din(new_new_n3709__), .dout(n10043));
  buf1  g2738(.din(n9800), .dout(n10046));
  buf1  g2739(.din(new_new_n3724__), .dout(n10049));
  buf1  g2740(.din(n9803), .dout(n10052));
  buf1  g2741(.din(new_new_n3733__), .dout(n10055));
  buf1  g2742(.din(new_new_n5482__), .dout(n10058));
  buf1  g2743(.din(n10058), .dout(n10061));
  buf1  g2744(.din(n9812), .dout(n10064));
  buf1  g2745(.din(n9815), .dout(n10067));
  buf1  g2746(.din(n9818), .dout(n10070));
  buf1  g2747(.din(n9821), .dout(n10073));
  buf1  g2748(.din(n9824), .dout(n10076));
  buf1  g2749(.din(n9827), .dout(n10079));
  buf1  g2750(.din(new_new_n3736__), .dout(n10082));
  not1  g2751(.din(new_new_n5508__), .dout(n10085));
  buf1  g2752(.din(n10085), .dout(n10088));
  not1  g2753(.din(new_new_n5510__), .dout(n10091));
  buf1  g2754(.din(n10091), .dout(n10094));
  not1  g2755(.din(new_new_n5511__), .dout(n10097));
  buf1  g2756(.din(n10097), .dout(n10100));
  not1  g2757(.din(new_new_n5513__), .dout(n10103));
  buf1  g2758(.din(n10103), .dout(n10106));
  not1  g2759(.din(new_new_n5514__), .dout(n10109));
  buf1  g2760(.din(n10109), .dout(n10112));
  not1  g2761(.din(new_new_n5519__), .dout(n10115));
  buf1  g2762(.din(n10115), .dout(n10118));
  not1  g2763(.din(new_new_n5521__), .dout(n10121));
  buf1  g2764(.din(n10121), .dout(n10124));
  not1  g2765(.din(new_new_n5522__), .dout(n10127));
  buf1  g2766(.din(n10127), .dout(n10130));
  not1  g2767(.din(new_new_n5524__), .dout(n10133));
  buf1  g2768(.din(n10133), .dout(n10136));
  not1  g2769(.din(new_new_n5525__), .dout(n10139));
  buf1  g2770(.din(n10139), .dout(n10142));
  not1  g2771(.din(new_new_n5530__), .dout(n10145));
  buf1  g2772(.din(n10145), .dout(n10148));
  not1  g2773(.din(new_new_n5532__), .dout(n10151));
  buf1  g2774(.din(n10151), .dout(n10154));
  not1  g2775(.din(new_new_n5533__), .dout(n10157));
  buf1  g2776(.din(n10157), .dout(n10160));
  not1  g2777(.din(new_new_n5535__), .dout(n10163));
  buf1  g2778(.din(n10163), .dout(n10166));
  not1  g2779(.din(new_new_n5536__), .dout(n10169));
  buf1  g2780(.din(n10169), .dout(n10172));
  not1  g2781(.din(new_new_n5541__), .dout(n10175));
  buf1  g2782(.din(n10175), .dout(n10178));
  not1  g2783(.din(new_new_n5543__), .dout(n10181));
  buf1  g2784(.din(n10181), .dout(n10184));
  not1  g2785(.din(new_new_n5544__), .dout(n10187));
  buf1  g2786(.din(n10187), .dout(n10190));
  not1  g2787(.din(new_new_n5546__), .dout(n10193));
  buf1  g2788(.din(n10193), .dout(n10196));
  not1  g2789(.din(new_new_n5547__), .dout(n10199));
  buf1  g2790(.din(n10199), .dout(n10202));
  buf1  g2791(.din(new_new_n5552__), .dout(n10205));
  buf1  g2792(.din(n10205), .dout(n10208));
  buf1  g2793(.din(new_new_n5554__), .dout(n10211));
  buf1  g2794(.din(n10211), .dout(n10214));
  buf1  g2795(.din(new_new_n5555__), .dout(n10217));
  buf1  g2796(.din(n10217), .dout(n10220));
  buf1  g2797(.din(new_new_n5557__), .dout(n10223));
  buf1  g2798(.din(n10223), .dout(n10226));
  buf1  g2799(.din(new_new_n5558__), .dout(n10229));
  buf1  g2800(.din(n10229), .dout(n10232));
  buf1  g2801(.din(new_new_n5563__), .dout(n10235));
  buf1  g2802(.din(n10235), .dout(n10238));
  buf1  g2803(.din(new_new_n5565__), .dout(n10241));
  buf1  g2804(.din(n10241), .dout(n10244));
  buf1  g2805(.din(new_new_n5566__), .dout(n10247));
  buf1  g2806(.din(n10247), .dout(n10250));
  buf1  g2807(.din(new_new_n5568__), .dout(n10253));
  buf1  g2808(.din(n10253), .dout(n10256));
  buf1  g2809(.din(new_new_n5569__), .dout(n10259));
  buf1  g2810(.din(n10259), .dout(n10262));
  not1  g2811(.din(new_new_n5574__), .dout(n10265));
  buf1  g2812(.din(n10265), .dout(n10268));
  not1  g2813(.din(new_new_n5576__), .dout(n10271));
  buf1  g2814(.din(n10271), .dout(n10274));
  not1  g2815(.din(new_new_n5577__), .dout(n10277));
  buf1  g2816(.din(n10277), .dout(n10280));
  not1  g2817(.din(new_new_n5579__), .dout(n10283));
  buf1  g2818(.din(n10283), .dout(n10286));
  not1  g2819(.din(new_new_n5580__), .dout(n10289));
  buf1  g2820(.din(n10289), .dout(n10292));
  not1  g2821(.din(new_new_n5585__), .dout(n10295));
  buf1  g2822(.din(n10295), .dout(n10298));
  not1  g2823(.din(new_new_n5587__), .dout(n10301));
  buf1  g2824(.din(n10301), .dout(n10304));
  not1  g2825(.din(new_new_n5588__), .dout(n10307));
  buf1  g2826(.din(n10307), .dout(n10310));
  not1  g2827(.din(new_new_n5590__), .dout(n10313));
  buf1  g2828(.din(n10313), .dout(n10316));
  not1  g2829(.din(new_new_n5591__), .dout(n10319));
  buf1  g2830(.din(n10319), .dout(n10322));
  not1  g2831(.din(new_new_n5469__), .dout(n10325));
  not1  g2832(.din(new_new_n5472__), .dout(n10328));
  buf1  g2833(.din(new_new_n5601__), .dout(n10331));
  not1  g2834(.din(new_new_n5465__), .dout(n10334));
  buf1  g2835(.din(n9878), .dout(n10337));
  buf1  g2836(.din(new_new_n5493__), .dout(n10340));
  buf1  g2837(.din(new_new_n5455__), .dout(n10343));
  buf1  g2838(.din(new_new_n5603__), .dout(n10346));
  buf1  g2839(.din(new_new_n5605__), .dout(n10349));
  buf1  g2840(.din(n9884), .dout(n10352));
  buf1  g2841(.din(n9887), .dout(n10355));
  buf1  g2842(.din(n9890), .dout(n10358));
  buf1  g2843(.din(n9605), .dout(n10361));
  not1  g2844(.din(new_new_n3772__), .dout(n10364));
  not1  g2845(.din(new_new_n3774__), .dout(n10367));
  not1  g2846(.din(new_new_n3775__), .dout(n10370));
  not1  g2847(.din(new_new_n3776__), .dout(n10373));
  buf1  g2848(.din(new_new_n5606__), .dout(n10376));
  buf1  g2849(.din(new_new_n5475__), .dout(n10379));
  buf1  g2850(.din(new_new_n5607__), .dout(n10382));
  buf1  g2851(.din(n10382), .dout(n10385));
  buf1  g2852(.din(n9992), .dout(n10388));
  buf1  g2853(.din(n9710), .dout(n10391));
  buf1  g2854(.din(new_new_n5446__), .dout(n10394));
  not1  g2855(.din(new_new_n3793__), .dout(n10397));
  not1  g2856(.din(new_new_n3794__), .dout(n10400));
  buf1  g2857(.din(new_new_n5608__), .dout(n10403));
  buf1  g2858(.din(new_new_n5478__), .dout(n10406));
  buf1  g2859(.din(new_new_n5477__), .dout(n10409));
  buf1  g2860(.din(new_new_n5473__), .dout(n10412));
  buf1  g2861(.din(new_new_n5609__), .dout(n10415));
  buf1  g2862(.din(n10415), .dout(n10418));
  not1  g2863(.din(new_new_n3807__), .dout(n10421));
  not1  g2864(.din(new_new_n5496__), .dout(n10424));
  not1  g2865(.din(new_new_n5471__), .dout(n10427));
  buf1  g2866(.din(n10331), .dout(n10430));
  buf1  g2867(.din(new_new_n5592__), .dout(n10433));
  buf1  g2868(.din(n10340), .dout(n10436));
  buf1  g2869(.din(n10346), .dout(n10439));
  buf1  g2870(.din(n10349), .dout(n10442));
  buf1  g2871(.din(new_new_n5463__), .dout(n10445));
  buf1  g2872(.din(new_new_n5596__), .dout(n10448));
  buf1  g2873(.din(new_new_n5599__), .dout(n10451));
  buf1  g2874(.din(new_new_n1143__), .dout(n10454));
  buf1  g2875(.din(new_new_n1157__), .dout(n10457));
  buf1  g2876(.din(new_new_n1187__), .dout(n10460));
  buf1  g2877(.din(new_new_n1195__), .dout(n10463));
  buf1  g2878(.din(new_new_n1197__), .dout(n10466));
  buf1  g2879(.din(new_new_n1199__), .dout(n10469));
  buf1  g2880(.din(new_new_n1205__), .dout(n10472));
  buf1  g2881(.din(new_new_n1207__), .dout(n10475));
  buf1  g2882(.din(new_new_n1209__), .dout(n10478));
  buf1  g2883(.din(new_new_n3808__), .dout(n10481));
  buf1  g2884(.din(new_new_n1149__), .dout(n10484));
  buf1  g2885(.din(new_new_n1189__), .dout(n10487));
  buf1  g2886(.din(new_new_n3809__), .dout(n10490));
  buf1  g2887(.din(n10376), .dout(n10493));
  buf1  g2888(.din(new_new_n5474__), .dout(n10496));
  buf1  g2889(.din(new_new_n3810__), .dout(n10499));
  buf1  g2890(.din(new_new_n1151__), .dout(n10502));
  buf1  g2891(.din(new_new_n1191__), .dout(n10505));
  buf1  g2892(.din(new_new_n1193__), .dout(n10508));
  buf1  g2893(.din(n10403), .dout(n10511));
  buf1  g2894(.din(new_new_n3811__), .dout(n10514));
  buf1  g2895(.din(new_new_n5476__), .dout(n10517));
  buf1  g2896(.din(new_new_n5602__), .dout(n10520));
  buf1  g2897(.din(new_new_n5604__), .dout(n10523));
  buf1  g2898(.din(n10445), .dout(n10526));
  buf1  g2899(.din(n10448), .dout(n10529));
  buf1  g2900(.din(n10451), .dout(n10532));
  buf1  g2901(.din(new_new_n1378__), .dout(new_new_n4363__));
  buf1  g2902(.din(new_new_n1377__), .dout(new_new_n4364__));
  buf1  g2903(.din(new_new_n1382__), .dout(new_new_n4365__));
  buf1  g2904(.din(new_new_n1381__), .dout(new_new_n4366__));
  buf1  g2905(.din(new_new_n2296__), .dout(new_new_n4367__));
  buf1  g2906(.din(new_new_n1298__), .dout(new_new_n4368__));
  buf1  g2907(.din(new_new_n1294__), .dout(new_new_n4369__));
  buf1  g2908(.din(new_new_n1292__), .dout(new_new_n4370__));
  buf1  g2909(.din(new_new_n2300__), .dout(new_new_n4371__));
  buf1  g2910(.din(new_new_n2301__), .dout(new_new_n4372__));
  buf1  g2911(.din(new_new_n2295__), .dout(new_new_n4373__));
  buf1  g2912(.din(new_new_n1366__), .dout(new_new_n4374__));
  buf1  g2913(.din(new_new_n1363__), .dout(new_new_n4375__));
  buf1  g2914(.din(new_new_n1365__), .dout(new_new_n4376__));
  buf1  g2915(.din(new_new_n1364__), .dout(new_new_n4377__));
  buf1  g2916(.din(new_new_n1357__), .dout(new_new_n4378__));
  buf1  g2917(.din(new_new_n1329__), .dout(new_new_n4379__));
  buf1  g2918(.din(new_new_n2349__), .dout(new_new_n4380__));
  buf1  g2919(.din(new_new_n2352__), .dout(new_new_n4381__));
  buf1  g2920(.din(new_new_n1746__), .dout(new_new_n4382__));
  buf1  g2921(.din(new_new_n1743__), .dout(new_new_n4383__));
  buf1  g2922(.din(new_new_n1745__), .dout(new_new_n4384__));
  buf1  g2923(.din(new_new_n1744__), .dout(new_new_n4385__));
  buf1  g2924(.din(new_new_n1369__), .dout(new_new_n4386__));
  buf1  g2925(.din(new_new_n1367__), .dout(new_new_n4387__));
  buf1  g2926(.din(new_new_n1370__), .dout(new_new_n4388__));
  buf1  g2927(.din(new_new_n1368__), .dout(new_new_n4389__));
  buf1  g2928(.din(new_new_n2389__), .dout(new_new_n4390__));
  buf1  g2929(.din(new_new_n2392__), .dout(new_new_n4391__));
  buf1  g2930(.din(new_new_n2395__), .dout(new_new_n4392__));
  buf1  g2931(.din(new_new_n2398__), .dout(new_new_n4393__));
  buf1  g2932(.din(new_new_n2404__), .dout(new_new_n4394__));
  buf1  g2933(.din(new_new_n2406__), .dout(new_new_n4395__));
  buf1  g2934(.din(new_new_n2412__), .dout(new_new_n4396__));
  buf1  g2935(.din(new_new_n2410__), .dout(new_new_n4397__));
  buf1  g2936(.din(new_new_n2420__), .dout(new_new_n4398__));
  buf1  g2937(.din(new_new_n2417__), .dout(new_new_n4399__));
  buf1  g2938(.din(new_new_n2419__), .dout(new_new_n4400__));
  buf1  g2939(.din(new_new_n2418__), .dout(new_new_n4401__));
  buf1  g2940(.din(new_new_n1687__), .dout(new_new_n4402__));
  buf1  g2941(.din(new_new_n1686__), .dout(new_new_n4403__));
  buf1  g2942(.din(new_new_n1688__), .dout(new_new_n4404__));
  buf1  g2943(.din(new_new_n1685__), .dout(new_new_n4405__));
  buf1  g2944(.din(new_new_n2438__), .dout(new_new_n4406__));
  buf1  g2945(.din(new_new_n2432__), .dout(new_new_n4407__));
  buf1  g2946(.din(new_new_n4407__), .dout(new_new_n4408__));
  buf1  g2947(.din(new_new_n4407__), .dout(new_new_n4409__));
  buf1  g2948(.din(new_new_n2437__), .dout(new_new_n4410__));
  buf1  g2949(.din(new_new_n2431__), .dout(new_new_n4411__));
  buf1  g2950(.din(new_new_n4411__), .dout(new_new_n4412__));
  buf1  g2951(.din(new_new_n4411__), .dout(new_new_n4413__));
  buf1  g2952(.din(new_new_n2439__), .dout(new_new_n4414__));
  buf1  g2953(.din(new_new_n4414__), .dout(new_new_n4415__));
  buf1  g2954(.din(new_new_n4414__), .dout(new_new_n4416__));
  buf1  g2955(.din(new_new_n2440__), .dout(new_new_n4417__));
  buf1  g2956(.din(new_new_n4417__), .dout(new_new_n4418__));
  buf1  g2957(.din(new_new_n4417__), .dout(new_new_n4419__));
  buf1  g2958(.din(new_new_n1793__), .dout(new_new_n4420__));
  buf1  g2959(.din(new_new_n1792__), .dout(new_new_n4421__));
  buf1  g2960(.din(new_new_n1794__), .dout(new_new_n4422__));
  buf1  g2961(.din(new_new_n1791__), .dout(new_new_n4423__));
  buf1  g2962(.din(new_new_n2449__), .dout(new_new_n4424__));
  buf1  g2963(.din(new_new_n2450__), .dout(new_new_n4425__));
  buf1  g2964(.din(new_new_n1777__), .dout(new_new_n4426__));
  buf1  g2965(.din(new_new_n1773__), .dout(new_new_n4427__));
  buf1  g2966(.din(new_new_n1778__), .dout(new_new_n4428__));
  buf1  g2967(.din(new_new_n1774__), .dout(new_new_n4429__));
  buf1  g2968(.din(new_new_n2459__), .dout(new_new_n4430__));
  buf1  g2969(.din(new_new_n2460__), .dout(new_new_n4431__));
  buf1  g2970(.din(new_new_n2426__), .dout(new_new_n4432__));
  buf1  g2971(.din(new_new_n2425__), .dout(new_new_n4433__));
  buf1  g2972(.din(new_new_n1768__), .dout(new_new_n4434__));
  buf1  g2973(.din(new_new_n1765__), .dout(new_new_n4435__));
  buf1  g2974(.din(new_new_n1767__), .dout(new_new_n4436__));
  buf1  g2975(.din(new_new_n1766__), .dout(new_new_n4437__));
  buf1  g2976(.din(new_new_n2483__), .dout(new_new_n4438__));
  buf1  g2977(.din(new_new_n2482__), .dout(new_new_n4439__));
  buf1  g2978(.din(new_new_n1635__), .dout(new_new_n4440__));
  buf1  g2979(.din(new_new_n1750__), .dout(new_new_n4441__));
  buf1  g2980(.din(new_new_n4441__), .dout(new_new_n4442__));
  buf1  g2981(.din(new_new_n1748__), .dout(new_new_n4443__));
  buf1  g2982(.din(new_new_n1749__), .dout(new_new_n4444__));
  buf1  g2983(.din(new_new_n4444__), .dout(new_new_n4445__));
  buf1  g2984(.din(new_new_n4444__), .dout(new_new_n4446__));
  buf1  g2985(.din(new_new_n1747__), .dout(new_new_n4447__));
  buf1  g2986(.din(new_new_n4447__), .dout(new_new_n4448__));
  buf1  g2987(.din(new_new_n1751__), .dout(new_new_n4449__));
  buf1  g2988(.din(new_new_n1449__), .dout(new_new_n4450__));
  buf1  g2989(.din(new_new_n4450__), .dout(new_new_n4451__));
  buf1  g2990(.din(new_new_n1450__), .dout(new_new_n4452__));
  buf1  g2991(.din(new_new_n4452__), .dout(new_new_n4453__));
  buf1  g2992(.din(new_new_n1470__), .dout(new_new_n4454__));
  buf1  g2993(.din(new_new_n1468__), .dout(new_new_n4455__));
  buf1  g2994(.din(new_new_n1469__), .dout(new_new_n4456__));
  buf1  g2995(.din(new_new_n1467__), .dout(new_new_n4457__));
  buf1  g2996(.din(new_new_n4457__), .dout(new_new_n4458__));
  buf1  g2997(.din(new_new_n1403__), .dout(new_new_n4459__));
  buf1  g2998(.din(new_new_n2523__), .dout(new_new_n4460__));
  buf1  g2999(.din(new_new_n4460__), .dout(new_new_n4461__));
  buf1  g3000(.din(new_new_n2517__), .dout(new_new_n4462__));
  buf1  g3001(.din(new_new_n2529__), .dout(new_new_n4463__));
  buf1  g3002(.din(new_new_n4463__), .dout(new_new_n4464__));
  buf1  g3003(.din(new_new_n2522__), .dout(new_new_n4465__));
  buf1  g3004(.din(new_new_n4465__), .dout(new_new_n4466__));
  buf1  g3005(.din(new_new_n4466__), .dout(new_new_n4467__));
  buf1  g3006(.din(new_new_n4466__), .dout(new_new_n4468__));
  buf1  g3007(.din(new_new_n4465__), .dout(new_new_n4469__));
  buf1  g3008(.din(new_new_n4469__), .dout(new_new_n4470__));
  buf1  g3009(.din(new_new_n1926__), .dout(new_new_n4471__));
  buf1  g3010(.din(new_new_n1924__), .dout(new_new_n4472__));
  buf1  g3011(.din(new_new_n1925__), .dout(new_new_n4473__));
  buf1  g3012(.din(new_new_n1923__), .dout(new_new_n4474__));
  buf1  g3013(.din(new_new_n2536__), .dout(new_new_n4475__));
  buf1  g3014(.din(new_new_n4475__), .dout(new_new_n4476__));
  buf1  g3015(.din(new_new_n2541__), .dout(new_new_n4477__));
  buf1  g3016(.din(new_new_n1862__), .dout(new_new_n4478__));
  buf1  g3017(.din(new_new_n4478__), .dout(new_new_n4479__));
  buf1  g3018(.din(new_new_n1885__), .dout(new_new_n4480__));
  buf1  g3019(.din(new_new_n4480__), .dout(new_new_n4481__));
  buf1  g3020(.din(new_new_n4481__), .dout(new_new_n4482__));
  buf1  g3021(.din(new_new_n4481__), .dout(new_new_n4483__));
  buf1  g3022(.din(new_new_n4480__), .dout(new_new_n4484__));
  buf1  g3023(.din(new_new_n1753__), .dout(new_new_n4485__));
  buf1  g3024(.din(new_new_n4485__), .dout(new_new_n4486__));
  buf1  g3025(.din(new_new_n4486__), .dout(new_new_n4487__));
  buf1  g3026(.din(new_new_n4486__), .dout(new_new_n4488__));
  buf1  g3027(.din(new_new_n4485__), .dout(new_new_n4489__));
  buf1  g3028(.din(new_new_n1452__), .dout(new_new_n4490__));
  buf1  g3029(.din(new_new_n4490__), .dout(new_new_n4491__));
  buf1  g3030(.din(new_new_n4491__), .dout(new_new_n4492__));
  buf1  g3031(.din(new_new_n4491__), .dout(new_new_n4493__));
  buf1  g3032(.din(new_new_n4490__), .dout(new_new_n4494__));
  buf1  g3033(.din(new_new_n1476__), .dout(new_new_n4495__));
  buf1  g3034(.din(new_new_n4495__), .dout(new_new_n4496__));
  buf1  g3035(.din(new_new_n4496__), .dout(new_new_n4497__));
  buf1  g3036(.din(new_new_n4496__), .dout(new_new_n4498__));
  buf1  g3037(.din(new_new_n4495__), .dout(new_new_n4499__));
  buf1  g3038(.din(new_new_n1868__), .dout(new_new_n4500__));
  buf1  g3039(.din(new_new_n4500__), .dout(new_new_n4501__));
  buf1  g3040(.din(new_new_n4501__), .dout(new_new_n4502__));
  buf1  g3041(.din(new_new_n4500__), .dout(new_new_n4503__));
  buf1  g3042(.din(new_new_n1866__), .dout(new_new_n4504__));
  buf1  g3043(.din(new_new_n4504__), .dout(new_new_n4505__));
  buf1  g3044(.din(new_new_n4505__), .dout(new_new_n4506__));
  buf1  g3045(.din(new_new_n4504__), .dout(new_new_n4507__));
  buf1  g3046(.din(new_new_n1864__), .dout(new_new_n4508__));
  buf1  g3047(.din(new_new_n4508__), .dout(new_new_n4509__));
  buf1  g3048(.din(new_new_n4508__), .dout(new_new_n4510__));
  buf1  g3049(.din(new_new_n1880__), .dout(new_new_n4511__));
  buf1  g3050(.din(new_new_n4511__), .dout(new_new_n4512__));
  buf1  g3051(.din(new_new_n4512__), .dout(new_new_n4513__));
  buf1  g3052(.din(new_new_n4513__), .dout(new_new_n4514__));
  buf1  g3053(.din(new_new_n4512__), .dout(new_new_n4515__));
  buf1  g3054(.din(new_new_n4511__), .dout(new_new_n4516__));
  buf1  g3055(.din(new_new_n4516__), .dout(new_new_n4517__));
  buf1  g3056(.din(new_new_n4516__), .dout(new_new_n4518__));
  buf1  g3057(.din(new_new_n1456__), .dout(new_new_n4519__));
  buf1  g3058(.din(new_new_n4519__), .dout(new_new_n4520__));
  buf1  g3059(.din(new_new_n4519__), .dout(new_new_n4521__));
  buf1  g3060(.din(new_new_n1895__), .dout(new_new_n4522__));
  buf1  g3061(.din(new_new_n4522__), .dout(new_new_n4523__));
  buf1  g3062(.din(new_new_n4523__), .dout(new_new_n4524__));
  buf1  g3063(.din(new_new_n4523__), .dout(new_new_n4525__));
  buf1  g3064(.din(new_new_n4522__), .dout(new_new_n4526__));
  buf1  g3065(.din(new_new_n1893__), .dout(new_new_n4527__));
  buf1  g3066(.din(new_new_n4527__), .dout(new_new_n4528__));
  buf1  g3067(.din(new_new_n4528__), .dout(new_new_n4529__));
  buf1  g3068(.din(new_new_n4528__), .dout(new_new_n4530__));
  buf1  g3069(.din(new_new_n4527__), .dout(new_new_n4531__));
  buf1  g3070(.din(new_new_n1889__), .dout(new_new_n4532__));
  buf1  g3071(.din(new_new_n4532__), .dout(new_new_n4533__));
  buf1  g3072(.din(new_new_n4533__), .dout(new_new_n4534__));
  buf1  g3073(.din(new_new_n4533__), .dout(new_new_n4535__));
  buf1  g3074(.din(new_new_n4532__), .dout(new_new_n4536__));
  buf1  g3075(.din(new_new_n4536__), .dout(new_new_n4537__));
  buf1  g3076(.din(new_new_n1883__), .dout(new_new_n4538__));
  buf1  g3077(.din(new_new_n4538__), .dout(new_new_n4539__));
  buf1  g3078(.din(new_new_n4539__), .dout(new_new_n4540__));
  buf1  g3079(.din(new_new_n4539__), .dout(new_new_n4541__));
  buf1  g3080(.din(new_new_n4538__), .dout(new_new_n4542__));
  buf1  g3081(.din(new_new_n1897__), .dout(new_new_n4543__));
  buf1  g3082(.din(new_new_n4543__), .dout(new_new_n4544__));
  buf1  g3083(.din(new_new_n4544__), .dout(new_new_n4545__));
  buf1  g3084(.din(new_new_n4544__), .dout(new_new_n4546__));
  buf1  g3085(.din(new_new_n4543__), .dout(new_new_n4547__));
  buf1  g3086(.din(new_new_n4547__), .dout(new_new_n4548__));
  buf1  g3087(.din(new_new_n1444__), .dout(new_new_n4549__));
  buf1  g3088(.din(new_new_n4549__), .dout(new_new_n4550__));
  buf1  g3089(.din(new_new_n4550__), .dout(new_new_n4551__));
  buf1  g3090(.din(new_new_n4550__), .dout(new_new_n4552__));
  buf1  g3091(.din(new_new_n4549__), .dout(new_new_n4553__));
  buf1  g3092(.din(new_new_n1446__), .dout(new_new_n4554__));
  buf1  g3093(.din(new_new_n4554__), .dout(new_new_n4555__));
  buf1  g3094(.din(new_new_n4555__), .dout(new_new_n4556__));
  buf1  g3095(.din(new_new_n4554__), .dout(new_new_n4557__));
  buf1  g3096(.din(new_new_n1879__), .dout(new_new_n4558__));
  buf1  g3097(.din(new_new_n4558__), .dout(new_new_n4559__));
  buf1  g3098(.din(new_new_n4559__), .dout(new_new_n4560__));
  buf1  g3099(.din(new_new_n4560__), .dout(new_new_n4561__));
  buf1  g3100(.din(new_new_n4559__), .dout(new_new_n4562__));
  buf1  g3101(.din(new_new_n4558__), .dout(new_new_n4563__));
  buf1  g3102(.din(new_new_n4563__), .dout(new_new_n4564__));
  buf1  g3103(.din(new_new_n4563__), .dout(new_new_n4565__));
  buf1  g3104(.din(new_new_n2581__), .dout(new_new_n4566__));
  buf1  g3105(.din(new_new_n4566__), .dout(new_new_n4567__));
  buf1  g3106(.din(new_new_n4567__), .dout(new_new_n4568__));
  buf1  g3107(.din(new_new_n4567__), .dout(new_new_n4569__));
  buf1  g3108(.din(new_new_n4566__), .dout(new_new_n4570__));
  buf1  g3109(.din(new_new_n4570__), .dout(new_new_n4571__));
  buf1  g3110(.din(new_new_n1397__), .dout(new_new_n4572__));
  buf1  g3111(.din(new_new_n4572__), .dout(new_new_n4573__));
  buf1  g3112(.din(new_new_n4572__), .dout(new_new_n4574__));
  buf1  g3113(.din(new_new_n1398__), .dout(new_new_n4575__));
  buf1  g3114(.din(new_new_n4575__), .dout(new_new_n4576__));
  buf1  g3115(.din(new_new_n4575__), .dout(new_new_n4577__));
  buf1  g3116(.din(new_new_n2586__), .dout(new_new_n4578__));
  buf1  g3117(.din(new_new_n4578__), .dout(new_new_n4579__));
  buf1  g3118(.din(new_new_n4578__), .dout(new_new_n4580__));
  buf1  g3119(.din(new_new_n2580__), .dout(new_new_n4581__));
  buf1  g3120(.din(new_new_n4581__), .dout(new_new_n4582__));
  buf1  g3121(.din(new_new_n4581__), .dout(new_new_n4583__));
  buf1  g3122(.din(new_new_n2589__), .dout(new_new_n4584__));
  buf1  g3123(.din(new_new_n4584__), .dout(new_new_n4585__));
  buf1  g3124(.din(new_new_n4584__), .dout(new_new_n4586__));
  buf1  g3125(.din(new_new_n2504__), .dout(new_new_n4587__));
  buf1  g3126(.din(new_new_n4587__), .dout(new_new_n4588__));
  buf1  g3127(.din(new_new_n4588__), .dout(new_new_n4589__));
  buf1  g3128(.din(new_new_n4588__), .dout(new_new_n4590__));
  buf1  g3129(.din(new_new_n4587__), .dout(new_new_n4591__));
  buf1  g3130(.din(new_new_n4591__), .dout(new_new_n4592__));
  buf1  g3131(.din(new_new_n4591__), .dout(new_new_n4593__));
  buf1  g3132(.din(new_new_n2505__), .dout(new_new_n4594__));
  buf1  g3133(.din(new_new_n4594__), .dout(new_new_n4595__));
  buf1  g3134(.din(new_new_n2594__), .dout(new_new_n4596__));
  buf1  g3135(.din(new_new_n4596__), .dout(new_new_n4597__));
  buf1  g3136(.din(new_new_n4597__), .dout(new_new_n4598__));
  buf1  g3137(.din(new_new_n4597__), .dout(new_new_n4599__));
  buf1  g3138(.din(new_new_n4596__), .dout(new_new_n4600__));
  buf1  g3139(.din(new_new_n1949__), .dout(new_new_n4601__));
  buf1  g3140(.din(new_new_n4601__), .dout(new_new_n4602__));
  buf1  g3141(.din(new_new_n2516__), .dout(new_new_n4603__));
  buf1  g3142(.din(new_new_n1950__), .dout(new_new_n4604__));
  buf1  g3143(.din(new_new_n4604__), .dout(new_new_n4605__));
  buf1  g3144(.din(new_new_n1661__), .dout(new_new_n4606__));
  buf1  g3145(.din(new_new_n4606__), .dout(new_new_n4607__));
  buf1  g3146(.din(new_new_n1662__), .dout(new_new_n4608__));
  buf1  g3147(.din(new_new_n2607__), .dout(new_new_n4609__));
  buf1  g3148(.din(new_new_n1881__), .dout(new_new_n4610__));
  buf1  g3149(.din(new_new_n4610__), .dout(new_new_n4611__));
  buf1  g3150(.din(new_new_n4611__), .dout(new_new_n4612__));
  buf1  g3151(.din(new_new_n4611__), .dout(new_new_n4613__));
  buf1  g3152(.din(new_new_n4610__), .dout(new_new_n4614__));
  buf1  g3153(.din(new_new_n1872__), .dout(new_new_n4615__));
  buf1  g3154(.din(new_new_n1870__), .dout(new_new_n4616__));
  buf1  g3155(.din(new_new_n4616__), .dout(new_new_n4617__));
  buf1  g3156(.din(new_new_n2655__), .dout(new_new_n4618__));
  buf1  g3157(.din(new_new_n4618__), .dout(new_new_n4619__));
  buf1  g3158(.din(new_new_n1946__), .dout(new_new_n4620__));
  buf1  g3159(.din(new_new_n1945__), .dout(new_new_n4621__));
  buf1  g3160(.din(new_new_n2658__), .dout(new_new_n4622__));
  buf1  g3161(.din(new_new_n4622__), .dout(new_new_n4623__));
  buf1  g3162(.din(new_new_n2496__), .dout(new_new_n4624__));
  buf1  g3163(.din(new_new_n2662__), .dout(new_new_n4625__));
  buf1  g3164(.din(new_new_n4625__), .dout(new_new_n4626__));
  buf1  g3165(.din(new_new_n2659__), .dout(new_new_n4627__));
  buf1  g3166(.din(new_new_n4627__), .dout(new_new_n4628__));
  buf1  g3167(.din(new_new_n2661__), .dout(new_new_n4629__));
  buf1  g3168(.din(new_new_n4629__), .dout(new_new_n4630__));
  buf1  g3169(.din(new_new_n2663__), .dout(new_new_n4631__));
  buf1  g3170(.din(new_new_n2656__), .dout(new_new_n4632__));
  buf1  g3171(.din(new_new_n4632__), .dout(new_new_n4633__));
  buf1  g3172(.din(new_new_n2668__), .dout(new_new_n4634__));
  buf1  g3173(.din(new_new_n1894__), .dout(new_new_n4635__));
  buf1  g3174(.din(new_new_n1896__), .dout(new_new_n4636__));
  buf1  g3175(.din(new_new_n1882__), .dout(new_new_n4637__));
  buf1  g3176(.din(new_new_n1886__), .dout(new_new_n4638__));
  buf1  g3177(.din(new_new_n1754__), .dout(new_new_n4639__));
  buf1  g3178(.din(new_new_n1451__), .dout(new_new_n4640__));
  buf1  g3179(.din(new_new_n1873__), .dout(new_new_n4641__));
  buf1  g3180(.din(new_new_n1884__), .dout(new_new_n4642__));
  buf1  g3181(.din(new_new_n1443__), .dout(new_new_n4643__));
  buf1  g3182(.din(new_new_n1445__), .dout(new_new_n4644__));
  buf1  g3183(.din(new_new_n1455__), .dout(new_new_n4645__));
  buf1  g3184(.din(new_new_n1869__), .dout(new_new_n4646__));
  buf1  g3185(.din(new_new_n1871__), .dout(new_new_n4647__));
  buf1  g3186(.din(new_new_n2499__), .dout(new_new_n4648__));
  buf1  g3187(.din(new_new_n2664__), .dout(new_new_n4649__));
  buf1  g3188(.din(new_new_n2669__), .dout(new_new_n4650__));
  buf1  g3189(.din(new_new_n2593__), .dout(new_new_n4651__));
  buf1  g3190(.din(new_new_n1639__), .dout(new_new_n4652__));
  buf1  g3191(.din(new_new_n1947__), .dout(new_new_n4653__));
  buf1  g3192(.din(new_new_n2493__), .dout(new_new_n4654__));
  buf1  g3193(.din(new_new_n1425__), .dout(new_new_n4655__));
  buf1  g3194(.din(new_new_n1956__), .dout(new_new_n4656__));
  buf1  g3195(.din(new_new_n4656__), .dout(new_new_n4657__));
  buf1  g3196(.din(new_new_n1955__), .dout(new_new_n4658__));
  buf1  g3197(.din(new_new_n4658__), .dout(new_new_n4659__));
  buf1  g3198(.din(new_new_n1723__), .dout(new_new_n4660__));
  buf1  g3199(.din(new_new_n2834__), .dout(new_new_n4661__));
  buf1  g3200(.din(new_new_n1725__), .dout(new_new_n4662__));
  buf1  g3201(.din(new_new_n2835__), .dout(new_new_n4663__));
  buf1  g3202(.din(new_new_n2837__), .dout(new_new_n4664__));
  buf1  g3203(.din(new_new_n4664__), .dout(new_new_n4665__));
  buf1  g3204(.din(new_new_n4665__), .dout(new_new_n4666__));
  buf1  g3205(.din(new_new_n4665__), .dout(new_new_n4667__));
  buf1  g3206(.din(new_new_n4664__), .dout(new_new_n4668__));
  buf1  g3207(.din(new_new_n4668__), .dout(new_new_n4669__));
  buf1  g3208(.din(new_new_n4668__), .dout(new_new_n4670__));
  buf1  g3209(.din(new_new_n2511__), .dout(new_new_n4671__));
  buf1  g3210(.din(new_new_n2836__), .dout(new_new_n4672__));
  buf1  g3211(.din(new_new_n4672__), .dout(new_new_n4673__));
  buf1  g3212(.din(new_new_n4673__), .dout(new_new_n4674__));
  buf1  g3213(.din(new_new_n4673__), .dout(new_new_n4675__));
  buf1  g3214(.din(new_new_n4672__), .dout(new_new_n4676__));
  buf1  g3215(.din(new_new_n4676__), .dout(new_new_n4677__));
  buf1  g3216(.din(new_new_n4676__), .dout(new_new_n4678__));
  buf1  g3217(.din(new_new_n2155__), .dout(new_new_n4679__));
  buf1  g3218(.din(new_new_n4679__), .dout(new_new_n4680__));
  buf1  g3219(.din(new_new_n4679__), .dout(new_new_n4681__));
  buf1  g3220(.din(new_new_n2149__), .dout(new_new_n4682__));
  buf1  g3221(.din(new_new_n4682__), .dout(new_new_n4683__));
  buf1  g3222(.din(new_new_n4682__), .dout(new_new_n4684__));
  buf1  g3223(.din(new_new_n2156__), .dout(new_new_n4685__));
  buf1  g3224(.din(new_new_n4685__), .dout(new_new_n4686__));
  buf1  g3225(.din(new_new_n2150__), .dout(new_new_n4687__));
  buf1  g3226(.din(new_new_n4687__), .dout(new_new_n4688__));
  buf1  g3227(.din(new_new_n2846__), .dout(new_new_n4689__));
  buf1  g3228(.din(new_new_n4689__), .dout(new_new_n4690__));
  buf1  g3229(.din(new_new_n4689__), .dout(new_new_n4691__));
  buf1  g3230(.din(new_new_n2847__), .dout(new_new_n4692__));
  buf1  g3231(.din(new_new_n4692__), .dout(new_new_n4693__));
  buf1  g3232(.din(new_new_n1962__), .dout(new_new_n4694__));
  buf1  g3233(.din(new_new_n1919__), .dout(new_new_n4695__));
  buf1  g3234(.din(new_new_n1961__), .dout(new_new_n4696__));
  buf1  g3235(.din(new_new_n1920__), .dout(new_new_n4697__));
  buf1  g3236(.din(new_new_n2864__), .dout(new_new_n4698__));
  buf1  g3237(.din(new_new_n4698__), .dout(new_new_n4699__));
  buf1  g3238(.din(new_new_n2187__), .dout(new_new_n4700__));
  buf1  g3239(.din(new_new_n4700__), .dout(new_new_n4701__));
  buf1  g3240(.din(new_new_n1667__), .dout(new_new_n4702__));
  buf1  g3241(.din(new_new_n2188__), .dout(new_new_n4703__));
  buf1  g3242(.din(new_new_n4703__), .dout(new_new_n4704__));
  buf1  g3243(.din(new_new_n2210__), .dout(new_new_n4705__));
  buf1  g3244(.din(new_new_n2209__), .dout(new_new_n4706__));
  buf1  g3245(.din(new_new_n1669__), .dout(new_new_n4707__));
  buf1  g3246(.din(new_new_n1670__), .dout(new_new_n4708__));
  buf1  g3247(.din(new_new_n2212__), .dout(new_new_n4709__));
  buf1  g3248(.din(new_new_n2211__), .dout(new_new_n4710__));
  buf1  g3249(.din(new_new_n2190__), .dout(new_new_n4711__));
  buf1  g3250(.din(new_new_n4711__), .dout(new_new_n4712__));
  buf1  g3251(.din(new_new_n1671__), .dout(new_new_n4713__));
  buf1  g3252(.din(new_new_n2189__), .dout(new_new_n4714__));
  buf1  g3253(.din(new_new_n4714__), .dout(new_new_n4715__));
  buf1  g3254(.din(new_new_n1672__), .dout(new_new_n4716__));
  buf1  g3255(.din(new_new_n1673__), .dout(new_new_n4717__));
  buf1  g3256(.din(new_new_n1674__), .dout(new_new_n4718__));
  buf1  g3257(.din(new_new_n4718__), .dout(new_new_n4719__));
  buf1  g3258(.din(new_new_n2876__), .dout(new_new_n4720__));
  buf1  g3259(.din(new_new_n2889__), .dout(new_new_n4721__));
  buf1  g3260(.din(new_new_n4721__), .dout(new_new_n4722__));
  buf1  g3261(.din(new_new_n4722__), .dout(new_new_n4723__));
  buf1  g3262(.din(new_new_n4722__), .dout(new_new_n4724__));
  buf1  g3263(.din(new_new_n4721__), .dout(new_new_n4725__));
  buf1  g3264(.din(new_new_n2153__), .dout(new_new_n4726__));
  buf1  g3265(.din(new_new_n2890__), .dout(new_new_n4727__));
  buf1  g3266(.din(new_new_n4727__), .dout(new_new_n4728__));
  buf1  g3267(.din(new_new_n2897__), .dout(new_new_n4729__));
  buf1  g3268(.din(new_new_n4729__), .dout(new_new_n4730__));
  buf1  g3269(.din(new_new_n2615__), .dout(new_new_n4731__));
  buf1  g3270(.din(new_new_n2524__), .dout(new_new_n4732__));
  buf1  g3271(.din(new_new_n2719__), .dout(new_new_n4733__));
  buf1  g3272(.din(new_new_n2833__), .dout(new_new_n4734__));
  buf1  g3273(.din(new_new_n2531__), .dout(new_new_n4735__));
  buf1  g3274(.din(new_new_n2770__), .dout(new_new_n4736__));
  buf1  g3275(.din(new_new_n2827__), .dout(new_new_n4737__));
  buf1  g3276(.din(new_new_n2538__), .dout(new_new_n4738__));
  buf1  g3277(.din(new_new_n2595__), .dout(new_new_n4739__));
  buf1  g3278(.din(new_new_n2604__), .dout(new_new_n4740__));
  buf1  g3279(.din(new_new_n2542__), .dout(new_new_n4741__));
  buf1  g3280(.din(new_new_n2673__), .dout(new_new_n4742__));
  buf1  g3281(.din(new_new_n1538__), .dout(new_new_n4743__));
  buf1  g3282(.din(new_new_n1523__), .dout(new_new_n4744__));
  buf1  g3283(.din(new_new_n1537__), .dout(new_new_n4745__));
  buf1  g3284(.din(new_new_n1524__), .dout(new_new_n4746__));
  buf1  g3285(.din(new_new_n2919__), .dout(new_new_n4747__));
  buf1  g3286(.din(new_new_n1839__), .dout(new_new_n4748__));
  buf1  g3287(.din(new_new_n4748__), .dout(new_new_n4749__));
  buf1  g3288(.din(new_new_n1843__), .dout(new_new_n4750__));
  buf1  g3289(.din(new_new_n4750__), .dout(new_new_n4751__));
  buf1  g3290(.din(new_new_n1828__), .dout(new_new_n4752__));
  buf1  g3291(.din(new_new_n4752__), .dout(new_new_n4753__));
  buf1  g3292(.din(new_new_n1831__), .dout(new_new_n4754__));
  buf1  g3293(.din(new_new_n4754__), .dout(new_new_n4755__));
  buf1  g3294(.din(new_new_n1847__), .dout(new_new_n4756__));
  buf1  g3295(.din(new_new_n4756__), .dout(new_new_n4757__));
  buf1  g3296(.din(new_new_n1819__), .dout(new_new_n4758__));
  buf1  g3297(.din(new_new_n4758__), .dout(new_new_n4759__));
  buf1  g3298(.din(new_new_n1836__), .dout(new_new_n4760__));
  buf1  g3299(.din(new_new_n4760__), .dout(new_new_n4761__));
  buf1  g3300(.din(new_new_n1823__), .dout(new_new_n4762__));
  buf1  g3301(.din(new_new_n4762__), .dout(new_new_n4763__));
  buf1  g3302(.din(new_new_n1248__), .dout(new_new_n4764__));
  buf1  g3303(.din(new_new_n1841__), .dout(new_new_n4765__));
  buf1  g3304(.din(new_new_n4765__), .dout(new_new_n4766__));
  buf1  g3305(.din(new_new_n1845__), .dout(new_new_n4767__));
  buf1  g3306(.din(new_new_n4767__), .dout(new_new_n4768__));
  buf1  g3307(.din(new_new_n1830__), .dout(new_new_n4769__));
  buf1  g3308(.din(new_new_n4769__), .dout(new_new_n4770__));
  buf1  g3309(.din(new_new_n1833__), .dout(new_new_n4771__));
  buf1  g3310(.din(new_new_n4771__), .dout(new_new_n4772__));
  buf1  g3311(.din(new_new_n1849__), .dout(new_new_n4773__));
  buf1  g3312(.din(new_new_n4773__), .dout(new_new_n4774__));
  buf1  g3313(.din(new_new_n1821__), .dout(new_new_n4775__));
  buf1  g3314(.din(new_new_n4775__), .dout(new_new_n4776__));
  buf1  g3315(.din(new_new_n1838__), .dout(new_new_n4777__));
  buf1  g3316(.din(new_new_n4777__), .dout(new_new_n4778__));
  buf1  g3317(.din(new_new_n1825__), .dout(new_new_n4779__));
  buf1  g3318(.din(new_new_n4779__), .dout(new_new_n4780__));
  buf1  g3319(.din(new_new_n1756__), .dout(new_new_n4781__));
  buf1  g3320(.din(new_new_n2609__), .dout(new_new_n4782__));
  buf1  g3321(.din(new_new_n2608__), .dout(new_new_n4783__));
  buf1  g3322(.din(new_new_n2821__), .dout(new_new_n4784__));
  buf1  g3323(.din(new_new_n1697__), .dout(new_new_n4785__));
  buf1  g3324(.din(new_new_n1695__), .dout(new_new_n4786__));
  buf1  g3325(.din(new_new_n1698__), .dout(new_new_n4787__));
  buf1  g3326(.din(new_new_n1696__), .dout(new_new_n4788__));
  buf1  g3327(.din(new_new_n1699__), .dout(new_new_n4789__));
  buf1  g3328(.din(new_new_n1700__), .dout(new_new_n4790__));
  buf1  g3329(.din(new_new_n1731__), .dout(new_new_n4791__));
  buf1  g3330(.din(new_new_n1732__), .dout(new_new_n4792__));
  buf1  g3331(.din(new_new_n2173__), .dout(new_new_n4793__));
  buf1  g3332(.din(new_new_n2174__), .dout(new_new_n4794__));
  buf1  g3333(.din(new_new_n2852__), .dout(new_new_n4795__));
  buf1  g3334(.din(new_new_n3065__), .dout(new_new_n4796__));
  buf1  g3335(.din(new_new_n2866__), .dout(new_new_n4797__));
  buf1  g3336(.din(new_new_n3011__), .dout(new_new_n4798__));
  buf1  g3337(.din(new_new_n3059__), .dout(new_new_n4799__));
  buf1  g3338(.din(new_new_n2898__), .dout(new_new_n4800__));
  buf1  g3339(.din(new_new_n2969__), .dout(new_new_n4801__));
  buf1  g3340(.din(new_new_n3066__), .dout(new_new_n4802__));
  buf1  g3341(.din(new_new_n2920__), .dout(new_new_n4803__));
  buf1  g3342(.din(new_new_n3053__), .dout(new_new_n4804__));
  buf1  g3343(.din(new_new_n3100__), .dout(new_new_n4805__));
  buf1  g3344(.din(new_new_n3103__), .dout(new_new_n4806__));
  buf1  g3345(.din(new_new_n3106__), .dout(new_new_n4807__));
  buf1  g3346(.din(new_new_n2218__), .dout(new_new_n4808__));
  buf1  g3347(.din(new_new_n2180__), .dout(new_new_n4809__));
  buf1  g3348(.din(new_new_n2217__), .dout(new_new_n4810__));
  buf1  g3349(.din(new_new_n4810__), .dout(new_new_n4811__));
  buf1  g3350(.din(new_new_n2179__), .dout(new_new_n4812__));
  buf1  g3351(.din(new_new_n4812__), .dout(new_new_n4813__));
  buf1  g3352(.din(new_new_n3122__), .dout(new_new_n4814__));
  buf1  g3353(.din(new_new_n3120__), .dout(new_new_n4815__));
  buf1  g3354(.din(new_new_n3121__), .dout(new_new_n4816__));
  buf1  g3355(.din(new_new_n4816__), .dout(new_new_n4817__));
  buf1  g3356(.din(new_new_n3119__), .dout(new_new_n4818__));
  buf1  g3357(.din(new_new_n4818__), .dout(new_new_n4819__));
  buf1  g3358(.din(new_new_n4818__), .dout(new_new_n4820__));
  buf1  g3359(.din(new_new_n3114__), .dout(new_new_n4821__));
  buf1  g3360(.din(new_new_n3123__), .dout(new_new_n4822__));
  buf1  g3361(.din(new_new_n3113__), .dout(new_new_n4823__));
  buf1  g3362(.din(new_new_n1605__), .dout(new_new_n4824__));
  buf1  g3363(.din(new_new_n4824__), .dout(new_new_n4825__));
  buf1  g3364(.din(new_new_n1600__), .dout(new_new_n4826__));
  buf1  g3365(.din(new_new_n1606__), .dout(new_new_n4827__));
  buf1  g3366(.din(new_new_n1599__), .dout(new_new_n4828__));
  buf1  g3367(.din(new_new_n4828__), .dout(new_new_n4829__));
  buf1  g3368(.din(new_new_n1624__), .dout(new_new_n4830__));
  buf1  g3369(.din(new_new_n1601__), .dout(new_new_n4831__));
  buf1  g3370(.din(new_new_n4831__), .dout(new_new_n4832__));
  buf1  g3371(.din(new_new_n1623__), .dout(new_new_n4833__));
  buf1  g3372(.din(new_new_n4833__), .dout(new_new_n4834__));
  buf1  g3373(.din(new_new_n1602__), .dout(new_new_n4835__));
  buf1  g3374(.din(new_new_n2894__), .dout(new_new_n4836__));
  buf1  g3375(.din(new_new_n4836__), .dout(new_new_n4837__));
  buf1  g3376(.din(new_new_n2839__), .dout(new_new_n4838__));
  buf1  g3377(.din(new_new_n4838__), .dout(new_new_n4839__));
  buf1  g3378(.din(new_new_n4839__), .dout(new_new_n4840__));
  buf1  g3379(.din(new_new_n4839__), .dout(new_new_n4841__));
  buf1  g3380(.din(new_new_n4838__), .dout(new_new_n4842__));
  buf1  g3381(.din(new_new_n3112__), .dout(new_new_n4843__));
  buf1  g3382(.din(new_new_n2220__), .dout(new_new_n4844__));
  buf1  g3383(.din(new_new_n2182__), .dout(new_new_n4845__));
  buf1  g3384(.din(new_new_n2219__), .dout(new_new_n4846__));
  buf1  g3385(.din(new_new_n4846__), .dout(new_new_n4847__));
  buf1  g3386(.din(new_new_n2181__), .dout(new_new_n4848__));
  buf1  g3387(.din(new_new_n4848__), .dout(new_new_n4849__));
  buf1  g3388(.din(new_new_n3149__), .dout(new_new_n4850__));
  buf1  g3389(.din(new_new_n3147__), .dout(new_new_n4851__));
  buf1  g3390(.din(new_new_n4851__), .dout(new_new_n4852__));
  buf1  g3391(.din(new_new_n3150__), .dout(new_new_n4853__));
  buf1  g3392(.din(new_new_n3148__), .dout(new_new_n4854__));
  buf1  g3393(.din(new_new_n4854__), .dout(new_new_n4855__));
  buf1  g3394(.din(new_new_n4854__), .dout(new_new_n4856__));
  buf1  g3395(.din(new_new_n2222__), .dout(new_new_n4857__));
  buf1  g3396(.din(new_new_n2192__), .dout(new_new_n4858__));
  buf1  g3397(.din(new_new_n2221__), .dout(new_new_n4859__));
  buf1  g3398(.din(new_new_n2191__), .dout(new_new_n4860__));
  buf1  g3399(.din(new_new_n3157__), .dout(new_new_n4861__));
  buf1  g3400(.din(new_new_n4861__), .dout(new_new_n4862__));
  buf1  g3401(.din(new_new_n4861__), .dout(new_new_n4863__));
  buf1  g3402(.din(new_new_n3158__), .dout(new_new_n4864__));
  buf1  g3403(.din(new_new_n4864__), .dout(new_new_n4865__));
  buf1  g3404(.din(new_new_n4865__), .dout(new_new_n4866__));
  buf1  g3405(.din(new_new_n4865__), .dout(new_new_n4867__));
  buf1  g3406(.din(new_new_n4864__), .dout(new_new_n4868__));
  buf1  g3407(.din(new_new_n3161__), .dout(new_new_n4869__));
  buf1  g3408(.din(new_new_n3160__), .dout(new_new_n4870__));
  buf1  g3409(.din(new_new_n4870__), .dout(new_new_n4871__));
  buf1  g3410(.din(new_new_n3162__), .dout(new_new_n4872__));
  buf1  g3411(.din(new_new_n3159__), .dout(new_new_n4873__));
  buf1  g3412(.din(new_new_n4873__), .dout(new_new_n4874__));
  buf1  g3413(.din(new_new_n2858__), .dout(new_new_n4875__));
  buf1  g3414(.din(new_new_n4875__), .dout(new_new_n4876__));
  buf1  g3415(.din(new_new_n4875__), .dout(new_new_n4877__));
  buf1  g3416(.din(new_new_n2859__), .dout(new_new_n4878__));
  buf1  g3417(.din(new_new_n4878__), .dout(new_new_n4879__));
  buf1  g3418(.din(new_new_n4879__), .dout(new_new_n4880__));
  buf1  g3419(.din(new_new_n4878__), .dout(new_new_n4881__));
  buf1  g3420(.din(new_new_n2838__), .dout(new_new_n4882__));
  buf1  g3421(.din(new_new_n4882__), .dout(new_new_n4883__));
  buf1  g3422(.din(new_new_n4883__), .dout(new_new_n4884__));
  buf1  g3423(.din(new_new_n4882__), .dout(new_new_n4885__));
  buf1  g3424(.din(new_new_n1479__), .dout(new_new_n4886__));
  buf1  g3425(.din(new_new_n1477__), .dout(new_new_n4887__));
  buf1  g3426(.din(new_new_n4887__), .dout(new_new_n4888__));
  buf1  g3427(.din(new_new_n3175__), .dout(new_new_n4889__));
  buf1  g3428(.din(new_new_n3094__), .dout(new_new_n4890__));
  buf1  g3429(.din(new_new_n4890__), .dout(new_new_n4891__));
  buf1  g3430(.din(new_new_n3096__), .dout(new_new_n4892__));
  buf1  g3431(.din(new_new_n4892__), .dout(new_new_n4893__));
  buf1  g3432(.din(new_new_n1931__), .dout(new_new_n4894__));
  buf1  g3433(.din(new_new_n1932__), .dout(new_new_n4895__));
  buf1  g3434(.din(new_new_n3179__), .dout(new_new_n4896__));
  buf1  g3435(.din(new_new_n3178__), .dout(new_new_n4897__));
  buf1  g3436(.din(new_new_n4897__), .dout(new_new_n4898__));
  buf1  g3437(.din(new_new_n2203__), .dout(new_new_n4899__));
  buf1  g3438(.din(new_new_n4899__), .dout(new_new_n4900__));
  buf1  g3439(.din(new_new_n4899__), .dout(new_new_n4901__));
  buf1  g3440(.din(new_new_n2201__), .dout(new_new_n4902__));
  buf1  g3441(.din(new_new_n4902__), .dout(new_new_n4903__));
  buf1  g3442(.din(new_new_n4903__), .dout(new_new_n4904__));
  buf1  g3443(.din(new_new_n4903__), .dout(new_new_n4905__));
  buf1  g3444(.din(new_new_n4902__), .dout(new_new_n4906__));
  buf1  g3445(.din(new_new_n4906__), .dout(new_new_n4907__));
  buf1  g3446(.din(new_new_n4906__), .dout(new_new_n4908__));
  buf1  g3447(.din(new_new_n2202__), .dout(new_new_n4909__));
  buf1  g3448(.din(new_new_n4909__), .dout(new_new_n4910__));
  buf1  g3449(.din(new_new_n4910__), .dout(new_new_n4911__));
  buf1  g3450(.din(new_new_n4910__), .dout(new_new_n4912__));
  buf1  g3451(.din(new_new_n4909__), .dout(new_new_n4913__));
  buf1  g3452(.din(new_new_n3186__), .dout(new_new_n4914__));
  buf1  g3453(.din(new_new_n4914__), .dout(new_new_n4915__));
  buf1  g3454(.din(new_new_n3187__), .dout(new_new_n4916__));
  buf1  g3455(.din(new_new_n4916__), .dout(new_new_n4917__));
  buf1  g3456(.din(new_new_n2208__), .dout(new_new_n4918__));
  buf1  g3457(.din(new_new_n2207__), .dout(new_new_n4919__));
  buf1  g3458(.din(new_new_n4919__), .dout(new_new_n4920__));
  buf1  g3459(.din(new_new_n3189__), .dout(new_new_n4921__));
  buf1  g3460(.din(new_new_n4921__), .dout(new_new_n4922__));
  buf1  g3461(.din(new_new_n4922__), .dout(new_new_n4923__));
  buf1  g3462(.din(new_new_n4923__), .dout(new_new_n4924__));
  buf1  g3463(.din(new_new_n4922__), .dout(new_new_n4925__));
  buf1  g3464(.din(new_new_n4921__), .dout(new_new_n4926__));
  buf1  g3465(.din(new_new_n4926__), .dout(new_new_n4927__));
  buf1  g3466(.din(new_new_n4926__), .dout(new_new_n4928__));
  buf1  g3467(.din(new_new_n2243__), .dout(new_new_n4929__));
  buf1  g3468(.din(new_new_n4929__), .dout(new_new_n4930__));
  buf1  g3469(.din(new_new_n4929__), .dout(new_new_n4931__));
  buf1  g3470(.din(new_new_n3188__), .dout(new_new_n4932__));
  buf1  g3471(.din(new_new_n4932__), .dout(new_new_n4933__));
  buf1  g3472(.din(new_new_n4933__), .dout(new_new_n4934__));
  buf1  g3473(.din(new_new_n4933__), .dout(new_new_n4935__));
  buf1  g3474(.din(new_new_n4932__), .dout(new_new_n4936__));
  buf1  g3475(.din(new_new_n4936__), .dout(new_new_n4937__));
  buf1  g3476(.din(new_new_n2244__), .dout(new_new_n4938__));
  buf1  g3477(.din(new_new_n4938__), .dout(new_new_n4939__));
  buf1  g3478(.din(new_new_n3191__), .dout(new_new_n4940__));
  buf1  g3479(.din(new_new_n3190__), .dout(new_new_n4941__));
  buf1  g3480(.din(new_new_n2247__), .dout(new_new_n4942__));
  buf1  g3481(.din(new_new_n2248__), .dout(new_new_n4943__));
  buf1  g3482(.din(new_new_n3196__), .dout(new_new_n4944__));
  buf1  g3483(.din(new_new_n3197__), .dout(new_new_n4945__));
  buf1  g3484(.din(new_new_n2237__), .dout(new_new_n4946__));
  buf1  g3485(.din(new_new_n4946__), .dout(new_new_n4947__));
  buf1  g3486(.din(new_new_n4947__), .dout(new_new_n4948__));
  buf1  g3487(.din(new_new_n4947__), .dout(new_new_n4949__));
  buf1  g3488(.din(new_new_n4946__), .dout(new_new_n4950__));
  buf1  g3489(.din(new_new_n2230__), .dout(new_new_n4951__));
  buf1  g3490(.din(new_new_n4951__), .dout(new_new_n4952__));
  buf1  g3491(.din(new_new_n4952__), .dout(new_new_n4953__));
  buf1  g3492(.din(new_new_n4952__), .dout(new_new_n4954__));
  buf1  g3493(.din(new_new_n4951__), .dout(new_new_n4955__));
  buf1  g3494(.din(new_new_n4955__), .dout(new_new_n4956__));
  buf1  g3495(.din(new_new_n4955__), .dout(new_new_n4957__));
  buf1  g3496(.din(new_new_n2238__), .dout(new_new_n4958__));
  buf1  g3497(.din(new_new_n4958__), .dout(new_new_n4959__));
  buf1  g3498(.din(new_new_n4959__), .dout(new_new_n4960__));
  buf1  g3499(.din(new_new_n4958__), .dout(new_new_n4961__));
  buf1  g3500(.din(new_new_n2229__), .dout(new_new_n4962__));
  buf1  g3501(.din(new_new_n4962__), .dout(new_new_n4963__));
  buf1  g3502(.din(new_new_n4963__), .dout(new_new_n4964__));
  buf1  g3503(.din(new_new_n4963__), .dout(new_new_n4965__));
  buf1  g3504(.din(new_new_n4962__), .dout(new_new_n4966__));
  buf1  g3505(.din(new_new_n2271__), .dout(new_new_n4967__));
  buf1  g3506(.din(new_new_n4967__), .dout(new_new_n4968__));
  buf1  g3507(.din(new_new_n4967__), .dout(new_new_n4969__));
  buf1  g3508(.din(new_new_n2186__), .dout(new_new_n4970__));
  buf1  g3509(.din(new_new_n4970__), .dout(new_new_n4971__));
  buf1  g3510(.din(new_new_n4971__), .dout(new_new_n4972__));
  buf1  g3511(.din(new_new_n4971__), .dout(new_new_n4973__));
  buf1  g3512(.din(new_new_n4970__), .dout(new_new_n4974__));
  buf1  g3513(.din(new_new_n4974__), .dout(new_new_n4975__));
  buf1  g3514(.din(new_new_n4974__), .dout(new_new_n4976__));
  buf1  g3515(.din(new_new_n2272__), .dout(new_new_n4977__));
  buf1  g3516(.din(new_new_n4977__), .dout(new_new_n4978__));
  buf1  g3517(.din(new_new_n2185__), .dout(new_new_n4979__));
  buf1  g3518(.din(new_new_n4979__), .dout(new_new_n4980__));
  buf1  g3519(.din(new_new_n4980__), .dout(new_new_n4981__));
  buf1  g3520(.din(new_new_n4980__), .dout(new_new_n4982__));
  buf1  g3521(.din(new_new_n4979__), .dout(new_new_n4983__));
  buf1  g3522(.din(new_new_n3204__), .dout(new_new_n4984__));
  buf1  g3523(.din(new_new_n4984__), .dout(new_new_n4985__));
  buf1  g3524(.din(new_new_n4985__), .dout(new_new_n4986__));
  buf1  g3525(.din(new_new_n4985__), .dout(new_new_n4987__));
  buf1  g3526(.din(new_new_n4984__), .dout(new_new_n4988__));
  buf1  g3527(.din(new_new_n4988__), .dout(new_new_n4989__));
  buf1  g3528(.din(new_new_n2241__), .dout(new_new_n4990__));
  buf1  g3529(.din(new_new_n4990__), .dout(new_new_n4991__));
  buf1  g3530(.din(new_new_n4990__), .dout(new_new_n4992__));
  buf1  g3531(.din(new_new_n3205__), .dout(new_new_n4993__));
  buf1  g3532(.din(new_new_n4993__), .dout(new_new_n4994__));
  buf1  g3533(.din(new_new_n4994__), .dout(new_new_n4995__));
  buf1  g3534(.din(new_new_n4993__), .dout(new_new_n4996__));
  buf1  g3535(.din(new_new_n2242__), .dout(new_new_n4997__));
  buf1  g3536(.din(new_new_n4997__), .dout(new_new_n4998__));
  buf1  g3537(.din(new_new_n2274__), .dout(new_new_n4999__));
  buf1  g3538(.din(new_new_n2273__), .dout(new_new_n5000__));
  buf1  g3539(.din(new_new_n2161__), .dout(new_new_n5001__));
  buf1  g3540(.din(new_new_n2245__), .dout(new_new_n5002__));
  buf1  g3541(.din(new_new_n5002__), .dout(new_new_n5003__));
  buf1  g3542(.din(new_new_n5002__), .dout(new_new_n5004__));
  buf1  g3543(.din(new_new_n2246__), .dout(new_new_n5005__));
  buf1  g3544(.din(new_new_n3221__), .dout(new_new_n5006__));
  buf1  g3545(.din(new_new_n5006__), .dout(new_new_n5007__));
  buf1  g3546(.din(new_new_n5006__), .dout(new_new_n5008__));
  buf1  g3547(.din(new_new_n3220__), .dout(new_new_n5009__));
  buf1  g3548(.din(new_new_n5009__), .dout(new_new_n5010__));
  buf1  g3549(.din(new_new_n2249__), .dout(new_new_n5011__));
  buf1  g3550(.din(new_new_n5011__), .dout(new_new_n5012__));
  buf1  g3551(.din(new_new_n2250__), .dout(new_new_n5013__));
  buf1  g3552(.din(new_new_n3227__), .dout(new_new_n5014__));
  buf1  g3553(.din(new_new_n3226__), .dout(new_new_n5015__));
  buf1  g3554(.din(new_new_n5015__), .dout(new_new_n5016__));
  buf1  g3555(.din(new_new_n1295__), .dout(new_new_n5017__));
  buf1  g3556(.din(new_new_n5017__), .dout(new_new_n5018__));
  buf1  g3557(.din(new_new_n2251__), .dout(new_new_n5019__));
  buf1  g3558(.din(new_new_n2277__), .dout(new_new_n5020__));
  buf1  g3559(.din(new_new_n5020__), .dout(new_new_n5021__));
  buf1  g3560(.din(new_new_n5021__), .dout(new_new_n5022__));
  buf1  g3561(.din(new_new_n5022__), .dout(new_new_n5023__));
  buf1  g3562(.din(new_new_n5021__), .dout(new_new_n5024__));
  buf1  g3563(.din(new_new_n5020__), .dout(new_new_n5025__));
  buf1  g3564(.din(new_new_n5025__), .dout(new_new_n5026__));
  buf1  g3565(.din(new_new_n5025__), .dout(new_new_n5027__));
  buf1  g3566(.din(new_new_n2255__), .dout(new_new_n5028__));
  buf1  g3567(.din(new_new_n5028__), .dout(new_new_n5029__));
  buf1  g3568(.din(new_new_n5029__), .dout(new_new_n5030__));
  buf1  g3569(.din(new_new_n5029__), .dout(new_new_n5031__));
  buf1  g3570(.din(new_new_n5028__), .dout(new_new_n5032__));
  buf1  g3571(.din(new_new_n5032__), .dout(new_new_n5033__));
  buf1  g3572(.din(new_new_n2278__), .dout(new_new_n5034__));
  buf1  g3573(.din(new_new_n5034__), .dout(new_new_n5035__));
  buf1  g3574(.din(new_new_n5035__), .dout(new_new_n5036__));
  buf1  g3575(.din(new_new_n5035__), .dout(new_new_n5037__));
  buf1  g3576(.din(new_new_n5034__), .dout(new_new_n5038__));
  buf1  g3577(.din(new_new_n5038__), .dout(new_new_n5039__));
  buf1  g3578(.din(new_new_n5038__), .dout(new_new_n5040__));
  buf1  g3579(.din(new_new_n2256__), .dout(new_new_n5041__));
  buf1  g3580(.din(new_new_n5041__), .dout(new_new_n5042__));
  buf1  g3581(.din(new_new_n5042__), .dout(new_new_n5043__));
  buf1  g3582(.din(new_new_n5041__), .dout(new_new_n5044__));
  buf1  g3583(.din(new_new_n2268__), .dout(new_new_n5045__));
  buf1  g3584(.din(new_new_n5045__), .dout(new_new_n5046__));
  buf1  g3585(.din(new_new_n5046__), .dout(new_new_n5047__));
  buf1  g3586(.din(new_new_n5046__), .dout(new_new_n5048__));
  buf1  g3587(.din(new_new_n5045__), .dout(new_new_n5049__));
  buf1  g3588(.din(new_new_n2259__), .dout(new_new_n5050__));
  buf1  g3589(.din(new_new_n5050__), .dout(new_new_n5051__));
  buf1  g3590(.din(new_new_n5051__), .dout(new_new_n5052__));
  buf1  g3591(.din(new_new_n5052__), .dout(new_new_n5053__));
  buf1  g3592(.din(new_new_n5051__), .dout(new_new_n5054__));
  buf1  g3593(.din(new_new_n5050__), .dout(new_new_n5055__));
  buf1  g3594(.din(new_new_n5055__), .dout(new_new_n5056__));
  buf1  g3595(.din(new_new_n5055__), .dout(new_new_n5057__));
  buf1  g3596(.din(new_new_n2267__), .dout(new_new_n5058__));
  buf1  g3597(.din(new_new_n5058__), .dout(new_new_n5059__));
  buf1  g3598(.din(new_new_n5059__), .dout(new_new_n5060__));
  buf1  g3599(.din(new_new_n5059__), .dout(new_new_n5061__));
  buf1  g3600(.din(new_new_n5058__), .dout(new_new_n5062__));
  buf1  g3601(.din(new_new_n5062__), .dout(new_new_n5063__));
  buf1  g3602(.din(new_new_n5062__), .dout(new_new_n5064__));
  buf1  g3603(.din(new_new_n2260__), .dout(new_new_n5065__));
  buf1  g3604(.din(new_new_n5065__), .dout(new_new_n5066__));
  buf1  g3605(.din(new_new_n5066__), .dout(new_new_n5067__));
  buf1  g3606(.din(new_new_n5066__), .dout(new_new_n5068__));
  buf1  g3607(.din(new_new_n5065__), .dout(new_new_n5069__));
  buf1  g3608(.din(new_new_n5069__), .dout(new_new_n5070__));
  buf1  g3609(.din(new_new_n5069__), .dout(new_new_n5071__));
  buf1  g3610(.din(new_new_n3268__), .dout(new_new_n5072__));
  buf1  g3611(.din(new_new_n5072__), .dout(new_new_n5073__));
  buf1  g3612(.din(new_new_n5073__), .dout(new_new_n5074__));
  buf1  g3613(.din(new_new_n5073__), .dout(new_new_n5075__));
  buf1  g3614(.din(new_new_n5072__), .dout(new_new_n5076__));
  buf1  g3615(.din(new_new_n5076__), .dout(new_new_n5077__));
  buf1  g3616(.din(new_new_n5076__), .dout(new_new_n5078__));
  buf1  g3617(.din(new_new_n2164__), .dout(new_new_n5079__));
  buf1  g3618(.din(new_new_n5079__), .dout(new_new_n5080__));
  buf1  g3619(.din(new_new_n5079__), .dout(new_new_n5081__));
  buf1  g3620(.din(new_new_n3269__), .dout(new_new_n5082__));
  buf1  g3621(.din(new_new_n5082__), .dout(new_new_n5083__));
  buf1  g3622(.din(new_new_n5083__), .dout(new_new_n5084__));
  buf1  g3623(.din(new_new_n5083__), .dout(new_new_n5085__));
  buf1  g3624(.din(new_new_n5082__), .dout(new_new_n5086__));
  buf1  g3625(.din(new_new_n5086__), .dout(new_new_n5087__));
  buf1  g3626(.din(new_new_n2163__), .dout(new_new_n5088__));
  buf1  g3627(.din(new_new_n5088__), .dout(new_new_n5089__));
  buf1  g3628(.din(new_new_n5089__), .dout(new_new_n5090__));
  buf1  g3629(.din(new_new_n5089__), .dout(new_new_n5091__));
  buf1  g3630(.din(new_new_n5088__), .dout(new_new_n5092__));
  buf1  g3631(.din(new_new_n2205__), .dout(new_new_n5093__));
  buf1  g3632(.din(new_new_n5093__), .dout(new_new_n5094__));
  buf1  g3633(.din(new_new_n5094__), .dout(new_new_n5095__));
  buf1  g3634(.din(new_new_n5093__), .dout(new_new_n5096__));
  buf1  g3635(.din(new_new_n2206__), .dout(new_new_n5097__));
  buf1  g3636(.din(new_new_n1855__), .dout(new_new_n5098__));
  buf1  g3637(.din(new_new_n5098__), .dout(new_new_n5099__));
  buf1  g3638(.din(new_new_n1856__), .dout(new_new_n5100__));
  buf1  g3639(.din(new_new_n3281__), .dout(new_new_n5101__));
  buf1  g3640(.din(new_new_n5101__), .dout(new_new_n5102__));
  buf1  g3641(.din(new_new_n5102__), .dout(new_new_n5103__));
  buf1  g3642(.din(new_new_n5103__), .dout(new_new_n5104__));
  buf1  g3643(.din(new_new_n5102__), .dout(new_new_n5105__));
  buf1  g3644(.din(new_new_n5101__), .dout(new_new_n5106__));
  buf1  g3645(.din(new_new_n5106__), .dout(new_new_n5107__));
  buf1  g3646(.din(new_new_n5106__), .dout(new_new_n5108__));
  buf1  g3647(.din(new_new_n3280__), .dout(new_new_n5109__));
  buf1  g3648(.din(new_new_n5109__), .dout(new_new_n5110__));
  buf1  g3649(.din(new_new_n5110__), .dout(new_new_n5111__));
  buf1  g3650(.din(new_new_n5110__), .dout(new_new_n5112__));
  buf1  g3651(.din(new_new_n5109__), .dout(new_new_n5113__));
  buf1  g3652(.din(new_new_n5113__), .dout(new_new_n5114__));
  buf1  g3653(.din(new_new_n5113__), .dout(new_new_n5115__));
  buf1  g3654(.din(new_new_n3284__), .dout(new_new_n5116__));
  buf1  g3655(.din(new_new_n5116__), .dout(new_new_n5117__));
  buf1  g3656(.din(new_new_n5117__), .dout(new_new_n5118__));
  buf1  g3657(.din(new_new_n5118__), .dout(new_new_n5119__));
  buf1  g3658(.din(new_new_n5117__), .dout(new_new_n5120__));
  buf1  g3659(.din(new_new_n5116__), .dout(new_new_n5121__));
  buf1  g3660(.din(new_new_n5121__), .dout(new_new_n5122__));
  buf1  g3661(.din(new_new_n5121__), .dout(new_new_n5123__));
  buf1  g3662(.din(new_new_n3285__), .dout(new_new_n5124__));
  buf1  g3663(.din(new_new_n5124__), .dout(new_new_n5125__));
  buf1  g3664(.din(new_new_n5125__), .dout(new_new_n5126__));
  buf1  g3665(.din(new_new_n5125__), .dout(new_new_n5127__));
  buf1  g3666(.din(new_new_n5124__), .dout(new_new_n5128__));
  buf1  g3667(.din(new_new_n5128__), .dout(new_new_n5129__));
  buf1  g3668(.din(new_new_n5128__), .dout(new_new_n5130__));
  buf1  g3669(.din(new_new_n3289__), .dout(new_new_n5131__));
  buf1  g3670(.din(new_new_n5131__), .dout(new_new_n5132__));
  buf1  g3671(.din(new_new_n5131__), .dout(new_new_n5133__));
  buf1  g3672(.din(new_new_n3288__), .dout(new_new_n5134__));
  buf1  g3673(.din(new_new_n5134__), .dout(new_new_n5135__));
  buf1  g3674(.din(new_new_n3290__), .dout(new_new_n5136__));
  buf1  g3675(.din(new_new_n5136__), .dout(new_new_n5137__));
  buf1  g3676(.din(new_new_n5137__), .dout(new_new_n5138__));
  buf1  g3677(.din(new_new_n5137__), .dout(new_new_n5139__));
  buf1  g3678(.din(new_new_n5136__), .dout(new_new_n5140__));
  buf1  g3679(.din(new_new_n5140__), .dout(new_new_n5141__));
  buf1  g3680(.din(new_new_n5140__), .dout(new_new_n5142__));
  buf1  g3681(.din(new_new_n3291__), .dout(new_new_n5143__));
  buf1  g3682(.din(new_new_n5143__), .dout(new_new_n5144__));
  buf1  g3683(.din(new_new_n5144__), .dout(new_new_n5145__));
  buf1  g3684(.din(new_new_n5144__), .dout(new_new_n5146__));
  buf1  g3685(.din(new_new_n5143__), .dout(new_new_n5147__));
  buf1  g3686(.din(new_new_n5147__), .dout(new_new_n5148__));
  buf1  g3687(.din(new_new_n3301__), .dout(new_new_n5149__));
  buf1  g3688(.din(new_new_n5149__), .dout(new_new_n5150__));
  buf1  g3689(.din(new_new_n5150__), .dout(new_new_n5151__));
  buf1  g3690(.din(new_new_n5151__), .dout(new_new_n5152__));
  buf1  g3691(.din(new_new_n5150__), .dout(new_new_n5153__));
  buf1  g3692(.din(new_new_n5149__), .dout(new_new_n5154__));
  buf1  g3693(.din(new_new_n5154__), .dout(new_new_n5155__));
  buf1  g3694(.din(new_new_n5154__), .dout(new_new_n5156__));
  buf1  g3695(.din(new_new_n3300__), .dout(new_new_n5157__));
  buf1  g3696(.din(new_new_n5157__), .dout(new_new_n5158__));
  buf1  g3697(.din(new_new_n5158__), .dout(new_new_n5159__));
  buf1  g3698(.din(new_new_n5158__), .dout(new_new_n5160__));
  buf1  g3699(.din(new_new_n5157__), .dout(new_new_n5161__));
  buf1  g3700(.din(new_new_n5161__), .dout(new_new_n5162__));
  buf1  g3701(.din(new_new_n3303__), .dout(new_new_n5163__));
  buf1  g3702(.din(new_new_n5163__), .dout(new_new_n5164__));
  buf1  g3703(.din(new_new_n5164__), .dout(new_new_n5165__));
  buf1  g3704(.din(new_new_n5163__), .dout(new_new_n5166__));
  buf1  g3705(.din(new_new_n3302__), .dout(new_new_n5167__));
  buf1  g3706(.din(new_new_n5167__), .dout(new_new_n5168__));
  buf1  g3707(.din(new_new_n5167__), .dout(new_new_n5169__));
  buf1  g3708(.din(new_new_n1859__), .dout(new_new_n5170__));
  buf1  g3709(.din(new_new_n5170__), .dout(new_new_n5171__));
  buf1  g3710(.din(new_new_n5171__), .dout(new_new_n5172__));
  buf1  g3711(.din(new_new_n5171__), .dout(new_new_n5173__));
  buf1  g3712(.din(new_new_n5170__), .dout(new_new_n5174__));
  buf1  g3713(.din(new_new_n5174__), .dout(new_new_n5175__));
  buf1  g3714(.din(new_new_n5174__), .dout(new_new_n5176__));
  buf1  g3715(.din(new_new_n1860__), .dout(new_new_n5177__));
  buf1  g3716(.din(new_new_n5177__), .dout(new_new_n5178__));
  buf1  g3717(.din(new_new_n5178__), .dout(new_new_n5179__));
  buf1  g3718(.din(new_new_n5178__), .dout(new_new_n5180__));
  buf1  g3719(.din(new_new_n5177__), .dout(new_new_n5181__));
  buf1  g3720(.din(new_new_n2269__), .dout(new_new_n5182__));
  buf1  g3721(.din(new_new_n5182__), .dout(new_new_n5183__));
  buf1  g3722(.din(new_new_n5182__), .dout(new_new_n5184__));
  buf1  g3723(.din(new_new_n2270__), .dout(new_new_n5185__));
  buf1  g3724(.din(new_new_n5185__), .dout(new_new_n5186__));
  buf1  g3725(.din(new_new_n3311__), .dout(new_new_n5187__));
  buf1  g3726(.din(new_new_n5187__), .dout(new_new_n5188__));
  buf1  g3727(.din(new_new_n3310__), .dout(new_new_n5189__));
  buf1  g3728(.din(new_new_n5189__), .dout(new_new_n5190__));
  buf1  g3729(.din(new_new_n5189__), .dout(new_new_n5191__));
  buf1  g3730(.din(new_new_n3298__), .dout(new_new_n5192__));
  buf1  g3731(.din(new_new_n5192__), .dout(new_new_n5193__));
  buf1  g3732(.din(new_new_n5193__), .dout(new_new_n5194__));
  buf1  g3733(.din(new_new_n5192__), .dout(new_new_n5195__));
  buf1  g3734(.din(new_new_n1270__), .dout(new_new_n5196__));
  buf1  g3735(.din(new_new_n5196__), .dout(new_new_n5197__));
  buf1  g3736(.din(new_new_n5197__), .dout(new_new_n5198__));
  buf1  g3737(.din(new_new_n5197__), .dout(new_new_n5199__));
  buf1  g3738(.din(new_new_n5196__), .dout(new_new_n5200__));
  buf1  g3739(.din(new_new_n3327__), .dout(new_new_n5201__));
  buf1  g3740(.din(new_new_n1272__), .dout(new_new_n5202__));
  buf1  g3741(.din(new_new_n5202__), .dout(new_new_n5203__));
  buf1  g3742(.din(new_new_n5203__), .dout(new_new_n5204__));
  buf1  g3743(.din(new_new_n5203__), .dout(new_new_n5205__));
  buf1  g3744(.din(new_new_n5202__), .dout(new_new_n5206__));
  buf1  g3745(.din(new_new_n3091__), .dout(new_new_n5207__));
  buf1  g3746(.din(new_new_n5207__), .dout(new_new_n5208__));
  buf1  g3747(.din(new_new_n1858__), .dout(new_new_n5209__));
  buf1  g3748(.din(new_new_n5209__), .dout(new_new_n5210__));
  buf1  g3749(.din(new_new_n5210__), .dout(new_new_n5211__));
  buf1  g3750(.din(new_new_n5209__), .dout(new_new_n5212__));
  buf1  g3751(.din(new_new_n1857__), .dout(new_new_n5213__));
  buf1  g3752(.din(new_new_n5213__), .dout(new_new_n5214__));
  buf1  g3753(.din(new_new_n5214__), .dout(new_new_n5215__));
  buf1  g3754(.din(new_new_n5214__), .dout(new_new_n5216__));
  buf1  g3755(.din(new_new_n5213__), .dout(new_new_n5217__));
  buf1  g3756(.din(new_new_n5217__), .dout(new_new_n5218__));
  buf1  g3757(.din(new_new_n5217__), .dout(new_new_n5219__));
  buf1  g3758(.din(new_new_n2235__), .dout(new_new_n5220__));
  buf1  g3759(.din(new_new_n5220__), .dout(new_new_n5221__));
  buf1  g3760(.din(new_new_n5221__), .dout(new_new_n5222__));
  buf1  g3761(.din(new_new_n5220__), .dout(new_new_n5223__));
  buf1  g3762(.din(new_new_n2236__), .dout(new_new_n5224__));
  buf1  g3763(.din(new_new_n2165__), .dout(new_new_n5225__));
  buf1  g3764(.din(new_new_n5225__), .dout(new_new_n5226__));
  buf1  g3765(.din(new_new_n5226__), .dout(new_new_n5227__));
  buf1  g3766(.din(new_new_n5226__), .dout(new_new_n5228__));
  buf1  g3767(.din(new_new_n5225__), .dout(new_new_n5229__));
  buf1  g3768(.din(new_new_n5229__), .dout(new_new_n5230__));
  buf1  g3769(.din(new_new_n5229__), .dout(new_new_n5231__));
  buf1  g3770(.din(new_new_n2166__), .dout(new_new_n5232__));
  buf1  g3771(.din(new_new_n5232__), .dout(new_new_n5233__));
  buf1  g3772(.din(new_new_n5233__), .dout(new_new_n5234__));
  buf1  g3773(.din(new_new_n5233__), .dout(new_new_n5235__));
  buf1  g3774(.din(new_new_n5232__), .dout(new_new_n5236__));
  buf1  g3775(.din(new_new_n2257__), .dout(new_new_n5237__));
  buf1  g3776(.din(new_new_n5237__), .dout(new_new_n5238__));
  buf1  g3777(.din(new_new_n5237__), .dout(new_new_n5239__));
  buf1  g3778(.din(new_new_n2258__), .dout(new_new_n5240__));
  buf1  g3779(.din(new_new_n3358__), .dout(new_new_n5241__));
  buf1  g3780(.din(new_new_n5241__), .dout(new_new_n5242__));
  buf1  g3781(.din(new_new_n5242__), .dout(new_new_n5243__));
  buf1  g3782(.din(new_new_n5241__), .dout(new_new_n5244__));
  buf1  g3783(.din(new_new_n3379__), .dout(new_new_n5245__));
  buf1  g3784(.din(new_new_n3405__), .dout(new_new_n5246__));
  buf1  g3785(.din(new_new_n5246__), .dout(new_new_n5247__));
  buf1  g3786(.din(new_new_n5246__), .dout(new_new_n5248__));
  buf1  g3787(.din(new_new_n3404__), .dout(new_new_n5249__));
  buf1  g3788(.din(new_new_n5249__), .dout(new_new_n5250__));
  buf1  g3789(.din(new_new_n5249__), .dout(new_new_n5251__));
  buf1  g3790(.din(new_new_n1299__), .dout(new_new_n5252__));
  buf1  g3791(.din(new_new_n1303__), .dout(new_new_n5253__));
  buf1  g3792(.din(new_new_n1267__), .dout(new_new_n5254__));
  buf1  g3793(.din(new_new_n2239__), .dout(new_new_n5255__));
  buf1  g3794(.din(new_new_n3476__), .dout(new_new_n5256__));
  buf1  g3795(.din(new_new_n5256__), .dout(new_new_n5257__));
  buf1  g3796(.din(new_new_n5257__), .dout(new_new_n5258__));
  buf1  g3797(.din(new_new_n5256__), .dout(new_new_n5259__));
  buf1  g3798(.din(new_new_n3497__), .dout(new_new_n5260__));
  buf1  g3799(.din(new_new_n3337__), .dout(new_new_n5261__));
  buf1  g3800(.din(new_new_n3502__), .dout(new_new_n5262__));
  buf1  g3801(.din(new_new_n5262__), .dout(new_new_n5263__));
  buf1  g3802(.din(new_new_n3331__), .dout(new_new_n5264__));
  buf1  g3803(.din(new_new_n3329__), .dout(new_new_n5265__));
  buf1  g3804(.din(new_new_n1273__), .dout(new_new_n5266__));
  buf1  g3805(.din(new_new_n5266__), .dout(new_new_n5267__));
  buf1  g3806(.din(new_new_n5266__), .dout(new_new_n5268__));
  buf1  g3807(.din(new_new_n3326__), .dout(new_new_n5269__));
  buf1  g3808(.din(new_new_n1275__), .dout(new_new_n5270__));
  buf1  g3809(.din(new_new_n5270__), .dout(new_new_n5271__));
  buf1  g3810(.din(new_new_n5270__), .dout(new_new_n5272__));
  buf1  g3811(.din(new_new_n3092__), .dout(new_new_n5273__));
  buf1  g3812(.din(new_new_n1328__), .dout(new_new_n5274__));
  buf1  g3813(.din(new_new_n5274__), .dout(new_new_n5275__));
  buf1  g3814(.din(new_new_n5275__), .dout(new_new_n5276__));
  buf1  g3815(.din(new_new_n5275__), .dout(new_new_n5277__));
  buf1  g3816(.din(new_new_n5274__), .dout(new_new_n5278__));
  buf1  g3817(.din(new_new_n5278__), .dout(new_new_n5279__));
  buf1  g3818(.din(new_new_n3333__), .dout(new_new_n5280__));
  buf1  g3819(.din(new_new_n1621__), .dout(new_new_n5281__));
  buf1  g3820(.din(new_new_n5281__), .dout(new_new_n5282__));
  buf1  g3821(.din(new_new_n5281__), .dout(new_new_n5283__));
  buf1  g3822(.din(new_new_n2908__), .dout(new_new_n5284__));
  buf1  g3823(.din(new_new_n5284__), .dout(new_new_n5285__));
  buf1  g3824(.din(new_new_n2902__), .dout(new_new_n5286__));
  buf1  g3825(.din(new_new_n5286__), .dout(new_new_n5287__));
  buf1  g3826(.din(new_new_n3068__), .dout(new_new_n5288__));
  buf1  g3827(.din(new_new_n5288__), .dout(new_new_n5289__));
  buf1  g3828(.din(new_new_n2904__), .dout(new_new_n5290__));
  buf1  g3829(.din(new_new_n5290__), .dout(new_new_n5291__));
  buf1  g3830(.din(new_new_n3545__), .dout(new_new_n5292__));
  buf1  g3831(.din(new_new_n3544__), .dout(new_new_n5293__));
  buf1  g3832(.din(new_new_n5293__), .dout(new_new_n5294__));
  buf1  g3833(.din(new_new_n3550__), .dout(new_new_n5295__));
  buf1  g3834(.din(new_new_n5295__), .dout(new_new_n5296__));
  buf1  g3835(.din(new_new_n5295__), .dout(new_new_n5297__));
  buf1  g3836(.din(new_new_n3334__), .dout(new_new_n5298__));
  buf1  g3837(.din(new_new_n5298__), .dout(new_new_n5299__));
  buf1  g3838(.din(new_new_n3524__), .dout(new_new_n5300__));
  buf1  g3839(.din(new_new_n3449__), .dout(new_new_n5301__));
  buf1  g3840(.din(new_new_n5301__), .dout(new_new_n5302__));
  buf1  g3841(.din(new_new_n5302__), .dout(new_new_n5303__));
  buf1  g3842(.din(new_new_n5301__), .dout(new_new_n5304__));
  buf1  g3843(.din(new_new_n3503__), .dout(new_new_n5305__));
  buf1  g3844(.din(new_new_n5305__), .dout(new_new_n5306__));
  buf1  g3845(.din(new_new_n5306__), .dout(new_new_n5307__));
  buf1  g3846(.din(new_new_n5305__), .dout(new_new_n5308__));
  buf1  g3847(.din(new_new_n3184__), .dout(new_new_n5309__));
  buf1  g3848(.din(new_new_n1625__), .dout(new_new_n5310__));
  buf1  g3849(.din(new_new_n1627__), .dout(new_new_n5311__));
  buf1  g3850(.din(new_new_n1657__), .dout(new_new_n5312__));
  buf1  g3851(.din(new_new_n1675__), .dout(new_new_n5313__));
  buf1  g3852(.din(new_new_n3551__), .dout(new_new_n5314__));
  buf1  g3853(.din(new_new_n5314__), .dout(new_new_n5315__));
  buf1  g3854(.din(new_new_n3125__), .dout(new_new_n5316__));
  buf1  g3855(.din(new_new_n1529__), .dout(new_new_n5317__));
  buf1  g3856(.din(new_new_n5317__), .dout(new_new_n5318__));
  buf1  g3857(.din(new_new_n1535__), .dout(new_new_n5319__));
  buf1  g3858(.din(new_new_n5319__), .dout(new_new_n5320__));
  buf1  g3859(.din(new_new_n5319__), .dout(new_new_n5321__));
  buf1  g3860(.din(new_new_n1597__), .dout(new_new_n5322__));
  buf1  g3861(.din(new_new_n5322__), .dout(new_new_n5323__));
  buf1  g3862(.din(new_new_n5322__), .dout(new_new_n5324__));
  buf1  g3863(.din(new_new_n3579__), .dout(new_new_n5325__));
  buf1  g3864(.din(new_new_n3578__), .dout(new_new_n5326__));
  buf1  g3865(.din(new_new_n5326__), .dout(new_new_n5327__));
  buf1  g3866(.din(new_new_n1549__), .dout(new_new_n5328__));
  buf1  g3867(.din(new_new_n5328__), .dout(new_new_n5329__));
  buf1  g3868(.din(new_new_n5329__), .dout(new_new_n5330__));
  buf1  g3869(.din(new_new_n5328__), .dout(new_new_n5331__));
  buf1  g3870(.din(new_new_n1550__), .dout(new_new_n5332__));
  buf1  g3871(.din(new_new_n5332__), .dout(new_new_n5333__));
  buf1  g3872(.din(new_new_n3603__), .dout(new_new_n5334__));
  buf1  g3873(.din(new_new_n5334__), .dout(new_new_n5335__));
  buf1  g3874(.din(new_new_n3605__), .dout(new_new_n5336__));
  buf1  g3875(.din(new_new_n3602__), .dout(new_new_n5337__));
  buf1  g3876(.din(new_new_n5337__), .dout(new_new_n5338__));
  buf1  g3877(.din(new_new_n5337__), .dout(new_new_n5339__));
  buf1  g3878(.din(new_new_n3601__), .dout(new_new_n5340__));
  buf1  g3879(.din(new_new_n5340__), .dout(new_new_n5341__));
  buf1  g3880(.din(new_new_n5340__), .dout(new_new_n5342__));
  buf1  g3881(.din(new_new_n3608__), .dout(new_new_n5343__));
  buf1  g3882(.din(new_new_n3609__), .dout(new_new_n5344__));
  buf1  g3883(.din(new_new_n3611__), .dout(new_new_n5345__));
  buf1  g3884(.din(new_new_n3613__), .dout(new_new_n5346__));
  buf1  g3885(.din(new_new_n3383__), .dout(new_new_n5347__));
  buf1  g3886(.din(new_new_n3381__), .dout(new_new_n5348__));
  buf1  g3887(.din(new_new_n3378__), .dout(new_new_n5349__));
  buf1  g3888(.din(new_new_n1604__), .dout(new_new_n5350__));
  buf1  g3889(.din(new_new_n5350__), .dout(new_new_n5351__));
  buf1  g3890(.din(new_new_n1528__), .dout(new_new_n5352__));
  buf1  g3891(.din(new_new_n5352__), .dout(new_new_n5353__));
  buf1  g3892(.din(new_new_n3539__), .dout(new_new_n5354__));
  buf1  g3893(.din(new_new_n1619__), .dout(new_new_n5355__));
  buf1  g3894(.din(new_new_n5355__), .dout(new_new_n5356__));
  buf1  g3895(.din(new_new_n5356__), .dout(new_new_n5357__));
  buf1  g3896(.din(new_new_n5355__), .dout(new_new_n5358__));
  buf1  g3897(.din(new_new_n1534__), .dout(new_new_n5359__));
  buf1  g3898(.din(new_new_n5359__), .dout(new_new_n5360__));
  buf1  g3899(.din(new_new_n3630__), .dout(new_new_n5361__));
  buf1  g3900(.din(new_new_n3536__), .dout(new_new_n5362__));
  buf1  g3901(.din(new_new_n3562__), .dout(new_new_n5363__));
  buf1  g3902(.din(new_new_n5363__), .dout(new_new_n5364__));
  buf1  g3903(.din(new_new_n5363__), .dout(new_new_n5365__));
  buf1  g3904(.din(new_new_n3560__), .dout(new_new_n5366__));
  buf1  g3905(.din(new_new_n5366__), .dout(new_new_n5367__));
  buf1  g3906(.din(new_new_n5366__), .dout(new_new_n5368__));
  buf1  g3907(.din(new_new_n3641__), .dout(new_new_n5369__));
  buf1  g3908(.din(new_new_n5369__), .dout(new_new_n5370__));
  buf1  g3909(.din(new_new_n3634__), .dout(new_new_n5371__));
  buf1  g3910(.din(new_new_n5371__), .dout(new_new_n5372__));
  buf1  g3911(.din(new_new_n3668__), .dout(new_new_n5373__));
  buf1  g3912(.din(new_new_n5373__), .dout(new_new_n5374__));
  buf1  g3913(.din(new_new_n5373__), .dout(new_new_n5375__));
  buf1  g3914(.din(new_new_n1269__), .dout(new_new_n5376__));
  buf1  g3915(.din(new_new_n5376__), .dout(new_new_n5377__));
  buf1  g3916(.din(new_new_n5376__), .dout(new_new_n5378__));
  buf1  g3917(.din(new_new_n3667__), .dout(new_new_n5379__));
  buf1  g3918(.din(new_new_n5379__), .dout(new_new_n5380__));
  buf1  g3919(.din(new_new_n5379__), .dout(new_new_n5381__));
  buf1  g3920(.din(new_new_n3262__), .dout(new_new_n5382__));
  buf1  g3921(.din(new_new_n3263__), .dout(new_new_n5383__));
  buf1  g3922(.din(new_new_n5383__), .dout(new_new_n5384__));
  buf1  g3923(.din(new_new_n5384__), .dout(new_new_n5385__));
  buf1  g3924(.din(new_new_n5383__), .dout(new_new_n5386__));
  buf1  g3925(.din(new_new_n1271__), .dout(new_new_n5387__));
  buf1  g3926(.din(new_new_n5387__), .dout(new_new_n5388__));
  buf1  g3927(.din(new_new_n5388__), .dout(new_new_n5389__));
  buf1  g3928(.din(new_new_n5387__), .dout(new_new_n5390__));
  buf1  g3929(.din(new_new_n3413__), .dout(new_new_n5391__));
  buf1  g3930(.din(new_new_n5391__), .dout(new_new_n5392__));
  buf1  g3931(.din(new_new_n5392__), .dout(new_new_n5393__));
  buf1  g3932(.din(new_new_n5391__), .dout(new_new_n5394__));
  buf1  g3933(.din(new_new_n3412__), .dout(new_new_n5395__));
  buf1  g3934(.din(new_new_n5395__), .dout(new_new_n5396__));
  buf1  g3935(.din(new_new_n3242__), .dout(new_new_n5397__));
  buf1  g3936(.din(new_new_n3243__), .dout(new_new_n5398__));
  buf1  g3937(.din(new_new_n5398__), .dout(new_new_n5399__));
  buf1  g3938(.din(new_new_n5399__), .dout(new_new_n5400__));
  buf1  g3939(.din(new_new_n5398__), .dout(new_new_n5401__));
  buf1  g3940(.din(new_new_n1547__), .dout(new_new_n5402__));
  buf1  g3941(.din(new_new_n1545__), .dout(new_new_n5403__));
  buf1  g3942(.din(new_new_n5403__), .dout(new_new_n5404__));
  buf1  g3943(.din(new_new_n1533__), .dout(new_new_n5405__));
  buf1  g3944(.din(new_new_n5405__), .dout(new_new_n5406__));
  buf1  g3945(.din(new_new_n5406__), .dout(new_new_n5407__));
  buf1  g3946(.din(new_new_n5406__), .dout(new_new_n5408__));
  buf1  g3947(.din(new_new_n5405__), .dout(new_new_n5409__));
  buf1  g3948(.din(new_new_n1527__), .dout(new_new_n5410__));
  buf1  g3949(.din(new_new_n5410__), .dout(new_new_n5411__));
  buf1  g3950(.din(new_new_n5411__), .dout(new_new_n5412__));
  buf1  g3951(.din(new_new_n5411__), .dout(new_new_n5413__));
  buf1  g3952(.din(new_new_n5410__), .dout(new_new_n5414__));
  buf1  g3953(.din(new_new_n1620__), .dout(new_new_n5415__));
  buf1  g3954(.din(new_new_n5415__), .dout(new_new_n5416__));
  buf1  g3955(.din(new_new_n3538__), .dout(new_new_n5417__));
  buf1  g3956(.din(new_new_n3335__), .dout(new_new_n5418__));
  buf1  g3957(.din(new_new_n1327__), .dout(new_new_n5419__));
  buf1  g3958(.din(new_new_n3140__), .dout(new_new_n5420__));
  buf1  g3959(.din(new_new_n3558__), .dout(new_new_n5421__));
  buf1  g3960(.din(new_new_n3556__), .dout(new_new_n5422__));
  buf1  g3961(.din(new_new_n1603__), .dout(new_new_n5423__));
  buf1  g3962(.din(new_new_n5423__), .dout(new_new_n5424__));
  buf1  g3963(.din(new_new_n5424__), .dout(new_new_n5425__));
  buf1  g3964(.din(new_new_n5423__), .dout(new_new_n5426__));
  buf1  g3965(.din(new_new_n2900__), .dout(new_new_n5427__));
  buf1  g3966(.din(new_new_n2899__), .dout(new_new_n5428__));
  buf1  g3967(.din(new_new_n5428__), .dout(new_new_n5429__));
  buf1  g3968(.din(new_new_n3174__), .dout(new_new_n5430__));
  buf1  g3969(.din(new_new_n3132__), .dout(new_new_n5431__));
  buf1  g3970(.din(new_new_n3138__), .dout(new_new_n5432__));
  buf1  g3971(.din(new_new_n3439__), .dout(new_new_n5433__));
  buf1  g3972(.din(new_new_n5433__), .dout(new_new_n5434__));
  buf1  g3973(.din(new_new_n5434__), .dout(new_new_n5435__));
  buf1  g3974(.din(new_new_n5433__), .dout(new_new_n5436__));
  buf1  g3975(.din(new_new_n3216__), .dout(new_new_n5437__));
  buf1  g3976(.din(new_new_n1274__), .dout(new_new_n5438__));
  buf1  g3977(.din(new_new_n5438__), .dout(new_new_n5439__));
  buf1  g3978(.din(new_new_n5438__), .dout(new_new_n5440__));
  buf1  g3979(.din(new_new_n3217__), .dout(new_new_n5441__));
  buf1  g3980(.din(new_new_n5441__), .dout(new_new_n5442__));
  buf1  g3981(.din(new_new_n1276__), .dout(new_new_n5443__));
  buf1  g3982(.din(new_new_n5443__), .dout(new_new_n5444__));
  buf1  g3983(.din(new_new_n5443__), .dout(new_new_n5445__));
  buf1  g3984(.din(new_new_n3741__), .dout(new_new_n5446__));
  buf1  g3985(.din(new_new_n3678__), .dout(new_new_n5447__));
  buf1  g3986(.din(new_new_n3501__), .dout(new_new_n5448__));
  buf1  g3987(.din(new_new_n3499__), .dout(new_new_n5449__));
  buf1  g3988(.din(new_new_n3496__), .dout(new_new_n5450__));
  buf1  g3989(.din(new_new_n3688__), .dout(new_new_n5451__));
  buf1  g3990(.din(new_new_n3525__), .dout(new_new_n5452__));
  buf1  g3991(.din(new_new_n5452__), .dout(new_new_n5453__));
  buf1  g3992(.din(new_new_n5452__), .dout(new_new_n5454__));
  buf1  g3993(.din(new_new_n1139__), .dout(new_new_n5455__));
  buf1  g3994(.din(new_new_n5455__), .dout(new_new_n5456__));
  buf1  g3995(.din(new_new_n1137__), .dout(new_new_n5457__));
  buf1  g3996(.din(new_new_n5457__), .dout(new_new_n5458__));
  buf1  g3997(.din(new_new_n5458__), .dout(new_new_n5459__));
  buf1  g3998(.din(new_new_n5458__), .dout(new_new_n5460__));
  buf1  g3999(.din(new_new_n5457__), .dout(new_new_n5461__));
  buf1  g4000(.din(new_new_n5461__), .dout(new_new_n5462__));
  buf1  g4001(.din(new_new_n5461__), .dout(new_new_n5463__));
  buf1  g4002(.din(new_new_n1265__), .dout(new_new_n5464__));
  buf1  g4003(.din(new_new_n3770__), .dout(new_new_n5465__));
  buf1  g4004(.din(new_new_n5465__), .dout(new_new_n5466__));
  buf1  g4005(.din(new_new_n3748__), .dout(new_new_n5467__));
  buf1  g4006(.din(new_new_n5467__), .dout(new_new_n5468__));
  buf1  g4007(.din(new_new_n5467__), .dout(new_new_n5469__));
  buf1  g4008(.din(new_new_n3696__), .dout(new_new_n5470__));
  buf1  g4009(.din(new_new_n3755__), .dout(new_new_n5471__));
  buf1  g4010(.din(new_new_n5471__), .dout(new_new_n5472__));
  buf1  g4011(.din(new_new_n1141__), .dout(new_new_n5473__));
  buf1  g4012(.din(new_new_n3778__), .dout(new_new_n5474__));
  buf1  g4013(.din(new_new_n5474__), .dout(new_new_n5475__));
  buf1  g4014(.din(new_new_n1135__), .dout(new_new_n5476__));
  buf1  g4015(.din(new_new_n5476__), .dout(new_new_n5477__));
  buf1  g4016(.din(new_new_n1133__), .dout(new_new_n5478__));
  buf1  g4017(.din(new_new_n1551__), .dout(new_new_n5479__));
  buf1  g4018(.din(new_new_n5479__), .dout(new_new_n5480__));
  buf1  g4019(.din(new_new_n5480__), .dout(new_new_n5481__));
  buf1  g4020(.din(new_new_n5479__), .dout(new_new_n5482__));
  buf1  g4021(.din(new_new_n2906__), .dout(new_new_n5483__));
  buf1  g4022(.din(new_new_n5483__), .dout(new_new_n5484__));
  buf1  g4023(.din(new_new_n5483__), .dout(new_new_n5485__));
  buf1  g4024(.din(new_new_n3098__), .dout(new_new_n5486__));
  buf1  g4025(.din(new_new_n5486__), .dout(new_new_n5487__));
  buf1  g4026(.din(new_new_n5486__), .dout(new_new_n5488__));
  buf1  g4027(.din(new_new_n3176__), .dout(new_new_n5489__));
  buf1  g4028(.din(new_new_n3177__), .dout(new_new_n5490__));
  buf1  g4029(.din(new_new_n3533__), .dout(new_new_n5491__));
  buf1  g4030(.din(new_new_n5491__), .dout(new_new_n5492__));
  buf1  g4031(.din(new_new_n5491__), .dout(new_new_n5493__));
  buf1  g4032(.din(new_new_n3553__), .dout(new_new_n5494__));
  buf1  g4033(.din(new_new_n3554__), .dout(new_new_n5495__));
  buf1  g4034(.din(new_new_n3559__), .dout(new_new_n5496__));
  buf1  g4035(.din(new_new_n5496__), .dout(new_new_n5497__));
  buf1  g4036(.din(new_new_n3565__), .dout(new_new_n5498__));
  buf1  g4037(.din(new_new_n3568__), .dout(new_new_n5499__));
  buf1  g4038(.din(new_new_n3571__), .dout(new_new_n5500__));
  buf1  g4039(.din(new_new_n3574__), .dout(new_new_n5501__));
  buf1  g4040(.din(new_new_n3577__), .dout(new_new_n5502__));
  buf1  g4041(.din(new_new_n3600__), .dout(new_new_n5503__));
  buf1  g4042(.din(new_new_n3606__), .dout(new_new_n5504__));
  buf1  g4043(.din(new_new_n5504__), .dout(new_new_n5505__));
  buf1  g4044(.din(new_new_n5505__), .dout(new_new_n5506__));
  buf1  g4045(.din(new_new_n5506__), .dout(new_new_n5507__));
  buf1  g4046(.din(new_new_n5506__), .dout(new_new_n5508__));
  buf1  g4047(.din(new_new_n5505__), .dout(new_new_n5509__));
  buf1  g4048(.din(new_new_n5509__), .dout(new_new_n5510__));
  buf1  g4049(.din(new_new_n5509__), .dout(new_new_n5511__));
  buf1  g4050(.din(new_new_n5504__), .dout(new_new_n5512__));
  buf1  g4051(.din(new_new_n5512__), .dout(new_new_n5513__));
  buf1  g4052(.din(new_new_n5512__), .dout(new_new_n5514__));
  buf1  g4053(.din(new_new_n3607__), .dout(new_new_n5515__));
  buf1  g4054(.din(new_new_n5515__), .dout(new_new_n5516__));
  buf1  g4055(.din(new_new_n5516__), .dout(new_new_n5517__));
  buf1  g4056(.din(new_new_n5517__), .dout(new_new_n5518__));
  buf1  g4057(.din(new_new_n5517__), .dout(new_new_n5519__));
  buf1  g4058(.din(new_new_n5516__), .dout(new_new_n5520__));
  buf1  g4059(.din(new_new_n5520__), .dout(new_new_n5521__));
  buf1  g4060(.din(new_new_n5520__), .dout(new_new_n5522__));
  buf1  g4061(.din(new_new_n5515__), .dout(new_new_n5523__));
  buf1  g4062(.din(new_new_n5523__), .dout(new_new_n5524__));
  buf1  g4063(.din(new_new_n5523__), .dout(new_new_n5525__));
  buf1  g4064(.din(new_new_n3610__), .dout(new_new_n5526__));
  buf1  g4065(.din(new_new_n5526__), .dout(new_new_n5527__));
  buf1  g4066(.din(new_new_n5527__), .dout(new_new_n5528__));
  buf1  g4067(.din(new_new_n5528__), .dout(new_new_n5529__));
  buf1  g4068(.din(new_new_n5528__), .dout(new_new_n5530__));
  buf1  g4069(.din(new_new_n5527__), .dout(new_new_n5531__));
  buf1  g4070(.din(new_new_n5531__), .dout(new_new_n5532__));
  buf1  g4071(.din(new_new_n5531__), .dout(new_new_n5533__));
  buf1  g4072(.din(new_new_n5526__), .dout(new_new_n5534__));
  buf1  g4073(.din(new_new_n5534__), .dout(new_new_n5535__));
  buf1  g4074(.din(new_new_n5534__), .dout(new_new_n5536__));
  buf1  g4075(.din(new_new_n3612__), .dout(new_new_n5537__));
  buf1  g4076(.din(new_new_n5537__), .dout(new_new_n5538__));
  buf1  g4077(.din(new_new_n5538__), .dout(new_new_n5539__));
  buf1  g4078(.din(new_new_n5539__), .dout(new_new_n5540__));
  buf1  g4079(.din(new_new_n5539__), .dout(new_new_n5541__));
  buf1  g4080(.din(new_new_n5538__), .dout(new_new_n5542__));
  buf1  g4081(.din(new_new_n5542__), .dout(new_new_n5543__));
  buf1  g4082(.din(new_new_n5542__), .dout(new_new_n5544__));
  buf1  g4083(.din(new_new_n5537__), .dout(new_new_n5545__));
  buf1  g4084(.din(new_new_n5545__), .dout(new_new_n5546__));
  buf1  g4085(.din(new_new_n5545__), .dout(new_new_n5547__));
  buf1  g4086(.din(new_new_n3614__), .dout(new_new_n5548__));
  buf1  g4087(.din(new_new_n5548__), .dout(new_new_n5549__));
  buf1  g4088(.din(new_new_n5549__), .dout(new_new_n5550__));
  buf1  g4089(.din(new_new_n5550__), .dout(new_new_n5551__));
  buf1  g4090(.din(new_new_n5550__), .dout(new_new_n5552__));
  buf1  g4091(.din(new_new_n5549__), .dout(new_new_n5553__));
  buf1  g4092(.din(new_new_n5553__), .dout(new_new_n5554__));
  buf1  g4093(.din(new_new_n5553__), .dout(new_new_n5555__));
  buf1  g4094(.din(new_new_n5548__), .dout(new_new_n5556__));
  buf1  g4095(.din(new_new_n5556__), .dout(new_new_n5557__));
  buf1  g4096(.din(new_new_n5556__), .dout(new_new_n5558__));
  buf1  g4097(.din(new_new_n3615__), .dout(new_new_n5559__));
  buf1  g4098(.din(new_new_n5559__), .dout(new_new_n5560__));
  buf1  g4099(.din(new_new_n5560__), .dout(new_new_n5561__));
  buf1  g4100(.din(new_new_n5561__), .dout(new_new_n5562__));
  buf1  g4101(.din(new_new_n5561__), .dout(new_new_n5563__));
  buf1  g4102(.din(new_new_n5560__), .dout(new_new_n5564__));
  buf1  g4103(.din(new_new_n5564__), .dout(new_new_n5565__));
  buf1  g4104(.din(new_new_n5564__), .dout(new_new_n5566__));
  buf1  g4105(.din(new_new_n5559__), .dout(new_new_n5567__));
  buf1  g4106(.din(new_new_n5567__), .dout(new_new_n5568__));
  buf1  g4107(.din(new_new_n5567__), .dout(new_new_n5569__));
  buf1  g4108(.din(new_new_n3616__), .dout(new_new_n5570__));
  buf1  g4109(.din(new_new_n5570__), .dout(new_new_n5571__));
  buf1  g4110(.din(new_new_n5571__), .dout(new_new_n5572__));
  buf1  g4111(.din(new_new_n5572__), .dout(new_new_n5573__));
  buf1  g4112(.din(new_new_n5572__), .dout(new_new_n5574__));
  buf1  g4113(.din(new_new_n5571__), .dout(new_new_n5575__));
  buf1  g4114(.din(new_new_n5575__), .dout(new_new_n5576__));
  buf1  g4115(.din(new_new_n5575__), .dout(new_new_n5577__));
  buf1  g4116(.din(new_new_n5570__), .dout(new_new_n5578__));
  buf1  g4117(.din(new_new_n5578__), .dout(new_new_n5579__));
  buf1  g4118(.din(new_new_n5578__), .dout(new_new_n5580__));
  buf1  g4119(.din(new_new_n3617__), .dout(new_new_n5581__));
  buf1  g4120(.din(new_new_n5581__), .dout(new_new_n5582__));
  buf1  g4121(.din(new_new_n5582__), .dout(new_new_n5583__));
  buf1  g4122(.din(new_new_n5583__), .dout(new_new_n5584__));
  buf1  g4123(.din(new_new_n5583__), .dout(new_new_n5585__));
  buf1  g4124(.din(new_new_n5582__), .dout(new_new_n5586__));
  buf1  g4125(.din(new_new_n5586__), .dout(new_new_n5587__));
  buf1  g4126(.din(new_new_n5586__), .dout(new_new_n5588__));
  buf1  g4127(.din(new_new_n5581__), .dout(new_new_n5589__));
  buf1  g4128(.din(new_new_n5589__), .dout(new_new_n5590__));
  buf1  g4129(.din(new_new_n5589__), .dout(new_new_n5591__));
  buf1  g4130(.din(new_new_n3625__), .dout(new_new_n5592__));
  buf1  g4131(.din(new_new_n5592__), .dout(new_new_n5593__));
  buf1  g4132(.din(new_new_n1147__), .dout(new_new_n5594__));
  buf1  g4133(.din(new_new_n5594__), .dout(new_new_n5595__));
  buf1  g4134(.din(new_new_n5594__), .dout(new_new_n5596__));
  buf1  g4135(.din(new_new_n1155__), .dout(new_new_n5597__));
  buf1  g4136(.din(new_new_n5597__), .dout(new_new_n5598__));
  buf1  g4137(.din(new_new_n5597__), .dout(new_new_n5599__));
  buf1  g4138(.din(new_new_n3642__), .dout(new_new_n5600__));
  buf1  g4139(.din(new_new_n3763__), .dout(new_new_n5601__));
  buf1  g4140(.din(new_new_n1145__), .dout(new_new_n5602__));
  buf1  g4141(.din(new_new_n5602__), .dout(new_new_n5603__));
  buf1  g4142(.din(new_new_n1153__), .dout(new_new_n5604__));
  buf1  g4143(.din(new_new_n5604__), .dout(new_new_n5605__));
  buf1  g4144(.din(new_new_n3777__), .dout(new_new_n5606__));
  buf1  g4145(.din(new_new_n3791__), .dout(new_new_n5607__));
  buf1  g4146(.din(new_new_n1131__), .dout(new_new_n5608__));
  buf1  g4147(.din(new_new_n3804__), .dout(new_new_n5609__));
  always @ (posedge clock) begin
    n1836_lo <= n8948;
    n1872_lo <= n8951;
    n1884_lo <= n8954;
    n1911_lo <= n8957;
    n1914_lo <= n8960;
    n1917_lo <= n8963;
    n1923_lo <= n8966;
    n1926_lo <= n8969;
    n1929_lo <= n8972;
    n1935_lo <= n8975;
    n1938_lo <= n8978;
    n1947_lo <= n8981;
    n1950_lo <= n8984;
    n1959_lo <= n8987;
    n1962_lo <= n8990;
    n1971_lo <= n8993;
    n1974_lo <= n8996;
    n1983_lo <= n8999;
    n1995_lo <= n9002;
    n2007_lo <= n9005;
    n2019_lo <= n9008;
    n2031_lo <= n9011;
    n2043_lo <= n9014;
    n2055_lo <= n9017;
    n2064_lo <= n9020;
    n2067_lo <= n9023;
    n2100_lo <= n9026;
    n2112_lo <= n9029;
    n2124_lo <= n9032;
    n2136_lo <= n9035;
    n2148_lo <= n9038;
    n2160_lo <= n9041;
    n2163_lo <= n9044;
    n2172_lo <= n9047;
    n2175_lo <= n9050;
    n2184_lo <= n9053;
    n2223_lo <= n9056;
    n2235_lo <= n9059;
    n2238_lo <= n9062;
    n2247_lo <= n9065;
    n2250_lo <= n9068;
    n2259_lo <= n9071;
    n2262_lo <= n9074;
    n2271_lo <= n9077;
    n2274_lo <= n9080;
    n2283_lo <= n9083;
    n2286_lo <= n9086;
    n2295_lo <= n9089;
    n2298_lo <= n9092;
    n2304_lo <= n9095;
    n2307_lo <= n9098;
    n2331_lo <= n9101;
    n2334_lo <= n9104;
    n2337_lo <= n9107;
    n2340_lo <= n9110;
    n3241_o2 <= n9113;
    n3242_o2 <= n9116;
    n3610_o2 <= n9119;
    n3980_o2 <= n9122;
    n3968_o2 <= n9125;
    n4298_o2 <= n9128;
    n4371_o2 <= n9131;
    n4413_o2 <= n9134;
    n4418_o2 <= n9137;
    n4628_o2 <= n9140;
    n4629_o2 <= n9143;
    n4633_o2 <= n9146;
    n4634_o2 <= n9149;
    n4732_o2 <= n9152;
    n4733_o2 <= n9155;
    n4884_o2 <= n9158;
    n4886_o2 <= n9161;
    n4890_o2 <= n9164;
    n5011_o2 <= n9167;
    n5012_o2 <= n9170;
    n5013_o2 <= n9173;
    n5014_o2 <= n9176;
    n5015_o2 <= n9179;
    n5021_o2 <= n9182;
    n5016_o2 <= n9185;
    n5026_o2 <= n9188;
    n4377_o2 <= n9191;
    n4378_o2 <= n9194;
    n4389_o2 <= n9197;
    n327_inv <= n9200;
    n330_inv <= n9203;
    n4398_o2 <= n9206;
    n4401_o2 <= n9209;
    n5117_o2 <= n9212;
    n5115_o2 <= n9215;
    n5122_o2 <= n9218;
    n5121_o2 <= n9221;
    n5119_o2 <= n9224;
    n5116_o2 <= n9227;
    n5123_o2 <= n9230;
    n5156_o2 <= n9233;
    n5167_o2 <= n9236;
    n4454_o2 <= n9239;
    n4455_o2 <= n9242;
    n4456_o2 <= n9245;
    n4505_o2 <= n9248;
    G742_o2 <= n9251;
    G727_o2 <= n9254;
    n4567_o2 <= n9257;
    n4568_o2 <= n9260;
    n4569_o2 <= n9263;
    n4571_o2 <= n9266;
    n4572_o2 <= n9269;
    n399_inv <= n9272;
    n4539_o2 <= n9275;
    n4651_o2 <= n9278;
    n4652_o2 <= n9281;
    n4653_o2 <= n9284;
    G1514_o2 <= n9287;
    G1823_o2 <= n9290;
    n4783_o2 <= n9293;
    n4787_o2 <= n9296;
    n426_inv <= n9299;
    n429_inv <= n9302;
    n4816_o2 <= n9305;
    n435_inv <= n9308;
    G572_o2 <= n9311;
    n4919_o2 <= n9314;
    n4920_o2 <= n9317;
    n4921_o2 <= n9320;
    G1048_o2 <= n9323;
    n5041_o2 <= n9326;
    n5094_o2 <= n9329;
    n5278_o2 <= n9332;
    n5301_o2 <= n9335;
    G2610_o2 <= n9338;
    G3174_o2 <= n9341;
    G3146_o2 <= n9344;
    G3217_o2 <= n9347;
    G3220_o2 <= n9350;
    G2839_o2 <= n9353;
    G3251_o2 <= n9356;
    G3042_o2 <= n9359;
    G3045_o2 <= n9362;
    G3262_o2 <= n9365;
    G2845_o2 <= n9368;
    G2929_o2 <= n9371;
    G2848_o2 <= n9374;
    G2851_o2 <= n9377;
    G3291_o2 <= n9380;
    G3254_o2 <= n9383;
    G2666_o2 <= n9386;
    n5099_o2 <= n9389;
    n5100_o2 <= n9392;
    n5101_o2 <= n9395;
    G2558_o2 <= n9398;
    n5266_o2 <= n9401;
    n5267_o2 <= n9404;
    G2759_o2 <= n9407;
    n537_inv <= n9410;
    n540_inv <= n9413;
    n543_inv <= n9416;
    n5292_o2 <= n9419;
    n5293_o2 <= n9422;
    n5294_o2 <= n9425;
    n5295_o2 <= n9428;
    G618_o2 <= n9431;
    G621_o2 <= n9434;
    G384_o2 <= n9437;
    G377_o2 <= n9440;
    n570_inv <= n9443;
    G3171_o2 <= n9446;
    G2552_o2 <= n9449;
    G3272_o2 <= n9452;
    G2015_o2 <= n9455;
    G3294_o2 <= n9458;
    G3281_o2 <= n9461;
    G3320_o2 <= n9464;
    G3275_o2 <= n9467;
    G3140_o2 <= n9470;
    G2836_o2 <= n9473;
    G2926_o2 <= n9476;
    G2842_o2 <= n9479;
    G3302_o2 <= n9482;
    G3288_o2 <= n9485;
    G3143_o2 <= n9488;
    G3100_o2 <= n9491;
    G2512_o2 <= n9494;
    n5325_o2 <= n9497;
    n5326_o2 <= n9500;
    n5327_o2 <= n9503;
    n1857_lo_buf_o2 <= n9506;
    n2097_lo_buf_o2 <= n9509;
    G2669_o2 <= n9512;
    n642_inv <= n9515;
    G568_o2 <= n9518;
    n648_inv <= n9521;
    G565_o2 <= n9524;
    G559_o2 <= n9527;
    n1821_lo_buf_o2 <= n9530;
    n1905_lo_buf_o2 <= n9533;
    n2133_lo_buf_o2 <= n9536;
    n2145_lo_buf_o2 <= n9539;
    n2157_lo_buf_o2 <= n9542;
    n2205_lo_buf_o2 <= n9545;
    n2217_lo_buf_o2 <= n9548;
    G447_o2 <= n9551;
    G434_o2 <= n9554;
    G422_o2 <= n9557;
    G461_o2 <= n9560;
    G3312_o2 <= n9563;
    G3332_o2 <= n9566;
    G3195_o2 <= n9569;
    G2607_o2 <= n9572;
    n702_inv <= n9575;
    G1005_o2 <= n9578;
    G1008_o2 <= n9581;
    n2001_lo_buf_o2 <= n9584;
    n2169_lo_buf_o2 <= n9587;
    n2229_lo_buf_o2 <= n9590;
    n2301_lo_buf_o2 <= n9593;
    n723_inv <= n9596;
    G2947_o2 <= n9599;
    n2013_lo_buf_o2 <= n9602;
    n2025_lo_buf_o2 <= n9605;
    n2037_lo_buf_o2 <= n9608;
    n2049_lo_buf_o2 <= n9611;
    n2181_lo_buf_o2 <= n9614;
    n744_inv <= n9617;
    n747_inv <= n9620;
    n750_inv <= n9623;
    n753_inv <= n9626;
    G3350_o2 <= n9629;
    G3360_o2 <= n9632;
    G3373_o2 <= n9635;
    G3237_o2 <= n9638;
    G2773_o2 <= n9641;
    G1733_o2 <= n9644;
    G1738_o2 <= n9647;
    G1751_o2 <= n9650;
    G2216_o2 <= n9653;
    G2219_o2 <= n9656;
    n786_inv <= n9659;
    n789_inv <= n9662;
    G787_o2 <= n9665;
    G2823_o2 <= n9668;
    G2796_o2 <= n9671;
    G875_o2 <= n9674;
    G2208_o2 <= n9677;
    G2211_o2 <= n9680;
    n1989_lo_buf_o2 <= n9683;
    n2061_lo_buf_o2 <= n9686;
    n2313_lo_buf_o2 <= n9689;
    G2232_o2 <= n9692;
    G1725_o2 <= n9695;
    G1764_o2 <= n9698;
    G2356_o2 <= n9701;
    G2359_o2 <= n9704;
    G1180_o2 <= n9707;
    G1756_o2 <= n9710;
    G2441_o2 <= n9713;
    G2887_o2 <= n9716;
    G2991_o2 <= n9719;
    n849_inv <= n9722;
    n852_inv <= n9725;
    n855_inv <= n9728;
    n858_inv <= n9731;
    n861_inv <= n9734;
    G2805_o2 <= n9737;
    G2906_o2 <= n9740;
    G2833_o2 <= n9743;
    n873_inv <= n9746;
    G3353_o2 <= n9749;
    G3367_o2 <= n9752;
    G3346_o2 <= n9755;
    G3340_o2 <= n9758;
    G3376_o2 <= n9761;
    G3359_o2 <= n9764;
    G3240_o2 <= n9767;
    G3344_o2 <= n9770;
    G2880_o2 <= n9773;
    G2939_o2 <= n9776;
    G2248_o2 <= n9779;
    G2251_o2 <= n9782;
    G2021_o2 <= n9785;
    G3383_o2 <= n9788;
    G3399_o2 <= n9791;
    G3404_o2 <= n9794;
    G3265_o2 <= n9797;
    G2866_o2 <= n9800;
    G2999_o2 <= n9803;
    G736_o2 <= n9806;
    G739_o2 <= n9809;
    G1200_o2 <= n9812;
    G1203_o2 <= n9815;
    G3027_o2 <= n9818;
    G1463_o2 <= n9821;
    G1460_o2 <= n9824;
    G3012_o2 <= n9827;
    G1574_o2 <= n9830;
    G1646_o2 <= n9833;
    G1592_o2 <= n9836;
    G1664_o2 <= n9839;
    G1547_o2 <= n9842;
    G1619_o2 <= n9845;
    G1556_o2 <= n9848;
    G1628_o2 <= n9851;
    G1583_o2 <= n9854;
    G1655_o2 <= n9857;
    G1529_o2 <= n9860;
    G1601_o2 <= n9863;
    G1538_o2 <= n9866;
    G1610_o2 <= n9869;
    G1565_o2 <= n9872;
    G1637_o2 <= n9875;
    G2437_o2 <= n9878;
    n1008_inv <= n9881;
    n1785_lo_buf_o2 <= n9884;
    n1845_lo_buf_o2 <= n9887;
    n1893_lo_buf_o2 <= n9890;
    n1941_lo_buf_o2 <= n9893;
    n1953_lo_buf_o2 <= n9896;
    n1965_lo_buf_o2 <= n9899;
    n1977_lo_buf_o2 <= n9902;
    n2241_lo_buf_o2 <= n9905;
    n2253_lo_buf_o2 <= n9908;
    n2265_lo_buf_o2 <= n9911;
    n2277_lo_buf_o2 <= n9914;
    n2289_lo_buf_o2 <= n9917;
    G519_o2 <= n9920;
    n1050_inv <= n9923;
    n1053_inv <= n9926;
    n1056_inv <= n9929;
    G1318_o2 <= n9932;
    n1062_inv <= n9935;
    G593_o2 <= n9938;
    n1068_inv <= n9941;
    n1071_inv <= n9944;
    n1074_inv <= n9947;
    G2284_o2 <= n9950;
    G2580_o2 <= n9953;
    G2302_o2 <= n9956;
    G2598_o2 <= n9959;
    G2497_o2 <= n9962;
    G2651_o2 <= n9965;
    G2296_o2 <= n9968;
    G2308_o2 <= n9971;
    G2592_o2 <= n9974;
    G2604_o2 <= n9977;
    G2902_o2 <= n9980;
    G2975_o2 <= n9983;
    G2962_o2 <= n9986;
    G3069_o2 <= n9989;
    G2018_o2 <= n9992;
    G1176_o2 <= n9995;
    G1189_o2 <= n9998;
    G3066_o2 <= n10001;
    G3137_o2 <= n10004;
    G3038_o2 <= n10007;
    G3117_o2 <= n10010;
    G2384_o2 <= n10013;
    G2472_o2 <= n10016;
    G772_o2 <= n10019;
    G935_o2 <= n10022;
    G2923_o2 <= n10025;
    G2971_o2 <= n10028;
    G2980_o2 <= n10031;
    G3039_o2 <= n10034;
    G2388_o2 <= n10037;
    G2287_o2 <= n10040;
    G3024_o2 <= n10043;
    G2916_o2 <= n10046;
    n1176_inv <= n10049;
    G3035_o2 <= n10052;
    G3107_o2 <= n10055;
    G1023_o2 <= n10058;
    G1024_o2 <= n10061;
    G1311_o2 <= n10064;
    G1312_o2 <= n10067;
    G3063_o2 <= n10070;
    G1520_o2 <= n10073;
    G1519_o2 <= n10076;
    G3078_o2 <= n10079;
    G2038_o2 <= n10082;
    G1848_o2 <= n10085;
    G1864_o2 <= n10088;
    G1872_o2 <= n10091;
    G1880_o2 <= n10094;
    G1888_o2 <= n10097;
    G1912_o2 <= n10100;
    G1928_o2 <= n10103;
    G1936_o2 <= n10106;
    G1944_o2 <= n10109;
    G1952_o2 <= n10112;
    G1850_o2 <= n10115;
    G1866_o2 <= n10118;
    G1874_o2 <= n10121;
    G1882_o2 <= n10124;
    G1890_o2 <= n10127;
    G1914_o2 <= n10130;
    G1930_o2 <= n10133;
    G1938_o2 <= n10136;
    G1946_o2 <= n10139;
    G1954_o2 <= n10142;
    G1845_o2 <= n10145;
    G1861_o2 <= n10148;
    G1869_o2 <= n10151;
    G1877_o2 <= n10154;
    G1885_o2 <= n10157;
    G1909_o2 <= n10160;
    G1925_o2 <= n10163;
    G1933_o2 <= n10166;
    G1941_o2 <= n10169;
    G1949_o2 <= n10172;
    G1846_o2 <= n10175;
    G1862_o2 <= n10178;
    G1870_o2 <= n10181;
    G1878_o2 <= n10184;
    G1886_o2 <= n10187;
    G1910_o2 <= n10190;
    G1926_o2 <= n10193;
    G1934_o2 <= n10196;
    G1942_o2 <= n10199;
    G1950_o2 <= n10202;
    G1849_o2 <= n10205;
    G1865_o2 <= n10208;
    G1873_o2 <= n10211;
    G1881_o2 <= n10214;
    G1889_o2 <= n10217;
    G1913_o2 <= n10220;
    G1929_o2 <= n10223;
    G1937_o2 <= n10226;
    G1945_o2 <= n10229;
    G1953_o2 <= n10232;
    G1843_o2 <= n10235;
    G1859_o2 <= n10238;
    G1867_o2 <= n10241;
    G1875_o2 <= n10244;
    G1883_o2 <= n10247;
    G1907_o2 <= n10250;
    G1923_o2 <= n10253;
    G1931_o2 <= n10256;
    G1939_o2 <= n10259;
    G1947_o2 <= n10262;
    G1844_o2 <= n10265;
    G1860_o2 <= n10268;
    G1868_o2 <= n10271;
    G1876_o2 <= n10274;
    G1884_o2 <= n10277;
    G1908_o2 <= n10280;
    G1924_o2 <= n10283;
    G1932_o2 <= n10286;
    G1940_o2 <= n10289;
    G1948_o2 <= n10292;
    G1847_o2 <= n10295;
    G1863_o2 <= n10298;
    G1871_o2 <= n10301;
    G1879_o2 <= n10304;
    G1887_o2 <= n10307;
    G1911_o2 <= n10310;
    G1927_o2 <= n10313;
    G1935_o2 <= n10316;
    G1943_o2 <= n10319;
    G1951_o2 <= n10322;
    G2444_o2 <= n10325;
    G2451_o2 <= n10328;
    G2502_o2 <= n10331;
    G2507_o2 <= n10334;
    n1464_inv <= n10337;
    G2583_o2 <= n10340;
    n1797_lo_buf_o2 <= n10343;
    n1833_lo_buf_o2 <= n10346;
    n1881_lo_buf_o2 <= n10349;
    n1479_inv <= n10352;
    n1482_inv <= n10355;
    n1485_inv <= n10358;
    G615_o2 <= n10361;
    G2254_o2 <= n10364;
    G2255_o2 <= n10367;
    G2027_o2 <= n10370;
    G2393_o2 <= n10373;
    G527_o2 <= n10376;
    G594_o2 <= n10379;
    G1689_o2 <= n10382;
    G1693_o2 <= n10385;
    G2281_o2 <= n10388;
    G2014_o2 <= n10391;
    G2459_o2 <= n10394;
    G2561_o2 <= n10397;
    G2533_o2 <= n10400;
    n1749_lo_buf_o2 <= n10403;
    n1761_lo_buf_o2 <= n10406;
    n1773_lo_buf_o2 <= n10409;
    n1809_lo_buf_o2 <= n10412;
    G1955_o2 <= n10415;
    G1958_o2 <= n10418;
    G2562_o2 <= n10421;
    G2398_o2 <= n10424;
    n1554_inv <= n10427;
    n1557_inv <= n10430;
    G2577_o2 <= n10433;
    G2627_o2 <= n10436;
    G654_o2 <= n10439;
    G660_o2 <= n10442;
    G831_o2 <= n10445;
    G919_o2 <= n10448;
    G925_o2 <= n10451;
    n1815_lo_buf_o2 <= n10454;
    n1899_lo_buf_o2 <= n10457;
    n2079_lo_buf_o2 <= n10460;
    n2127_lo_buf_o2 <= n10463;
    n2139_lo_buf_o2 <= n10466;
    n2151_lo_buf_o2 <= n10469;
    n2187_lo_buf_o2 <= n10472;
    n2199_lo_buf_o2 <= n10475;
    n2211_lo_buf_o2 <= n10478;
    G533_o2 <= n10481;
    n1854_lo_buf_o2 <= n10484;
    n2094_lo_buf_o2 <= n10487;
    G667_o2 <= n10490;
    G874_o2 <= n10493;
    G851_o2 <= n10496;
    G1127_o2 <= n10499;
    n1869_lo_buf_o2 <= n10502;
    n2109_lo_buf_o2 <= n10505;
    n2121_lo_buf_o2 <= n10508;
    G477_o2 <= n10511;
    G491_o2 <= n10514;
    G501_o2 <= n10517;
    G786_o2 <= n10520;
    G791_o2 <= n10523;
    G1126_o2 <= n10526;
    G1052_o2 <= n10529;
    G1054_o2 <= n10532;
  end
  initial begin
    n1836_lo <= 1'b0;
    n1872_lo <= 1'b0;
    n1884_lo <= 1'b0;
    n1911_lo <= 1'b0;
    n1914_lo <= 1'b0;
    n1917_lo <= 1'b0;
    n1923_lo <= 1'b0;
    n1926_lo <= 1'b0;
    n1929_lo <= 1'b0;
    n1935_lo <= 1'b0;
    n1938_lo <= 1'b0;
    n1947_lo <= 1'b0;
    n1950_lo <= 1'b0;
    n1959_lo <= 1'b0;
    n1962_lo <= 1'b0;
    n1971_lo <= 1'b0;
    n1974_lo <= 1'b0;
    n1983_lo <= 1'b0;
    n1995_lo <= 1'b0;
    n2007_lo <= 1'b0;
    n2019_lo <= 1'b0;
    n2031_lo <= 1'b0;
    n2043_lo <= 1'b0;
    n2055_lo <= 1'b0;
    n2064_lo <= 1'b0;
    n2067_lo <= 1'b0;
    n2100_lo <= 1'b0;
    n2112_lo <= 1'b0;
    n2124_lo <= 1'b0;
    n2136_lo <= 1'b0;
    n2148_lo <= 1'b0;
    n2160_lo <= 1'b0;
    n2163_lo <= 1'b0;
    n2172_lo <= 1'b0;
    n2175_lo <= 1'b0;
    n2184_lo <= 1'b0;
    n2223_lo <= 1'b0;
    n2235_lo <= 1'b0;
    n2238_lo <= 1'b0;
    n2247_lo <= 1'b0;
    n2250_lo <= 1'b0;
    n2259_lo <= 1'b0;
    n2262_lo <= 1'b0;
    n2271_lo <= 1'b0;
    n2274_lo <= 1'b0;
    n2283_lo <= 1'b0;
    n2286_lo <= 1'b0;
    n2295_lo <= 1'b0;
    n2298_lo <= 1'b0;
    n2304_lo <= 1'b0;
    n2307_lo <= 1'b0;
    n2331_lo <= 1'b0;
    n2334_lo <= 1'b0;
    n2337_lo <= 1'b0;
    n2340_lo <= 1'b0;
    n3241_o2 <= 1'b0;
    n3242_o2 <= 1'b0;
    n3610_o2 <= 1'b0;
    n3980_o2 <= 1'b0;
    n3968_o2 <= 1'b0;
    n4298_o2 <= 1'b0;
    n4371_o2 <= 1'b0;
    n4413_o2 <= 1'b0;
    n4418_o2 <= 1'b0;
    n4628_o2 <= 1'b0;
    n4629_o2 <= 1'b0;
    n4633_o2 <= 1'b0;
    n4634_o2 <= 1'b0;
    n4732_o2 <= 1'b0;
    n4733_o2 <= 1'b0;
    n4884_o2 <= 1'b0;
    n4886_o2 <= 1'b0;
    n4890_o2 <= 1'b0;
    n5011_o2 <= 1'b0;
    n5012_o2 <= 1'b0;
    n5013_o2 <= 1'b0;
    n5014_o2 <= 1'b0;
    n5015_o2 <= 1'b0;
    n5021_o2 <= 1'b0;
    n5016_o2 <= 1'b0;
    n5026_o2 <= 1'b0;
    n4377_o2 <= 1'b0;
    n4378_o2 <= 1'b0;
    n4389_o2 <= 1'b0;
    n327_inv <= 1'b0;
    n330_inv <= 1'b0;
    n4398_o2 <= 1'b0;
    n4401_o2 <= 1'b0;
    n5117_o2 <= 1'b0;
    n5115_o2 <= 1'b0;
    n5122_o2 <= 1'b0;
    n5121_o2 <= 1'b0;
    n5119_o2 <= 1'b0;
    n5116_o2 <= 1'b0;
    n5123_o2 <= 1'b0;
    n5156_o2 <= 1'b0;
    n5167_o2 <= 1'b0;
    n4454_o2 <= 1'b0;
    n4455_o2 <= 1'b0;
    n4456_o2 <= 1'b0;
    n4505_o2 <= 1'b0;
    G742_o2 <= 1'b0;
    G727_o2 <= 1'b0;
    n4567_o2 <= 1'b0;
    n4568_o2 <= 1'b0;
    n4569_o2 <= 1'b0;
    n4571_o2 <= 1'b0;
    n4572_o2 <= 1'b0;
    n399_inv <= 1'b0;
    n4539_o2 <= 1'b0;
    n4651_o2 <= 1'b0;
    n4652_o2 <= 1'b0;
    n4653_o2 <= 1'b0;
    G1514_o2 <= 1'b0;
    G1823_o2 <= 1'b0;
    n4783_o2 <= 1'b0;
    n4787_o2 <= 1'b0;
    n426_inv <= 1'b0;
    n429_inv <= 1'b0;
    n4816_o2 <= 1'b0;
    n435_inv <= 1'b0;
    G572_o2 <= 1'b0;
    n4919_o2 <= 1'b0;
    n4920_o2 <= 1'b0;
    n4921_o2 <= 1'b0;
    G1048_o2 <= 1'b0;
    n5041_o2 <= 1'b0;
    n5094_o2 <= 1'b0;
    n5278_o2 <= 1'b0;
    n5301_o2 <= 1'b0;
    G2610_o2 <= 1'b0;
    G3174_o2 <= 1'b0;
    G3146_o2 <= 1'b0;
    G3217_o2 <= 1'b0;
    G3220_o2 <= 1'b0;
    G2839_o2 <= 1'b0;
    G3251_o2 <= 1'b0;
    G3042_o2 <= 1'b0;
    G3045_o2 <= 1'b0;
    G3262_o2 <= 1'b0;
    G2845_o2 <= 1'b0;
    G2929_o2 <= 1'b0;
    G2848_o2 <= 1'b0;
    G2851_o2 <= 1'b0;
    G3291_o2 <= 1'b0;
    G3254_o2 <= 1'b0;
    G2666_o2 <= 1'b0;
    n5099_o2 <= 1'b0;
    n5100_o2 <= 1'b0;
    n5101_o2 <= 1'b0;
    G2558_o2 <= 1'b0;
    n5266_o2 <= 1'b0;
    n5267_o2 <= 1'b0;
    G2759_o2 <= 1'b0;
    n537_inv <= 1'b0;
    n540_inv <= 1'b0;
    n543_inv <= 1'b0;
    n5292_o2 <= 1'b0;
    n5293_o2 <= 1'b0;
    n5294_o2 <= 1'b0;
    n5295_o2 <= 1'b0;
    G618_o2 <= 1'b0;
    G621_o2 <= 1'b0;
    G384_o2 <= 1'b0;
    G377_o2 <= 1'b0;
    n570_inv <= 1'b0;
    G3171_o2 <= 1'b0;
    G2552_o2 <= 1'b0;
    G3272_o2 <= 1'b0;
    G2015_o2 <= 1'b0;
    G3294_o2 <= 1'b0;
    G3281_o2 <= 1'b0;
    G3320_o2 <= 1'b0;
    G3275_o2 <= 1'b0;
    G3140_o2 <= 1'b0;
    G2836_o2 <= 1'b0;
    G2926_o2 <= 1'b0;
    G2842_o2 <= 1'b0;
    G3302_o2 <= 1'b0;
    G3288_o2 <= 1'b0;
    G3143_o2 <= 1'b0;
    G3100_o2 <= 1'b0;
    G2512_o2 <= 1'b0;
    n5325_o2 <= 1'b0;
    n5326_o2 <= 1'b0;
    n5327_o2 <= 1'b0;
    n1857_lo_buf_o2 <= 1'b0;
    n2097_lo_buf_o2 <= 1'b0;
    G2669_o2 <= 1'b0;
    n642_inv <= 1'b0;
    G568_o2 <= 1'b0;
    n648_inv <= 1'b0;
    G565_o2 <= 1'b0;
    G559_o2 <= 1'b0;
    n1821_lo_buf_o2 <= 1'b0;
    n1905_lo_buf_o2 <= 1'b0;
    n2133_lo_buf_o2 <= 1'b0;
    n2145_lo_buf_o2 <= 1'b0;
    n2157_lo_buf_o2 <= 1'b0;
    n2205_lo_buf_o2 <= 1'b0;
    n2217_lo_buf_o2 <= 1'b0;
    G447_o2 <= 1'b0;
    G434_o2 <= 1'b0;
    G422_o2 <= 1'b0;
    G461_o2 <= 1'b0;
    G3312_o2 <= 1'b0;
    G3332_o2 <= 1'b0;
    G3195_o2 <= 1'b0;
    G2607_o2 <= 1'b0;
    n702_inv <= 1'b0;
    G1005_o2 <= 1'b0;
    G1008_o2 <= 1'b0;
    n2001_lo_buf_o2 <= 1'b0;
    n2169_lo_buf_o2 <= 1'b0;
    n2229_lo_buf_o2 <= 1'b0;
    n2301_lo_buf_o2 <= 1'b0;
    n723_inv <= 1'b0;
    G2947_o2 <= 1'b0;
    n2013_lo_buf_o2 <= 1'b0;
    n2025_lo_buf_o2 <= 1'b0;
    n2037_lo_buf_o2 <= 1'b0;
    n2049_lo_buf_o2 <= 1'b0;
    n2181_lo_buf_o2 <= 1'b0;
    n744_inv <= 1'b0;
    n747_inv <= 1'b0;
    n750_inv <= 1'b0;
    n753_inv <= 1'b0;
    G3350_o2 <= 1'b0;
    G3360_o2 <= 1'b0;
    G3373_o2 <= 1'b0;
    G3237_o2 <= 1'b0;
    G2773_o2 <= 1'b0;
    G1733_o2 <= 1'b0;
    G1738_o2 <= 1'b0;
    G1751_o2 <= 1'b0;
    G2216_o2 <= 1'b0;
    G2219_o2 <= 1'b0;
    n786_inv <= 1'b0;
    n789_inv <= 1'b0;
    G787_o2 <= 1'b0;
    G2823_o2 <= 1'b0;
    G2796_o2 <= 1'b0;
    G875_o2 <= 1'b0;
    G2208_o2 <= 1'b0;
    G2211_o2 <= 1'b0;
    n1989_lo_buf_o2 <= 1'b0;
    n2061_lo_buf_o2 <= 1'b0;
    n2313_lo_buf_o2 <= 1'b0;
    G2232_o2 <= 1'b0;
    G1725_o2 <= 1'b0;
    G1764_o2 <= 1'b0;
    G2356_o2 <= 1'b0;
    G2359_o2 <= 1'b0;
    G1180_o2 <= 1'b0;
    G1756_o2 <= 1'b0;
    G2441_o2 <= 1'b0;
    G2887_o2 <= 1'b0;
    G2991_o2 <= 1'b0;
    n849_inv <= 1'b0;
    n852_inv <= 1'b0;
    n855_inv <= 1'b0;
    n858_inv <= 1'b0;
    n861_inv <= 1'b0;
    G2805_o2 <= 1'b0;
    G2906_o2 <= 1'b0;
    G2833_o2 <= 1'b0;
    n873_inv <= 1'b0;
    G3353_o2 <= 1'b0;
    G3367_o2 <= 1'b0;
    G3346_o2 <= 1'b0;
    G3340_o2 <= 1'b0;
    G3376_o2 <= 1'b0;
    G3359_o2 <= 1'b0;
    G3240_o2 <= 1'b0;
    G3344_o2 <= 1'b0;
    G2880_o2 <= 1'b0;
    G2939_o2 <= 1'b0;
    G2248_o2 <= 1'b0;
    G2251_o2 <= 1'b0;
    G2021_o2 <= 1'b0;
    G3383_o2 <= 1'b0;
    G3399_o2 <= 1'b0;
    G3404_o2 <= 1'b0;
    G3265_o2 <= 1'b0;
    G2866_o2 <= 1'b0;
    G2999_o2 <= 1'b0;
    G736_o2 <= 1'b0;
    G739_o2 <= 1'b0;
    G1200_o2 <= 1'b0;
    G1203_o2 <= 1'b0;
    G3027_o2 <= 1'b0;
    G1463_o2 <= 1'b0;
    G1460_o2 <= 1'b0;
    G3012_o2 <= 1'b0;
    G1574_o2 <= 1'b0;
    G1646_o2 <= 1'b0;
    G1592_o2 <= 1'b0;
    G1664_o2 <= 1'b0;
    G1547_o2 <= 1'b0;
    G1619_o2 <= 1'b0;
    G1556_o2 <= 1'b0;
    G1628_o2 <= 1'b0;
    G1583_o2 <= 1'b0;
    G1655_o2 <= 1'b0;
    G1529_o2 <= 1'b0;
    G1601_o2 <= 1'b0;
    G1538_o2 <= 1'b0;
    G1610_o2 <= 1'b0;
    G1565_o2 <= 1'b0;
    G1637_o2 <= 1'b0;
    G2437_o2 <= 1'b0;
    n1008_inv <= 1'b0;
    n1785_lo_buf_o2 <= 1'b0;
    n1845_lo_buf_o2 <= 1'b0;
    n1893_lo_buf_o2 <= 1'b0;
    n1941_lo_buf_o2 <= 1'b0;
    n1953_lo_buf_o2 <= 1'b0;
    n1965_lo_buf_o2 <= 1'b0;
    n1977_lo_buf_o2 <= 1'b0;
    n2241_lo_buf_o2 <= 1'b0;
    n2253_lo_buf_o2 <= 1'b0;
    n2265_lo_buf_o2 <= 1'b0;
    n2277_lo_buf_o2 <= 1'b0;
    n2289_lo_buf_o2 <= 1'b0;
    G519_o2 <= 1'b0;
    n1050_inv <= 1'b0;
    n1053_inv <= 1'b0;
    n1056_inv <= 1'b0;
    G1318_o2 <= 1'b0;
    n1062_inv <= 1'b0;
    G593_o2 <= 1'b0;
    n1068_inv <= 1'b0;
    n1071_inv <= 1'b0;
    n1074_inv <= 1'b0;
    G2284_o2 <= 1'b0;
    G2580_o2 <= 1'b0;
    G2302_o2 <= 1'b0;
    G2598_o2 <= 1'b0;
    G2497_o2 <= 1'b0;
    G2651_o2 <= 1'b0;
    G2296_o2 <= 1'b0;
    G2308_o2 <= 1'b0;
    G2592_o2 <= 1'b0;
    G2604_o2 <= 1'b0;
    G2902_o2 <= 1'b0;
    G2975_o2 <= 1'b0;
    G2962_o2 <= 1'b0;
    G3069_o2 <= 1'b0;
    G2018_o2 <= 1'b0;
    G1176_o2 <= 1'b0;
    G1189_o2 <= 1'b0;
    G3066_o2 <= 1'b0;
    G3137_o2 <= 1'b0;
    G3038_o2 <= 1'b0;
    G3117_o2 <= 1'b0;
    G2384_o2 <= 1'b0;
    G2472_o2 <= 1'b0;
    G772_o2 <= 1'b0;
    G935_o2 <= 1'b0;
    G2923_o2 <= 1'b0;
    G2971_o2 <= 1'b0;
    G2980_o2 <= 1'b0;
    G3039_o2 <= 1'b0;
    G2388_o2 <= 1'b0;
    G2287_o2 <= 1'b0;
    G3024_o2 <= 1'b0;
    G2916_o2 <= 1'b0;
    n1176_inv <= 1'b0;
    G3035_o2 <= 1'b0;
    G3107_o2 <= 1'b0;
    G1023_o2 <= 1'b0;
    G1024_o2 <= 1'b0;
    G1311_o2 <= 1'b0;
    G1312_o2 <= 1'b0;
    G3063_o2 <= 1'b0;
    G1520_o2 <= 1'b0;
    G1519_o2 <= 1'b0;
    G3078_o2 <= 1'b0;
    G2038_o2 <= 1'b0;
    G1848_o2 <= 1'b0;
    G1864_o2 <= 1'b0;
    G1872_o2 <= 1'b0;
    G1880_o2 <= 1'b0;
    G1888_o2 <= 1'b0;
    G1912_o2 <= 1'b0;
    G1928_o2 <= 1'b0;
    G1936_o2 <= 1'b0;
    G1944_o2 <= 1'b0;
    G1952_o2 <= 1'b0;
    G1850_o2 <= 1'b0;
    G1866_o2 <= 1'b0;
    G1874_o2 <= 1'b0;
    G1882_o2 <= 1'b0;
    G1890_o2 <= 1'b0;
    G1914_o2 <= 1'b0;
    G1930_o2 <= 1'b0;
    G1938_o2 <= 1'b0;
    G1946_o2 <= 1'b0;
    G1954_o2 <= 1'b0;
    G1845_o2 <= 1'b0;
    G1861_o2 <= 1'b0;
    G1869_o2 <= 1'b0;
    G1877_o2 <= 1'b0;
    G1885_o2 <= 1'b0;
    G1909_o2 <= 1'b0;
    G1925_o2 <= 1'b0;
    G1933_o2 <= 1'b0;
    G1941_o2 <= 1'b0;
    G1949_o2 <= 1'b0;
    G1846_o2 <= 1'b0;
    G1862_o2 <= 1'b0;
    G1870_o2 <= 1'b0;
    G1878_o2 <= 1'b0;
    G1886_o2 <= 1'b0;
    G1910_o2 <= 1'b0;
    G1926_o2 <= 1'b0;
    G1934_o2 <= 1'b0;
    G1942_o2 <= 1'b0;
    G1950_o2 <= 1'b0;
    G1849_o2 <= 1'b0;
    G1865_o2 <= 1'b0;
    G1873_o2 <= 1'b0;
    G1881_o2 <= 1'b0;
    G1889_o2 <= 1'b0;
    G1913_o2 <= 1'b0;
    G1929_o2 <= 1'b0;
    G1937_o2 <= 1'b0;
    G1945_o2 <= 1'b0;
    G1953_o2 <= 1'b0;
    G1843_o2 <= 1'b0;
    G1859_o2 <= 1'b0;
    G1867_o2 <= 1'b0;
    G1875_o2 <= 1'b0;
    G1883_o2 <= 1'b0;
    G1907_o2 <= 1'b0;
    G1923_o2 <= 1'b0;
    G1931_o2 <= 1'b0;
    G1939_o2 <= 1'b0;
    G1947_o2 <= 1'b0;
    G1844_o2 <= 1'b0;
    G1860_o2 <= 1'b0;
    G1868_o2 <= 1'b0;
    G1876_o2 <= 1'b0;
    G1884_o2 <= 1'b0;
    G1908_o2 <= 1'b0;
    G1924_o2 <= 1'b0;
    G1932_o2 <= 1'b0;
    G1940_o2 <= 1'b0;
    G1948_o2 <= 1'b0;
    G1847_o2 <= 1'b0;
    G1863_o2 <= 1'b0;
    G1871_o2 <= 1'b0;
    G1879_o2 <= 1'b0;
    G1887_o2 <= 1'b0;
    G1911_o2 <= 1'b0;
    G1927_o2 <= 1'b0;
    G1935_o2 <= 1'b0;
    G1943_o2 <= 1'b0;
    G1951_o2 <= 1'b0;
    G2444_o2 <= 1'b0;
    G2451_o2 <= 1'b0;
    G2502_o2 <= 1'b0;
    G2507_o2 <= 1'b0;
    n1464_inv <= 1'b0;
    G2583_o2 <= 1'b0;
    n1797_lo_buf_o2 <= 1'b0;
    n1833_lo_buf_o2 <= 1'b0;
    n1881_lo_buf_o2 <= 1'b0;
    n1479_inv <= 1'b0;
    n1482_inv <= 1'b0;
    n1485_inv <= 1'b0;
    G615_o2 <= 1'b0;
    G2254_o2 <= 1'b0;
    G2255_o2 <= 1'b0;
    G2027_o2 <= 1'b0;
    G2393_o2 <= 1'b0;
    G527_o2 <= 1'b0;
    G594_o2 <= 1'b0;
    G1689_o2 <= 1'b0;
    G1693_o2 <= 1'b0;
    G2281_o2 <= 1'b0;
    G2014_o2 <= 1'b0;
    G2459_o2 <= 1'b0;
    G2561_o2 <= 1'b0;
    G2533_o2 <= 1'b0;
    n1749_lo_buf_o2 <= 1'b0;
    n1761_lo_buf_o2 <= 1'b0;
    n1773_lo_buf_o2 <= 1'b0;
    n1809_lo_buf_o2 <= 1'b0;
    G1955_o2 <= 1'b0;
    G1958_o2 <= 1'b0;
    G2562_o2 <= 1'b0;
    G2398_o2 <= 1'b0;
    n1554_inv <= 1'b0;
    n1557_inv <= 1'b0;
    G2577_o2 <= 1'b0;
    G2627_o2 <= 1'b0;
    G654_o2 <= 1'b0;
    G660_o2 <= 1'b0;
    G831_o2 <= 1'b0;
    G919_o2 <= 1'b0;
    G925_o2 <= 1'b0;
    n1815_lo_buf_o2 <= 1'b0;
    n1899_lo_buf_o2 <= 1'b0;
    n2079_lo_buf_o2 <= 1'b0;
    n2127_lo_buf_o2 <= 1'b0;
    n2139_lo_buf_o2 <= 1'b0;
    n2151_lo_buf_o2 <= 1'b0;
    n2187_lo_buf_o2 <= 1'b0;
    n2199_lo_buf_o2 <= 1'b0;
    n2211_lo_buf_o2 <= 1'b0;
    G533_o2 <= 1'b0;
    n1854_lo_buf_o2 <= 1'b0;
    n2094_lo_buf_o2 <= 1'b0;
    G667_o2 <= 1'b0;
    G874_o2 <= 1'b0;
    G851_o2 <= 1'b0;
    G1127_o2 <= 1'b0;
    n1869_lo_buf_o2 <= 1'b0;
    n2109_lo_buf_o2 <= 1'b0;
    n2121_lo_buf_o2 <= 1'b0;
    G477_o2 <= 1'b0;
    G491_o2 <= 1'b0;
    G501_o2 <= 1'b0;
    G786_o2 <= 1'b0;
    G791_o2 <= 1'b0;
    G1126_o2 <= 1'b0;
    G1052_o2 <= 1'b0;
    G1054_o2 <= 1'b0;
  end
endmodule


