// Benchmark "c6288" written by ABC on Sun Oct 29 16:27:02 2023

module c6288_pclk (  clk,
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32,
    G6257, G6258, G6259, G6260, G6261, G6262, G6263, G6264, G6265, G6266,
    G6267, G6268, G6269, G6270, G6271, G6272, G6273, G6274, G6275, G6276,
    G6277, G6278, G6279, G6280, G6281, G6282, G6283, G6284, G6285, G6286,
    G6287, G6288  );
  
  input clk, G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32;
  output G6257, G6258, G6259, G6260, G6261, G6262, G6263, G6264, G6265, G6266,
    G6267, G6268, G6269, G6270, G6271, G6272, G6273, G6274, G6275, G6276,
    G6277, G6278, G6279, G6280, G6281, G6282, G6283, G6284, G6285, G6286,
    G6287, G6288;
  reg n2482_lo, n2485_lo, n2488_lo, n2491_lo, n2494_lo, n2497_lo, n2500_lo,
    n2503_lo, n2506_lo, n2509_lo, n2512_lo, n2515_lo, n2518_lo, n2521_lo,
    n2524_lo, n2527_lo, n2530_lo, n2533_lo, n2536_lo, n2539_lo, n2542_lo,
    n2545_lo, n2548_lo, n2551_lo, n2554_lo, n2557_lo, n2560_lo, n2563_lo,
    n2566_lo, n2569_lo, n2572_lo, n2575_lo, n2578_lo, n2581_lo, n2584_lo,
    n2587_lo, n2590_lo, n2593_lo, n2596_lo, n2599_lo, n2602_lo, n2605_lo,
    n2608_lo, n2611_lo, n2614_lo, n2617_lo, n2620_lo, n2623_lo, n2626_lo,
    n2629_lo, n2632_lo, n2635_lo, n2638_lo, n2641_lo, n2644_lo, n2647_lo,
    n2650_lo, n2653_lo, n2656_lo, n2659_lo, n2662_lo, n2665_lo, n2668_lo,
    n2671_lo, n2674_lo, n2677_lo, n2680_lo, n2683_lo, n2686_lo, n2689_lo,
    n2692_lo, n2695_lo, n2698_lo, n2701_lo, n2704_lo, n2707_lo, n2710_lo,
    n2713_lo, n2716_lo, n2719_lo, n2722_lo, n2725_lo, n2728_lo, n2731_lo,
    n2734_lo, n2737_lo, n2740_lo, n2743_lo, n2746_lo, n2749_lo, n2752_lo,
    n2755_lo, n2758_lo, n2761_lo, n2764_lo, n2767_lo, n2770_lo, n2773_lo,
    n2776_lo, n2779_lo, n2782_lo, n2785_lo, n2788_lo, n2791_lo, n2794_lo,
    n2797_lo, n2800_lo, n2803_lo, n2806_lo, n2809_lo, n2812_lo, n2815_lo,
    n2818_lo, n2821_lo, n2824_lo, n2827_lo, n2830_lo, n2833_lo, n2836_lo,
    n2839_lo, n2842_lo, n2845_lo, n2848_lo, n2851_lo, n2854_lo, n2857_lo,
    n2860_lo, n2863_lo;
  wire new_G545_, new_G548_, new_G551_, new_G554_, new_G557_, new_G560_,
    new_G563_, new_G566_, new_G569_, new_G572_, new_G575_, new_G578_,
    new_G581_, new_G584_, new_G587_, new_G590_, new_G593_, new_G596_,
    new_G599_, new_G602_, new_G605_, new_G608_, new_G611_, new_G614_,
    new_G617_, new_G620_, new_G623_, new_G626_, new_G629_, new_G632_,
    new_G635_, new_G638_, new_G641_, new_G644_, new_G647_, new_G650_,
    new_G653_, new_G656_, new_G659_, new_G662_, new_G665_, new_G668_,
    new_G671_, new_G674_, new_G677_, new_G680_, new_G683_, new_G686_,
    new_G689_, new_G692_, new_G695_, new_G698_, new_G701_, new_G704_,
    new_G707_, new_G710_, new_G713_, new_G716_, new_G719_, new_G722_,
    new_G725_, new_G728_, new_G731_, new_G734_, new_G737_, new_G740_,
    new_G743_, new_G746_, new_G749_, new_G752_, new_G755_, new_G758_,
    new_G761_, new_G764_, new_G767_, new_G770_, new_G773_, new_G776_,
    new_G779_, new_G782_, new_G785_, new_G788_, new_G791_, new_G794_,
    new_G797_, new_G800_, new_G803_, new_G806_, new_G809_, new_G812_,
    new_G815_, new_G818_, new_G821_, new_G824_, new_G827_, new_G830_,
    new_G833_, new_G836_, new_G839_, new_G842_, new_G845_, new_G848_,
    new_G851_, new_G854_, new_G857_, new_G860_, new_G863_, new_G866_,
    new_G869_, new_G872_, new_G875_, new_G878_, new_G881_, new_G884_,
    new_G887_, new_G890_, new_G893_, new_G896_, new_G899_, new_G902_,
    new_G905_, new_G908_, new_G911_, new_G914_, new_G917_, new_G920_,
    new_G923_, new_G926_, new_G929_, new_G932_, new_G935_, new_G938_,
    new_G941_, new_G944_, new_G947_, new_G950_, new_G953_, new_G956_,
    new_G959_, new_G962_, new_G965_, new_G968_, new_G971_, new_G974_,
    new_G977_, new_G980_, new_G983_, new_G986_, new_G989_, new_G992_,
    new_G995_, new_G998_, new_G1001_, new_G1004_, new_G1007_, new_G1010_,
    new_G1013_, new_G1016_, new_G1019_, new_G1022_, new_G1025_, new_G1028_,
    new_G1031_, new_G1034_, new_G1037_, new_G1040_, new_G1043_, new_G1046_,
    new_G1049_, new_G1052_, new_G1055_, new_G1058_, new_G1061_, new_G1064_,
    new_G1067_, new_G1070_, new_G1073_, new_G1076_, new_G1079_, new_G1082_,
    new_G1085_, new_G1088_, new_G1091_, new_G1094_, new_G1097_, new_G1100_,
    new_G1103_, new_G1106_, new_G1109_, new_G1112_, new_G1115_, new_G1118_,
    new_G1121_, new_G1124_, new_G1127_, new_G1130_, new_G1133_, new_G1136_,
    new_G1139_, new_G1142_, new_G1145_, new_G1148_, new_G1151_, new_G1154_,
    new_G1157_, new_G1160_, new_G1163_, new_G1166_, new_G1169_, new_G1172_,
    new_G1175_, new_G1178_, new_G1181_, new_G1184_, new_G1187_, new_G1190_,
    new_G1193_, new_G1196_, new_G1199_, new_G1202_, new_G1205_, new_G1208_,
    new_G1211_, new_G1214_, new_G1217_, new_G1220_, new_G1223_, new_G1226_,
    new_G1229_, new_G1232_, new_G1235_, new_G1238_, new_G1241_, new_G1244_,
    new_G1247_, new_G1250_, new_G1253_, new_G1256_, new_G1259_, new_G1262_,
    new_G1265_, new_G1268_, new_G1271_, new_G1274_, new_G1277_, new_G1280_,
    new_G1283_, new_G1286_, new_G1289_, new_G1292_, new_G1295_, new_G1298_,
    new_G1301_, new_G1304_, new_G1307_, new_G1310_, new_G1314_, new_G1318_,
    new_G1322_, new_G1326_, new_G1330_, new_G1334_, new_G1338_, new_G1342_,
    new_G1346_, new_G1350_, new_G1354_, new_G1358_, new_G1362_, new_G1366_,
    new_G1370_, new_G1371_, new_G1372_, new_G1373_, new_G1374_, new_G1375_,
    new_G1376_, new_G1377_, new_G1378_, new_G1379_, new_G1380_, new_G1381_,
    new_G1382_, new_G1383_, new_G1384_, new_G1385_, new_G1386_, new_G1387_,
    new_G1388_, new_G1389_, new_G1390_, new_G1391_, new_G1392_, new_G1393_,
    new_G1394_, new_G1395_, new_G1396_, new_G1397_, new_G1398_, new_G1399_,
    new_G1400_, new_G1403_, new_G1406_, new_G1409_, new_G1412_, new_G1415_,
    new_G1418_, new_G1421_, new_G1424_, new_G1427_, new_G1430_, new_G1433_,
    new_G1436_, new_G1439_, new_G1442_, new_G1445_, new_G1449_, new_G1453_,
    new_G1457_, new_G1461_, new_G1465_, new_G1469_, new_G1473_, new_G1477_,
    new_G1481_, new_G1485_, new_G1489_, new_G1493_, new_G1497_, new_G1501_,
    new_G1505_, new_G1506_, new_G1507_, new_G1510_, new_G1511_, new_G1512_,
    new_G1515_, new_G1516_, new_G1517_, new_G1520_, new_G1521_, new_G1522_,
    new_G1525_, new_G1526_, new_G1527_, new_G1530_, new_G1531_, new_G1532_,
    new_G1535_, new_G1536_, new_G1537_, new_G1540_, new_G1541_, new_G1542_,
    new_G1545_, new_G1546_, new_G1547_, new_G1550_, new_G1551_, new_G1552_,
    new_G1555_, new_G1556_, new_G1557_, new_G1560_, new_G1561_, new_G1562_,
    new_G1565_, new_G1566_, new_G1567_, new_G1570_, new_G1571_, new_G1572_,
    new_G1575_, new_G1576_, new_G1577_, new_G1580_, new_G1583_, new_G1586_,
    new_G1589_, new_G1592_, new_G1595_, new_G1598_, new_G1601_, new_G1604_,
    new_G1607_, new_G1610_, new_G1613_, new_G1616_, new_G1619_, new_G1622_,
    new_G1626_, new_G1630_, new_G1634_, new_G1638_, new_G1642_, new_G1646_,
    new_G1650_, new_G1654_, new_G1658_, new_G1662_, new_G1666_, new_G1670_,
    new_G1674_, new_G1678_, new_G1682_, new_G1683_, new_G1684_, new_G1685_,
    new_G1686_, new_G1687_, new_G1688_, new_G1689_, new_G1690_, new_G1691_,
    new_G1692_, new_G1693_, new_G1694_, new_G1695_, new_G1696_, new_G1697_,
    new_G1698_, new_G1699_, new_G1700_, new_G1701_, new_G1702_, new_G1703_,
    new_G1704_, new_G1705_, new_G1706_, new_G1707_, new_G1708_, new_G1709_,
    new_G1710_, new_G1711_, new_G1712_, new_G1715_, new_G1718_, new_G1721_,
    new_G1724_, new_G1727_, new_G1730_, new_G1733_, new_G1736_, new_G1739_,
    new_G1742_, new_G1745_, new_G1748_, new_G1751_, new_G1754_, new_G1757_,
    new_G1761_, new_G1765_, new_G1769_, new_G1773_, new_G1777_, new_G1781_,
    new_G1785_, new_G1789_, new_G1793_, new_G1797_, new_G1801_, new_G1805_,
    new_G1809_, new_G1813_, new_G1817_, new_G1818_, new_G1819_, new_G1822_,
    new_G1823_, new_G1824_, new_G1827_, new_G1828_, new_G1829_, new_G1832_,
    new_G1833_, new_G1834_, new_G1837_, new_G1838_, new_G1839_, new_G1842_,
    new_G1843_, new_G1844_, new_G1847_, new_G1848_, new_G1849_, new_G1852_,
    new_G1853_, new_G1854_, new_G1857_, new_G1858_, new_G1859_, new_G1862_,
    new_G1863_, new_G1864_, new_G1867_, new_G1868_, new_G1869_, new_G1872_,
    new_G1873_, new_G1874_, new_G1877_, new_G1878_, new_G1879_, new_G1882_,
    new_G1883_, new_G1884_, new_G1887_, new_G1888_, new_G1889_, new_G1892_,
    new_G1895_, new_G1899_, new_G1902_, new_G1905_, new_G1908_, new_G1911_,
    new_G1914_, new_G1917_, new_G1920_, new_G1923_, new_G1926_, new_G1929_,
    new_G1932_, new_G1935_, new_G1938_, new_G1942_, new_G1943_, new_G1944_,
    new_G1948_, new_G1952_, new_G1956_, new_G1960_, new_G1964_, new_G1968_,
    new_G1972_, new_G1976_, new_G1980_, new_G1984_, new_G1988_, new_G1992_,
    new_G1996_, new_G1997_, new_G1998_, new_G2001_, new_G2002_, new_G2003_,
    new_G2004_, new_G2005_, new_G2006_, new_G2007_, new_G2008_, new_G2009_,
    new_G2010_, new_G2011_, new_G2012_, new_G2013_, new_G2014_, new_G2015_,
    new_G2016_, new_G2017_, new_G2018_, new_G2019_, new_G2020_, new_G2021_,
    new_G2022_, new_G2023_, new_G2024_, new_G2025_, new_G2026_, new_G2027_,
    new_G2030_, new_G2034_, new_G2037_, new_G2040_, new_G2043_, new_G2046_,
    new_G2049_, new_G2052_, new_G2055_, new_G2058_, new_G2061_, new_G2064_,
    new_G2067_, new_G2070_, new_G2073_, new_G2077_, new_G2078_, new_G2079_,
    new_G2082_, new_G2086_, new_G2090_, new_G2094_, new_G2098_, new_G2102_,
    new_G2106_, new_G2110_, new_G2114_, new_G2118_, new_G2122_, new_G2126_,
    new_G2130_, new_G2134_, new_G2135_, new_G2136_, new_G2139_, new_G2142_,
    new_G2146_, new_G2147_, new_G2148_, new_G2151_, new_G2152_, new_G2153_,
    new_G2156_, new_G2157_, new_G2158_, new_G2161_, new_G2162_, new_G2163_,
    new_G2166_, new_G2167_, new_G2168_, new_G2171_, new_G2172_, new_G2173_,
    new_G2176_, new_G2177_, new_G2178_, new_G2181_, new_G2182_, new_G2183_,
    new_G2186_, new_G2187_, new_G2188_, new_G2191_, new_G2192_, new_G2193_,
    new_G2196_, new_G2197_, new_G2198_, new_G2201_, new_G2202_, new_G2203_,
    new_G2206_, new_G2207_, new_G2208_, new_G2211_, new_G2214_, new_G2218_,
    new_G2219_, new_G2220_, new_G2223_, new_G2226_, new_G2229_, new_G2232_,
    new_G2235_, new_G2238_, new_G2241_, new_G2244_, new_G2247_, new_G2250_,
    new_G2253_, new_G2256_, new_G2260_, new_G2261_, new_G2262_, new_G2265_,
    new_G2269_, new_G2273_, new_G2277_, new_G2281_, new_G2285_, new_G2289_,
    new_G2293_, new_G2297_, new_G2301_, new_G2305_, new_G2309_, new_G2313_,
    new_G2314_, new_G2315_, new_G2318_, new_G2322_, new_G2323_, new_G2324_,
    new_G2325_, new_G2326_, new_G2327_, new_G2328_, new_G2329_, new_G2330_,
    new_G2331_, new_G2332_, new_G2333_, new_G2334_, new_G2335_, new_G2336_,
    new_G2337_, new_G2338_, new_G2339_, new_G2340_, new_G2341_, new_G2342_,
    new_G2343_, new_G2344_, new_G2345_, new_G2346_, new_G2349_, new_G2353_,
    new_G2354_, new_G2355_, new_G2358_, new_G2361_, new_G2364_, new_G2367_,
    new_G2370_, new_G2373_, new_G2376_, new_G2379_, new_G2382_, new_G2385_,
    new_G2388_, new_G2391_, new_G2394_, new_G2398_, new_G2399_, new_G2400_,
    new_G2403_, new_G2406_, new_G2410_, new_G2414_, new_G2418_, new_G2422_,
    new_G2426_, new_G2430_, new_G2434_, new_G2438_, new_G2442_, new_G2446_,
    new_G2450_, new_G2454_, new_G2458_, new_G2459_, new_G2460_, new_G2463_,
    new_G2466_, new_G2470_, new_G2471_, new_G2472_, new_G2473_, new_G2474_,
    new_G2477_, new_G2478_, new_G2479_, new_G2482_, new_G2483_, new_G2484_,
    new_G2487_, new_G2488_, new_G2489_, new_G2492_, new_G2493_, new_G2494_,
    new_G2497_, new_G2498_, new_G2499_, new_G2502_, new_G2503_, new_G2504_,
    new_G2507_, new_G2508_, new_G2509_, new_G2512_, new_G2513_, new_G2514_,
    new_G2517_, new_G2518_, new_G2519_, new_G2522_, new_G2523_, new_G2524_,
    new_G2527_, new_G2528_, new_G2529_, new_G2532_, new_G2535_, new_G2539_,
    new_G2540_, new_G2541_, new_G2544_, new_G2547_, new_G2550_, new_G2553_,
    new_G2556_, new_G2559_, new_G2562_, new_G2565_, new_G2568_, new_G2571_,
    new_G2574_, new_G2577_, new_G2581_, new_G2582_, new_G2583_, new_G2586_,
    new_G2590_, new_G2594_, new_G2598_, new_G2602_, new_G2606_, new_G2610_,
    new_G2614_, new_G2618_, new_G2622_, new_G2626_, new_G2630_, new_G2634_,
    new_G2635_, new_G2636_, new_G2639_, new_G2643_, new_G2644_, new_G2645_,
    new_G2648_, new_G2649_, new_G2650_, new_G2651_, new_G2652_, new_G2653_,
    new_G2654_, new_G2655_, new_G2656_, new_G2657_, new_G2658_, new_G2659_,
    new_G2660_, new_G2661_, new_G2662_, new_G2663_, new_G2664_, new_G2665_,
    new_G2666_, new_G2667_, new_G2668_, new_G2669_, new_G2670_, new_G2673_,
    new_G2677_, new_G2678_, new_G2679_, new_G2682_, new_G2685_, new_G2689_,
    new_G2692_, new_G2695_, new_G2698_, new_G2701_, new_G2704_, new_G2707_,
    new_G2710_, new_G2713_, new_G2716_, new_G2719_, new_G2722_, new_G2726_,
    new_G2727_, new_G2728_, new_G2731_, new_G2734_, new_G2738_, new_G2739_,
    new_G2740_, new_G2744_, new_G2748_, new_G2752_, new_G2756_, new_G2760_,
    new_G2764_, new_G2768_, new_G2772_, new_G2776_, new_G2780_, new_G2784_,
    new_G2785_, new_G2786_, new_G2789_, new_G2792_, new_G2796_, new_G2797_,
    new_G2798_, new_G2801_, new_G2802_, new_G2803_, new_G2806_, new_G2807_,
    new_G2808_, new_G2811_, new_G2812_, new_G2813_, new_G2816_, new_G2817_,
    new_G2818_, new_G2821_, new_G2822_, new_G2823_, new_G2826_, new_G2827_,
    new_G2828_, new_G2831_, new_G2832_, new_G2833_, new_G2836_, new_G2837_,
    new_G2838_, new_G2841_, new_G2842_, new_G2843_, new_G2846_, new_G2847_,
    new_G2848_, new_G2851_, new_G2852_, new_G2853_, new_G2856_, new_G2859_,
    new_G2863_, new_G2864_, new_G2865_, new_G2868_, new_G2872_, new_G2875_,
    new_G2878_, new_G2881_, new_G2884_, new_G2887_, new_G2890_, new_G2893_,
    new_G2896_, new_G2899_, new_G2902_, new_G2906_, new_G2907_, new_G2908_,
    new_G2911_, new_G2915_, new_G2916_, new_G2917_, new_G2920_, new_G2924_,
    new_G2928_, new_G2932_, new_G2936_, new_G2940_, new_G2944_, new_G2948_,
    new_G2952_, new_G2956_, new_G2960_, new_G2961_, new_G2962_, new_G2965_,
    new_G2969_, new_G2970_, new_G2971_, new_G2974_, new_G2977_, new_G2981_,
    new_G2982_, new_G2983_, new_G2984_, new_G2985_, new_G2986_, new_G2987_,
    new_G2988_, new_G2989_, new_G2990_, new_G2991_, new_G2992_, new_G2993_,
    new_G2994_, new_G2995_, new_G2996_, new_G2997_, new_G2998_, new_G2999_,
    new_G3000_, new_G3001_, new_G3004_, new_G3008_, new_G3009_, new_G3010_,
    new_G3013_, new_G3016_, new_G3020_, new_G3021_, new_G3022_, new_G3025_,
    new_G3028_, new_G3031_, new_G3034_, new_G3037_, new_G3040_, new_G3043_,
    new_G3046_, new_G3049_, new_G3052_, new_G3056_, new_G3057_, new_G3058_,
    new_G3061_, new_G3064_, new_G3068_, new_G3069_, new_G3070_, new_G3073_,
    new_G3077_, new_G3081_, new_G3085_, new_G3089_, new_G3093_, new_G3097_,
    new_G3101_, new_G3105_, new_G3109_, new_G3113_, new_G3114_, new_G3115_,
    new_G3118_, new_G3121_, new_G3125_, new_G3126_, new_G3127_, new_G3130_,
    new_G3134_, new_G3135_, new_G3136_, new_G3139_, new_G3140_, new_G3141_,
    new_G3144_, new_G3145_, new_G3146_, new_G3149_, new_G3150_, new_G3151_,
    new_G3154_, new_G3155_, new_G3156_, new_G3159_, new_G3160_, new_G3161_,
    new_G3164_, new_G3165_, new_G3166_, new_G3169_, new_G3170_, new_G3171_,
    new_G3174_, new_G3175_, new_G3176_, new_G3179_, new_G3180_, new_G3181_,
    new_G3184_, new_G3187_, new_G3191_, new_G3192_, new_G3193_, new_G3196_,
    new_G3200_, new_G3201_, new_G3202_, new_G3205_, new_G3208_, new_G3211_,
    new_G3214_, new_G3217_, new_G3220_, new_G3223_, new_G3226_, new_G3229_,
    new_G3232_, new_G3236_, new_G3237_, new_G3238_, new_G3241_, new_G3245_,
    new_G3246_, new_G3247_, new_G3250_, new_G3253_, new_G3257_, new_G3261_,
    new_G3265_, new_G3269_, new_G3273_, new_G3277_, new_G3281_, new_G3285_,
    new_G3289_, new_G3293_, new_G3294_, new_G3295_, new_G3298_, new_G3302_,
    new_G3303_, new_G3304_, new_G3307_, new_G3310_, new_G3314_, new_G3315_,
    new_G3316_, new_G3317_, new_G3318_, new_G3319_, new_G3320_, new_G3321_,
    new_G3322_, new_G3323_, new_G3324_, new_G3325_, new_G3326_, new_G3327_,
    new_G3328_, new_G3329_, new_G3330_, new_G3331_, new_G3332_, new_G3333_,
    new_G3334_, new_G3337_, new_G3341_, new_G3342_, new_G3343_, new_G3346_,
    new_G3349_, new_G3353_, new_G3354_, new_G3355_, new_G3358_, new_G3361_,
    new_G3364_, new_G3367_, new_G3370_, new_G3373_, new_G3376_, new_G3379_,
    new_G3382_, new_G3385_, new_G3389_, new_G3390_, new_G3391_, new_G3394_,
    new_G3397_, new_G3401_, new_G3402_, new_G3403_, new_G3406_, new_G3410_,
    new_G3414_, new_G3418_, new_G3422_, new_G3426_, new_G3430_, new_G3434_,
    new_G3438_, new_G3442_, new_G3446_, new_G3447_, new_G3448_, new_G3451_,
    new_G3454_, new_G3458_, new_G3459_, new_G3460_, new_G3463_, new_G3467_,
    new_G3468_, new_G3469_, new_G3472_, new_G3473_, new_G3474_, new_G3477_,
    new_G3478_, new_G3479_, new_G3482_, new_G3483_, new_G3484_, new_G3487_,
    new_G3488_, new_G3489_, new_G3492_, new_G3493_, new_G3494_, new_G3497_,
    new_G3498_, new_G3499_, new_G3502_, new_G3503_, new_G3504_, new_G3507_,
    new_G3508_, new_G3509_, new_G3512_, new_G3513_, new_G3514_, new_G3517_,
    new_G3520_, new_G3524_, new_G3525_, new_G3526_, new_G3529_, new_G3533_,
    new_G3534_, new_G3535_, new_G3538_, new_G3541_, new_G3545_, new_G3548_,
    new_G3551_, new_G3554_, new_G3557_, new_G3560_, new_G3563_, new_G3566_,
    new_G3569_, new_G3573_, new_G3574_, new_G3575_, new_G3578_, new_G3582_,
    new_G3583_, new_G3584_, new_G3587_, new_G3590_, new_G3594_, new_G3595_,
    new_G3596_, new_G3600_, new_G3604_, new_G3608_, new_G3612_, new_G3616_,
    new_G3620_, new_G3624_, new_G3628_, new_G3629_, new_G3630_, new_G3633_,
    new_G3637_, new_G3638_, new_G3639_, new_G3642_, new_G3645_, new_G3649_,
    new_G3650_, new_G3651_, new_G3654_, new_G3655_, new_G3656_, new_G3657_,
    new_G3658_, new_G3659_, new_G3660_, new_G3661_, new_G3662_, new_G3663_,
    new_G3664_, new_G3665_, new_G3666_, new_G3667_, new_G3668_, new_G3669_,
    new_G3670_, new_G3673_, new_G3677_, new_G3678_, new_G3679_, new_G3682_,
    new_G3685_, new_G3689_, new_G3690_, new_G3691_, new_G3694_, new_G3698_,
    new_G3701_, new_G3704_, new_G3707_, new_G3710_, new_G3713_, new_G3716_,
    new_G3719_, new_G3722_, new_G3726_, new_G3727_, new_G3728_, new_G3731_,
    new_G3734_, new_G3738_, new_G3739_, new_G3740_, new_G3743_, new_G3747_,
    new_G3748_, new_G3749_, new_G3752_, new_G3756_, new_G3760_, new_G3764_,
    new_G3768_, new_G3772_, new_G3776_, new_G3780_, new_G3784_, new_G3785_,
    new_G3786_, new_G3789_, new_G3792_, new_G3796_, new_G3797_, new_G3798_,
    new_G3801_, new_G3805_, new_G3806_, new_G3807_, new_G3810_, new_G3813_,
    new_G3817_, new_G3818_, new_G3819_, new_G3822_, new_G3823_, new_G3824_,
    new_G3827_, new_G3828_, new_G3829_, new_G3832_, new_G3833_, new_G3834_,
    new_G3837_, new_G3838_, new_G3839_, new_G3842_, new_G3843_, new_G3844_,
    new_G3847_, new_G3848_, new_G3849_, new_G3852_, new_G3853_, new_G3854_,
    new_G3857_, new_G3860_, new_G3864_, new_G3865_, new_G3866_, new_G3869_,
    new_G3873_, new_G3874_, new_G3875_, new_G3878_, new_G3881_, new_G3885_,
    new_G3886_, new_G3887_, new_G3890_, new_G3893_, new_G3896_, new_G3899_,
    new_G3902_, new_G3905_, new_G3908_, new_G3912_, new_G3913_, new_G3914_,
    new_G3917_, new_G3921_, new_G3922_, new_G3923_, new_G3926_, new_G3929_,
    new_G3933_, new_G3934_, new_G3935_, new_G3938_, new_G3942_, new_G3946_,
    new_G3950_, new_G3954_, new_G3958_, new_G3962_, new_G3966_, new_G3967_,
    new_G3968_, new_G3971_, new_G3975_, new_G3976_, new_G3977_, new_G3980_,
    new_G3983_, new_G3987_, new_G3988_, new_G3989_, new_G3992_, new_G3996_,
    new_G3997_, new_G3998_, new_G3999_, new_G4000_, new_G4001_, new_G4002_,
    new_G4003_, new_G4004_, new_G4005_, new_G4006_, new_G4007_, new_G4008_,
    new_G4009_, new_G4010_, new_G4013_, new_G4017_, new_G4018_, new_G4019_,
    new_G4022_, new_G4025_, new_G4029_, new_G4030_, new_G4031_, new_G4034_,
    new_G4038_, new_G4039_, new_G4040_, new_G4043_, new_G4046_, new_G4049_,
    new_G4052_, new_G4055_, new_G4058_, new_G4061_, new_G4064_, new_G4068_,
    new_G4069_, new_G4070_, new_G4073_, new_G4076_, new_G4080_, new_G4081_,
    new_G4082_, new_G4085_, new_G4089_, new_G4090_, new_G4091_, new_G4094_,
    new_G4097_, new_G4101_, new_G4105_, new_G4109_, new_G4113_, new_G4117_,
    new_G4121_, new_G4125_, new_G4129_, new_G4130_, new_G4131_, new_G4134_,
    new_G4137_, new_G4141_, new_G4142_, new_G4143_, new_G4146_, new_G4150_,
    new_G4151_, new_G4152_, new_G4155_, new_G4158_, new_G4162_, new_G4163_,
    new_G4164_, new_G4165_, new_G4166_, new_G4169_, new_G4170_, new_G4171_,
    new_G4174_, new_G4175_, new_G4176_, new_G4179_, new_G4180_, new_G4181_,
    new_G4184_, new_G4185_, new_G4186_, new_G4189_, new_G4190_, new_G4191_,
    new_G4194_, new_G4195_, new_G4196_, new_G4199_, new_G4202_, new_G4206_,
    new_G4207_, new_G4208_, new_G4211_, new_G4215_, new_G4216_, new_G4217_,
    new_G4220_, new_G4223_, new_G4227_, new_G4228_, new_G4229_, new_G4232_,
    new_G4235_, new_G4238_, new_G4241_, new_G4244_, new_G4247_, new_G4250_,
    new_G4254_, new_G4255_, new_G4256_, new_G4259_, new_G4263_, new_G4264_,
    new_G4265_, new_G4268_, new_G4271_, new_G4275_, new_G4276_, new_G4277_,
    new_G4280_, new_G4284_, new_G4288_, new_G4292_, new_G4296_, new_G4300_,
    new_G4304_, new_G4308_, new_G4309_, new_G4310_, new_G4313_, new_G4317_,
    new_G4318_, new_G4319_, new_G4322_, new_G4325_, new_G4329_, new_G4330_,
    new_G4331_, new_G4334_, new_G4338_, new_G4339_, new_G4340_, new_G4343_,
    new_G4344_, new_G4345_, new_G4346_, new_G4347_, new_G4348_, new_G4349_,
    new_G4350_, new_G4351_, new_G4352_, new_G4353_, new_G4354_, new_G4355_,
    new_G4358_, new_G4362_, new_G4363_, new_G4364_, new_G4367_, new_G4370_,
    new_G4374_, new_G4375_, new_G4376_, new_G4379_, new_G4383_, new_G4384_,
    new_G4385_, new_G4388_, new_G4391_, new_G4395_, new_G4398_, new_G4401_,
    new_G4404_, new_G4407_, new_G4410_, new_G4413_, new_G4417_, new_G4418_,
    new_G4419_, new_G4422_, new_G4425_, new_G4429_, new_G4430_, new_G4431_,
    new_G4434_, new_G4438_, new_G4439_, new_G4440_, new_G4443_, new_G4446_,
    new_G4450_, new_G4451_, new_G4452_, new_G4456_, new_G4460_, new_G4464_,
    new_G4468_, new_G4472_, new_G4476_, new_G4477_, new_G4478_, new_G4481_,
    new_G4484_, new_G4488_, new_G4489_, new_G4490_, new_G4493_, new_G4497_,
    new_G4498_, new_G4499_, new_G4502_, new_G4505_, new_G4509_, new_G4510_,
    new_G4511_, new_G4514_, new_G4515_, new_G4516_, new_G4519_, new_G4520_,
    new_G4521_, new_G4524_, new_G4525_, new_G4526_, new_G4529_, new_G4530_,
    new_G4531_, new_G4534_, new_G4535_, new_G4536_, new_G4539_, new_G4540_,
    new_G4541_, new_G4544_, new_G4547_, new_G4551_, new_G4552_, new_G4553_,
    new_G4556_, new_G4560_, new_G4561_, new_G4562_, new_G4565_, new_G4568_,
    new_G4572_, new_G4573_, new_G4574_, new_G4577_, new_G4581_, new_G4584_,
    new_G4587_, new_G4590_, new_G4593_, new_G4596_, new_G4600_, new_G4601_,
    new_G4602_, new_G4605_, new_G4609_, new_G4610_, new_G4611_, new_G4614_,
    new_G4617_, new_G4621_, new_G4622_, new_G4623_, new_G4626_, new_G4630_,
    new_G4631_, new_G4632_, new_G4635_, new_G4639_, new_G4643_, new_G4647_,
    new_G4651_, new_G4655_, new_G4656_, new_G4657_, new_G4660_, new_G4664_,
    new_G4665_, new_G4666_, new_G4669_, new_G4672_, new_G4676_, new_G4677_,
    new_G4678_, new_G4681_, new_G4685_, new_G4686_, new_G4687_, new_G4690_,
    new_G4693_, new_G4697_, new_G4698_, new_G4699_, new_G4700_, new_G4701_,
    new_G4702_, new_G4703_, new_G4704_, new_G4705_, new_G4706_, new_G4707_,
    new_G4710_, new_G4714_, new_G4715_, new_G4716_, new_G4719_, new_G4722_,
    new_G4726_, new_G4727_, new_G4728_, new_G4731_, new_G4735_, new_G4736_,
    new_G4737_, new_G4740_, new_G4743_, new_G4747_, new_G4748_, new_G4749_,
    new_G4752_, new_G4755_, new_G4758_, new_G4761_, new_G4764_, new_G4768_,
    new_G4769_, new_G4770_, new_G4773_, new_G4776_, new_G4780_, new_G4781_,
    new_G4782_, new_G4785_, new_G4789_, new_G4790_, new_G4791_, new_G4794_,
    new_G4797_, new_G4801_, new_G4802_, new_G4803_, new_G4806_, new_G4810_,
    new_G4814_, new_G4818_, new_G4822_, new_G4826_, new_G4827_, new_G4828_,
    new_G4831_, new_G4834_, new_G4838_, new_G4839_, new_G4840_, new_G4843_,
    new_G4847_, new_G4848_, new_G4849_, new_G4852_, new_G4855_, new_G4859_,
    new_G4860_, new_G4861_, new_G4864_, new_G4868_, new_G4869_, new_G4870_,
    new_G4873_, new_G4874_, new_G4875_, new_G4878_, new_G4879_, new_G4880_,
    new_G4883_, new_G4884_, new_G4885_, new_G4888_, new_G4889_, new_G4890_,
    new_G4893_, new_G4896_, new_G4900_, new_G4901_, new_G4902_, new_G4905_,
    new_G4909_, new_G4910_, new_G4911_, new_G4914_, new_G4917_, new_G4921_,
    new_G4922_, new_G4923_, new_G4926_, new_G4930_, new_G4931_, new_G4932_,
    new_G4935_, new_G4938_, new_G4941_, new_G4944_, new_G4947_, new_G4951_,
    new_G4952_, new_G4953_, new_G4956_, new_G4960_, new_G4961_, new_G4962_,
    new_G4965_, new_G4968_, new_G4972_, new_G4973_, new_G4974_, new_G4977_,
    new_G4981_, new_G4982_, new_G4983_, new_G4986_, new_G4989_, new_G4993_,
    new_G4997_, new_G5001_, new_G5005_, new_G5009_, new_G5010_, new_G5011_,
    new_G5014_, new_G5018_, new_G5019_, new_G5020_, new_G5023_, new_G5026_,
    new_G5030_, new_G5031_, new_G5032_, new_G5035_, new_G5039_, new_G5040_,
    new_G5041_, new_G5044_, new_G5047_, new_G5051_, new_G5052_, new_G5053_,
    new_G5054_, new_G5055_, new_G5056_, new_G5057_, new_G5058_, new_G5059_,
    new_G5060_, new_G5061_, new_G5064_, new_G5068_, new_G5069_, new_G5070_,
    new_G5073_, new_G5076_, new_G5080_, new_G5081_, new_G5082_, new_G5085_,
    new_G5089_, new_G5090_, new_G5091_, new_G5094_, new_G5097_, new_G5101_,
    new_G5102_, new_G5103_, new_G5106_, new_G5109_, new_G5112_, new_G5115_,
    new_G5118_, new_G5122_, new_G5123_, new_G5124_, new_G5127_, new_G5130_,
    new_G5134_, new_G5135_, new_G5136_, new_G5139_, new_G5143_, new_G5144_,
    new_G5145_, new_G5148_, new_G5151_, new_G5155_, new_G5156_, new_G5157_,
    new_G5160_, new_G5164_, new_G5168_, new_G5172_, new_G5176_, new_G5180_,
    new_G5181_, new_G5182_, new_G5185_, new_G5188_, new_G5192_, new_G5193_,
    new_G5194_, new_G5197_, new_G5201_, new_G5202_, new_G5203_, new_G5206_,
    new_G5209_, new_G5213_, new_G5214_, new_G5215_, new_G5218_, new_G5222_,
    new_G5223_, new_G5224_, new_G5227_, new_G5228_, new_G5229_, new_G5232_,
    new_G5233_, new_G5234_, new_G5237_, new_G5238_, new_G5239_, new_G5242_,
    new_G5243_, new_G5244_, new_G5247_, new_G5250_, new_G5254_, new_G5255_,
    new_G5256_, new_G5259_, new_G5263_, new_G5264_, new_G5265_, new_G5268_,
    new_G5271_, new_G5275_, new_G5276_, new_G5277_, new_G5280_, new_G5284_,
    new_G5285_, new_G5286_, new_G5289_, new_G5292_, new_G5296_, new_G5299_,
    new_G5302_, new_G5305_, new_G5309_, new_G5310_, new_G5311_, new_G5314_,
    new_G5318_, new_G5319_, new_G5320_, new_G5323_, new_G5326_, new_G5330_,
    new_G5331_, new_G5332_, new_G5335_, new_G5339_, new_G5340_, new_G5341_,
    new_G5344_, new_G5347_, new_G5351_, new_G5352_, new_G5353_, new_G5357_,
    new_G5361_, new_G5365_, new_G5366_, new_G5367_, new_G5370_, new_G5374_,
    new_G5375_, new_G5376_, new_G5379_, new_G5382_, new_G5386_, new_G5387_,
    new_G5388_, new_G5391_, new_G5395_, new_G5396_, new_G5397_, new_G5400_,
    new_G5403_, new_G5407_, new_G5408_, new_G5409_, new_G5412_, new_G5413_,
    new_G5414_, new_G5415_, new_G5416_, new_G5417_, new_G5418_, new_G5421_,
    new_G5425_, new_G5426_, new_G5427_, new_G5430_, new_G5433_, new_G5437_,
    new_G5438_, new_G5439_, new_G5442_, new_G5446_, new_G5447_, new_G5448_,
    new_G5451_, new_G5454_, new_G5458_, new_G5459_, new_G5460_, new_G5463_,
    new_G5467_, new_G5470_, new_G5473_, new_G5476_, new_G5480_, new_G5481_,
    new_G5482_, new_G5485_, new_G5488_, new_G5492_, new_G5493_, new_G5494_,
    new_G5497_, new_G5501_, new_G5502_, new_G5503_, new_G5506_, new_G5509_,
    new_G5513_, new_G5514_, new_G5515_, new_G5518_, new_G5522_, new_G5523_,
    new_G5524_, new_G5527_, new_G5531_, new_G5535_, new_G5539_, new_G5540_,
    new_G5541_, new_G5544_, new_G5547_, new_G5551_, new_G5552_, new_G5553_,
    new_G5556_, new_G5560_, new_G5561_, new_G5562_, new_G5565_, new_G5568_,
    new_G5572_, new_G5573_, new_G5574_, new_G5577_, new_G5581_, new_G5582_,
    new_G5583_, new_G5586_, new_G5589_, new_G5593_, new_G5594_, new_G5595_,
    new_G5598_, new_G5599_, new_G5600_, new_G5603_, new_G5604_, new_G5605_,
    new_G5608_, new_G5611_, new_G5615_, new_G5616_, new_G5617_, new_G5620_,
    new_G5624_, new_G5625_, new_G5626_, new_G5629_, new_G5632_, new_G5636_,
    new_G5637_, new_G5638_, new_G5641_, new_G5645_, new_G5646_, new_G5647_,
    new_G5650_, new_G5653_, new_G5657_, new_G5658_, new_G5659_, new_G5662_,
    new_G5665_, new_G5669_, new_G5670_, new_G5671_, new_G5674_, new_G5678_,
    new_G5679_, new_G5680_, new_G5683_, new_G5686_, new_G5690_, new_G5691_,
    new_G5692_, new_G5695_, new_G5699_, new_G5700_, new_G5701_, new_G5704_,
    new_G5707_, new_G5711_, new_G5712_, new_G5713_, new_G5716_, new_G5720_,
    new_G5724_, new_G5725_, new_G5726_, new_G5729_, new_G5733_, new_G5734_,
    new_G5735_, new_G5738_, new_G5741_, new_G5745_, new_G5746_, new_G5747_,
    new_G5750_, new_G5754_, new_G5755_, new_G5756_, new_G5759_, new_G5762_,
    new_G5766_, new_G5767_, new_G5768_, new_G5771_, new_G5772_, new_G5773_,
    new_G5774_, new_G5775_, new_G5778_, new_G5782_, new_G5783_, new_G5784_,
    new_G5787_, new_G5790_, new_G5794_, new_G5795_, new_G5796_, new_G5799_,
    new_G5803_, new_G5804_, new_G5805_, new_G5808_, new_G5811_, new_G5815_,
    new_G5816_, new_G5817_, new_G5820_, new_G5823_, new_G5826_, new_G5830_,
    new_G5831_, new_G5832_, new_G5835_, new_G5838_, new_G5842_, new_G5843_,
    new_G5844_, new_G5847_, new_G5851_, new_G5852_, new_G5853_, new_G5856_,
    new_G5859_, new_G5863_, new_G5864_, new_G5865_, new_G5868_, new_G5872_,
    new_G5876_, new_G5877_, new_G5878_, new_G5881_, new_G5884_, new_G5888_,
    new_G5889_, new_G5890_, new_G5893_, new_G5897_, new_G5898_, new_G5899_,
    new_G5902_, new_G5905_, new_G5909_, new_G5910_, new_G5911_, new_G5914_,
    new_G5915_, new_G5916_, new_G5919_, new_G5920_, new_G5921_, new_G5924_,
    new_G5927_, new_G5931_, new_G5932_, new_G5933_, new_G5936_, new_G5940_,
    new_G5941_, new_G5942_, new_G5945_, new_G5948_, new_G5952_, new_G5953_,
    new_G5954_, new_G5957_, new_G5960_, new_G5964_, new_G5965_, new_G5966_,
    new_G5969_, new_G5973_, new_G5974_, new_G5975_, new_G5978_, new_G5981_,
    new_G5985_, new_G5986_, new_G5987_, new_G5990_, new_G5994_, new_G5995_,
    new_G5996_, new_G5999_, new_G6003_, new_G6004_, new_G6005_, new_G6008_,
    new_G6011_, new_G6015_, new_G6016_, new_G6017_, new_G6020_, new_G6021_,
    new_G6022_, new_G6025_, new_G6029_, new_G6030_, new_G6031_, new_G6034_,
    new_G6037_, new_G6041_, new_G6042_, new_G6043_, new_G6046_, new_G6049_,
    new_G6053_, new_G6054_, new_G6055_, new_G6058_, new_G6061_, new_G6065_,
    new_G6066_, new_G6067_, new_G6070_, new_G6074_, new_G6075_, new_G6076_,
    new_G6079_, new_G6082_, new_G6086_, new_G6087_, new_G6088_, new_G6091_,
    new_G6092_, new_G6093_, new_G6096_, new_G6099_, new_G6103_, new_G6104_,
    new_G6105_, new_G6108_, new_G6112_, new_G6113_, new_G6114_, new_G6117_,
    new_G6118_, new_G6119_, new_G6122_, new_G6125_, new_G6129_, new_G6130_,
    new_G6131_, new_G6134_, new_G6138_, new_G6139_, new_G6140_, new_G6143_,
    new_G6147_, new_G6148_, new_G6149_, new_G6152_, new_G6156_, new_G6157_,
    new_G6158_, new_G6161_, new_G6165_, new_G6166_, new_G6167_, new_G6170_,
    new_G6174_, new_G6175_, new_G6176_, new_G6179_, new_G6183_, new_G6184_,
    new_G6185_, new_G6188_, new_G6192_, new_G6193_, new_G6194_, new_G6197_,
    new_G6201_, new_G6202_, new_G6203_, new_G6206_, new_G6210_, new_G6211_,
    new_G6212_, new_G6215_, new_G6219_, new_G6220_, new_G6221_, new_G6224_,
    new_G6228_, new_G6229_, new_G6230_, new_G6233_, new_G6237_, new_G6238_,
    new_G6239_, new_G6242_, new_G6246_, new_G6247_, new_G6248_, new_G6251_,
    new_G6255_, new_G6256_, n2482_li, n2485_li, n2488_li, n2491_li,
    n2494_li, n2497_li, n2500_li, n2503_li, n2506_li, n2509_li, n2512_li,
    n2515_li, n2518_li, n2521_li, n2524_li, n2527_li, n2530_li, n2533_li,
    n2536_li, n2539_li, n2542_li, n2545_li, n2548_li, n2551_li, n2554_li,
    n2557_li, n2560_li, n2563_li, n2566_li, n2569_li, n2572_li, n2575_li,
    n2578_li, n2581_li, n2584_li, n2587_li, n2590_li, n2593_li, n2596_li,
    n2599_li, n2602_li, n2605_li, n2608_li, n2611_li, n2614_li, n2617_li,
    n2620_li, n2623_li, n2626_li, n2629_li, n2632_li, n2635_li, n2638_li,
    n2641_li, n2644_li, n2647_li, n2650_li, n2653_li, n2656_li, n2659_li,
    n2662_li, n2665_li, n2668_li, n2671_li, n2674_li, n2677_li, n2680_li,
    n2683_li, n2686_li, n2689_li, n2692_li, n2695_li, n2698_li, n2701_li,
    n2704_li, n2707_li, n2710_li, n2713_li, n2716_li, n2719_li, n2722_li,
    n2725_li, n2728_li, n2731_li, n2734_li, n2737_li, n2740_li, n2743_li,
    n2746_li, n2749_li, n2752_li, n2755_li, n2758_li, n2761_li, n2764_li,
    n2767_li, n2770_li, n2773_li, n2776_li, n2779_li, n2782_li, n2785_li,
    n2788_li, n2791_li, n2794_li, n2797_li, n2800_li, n2803_li, n2806_li,
    n2809_li, n2812_li, n2815_li, n2818_li, n2821_li, n2824_li, n2827_li,
    n2830_li, n2833_li, n2836_li, n2839_li, n2842_li, n2845_li, n2848_li,
    n2851_li, n2854_li, n2857_li, n2860_li, n2863_li;
  assign new_G545_ = n2491_lo & n2695_lo;
  assign new_G548_ = n2491_lo & n2707_lo;
  assign new_G551_ = n2491_lo & n2719_lo;
  assign new_G554_ = n2491_lo & n2731_lo;
  assign new_G557_ = n2491_lo & n2743_lo;
  assign new_G560_ = n2491_lo & n2755_lo;
  assign new_G563_ = n2491_lo & n2767_lo;
  assign new_G566_ = n2491_lo & n2779_lo;
  assign new_G569_ = n2491_lo & n2791_lo;
  assign new_G572_ = n2491_lo & n2803_lo;
  assign new_G575_ = n2491_lo & n2815_lo;
  assign new_G578_ = n2491_lo & n2827_lo;
  assign new_G581_ = n2491_lo & n2839_lo;
  assign new_G584_ = n2491_lo & n2851_lo;
  assign new_G587_ = n2491_lo & n2863_lo;
  assign new_G590_ = n2503_lo & n2683_lo;
  assign new_G593_ = n2503_lo & n2695_lo;
  assign new_G596_ = n2503_lo & n2707_lo;
  assign new_G599_ = n2503_lo & n2719_lo;
  assign new_G602_ = n2503_lo & n2731_lo;
  assign new_G605_ = n2503_lo & n2743_lo;
  assign new_G608_ = n2503_lo & n2755_lo;
  assign new_G611_ = n2503_lo & n2767_lo;
  assign new_G614_ = n2503_lo & n2779_lo;
  assign new_G617_ = n2503_lo & n2791_lo;
  assign new_G620_ = n2503_lo & n2803_lo;
  assign new_G623_ = n2503_lo & n2815_lo;
  assign new_G626_ = n2503_lo & n2827_lo;
  assign new_G629_ = n2503_lo & n2839_lo;
  assign new_G632_ = n2503_lo & n2851_lo;
  assign new_G635_ = n2503_lo & n2863_lo;
  assign new_G638_ = n2515_lo & n2683_lo;
  assign new_G641_ = n2515_lo & n2695_lo;
  assign new_G644_ = n2515_lo & n2707_lo;
  assign new_G647_ = n2515_lo & n2719_lo;
  assign new_G650_ = n2515_lo & n2731_lo;
  assign new_G653_ = n2515_lo & n2743_lo;
  assign new_G656_ = n2515_lo & n2755_lo;
  assign new_G659_ = n2515_lo & n2767_lo;
  assign new_G662_ = n2515_lo & n2779_lo;
  assign new_G665_ = n2515_lo & n2791_lo;
  assign new_G668_ = n2515_lo & n2803_lo;
  assign new_G671_ = n2515_lo & n2815_lo;
  assign new_G674_ = n2515_lo & n2827_lo;
  assign new_G677_ = n2515_lo & n2839_lo;
  assign new_G680_ = n2515_lo & n2851_lo;
  assign new_G683_ = n2515_lo & n2863_lo;
  assign new_G686_ = n2527_lo & n2683_lo;
  assign new_G689_ = n2527_lo & n2695_lo;
  assign new_G692_ = n2527_lo & n2707_lo;
  assign new_G695_ = n2527_lo & n2719_lo;
  assign new_G698_ = n2527_lo & n2731_lo;
  assign new_G701_ = n2527_lo & n2743_lo;
  assign new_G704_ = n2527_lo & n2755_lo;
  assign new_G707_ = n2527_lo & n2767_lo;
  assign new_G710_ = n2527_lo & n2779_lo;
  assign new_G713_ = n2527_lo & n2791_lo;
  assign new_G716_ = n2527_lo & n2803_lo;
  assign new_G719_ = n2527_lo & n2815_lo;
  assign new_G722_ = n2527_lo & n2827_lo;
  assign new_G725_ = n2527_lo & n2839_lo;
  assign new_G728_ = n2527_lo & n2851_lo;
  assign new_G731_ = n2527_lo & n2863_lo;
  assign new_G734_ = n2539_lo & n2683_lo;
  assign new_G737_ = n2539_lo & n2695_lo;
  assign new_G740_ = n2539_lo & n2707_lo;
  assign new_G743_ = n2539_lo & n2719_lo;
  assign new_G746_ = n2539_lo & n2731_lo;
  assign new_G749_ = n2539_lo & n2743_lo;
  assign new_G752_ = n2539_lo & n2755_lo;
  assign new_G755_ = n2539_lo & n2767_lo;
  assign new_G758_ = n2539_lo & n2779_lo;
  assign new_G761_ = n2539_lo & n2791_lo;
  assign new_G764_ = n2539_lo & n2803_lo;
  assign new_G767_ = n2539_lo & n2815_lo;
  assign new_G770_ = n2539_lo & n2827_lo;
  assign new_G773_ = n2539_lo & n2839_lo;
  assign new_G776_ = n2539_lo & n2851_lo;
  assign new_G779_ = n2539_lo & n2863_lo;
  assign new_G782_ = n2551_lo & n2683_lo;
  assign new_G785_ = n2551_lo & n2695_lo;
  assign new_G788_ = n2551_lo & n2707_lo;
  assign new_G791_ = n2551_lo & n2719_lo;
  assign new_G794_ = n2551_lo & n2731_lo;
  assign new_G797_ = n2551_lo & n2743_lo;
  assign new_G800_ = n2551_lo & n2755_lo;
  assign new_G803_ = n2551_lo & n2767_lo;
  assign new_G806_ = n2551_lo & n2779_lo;
  assign new_G809_ = n2551_lo & n2791_lo;
  assign new_G812_ = n2551_lo & n2803_lo;
  assign new_G815_ = n2551_lo & n2815_lo;
  assign new_G818_ = n2551_lo & n2827_lo;
  assign new_G821_ = n2551_lo & n2839_lo;
  assign new_G824_ = n2551_lo & n2851_lo;
  assign new_G827_ = n2551_lo & n2863_lo;
  assign new_G830_ = n2563_lo & n2683_lo;
  assign new_G833_ = n2563_lo & n2695_lo;
  assign new_G836_ = n2563_lo & n2707_lo;
  assign new_G839_ = n2563_lo & n2719_lo;
  assign new_G842_ = n2563_lo & n2731_lo;
  assign new_G845_ = n2563_lo & n2743_lo;
  assign new_G848_ = n2563_lo & n2755_lo;
  assign new_G851_ = n2563_lo & n2767_lo;
  assign new_G854_ = n2563_lo & n2779_lo;
  assign new_G857_ = n2563_lo & n2791_lo;
  assign new_G860_ = n2563_lo & n2803_lo;
  assign new_G863_ = n2563_lo & n2815_lo;
  assign new_G866_ = n2563_lo & n2827_lo;
  assign new_G869_ = n2563_lo & n2839_lo;
  assign new_G872_ = n2563_lo & n2851_lo;
  assign new_G875_ = n2563_lo & n2863_lo;
  assign new_G878_ = n2575_lo & n2683_lo;
  assign new_G881_ = n2575_lo & n2695_lo;
  assign new_G884_ = n2575_lo & n2707_lo;
  assign new_G887_ = n2575_lo & n2719_lo;
  assign new_G890_ = n2575_lo & n2731_lo;
  assign new_G893_ = n2575_lo & n2743_lo;
  assign new_G896_ = n2575_lo & n2755_lo;
  assign new_G899_ = n2575_lo & n2767_lo;
  assign new_G902_ = n2575_lo & n2779_lo;
  assign new_G905_ = n2575_lo & n2791_lo;
  assign new_G908_ = n2575_lo & n2803_lo;
  assign new_G911_ = n2575_lo & n2815_lo;
  assign new_G914_ = n2575_lo & n2827_lo;
  assign new_G917_ = n2575_lo & n2839_lo;
  assign new_G920_ = n2575_lo & n2851_lo;
  assign new_G923_ = n2575_lo & n2863_lo;
  assign new_G926_ = n2587_lo & n2683_lo;
  assign new_G929_ = n2587_lo & n2695_lo;
  assign new_G932_ = n2587_lo & n2707_lo;
  assign new_G935_ = n2587_lo & n2719_lo;
  assign new_G938_ = n2587_lo & n2731_lo;
  assign new_G941_ = n2587_lo & n2743_lo;
  assign new_G944_ = n2587_lo & n2755_lo;
  assign new_G947_ = n2587_lo & n2767_lo;
  assign new_G950_ = n2587_lo & n2779_lo;
  assign new_G953_ = n2587_lo & n2791_lo;
  assign new_G956_ = n2587_lo & n2803_lo;
  assign new_G959_ = n2587_lo & n2815_lo;
  assign new_G962_ = n2587_lo & n2827_lo;
  assign new_G965_ = n2587_lo & n2839_lo;
  assign new_G968_ = n2587_lo & n2851_lo;
  assign new_G971_ = n2587_lo & n2863_lo;
  assign new_G974_ = n2599_lo & n2683_lo;
  assign new_G977_ = n2599_lo & n2695_lo;
  assign new_G980_ = n2599_lo & n2707_lo;
  assign new_G983_ = n2599_lo & n2719_lo;
  assign new_G986_ = n2599_lo & n2731_lo;
  assign new_G989_ = n2599_lo & n2743_lo;
  assign new_G992_ = n2599_lo & n2755_lo;
  assign new_G995_ = n2599_lo & n2767_lo;
  assign new_G998_ = n2599_lo & n2779_lo;
  assign new_G1001_ = n2599_lo & n2791_lo;
  assign new_G1004_ = n2599_lo & n2803_lo;
  assign new_G1007_ = n2599_lo & n2815_lo;
  assign new_G1010_ = n2599_lo & n2827_lo;
  assign new_G1013_ = n2599_lo & n2839_lo;
  assign new_G1016_ = n2599_lo & n2851_lo;
  assign new_G1019_ = n2599_lo & n2863_lo;
  assign new_G1022_ = n2611_lo & n2683_lo;
  assign new_G1025_ = n2611_lo & n2695_lo;
  assign new_G1028_ = n2611_lo & n2707_lo;
  assign new_G1031_ = n2611_lo & n2719_lo;
  assign new_G1034_ = n2611_lo & n2731_lo;
  assign new_G1037_ = n2611_lo & n2743_lo;
  assign new_G1040_ = n2611_lo & n2755_lo;
  assign new_G1043_ = n2611_lo & n2767_lo;
  assign new_G1046_ = n2611_lo & n2779_lo;
  assign new_G1049_ = n2611_lo & n2791_lo;
  assign new_G1052_ = n2611_lo & n2803_lo;
  assign new_G1055_ = n2611_lo & n2815_lo;
  assign new_G1058_ = n2611_lo & n2827_lo;
  assign new_G1061_ = n2611_lo & n2839_lo;
  assign new_G1064_ = n2611_lo & n2851_lo;
  assign new_G1067_ = n2611_lo & n2863_lo;
  assign new_G1070_ = n2623_lo & n2683_lo;
  assign new_G1073_ = n2623_lo & n2695_lo;
  assign new_G1076_ = n2623_lo & n2707_lo;
  assign new_G1079_ = n2623_lo & n2719_lo;
  assign new_G1082_ = n2623_lo & n2731_lo;
  assign new_G1085_ = n2623_lo & n2743_lo;
  assign new_G1088_ = n2623_lo & n2755_lo;
  assign new_G1091_ = n2623_lo & n2767_lo;
  assign new_G1094_ = n2623_lo & n2779_lo;
  assign new_G1097_ = n2623_lo & n2791_lo;
  assign new_G1100_ = n2623_lo & n2803_lo;
  assign new_G1103_ = n2623_lo & n2815_lo;
  assign new_G1106_ = n2623_lo & n2827_lo;
  assign new_G1109_ = n2623_lo & n2839_lo;
  assign new_G1112_ = n2623_lo & n2851_lo;
  assign new_G1115_ = n2623_lo & n2863_lo;
  assign new_G1118_ = n2635_lo & n2683_lo;
  assign new_G1121_ = n2635_lo & n2695_lo;
  assign new_G1124_ = n2635_lo & n2707_lo;
  assign new_G1127_ = n2635_lo & n2719_lo;
  assign new_G1130_ = n2635_lo & n2731_lo;
  assign new_G1133_ = n2635_lo & n2743_lo;
  assign new_G1136_ = n2635_lo & n2755_lo;
  assign new_G1139_ = n2635_lo & n2767_lo;
  assign new_G1142_ = n2635_lo & n2779_lo;
  assign new_G1145_ = n2635_lo & n2791_lo;
  assign new_G1148_ = n2635_lo & n2803_lo;
  assign new_G1151_ = n2635_lo & n2815_lo;
  assign new_G1154_ = n2635_lo & n2827_lo;
  assign new_G1157_ = n2635_lo & n2839_lo;
  assign new_G1160_ = n2635_lo & n2851_lo;
  assign new_G1163_ = n2635_lo & n2863_lo;
  assign new_G1166_ = n2647_lo & n2683_lo;
  assign new_G1169_ = n2647_lo & n2695_lo;
  assign new_G1172_ = n2647_lo & n2707_lo;
  assign new_G1175_ = n2647_lo & n2719_lo;
  assign new_G1178_ = n2647_lo & n2731_lo;
  assign new_G1181_ = n2647_lo & n2743_lo;
  assign new_G1184_ = n2647_lo & n2755_lo;
  assign new_G1187_ = n2647_lo & n2767_lo;
  assign new_G1190_ = n2647_lo & n2779_lo;
  assign new_G1193_ = n2647_lo & n2791_lo;
  assign new_G1196_ = n2647_lo & n2803_lo;
  assign new_G1199_ = n2647_lo & n2815_lo;
  assign new_G1202_ = n2647_lo & n2827_lo;
  assign new_G1205_ = n2647_lo & n2839_lo;
  assign new_G1208_ = n2647_lo & n2851_lo;
  assign new_G1211_ = n2647_lo & n2863_lo;
  assign new_G1214_ = n2659_lo & n2683_lo;
  assign new_G1217_ = n2659_lo & n2695_lo;
  assign new_G1220_ = n2659_lo & n2707_lo;
  assign new_G1223_ = n2659_lo & n2719_lo;
  assign new_G1226_ = n2659_lo & n2731_lo;
  assign new_G1229_ = n2659_lo & n2743_lo;
  assign new_G1232_ = n2659_lo & n2755_lo;
  assign new_G1235_ = n2659_lo & n2767_lo;
  assign new_G1238_ = n2659_lo & n2779_lo;
  assign new_G1241_ = n2659_lo & n2791_lo;
  assign new_G1244_ = n2659_lo & n2803_lo;
  assign new_G1247_ = n2659_lo & n2815_lo;
  assign new_G1250_ = n2659_lo & n2827_lo;
  assign new_G1253_ = n2659_lo & n2839_lo;
  assign new_G1256_ = n2659_lo & n2851_lo;
  assign new_G1259_ = n2659_lo & n2863_lo;
  assign new_G1262_ = n2671_lo & n2683_lo;
  assign new_G1265_ = n2671_lo & n2695_lo;
  assign new_G1268_ = n2671_lo & n2707_lo;
  assign new_G1271_ = n2671_lo & n2719_lo;
  assign new_G1274_ = n2671_lo & n2731_lo;
  assign new_G1277_ = n2671_lo & n2743_lo;
  assign new_G1280_ = n2671_lo & n2755_lo;
  assign new_G1283_ = n2671_lo & n2767_lo;
  assign new_G1286_ = n2671_lo & n2779_lo;
  assign new_G1289_ = n2671_lo & n2791_lo;
  assign new_G1292_ = n2671_lo & n2803_lo;
  assign new_G1295_ = n2671_lo & n2815_lo;
  assign new_G1298_ = n2671_lo & n2827_lo;
  assign new_G1301_ = n2671_lo & n2839_lo;
  assign new_G1304_ = n2671_lo & n2851_lo;
  assign new_G1307_ = n2671_lo & n2863_lo;
  assign new_G1310_ = ~new_G590_;
  assign new_G1314_ = ~new_G638_;
  assign new_G1318_ = ~new_G686_;
  assign new_G1322_ = ~new_G734_;
  assign new_G1326_ = ~new_G782_;
  assign new_G1330_ = ~new_G830_;
  assign new_G1334_ = ~new_G878_;
  assign new_G1338_ = ~new_G926_;
  assign new_G1342_ = ~new_G974_;
  assign new_G1346_ = ~new_G1022_;
  assign new_G1350_ = ~new_G1070_;
  assign new_G1354_ = ~new_G1118_;
  assign new_G1358_ = ~new_G1166_;
  assign new_G1362_ = ~new_G1214_;
  assign new_G1366_ = ~new_G1262_;
  assign new_G1370_ = ~new_G590_ & ~new_G1310_;
  assign new_G1371_ = ~new_G1310_;
  assign new_G1372_ = ~new_G638_ & ~new_G1314_;
  assign new_G1373_ = ~new_G1314_;
  assign new_G1374_ = ~new_G686_ & ~new_G1318_;
  assign new_G1375_ = ~new_G1318_;
  assign new_G1376_ = ~new_G734_ & ~new_G1322_;
  assign new_G1377_ = ~new_G1322_;
  assign new_G1378_ = ~new_G782_ & ~new_G1326_;
  assign new_G1379_ = ~new_G1326_;
  assign new_G1380_ = ~new_G830_ & ~new_G1330_;
  assign new_G1381_ = ~new_G1330_;
  assign new_G1382_ = ~new_G878_ & ~new_G1334_;
  assign new_G1383_ = ~new_G1334_;
  assign new_G1384_ = ~new_G926_ & ~new_G1338_;
  assign new_G1385_ = ~new_G1338_;
  assign new_G1386_ = ~new_G974_ & ~new_G1342_;
  assign new_G1387_ = ~new_G1342_;
  assign new_G1388_ = ~new_G1022_ & ~new_G1346_;
  assign new_G1389_ = ~new_G1346_;
  assign new_G1390_ = ~new_G1070_ & ~new_G1350_;
  assign new_G1391_ = ~new_G1350_;
  assign new_G1392_ = ~new_G1118_ & ~new_G1354_;
  assign new_G1393_ = ~new_G1354_;
  assign new_G1394_ = ~new_G1166_ & ~new_G1358_;
  assign new_G1395_ = ~new_G1358_;
  assign new_G1396_ = ~new_G1214_ & ~new_G1362_;
  assign new_G1397_ = ~new_G1362_;
  assign new_G1398_ = ~new_G1262_ & ~new_G1366_;
  assign new_G1399_ = ~new_G1366_;
  assign new_G1400_ = ~new_G1370_ & ~new_G1371_;
  assign new_G1403_ = ~new_G1372_ & ~new_G1373_;
  assign new_G1406_ = ~new_G1374_ & ~new_G1375_;
  assign new_G1409_ = ~new_G1376_ & ~new_G1377_;
  assign new_G1412_ = ~new_G1378_ & ~new_G1379_;
  assign new_G1415_ = ~new_G1380_ & ~new_G1381_;
  assign new_G1418_ = ~new_G1382_ & ~new_G1383_;
  assign new_G1421_ = ~new_G1384_ & ~new_G1385_;
  assign new_G1424_ = ~new_G1386_ & ~new_G1387_;
  assign new_G1427_ = ~new_G1388_ & ~new_G1389_;
  assign new_G1430_ = ~new_G1390_ & ~new_G1391_;
  assign new_G1433_ = ~new_G1392_ & ~new_G1393_;
  assign new_G1436_ = ~new_G1394_ & ~new_G1395_;
  assign new_G1439_ = ~new_G1396_ & ~new_G1397_;
  assign new_G1442_ = ~new_G1398_ & ~new_G1399_;
  assign new_G1445_ = ~new_G1400_ & ~new_G545_;
  assign new_G1449_ = ~new_G1403_ & ~new_G593_;
  assign new_G1453_ = ~new_G1406_ & ~new_G641_;
  assign new_G1457_ = ~new_G1409_ & ~new_G689_;
  assign new_G1461_ = ~new_G1412_ & ~new_G737_;
  assign new_G1465_ = ~new_G1415_ & ~new_G785_;
  assign new_G1469_ = ~new_G1418_ & ~new_G833_;
  assign new_G1473_ = ~new_G1421_ & ~new_G881_;
  assign new_G1477_ = ~new_G1424_ & ~new_G929_;
  assign new_G1481_ = ~new_G1427_ & ~new_G977_;
  assign new_G1485_ = ~new_G1430_ & ~new_G1025_;
  assign new_G1489_ = ~new_G1433_ & ~new_G1073_;
  assign new_G1493_ = ~new_G1436_ & ~new_G1121_;
  assign new_G1497_ = ~new_G1439_ & ~new_G1169_;
  assign new_G1501_ = ~new_G1442_ & ~new_G1217_;
  assign new_G1505_ = ~new_G1400_ & ~new_G1445_;
  assign new_G1506_ = ~new_G1445_ & ~new_G545_;
  assign new_G1507_ = ~new_G1310_ & ~new_G1445_;
  assign new_G1510_ = ~new_G1403_ & ~new_G1449_;
  assign new_G1511_ = ~new_G1449_ & ~new_G593_;
  assign new_G1512_ = ~new_G1314_ & ~new_G1449_;
  assign new_G1515_ = ~new_G1406_ & ~new_G1453_;
  assign new_G1516_ = ~new_G1453_ & ~new_G641_;
  assign new_G1517_ = ~new_G1318_ & ~new_G1453_;
  assign new_G1520_ = ~new_G1409_ & ~new_G1457_;
  assign new_G1521_ = ~new_G1457_ & ~new_G689_;
  assign new_G1522_ = ~new_G1322_ & ~new_G1457_;
  assign new_G1525_ = ~new_G1412_ & ~new_G1461_;
  assign new_G1526_ = ~new_G1461_ & ~new_G737_;
  assign new_G1527_ = ~new_G1326_ & ~new_G1461_;
  assign new_G1530_ = ~new_G1415_ & ~new_G1465_;
  assign new_G1531_ = ~new_G1465_ & ~new_G785_;
  assign new_G1532_ = ~new_G1330_ & ~new_G1465_;
  assign new_G1535_ = ~new_G1418_ & ~new_G1469_;
  assign new_G1536_ = ~new_G1469_ & ~new_G833_;
  assign new_G1537_ = ~new_G1334_ & ~new_G1469_;
  assign new_G1540_ = ~new_G1421_ & ~new_G1473_;
  assign new_G1541_ = ~new_G1473_ & ~new_G881_;
  assign new_G1542_ = ~new_G1338_ & ~new_G1473_;
  assign new_G1545_ = ~new_G1424_ & ~new_G1477_;
  assign new_G1546_ = ~new_G1477_ & ~new_G929_;
  assign new_G1547_ = ~new_G1342_ & ~new_G1477_;
  assign new_G1550_ = ~new_G1427_ & ~new_G1481_;
  assign new_G1551_ = ~new_G1481_ & ~new_G977_;
  assign new_G1552_ = ~new_G1346_ & ~new_G1481_;
  assign new_G1555_ = ~new_G1430_ & ~new_G1485_;
  assign new_G1556_ = ~new_G1485_ & ~new_G1025_;
  assign new_G1557_ = ~new_G1350_ & ~new_G1485_;
  assign new_G1560_ = ~new_G1433_ & ~new_G1489_;
  assign new_G1561_ = ~new_G1489_ & ~new_G1073_;
  assign new_G1562_ = ~new_G1354_ & ~new_G1489_;
  assign new_G1565_ = ~new_G1436_ & ~new_G1493_;
  assign new_G1566_ = ~new_G1493_ & ~new_G1121_;
  assign new_G1567_ = ~new_G1358_ & ~new_G1493_;
  assign new_G1570_ = ~new_G1439_ & ~new_G1497_;
  assign new_G1571_ = ~new_G1497_ & ~new_G1169_;
  assign new_G1572_ = ~new_G1362_ & ~new_G1497_;
  assign new_G1575_ = ~new_G1442_ & ~new_G1501_;
  assign new_G1576_ = ~new_G1501_ & ~new_G1217_;
  assign new_G1577_ = ~new_G1366_ & ~new_G1501_;
  assign new_G1580_ = ~new_G1510_ & ~new_G1511_;
  assign new_G1583_ = ~new_G1515_ & ~new_G1516_;
  assign new_G1586_ = ~new_G1520_ & ~new_G1521_;
  assign new_G1589_ = ~new_G1525_ & ~new_G1526_;
  assign new_G1592_ = ~new_G1530_ & ~new_G1531_;
  assign new_G1595_ = ~new_G1535_ & ~new_G1536_;
  assign new_G1598_ = ~new_G1540_ & ~new_G1541_;
  assign new_G1601_ = ~new_G1545_ & ~new_G1546_;
  assign new_G1604_ = ~new_G1550_ & ~new_G1551_;
  assign new_G1607_ = ~new_G1555_ & ~new_G1556_;
  assign new_G1610_ = ~new_G1560_ & ~new_G1561_;
  assign new_G1613_ = ~new_G1565_ & ~new_G1566_;
  assign new_G1616_ = ~new_G1570_ & ~new_G1571_;
  assign new_G1619_ = ~new_G1575_ & ~new_G1576_;
  assign new_G1622_ = ~new_G1265_ & ~new_G1577_;
  assign new_G1626_ = ~new_G1580_ & ~new_G1507_;
  assign new_G1630_ = ~new_G1583_ & ~new_G1512_;
  assign new_G1634_ = ~new_G1586_ & ~new_G1517_;
  assign new_G1638_ = ~new_G1589_ & ~new_G1522_;
  assign new_G1642_ = ~new_G1592_ & ~new_G1527_;
  assign new_G1646_ = ~new_G1595_ & ~new_G1532_;
  assign new_G1650_ = ~new_G1598_ & ~new_G1537_;
  assign new_G1654_ = ~new_G1601_ & ~new_G1542_;
  assign new_G1658_ = ~new_G1604_ & ~new_G1547_;
  assign new_G1662_ = ~new_G1607_ & ~new_G1552_;
  assign new_G1666_ = ~new_G1610_ & ~new_G1557_;
  assign new_G1670_ = ~new_G1613_ & ~new_G1562_;
  assign new_G1674_ = ~new_G1616_ & ~new_G1567_;
  assign new_G1678_ = ~new_G1619_ & ~new_G1572_;
  assign new_G1682_ = ~new_G1265_ & ~new_G1622_;
  assign new_G1683_ = ~new_G1622_ & ~new_G1577_;
  assign new_G1684_ = ~new_G1580_ & ~new_G1626_;
  assign new_G1685_ = ~new_G1626_ & ~new_G1507_;
  assign new_G1686_ = ~new_G1583_ & ~new_G1630_;
  assign new_G1687_ = ~new_G1630_ & ~new_G1512_;
  assign new_G1688_ = ~new_G1586_ & ~new_G1634_;
  assign new_G1689_ = ~new_G1634_ & ~new_G1517_;
  assign new_G1690_ = ~new_G1589_ & ~new_G1638_;
  assign new_G1691_ = ~new_G1638_ & ~new_G1522_;
  assign new_G1692_ = ~new_G1592_ & ~new_G1642_;
  assign new_G1693_ = ~new_G1642_ & ~new_G1527_;
  assign new_G1694_ = ~new_G1595_ & ~new_G1646_;
  assign new_G1695_ = ~new_G1646_ & ~new_G1532_;
  assign new_G1696_ = ~new_G1598_ & ~new_G1650_;
  assign new_G1697_ = ~new_G1650_ & ~new_G1537_;
  assign new_G1698_ = ~new_G1601_ & ~new_G1654_;
  assign new_G1699_ = ~new_G1654_ & ~new_G1542_;
  assign new_G1700_ = ~new_G1604_ & ~new_G1658_;
  assign new_G1701_ = ~new_G1658_ & ~new_G1547_;
  assign new_G1702_ = ~new_G1607_ & ~new_G1662_;
  assign new_G1703_ = ~new_G1662_ & ~new_G1552_;
  assign new_G1704_ = ~new_G1610_ & ~new_G1666_;
  assign new_G1705_ = ~new_G1666_ & ~new_G1557_;
  assign new_G1706_ = ~new_G1613_ & ~new_G1670_;
  assign new_G1707_ = ~new_G1670_ & ~new_G1562_;
  assign new_G1708_ = ~new_G1616_ & ~new_G1674_;
  assign new_G1709_ = ~new_G1674_ & ~new_G1567_;
  assign new_G1710_ = ~new_G1619_ & ~new_G1678_;
  assign new_G1711_ = ~new_G1678_ & ~new_G1572_;
  assign new_G1712_ = ~new_G1682_ & ~new_G1683_;
  assign new_G1715_ = ~new_G1684_ & ~new_G1685_;
  assign new_G1718_ = ~new_G1686_ & ~new_G1687_;
  assign new_G1721_ = ~new_G1688_ & ~new_G1689_;
  assign new_G1724_ = ~new_G1690_ & ~new_G1691_;
  assign new_G1727_ = ~new_G1692_ & ~new_G1693_;
  assign new_G1730_ = ~new_G1694_ & ~new_G1695_;
  assign new_G1733_ = ~new_G1696_ & ~new_G1697_;
  assign new_G1736_ = ~new_G1698_ & ~new_G1699_;
  assign new_G1739_ = ~new_G1700_ & ~new_G1701_;
  assign new_G1742_ = ~new_G1702_ & ~new_G1703_;
  assign new_G1745_ = ~new_G1704_ & ~new_G1705_;
  assign new_G1748_ = ~new_G1706_ & ~new_G1707_;
  assign new_G1751_ = ~new_G1708_ & ~new_G1709_;
  assign new_G1754_ = ~new_G1710_ & ~new_G1711_;
  assign new_G1757_ = ~new_G1712_ & ~new_G1220_;
  assign new_G1761_ = ~new_G1715_ & ~new_G548_;
  assign new_G1765_ = ~new_G1718_ & ~new_G596_;
  assign new_G1769_ = ~new_G1721_ & ~new_G644_;
  assign new_G1773_ = ~new_G1724_ & ~new_G692_;
  assign new_G1777_ = ~new_G1727_ & ~new_G740_;
  assign new_G1781_ = ~new_G1730_ & ~new_G788_;
  assign new_G1785_ = ~new_G1733_ & ~new_G836_;
  assign new_G1789_ = ~new_G1736_ & ~new_G884_;
  assign new_G1793_ = ~new_G1739_ & ~new_G932_;
  assign new_G1797_ = ~new_G1742_ & ~new_G980_;
  assign new_G1801_ = ~new_G1745_ & ~new_G1028_;
  assign new_G1805_ = ~new_G1748_ & ~new_G1076_;
  assign new_G1809_ = ~new_G1751_ & ~new_G1124_;
  assign new_G1813_ = ~new_G1754_ & ~new_G1172_;
  assign new_G1817_ = ~new_G1712_ & ~new_G1757_;
  assign new_G1818_ = ~new_G1757_ & ~new_G1220_;
  assign new_G1819_ = ~new_G1622_ & ~new_G1757_;
  assign new_G1822_ = ~new_G1715_ & ~new_G1761_;
  assign new_G1823_ = ~new_G1761_ & ~new_G548_;
  assign new_G1824_ = ~new_G1626_ & ~new_G1761_;
  assign new_G1827_ = ~new_G1718_ & ~new_G1765_;
  assign new_G1828_ = ~new_G1765_ & ~new_G596_;
  assign new_G1829_ = ~new_G1630_ & ~new_G1765_;
  assign new_G1832_ = ~new_G1721_ & ~new_G1769_;
  assign new_G1833_ = ~new_G1769_ & ~new_G644_;
  assign new_G1834_ = ~new_G1634_ & ~new_G1769_;
  assign new_G1837_ = ~new_G1724_ & ~new_G1773_;
  assign new_G1838_ = ~new_G1773_ & ~new_G692_;
  assign new_G1839_ = ~new_G1638_ & ~new_G1773_;
  assign new_G1842_ = ~new_G1727_ & ~new_G1777_;
  assign new_G1843_ = ~new_G1777_ & ~new_G740_;
  assign new_G1844_ = ~new_G1642_ & ~new_G1777_;
  assign new_G1847_ = ~new_G1730_ & ~new_G1781_;
  assign new_G1848_ = ~new_G1781_ & ~new_G788_;
  assign new_G1849_ = ~new_G1646_ & ~new_G1781_;
  assign new_G1852_ = ~new_G1733_ & ~new_G1785_;
  assign new_G1853_ = ~new_G1785_ & ~new_G836_;
  assign new_G1854_ = ~new_G1650_ & ~new_G1785_;
  assign new_G1857_ = ~new_G1736_ & ~new_G1789_;
  assign new_G1858_ = ~new_G1789_ & ~new_G884_;
  assign new_G1859_ = ~new_G1654_ & ~new_G1789_;
  assign new_G1862_ = ~new_G1739_ & ~new_G1793_;
  assign new_G1863_ = ~new_G1793_ & ~new_G932_;
  assign new_G1864_ = ~new_G1658_ & ~new_G1793_;
  assign new_G1867_ = ~new_G1742_ & ~new_G1797_;
  assign new_G1868_ = ~new_G1797_ & ~new_G980_;
  assign new_G1869_ = ~new_G1662_ & ~new_G1797_;
  assign new_G1872_ = ~new_G1745_ & ~new_G1801_;
  assign new_G1873_ = ~new_G1801_ & ~new_G1028_;
  assign new_G1874_ = ~new_G1666_ & ~new_G1801_;
  assign new_G1877_ = ~new_G1748_ & ~new_G1805_;
  assign new_G1878_ = ~new_G1805_ & ~new_G1076_;
  assign new_G1879_ = ~new_G1670_ & ~new_G1805_;
  assign new_G1882_ = ~new_G1751_ & ~new_G1809_;
  assign new_G1883_ = ~new_G1809_ & ~new_G1124_;
  assign new_G1884_ = ~new_G1674_ & ~new_G1809_;
  assign new_G1887_ = ~new_G1754_ & ~new_G1813_;
  assign new_G1888_ = ~new_G1813_ & ~new_G1172_;
  assign new_G1889_ = ~new_G1678_ & ~new_G1813_;
  assign new_G1892_ = ~new_G1817_ & ~new_G1818_;
  assign new_G1895_ = ~new_G1268_ & ~new_G1819_;
  assign new_G1899_ = ~new_G1827_ & ~new_G1828_;
  assign new_G1902_ = ~new_G1832_ & ~new_G1833_;
  assign new_G1905_ = ~new_G1837_ & ~new_G1838_;
  assign new_G1908_ = ~new_G1842_ & ~new_G1843_;
  assign new_G1911_ = ~new_G1847_ & ~new_G1848_;
  assign new_G1914_ = ~new_G1852_ & ~new_G1853_;
  assign new_G1917_ = ~new_G1857_ & ~new_G1858_;
  assign new_G1920_ = ~new_G1862_ & ~new_G1863_;
  assign new_G1923_ = ~new_G1867_ & ~new_G1868_;
  assign new_G1926_ = ~new_G1872_ & ~new_G1873_;
  assign new_G1929_ = ~new_G1877_ & ~new_G1878_;
  assign new_G1932_ = ~new_G1882_ & ~new_G1883_;
  assign new_G1935_ = ~new_G1887_ & ~new_G1888_;
  assign new_G1938_ = ~new_G1892_ & ~new_G1889_;
  assign new_G1942_ = ~new_G1268_ & ~new_G1895_;
  assign new_G1943_ = ~new_G1895_ & ~new_G1819_;
  assign new_G1944_ = ~new_G1899_ & ~new_G1824_;
  assign new_G1948_ = ~new_G1902_ & ~new_G1829_;
  assign new_G1952_ = ~new_G1905_ & ~new_G1834_;
  assign new_G1956_ = ~new_G1908_ & ~new_G1839_;
  assign new_G1960_ = ~new_G1911_ & ~new_G1844_;
  assign new_G1964_ = ~new_G1914_ & ~new_G1849_;
  assign new_G1968_ = ~new_G1917_ & ~new_G1854_;
  assign new_G1972_ = ~new_G1920_ & ~new_G1859_;
  assign new_G1976_ = ~new_G1923_ & ~new_G1864_;
  assign new_G1980_ = ~new_G1926_ & ~new_G1869_;
  assign new_G1984_ = ~new_G1929_ & ~new_G1874_;
  assign new_G1988_ = ~new_G1932_ & ~new_G1879_;
  assign new_G1992_ = ~new_G1935_ & ~new_G1884_;
  assign new_G1996_ = ~new_G1892_ & ~new_G1938_;
  assign new_G1997_ = ~new_G1938_ & ~new_G1889_;
  assign new_G1998_ = ~new_G1942_ & ~new_G1943_;
  assign new_G2001_ = ~new_G1899_ & ~new_G1944_;
  assign new_G2002_ = ~new_G1944_ & ~new_G1824_;
  assign new_G2003_ = ~new_G1902_ & ~new_G1948_;
  assign new_G2004_ = ~new_G1948_ & ~new_G1829_;
  assign new_G2005_ = ~new_G1905_ & ~new_G1952_;
  assign new_G2006_ = ~new_G1952_ & ~new_G1834_;
  assign new_G2007_ = ~new_G1908_ & ~new_G1956_;
  assign new_G2008_ = ~new_G1956_ & ~new_G1839_;
  assign new_G2009_ = ~new_G1911_ & ~new_G1960_;
  assign new_G2010_ = ~new_G1960_ & ~new_G1844_;
  assign new_G2011_ = ~new_G1914_ & ~new_G1964_;
  assign new_G2012_ = ~new_G1964_ & ~new_G1849_;
  assign new_G2013_ = ~new_G1917_ & ~new_G1968_;
  assign new_G2014_ = ~new_G1968_ & ~new_G1854_;
  assign new_G2015_ = ~new_G1920_ & ~new_G1972_;
  assign new_G2016_ = ~new_G1972_ & ~new_G1859_;
  assign new_G2017_ = ~new_G1923_ & ~new_G1976_;
  assign new_G2018_ = ~new_G1976_ & ~new_G1864_;
  assign new_G2019_ = ~new_G1926_ & ~new_G1980_;
  assign new_G2020_ = ~new_G1980_ & ~new_G1869_;
  assign new_G2021_ = ~new_G1929_ & ~new_G1984_;
  assign new_G2022_ = ~new_G1984_ & ~new_G1874_;
  assign new_G2023_ = ~new_G1932_ & ~new_G1988_;
  assign new_G2024_ = ~new_G1988_ & ~new_G1879_;
  assign new_G2025_ = ~new_G1935_ & ~new_G1992_;
  assign new_G2026_ = ~new_G1992_ & ~new_G1884_;
  assign new_G2027_ = ~new_G1996_ & ~new_G1997_;
  assign new_G2030_ = ~new_G1998_ & ~new_G1223_;
  assign new_G2034_ = ~new_G2001_ & ~new_G2002_;
  assign new_G2037_ = ~new_G2003_ & ~new_G2004_;
  assign new_G2040_ = ~new_G2005_ & ~new_G2006_;
  assign new_G2043_ = ~new_G2007_ & ~new_G2008_;
  assign new_G2046_ = ~new_G2009_ & ~new_G2010_;
  assign new_G2049_ = ~new_G2011_ & ~new_G2012_;
  assign new_G2052_ = ~new_G2013_ & ~new_G2014_;
  assign new_G2055_ = ~new_G2015_ & ~new_G2016_;
  assign new_G2058_ = ~new_G2017_ & ~new_G2018_;
  assign new_G2061_ = ~new_G2019_ & ~new_G2020_;
  assign new_G2064_ = ~new_G2021_ & ~new_G2022_;
  assign new_G2067_ = ~new_G2023_ & ~new_G2024_;
  assign new_G2070_ = ~new_G2025_ & ~new_G2026_;
  assign new_G2073_ = ~new_G2027_ & ~new_G1175_;
  assign new_G2077_ = ~new_G1998_ & ~new_G2030_;
  assign new_G2078_ = ~new_G2030_ & ~new_G1223_;
  assign new_G2079_ = ~new_G1895_ & ~new_G2030_;
  assign new_G2082_ = ~new_G2034_ & ~new_G551_;
  assign new_G2086_ = ~new_G2037_ & ~new_G599_;
  assign new_G2090_ = ~new_G2040_ & ~new_G647_;
  assign new_G2094_ = ~new_G2043_ & ~new_G695_;
  assign new_G2098_ = ~new_G2046_ & ~new_G743_;
  assign new_G2102_ = ~new_G2049_ & ~new_G791_;
  assign new_G2106_ = ~new_G2052_ & ~new_G839_;
  assign new_G2110_ = ~new_G2055_ & ~new_G887_;
  assign new_G2114_ = ~new_G2058_ & ~new_G935_;
  assign new_G2118_ = ~new_G2061_ & ~new_G983_;
  assign new_G2122_ = ~new_G2064_ & ~new_G1031_;
  assign new_G2126_ = ~new_G2067_ & ~new_G1079_;
  assign new_G2130_ = ~new_G2070_ & ~new_G1127_;
  assign new_G2134_ = ~new_G2027_ & ~new_G2073_;
  assign new_G2135_ = ~new_G2073_ & ~new_G1175_;
  assign new_G2136_ = ~new_G1938_ & ~new_G2073_;
  assign new_G2139_ = ~new_G2077_ & ~new_G2078_;
  assign new_G2142_ = ~new_G1271_ & ~new_G2079_;
  assign new_G2146_ = ~new_G2034_ & ~new_G2082_;
  assign new_G2147_ = ~new_G2082_ & ~new_G551_;
  assign new_G2148_ = ~new_G1944_ & ~new_G2082_;
  assign new_G2151_ = ~new_G2037_ & ~new_G2086_;
  assign new_G2152_ = ~new_G2086_ & ~new_G599_;
  assign new_G2153_ = ~new_G1948_ & ~new_G2086_;
  assign new_G2156_ = ~new_G2040_ & ~new_G2090_;
  assign new_G2157_ = ~new_G2090_ & ~new_G647_;
  assign new_G2158_ = ~new_G1952_ & ~new_G2090_;
  assign new_G2161_ = ~new_G2043_ & ~new_G2094_;
  assign new_G2162_ = ~new_G2094_ & ~new_G695_;
  assign new_G2163_ = ~new_G1956_ & ~new_G2094_;
  assign new_G2166_ = ~new_G2046_ & ~new_G2098_;
  assign new_G2167_ = ~new_G2098_ & ~new_G743_;
  assign new_G2168_ = ~new_G1960_ & ~new_G2098_;
  assign new_G2171_ = ~new_G2049_ & ~new_G2102_;
  assign new_G2172_ = ~new_G2102_ & ~new_G791_;
  assign new_G2173_ = ~new_G1964_ & ~new_G2102_;
  assign new_G2176_ = ~new_G2052_ & ~new_G2106_;
  assign new_G2177_ = ~new_G2106_ & ~new_G839_;
  assign new_G2178_ = ~new_G1968_ & ~new_G2106_;
  assign new_G2181_ = ~new_G2055_ & ~new_G2110_;
  assign new_G2182_ = ~new_G2110_ & ~new_G887_;
  assign new_G2183_ = ~new_G1972_ & ~new_G2110_;
  assign new_G2186_ = ~new_G2058_ & ~new_G2114_;
  assign new_G2187_ = ~new_G2114_ & ~new_G935_;
  assign new_G2188_ = ~new_G1976_ & ~new_G2114_;
  assign new_G2191_ = ~new_G2061_ & ~new_G2118_;
  assign new_G2192_ = ~new_G2118_ & ~new_G983_;
  assign new_G2193_ = ~new_G1980_ & ~new_G2118_;
  assign new_G2196_ = ~new_G2064_ & ~new_G2122_;
  assign new_G2197_ = ~new_G2122_ & ~new_G1031_;
  assign new_G2198_ = ~new_G1984_ & ~new_G2122_;
  assign new_G2201_ = ~new_G2067_ & ~new_G2126_;
  assign new_G2202_ = ~new_G2126_ & ~new_G1079_;
  assign new_G2203_ = ~new_G1988_ & ~new_G2126_;
  assign new_G2206_ = ~new_G2070_ & ~new_G2130_;
  assign new_G2207_ = ~new_G2130_ & ~new_G1127_;
  assign new_G2208_ = ~new_G1992_ & ~new_G2130_;
  assign new_G2211_ = ~new_G2134_ & ~new_G2135_;
  assign new_G2214_ = ~new_G2139_ & ~new_G2136_;
  assign new_G2218_ = ~new_G1271_ & ~new_G2142_;
  assign new_G2219_ = ~new_G2142_ & ~new_G2079_;
  assign new_G2220_ = ~new_G2151_ & ~new_G2152_;
  assign new_G2223_ = ~new_G2156_ & ~new_G2157_;
  assign new_G2226_ = ~new_G2161_ & ~new_G2162_;
  assign new_G2229_ = ~new_G2166_ & ~new_G2167_;
  assign new_G2232_ = ~new_G2171_ & ~new_G2172_;
  assign new_G2235_ = ~new_G2176_ & ~new_G2177_;
  assign new_G2238_ = ~new_G2181_ & ~new_G2182_;
  assign new_G2241_ = ~new_G2186_ & ~new_G2187_;
  assign new_G2244_ = ~new_G2191_ & ~new_G2192_;
  assign new_G2247_ = ~new_G2196_ & ~new_G2197_;
  assign new_G2250_ = ~new_G2201_ & ~new_G2202_;
  assign new_G2253_ = ~new_G2206_ & ~new_G2207_;
  assign new_G2256_ = ~new_G2211_ & ~new_G2208_;
  assign new_G2260_ = ~new_G2139_ & ~new_G2214_;
  assign new_G2261_ = ~new_G2214_ & ~new_G2136_;
  assign new_G2262_ = ~new_G2218_ & ~new_G2219_;
  assign new_G2265_ = ~new_G2220_ & ~new_G2148_;
  assign new_G2269_ = ~new_G2223_ & ~new_G2153_;
  assign new_G2273_ = ~new_G2226_ & ~new_G2158_;
  assign new_G2277_ = ~new_G2229_ & ~new_G2163_;
  assign new_G2281_ = ~new_G2232_ & ~new_G2168_;
  assign new_G2285_ = ~new_G2235_ & ~new_G2173_;
  assign new_G2289_ = ~new_G2238_ & ~new_G2178_;
  assign new_G2293_ = ~new_G2241_ & ~new_G2183_;
  assign new_G2297_ = ~new_G2244_ & ~new_G2188_;
  assign new_G2301_ = ~new_G2247_ & ~new_G2193_;
  assign new_G2305_ = ~new_G2250_ & ~new_G2198_;
  assign new_G2309_ = ~new_G2253_ & ~new_G2203_;
  assign new_G2313_ = ~new_G2211_ & ~new_G2256_;
  assign new_G2314_ = ~new_G2256_ & ~new_G2208_;
  assign new_G2315_ = ~new_G2260_ & ~new_G2261_;
  assign new_G2318_ = ~new_G2262_ & ~new_G1226_;
  assign new_G2322_ = ~new_G2220_ & ~new_G2265_;
  assign new_G2323_ = ~new_G2265_ & ~new_G2148_;
  assign new_G2324_ = ~new_G2223_ & ~new_G2269_;
  assign new_G2325_ = ~new_G2269_ & ~new_G2153_;
  assign new_G2326_ = ~new_G2226_ & ~new_G2273_;
  assign new_G2327_ = ~new_G2273_ & ~new_G2158_;
  assign new_G2328_ = ~new_G2229_ & ~new_G2277_;
  assign new_G2329_ = ~new_G2277_ & ~new_G2163_;
  assign new_G2330_ = ~new_G2232_ & ~new_G2281_;
  assign new_G2331_ = ~new_G2281_ & ~new_G2168_;
  assign new_G2332_ = ~new_G2235_ & ~new_G2285_;
  assign new_G2333_ = ~new_G2285_ & ~new_G2173_;
  assign new_G2334_ = ~new_G2238_ & ~new_G2289_;
  assign new_G2335_ = ~new_G2289_ & ~new_G2178_;
  assign new_G2336_ = ~new_G2241_ & ~new_G2293_;
  assign new_G2337_ = ~new_G2293_ & ~new_G2183_;
  assign new_G2338_ = ~new_G2244_ & ~new_G2297_;
  assign new_G2339_ = ~new_G2297_ & ~new_G2188_;
  assign new_G2340_ = ~new_G2247_ & ~new_G2301_;
  assign new_G2341_ = ~new_G2301_ & ~new_G2193_;
  assign new_G2342_ = ~new_G2250_ & ~new_G2305_;
  assign new_G2343_ = ~new_G2305_ & ~new_G2198_;
  assign new_G2344_ = ~new_G2253_ & ~new_G2309_;
  assign new_G2345_ = ~new_G2309_ & ~new_G2203_;
  assign new_G2346_ = ~new_G2313_ & ~new_G2314_;
  assign new_G2349_ = ~new_G2315_ & ~new_G1178_;
  assign new_G2353_ = ~new_G2262_ & ~new_G2318_;
  assign new_G2354_ = ~new_G2318_ & ~new_G1226_;
  assign new_G2355_ = ~new_G2142_ & ~new_G2318_;
  assign new_G2358_ = ~new_G2322_ & ~new_G2323_;
  assign new_G2361_ = ~new_G2324_ & ~new_G2325_;
  assign new_G2364_ = ~new_G2326_ & ~new_G2327_;
  assign new_G2367_ = ~new_G2328_ & ~new_G2329_;
  assign new_G2370_ = ~new_G2330_ & ~new_G2331_;
  assign new_G2373_ = ~new_G2332_ & ~new_G2333_;
  assign new_G2376_ = ~new_G2334_ & ~new_G2335_;
  assign new_G2379_ = ~new_G2336_ & ~new_G2337_;
  assign new_G2382_ = ~new_G2338_ & ~new_G2339_;
  assign new_G2385_ = ~new_G2340_ & ~new_G2341_;
  assign new_G2388_ = ~new_G2342_ & ~new_G2343_;
  assign new_G2391_ = ~new_G2344_ & ~new_G2345_;
  assign new_G2394_ = ~new_G2346_ & ~new_G1130_;
  assign new_G2398_ = ~new_G2315_ & ~new_G2349_;
  assign new_G2399_ = ~new_G2349_ & ~new_G1178_;
  assign new_G2400_ = ~new_G2214_ & ~new_G2349_;
  assign new_G2403_ = ~new_G2353_ & ~new_G2354_;
  assign new_G2406_ = ~new_G1274_ & ~new_G2355_;
  assign new_G2410_ = ~new_G2358_ & ~new_G554_;
  assign new_G2414_ = ~new_G2361_ & ~new_G602_;
  assign new_G2418_ = ~new_G2364_ & ~new_G650_;
  assign new_G2422_ = ~new_G2367_ & ~new_G698_;
  assign new_G2426_ = ~new_G2370_ & ~new_G746_;
  assign new_G2430_ = ~new_G2373_ & ~new_G794_;
  assign new_G2434_ = ~new_G2376_ & ~new_G842_;
  assign new_G2438_ = ~new_G2379_ & ~new_G890_;
  assign new_G2442_ = ~new_G2382_ & ~new_G938_;
  assign new_G2446_ = ~new_G2385_ & ~new_G986_;
  assign new_G2450_ = ~new_G2388_ & ~new_G1034_;
  assign new_G2454_ = ~new_G2391_ & ~new_G1082_;
  assign new_G2458_ = ~new_G2346_ & ~new_G2394_;
  assign new_G2459_ = ~new_G2394_ & ~new_G1130_;
  assign new_G2460_ = ~new_G2256_ & ~new_G2394_;
  assign new_G2463_ = ~new_G2398_ & ~new_G2399_;
  assign new_G2466_ = ~new_G2403_ & ~new_G2400_;
  assign new_G2470_ = ~new_G1274_ & ~new_G2406_;
  assign new_G2471_ = ~new_G2406_ & ~new_G2355_;
  assign new_G2472_ = ~new_G2358_ & ~new_G2410_;
  assign new_G2473_ = ~new_G2410_ & ~new_G554_;
  assign new_G2474_ = ~new_G2265_ & ~new_G2410_;
  assign new_G2477_ = ~new_G2361_ & ~new_G2414_;
  assign new_G2478_ = ~new_G2414_ & ~new_G602_;
  assign new_G2479_ = ~new_G2269_ & ~new_G2414_;
  assign new_G2482_ = ~new_G2364_ & ~new_G2418_;
  assign new_G2483_ = ~new_G2418_ & ~new_G650_;
  assign new_G2484_ = ~new_G2273_ & ~new_G2418_;
  assign new_G2487_ = ~new_G2367_ & ~new_G2422_;
  assign new_G2488_ = ~new_G2422_ & ~new_G698_;
  assign new_G2489_ = ~new_G2277_ & ~new_G2422_;
  assign new_G2492_ = ~new_G2370_ & ~new_G2426_;
  assign new_G2493_ = ~new_G2426_ & ~new_G746_;
  assign new_G2494_ = ~new_G2281_ & ~new_G2426_;
  assign new_G2497_ = ~new_G2373_ & ~new_G2430_;
  assign new_G2498_ = ~new_G2430_ & ~new_G794_;
  assign new_G2499_ = ~new_G2285_ & ~new_G2430_;
  assign new_G2502_ = ~new_G2376_ & ~new_G2434_;
  assign new_G2503_ = ~new_G2434_ & ~new_G842_;
  assign new_G2504_ = ~new_G2289_ & ~new_G2434_;
  assign new_G2507_ = ~new_G2379_ & ~new_G2438_;
  assign new_G2508_ = ~new_G2438_ & ~new_G890_;
  assign new_G2509_ = ~new_G2293_ & ~new_G2438_;
  assign new_G2512_ = ~new_G2382_ & ~new_G2442_;
  assign new_G2513_ = ~new_G2442_ & ~new_G938_;
  assign new_G2514_ = ~new_G2297_ & ~new_G2442_;
  assign new_G2517_ = ~new_G2385_ & ~new_G2446_;
  assign new_G2518_ = ~new_G2446_ & ~new_G986_;
  assign new_G2519_ = ~new_G2301_ & ~new_G2446_;
  assign new_G2522_ = ~new_G2388_ & ~new_G2450_;
  assign new_G2523_ = ~new_G2450_ & ~new_G1034_;
  assign new_G2524_ = ~new_G2305_ & ~new_G2450_;
  assign new_G2527_ = ~new_G2391_ & ~new_G2454_;
  assign new_G2528_ = ~new_G2454_ & ~new_G1082_;
  assign new_G2529_ = ~new_G2309_ & ~new_G2454_;
  assign new_G2532_ = ~new_G2458_ & ~new_G2459_;
  assign new_G2535_ = ~new_G2463_ & ~new_G2460_;
  assign new_G2539_ = ~new_G2403_ & ~new_G2466_;
  assign new_G2540_ = ~new_G2466_ & ~new_G2400_;
  assign new_G2541_ = ~new_G2470_ & ~new_G2471_;
  assign new_G2544_ = ~new_G2477_ & ~new_G2478_;
  assign new_G2547_ = ~new_G2482_ & ~new_G2483_;
  assign new_G2550_ = ~new_G2487_ & ~new_G2488_;
  assign new_G2553_ = ~new_G2492_ & ~new_G2493_;
  assign new_G2556_ = ~new_G2497_ & ~new_G2498_;
  assign new_G2559_ = ~new_G2502_ & ~new_G2503_;
  assign new_G2562_ = ~new_G2507_ & ~new_G2508_;
  assign new_G2565_ = ~new_G2512_ & ~new_G2513_;
  assign new_G2568_ = ~new_G2517_ & ~new_G2518_;
  assign new_G2571_ = ~new_G2522_ & ~new_G2523_;
  assign new_G2574_ = ~new_G2527_ & ~new_G2528_;
  assign new_G2577_ = ~new_G2532_ & ~new_G2529_;
  assign new_G2581_ = ~new_G2463_ & ~new_G2535_;
  assign new_G2582_ = ~new_G2535_ & ~new_G2460_;
  assign new_G2583_ = ~new_G2539_ & ~new_G2540_;
  assign new_G2586_ = ~new_G2541_ & ~new_G1229_;
  assign new_G2590_ = ~new_G2544_ & ~new_G2474_;
  assign new_G2594_ = ~new_G2547_ & ~new_G2479_;
  assign new_G2598_ = ~new_G2550_ & ~new_G2484_;
  assign new_G2602_ = ~new_G2553_ & ~new_G2489_;
  assign new_G2606_ = ~new_G2556_ & ~new_G2494_;
  assign new_G2610_ = ~new_G2559_ & ~new_G2499_;
  assign new_G2614_ = ~new_G2562_ & ~new_G2504_;
  assign new_G2618_ = ~new_G2565_ & ~new_G2509_;
  assign new_G2622_ = ~new_G2568_ & ~new_G2514_;
  assign new_G2626_ = ~new_G2571_ & ~new_G2519_;
  assign new_G2630_ = ~new_G2574_ & ~new_G2524_;
  assign new_G2634_ = ~new_G2532_ & ~new_G2577_;
  assign new_G2635_ = ~new_G2577_ & ~new_G2529_;
  assign new_G2636_ = ~new_G2581_ & ~new_G2582_;
  assign new_G2639_ = ~new_G2583_ & ~new_G1181_;
  assign new_G2643_ = ~new_G2541_ & ~new_G2586_;
  assign new_G2644_ = ~new_G2586_ & ~new_G1229_;
  assign new_G2645_ = ~new_G2406_ & ~new_G2586_;
  assign new_G2648_ = ~new_G2544_ & ~new_G2590_;
  assign new_G2649_ = ~new_G2590_ & ~new_G2474_;
  assign new_G2650_ = ~new_G2547_ & ~new_G2594_;
  assign new_G2651_ = ~new_G2594_ & ~new_G2479_;
  assign new_G2652_ = ~new_G2550_ & ~new_G2598_;
  assign new_G2653_ = ~new_G2598_ & ~new_G2484_;
  assign new_G2654_ = ~new_G2553_ & ~new_G2602_;
  assign new_G2655_ = ~new_G2602_ & ~new_G2489_;
  assign new_G2656_ = ~new_G2556_ & ~new_G2606_;
  assign new_G2657_ = ~new_G2606_ & ~new_G2494_;
  assign new_G2658_ = ~new_G2559_ & ~new_G2610_;
  assign new_G2659_ = ~new_G2610_ & ~new_G2499_;
  assign new_G2660_ = ~new_G2562_ & ~new_G2614_;
  assign new_G2661_ = ~new_G2614_ & ~new_G2504_;
  assign new_G2662_ = ~new_G2565_ & ~new_G2618_;
  assign new_G2663_ = ~new_G2618_ & ~new_G2509_;
  assign new_G2664_ = ~new_G2568_ & ~new_G2622_;
  assign new_G2665_ = ~new_G2622_ & ~new_G2514_;
  assign new_G2666_ = ~new_G2571_ & ~new_G2626_;
  assign new_G2667_ = ~new_G2626_ & ~new_G2519_;
  assign new_G2668_ = ~new_G2574_ & ~new_G2630_;
  assign new_G2669_ = ~new_G2630_ & ~new_G2524_;
  assign new_G2670_ = ~new_G2634_ & ~new_G2635_;
  assign new_G2673_ = ~new_G2636_ & ~new_G1133_;
  assign new_G2677_ = ~new_G2583_ & ~new_G2639_;
  assign new_G2678_ = ~new_G2639_ & ~new_G1181_;
  assign new_G2679_ = ~new_G2466_ & ~new_G2639_;
  assign new_G2682_ = ~new_G2643_ & ~new_G2644_;
  assign new_G2685_ = ~new_G1277_ & ~new_G2645_;
  assign new_G2689_ = ~new_G2648_ & ~new_G2649_;
  assign new_G2692_ = ~new_G2650_ & ~new_G2651_;
  assign new_G2695_ = ~new_G2652_ & ~new_G2653_;
  assign new_G2698_ = ~new_G2654_ & ~new_G2655_;
  assign new_G2701_ = ~new_G2656_ & ~new_G2657_;
  assign new_G2704_ = ~new_G2658_ & ~new_G2659_;
  assign new_G2707_ = ~new_G2660_ & ~new_G2661_;
  assign new_G2710_ = ~new_G2662_ & ~new_G2663_;
  assign new_G2713_ = ~new_G2664_ & ~new_G2665_;
  assign new_G2716_ = ~new_G2666_ & ~new_G2667_;
  assign new_G2719_ = ~new_G2668_ & ~new_G2669_;
  assign new_G2722_ = ~new_G2670_ & ~new_G1085_;
  assign new_G2726_ = ~new_G2636_ & ~new_G2673_;
  assign new_G2727_ = ~new_G2673_ & ~new_G1133_;
  assign new_G2728_ = ~new_G2535_ & ~new_G2673_;
  assign new_G2731_ = ~new_G2677_ & ~new_G2678_;
  assign new_G2734_ = ~new_G2682_ & ~new_G2679_;
  assign new_G2738_ = ~new_G1277_ & ~new_G2685_;
  assign new_G2739_ = ~new_G2685_ & ~new_G2645_;
  assign new_G2740_ = ~new_G2689_ & ~new_G557_;
  assign new_G2744_ = ~new_G2692_ & ~new_G605_;
  assign new_G2748_ = ~new_G2695_ & ~new_G653_;
  assign new_G2752_ = ~new_G2698_ & ~new_G701_;
  assign new_G2756_ = ~new_G2701_ & ~new_G749_;
  assign new_G2760_ = ~new_G2704_ & ~new_G797_;
  assign new_G2764_ = ~new_G2707_ & ~new_G845_;
  assign new_G2768_ = ~new_G2710_ & ~new_G893_;
  assign new_G2772_ = ~new_G2713_ & ~new_G941_;
  assign new_G2776_ = ~new_G2716_ & ~new_G989_;
  assign new_G2780_ = ~new_G2719_ & ~new_G1037_;
  assign new_G2784_ = ~new_G2670_ & ~new_G2722_;
  assign new_G2785_ = ~new_G2722_ & ~new_G1085_;
  assign new_G2786_ = ~new_G2577_ & ~new_G2722_;
  assign new_G2789_ = ~new_G2726_ & ~new_G2727_;
  assign new_G2792_ = ~new_G2731_ & ~new_G2728_;
  assign new_G2796_ = ~new_G2682_ & ~new_G2734_;
  assign new_G2797_ = ~new_G2734_ & ~new_G2679_;
  assign new_G2798_ = ~new_G2738_ & ~new_G2739_;
  assign new_G2801_ = ~new_G2689_ & ~new_G2740_;
  assign new_G2802_ = ~new_G2740_ & ~new_G557_;
  assign new_G2803_ = ~new_G2590_ & ~new_G2740_;
  assign new_G2806_ = ~new_G2692_ & ~new_G2744_;
  assign new_G2807_ = ~new_G2744_ & ~new_G605_;
  assign new_G2808_ = ~new_G2594_ & ~new_G2744_;
  assign new_G2811_ = ~new_G2695_ & ~new_G2748_;
  assign new_G2812_ = ~new_G2748_ & ~new_G653_;
  assign new_G2813_ = ~new_G2598_ & ~new_G2748_;
  assign new_G2816_ = ~new_G2698_ & ~new_G2752_;
  assign new_G2817_ = ~new_G2752_ & ~new_G701_;
  assign new_G2818_ = ~new_G2602_ & ~new_G2752_;
  assign new_G2821_ = ~new_G2701_ & ~new_G2756_;
  assign new_G2822_ = ~new_G2756_ & ~new_G749_;
  assign new_G2823_ = ~new_G2606_ & ~new_G2756_;
  assign new_G2826_ = ~new_G2704_ & ~new_G2760_;
  assign new_G2827_ = ~new_G2760_ & ~new_G797_;
  assign new_G2828_ = ~new_G2610_ & ~new_G2760_;
  assign new_G2831_ = ~new_G2707_ & ~new_G2764_;
  assign new_G2832_ = ~new_G2764_ & ~new_G845_;
  assign new_G2833_ = ~new_G2614_ & ~new_G2764_;
  assign new_G2836_ = ~new_G2710_ & ~new_G2768_;
  assign new_G2837_ = ~new_G2768_ & ~new_G893_;
  assign new_G2838_ = ~new_G2618_ & ~new_G2768_;
  assign new_G2841_ = ~new_G2713_ & ~new_G2772_;
  assign new_G2842_ = ~new_G2772_ & ~new_G941_;
  assign new_G2843_ = ~new_G2622_ & ~new_G2772_;
  assign new_G2846_ = ~new_G2716_ & ~new_G2776_;
  assign new_G2847_ = ~new_G2776_ & ~new_G989_;
  assign new_G2848_ = ~new_G2626_ & ~new_G2776_;
  assign new_G2851_ = ~new_G2719_ & ~new_G2780_;
  assign new_G2852_ = ~new_G2780_ & ~new_G1037_;
  assign new_G2853_ = ~new_G2630_ & ~new_G2780_;
  assign new_G2856_ = ~new_G2784_ & ~new_G2785_;
  assign new_G2859_ = ~new_G2789_ & ~new_G2786_;
  assign new_G2863_ = ~new_G2731_ & ~new_G2792_;
  assign new_G2864_ = ~new_G2792_ & ~new_G2728_;
  assign new_G2865_ = ~new_G2796_ & ~new_G2797_;
  assign new_G2868_ = ~new_G2798_ & ~new_G1232_;
  assign new_G2872_ = ~new_G2806_ & ~new_G2807_;
  assign new_G2875_ = ~new_G2811_ & ~new_G2812_;
  assign new_G2878_ = ~new_G2816_ & ~new_G2817_;
  assign new_G2881_ = ~new_G2821_ & ~new_G2822_;
  assign new_G2884_ = ~new_G2826_ & ~new_G2827_;
  assign new_G2887_ = ~new_G2831_ & ~new_G2832_;
  assign new_G2890_ = ~new_G2836_ & ~new_G2837_;
  assign new_G2893_ = ~new_G2841_ & ~new_G2842_;
  assign new_G2896_ = ~new_G2846_ & ~new_G2847_;
  assign new_G2899_ = ~new_G2851_ & ~new_G2852_;
  assign new_G2902_ = ~new_G2856_ & ~new_G2853_;
  assign new_G2906_ = ~new_G2789_ & ~new_G2859_;
  assign new_G2907_ = ~new_G2859_ & ~new_G2786_;
  assign new_G2908_ = ~new_G2863_ & ~new_G2864_;
  assign new_G2911_ = ~new_G2865_ & ~new_G1184_;
  assign new_G2915_ = ~new_G2798_ & ~new_G2868_;
  assign new_G2916_ = ~new_G2868_ & ~new_G1232_;
  assign new_G2917_ = ~new_G2685_ & ~new_G2868_;
  assign new_G2920_ = ~new_G2872_ & ~new_G2803_;
  assign new_G2924_ = ~new_G2875_ & ~new_G2808_;
  assign new_G2928_ = ~new_G2878_ & ~new_G2813_;
  assign new_G2932_ = ~new_G2881_ & ~new_G2818_;
  assign new_G2936_ = ~new_G2884_ & ~new_G2823_;
  assign new_G2940_ = ~new_G2887_ & ~new_G2828_;
  assign new_G2944_ = ~new_G2890_ & ~new_G2833_;
  assign new_G2948_ = ~new_G2893_ & ~new_G2838_;
  assign new_G2952_ = ~new_G2896_ & ~new_G2843_;
  assign new_G2956_ = ~new_G2899_ & ~new_G2848_;
  assign new_G2960_ = ~new_G2856_ & ~new_G2902_;
  assign new_G2961_ = ~new_G2902_ & ~new_G2853_;
  assign new_G2962_ = ~new_G2906_ & ~new_G2907_;
  assign new_G2965_ = ~new_G2908_ & ~new_G1136_;
  assign new_G2969_ = ~new_G2865_ & ~new_G2911_;
  assign new_G2970_ = ~new_G2911_ & ~new_G1184_;
  assign new_G2971_ = ~new_G2734_ & ~new_G2911_;
  assign new_G2974_ = ~new_G2915_ & ~new_G2916_;
  assign new_G2977_ = ~new_G1280_ & ~new_G2917_;
  assign new_G2981_ = ~new_G2872_ & ~new_G2920_;
  assign new_G2982_ = ~new_G2920_ & ~new_G2803_;
  assign new_G2983_ = ~new_G2875_ & ~new_G2924_;
  assign new_G2984_ = ~new_G2924_ & ~new_G2808_;
  assign new_G2985_ = ~new_G2878_ & ~new_G2928_;
  assign new_G2986_ = ~new_G2928_ & ~new_G2813_;
  assign new_G2987_ = ~new_G2881_ & ~new_G2932_;
  assign new_G2988_ = ~new_G2932_ & ~new_G2818_;
  assign new_G2989_ = ~new_G2884_ & ~new_G2936_;
  assign new_G2990_ = ~new_G2936_ & ~new_G2823_;
  assign new_G2991_ = ~new_G2887_ & ~new_G2940_;
  assign new_G2992_ = ~new_G2940_ & ~new_G2828_;
  assign new_G2993_ = ~new_G2890_ & ~new_G2944_;
  assign new_G2994_ = ~new_G2944_ & ~new_G2833_;
  assign new_G2995_ = ~new_G2893_ & ~new_G2948_;
  assign new_G2996_ = ~new_G2948_ & ~new_G2838_;
  assign new_G2997_ = ~new_G2896_ & ~new_G2952_;
  assign new_G2998_ = ~new_G2952_ & ~new_G2843_;
  assign new_G2999_ = ~new_G2899_ & ~new_G2956_;
  assign new_G3000_ = ~new_G2956_ & ~new_G2848_;
  assign new_G3001_ = ~new_G2960_ & ~new_G2961_;
  assign new_G3004_ = ~new_G2962_ & ~new_G1088_;
  assign new_G3008_ = ~new_G2908_ & ~new_G2965_;
  assign new_G3009_ = ~new_G2965_ & ~new_G1136_;
  assign new_G3010_ = ~new_G2792_ & ~new_G2965_;
  assign new_G3013_ = ~new_G2969_ & ~new_G2970_;
  assign new_G3016_ = ~new_G2974_ & ~new_G2971_;
  assign new_G3020_ = ~new_G1280_ & ~new_G2977_;
  assign new_G3021_ = ~new_G2977_ & ~new_G2917_;
  assign new_G3022_ = ~new_G2981_ & ~new_G2982_;
  assign new_G3025_ = ~new_G2983_ & ~new_G2984_;
  assign new_G3028_ = ~new_G2985_ & ~new_G2986_;
  assign new_G3031_ = ~new_G2987_ & ~new_G2988_;
  assign new_G3034_ = ~new_G2989_ & ~new_G2990_;
  assign new_G3037_ = ~new_G2991_ & ~new_G2992_;
  assign new_G3040_ = ~new_G2993_ & ~new_G2994_;
  assign new_G3043_ = ~new_G2995_ & ~new_G2996_;
  assign new_G3046_ = ~new_G2997_ & ~new_G2998_;
  assign new_G3049_ = ~new_G2999_ & ~new_G3000_;
  assign new_G3052_ = ~new_G3001_ & ~new_G1040_;
  assign new_G3056_ = ~new_G2962_ & ~new_G3004_;
  assign new_G3057_ = ~new_G3004_ & ~new_G1088_;
  assign new_G3058_ = ~new_G2859_ & ~new_G3004_;
  assign new_G3061_ = ~new_G3008_ & ~new_G3009_;
  assign new_G3064_ = ~new_G3013_ & ~new_G3010_;
  assign new_G3068_ = ~new_G2974_ & ~new_G3016_;
  assign new_G3069_ = ~new_G3016_ & ~new_G2971_;
  assign new_G3070_ = ~new_G3020_ & ~new_G3021_;
  assign new_G3073_ = ~new_G3022_ & ~new_G560_;
  assign new_G3077_ = ~new_G3025_ & ~new_G608_;
  assign new_G3081_ = ~new_G3028_ & ~new_G656_;
  assign new_G3085_ = ~new_G3031_ & ~new_G704_;
  assign new_G3089_ = ~new_G3034_ & ~new_G752_;
  assign new_G3093_ = ~new_G3037_ & ~new_G800_;
  assign new_G3097_ = ~new_G3040_ & ~new_G848_;
  assign new_G3101_ = ~new_G3043_ & ~new_G896_;
  assign new_G3105_ = ~new_G3046_ & ~new_G944_;
  assign new_G3109_ = ~new_G3049_ & ~new_G992_;
  assign new_G3113_ = ~new_G3001_ & ~new_G3052_;
  assign new_G3114_ = ~new_G3052_ & ~new_G1040_;
  assign new_G3115_ = ~new_G2902_ & ~new_G3052_;
  assign new_G3118_ = ~new_G3056_ & ~new_G3057_;
  assign new_G3121_ = ~new_G3061_ & ~new_G3058_;
  assign new_G3125_ = ~new_G3013_ & ~new_G3064_;
  assign new_G3126_ = ~new_G3064_ & ~new_G3010_;
  assign new_G3127_ = ~new_G3068_ & ~new_G3069_;
  assign new_G3130_ = ~new_G3070_ & ~new_G1235_;
  assign new_G3134_ = ~new_G3022_ & ~new_G3073_;
  assign new_G3135_ = ~new_G3073_ & ~new_G560_;
  assign new_G3136_ = ~new_G2920_ & ~new_G3073_;
  assign new_G3139_ = ~new_G3025_ & ~new_G3077_;
  assign new_G3140_ = ~new_G3077_ & ~new_G608_;
  assign new_G3141_ = ~new_G2924_ & ~new_G3077_;
  assign new_G3144_ = ~new_G3028_ & ~new_G3081_;
  assign new_G3145_ = ~new_G3081_ & ~new_G656_;
  assign new_G3146_ = ~new_G2928_ & ~new_G3081_;
  assign new_G3149_ = ~new_G3031_ & ~new_G3085_;
  assign new_G3150_ = ~new_G3085_ & ~new_G704_;
  assign new_G3151_ = ~new_G2932_ & ~new_G3085_;
  assign new_G3154_ = ~new_G3034_ & ~new_G3089_;
  assign new_G3155_ = ~new_G3089_ & ~new_G752_;
  assign new_G3156_ = ~new_G2936_ & ~new_G3089_;
  assign new_G3159_ = ~new_G3037_ & ~new_G3093_;
  assign new_G3160_ = ~new_G3093_ & ~new_G800_;
  assign new_G3161_ = ~new_G2940_ & ~new_G3093_;
  assign new_G3164_ = ~new_G3040_ & ~new_G3097_;
  assign new_G3165_ = ~new_G3097_ & ~new_G848_;
  assign new_G3166_ = ~new_G2944_ & ~new_G3097_;
  assign new_G3169_ = ~new_G3043_ & ~new_G3101_;
  assign new_G3170_ = ~new_G3101_ & ~new_G896_;
  assign new_G3171_ = ~new_G2948_ & ~new_G3101_;
  assign new_G3174_ = ~new_G3046_ & ~new_G3105_;
  assign new_G3175_ = ~new_G3105_ & ~new_G944_;
  assign new_G3176_ = ~new_G2952_ & ~new_G3105_;
  assign new_G3179_ = ~new_G3049_ & ~new_G3109_;
  assign new_G3180_ = ~new_G3109_ & ~new_G992_;
  assign new_G3181_ = ~new_G2956_ & ~new_G3109_;
  assign new_G3184_ = ~new_G3113_ & ~new_G3114_;
  assign new_G3187_ = ~new_G3118_ & ~new_G3115_;
  assign new_G3191_ = ~new_G3061_ & ~new_G3121_;
  assign new_G3192_ = ~new_G3121_ & ~new_G3058_;
  assign new_G3193_ = ~new_G3125_ & ~new_G3126_;
  assign new_G3196_ = ~new_G3127_ & ~new_G1187_;
  assign new_G3200_ = ~new_G3070_ & ~new_G3130_;
  assign new_G3201_ = ~new_G3130_ & ~new_G1235_;
  assign new_G3202_ = ~new_G2977_ & ~new_G3130_;
  assign new_G3205_ = ~new_G3139_ & ~new_G3140_;
  assign new_G3208_ = ~new_G3144_ & ~new_G3145_;
  assign new_G3211_ = ~new_G3149_ & ~new_G3150_;
  assign new_G3214_ = ~new_G3154_ & ~new_G3155_;
  assign new_G3217_ = ~new_G3159_ & ~new_G3160_;
  assign new_G3220_ = ~new_G3164_ & ~new_G3165_;
  assign new_G3223_ = ~new_G3169_ & ~new_G3170_;
  assign new_G3226_ = ~new_G3174_ & ~new_G3175_;
  assign new_G3229_ = ~new_G3179_ & ~new_G3180_;
  assign new_G3232_ = ~new_G3184_ & ~new_G3181_;
  assign new_G3236_ = ~new_G3118_ & ~new_G3187_;
  assign new_G3237_ = ~new_G3187_ & ~new_G3115_;
  assign new_G3238_ = ~new_G3191_ & ~new_G3192_;
  assign new_G3241_ = ~new_G3193_ & ~new_G1139_;
  assign new_G3245_ = ~new_G3127_ & ~new_G3196_;
  assign new_G3246_ = ~new_G3196_ & ~new_G1187_;
  assign new_G3247_ = ~new_G3016_ & ~new_G3196_;
  assign new_G3250_ = ~new_G3200_ & ~new_G3201_;
  assign new_G3253_ = ~new_G1283_ & ~new_G3202_;
  assign new_G3257_ = ~new_G3205_ & ~new_G3136_;
  assign new_G3261_ = ~new_G3208_ & ~new_G3141_;
  assign new_G3265_ = ~new_G3211_ & ~new_G3146_;
  assign new_G3269_ = ~new_G3214_ & ~new_G3151_;
  assign new_G3273_ = ~new_G3217_ & ~new_G3156_;
  assign new_G3277_ = ~new_G3220_ & ~new_G3161_;
  assign new_G3281_ = ~new_G3223_ & ~new_G3166_;
  assign new_G3285_ = ~new_G3226_ & ~new_G3171_;
  assign new_G3289_ = ~new_G3229_ & ~new_G3176_;
  assign new_G3293_ = ~new_G3184_ & ~new_G3232_;
  assign new_G3294_ = ~new_G3232_ & ~new_G3181_;
  assign new_G3295_ = ~new_G3236_ & ~new_G3237_;
  assign new_G3298_ = ~new_G3238_ & ~new_G1091_;
  assign new_G3302_ = ~new_G3193_ & ~new_G3241_;
  assign new_G3303_ = ~new_G3241_ & ~new_G1139_;
  assign new_G3304_ = ~new_G3064_ & ~new_G3241_;
  assign new_G3307_ = ~new_G3245_ & ~new_G3246_;
  assign new_G3310_ = ~new_G3250_ & ~new_G3247_;
  assign new_G3314_ = ~new_G1283_ & ~new_G3253_;
  assign new_G3315_ = ~new_G3253_ & ~new_G3202_;
  assign new_G3316_ = ~new_G3205_ & ~new_G3257_;
  assign new_G3317_ = ~new_G3257_ & ~new_G3136_;
  assign new_G3318_ = ~new_G3208_ & ~new_G3261_;
  assign new_G3319_ = ~new_G3261_ & ~new_G3141_;
  assign new_G3320_ = ~new_G3211_ & ~new_G3265_;
  assign new_G3321_ = ~new_G3265_ & ~new_G3146_;
  assign new_G3322_ = ~new_G3214_ & ~new_G3269_;
  assign new_G3323_ = ~new_G3269_ & ~new_G3151_;
  assign new_G3324_ = ~new_G3217_ & ~new_G3273_;
  assign new_G3325_ = ~new_G3273_ & ~new_G3156_;
  assign new_G3326_ = ~new_G3220_ & ~new_G3277_;
  assign new_G3327_ = ~new_G3277_ & ~new_G3161_;
  assign new_G3328_ = ~new_G3223_ & ~new_G3281_;
  assign new_G3329_ = ~new_G3281_ & ~new_G3166_;
  assign new_G3330_ = ~new_G3226_ & ~new_G3285_;
  assign new_G3331_ = ~new_G3285_ & ~new_G3171_;
  assign new_G3332_ = ~new_G3229_ & ~new_G3289_;
  assign new_G3333_ = ~new_G3289_ & ~new_G3176_;
  assign new_G3334_ = ~new_G3293_ & ~new_G3294_;
  assign new_G3337_ = ~new_G3295_ & ~new_G1043_;
  assign new_G3341_ = ~new_G3238_ & ~new_G3298_;
  assign new_G3342_ = ~new_G3298_ & ~new_G1091_;
  assign new_G3343_ = ~new_G3121_ & ~new_G3298_;
  assign new_G3346_ = ~new_G3302_ & ~new_G3303_;
  assign new_G3349_ = ~new_G3307_ & ~new_G3304_;
  assign new_G3353_ = ~new_G3250_ & ~new_G3310_;
  assign new_G3354_ = ~new_G3310_ & ~new_G3247_;
  assign new_G3355_ = ~new_G3314_ & ~new_G3315_;
  assign new_G3358_ = ~new_G3316_ & ~new_G3317_;
  assign new_G3361_ = ~new_G3318_ & ~new_G3319_;
  assign new_G3364_ = ~new_G3320_ & ~new_G3321_;
  assign new_G3367_ = ~new_G3322_ & ~new_G3323_;
  assign new_G3370_ = ~new_G3324_ & ~new_G3325_;
  assign new_G3373_ = ~new_G3326_ & ~new_G3327_;
  assign new_G3376_ = ~new_G3328_ & ~new_G3329_;
  assign new_G3379_ = ~new_G3330_ & ~new_G3331_;
  assign new_G3382_ = ~new_G3332_ & ~new_G3333_;
  assign new_G3385_ = ~new_G3334_ & ~new_G995_;
  assign new_G3389_ = ~new_G3295_ & ~new_G3337_;
  assign new_G3390_ = ~new_G3337_ & ~new_G1043_;
  assign new_G3391_ = ~new_G3187_ & ~new_G3337_;
  assign new_G3394_ = ~new_G3341_ & ~new_G3342_;
  assign new_G3397_ = ~new_G3346_ & ~new_G3343_;
  assign new_G3401_ = ~new_G3307_ & ~new_G3349_;
  assign new_G3402_ = ~new_G3349_ & ~new_G3304_;
  assign new_G3403_ = ~new_G3353_ & ~new_G3354_;
  assign new_G3406_ = ~new_G3355_ & ~new_G1238_;
  assign new_G3410_ = ~new_G3358_ & ~new_G563_;
  assign new_G3414_ = ~new_G3361_ & ~new_G611_;
  assign new_G3418_ = ~new_G3364_ & ~new_G659_;
  assign new_G3422_ = ~new_G3367_ & ~new_G707_;
  assign new_G3426_ = ~new_G3370_ & ~new_G755_;
  assign new_G3430_ = ~new_G3373_ & ~new_G803_;
  assign new_G3434_ = ~new_G3376_ & ~new_G851_;
  assign new_G3438_ = ~new_G3379_ & ~new_G899_;
  assign new_G3442_ = ~new_G3382_ & ~new_G947_;
  assign new_G3446_ = ~new_G3334_ & ~new_G3385_;
  assign new_G3447_ = ~new_G3385_ & ~new_G995_;
  assign new_G3448_ = ~new_G3232_ & ~new_G3385_;
  assign new_G3451_ = ~new_G3389_ & ~new_G3390_;
  assign new_G3454_ = ~new_G3394_ & ~new_G3391_;
  assign new_G3458_ = ~new_G3346_ & ~new_G3397_;
  assign new_G3459_ = ~new_G3397_ & ~new_G3343_;
  assign new_G3460_ = ~new_G3401_ & ~new_G3402_;
  assign new_G3463_ = ~new_G3403_ & ~new_G1190_;
  assign new_G3467_ = ~new_G3355_ & ~new_G3406_;
  assign new_G3468_ = ~new_G3406_ & ~new_G1238_;
  assign new_G3469_ = ~new_G3253_ & ~new_G3406_;
  assign new_G3472_ = ~new_G3358_ & ~new_G3410_;
  assign new_G3473_ = ~new_G3410_ & ~new_G563_;
  assign new_G3474_ = ~new_G3257_ & ~new_G3410_;
  assign new_G3477_ = ~new_G3361_ & ~new_G3414_;
  assign new_G3478_ = ~new_G3414_ & ~new_G611_;
  assign new_G3479_ = ~new_G3261_ & ~new_G3414_;
  assign new_G3482_ = ~new_G3364_ & ~new_G3418_;
  assign new_G3483_ = ~new_G3418_ & ~new_G659_;
  assign new_G3484_ = ~new_G3265_ & ~new_G3418_;
  assign new_G3487_ = ~new_G3367_ & ~new_G3422_;
  assign new_G3488_ = ~new_G3422_ & ~new_G707_;
  assign new_G3489_ = ~new_G3269_ & ~new_G3422_;
  assign new_G3492_ = ~new_G3370_ & ~new_G3426_;
  assign new_G3493_ = ~new_G3426_ & ~new_G755_;
  assign new_G3494_ = ~new_G3273_ & ~new_G3426_;
  assign new_G3497_ = ~new_G3373_ & ~new_G3430_;
  assign new_G3498_ = ~new_G3430_ & ~new_G803_;
  assign new_G3499_ = ~new_G3277_ & ~new_G3430_;
  assign new_G3502_ = ~new_G3376_ & ~new_G3434_;
  assign new_G3503_ = ~new_G3434_ & ~new_G851_;
  assign new_G3504_ = ~new_G3281_ & ~new_G3434_;
  assign new_G3507_ = ~new_G3379_ & ~new_G3438_;
  assign new_G3508_ = ~new_G3438_ & ~new_G899_;
  assign new_G3509_ = ~new_G3285_ & ~new_G3438_;
  assign new_G3512_ = ~new_G3382_ & ~new_G3442_;
  assign new_G3513_ = ~new_G3442_ & ~new_G947_;
  assign new_G3514_ = ~new_G3289_ & ~new_G3442_;
  assign new_G3517_ = ~new_G3446_ & ~new_G3447_;
  assign new_G3520_ = ~new_G3451_ & ~new_G3448_;
  assign new_G3524_ = ~new_G3394_ & ~new_G3454_;
  assign new_G3525_ = ~new_G3454_ & ~new_G3391_;
  assign new_G3526_ = ~new_G3458_ & ~new_G3459_;
  assign new_G3529_ = ~new_G3460_ & ~new_G1142_;
  assign new_G3533_ = ~new_G3403_ & ~new_G3463_;
  assign new_G3534_ = ~new_G3463_ & ~new_G1190_;
  assign new_G3535_ = ~new_G3310_ & ~new_G3463_;
  assign new_G3538_ = ~new_G3467_ & ~new_G3468_;
  assign new_G3541_ = ~new_G1286_ & ~new_G3469_;
  assign new_G3545_ = ~new_G3477_ & ~new_G3478_;
  assign new_G3548_ = ~new_G3482_ & ~new_G3483_;
  assign new_G3551_ = ~new_G3487_ & ~new_G3488_;
  assign new_G3554_ = ~new_G3492_ & ~new_G3493_;
  assign new_G3557_ = ~new_G3497_ & ~new_G3498_;
  assign new_G3560_ = ~new_G3502_ & ~new_G3503_;
  assign new_G3563_ = ~new_G3507_ & ~new_G3508_;
  assign new_G3566_ = ~new_G3512_ & ~new_G3513_;
  assign new_G3569_ = ~new_G3517_ & ~new_G3514_;
  assign new_G3573_ = ~new_G3451_ & ~new_G3520_;
  assign new_G3574_ = ~new_G3520_ & ~new_G3448_;
  assign new_G3575_ = ~new_G3524_ & ~new_G3525_;
  assign new_G3578_ = ~new_G3526_ & ~new_G1094_;
  assign new_G3582_ = ~new_G3460_ & ~new_G3529_;
  assign new_G3583_ = ~new_G3529_ & ~new_G1142_;
  assign new_G3584_ = ~new_G3349_ & ~new_G3529_;
  assign new_G3587_ = ~new_G3533_ & ~new_G3534_;
  assign new_G3590_ = ~new_G3538_ & ~new_G3535_;
  assign new_G3594_ = ~new_G1286_ & ~new_G3541_;
  assign new_G3595_ = ~new_G3541_ & ~new_G3469_;
  assign new_G3596_ = ~new_G3545_ & ~new_G3474_;
  assign new_G3600_ = ~new_G3548_ & ~new_G3479_;
  assign new_G3604_ = ~new_G3551_ & ~new_G3484_;
  assign new_G3608_ = ~new_G3554_ & ~new_G3489_;
  assign new_G3612_ = ~new_G3557_ & ~new_G3494_;
  assign new_G3616_ = ~new_G3560_ & ~new_G3499_;
  assign new_G3620_ = ~new_G3563_ & ~new_G3504_;
  assign new_G3624_ = ~new_G3566_ & ~new_G3509_;
  assign new_G3628_ = ~new_G3517_ & ~new_G3569_;
  assign new_G3629_ = ~new_G3569_ & ~new_G3514_;
  assign new_G3630_ = ~new_G3573_ & ~new_G3574_;
  assign new_G3633_ = ~new_G3575_ & ~new_G1046_;
  assign new_G3637_ = ~new_G3526_ & ~new_G3578_;
  assign new_G3638_ = ~new_G3578_ & ~new_G1094_;
  assign new_G3639_ = ~new_G3397_ & ~new_G3578_;
  assign new_G3642_ = ~new_G3582_ & ~new_G3583_;
  assign new_G3645_ = ~new_G3587_ & ~new_G3584_;
  assign new_G3649_ = ~new_G3538_ & ~new_G3590_;
  assign new_G3650_ = ~new_G3590_ & ~new_G3535_;
  assign new_G3651_ = ~new_G3594_ & ~new_G3595_;
  assign new_G3654_ = ~new_G3545_ & ~new_G3596_;
  assign new_G3655_ = ~new_G3596_ & ~new_G3474_;
  assign new_G3656_ = ~new_G3548_ & ~new_G3600_;
  assign new_G3657_ = ~new_G3600_ & ~new_G3479_;
  assign new_G3658_ = ~new_G3551_ & ~new_G3604_;
  assign new_G3659_ = ~new_G3604_ & ~new_G3484_;
  assign new_G3660_ = ~new_G3554_ & ~new_G3608_;
  assign new_G3661_ = ~new_G3608_ & ~new_G3489_;
  assign new_G3662_ = ~new_G3557_ & ~new_G3612_;
  assign new_G3663_ = ~new_G3612_ & ~new_G3494_;
  assign new_G3664_ = ~new_G3560_ & ~new_G3616_;
  assign new_G3665_ = ~new_G3616_ & ~new_G3499_;
  assign new_G3666_ = ~new_G3563_ & ~new_G3620_;
  assign new_G3667_ = ~new_G3620_ & ~new_G3504_;
  assign new_G3668_ = ~new_G3566_ & ~new_G3624_;
  assign new_G3669_ = ~new_G3624_ & ~new_G3509_;
  assign new_G3670_ = ~new_G3628_ & ~new_G3629_;
  assign new_G3673_ = ~new_G3630_ & ~new_G998_;
  assign new_G3677_ = ~new_G3575_ & ~new_G3633_;
  assign new_G3678_ = ~new_G3633_ & ~new_G1046_;
  assign new_G3679_ = ~new_G3454_ & ~new_G3633_;
  assign new_G3682_ = ~new_G3637_ & ~new_G3638_;
  assign new_G3685_ = ~new_G3642_ & ~new_G3639_;
  assign new_G3689_ = ~new_G3587_ & ~new_G3645_;
  assign new_G3690_ = ~new_G3645_ & ~new_G3584_;
  assign new_G3691_ = ~new_G3649_ & ~new_G3650_;
  assign new_G3694_ = ~new_G3651_ & ~new_G1241_;
  assign new_G3698_ = ~new_G3654_ & ~new_G3655_;
  assign new_G3701_ = ~new_G3656_ & ~new_G3657_;
  assign new_G3704_ = ~new_G3658_ & ~new_G3659_;
  assign new_G3707_ = ~new_G3660_ & ~new_G3661_;
  assign new_G3710_ = ~new_G3662_ & ~new_G3663_;
  assign new_G3713_ = ~new_G3664_ & ~new_G3665_;
  assign new_G3716_ = ~new_G3666_ & ~new_G3667_;
  assign new_G3719_ = ~new_G3668_ & ~new_G3669_;
  assign new_G3722_ = ~new_G3670_ & ~new_G950_;
  assign new_G3726_ = ~new_G3630_ & ~new_G3673_;
  assign new_G3727_ = ~new_G3673_ & ~new_G998_;
  assign new_G3728_ = ~new_G3520_ & ~new_G3673_;
  assign new_G3731_ = ~new_G3677_ & ~new_G3678_;
  assign new_G3734_ = ~new_G3682_ & ~new_G3679_;
  assign new_G3738_ = ~new_G3642_ & ~new_G3685_;
  assign new_G3739_ = ~new_G3685_ & ~new_G3639_;
  assign new_G3740_ = ~new_G3689_ & ~new_G3690_;
  assign new_G3743_ = ~new_G3691_ & ~new_G1193_;
  assign new_G3747_ = ~new_G3651_ & ~new_G3694_;
  assign new_G3748_ = ~new_G3694_ & ~new_G1241_;
  assign new_G3749_ = ~new_G3541_ & ~new_G3694_;
  assign new_G3752_ = ~new_G3698_ & ~new_G566_;
  assign new_G3756_ = ~new_G3701_ & ~new_G614_;
  assign new_G3760_ = ~new_G3704_ & ~new_G662_;
  assign new_G3764_ = ~new_G3707_ & ~new_G710_;
  assign new_G3768_ = ~new_G3710_ & ~new_G758_;
  assign new_G3772_ = ~new_G3713_ & ~new_G806_;
  assign new_G3776_ = ~new_G3716_ & ~new_G854_;
  assign new_G3780_ = ~new_G3719_ & ~new_G902_;
  assign new_G3784_ = ~new_G3670_ & ~new_G3722_;
  assign new_G3785_ = ~new_G3722_ & ~new_G950_;
  assign new_G3786_ = ~new_G3569_ & ~new_G3722_;
  assign new_G3789_ = ~new_G3726_ & ~new_G3727_;
  assign new_G3792_ = ~new_G3731_ & ~new_G3728_;
  assign new_G3796_ = ~new_G3682_ & ~new_G3734_;
  assign new_G3797_ = ~new_G3734_ & ~new_G3679_;
  assign new_G3798_ = ~new_G3738_ & ~new_G3739_;
  assign new_G3801_ = ~new_G3740_ & ~new_G1145_;
  assign new_G3805_ = ~new_G3691_ & ~new_G3743_;
  assign new_G3806_ = ~new_G3743_ & ~new_G1193_;
  assign new_G3807_ = ~new_G3590_ & ~new_G3743_;
  assign new_G3810_ = ~new_G3747_ & ~new_G3748_;
  assign new_G3813_ = ~new_G1289_ & ~new_G3749_;
  assign new_G3817_ = ~new_G3698_ & ~new_G3752_;
  assign new_G3818_ = ~new_G3752_ & ~new_G566_;
  assign new_G3819_ = ~new_G3596_ & ~new_G3752_;
  assign new_G3822_ = ~new_G3701_ & ~new_G3756_;
  assign new_G3823_ = ~new_G3756_ & ~new_G614_;
  assign new_G3824_ = ~new_G3600_ & ~new_G3756_;
  assign new_G3827_ = ~new_G3704_ & ~new_G3760_;
  assign new_G3828_ = ~new_G3760_ & ~new_G662_;
  assign new_G3829_ = ~new_G3604_ & ~new_G3760_;
  assign new_G3832_ = ~new_G3707_ & ~new_G3764_;
  assign new_G3833_ = ~new_G3764_ & ~new_G710_;
  assign new_G3834_ = ~new_G3608_ & ~new_G3764_;
  assign new_G3837_ = ~new_G3710_ & ~new_G3768_;
  assign new_G3838_ = ~new_G3768_ & ~new_G758_;
  assign new_G3839_ = ~new_G3612_ & ~new_G3768_;
  assign new_G3842_ = ~new_G3713_ & ~new_G3772_;
  assign new_G3843_ = ~new_G3772_ & ~new_G806_;
  assign new_G3844_ = ~new_G3616_ & ~new_G3772_;
  assign new_G3847_ = ~new_G3716_ & ~new_G3776_;
  assign new_G3848_ = ~new_G3776_ & ~new_G854_;
  assign new_G3849_ = ~new_G3620_ & ~new_G3776_;
  assign new_G3852_ = ~new_G3719_ & ~new_G3780_;
  assign new_G3853_ = ~new_G3780_ & ~new_G902_;
  assign new_G3854_ = ~new_G3624_ & ~new_G3780_;
  assign new_G3857_ = ~new_G3784_ & ~new_G3785_;
  assign new_G3860_ = ~new_G3789_ & ~new_G3786_;
  assign new_G3864_ = ~new_G3731_ & ~new_G3792_;
  assign new_G3865_ = ~new_G3792_ & ~new_G3728_;
  assign new_G3866_ = ~new_G3796_ & ~new_G3797_;
  assign new_G3869_ = ~new_G3798_ & ~new_G1097_;
  assign new_G3873_ = ~new_G3740_ & ~new_G3801_;
  assign new_G3874_ = ~new_G3801_ & ~new_G1145_;
  assign new_G3875_ = ~new_G3645_ & ~new_G3801_;
  assign new_G3878_ = ~new_G3805_ & ~new_G3806_;
  assign new_G3881_ = ~new_G3810_ & ~new_G3807_;
  assign new_G3885_ = ~new_G1289_ & ~new_G3813_;
  assign new_G3886_ = ~new_G3813_ & ~new_G3749_;
  assign new_G3887_ = ~new_G3822_ & ~new_G3823_;
  assign new_G3890_ = ~new_G3827_ & ~new_G3828_;
  assign new_G3893_ = ~new_G3832_ & ~new_G3833_;
  assign new_G3896_ = ~new_G3837_ & ~new_G3838_;
  assign new_G3899_ = ~new_G3842_ & ~new_G3843_;
  assign new_G3902_ = ~new_G3847_ & ~new_G3848_;
  assign new_G3905_ = ~new_G3852_ & ~new_G3853_;
  assign new_G3908_ = ~new_G3857_ & ~new_G3854_;
  assign new_G3912_ = ~new_G3789_ & ~new_G3860_;
  assign new_G3913_ = ~new_G3860_ & ~new_G3786_;
  assign new_G3914_ = ~new_G3864_ & ~new_G3865_;
  assign new_G3917_ = ~new_G3866_ & ~new_G1049_;
  assign new_G3921_ = ~new_G3798_ & ~new_G3869_;
  assign new_G3922_ = ~new_G3869_ & ~new_G1097_;
  assign new_G3923_ = ~new_G3685_ & ~new_G3869_;
  assign new_G3926_ = ~new_G3873_ & ~new_G3874_;
  assign new_G3929_ = ~new_G3878_ & ~new_G3875_;
  assign new_G3933_ = ~new_G3810_ & ~new_G3881_;
  assign new_G3934_ = ~new_G3881_ & ~new_G3807_;
  assign new_G3935_ = ~new_G3885_ & ~new_G3886_;
  assign new_G3938_ = ~new_G3887_ & ~new_G3819_;
  assign new_G3942_ = ~new_G3890_ & ~new_G3824_;
  assign new_G3946_ = ~new_G3893_ & ~new_G3829_;
  assign new_G3950_ = ~new_G3896_ & ~new_G3834_;
  assign new_G3954_ = ~new_G3899_ & ~new_G3839_;
  assign new_G3958_ = ~new_G3902_ & ~new_G3844_;
  assign new_G3962_ = ~new_G3905_ & ~new_G3849_;
  assign new_G3966_ = ~new_G3857_ & ~new_G3908_;
  assign new_G3967_ = ~new_G3908_ & ~new_G3854_;
  assign new_G3968_ = ~new_G3912_ & ~new_G3913_;
  assign new_G3971_ = ~new_G3914_ & ~new_G1001_;
  assign new_G3975_ = ~new_G3866_ & ~new_G3917_;
  assign new_G3976_ = ~new_G3917_ & ~new_G1049_;
  assign new_G3977_ = ~new_G3734_ & ~new_G3917_;
  assign new_G3980_ = ~new_G3921_ & ~new_G3922_;
  assign new_G3983_ = ~new_G3926_ & ~new_G3923_;
  assign new_G3987_ = ~new_G3878_ & ~new_G3929_;
  assign new_G3988_ = ~new_G3929_ & ~new_G3875_;
  assign new_G3989_ = ~new_G3933_ & ~new_G3934_;
  assign new_G3992_ = ~new_G3935_ & ~new_G1244_;
  assign new_G3996_ = ~new_G3887_ & ~new_G3938_;
  assign new_G3997_ = ~new_G3938_ & ~new_G3819_;
  assign new_G3998_ = ~new_G3890_ & ~new_G3942_;
  assign new_G3999_ = ~new_G3942_ & ~new_G3824_;
  assign new_G4000_ = ~new_G3893_ & ~new_G3946_;
  assign new_G4001_ = ~new_G3946_ & ~new_G3829_;
  assign new_G4002_ = ~new_G3896_ & ~new_G3950_;
  assign new_G4003_ = ~new_G3950_ & ~new_G3834_;
  assign new_G4004_ = ~new_G3899_ & ~new_G3954_;
  assign new_G4005_ = ~new_G3954_ & ~new_G3839_;
  assign new_G4006_ = ~new_G3902_ & ~new_G3958_;
  assign new_G4007_ = ~new_G3958_ & ~new_G3844_;
  assign new_G4008_ = ~new_G3905_ & ~new_G3962_;
  assign new_G4009_ = ~new_G3962_ & ~new_G3849_;
  assign new_G4010_ = ~new_G3966_ & ~new_G3967_;
  assign new_G4013_ = ~new_G3968_ & ~new_G953_;
  assign new_G4017_ = ~new_G3914_ & ~new_G3971_;
  assign new_G4018_ = ~new_G3971_ & ~new_G1001_;
  assign new_G4019_ = ~new_G3792_ & ~new_G3971_;
  assign new_G4022_ = ~new_G3975_ & ~new_G3976_;
  assign new_G4025_ = ~new_G3980_ & ~new_G3977_;
  assign new_G4029_ = ~new_G3926_ & ~new_G3983_;
  assign new_G4030_ = ~new_G3983_ & ~new_G3923_;
  assign new_G4031_ = ~new_G3987_ & ~new_G3988_;
  assign new_G4034_ = ~new_G3989_ & ~new_G1196_;
  assign new_G4038_ = ~new_G3935_ & ~new_G3992_;
  assign new_G4039_ = ~new_G3992_ & ~new_G1244_;
  assign new_G4040_ = ~new_G3813_ & ~new_G3992_;
  assign new_G4043_ = ~new_G3996_ & ~new_G3997_;
  assign new_G4046_ = ~new_G3998_ & ~new_G3999_;
  assign new_G4049_ = ~new_G4000_ & ~new_G4001_;
  assign new_G4052_ = ~new_G4002_ & ~new_G4003_;
  assign new_G4055_ = ~new_G4004_ & ~new_G4005_;
  assign new_G4058_ = ~new_G4006_ & ~new_G4007_;
  assign new_G4061_ = ~new_G4008_ & ~new_G4009_;
  assign new_G4064_ = ~new_G4010_ & ~new_G905_;
  assign new_G4068_ = ~new_G3968_ & ~new_G4013_;
  assign new_G4069_ = ~new_G4013_ & ~new_G953_;
  assign new_G4070_ = ~new_G3860_ & ~new_G4013_;
  assign new_G4073_ = ~new_G4017_ & ~new_G4018_;
  assign new_G4076_ = ~new_G4022_ & ~new_G4019_;
  assign new_G4080_ = ~new_G3980_ & ~new_G4025_;
  assign new_G4081_ = ~new_G4025_ & ~new_G3977_;
  assign new_G4082_ = ~new_G4029_ & ~new_G4030_;
  assign new_G4085_ = ~new_G4031_ & ~new_G1148_;
  assign new_G4089_ = ~new_G3989_ & ~new_G4034_;
  assign new_G4090_ = ~new_G4034_ & ~new_G1196_;
  assign new_G4091_ = ~new_G3881_ & ~new_G4034_;
  assign new_G4094_ = ~new_G4038_ & ~new_G4039_;
  assign new_G4097_ = ~new_G1292_ & ~new_G4040_;
  assign new_G4101_ = ~new_G4043_ & ~new_G569_;
  assign new_G4105_ = ~new_G4046_ & ~new_G617_;
  assign new_G4109_ = ~new_G4049_ & ~new_G665_;
  assign new_G4113_ = ~new_G4052_ & ~new_G713_;
  assign new_G4117_ = ~new_G4055_ & ~new_G761_;
  assign new_G4121_ = ~new_G4058_ & ~new_G809_;
  assign new_G4125_ = ~new_G4061_ & ~new_G857_;
  assign new_G4129_ = ~new_G4010_ & ~new_G4064_;
  assign new_G4130_ = ~new_G4064_ & ~new_G905_;
  assign new_G4131_ = ~new_G3908_ & ~new_G4064_;
  assign new_G4134_ = ~new_G4068_ & ~new_G4069_;
  assign new_G4137_ = ~new_G4073_ & ~new_G4070_;
  assign new_G4141_ = ~new_G4022_ & ~new_G4076_;
  assign new_G4142_ = ~new_G4076_ & ~new_G4019_;
  assign new_G4143_ = ~new_G4080_ & ~new_G4081_;
  assign new_G4146_ = ~new_G4082_ & ~new_G1100_;
  assign new_G4150_ = ~new_G4031_ & ~new_G4085_;
  assign new_G4151_ = ~new_G4085_ & ~new_G1148_;
  assign new_G4152_ = ~new_G3929_ & ~new_G4085_;
  assign new_G4155_ = ~new_G4089_ & ~new_G4090_;
  assign new_G4158_ = ~new_G4094_ & ~new_G4091_;
  assign new_G4162_ = ~new_G1292_ & ~new_G4097_;
  assign new_G4163_ = ~new_G4097_ & ~new_G4040_;
  assign new_G4164_ = ~new_G4043_ & ~new_G4101_;
  assign new_G4165_ = ~new_G4101_ & ~new_G569_;
  assign new_G4166_ = ~new_G3938_ & ~new_G4101_;
  assign new_G4169_ = ~new_G4046_ & ~new_G4105_;
  assign new_G4170_ = ~new_G4105_ & ~new_G617_;
  assign new_G4171_ = ~new_G3942_ & ~new_G4105_;
  assign new_G4174_ = ~new_G4049_ & ~new_G4109_;
  assign new_G4175_ = ~new_G4109_ & ~new_G665_;
  assign new_G4176_ = ~new_G3946_ & ~new_G4109_;
  assign new_G4179_ = ~new_G4052_ & ~new_G4113_;
  assign new_G4180_ = ~new_G4113_ & ~new_G713_;
  assign new_G4181_ = ~new_G3950_ & ~new_G4113_;
  assign new_G4184_ = ~new_G4055_ & ~new_G4117_;
  assign new_G4185_ = ~new_G4117_ & ~new_G761_;
  assign new_G4186_ = ~new_G3954_ & ~new_G4117_;
  assign new_G4189_ = ~new_G4058_ & ~new_G4121_;
  assign new_G4190_ = ~new_G4121_ & ~new_G809_;
  assign new_G4191_ = ~new_G3958_ & ~new_G4121_;
  assign new_G4194_ = ~new_G4061_ & ~new_G4125_;
  assign new_G4195_ = ~new_G4125_ & ~new_G857_;
  assign new_G4196_ = ~new_G3962_ & ~new_G4125_;
  assign new_G4199_ = ~new_G4129_ & ~new_G4130_;
  assign new_G4202_ = ~new_G4134_ & ~new_G4131_;
  assign new_G4206_ = ~new_G4073_ & ~new_G4137_;
  assign new_G4207_ = ~new_G4137_ & ~new_G4070_;
  assign new_G4208_ = ~new_G4141_ & ~new_G4142_;
  assign new_G4211_ = ~new_G4143_ & ~new_G1052_;
  assign new_G4215_ = ~new_G4082_ & ~new_G4146_;
  assign new_G4216_ = ~new_G4146_ & ~new_G1100_;
  assign new_G4217_ = ~new_G3983_ & ~new_G4146_;
  assign new_G4220_ = ~new_G4150_ & ~new_G4151_;
  assign new_G4223_ = ~new_G4155_ & ~new_G4152_;
  assign new_G4227_ = ~new_G4094_ & ~new_G4158_;
  assign new_G4228_ = ~new_G4158_ & ~new_G4091_;
  assign new_G4229_ = ~new_G4162_ & ~new_G4163_;
  assign new_G4232_ = ~new_G4169_ & ~new_G4170_;
  assign new_G4235_ = ~new_G4174_ & ~new_G4175_;
  assign new_G4238_ = ~new_G4179_ & ~new_G4180_;
  assign new_G4241_ = ~new_G4184_ & ~new_G4185_;
  assign new_G4244_ = ~new_G4189_ & ~new_G4190_;
  assign new_G4247_ = ~new_G4194_ & ~new_G4195_;
  assign new_G4250_ = ~new_G4199_ & ~new_G4196_;
  assign new_G4254_ = ~new_G4134_ & ~new_G4202_;
  assign new_G4255_ = ~new_G4202_ & ~new_G4131_;
  assign new_G4256_ = ~new_G4206_ & ~new_G4207_;
  assign new_G4259_ = ~new_G4208_ & ~new_G1004_;
  assign new_G4263_ = ~new_G4143_ & ~new_G4211_;
  assign new_G4264_ = ~new_G4211_ & ~new_G1052_;
  assign new_G4265_ = ~new_G4025_ & ~new_G4211_;
  assign new_G4268_ = ~new_G4215_ & ~new_G4216_;
  assign new_G4271_ = ~new_G4220_ & ~new_G4217_;
  assign new_G4275_ = ~new_G4155_ & ~new_G4223_;
  assign new_G4276_ = ~new_G4223_ & ~new_G4152_;
  assign new_G4277_ = ~new_G4227_ & ~new_G4228_;
  assign new_G4280_ = ~new_G4229_ & ~new_G1247_;
  assign new_G4284_ = ~new_G4232_ & ~new_G4166_;
  assign new_G4288_ = ~new_G4235_ & ~new_G4171_;
  assign new_G4292_ = ~new_G4238_ & ~new_G4176_;
  assign new_G4296_ = ~new_G4241_ & ~new_G4181_;
  assign new_G4300_ = ~new_G4244_ & ~new_G4186_;
  assign new_G4304_ = ~new_G4247_ & ~new_G4191_;
  assign new_G4308_ = ~new_G4199_ & ~new_G4250_;
  assign new_G4309_ = ~new_G4250_ & ~new_G4196_;
  assign new_G4310_ = ~new_G4254_ & ~new_G4255_;
  assign new_G4313_ = ~new_G4256_ & ~new_G956_;
  assign new_G4317_ = ~new_G4208_ & ~new_G4259_;
  assign new_G4318_ = ~new_G4259_ & ~new_G1004_;
  assign new_G4319_ = ~new_G4076_ & ~new_G4259_;
  assign new_G4322_ = ~new_G4263_ & ~new_G4264_;
  assign new_G4325_ = ~new_G4268_ & ~new_G4265_;
  assign new_G4329_ = ~new_G4220_ & ~new_G4271_;
  assign new_G4330_ = ~new_G4271_ & ~new_G4217_;
  assign new_G4331_ = ~new_G4275_ & ~new_G4276_;
  assign new_G4334_ = ~new_G4277_ & ~new_G1199_;
  assign new_G4338_ = ~new_G4229_ & ~new_G4280_;
  assign new_G4339_ = ~new_G4280_ & ~new_G1247_;
  assign new_G4340_ = ~new_G4097_ & ~new_G4280_;
  assign new_G4343_ = ~new_G4232_ & ~new_G4284_;
  assign new_G4344_ = ~new_G4284_ & ~new_G4166_;
  assign new_G4345_ = ~new_G4235_ & ~new_G4288_;
  assign new_G4346_ = ~new_G4288_ & ~new_G4171_;
  assign new_G4347_ = ~new_G4238_ & ~new_G4292_;
  assign new_G4348_ = ~new_G4292_ & ~new_G4176_;
  assign new_G4349_ = ~new_G4241_ & ~new_G4296_;
  assign new_G4350_ = ~new_G4296_ & ~new_G4181_;
  assign new_G4351_ = ~new_G4244_ & ~new_G4300_;
  assign new_G4352_ = ~new_G4300_ & ~new_G4186_;
  assign new_G4353_ = ~new_G4247_ & ~new_G4304_;
  assign new_G4354_ = ~new_G4304_ & ~new_G4191_;
  assign new_G4355_ = ~new_G4308_ & ~new_G4309_;
  assign new_G4358_ = ~new_G4310_ & ~new_G908_;
  assign new_G4362_ = ~new_G4256_ & ~new_G4313_;
  assign new_G4363_ = ~new_G4313_ & ~new_G956_;
  assign new_G4364_ = ~new_G4137_ & ~new_G4313_;
  assign new_G4367_ = ~new_G4317_ & ~new_G4318_;
  assign new_G4370_ = ~new_G4322_ & ~new_G4319_;
  assign new_G4374_ = ~new_G4268_ & ~new_G4325_;
  assign new_G4375_ = ~new_G4325_ & ~new_G4265_;
  assign new_G4376_ = ~new_G4329_ & ~new_G4330_;
  assign new_G4379_ = ~new_G4331_ & ~new_G1151_;
  assign new_G4383_ = ~new_G4277_ & ~new_G4334_;
  assign new_G4384_ = ~new_G4334_ & ~new_G1199_;
  assign new_G4385_ = ~new_G4158_ & ~new_G4334_;
  assign new_G4388_ = ~new_G4338_ & ~new_G4339_;
  assign new_G4391_ = ~new_G1295_ & ~new_G4340_;
  assign new_G4395_ = ~new_G4343_ & ~new_G4344_;
  assign new_G4398_ = ~new_G4345_ & ~new_G4346_;
  assign new_G4401_ = ~new_G4347_ & ~new_G4348_;
  assign new_G4404_ = ~new_G4349_ & ~new_G4350_;
  assign new_G4407_ = ~new_G4351_ & ~new_G4352_;
  assign new_G4410_ = ~new_G4353_ & ~new_G4354_;
  assign new_G4413_ = ~new_G4355_ & ~new_G860_;
  assign new_G4417_ = ~new_G4310_ & ~new_G4358_;
  assign new_G4418_ = ~new_G4358_ & ~new_G908_;
  assign new_G4419_ = ~new_G4202_ & ~new_G4358_;
  assign new_G4422_ = ~new_G4362_ & ~new_G4363_;
  assign new_G4425_ = ~new_G4367_ & ~new_G4364_;
  assign new_G4429_ = ~new_G4322_ & ~new_G4370_;
  assign new_G4430_ = ~new_G4370_ & ~new_G4319_;
  assign new_G4431_ = ~new_G4374_ & ~new_G4375_;
  assign new_G4434_ = ~new_G4376_ & ~new_G1103_;
  assign new_G4438_ = ~new_G4331_ & ~new_G4379_;
  assign new_G4439_ = ~new_G4379_ & ~new_G1151_;
  assign new_G4440_ = ~new_G4223_ & ~new_G4379_;
  assign new_G4443_ = ~new_G4383_ & ~new_G4384_;
  assign new_G4446_ = ~new_G4388_ & ~new_G4385_;
  assign new_G4450_ = ~new_G1295_ & ~new_G4391_;
  assign new_G4451_ = ~new_G4391_ & ~new_G4340_;
  assign new_G4452_ = ~new_G4395_ & ~new_G572_;
  assign new_G4456_ = ~new_G4398_ & ~new_G620_;
  assign new_G4460_ = ~new_G4401_ & ~new_G668_;
  assign new_G4464_ = ~new_G4404_ & ~new_G716_;
  assign new_G4468_ = ~new_G4407_ & ~new_G764_;
  assign new_G4472_ = ~new_G4410_ & ~new_G812_;
  assign new_G4476_ = ~new_G4355_ & ~new_G4413_;
  assign new_G4477_ = ~new_G4413_ & ~new_G860_;
  assign new_G4478_ = ~new_G4250_ & ~new_G4413_;
  assign new_G4481_ = ~new_G4417_ & ~new_G4418_;
  assign new_G4484_ = ~new_G4422_ & ~new_G4419_;
  assign new_G4488_ = ~new_G4367_ & ~new_G4425_;
  assign new_G4489_ = ~new_G4425_ & ~new_G4364_;
  assign new_G4490_ = ~new_G4429_ & ~new_G4430_;
  assign new_G4493_ = ~new_G4431_ & ~new_G1055_;
  assign new_G4497_ = ~new_G4376_ & ~new_G4434_;
  assign new_G4498_ = ~new_G4434_ & ~new_G1103_;
  assign new_G4499_ = ~new_G4271_ & ~new_G4434_;
  assign new_G4502_ = ~new_G4438_ & ~new_G4439_;
  assign new_G4505_ = ~new_G4443_ & ~new_G4440_;
  assign new_G4509_ = ~new_G4388_ & ~new_G4446_;
  assign new_G4510_ = ~new_G4446_ & ~new_G4385_;
  assign new_G4511_ = ~new_G4450_ & ~new_G4451_;
  assign new_G4514_ = ~new_G4395_ & ~new_G4452_;
  assign new_G4515_ = ~new_G4452_ & ~new_G572_;
  assign new_G4516_ = ~new_G4284_ & ~new_G4452_;
  assign new_G4519_ = ~new_G4398_ & ~new_G4456_;
  assign new_G4520_ = ~new_G4456_ & ~new_G620_;
  assign new_G4521_ = ~new_G4288_ & ~new_G4456_;
  assign new_G4524_ = ~new_G4401_ & ~new_G4460_;
  assign new_G4525_ = ~new_G4460_ & ~new_G668_;
  assign new_G4526_ = ~new_G4292_ & ~new_G4460_;
  assign new_G4529_ = ~new_G4404_ & ~new_G4464_;
  assign new_G4530_ = ~new_G4464_ & ~new_G716_;
  assign new_G4531_ = ~new_G4296_ & ~new_G4464_;
  assign new_G4534_ = ~new_G4407_ & ~new_G4468_;
  assign new_G4535_ = ~new_G4468_ & ~new_G764_;
  assign new_G4536_ = ~new_G4300_ & ~new_G4468_;
  assign new_G4539_ = ~new_G4410_ & ~new_G4472_;
  assign new_G4540_ = ~new_G4472_ & ~new_G812_;
  assign new_G4541_ = ~new_G4304_ & ~new_G4472_;
  assign new_G4544_ = ~new_G4476_ & ~new_G4477_;
  assign new_G4547_ = ~new_G4481_ & ~new_G4478_;
  assign new_G4551_ = ~new_G4422_ & ~new_G4484_;
  assign new_G4552_ = ~new_G4484_ & ~new_G4419_;
  assign new_G4553_ = ~new_G4488_ & ~new_G4489_;
  assign new_G4556_ = ~new_G4490_ & ~new_G1007_;
  assign new_G4560_ = ~new_G4431_ & ~new_G4493_;
  assign new_G4561_ = ~new_G4493_ & ~new_G1055_;
  assign new_G4562_ = ~new_G4325_ & ~new_G4493_;
  assign new_G4565_ = ~new_G4497_ & ~new_G4498_;
  assign new_G4568_ = ~new_G4502_ & ~new_G4499_;
  assign new_G4572_ = ~new_G4443_ & ~new_G4505_;
  assign new_G4573_ = ~new_G4505_ & ~new_G4440_;
  assign new_G4574_ = ~new_G4509_ & ~new_G4510_;
  assign new_G4577_ = ~new_G4511_ & ~new_G1250_;
  assign new_G4581_ = ~new_G4519_ & ~new_G4520_;
  assign new_G4584_ = ~new_G4524_ & ~new_G4525_;
  assign new_G4587_ = ~new_G4529_ & ~new_G4530_;
  assign new_G4590_ = ~new_G4534_ & ~new_G4535_;
  assign new_G4593_ = ~new_G4539_ & ~new_G4540_;
  assign new_G4596_ = ~new_G4544_ & ~new_G4541_;
  assign new_G4600_ = ~new_G4481_ & ~new_G4547_;
  assign new_G4601_ = ~new_G4547_ & ~new_G4478_;
  assign new_G4602_ = ~new_G4551_ & ~new_G4552_;
  assign new_G4605_ = ~new_G4553_ & ~new_G959_;
  assign new_G4609_ = ~new_G4490_ & ~new_G4556_;
  assign new_G4610_ = ~new_G4556_ & ~new_G1007_;
  assign new_G4611_ = ~new_G4370_ & ~new_G4556_;
  assign new_G4614_ = ~new_G4560_ & ~new_G4561_;
  assign new_G4617_ = ~new_G4565_ & ~new_G4562_;
  assign new_G4621_ = ~new_G4502_ & ~new_G4568_;
  assign new_G4622_ = ~new_G4568_ & ~new_G4499_;
  assign new_G4623_ = ~new_G4572_ & ~new_G4573_;
  assign new_G4626_ = ~new_G4574_ & ~new_G1202_;
  assign new_G4630_ = ~new_G4511_ & ~new_G4577_;
  assign new_G4631_ = ~new_G4577_ & ~new_G1250_;
  assign new_G4632_ = ~new_G4391_ & ~new_G4577_;
  assign new_G4635_ = ~new_G4581_ & ~new_G4516_;
  assign new_G4639_ = ~new_G4584_ & ~new_G4521_;
  assign new_G4643_ = ~new_G4587_ & ~new_G4526_;
  assign new_G4647_ = ~new_G4590_ & ~new_G4531_;
  assign new_G4651_ = ~new_G4593_ & ~new_G4536_;
  assign new_G4655_ = ~new_G4544_ & ~new_G4596_;
  assign new_G4656_ = ~new_G4596_ & ~new_G4541_;
  assign new_G4657_ = ~new_G4600_ & ~new_G4601_;
  assign new_G4660_ = ~new_G4602_ & ~new_G911_;
  assign new_G4664_ = ~new_G4553_ & ~new_G4605_;
  assign new_G4665_ = ~new_G4605_ & ~new_G959_;
  assign new_G4666_ = ~new_G4425_ & ~new_G4605_;
  assign new_G4669_ = ~new_G4609_ & ~new_G4610_;
  assign new_G4672_ = ~new_G4614_ & ~new_G4611_;
  assign new_G4676_ = ~new_G4565_ & ~new_G4617_;
  assign new_G4677_ = ~new_G4617_ & ~new_G4562_;
  assign new_G4678_ = ~new_G4621_ & ~new_G4622_;
  assign new_G4681_ = ~new_G4623_ & ~new_G1154_;
  assign new_G4685_ = ~new_G4574_ & ~new_G4626_;
  assign new_G4686_ = ~new_G4626_ & ~new_G1202_;
  assign new_G4687_ = ~new_G4446_ & ~new_G4626_;
  assign new_G4690_ = ~new_G4630_ & ~new_G4631_;
  assign new_G4693_ = ~new_G1298_ & ~new_G4632_;
  assign new_G4697_ = ~new_G4581_ & ~new_G4635_;
  assign new_G4698_ = ~new_G4635_ & ~new_G4516_;
  assign new_G4699_ = ~new_G4584_ & ~new_G4639_;
  assign new_G4700_ = ~new_G4639_ & ~new_G4521_;
  assign new_G4701_ = ~new_G4587_ & ~new_G4643_;
  assign new_G4702_ = ~new_G4643_ & ~new_G4526_;
  assign new_G4703_ = ~new_G4590_ & ~new_G4647_;
  assign new_G4704_ = ~new_G4647_ & ~new_G4531_;
  assign new_G4705_ = ~new_G4593_ & ~new_G4651_;
  assign new_G4706_ = ~new_G4651_ & ~new_G4536_;
  assign new_G4707_ = ~new_G4655_ & ~new_G4656_;
  assign new_G4710_ = ~new_G4657_ & ~new_G863_;
  assign new_G4714_ = ~new_G4602_ & ~new_G4660_;
  assign new_G4715_ = ~new_G4660_ & ~new_G911_;
  assign new_G4716_ = ~new_G4484_ & ~new_G4660_;
  assign new_G4719_ = ~new_G4664_ & ~new_G4665_;
  assign new_G4722_ = ~new_G4669_ & ~new_G4666_;
  assign new_G4726_ = ~new_G4614_ & ~new_G4672_;
  assign new_G4727_ = ~new_G4672_ & ~new_G4611_;
  assign new_G4728_ = ~new_G4676_ & ~new_G4677_;
  assign new_G4731_ = ~new_G4678_ & ~new_G1106_;
  assign new_G4735_ = ~new_G4623_ & ~new_G4681_;
  assign new_G4736_ = ~new_G4681_ & ~new_G1154_;
  assign new_G4737_ = ~new_G4505_ & ~new_G4681_;
  assign new_G4740_ = ~new_G4685_ & ~new_G4686_;
  assign new_G4743_ = ~new_G4690_ & ~new_G4687_;
  assign new_G4747_ = ~new_G1298_ & ~new_G4693_;
  assign new_G4748_ = ~new_G4693_ & ~new_G4632_;
  assign new_G4749_ = ~new_G4697_ & ~new_G4698_;
  assign new_G4752_ = ~new_G4699_ & ~new_G4700_;
  assign new_G4755_ = ~new_G4701_ & ~new_G4702_;
  assign new_G4758_ = ~new_G4703_ & ~new_G4704_;
  assign new_G4761_ = ~new_G4705_ & ~new_G4706_;
  assign new_G4764_ = ~new_G4707_ & ~new_G815_;
  assign new_G4768_ = ~new_G4657_ & ~new_G4710_;
  assign new_G4769_ = ~new_G4710_ & ~new_G863_;
  assign new_G4770_ = ~new_G4547_ & ~new_G4710_;
  assign new_G4773_ = ~new_G4714_ & ~new_G4715_;
  assign new_G4776_ = ~new_G4719_ & ~new_G4716_;
  assign new_G4780_ = ~new_G4669_ & ~new_G4722_;
  assign new_G4781_ = ~new_G4722_ & ~new_G4666_;
  assign new_G4782_ = ~new_G4726_ & ~new_G4727_;
  assign new_G4785_ = ~new_G4728_ & ~new_G1058_;
  assign new_G4789_ = ~new_G4678_ & ~new_G4731_;
  assign new_G4790_ = ~new_G4731_ & ~new_G1106_;
  assign new_G4791_ = ~new_G4568_ & ~new_G4731_;
  assign new_G4794_ = ~new_G4735_ & ~new_G4736_;
  assign new_G4797_ = ~new_G4740_ & ~new_G4737_;
  assign new_G4801_ = ~new_G4690_ & ~new_G4743_;
  assign new_G4802_ = ~new_G4743_ & ~new_G4687_;
  assign new_G4803_ = ~new_G4747_ & ~new_G4748_;
  assign new_G4806_ = ~new_G4749_ & ~new_G575_;
  assign new_G4810_ = ~new_G4752_ & ~new_G623_;
  assign new_G4814_ = ~new_G4755_ & ~new_G671_;
  assign new_G4818_ = ~new_G4758_ & ~new_G719_;
  assign new_G4822_ = ~new_G4761_ & ~new_G767_;
  assign new_G4826_ = ~new_G4707_ & ~new_G4764_;
  assign new_G4827_ = ~new_G4764_ & ~new_G815_;
  assign new_G4828_ = ~new_G4596_ & ~new_G4764_;
  assign new_G4831_ = ~new_G4768_ & ~new_G4769_;
  assign new_G4834_ = ~new_G4773_ & ~new_G4770_;
  assign new_G4838_ = ~new_G4719_ & ~new_G4776_;
  assign new_G4839_ = ~new_G4776_ & ~new_G4716_;
  assign new_G4840_ = ~new_G4780_ & ~new_G4781_;
  assign new_G4843_ = ~new_G4782_ & ~new_G1010_;
  assign new_G4847_ = ~new_G4728_ & ~new_G4785_;
  assign new_G4848_ = ~new_G4785_ & ~new_G1058_;
  assign new_G4849_ = ~new_G4617_ & ~new_G4785_;
  assign new_G4852_ = ~new_G4789_ & ~new_G4790_;
  assign new_G4855_ = ~new_G4794_ & ~new_G4791_;
  assign new_G4859_ = ~new_G4740_ & ~new_G4797_;
  assign new_G4860_ = ~new_G4797_ & ~new_G4737_;
  assign new_G4861_ = ~new_G4801_ & ~new_G4802_;
  assign new_G4864_ = ~new_G4803_ & ~new_G1253_;
  assign new_G4868_ = ~new_G4749_ & ~new_G4806_;
  assign new_G4869_ = ~new_G4806_ & ~new_G575_;
  assign new_G4870_ = ~new_G4635_ & ~new_G4806_;
  assign new_G4873_ = ~new_G4752_ & ~new_G4810_;
  assign new_G4874_ = ~new_G4810_ & ~new_G623_;
  assign new_G4875_ = ~new_G4639_ & ~new_G4810_;
  assign new_G4878_ = ~new_G4755_ & ~new_G4814_;
  assign new_G4879_ = ~new_G4814_ & ~new_G671_;
  assign new_G4880_ = ~new_G4643_ & ~new_G4814_;
  assign new_G4883_ = ~new_G4758_ & ~new_G4818_;
  assign new_G4884_ = ~new_G4818_ & ~new_G719_;
  assign new_G4885_ = ~new_G4647_ & ~new_G4818_;
  assign new_G4888_ = ~new_G4761_ & ~new_G4822_;
  assign new_G4889_ = ~new_G4822_ & ~new_G767_;
  assign new_G4890_ = ~new_G4651_ & ~new_G4822_;
  assign new_G4893_ = ~new_G4826_ & ~new_G4827_;
  assign new_G4896_ = ~new_G4831_ & ~new_G4828_;
  assign new_G4900_ = ~new_G4773_ & ~new_G4834_;
  assign new_G4901_ = ~new_G4834_ & ~new_G4770_;
  assign new_G4902_ = ~new_G4838_ & ~new_G4839_;
  assign new_G4905_ = ~new_G4840_ & ~new_G962_;
  assign new_G4909_ = ~new_G4782_ & ~new_G4843_;
  assign new_G4910_ = ~new_G4843_ & ~new_G1010_;
  assign new_G4911_ = ~new_G4672_ & ~new_G4843_;
  assign new_G4914_ = ~new_G4847_ & ~new_G4848_;
  assign new_G4917_ = ~new_G4852_ & ~new_G4849_;
  assign new_G4921_ = ~new_G4794_ & ~new_G4855_;
  assign new_G4922_ = ~new_G4855_ & ~new_G4791_;
  assign new_G4923_ = ~new_G4859_ & ~new_G4860_;
  assign new_G4926_ = ~new_G4861_ & ~new_G1205_;
  assign new_G4930_ = ~new_G4803_ & ~new_G4864_;
  assign new_G4931_ = ~new_G4864_ & ~new_G1253_;
  assign new_G4932_ = ~new_G4693_ & ~new_G4864_;
  assign new_G4935_ = ~new_G4873_ & ~new_G4874_;
  assign new_G4938_ = ~new_G4878_ & ~new_G4879_;
  assign new_G4941_ = ~new_G4883_ & ~new_G4884_;
  assign new_G4944_ = ~new_G4888_ & ~new_G4889_;
  assign new_G4947_ = ~new_G4893_ & ~new_G4890_;
  assign new_G4951_ = ~new_G4831_ & ~new_G4896_;
  assign new_G4952_ = ~new_G4896_ & ~new_G4828_;
  assign new_G4953_ = ~new_G4900_ & ~new_G4901_;
  assign new_G4956_ = ~new_G4902_ & ~new_G914_;
  assign new_G4960_ = ~new_G4840_ & ~new_G4905_;
  assign new_G4961_ = ~new_G4905_ & ~new_G962_;
  assign new_G4962_ = ~new_G4722_ & ~new_G4905_;
  assign new_G4965_ = ~new_G4909_ & ~new_G4910_;
  assign new_G4968_ = ~new_G4914_ & ~new_G4911_;
  assign new_G4972_ = ~new_G4852_ & ~new_G4917_;
  assign new_G4973_ = ~new_G4917_ & ~new_G4849_;
  assign new_G4974_ = ~new_G4921_ & ~new_G4922_;
  assign new_G4977_ = ~new_G4923_ & ~new_G1157_;
  assign new_G4981_ = ~new_G4861_ & ~new_G4926_;
  assign new_G4982_ = ~new_G4926_ & ~new_G1205_;
  assign new_G4983_ = ~new_G4743_ & ~new_G4926_;
  assign new_G4986_ = ~new_G4930_ & ~new_G4931_;
  assign new_G4989_ = ~new_G1301_ & ~new_G4932_;
  assign new_G4993_ = ~new_G4935_ & ~new_G4870_;
  assign new_G4997_ = ~new_G4938_ & ~new_G4875_;
  assign new_G5001_ = ~new_G4941_ & ~new_G4880_;
  assign new_G5005_ = ~new_G4944_ & ~new_G4885_;
  assign new_G5009_ = ~new_G4893_ & ~new_G4947_;
  assign new_G5010_ = ~new_G4947_ & ~new_G4890_;
  assign new_G5011_ = ~new_G4951_ & ~new_G4952_;
  assign new_G5014_ = ~new_G4953_ & ~new_G866_;
  assign new_G5018_ = ~new_G4902_ & ~new_G4956_;
  assign new_G5019_ = ~new_G4956_ & ~new_G914_;
  assign new_G5020_ = ~new_G4776_ & ~new_G4956_;
  assign new_G5023_ = ~new_G4960_ & ~new_G4961_;
  assign new_G5026_ = ~new_G4965_ & ~new_G4962_;
  assign new_G5030_ = ~new_G4914_ & ~new_G4968_;
  assign new_G5031_ = ~new_G4968_ & ~new_G4911_;
  assign new_G5032_ = ~new_G4972_ & ~new_G4973_;
  assign new_G5035_ = ~new_G4974_ & ~new_G1109_;
  assign new_G5039_ = ~new_G4923_ & ~new_G4977_;
  assign new_G5040_ = ~new_G4977_ & ~new_G1157_;
  assign new_G5041_ = ~new_G4797_ & ~new_G4977_;
  assign new_G5044_ = ~new_G4981_ & ~new_G4982_;
  assign new_G5047_ = ~new_G4986_ & ~new_G4983_;
  assign new_G5051_ = ~new_G1301_ & ~new_G4989_;
  assign new_G5052_ = ~new_G4989_ & ~new_G4932_;
  assign new_G5053_ = ~new_G4935_ & ~new_G4993_;
  assign new_G5054_ = ~new_G4993_ & ~new_G4870_;
  assign new_G5055_ = ~new_G4938_ & ~new_G4997_;
  assign new_G5056_ = ~new_G4997_ & ~new_G4875_;
  assign new_G5057_ = ~new_G4941_ & ~new_G5001_;
  assign new_G5058_ = ~new_G5001_ & ~new_G4880_;
  assign new_G5059_ = ~new_G4944_ & ~new_G5005_;
  assign new_G5060_ = ~new_G5005_ & ~new_G4885_;
  assign new_G5061_ = ~new_G5009_ & ~new_G5010_;
  assign new_G5064_ = ~new_G5011_ & ~new_G818_;
  assign new_G5068_ = ~new_G4953_ & ~new_G5014_;
  assign new_G5069_ = ~new_G5014_ & ~new_G866_;
  assign new_G5070_ = ~new_G4834_ & ~new_G5014_;
  assign new_G5073_ = ~new_G5018_ & ~new_G5019_;
  assign new_G5076_ = ~new_G5023_ & ~new_G5020_;
  assign new_G5080_ = ~new_G4965_ & ~new_G5026_;
  assign new_G5081_ = ~new_G5026_ & ~new_G4962_;
  assign new_G5082_ = ~new_G5030_ & ~new_G5031_;
  assign new_G5085_ = ~new_G5032_ & ~new_G1061_;
  assign new_G5089_ = ~new_G4974_ & ~new_G5035_;
  assign new_G5090_ = ~new_G5035_ & ~new_G1109_;
  assign new_G5091_ = ~new_G4855_ & ~new_G5035_;
  assign new_G5094_ = ~new_G5039_ & ~new_G5040_;
  assign new_G5097_ = ~new_G5044_ & ~new_G5041_;
  assign new_G5101_ = ~new_G4986_ & ~new_G5047_;
  assign new_G5102_ = ~new_G5047_ & ~new_G4983_;
  assign new_G5103_ = ~new_G5051_ & ~new_G5052_;
  assign new_G5106_ = ~new_G5053_ & ~new_G5054_;
  assign new_G5109_ = ~new_G5055_ & ~new_G5056_;
  assign new_G5112_ = ~new_G5057_ & ~new_G5058_;
  assign new_G5115_ = ~new_G5059_ & ~new_G5060_;
  assign new_G5118_ = ~new_G5061_ & ~new_G770_;
  assign new_G5122_ = ~new_G5011_ & ~new_G5064_;
  assign new_G5123_ = ~new_G5064_ & ~new_G818_;
  assign new_G5124_ = ~new_G4896_ & ~new_G5064_;
  assign new_G5127_ = ~new_G5068_ & ~new_G5069_;
  assign new_G5130_ = ~new_G5073_ & ~new_G5070_;
  assign new_G5134_ = ~new_G5023_ & ~new_G5076_;
  assign new_G5135_ = ~new_G5076_ & ~new_G5020_;
  assign new_G5136_ = ~new_G5080_ & ~new_G5081_;
  assign new_G5139_ = ~new_G5082_ & ~new_G1013_;
  assign new_G5143_ = ~new_G5032_ & ~new_G5085_;
  assign new_G5144_ = ~new_G5085_ & ~new_G1061_;
  assign new_G5145_ = ~new_G4917_ & ~new_G5085_;
  assign new_G5148_ = ~new_G5089_ & ~new_G5090_;
  assign new_G5151_ = ~new_G5094_ & ~new_G5091_;
  assign new_G5155_ = ~new_G5044_ & ~new_G5097_;
  assign new_G5156_ = ~new_G5097_ & ~new_G5041_;
  assign new_G5157_ = ~new_G5101_ & ~new_G5102_;
  assign new_G5160_ = ~new_G5103_ & ~new_G1256_;
  assign new_G5164_ = ~new_G5106_ & ~new_G578_;
  assign new_G5168_ = ~new_G5109_ & ~new_G626_;
  assign new_G5172_ = ~new_G5112_ & ~new_G674_;
  assign new_G5176_ = ~new_G5115_ & ~new_G722_;
  assign new_G5180_ = ~new_G5061_ & ~new_G5118_;
  assign new_G5181_ = ~new_G5118_ & ~new_G770_;
  assign new_G5182_ = ~new_G4947_ & ~new_G5118_;
  assign new_G5185_ = ~new_G5122_ & ~new_G5123_;
  assign new_G5188_ = ~new_G5127_ & ~new_G5124_;
  assign new_G5192_ = ~new_G5073_ & ~new_G5130_;
  assign new_G5193_ = ~new_G5130_ & ~new_G5070_;
  assign new_G5194_ = ~new_G5134_ & ~new_G5135_;
  assign new_G5197_ = ~new_G5136_ & ~new_G965_;
  assign new_G5201_ = ~new_G5082_ & ~new_G5139_;
  assign new_G5202_ = ~new_G5139_ & ~new_G1013_;
  assign new_G5203_ = ~new_G4968_ & ~new_G5139_;
  assign new_G5206_ = ~new_G5143_ & ~new_G5144_;
  assign new_G5209_ = ~new_G5148_ & ~new_G5145_;
  assign new_G5213_ = ~new_G5094_ & ~new_G5151_;
  assign new_G5214_ = ~new_G5151_ & ~new_G5091_;
  assign new_G5215_ = ~new_G5155_ & ~new_G5156_;
  assign new_G5218_ = ~new_G5157_ & ~new_G1208_;
  assign new_G5222_ = ~new_G5103_ & ~new_G5160_;
  assign new_G5223_ = ~new_G5160_ & ~new_G1256_;
  assign new_G5224_ = ~new_G4989_ & ~new_G5160_;
  assign new_G5227_ = ~new_G5106_ & ~new_G5164_;
  assign new_G5228_ = ~new_G5164_ & ~new_G578_;
  assign new_G5229_ = ~new_G4993_ & ~new_G5164_;
  assign new_G5232_ = ~new_G5109_ & ~new_G5168_;
  assign new_G5233_ = ~new_G5168_ & ~new_G626_;
  assign new_G5234_ = ~new_G4997_ & ~new_G5168_;
  assign new_G5237_ = ~new_G5112_ & ~new_G5172_;
  assign new_G5238_ = ~new_G5172_ & ~new_G674_;
  assign new_G5239_ = ~new_G5001_ & ~new_G5172_;
  assign new_G5242_ = ~new_G5115_ & ~new_G5176_;
  assign new_G5243_ = ~new_G5176_ & ~new_G722_;
  assign new_G5244_ = ~new_G5005_ & ~new_G5176_;
  assign new_G5247_ = ~new_G5180_ & ~new_G5181_;
  assign new_G5250_ = ~new_G5185_ & ~new_G5182_;
  assign new_G5254_ = ~new_G5127_ & ~new_G5188_;
  assign new_G5255_ = ~new_G5188_ & ~new_G5124_;
  assign new_G5256_ = ~new_G5192_ & ~new_G5193_;
  assign new_G5259_ = ~new_G5194_ & ~new_G917_;
  assign new_G5263_ = ~new_G5136_ & ~new_G5197_;
  assign new_G5264_ = ~new_G5197_ & ~new_G965_;
  assign new_G5265_ = ~new_G5026_ & ~new_G5197_;
  assign new_G5268_ = ~new_G5201_ & ~new_G5202_;
  assign new_G5271_ = ~new_G5206_ & ~new_G5203_;
  assign new_G5275_ = ~new_G5148_ & ~new_G5209_;
  assign new_G5276_ = ~new_G5209_ & ~new_G5145_;
  assign new_G5277_ = ~new_G5213_ & ~new_G5214_;
  assign new_G5280_ = ~new_G5215_ & ~new_G1160_;
  assign new_G5284_ = ~new_G5157_ & ~new_G5218_;
  assign new_G5285_ = ~new_G5218_ & ~new_G1208_;
  assign new_G5286_ = ~new_G5047_ & ~new_G5218_;
  assign new_G5289_ = ~new_G5222_ & ~new_G5223_;
  assign new_G5292_ = ~new_G1304_ & ~new_G5224_;
  assign new_G5296_ = ~new_G5232_ & ~new_G5233_;
  assign new_G5299_ = ~new_G5237_ & ~new_G5238_;
  assign new_G5302_ = ~new_G5242_ & ~new_G5243_;
  assign new_G5305_ = ~new_G5247_ & ~new_G5244_;
  assign new_G5309_ = ~new_G5185_ & ~new_G5250_;
  assign new_G5310_ = ~new_G5250_ & ~new_G5182_;
  assign new_G5311_ = ~new_G5254_ & ~new_G5255_;
  assign new_G5314_ = ~new_G5256_ & ~new_G869_;
  assign new_G5318_ = ~new_G5194_ & ~new_G5259_;
  assign new_G5319_ = ~new_G5259_ & ~new_G917_;
  assign new_G5320_ = ~new_G5076_ & ~new_G5259_;
  assign new_G5323_ = ~new_G5263_ & ~new_G5264_;
  assign new_G5326_ = ~new_G5268_ & ~new_G5265_;
  assign new_G5330_ = ~new_G5206_ & ~new_G5271_;
  assign new_G5331_ = ~new_G5271_ & ~new_G5203_;
  assign new_G5332_ = ~new_G5275_ & ~new_G5276_;
  assign new_G5335_ = ~new_G5277_ & ~new_G1112_;
  assign new_G5339_ = ~new_G5215_ & ~new_G5280_;
  assign new_G5340_ = ~new_G5280_ & ~new_G1160_;
  assign new_G5341_ = ~new_G5097_ & ~new_G5280_;
  assign new_G5344_ = ~new_G5284_ & ~new_G5285_;
  assign new_G5347_ = ~new_G5289_ & ~new_G5286_;
  assign new_G5351_ = ~new_G1304_ & ~new_G5292_;
  assign new_G5352_ = ~new_G5292_ & ~new_G5224_;
  assign new_G5353_ = ~new_G5296_ & ~new_G5229_;
  assign new_G5357_ = ~new_G5299_ & ~new_G5234_;
  assign new_G5361_ = ~new_G5302_ & ~new_G5239_;
  assign new_G5365_ = ~new_G5247_ & ~new_G5305_;
  assign new_G5366_ = ~new_G5305_ & ~new_G5244_;
  assign new_G5367_ = ~new_G5309_ & ~new_G5310_;
  assign new_G5370_ = ~new_G5311_ & ~new_G821_;
  assign new_G5374_ = ~new_G5256_ & ~new_G5314_;
  assign new_G5375_ = ~new_G5314_ & ~new_G869_;
  assign new_G5376_ = ~new_G5130_ & ~new_G5314_;
  assign new_G5379_ = ~new_G5318_ & ~new_G5319_;
  assign new_G5382_ = ~new_G5323_ & ~new_G5320_;
  assign new_G5386_ = ~new_G5268_ & ~new_G5326_;
  assign new_G5387_ = ~new_G5326_ & ~new_G5265_;
  assign new_G5388_ = ~new_G5330_ & ~new_G5331_;
  assign new_G5391_ = ~new_G5332_ & ~new_G1064_;
  assign new_G5395_ = ~new_G5277_ & ~new_G5335_;
  assign new_G5396_ = ~new_G5335_ & ~new_G1112_;
  assign new_G5397_ = ~new_G5151_ & ~new_G5335_;
  assign new_G5400_ = ~new_G5339_ & ~new_G5340_;
  assign new_G5403_ = ~new_G5344_ & ~new_G5341_;
  assign new_G5407_ = ~new_G5289_ & ~new_G5347_;
  assign new_G5408_ = ~new_G5347_ & ~new_G5286_;
  assign new_G5409_ = ~new_G5351_ & ~new_G5352_;
  assign new_G5412_ = ~new_G5296_ & ~new_G5353_;
  assign new_G5413_ = ~new_G5353_ & ~new_G5229_;
  assign new_G5414_ = ~new_G5299_ & ~new_G5357_;
  assign new_G5415_ = ~new_G5357_ & ~new_G5234_;
  assign new_G5416_ = ~new_G5302_ & ~new_G5361_;
  assign new_G5417_ = ~new_G5361_ & ~new_G5239_;
  assign new_G5418_ = ~new_G5365_ & ~new_G5366_;
  assign new_G5421_ = ~new_G5367_ & ~new_G773_;
  assign new_G5425_ = ~new_G5311_ & ~new_G5370_;
  assign new_G5426_ = ~new_G5370_ & ~new_G821_;
  assign new_G5427_ = ~new_G5188_ & ~new_G5370_;
  assign new_G5430_ = ~new_G5374_ & ~new_G5375_;
  assign new_G5433_ = ~new_G5379_ & ~new_G5376_;
  assign new_G5437_ = ~new_G5323_ & ~new_G5382_;
  assign new_G5438_ = ~new_G5382_ & ~new_G5320_;
  assign new_G5439_ = ~new_G5386_ & ~new_G5387_;
  assign new_G5442_ = ~new_G5388_ & ~new_G1016_;
  assign new_G5446_ = ~new_G5332_ & ~new_G5391_;
  assign new_G5447_ = ~new_G5391_ & ~new_G1064_;
  assign new_G5448_ = ~new_G5209_ & ~new_G5391_;
  assign new_G5451_ = ~new_G5395_ & ~new_G5396_;
  assign new_G5454_ = ~new_G5400_ & ~new_G5397_;
  assign new_G5458_ = ~new_G5344_ & ~new_G5403_;
  assign new_G5459_ = ~new_G5403_ & ~new_G5341_;
  assign new_G5460_ = ~new_G5407_ & ~new_G5408_;
  assign new_G5463_ = ~new_G5409_ & ~new_G1259_;
  assign new_G5467_ = ~new_G5412_ & ~new_G5413_;
  assign new_G5470_ = ~new_G5414_ & ~new_G5415_;
  assign new_G5473_ = ~new_G5416_ & ~new_G5417_;
  assign new_G5476_ = ~new_G5418_ & ~new_G725_;
  assign new_G5480_ = ~new_G5367_ & ~new_G5421_;
  assign new_G5481_ = ~new_G5421_ & ~new_G773_;
  assign new_G5482_ = ~new_G5250_ & ~new_G5421_;
  assign new_G5485_ = ~new_G5425_ & ~new_G5426_;
  assign new_G5488_ = ~new_G5430_ & ~new_G5427_;
  assign new_G5492_ = ~new_G5379_ & ~new_G5433_;
  assign new_G5493_ = ~new_G5433_ & ~new_G5376_;
  assign new_G5494_ = ~new_G5437_ & ~new_G5438_;
  assign new_G5497_ = ~new_G5439_ & ~new_G968_;
  assign new_G5501_ = ~new_G5388_ & ~new_G5442_;
  assign new_G5502_ = ~new_G5442_ & ~new_G1016_;
  assign new_G5503_ = ~new_G5271_ & ~new_G5442_;
  assign new_G5506_ = ~new_G5446_ & ~new_G5447_;
  assign new_G5509_ = ~new_G5451_ & ~new_G5448_;
  assign new_G5513_ = ~new_G5400_ & ~new_G5454_;
  assign new_G5514_ = ~new_G5454_ & ~new_G5397_;
  assign new_G5515_ = ~new_G5458_ & ~new_G5459_;
  assign new_G5518_ = ~new_G5460_ & ~new_G1211_;
  assign new_G5522_ = ~new_G5409_ & ~new_G5463_;
  assign new_G5523_ = ~new_G5463_ & ~new_G1259_;
  assign new_G5524_ = ~new_G5292_ & ~new_G5463_;
  assign new_G5527_ = ~new_G5467_ & ~new_G581_;
  assign new_G5531_ = ~new_G5470_ & ~new_G629_;
  assign new_G5535_ = ~new_G5473_ & ~new_G677_;
  assign new_G5539_ = ~new_G5418_ & ~new_G5476_;
  assign new_G5540_ = ~new_G5476_ & ~new_G725_;
  assign new_G5541_ = ~new_G5305_ & ~new_G5476_;
  assign new_G5544_ = ~new_G5480_ & ~new_G5481_;
  assign new_G5547_ = ~new_G5485_ & ~new_G5482_;
  assign new_G5551_ = ~new_G5430_ & ~new_G5488_;
  assign new_G5552_ = ~new_G5488_ & ~new_G5427_;
  assign new_G5553_ = ~new_G5492_ & ~new_G5493_;
  assign new_G5556_ = ~new_G5494_ & ~new_G920_;
  assign new_G5560_ = ~new_G5439_ & ~new_G5497_;
  assign new_G5561_ = ~new_G5497_ & ~new_G968_;
  assign new_G5562_ = ~new_G5326_ & ~new_G5497_;
  assign new_G5565_ = ~new_G5501_ & ~new_G5502_;
  assign new_G5568_ = ~new_G5506_ & ~new_G5503_;
  assign new_G5572_ = ~new_G5451_ & ~new_G5509_;
  assign new_G5573_ = ~new_G5509_ & ~new_G5448_;
  assign new_G5574_ = ~new_G5513_ & ~new_G5514_;
  assign new_G5577_ = ~new_G5515_ & ~new_G1163_;
  assign new_G5581_ = ~new_G5460_ & ~new_G5518_;
  assign new_G5582_ = ~new_G5518_ & ~new_G1211_;
  assign new_G5583_ = ~new_G5347_ & ~new_G5518_;
  assign new_G5586_ = ~new_G5522_ & ~new_G5523_;
  assign new_G5589_ = ~new_G1307_ & ~new_G5524_;
  assign new_G5593_ = ~new_G5467_ & ~new_G5527_;
  assign new_G5594_ = ~new_G5527_ & ~new_G581_;
  assign new_G5595_ = ~new_G5353_ & ~new_G5527_;
  assign new_G5598_ = ~new_G5470_ & ~new_G5531_;
  assign new_G5599_ = ~new_G5531_ & ~new_G629_;
  assign new_G5600_ = ~new_G5357_ & ~new_G5531_;
  assign new_G5603_ = ~new_G5473_ & ~new_G5535_;
  assign new_G5604_ = ~new_G5535_ & ~new_G677_;
  assign new_G5605_ = ~new_G5361_ & ~new_G5535_;
  assign new_G5608_ = ~new_G5539_ & ~new_G5540_;
  assign new_G5611_ = ~new_G5544_ & ~new_G5541_;
  assign new_G5615_ = ~new_G5485_ & ~new_G5547_;
  assign new_G5616_ = ~new_G5547_ & ~new_G5482_;
  assign new_G5617_ = ~new_G5551_ & ~new_G5552_;
  assign new_G5620_ = ~new_G5553_ & ~new_G872_;
  assign new_G5624_ = ~new_G5494_ & ~new_G5556_;
  assign new_G5625_ = ~new_G5556_ & ~new_G920_;
  assign new_G5626_ = ~new_G5382_ & ~new_G5556_;
  assign new_G5629_ = ~new_G5560_ & ~new_G5561_;
  assign new_G5632_ = ~new_G5565_ & ~new_G5562_;
  assign new_G5636_ = ~new_G5506_ & ~new_G5568_;
  assign new_G5637_ = ~new_G5568_ & ~new_G5503_;
  assign new_G5638_ = ~new_G5572_ & ~new_G5573_;
  assign new_G5641_ = ~new_G5574_ & ~new_G1115_;
  assign new_G5645_ = ~new_G5515_ & ~new_G5577_;
  assign new_G5646_ = ~new_G5577_ & ~new_G1163_;
  assign new_G5647_ = ~new_G5403_ & ~new_G5577_;
  assign new_G5650_ = ~new_G5581_ & ~new_G5582_;
  assign new_G5653_ = ~new_G5586_ & ~new_G5583_;
  assign new_G5657_ = ~new_G1307_ & ~new_G5589_;
  assign new_G5658_ = ~new_G5589_ & ~new_G5524_;
  assign new_G5659_ = ~new_G5598_ & ~new_G5599_;
  assign new_G5662_ = ~new_G5603_ & ~new_G5604_;
  assign new_G5665_ = ~new_G5608_ & ~new_G5605_;
  assign new_G5669_ = ~new_G5544_ & ~new_G5611_;
  assign new_G5670_ = ~new_G5611_ & ~new_G5541_;
  assign new_G5671_ = ~new_G5615_ & ~new_G5616_;
  assign new_G5674_ = ~new_G5617_ & ~new_G824_;
  assign new_G5678_ = ~new_G5553_ & ~new_G5620_;
  assign new_G5679_ = ~new_G5620_ & ~new_G872_;
  assign new_G5680_ = ~new_G5433_ & ~new_G5620_;
  assign new_G5683_ = ~new_G5624_ & ~new_G5625_;
  assign new_G5686_ = ~new_G5629_ & ~new_G5626_;
  assign new_G5690_ = ~new_G5565_ & ~new_G5632_;
  assign new_G5691_ = ~new_G5632_ & ~new_G5562_;
  assign new_G5692_ = ~new_G5636_ & ~new_G5637_;
  assign new_G5695_ = ~new_G5638_ & ~new_G1067_;
  assign new_G5699_ = ~new_G5574_ & ~new_G5641_;
  assign new_G5700_ = ~new_G5641_ & ~new_G1115_;
  assign new_G5701_ = ~new_G5454_ & ~new_G5641_;
  assign new_G5704_ = ~new_G5645_ & ~new_G5646_;
  assign new_G5707_ = ~new_G5650_ & ~new_G5647_;
  assign new_G5711_ = ~new_G5586_ & ~new_G5653_;
  assign new_G5712_ = ~new_G5653_ & ~new_G5583_;
  assign new_G5713_ = ~new_G5657_ & ~new_G5658_;
  assign new_G5716_ = ~new_G5659_ & ~new_G5595_;
  assign new_G5720_ = ~new_G5662_ & ~new_G5600_;
  assign new_G5724_ = ~new_G5608_ & ~new_G5665_;
  assign new_G5725_ = ~new_G5665_ & ~new_G5605_;
  assign new_G5726_ = ~new_G5669_ & ~new_G5670_;
  assign new_G5729_ = ~new_G5671_ & ~new_G776_;
  assign new_G5733_ = ~new_G5617_ & ~new_G5674_;
  assign new_G5734_ = ~new_G5674_ & ~new_G824_;
  assign new_G5735_ = ~new_G5488_ & ~new_G5674_;
  assign new_G5738_ = ~new_G5678_ & ~new_G5679_;
  assign new_G5741_ = ~new_G5683_ & ~new_G5680_;
  assign new_G5745_ = ~new_G5629_ & ~new_G5686_;
  assign new_G5746_ = ~new_G5686_ & ~new_G5626_;
  assign new_G5747_ = ~new_G5690_ & ~new_G5691_;
  assign new_G5750_ = ~new_G5692_ & ~new_G1019_;
  assign new_G5754_ = ~new_G5638_ & ~new_G5695_;
  assign new_G5755_ = ~new_G5695_ & ~new_G1067_;
  assign new_G5756_ = ~new_G5509_ & ~new_G5695_;
  assign new_G5759_ = ~new_G5699_ & ~new_G5700_;
  assign new_G5762_ = ~new_G5704_ & ~new_G5701_;
  assign new_G5766_ = ~new_G5650_ & ~new_G5707_;
  assign new_G5767_ = ~new_G5707_ & ~new_G5647_;
  assign new_G5768_ = ~new_G5711_ & ~new_G5712_;
  assign new_G5771_ = ~new_G5659_ & ~new_G5716_;
  assign new_G5772_ = ~new_G5716_ & ~new_G5595_;
  assign new_G5773_ = ~new_G5662_ & ~new_G5720_;
  assign new_G5774_ = ~new_G5720_ & ~new_G5600_;
  assign new_G5775_ = ~new_G5724_ & ~new_G5725_;
  assign new_G5778_ = ~new_G5726_ & ~new_G728_;
  assign new_G5782_ = ~new_G5671_ & ~new_G5729_;
  assign new_G5783_ = ~new_G5729_ & ~new_G776_;
  assign new_G5784_ = ~new_G5547_ & ~new_G5729_;
  assign new_G5787_ = ~new_G5733_ & ~new_G5734_;
  assign new_G5790_ = ~new_G5738_ & ~new_G5735_;
  assign new_G5794_ = ~new_G5683_ & ~new_G5741_;
  assign new_G5795_ = ~new_G5741_ & ~new_G5680_;
  assign new_G5796_ = ~new_G5745_ & ~new_G5746_;
  assign new_G5799_ = ~new_G5747_ & ~new_G971_;
  assign new_G5803_ = ~new_G5692_ & ~new_G5750_;
  assign new_G5804_ = ~new_G5750_ & ~new_G1019_;
  assign new_G5805_ = ~new_G5568_ & ~new_G5750_;
  assign new_G5808_ = ~new_G5754_ & ~new_G5755_;
  assign new_G5811_ = ~new_G5759_ & ~new_G5756_;
  assign new_G5815_ = ~new_G5704_ & ~new_G5762_;
  assign new_G5816_ = ~new_G5762_ & ~new_G5701_;
  assign new_G5817_ = ~new_G5766_ & ~new_G5767_;
  assign new_G5820_ = ~new_G5771_ & ~new_G5772_;
  assign new_G5823_ = ~new_G5773_ & ~new_G5774_;
  assign new_G5826_ = ~new_G5775_ & ~new_G680_;
  assign new_G5830_ = ~new_G5726_ & ~new_G5778_;
  assign new_G5831_ = ~new_G5778_ & ~new_G728_;
  assign new_G5832_ = ~new_G5611_ & ~new_G5778_;
  assign new_G5835_ = ~new_G5782_ & ~new_G5783_;
  assign new_G5838_ = ~new_G5787_ & ~new_G5784_;
  assign new_G5842_ = ~new_G5738_ & ~new_G5790_;
  assign new_G5843_ = ~new_G5790_ & ~new_G5735_;
  assign new_G5844_ = ~new_G5794_ & ~new_G5795_;
  assign new_G5847_ = ~new_G5796_ & ~new_G923_;
  assign new_G5851_ = ~new_G5747_ & ~new_G5799_;
  assign new_G5852_ = ~new_G5799_ & ~new_G971_;
  assign new_G5853_ = ~new_G5632_ & ~new_G5799_;
  assign new_G5856_ = ~new_G5803_ & ~new_G5804_;
  assign new_G5859_ = ~new_G5808_ & ~new_G5805_;
  assign new_G5863_ = ~new_G5759_ & ~new_G5811_;
  assign new_G5864_ = ~new_G5811_ & ~new_G5756_;
  assign new_G5865_ = ~new_G5815_ & ~new_G5816_;
  assign new_G5868_ = ~new_G5820_ & ~new_G584_;
  assign new_G5872_ = ~new_G5823_ & ~new_G632_;
  assign new_G5876_ = ~new_G5775_ & ~new_G5826_;
  assign new_G5877_ = ~new_G5826_ & ~new_G680_;
  assign new_G5878_ = ~new_G5665_ & ~new_G5826_;
  assign new_G5881_ = ~new_G5830_ & ~new_G5831_;
  assign new_G5884_ = ~new_G5835_ & ~new_G5832_;
  assign new_G5888_ = ~new_G5787_ & ~new_G5838_;
  assign new_G5889_ = ~new_G5838_ & ~new_G5784_;
  assign new_G5890_ = ~new_G5842_ & ~new_G5843_;
  assign new_G5893_ = ~new_G5844_ & ~new_G875_;
  assign new_G5897_ = ~new_G5796_ & ~new_G5847_;
  assign new_G5898_ = ~new_G5847_ & ~new_G923_;
  assign new_G5899_ = ~new_G5686_ & ~new_G5847_;
  assign new_G5902_ = ~new_G5851_ & ~new_G5852_;
  assign new_G5905_ = ~new_G5856_ & ~new_G5853_;
  assign new_G5909_ = ~new_G5808_ & ~new_G5859_;
  assign new_G5910_ = ~new_G5859_ & ~new_G5805_;
  assign new_G5911_ = ~new_G5863_ & ~new_G5864_;
  assign new_G5914_ = ~new_G5820_ & ~new_G5868_;
  assign new_G5915_ = ~new_G5868_ & ~new_G584_;
  assign new_G5916_ = ~new_G5716_ & ~new_G5868_;
  assign new_G5919_ = ~new_G5823_ & ~new_G5872_;
  assign new_G5920_ = ~new_G5872_ & ~new_G632_;
  assign new_G5921_ = ~new_G5720_ & ~new_G5872_;
  assign new_G5924_ = ~new_G5876_ & ~new_G5877_;
  assign new_G5927_ = ~new_G5881_ & ~new_G5878_;
  assign new_G5931_ = ~new_G5835_ & ~new_G5884_;
  assign new_G5932_ = ~new_G5884_ & ~new_G5832_;
  assign new_G5933_ = ~new_G5888_ & ~new_G5889_;
  assign new_G5936_ = ~new_G5890_ & ~new_G827_;
  assign new_G5940_ = ~new_G5844_ & ~new_G5893_;
  assign new_G5941_ = ~new_G5893_ & ~new_G875_;
  assign new_G5942_ = ~new_G5741_ & ~new_G5893_;
  assign new_G5945_ = ~new_G5897_ & ~new_G5898_;
  assign new_G5948_ = ~new_G5902_ & ~new_G5899_;
  assign new_G5952_ = ~new_G5856_ & ~new_G5905_;
  assign new_G5953_ = ~new_G5905_ & ~new_G5853_;
  assign new_G5954_ = ~new_G5909_ & ~new_G5910_;
  assign new_G5957_ = ~new_G5919_ & ~new_G5920_;
  assign new_G5960_ = ~new_G5924_ & ~new_G5921_;
  assign new_G5964_ = ~new_G5881_ & ~new_G5927_;
  assign new_G5965_ = ~new_G5927_ & ~new_G5878_;
  assign new_G5966_ = ~new_G5931_ & ~new_G5932_;
  assign new_G5969_ = ~new_G5933_ & ~new_G779_;
  assign new_G5973_ = ~new_G5890_ & ~new_G5936_;
  assign new_G5974_ = ~new_G5936_ & ~new_G827_;
  assign new_G5975_ = ~new_G5790_ & ~new_G5936_;
  assign new_G5978_ = ~new_G5940_ & ~new_G5941_;
  assign new_G5981_ = ~new_G5945_ & ~new_G5942_;
  assign new_G5985_ = ~new_G5902_ & ~new_G5948_;
  assign new_G5986_ = ~new_G5948_ & ~new_G5899_;
  assign new_G5987_ = ~new_G5952_ & ~new_G5953_;
  assign new_G5990_ = ~new_G5957_ & ~new_G5916_;
  assign new_G5994_ = ~new_G5924_ & ~new_G5960_;
  assign new_G5995_ = ~new_G5960_ & ~new_G5921_;
  assign new_G5996_ = ~new_G5964_ & ~new_G5965_;
  assign new_G5999_ = ~new_G5966_ & ~new_G731_;
  assign new_G6003_ = ~new_G5933_ & ~new_G5969_;
  assign new_G6004_ = ~new_G5969_ & ~new_G779_;
  assign new_G6005_ = ~new_G5838_ & ~new_G5969_;
  assign new_G6008_ = ~new_G5973_ & ~new_G5974_;
  assign new_G6011_ = ~new_G5978_ & ~new_G5975_;
  assign new_G6015_ = ~new_G5945_ & ~new_G5981_;
  assign new_G6016_ = ~new_G5981_ & ~new_G5942_;
  assign new_G6017_ = ~new_G5985_ & ~new_G5986_;
  assign new_G6020_ = ~new_G5957_ & ~new_G5990_;
  assign new_G6021_ = ~new_G5990_ & ~new_G5916_;
  assign new_G6022_ = ~new_G5994_ & ~new_G5995_;
  assign new_G6025_ = ~new_G5996_ & ~new_G683_;
  assign new_G6029_ = ~new_G5966_ & ~new_G5999_;
  assign new_G6030_ = ~new_G5999_ & ~new_G731_;
  assign new_G6031_ = ~new_G5884_ & ~new_G5999_;
  assign new_G6034_ = ~new_G6003_ & ~new_G6004_;
  assign new_G6037_ = ~new_G6008_ & ~new_G6005_;
  assign new_G6041_ = ~new_G5978_ & ~new_G6011_;
  assign new_G6042_ = ~new_G6011_ & ~new_G5975_;
  assign new_G6043_ = ~new_G6015_ & ~new_G6016_;
  assign new_G6046_ = ~new_G6020_ & ~new_G6021_;
  assign new_G6049_ = ~new_G6022_ & ~new_G635_;
  assign new_G6053_ = ~new_G5996_ & ~new_G6025_;
  assign new_G6054_ = ~new_G6025_ & ~new_G683_;
  assign new_G6055_ = ~new_G5927_ & ~new_G6025_;
  assign new_G6058_ = ~new_G6029_ & ~new_G6030_;
  assign new_G6061_ = ~new_G6034_ & ~new_G6031_;
  assign new_G6065_ = ~new_G6008_ & ~new_G6037_;
  assign new_G6066_ = ~new_G6037_ & ~new_G6005_;
  assign new_G6067_ = ~new_G6041_ & ~new_G6042_;
  assign new_G6070_ = ~new_G6046_ & ~new_G587_;
  assign new_G6074_ = ~new_G6022_ & ~new_G6049_;
  assign new_G6075_ = ~new_G6049_ & ~new_G635_;
  assign new_G6076_ = ~new_G5960_ & ~new_G6049_;
  assign new_G6079_ = ~new_G6053_ & ~new_G6054_;
  assign new_G6082_ = ~new_G6058_ & ~new_G6055_;
  assign new_G6086_ = ~new_G6034_ & ~new_G6061_;
  assign new_G6087_ = ~new_G6061_ & ~new_G6031_;
  assign new_G6088_ = ~new_G6065_ & ~new_G6066_;
  assign new_G6091_ = ~new_G6046_ & ~new_G6070_;
  assign new_G6092_ = ~new_G6070_ & ~new_G587_;
  assign new_G6093_ = ~new_G5990_ & ~new_G6070_;
  assign new_G6096_ = ~new_G6074_ & ~new_G6075_;
  assign new_G6099_ = ~new_G6079_ & ~new_G6076_;
  assign new_G6103_ = ~new_G6058_ & ~new_G6082_;
  assign new_G6104_ = ~new_G6082_ & ~new_G6055_;
  assign new_G6105_ = ~new_G6086_ & ~new_G6087_;
  assign new_G6108_ = ~new_G6096_ & ~new_G6093_;
  assign new_G6112_ = ~new_G6079_ & ~new_G6099_;
  assign new_G6113_ = ~new_G6099_ & ~new_G6076_;
  assign new_G6114_ = ~new_G6103_ & ~new_G6104_;
  assign new_G6117_ = ~new_G6096_ & ~new_G6108_;
  assign new_G6118_ = ~new_G6108_ & ~new_G6093_;
  assign new_G6119_ = ~new_G6112_ & ~new_G6113_;
  assign new_G6122_ = ~new_G6117_ & ~new_G6118_;
  assign new_G6125_ = ~new_G6122_;
  assign new_G6129_ = ~new_G6122_ & ~new_G6125_;
  assign new_G6130_ = ~new_G6125_;
  assign new_G6131_ = ~new_G6108_ & ~new_G6125_;
  assign new_G6134_ = ~new_G6119_ & ~new_G6131_;
  assign new_G6138_ = ~new_G6119_ & ~new_G6134_;
  assign new_G6139_ = ~new_G6134_ & ~new_G6131_;
  assign new_G6140_ = ~new_G6099_ & ~new_G6134_;
  assign new_G6143_ = ~new_G6114_ & ~new_G6140_;
  assign new_G6147_ = ~new_G6114_ & ~new_G6143_;
  assign new_G6148_ = ~new_G6143_ & ~new_G6140_;
  assign new_G6149_ = ~new_G6082_ & ~new_G6143_;
  assign new_G6152_ = ~new_G6105_ & ~new_G6149_;
  assign new_G6156_ = ~new_G6105_ & ~new_G6152_;
  assign new_G6157_ = ~new_G6152_ & ~new_G6149_;
  assign new_G6158_ = ~new_G6061_ & ~new_G6152_;
  assign new_G6161_ = ~new_G6088_ & ~new_G6158_;
  assign new_G6165_ = ~new_G6088_ & ~new_G6161_;
  assign new_G6166_ = ~new_G6161_ & ~new_G6158_;
  assign new_G6167_ = ~new_G6037_ & ~new_G6161_;
  assign new_G6170_ = ~new_G6067_ & ~new_G6167_;
  assign new_G6174_ = ~new_G6067_ & ~new_G6170_;
  assign new_G6175_ = ~new_G6170_ & ~new_G6167_;
  assign new_G6176_ = ~new_G6011_ & ~new_G6170_;
  assign new_G6179_ = ~new_G6043_ & ~new_G6176_;
  assign new_G6183_ = ~new_G6043_ & ~new_G6179_;
  assign new_G6184_ = ~new_G6179_ & ~new_G6176_;
  assign new_G6185_ = ~new_G5981_ & ~new_G6179_;
  assign new_G6188_ = ~new_G6017_ & ~new_G6185_;
  assign new_G6192_ = ~new_G6017_ & ~new_G6188_;
  assign new_G6193_ = ~new_G6188_ & ~new_G6185_;
  assign new_G6194_ = ~new_G5948_ & ~new_G6188_;
  assign new_G6197_ = ~new_G5987_ & ~new_G6194_;
  assign new_G6201_ = ~new_G5987_ & ~new_G6197_;
  assign new_G6202_ = ~new_G6197_ & ~new_G6194_;
  assign new_G6203_ = ~new_G5905_ & ~new_G6197_;
  assign new_G6206_ = ~new_G5954_ & ~new_G6203_;
  assign new_G6210_ = ~new_G5954_ & ~new_G6206_;
  assign new_G6211_ = ~new_G6206_ & ~new_G6203_;
  assign new_G6212_ = ~new_G5859_ & ~new_G6206_;
  assign new_G6215_ = ~new_G5911_ & ~new_G6212_;
  assign new_G6219_ = ~new_G5911_ & ~new_G6215_;
  assign new_G6220_ = ~new_G6215_ & ~new_G6212_;
  assign new_G6221_ = ~new_G5811_ & ~new_G6215_;
  assign new_G6224_ = ~new_G5865_ & ~new_G6221_;
  assign new_G6228_ = ~new_G5865_ & ~new_G6224_;
  assign new_G6229_ = ~new_G6224_ & ~new_G6221_;
  assign new_G6230_ = ~new_G5762_ & ~new_G6224_;
  assign new_G6233_ = ~new_G5817_ & ~new_G6230_;
  assign new_G6237_ = ~new_G5817_ & ~new_G6233_;
  assign new_G6238_ = ~new_G6233_ & ~new_G6230_;
  assign new_G6239_ = ~new_G5707_ & ~new_G6233_;
  assign new_G6242_ = ~new_G5768_ & ~new_G6239_;
  assign new_G6246_ = ~new_G5768_ & ~new_G6242_;
  assign new_G6247_ = ~new_G6242_ & ~new_G6239_;
  assign new_G6248_ = ~new_G5653_ & ~new_G6242_;
  assign new_G6251_ = ~new_G5713_ & ~new_G6248_;
  assign new_G6255_ = ~new_G5713_ & ~new_G6251_;
  assign new_G6256_ = ~new_G6251_ & ~new_G6248_;
  assign G6257 = n2491_lo & n2683_lo;
  assign G6258 = ~new_G1505_ & ~new_G1506_;
  assign G6259 = ~new_G1822_ & ~new_G1823_;
  assign G6260 = ~new_G2146_ & ~new_G2147_;
  assign G6261 = ~new_G2472_ & ~new_G2473_;
  assign G6262 = ~new_G2801_ & ~new_G2802_;
  assign G6263 = ~new_G3134_ & ~new_G3135_;
  assign G6264 = ~new_G3472_ & ~new_G3473_;
  assign G6265 = ~new_G3817_ & ~new_G3818_;
  assign G6266 = ~new_G4164_ & ~new_G4165_;
  assign G6267 = ~new_G4514_ & ~new_G4515_;
  assign G6268 = ~new_G4868_ & ~new_G4869_;
  assign G6269 = ~new_G5227_ & ~new_G5228_;
  assign G6270 = ~new_G5593_ & ~new_G5594_;
  assign G6271 = ~new_G5914_ & ~new_G5915_;
  assign G6272 = ~new_G6091_ & ~new_G6092_;
  assign G6273 = ~new_G6129_ & ~new_G6130_;
  assign G6274 = ~new_G6138_ & ~new_G6139_;
  assign G6275 = ~new_G6147_ & ~new_G6148_;
  assign G6276 = ~new_G6156_ & ~new_G6157_;
  assign G6277 = ~new_G6165_ & ~new_G6166_;
  assign G6278 = ~new_G6174_ & ~new_G6175_;
  assign G6279 = ~new_G6183_ & ~new_G6184_;
  assign G6280 = ~new_G6192_ & ~new_G6193_;
  assign G6281 = ~new_G6201_ & ~new_G6202_;
  assign G6282 = ~new_G6210_ & ~new_G6211_;
  assign G6283 = ~new_G6219_ & ~new_G6220_;
  assign G6284 = ~new_G6228_ & ~new_G6229_;
  assign G6285 = ~new_G6237_ & ~new_G6238_;
  assign G6286 = ~new_G6246_ & ~new_G6247_;
  assign G6287 = ~new_G5589_ & ~new_G6251_;
  assign G6288 = ~new_G6255_ & ~new_G6256_;
  assign n2482_li = G1;
  assign n2485_li = n2482_lo;
  assign n2488_li = n2485_lo;
  assign n2491_li = n2488_lo;
  assign n2494_li = G2;
  assign n2497_li = n2494_lo;
  assign n2500_li = n2497_lo;
  assign n2503_li = n2500_lo;
  assign n2506_li = G3;
  assign n2509_li = n2506_lo;
  assign n2512_li = n2509_lo;
  assign n2515_li = n2512_lo;
  assign n2518_li = G4;
  assign n2521_li = n2518_lo;
  assign n2524_li = n2521_lo;
  assign n2527_li = n2524_lo;
  assign n2530_li = G5;
  assign n2533_li = n2530_lo;
  assign n2536_li = n2533_lo;
  assign n2539_li = n2536_lo;
  assign n2542_li = G6;
  assign n2545_li = n2542_lo;
  assign n2548_li = n2545_lo;
  assign n2551_li = n2548_lo;
  assign n2554_li = G7;
  assign n2557_li = n2554_lo;
  assign n2560_li = n2557_lo;
  assign n2563_li = n2560_lo;
  assign n2566_li = G8;
  assign n2569_li = n2566_lo;
  assign n2572_li = n2569_lo;
  assign n2575_li = n2572_lo;
  assign n2578_li = G9;
  assign n2581_li = n2578_lo;
  assign n2584_li = n2581_lo;
  assign n2587_li = n2584_lo;
  assign n2590_li = G10;
  assign n2593_li = n2590_lo;
  assign n2596_li = n2593_lo;
  assign n2599_li = n2596_lo;
  assign n2602_li = G11;
  assign n2605_li = n2602_lo;
  assign n2608_li = n2605_lo;
  assign n2611_li = n2608_lo;
  assign n2614_li = G12;
  assign n2617_li = n2614_lo;
  assign n2620_li = n2617_lo;
  assign n2623_li = n2620_lo;
  assign n2626_li = G13;
  assign n2629_li = n2626_lo;
  assign n2632_li = n2629_lo;
  assign n2635_li = n2632_lo;
  assign n2638_li = G14;
  assign n2641_li = n2638_lo;
  assign n2644_li = n2641_lo;
  assign n2647_li = n2644_lo;
  assign n2650_li = G15;
  assign n2653_li = n2650_lo;
  assign n2656_li = n2653_lo;
  assign n2659_li = n2656_lo;
  assign n2662_li = G16;
  assign n2665_li = n2662_lo;
  assign n2668_li = n2665_lo;
  assign n2671_li = n2668_lo;
  assign n2674_li = G17;
  assign n2677_li = n2674_lo;
  assign n2680_li = n2677_lo;
  assign n2683_li = n2680_lo;
  assign n2686_li = G18;
  assign n2689_li = n2686_lo;
  assign n2692_li = n2689_lo;
  assign n2695_li = n2692_lo;
  assign n2698_li = G19;
  assign n2701_li = n2698_lo;
  assign n2704_li = n2701_lo;
  assign n2707_li = n2704_lo;
  assign n2710_li = G20;
  assign n2713_li = n2710_lo;
  assign n2716_li = n2713_lo;
  assign n2719_li = n2716_lo;
  assign n2722_li = G21;
  assign n2725_li = n2722_lo;
  assign n2728_li = n2725_lo;
  assign n2731_li = n2728_lo;
  assign n2734_li = G22;
  assign n2737_li = n2734_lo;
  assign n2740_li = n2737_lo;
  assign n2743_li = n2740_lo;
  assign n2746_li = G23;
  assign n2749_li = n2746_lo;
  assign n2752_li = n2749_lo;
  assign n2755_li = n2752_lo;
  assign n2758_li = G24;
  assign n2761_li = n2758_lo;
  assign n2764_li = n2761_lo;
  assign n2767_li = n2764_lo;
  assign n2770_li = G25;
  assign n2773_li = n2770_lo;
  assign n2776_li = n2773_lo;
  assign n2779_li = n2776_lo;
  assign n2782_li = G26;
  assign n2785_li = n2782_lo;
  assign n2788_li = n2785_lo;
  assign n2791_li = n2788_lo;
  assign n2794_li = G27;
  assign n2797_li = n2794_lo;
  assign n2800_li = n2797_lo;
  assign n2803_li = n2800_lo;
  assign n2806_li = G28;
  assign n2809_li = n2806_lo;
  assign n2812_li = n2809_lo;
  assign n2815_li = n2812_lo;
  assign n2818_li = G29;
  assign n2821_li = n2818_lo;
  assign n2824_li = n2821_lo;
  assign n2827_li = n2824_lo;
  assign n2830_li = G30;
  assign n2833_li = n2830_lo;
  assign n2836_li = n2833_lo;
  assign n2839_li = n2836_lo;
  assign n2842_li = G31;
  assign n2845_li = n2842_lo;
  assign n2848_li = n2845_lo;
  assign n2851_li = n2848_lo;
  assign n2854_li = G32;
  assign n2857_li = n2854_lo;
  assign n2860_li = n2857_lo;
  assign n2863_li = n2860_lo;
  always @ (posedge clk) begin
    n2482_lo <= n2482_li;
    n2485_lo <= n2485_li;
    n2488_lo <= n2488_li;
    n2491_lo <= n2491_li;
    n2494_lo <= n2494_li;
    n2497_lo <= n2497_li;
    n2500_lo <= n2500_li;
    n2503_lo <= n2503_li;
    n2506_lo <= n2506_li;
    n2509_lo <= n2509_li;
    n2512_lo <= n2512_li;
    n2515_lo <= n2515_li;
    n2518_lo <= n2518_li;
    n2521_lo <= n2521_li;
    n2524_lo <= n2524_li;
    n2527_lo <= n2527_li;
    n2530_lo <= n2530_li;
    n2533_lo <= n2533_li;
    n2536_lo <= n2536_li;
    n2539_lo <= n2539_li;
    n2542_lo <= n2542_li;
    n2545_lo <= n2545_li;
    n2548_lo <= n2548_li;
    n2551_lo <= n2551_li;
    n2554_lo <= n2554_li;
    n2557_lo <= n2557_li;
    n2560_lo <= n2560_li;
    n2563_lo <= n2563_li;
    n2566_lo <= n2566_li;
    n2569_lo <= n2569_li;
    n2572_lo <= n2572_li;
    n2575_lo <= n2575_li;
    n2578_lo <= n2578_li;
    n2581_lo <= n2581_li;
    n2584_lo <= n2584_li;
    n2587_lo <= n2587_li;
    n2590_lo <= n2590_li;
    n2593_lo <= n2593_li;
    n2596_lo <= n2596_li;
    n2599_lo <= n2599_li;
    n2602_lo <= n2602_li;
    n2605_lo <= n2605_li;
    n2608_lo <= n2608_li;
    n2611_lo <= n2611_li;
    n2614_lo <= n2614_li;
    n2617_lo <= n2617_li;
    n2620_lo <= n2620_li;
    n2623_lo <= n2623_li;
    n2626_lo <= n2626_li;
    n2629_lo <= n2629_li;
    n2632_lo <= n2632_li;
    n2635_lo <= n2635_li;
    n2638_lo <= n2638_li;
    n2641_lo <= n2641_li;
    n2644_lo <= n2644_li;
    n2647_lo <= n2647_li;
    n2650_lo <= n2650_li;
    n2653_lo <= n2653_li;
    n2656_lo <= n2656_li;
    n2659_lo <= n2659_li;
    n2662_lo <= n2662_li;
    n2665_lo <= n2665_li;
    n2668_lo <= n2668_li;
    n2671_lo <= n2671_li;
    n2674_lo <= n2674_li;
    n2677_lo <= n2677_li;
    n2680_lo <= n2680_li;
    n2683_lo <= n2683_li;
    n2686_lo <= n2686_li;
    n2689_lo <= n2689_li;
    n2692_lo <= n2692_li;
    n2695_lo <= n2695_li;
    n2698_lo <= n2698_li;
    n2701_lo <= n2701_li;
    n2704_lo <= n2704_li;
    n2707_lo <= n2707_li;
    n2710_lo <= n2710_li;
    n2713_lo <= n2713_li;
    n2716_lo <= n2716_li;
    n2719_lo <= n2719_li;
    n2722_lo <= n2722_li;
    n2725_lo <= n2725_li;
    n2728_lo <= n2728_li;
    n2731_lo <= n2731_li;
    n2734_lo <= n2734_li;
    n2737_lo <= n2737_li;
    n2740_lo <= n2740_li;
    n2743_lo <= n2743_li;
    n2746_lo <= n2746_li;
    n2749_lo <= n2749_li;
    n2752_lo <= n2752_li;
    n2755_lo <= n2755_li;
    n2758_lo <= n2758_li;
    n2761_lo <= n2761_li;
    n2764_lo <= n2764_li;
    n2767_lo <= n2767_li;
    n2770_lo <= n2770_li;
    n2773_lo <= n2773_li;
    n2776_lo <= n2776_li;
    n2779_lo <= n2779_li;
    n2782_lo <= n2782_li;
    n2785_lo <= n2785_li;
    n2788_lo <= n2788_li;
    n2791_lo <= n2791_li;
    n2794_lo <= n2794_li;
    n2797_lo <= n2797_li;
    n2800_lo <= n2800_li;
    n2803_lo <= n2803_li;
    n2806_lo <= n2806_li;
    n2809_lo <= n2809_li;
    n2812_lo <= n2812_li;
    n2815_lo <= n2815_li;
    n2818_lo <= n2818_li;
    n2821_lo <= n2821_li;
    n2824_lo <= n2824_li;
    n2827_lo <= n2827_li;
    n2830_lo <= n2830_li;
    n2833_lo <= n2833_li;
    n2836_lo <= n2836_li;
    n2839_lo <= n2839_li;
    n2842_lo <= n2842_li;
    n2845_lo <= n2845_li;
    n2848_lo <= n2848_li;
    n2851_lo <= n2851_li;
    n2854_lo <= n2854_li;
    n2857_lo <= n2857_li;
    n2860_lo <= n2860_li;
    n2863_lo <= n2863_li;
  end
  initial begin
    n2482_lo <= 1'b0;
    n2485_lo <= 1'b0;
    n2488_lo <= 1'b0;
    n2491_lo <= 1'b0;
    n2494_lo <= 1'b0;
    n2497_lo <= 1'b0;
    n2500_lo <= 1'b0;
    n2503_lo <= 1'b0;
    n2506_lo <= 1'b0;
    n2509_lo <= 1'b0;
    n2512_lo <= 1'b0;
    n2515_lo <= 1'b0;
    n2518_lo <= 1'b0;
    n2521_lo <= 1'b0;
    n2524_lo <= 1'b0;
    n2527_lo <= 1'b0;
    n2530_lo <= 1'b0;
    n2533_lo <= 1'b0;
    n2536_lo <= 1'b0;
    n2539_lo <= 1'b0;
    n2542_lo <= 1'b0;
    n2545_lo <= 1'b0;
    n2548_lo <= 1'b0;
    n2551_lo <= 1'b0;
    n2554_lo <= 1'b0;
    n2557_lo <= 1'b0;
    n2560_lo <= 1'b0;
    n2563_lo <= 1'b0;
    n2566_lo <= 1'b0;
    n2569_lo <= 1'b0;
    n2572_lo <= 1'b0;
    n2575_lo <= 1'b0;
    n2578_lo <= 1'b0;
    n2581_lo <= 1'b0;
    n2584_lo <= 1'b0;
    n2587_lo <= 1'b0;
    n2590_lo <= 1'b0;
    n2593_lo <= 1'b0;
    n2596_lo <= 1'b0;
    n2599_lo <= 1'b0;
    n2602_lo <= 1'b0;
    n2605_lo <= 1'b0;
    n2608_lo <= 1'b0;
    n2611_lo <= 1'b0;
    n2614_lo <= 1'b0;
    n2617_lo <= 1'b0;
    n2620_lo <= 1'b0;
    n2623_lo <= 1'b0;
    n2626_lo <= 1'b0;
    n2629_lo <= 1'b0;
    n2632_lo <= 1'b0;
    n2635_lo <= 1'b0;
    n2638_lo <= 1'b0;
    n2641_lo <= 1'b0;
    n2644_lo <= 1'b0;
    n2647_lo <= 1'b0;
    n2650_lo <= 1'b0;
    n2653_lo <= 1'b0;
    n2656_lo <= 1'b0;
    n2659_lo <= 1'b0;
    n2662_lo <= 1'b0;
    n2665_lo <= 1'b0;
    n2668_lo <= 1'b0;
    n2671_lo <= 1'b0;
    n2674_lo <= 1'b0;
    n2677_lo <= 1'b0;
    n2680_lo <= 1'b0;
    n2683_lo <= 1'b0;
    n2686_lo <= 1'b0;
    n2689_lo <= 1'b0;
    n2692_lo <= 1'b0;
    n2695_lo <= 1'b0;
    n2698_lo <= 1'b0;
    n2701_lo <= 1'b0;
    n2704_lo <= 1'b0;
    n2707_lo <= 1'b0;
    n2710_lo <= 1'b0;
    n2713_lo <= 1'b0;
    n2716_lo <= 1'b0;
    n2719_lo <= 1'b0;
    n2722_lo <= 1'b0;
    n2725_lo <= 1'b0;
    n2728_lo <= 1'b0;
    n2731_lo <= 1'b0;
    n2734_lo <= 1'b0;
    n2737_lo <= 1'b0;
    n2740_lo <= 1'b0;
    n2743_lo <= 1'b0;
    n2746_lo <= 1'b0;
    n2749_lo <= 1'b0;
    n2752_lo <= 1'b0;
    n2755_lo <= 1'b0;
    n2758_lo <= 1'b0;
    n2761_lo <= 1'b0;
    n2764_lo <= 1'b0;
    n2767_lo <= 1'b0;
    n2770_lo <= 1'b0;
    n2773_lo <= 1'b0;
    n2776_lo <= 1'b0;
    n2779_lo <= 1'b0;
    n2782_lo <= 1'b0;
    n2785_lo <= 1'b0;
    n2788_lo <= 1'b0;
    n2791_lo <= 1'b0;
    n2794_lo <= 1'b0;
    n2797_lo <= 1'b0;
    n2800_lo <= 1'b0;
    n2803_lo <= 1'b0;
    n2806_lo <= 1'b0;
    n2809_lo <= 1'b0;
    n2812_lo <= 1'b0;
    n2815_lo <= 1'b0;
    n2818_lo <= 1'b0;
    n2821_lo <= 1'b0;
    n2824_lo <= 1'b0;
    n2827_lo <= 1'b0;
    n2830_lo <= 1'b0;
    n2833_lo <= 1'b0;
    n2836_lo <= 1'b0;
    n2839_lo <= 1'b0;
    n2842_lo <= 1'b0;
    n2845_lo <= 1'b0;
    n2848_lo <= 1'b0;
    n2851_lo <= 1'b0;
    n2854_lo <= 1'b0;
    n2857_lo <= 1'b0;
    n2860_lo <= 1'b0;
    n2863_lo <= 1'b0;
  end
endmodule


