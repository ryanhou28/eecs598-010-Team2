
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  G42,
  G43,
  G44,
  G45,
  G46,
  G47,
  G48,
  G49,
  G50,
  G3519,
  G3520,
  G3521,
  G3522,
  G3523,
  G3524,
  G3525,
  G3526,
  G3527,
  G3528,
  G3529,
  G3530,
  G3531,
  G3532,
  G3533,
  G3534,
  G3535,
  G3536,
  G3537,
  G3538,
  G3539,
  G3540
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input G42;input G43;input G44;input G45;input G46;input G47;input G48;input G49;input G50;
  output G3519;output G3520;output G3521;output G3522;output G3523;output G3524;output G3525;output G3526;output G3527;output G3528;output G3529;output G3530;output G3531;output G3532;output G3533;output G3534;output G3535;output G3536;output G3537;output G3538;output G3539;output G3540;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire g51_p;
  wire g51_n;
  wire g52_p;
  wire g52_n;
  wire g53_p;
  wire g53_n;
  wire g54_p;
  wire g54_n;
  wire g55_p;
  wire g55_n;
  wire g56_p;
  wire g56_n;
  wire g57_p;
  wire g57_n;
  wire g58_p;
  wire g58_n;
  wire g59_p;
  wire g59_n;
  wire g60_p;
  wire g60_n;
  wire g61_p;
  wire g61_n;
  wire g62_p;
  wire g62_n;
  wire g63_p;
  wire g63_n;
  wire g64_p;
  wire g64_n;
  wire g65_p;
  wire g65_n;
  wire g66_p;
  wire g66_n;
  wire g67_p;
  wire g67_n;
  wire g68_p;
  wire g68_n;
  wire g69_p;
  wire g69_n;
  wire g70_p;
  wire g70_n;
  wire g71_p;
  wire g71_n;
  wire g72_p;
  wire g72_n;
  wire g73_p;
  wire g73_n;
  wire g74_p;
  wire g74_n;
  wire g75_p;
  wire g75_n;
  wire g76_p;
  wire g76_n;
  wire g77_p;
  wire g77_n;
  wire g78_p;
  wire g78_n;
  wire g79_p;
  wire g79_n;
  wire g80_p;
  wire g80_n;
  wire g81_p;
  wire g81_n;
  wire g82_p;
  wire g82_n;
  wire g83_p;
  wire g83_n;
  wire g84_p;
  wire g84_n;
  wire g85_p;
  wire g85_n;
  wire g86_p;
  wire g86_n;
  wire g87_p;
  wire g87_n;
  wire g88_p;
  wire g88_n;
  wire g89_p;
  wire g89_n;
  wire g90_p;
  wire g90_n;
  wire g91_p;
  wire g91_n;
  wire g92_p;
  wire g92_n;
  wire g93_p;
  wire g93_n;
  wire g94_p;
  wire g94_n;
  wire g95_p;
  wire g95_n;
  wire g96_p;
  wire g96_n;
  wire g97_p;
  wire g97_n;
  wire g98_p;
  wire g98_n;
  wire g99_p;
  wire g99_n;
  wire g100_p;
  wire g100_n;
  wire g101_p;
  wire g101_n;
  wire g102_p;
  wire g102_n;
  wire g103_p;
  wire g103_n;
  wire g104_p;
  wire g104_n;
  wire g105_p;
  wire g105_n;
  wire g106_p;
  wire g106_n;
  wire g107_p;
  wire g107_n;
  wire g108_p;
  wire g108_n;
  wire g109_p;
  wire g109_n;
  wire g110_p;
  wire g110_n;
  wire g111_p;
  wire g111_n;
  wire g112_p;
  wire g112_n;
  wire g113_p;
  wire g113_n;
  wire g114_p;
  wire g114_n;
  wire g115_p;
  wire g115_n;
  wire g116_p;
  wire g116_n;
  wire g117_p;
  wire g117_n;
  wire g118_p;
  wire g118_n;
  wire g119_p;
  wire g119_n;
  wire g120_p;
  wire g120_n;
  wire g121_p;
  wire g121_n;
  wire g122_p;
  wire g122_n;
  wire g123_p;
  wire g123_n;
  wire g124_p;
  wire g124_n;
  wire g125_p;
  wire g125_n;
  wire g126_p;
  wire g126_n;
  wire g127_p;
  wire g127_n;
  wire g128_p;
  wire g128_n;
  wire g129_p;
  wire g129_n;
  wire g130_p;
  wire g130_n;
  wire g131_p;
  wire g131_n;
  wire g132_p;
  wire g132_n;
  wire g133_p;
  wire g133_n;
  wire g134_p;
  wire g134_n;
  wire g135_p;
  wire g135_n;
  wire g136_p;
  wire g136_n;
  wire g137_p;
  wire g137_n;
  wire g138_p;
  wire g138_n;
  wire g139_p;
  wire g139_n;
  wire g140_p;
  wire g140_n;
  wire g141_p;
  wire g141_n;
  wire g142_p;
  wire g142_n;
  wire g143_p;
  wire g143_n;
  wire g144_p;
  wire g144_n;
  wire g145_p;
  wire g145_n;
  wire g146_p;
  wire g146_n;
  wire g147_p;
  wire g147_n;
  wire g148_p;
  wire g148_n;
  wire g149_p;
  wire g149_n;
  wire g150_p;
  wire g150_n;
  wire g151_p;
  wire g151_n;
  wire g152_p;
  wire g152_n;
  wire g153_p;
  wire g153_n;
  wire g154_p;
  wire g154_n;
  wire g155_p;
  wire g155_n;
  wire g156_p;
  wire g156_n;
  wire g157_p;
  wire g157_n;
  wire g158_p;
  wire g158_n;
  wire g159_p;
  wire g159_n;
  wire g160_p;
  wire g160_n;
  wire g161_p;
  wire g161_n;
  wire g162_p;
  wire g162_n;
  wire g163_p;
  wire g163_n;
  wire g164_p;
  wire g164_n;
  wire g165_p;
  wire g165_n;
  wire g166_p;
  wire g166_n;
  wire g167_p;
  wire g167_n;
  wire g168_p;
  wire g168_n;
  wire g169_p;
  wire g169_n;
  wire g170_p;
  wire g170_n;
  wire g171_p;
  wire g171_n;
  wire g172_p;
  wire g172_n;
  wire g173_p;
  wire g173_n;
  wire g174_p;
  wire g174_n;
  wire g175_p;
  wire g175_n;
  wire g176_p;
  wire g176_n;
  wire g177_p;
  wire g177_n;
  wire g178_p;
  wire g178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire g693_p;
  wire g693_n;
  wire g694_p;
  wire g694_n;
  wire g695_p;
  wire g695_n;
  wire g696_p;
  wire g696_n;
  wire g697_p;
  wire g697_n;
  wire g698_p;
  wire g698_n;
  wire g699_p;
  wire g699_n;
  wire g700_p;
  wire g700_n;
  wire g701_p;
  wire g701_n;
  wire g702_p;
  wire g702_n;
  wire g703_p;
  wire g703_n;
  wire g704_p;
  wire g704_n;
  wire g705_p;
  wire g705_n;
  wire g706_p;
  wire g706_n;
  wire g707_p;
  wire g707_n;
  wire g708_p;
  wire g708_n;
  wire g709_p;
  wire g709_n;
  wire g710_p;
  wire g710_n;
  wire g711_p;
  wire g711_n;
  wire g712_p;
  wire g712_n;
  wire g713_p;
  wire g713_n;
  wire g714_p;
  wire g714_n;
  wire g715_p;
  wire g715_n;
  wire g716_p;
  wire g716_n;
  wire g717_p;
  wire g717_n;
  wire g718_p;
  wire g718_n;
  wire g719_p;
  wire g719_n;
  wire g720_p;
  wire g720_n;
  wire g721_p;
  wire g721_n;
  wire g722_p;
  wire g722_n;
  wire g723_p;
  wire g723_n;
  wire g724_p;
  wire g724_n;
  wire g725_p;
  wire g725_n;
  wire g726_p;
  wire g726_n;
  wire g727_p;
  wire g727_n;
  wire g728_p;
  wire g728_n;
  wire g729_p;
  wire g729_n;
  wire g730_p;
  wire g730_n;
  wire g731_p;
  wire g731_n;
  wire g732_p;
  wire g732_n;
  wire g733_p;
  wire g733_n;
  wire g734_p;
  wire g734_n;
  wire g735_p;
  wire g735_n;
  wire g736_p;
  wire g736_n;
  wire g737_p;
  wire g737_n;
  wire g738_p;
  wire g738_n;
  wire g739_p;
  wire g739_n;
  wire g740_p;
  wire g740_n;
  wire g741_p;
  wire g741_n;
  wire g742_p;
  wire g742_n;
  wire g743_p;
  wire g743_n;
  wire g744_p;
  wire g744_n;
  wire g745_p;
  wire g745_n;
  wire g746_p;
  wire g746_n;
  wire g747_p;
  wire g747_n;
  wire g748_p;
  wire g748_n;
  wire g749_p;
  wire g749_n;
  wire g750_p;
  wire g750_n;
  wire g751_p;
  wire g751_n;
  wire g752_p;
  wire g752_n;
  wire g753_p;
  wire g753_n;
  wire g754_p;
  wire g754_n;
  wire g755_p;
  wire g755_n;
  wire g756_p;
  wire g756_n;
  wire g757_p;
  wire g757_n;
  wire g758_p;
  wire g758_n;
  wire g759_p;
  wire g759_n;
  wire g760_p;
  wire g760_n;
  wire g761_p;
  wire g761_n;
  wire g762_p;
  wire g762_n;
  wire g763_p;
  wire g763_n;
  wire g764_p;
  wire g764_n;
  wire g765_p;
  wire g765_n;
  wire g766_p;
  wire g766_n;
  wire g767_p;
  wire g767_n;
  wire g768_p;
  wire g768_n;
  wire g769_p;
  wire g769_n;
  wire g770_p;
  wire g770_n;
  wire g771_p;
  wire g771_n;
  wire g772_p;
  wire g772_n;
  wire g773_p;
  wire g773_n;
  wire g774_p;
  wire g774_n;
  wire g775_p;
  wire g775_n;
  wire g776_p;
  wire g776_n;
  wire g777_p;
  wire g777_n;
  wire g778_p;
  wire g778_n;
  wire g779_p;
  wire g779_n;
  wire g780_p;
  wire g780_n;
  wire g781_p;
  wire g781_n;
  wire g782_p;
  wire g782_n;
  wire g783_p;
  wire g783_n;
  wire g784_p;
  wire g784_n;
  wire g785_p;
  wire g785_n;
  wire g786_p;
  wire g786_n;
  wire g787_p;
  wire g787_n;
  wire g788_p;
  wire g788_n;
  wire g789_p;
  wire g789_n;
  wire g790_p;
  wire g790_n;
  wire g791_p;
  wire g791_n;
  wire g792_p;
  wire g792_n;
  wire g793_p;
  wire g793_n;
  wire g794_p;
  wire g794_n;
  wire g795_p;
  wire g795_n;
  wire g796_p;
  wire g796_n;
  wire g797_p;
  wire g797_n;
  wire g798_p;
  wire g798_n;
  wire g799_p;
  wire g799_n;
  wire g800_p;
  wire g800_n;
  wire g801_p;
  wire g801_n;
  wire g802_p;
  wire g802_n;
  wire g803_p;
  wire g803_n;
  wire g804_p;
  wire g804_n;
  wire g805_p;
  wire g805_n;
  wire g806_p;
  wire g806_n;
  wire g807_p;
  wire g807_n;
  wire g808_p;
  wire g808_n;
  wire g809_p;
  wire g809_n;
  wire g810_p;
  wire g810_n;
  wire g811_p;
  wire g811_n;
  wire g812_p;
  wire g812_n;
  wire g813_p;
  wire g813_n;
  wire g814_p;
  wire g814_n;
  wire g815_p;
  wire g815_n;
  wire g816_p;
  wire g816_n;
  wire g817_p;
  wire g817_n;
  wire g818_p;
  wire g818_n;
  wire g819_p;
  wire g819_n;
  wire g820_p;
  wire g820_n;
  wire g821_p;
  wire g821_n;
  wire g822_p;
  wire g822_n;
  wire g823_p;
  wire g823_n;
  wire g824_p;
  wire g824_n;
  wire g825_p;
  wire g825_n;
  wire g826_p;
  wire g826_n;
  wire g827_p;
  wire g827_n;
  wire g828_p;
  wire g828_n;
  wire g829_p;
  wire g829_n;
  wire g830_p;
  wire g830_n;
  wire g831_p;
  wire g831_n;
  wire g832_p;
  wire g832_n;
  wire g833_p;
  wire g833_n;
  wire g834_p;
  wire g834_n;
  wire g835_p;
  wire g835_n;
  wire g836_p;
  wire g836_n;
  wire g837_p;
  wire g837_n;
  wire g838_p;
  wire g838_n;
  wire g839_p;
  wire g839_n;
  wire g840_p;
  wire g840_n;
  wire g841_p;
  wire g841_n;
  wire g842_p;
  wire g842_n;
  wire g843_p;
  wire g843_n;
  wire g844_p;
  wire g844_n;
  wire g845_p;
  wire g845_n;
  wire g846_p;
  wire g846_n;
  wire g847_p;
  wire g847_n;
  wire g848_p;
  wire g848_n;
  wire g849_p;
  wire g849_n;
  wire g850_p;
  wire g850_n;
  wire g851_p;
  wire g851_n;
  wire g852_p;
  wire g852_n;
  wire g853_p;
  wire g853_n;
  wire g854_p;
  wire g854_n;
  wire g855_p;
  wire g855_n;
  wire g856_p;
  wire g856_n;
  wire g857_p;
  wire g857_n;
  wire g858_p;
  wire g858_n;
  wire g859_p;
  wire g859_n;
  wire g860_p;
  wire g860_n;
  wire g861_p;
  wire g861_n;
  wire g862_p;
  wire g862_n;
  wire g863_p;
  wire g863_n;
  wire g864_p;
  wire g864_n;
  wire g865_p;
  wire g865_n;
  wire g866_p;
  wire g866_n;
  wire g867_p;
  wire g867_n;
  wire g868_p;
  wire g868_n;
  wire g869_p;
  wire g869_n;
  wire g870_p;
  wire g870_n;
  wire g871_p;
  wire g871_n;
  wire g872_p;
  wire g872_n;
  wire g873_p;
  wire g873_n;
  wire g874_p;
  wire g874_n;
  wire g875_p;
  wire g875_n;
  wire g876_p;
  wire g876_n;
  wire g877_p;
  wire g877_n;
  wire g878_p;
  wire g878_n;
  wire g879_p;
  wire g879_n;
  wire g880_p;
  wire g880_n;
  wire g881_p;
  wire g881_n;
  wire g882_p;
  wire g882_n;
  wire g883_p;
  wire g883_n;
  wire g884_p;
  wire g884_n;
  wire g885_p;
  wire g885_n;
  wire g886_p;
  wire g886_n;
  wire g887_p;
  wire g887_n;
  wire g888_p;
  wire g888_n;
  wire g889_p;
  wire g889_n;
  wire g890_p;
  wire g890_n;
  wire g891_p;
  wire g891_n;
  wire g892_p;
  wire g892_n;
  wire g893_p;
  wire g893_n;
  wire g894_p;
  wire g894_n;
  wire g895_p;
  wire g895_n;
  wire g896_p;
  wire g896_n;
  wire g897_p;
  wire g897_n;
  wire g898_p;
  wire g898_n;
  wire g899_p;
  wire g899_n;
  wire g900_p;
  wire g900_n;
  wire g901_p;
  wire g901_n;
  wire g902_p;
  wire g902_n;
  wire g903_p;
  wire g903_n;
  wire g904_p;
  wire g904_n;
  wire G7_n_spl_;
  wire G7_n_spl_0;
  wire G7_n_spl_00;
  wire G7_n_spl_000;
  wire G7_n_spl_0000;
  wire G7_n_spl_001;
  wire G7_n_spl_01;
  wire G7_n_spl_010;
  wire G7_n_spl_011;
  wire G7_n_spl_1;
  wire G7_n_spl_10;
  wire G7_n_spl_100;
  wire G7_n_spl_101;
  wire G7_n_spl_11;
  wire G7_n_spl_110;
  wire G7_n_spl_111;
  wire G8_n_spl_;
  wire G8_n_spl_0;
  wire G8_n_spl_00;
  wire G8_n_spl_000;
  wire G8_n_spl_001;
  wire G8_n_spl_01;
  wire G8_n_spl_010;
  wire G8_n_spl_011;
  wire G8_n_spl_1;
  wire G8_n_spl_10;
  wire G8_n_spl_100;
  wire G8_n_spl_101;
  wire G8_n_spl_11;
  wire G8_n_spl_110;
  wire G7_p_spl_;
  wire G7_p_spl_0;
  wire G7_p_spl_00;
  wire G7_p_spl_000;
  wire G7_p_spl_0000;
  wire G7_p_spl_0001;
  wire G7_p_spl_001;
  wire G7_p_spl_01;
  wire G7_p_spl_010;
  wire G7_p_spl_011;
  wire G7_p_spl_1;
  wire G7_p_spl_10;
  wire G7_p_spl_100;
  wire G7_p_spl_101;
  wire G7_p_spl_11;
  wire G7_p_spl_110;
  wire G7_p_spl_111;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire G8_p_spl_00;
  wire G8_p_spl_000;
  wire G8_p_spl_001;
  wire G8_p_spl_01;
  wire G8_p_spl_010;
  wire G8_p_spl_011;
  wire G8_p_spl_1;
  wire G8_p_spl_10;
  wire G8_p_spl_100;
  wire G8_p_spl_101;
  wire G8_p_spl_11;
  wire G8_p_spl_110;
  wire G8_p_spl_111;
  wire G9_n_spl_;
  wire G9_n_spl_0;
  wire G9_n_spl_00;
  wire G9_n_spl_000;
  wire G9_n_spl_001;
  wire G9_n_spl_01;
  wire G9_n_spl_010;
  wire G9_n_spl_011;
  wire G9_n_spl_1;
  wire G9_n_spl_10;
  wire G9_n_spl_100;
  wire G9_n_spl_101;
  wire G9_n_spl_11;
  wire G9_n_spl_110;
  wire g51_p_spl_;
  wire G9_p_spl_;
  wire G9_p_spl_0;
  wire G9_p_spl_00;
  wire G9_p_spl_000;
  wire G9_p_spl_001;
  wire G9_p_spl_01;
  wire G9_p_spl_010;
  wire G9_p_spl_011;
  wire G9_p_spl_1;
  wire G9_p_spl_10;
  wire G9_p_spl_100;
  wire G9_p_spl_101;
  wire G9_p_spl_11;
  wire G9_p_spl_110;
  wire g51_n_spl_;
  wire G10_n_spl_;
  wire G10_n_spl_0;
  wire G10_n_spl_00;
  wire G10_n_spl_000;
  wire G10_n_spl_001;
  wire G10_n_spl_01;
  wire G10_n_spl_010;
  wire G10_n_spl_011;
  wire G10_n_spl_1;
  wire G10_n_spl_10;
  wire G10_n_spl_100;
  wire G10_n_spl_101;
  wire G10_n_spl_11;
  wire G10_n_spl_110;
  wire g52_p_spl_;
  wire G12_n_spl_;
  wire G12_n_spl_0;
  wire G12_n_spl_00;
  wire G12_n_spl_000;
  wire G12_n_spl_001;
  wire G12_n_spl_01;
  wire G12_n_spl_010;
  wire G12_n_spl_011;
  wire G12_n_spl_1;
  wire G12_n_spl_10;
  wire G12_n_spl_100;
  wire G12_n_spl_101;
  wire G12_n_spl_11;
  wire G13_n_spl_;
  wire G13_n_spl_0;
  wire G13_n_spl_00;
  wire G13_n_spl_000;
  wire G13_n_spl_001;
  wire G13_n_spl_01;
  wire G13_n_spl_010;
  wire G13_n_spl_011;
  wire G13_n_spl_1;
  wire G13_n_spl_10;
  wire G13_n_spl_100;
  wire G13_n_spl_101;
  wire G13_n_spl_11;
  wire G13_n_spl_110;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire G12_p_spl_00;
  wire G12_p_spl_000;
  wire G12_p_spl_001;
  wire G12_p_spl_01;
  wire G12_p_spl_010;
  wire G12_p_spl_011;
  wire G12_p_spl_1;
  wire G12_p_spl_10;
  wire G12_p_spl_100;
  wire G12_p_spl_101;
  wire G12_p_spl_11;
  wire G12_p_spl_110;
  wire G13_p_spl_;
  wire G13_p_spl_0;
  wire G13_p_spl_00;
  wire G13_p_spl_000;
  wire G13_p_spl_001;
  wire G13_p_spl_01;
  wire G13_p_spl_010;
  wire G13_p_spl_011;
  wire G13_p_spl_1;
  wire G13_p_spl_10;
  wire G13_p_spl_100;
  wire G13_p_spl_101;
  wire G13_p_spl_11;
  wire G13_p_spl_110;
  wire G13_p_spl_111;
  wire G11_p_spl_;
  wire G11_p_spl_0;
  wire G11_p_spl_00;
  wire G11_p_spl_000;
  wire G11_p_spl_001;
  wire G11_p_spl_01;
  wire G11_p_spl_010;
  wire G11_p_spl_011;
  wire G11_p_spl_1;
  wire G11_p_spl_10;
  wire G11_p_spl_100;
  wire G11_p_spl_101;
  wire G11_p_spl_11;
  wire g54_n_spl_;
  wire G11_n_spl_;
  wire G11_n_spl_0;
  wire G11_n_spl_00;
  wire G11_n_spl_000;
  wire G11_n_spl_001;
  wire G11_n_spl_01;
  wire G11_n_spl_010;
  wire G11_n_spl_011;
  wire G11_n_spl_1;
  wire G11_n_spl_10;
  wire G11_n_spl_100;
  wire G11_n_spl_11;
  wire g54_p_spl_;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire G1_n_spl_00;
  wire G1_n_spl_000;
  wire G1_n_spl_001;
  wire G1_n_spl_01;
  wire G1_n_spl_010;
  wire G1_n_spl_1;
  wire G1_n_spl_10;
  wire G1_n_spl_11;
  wire G3_n_spl_;
  wire G3_n_spl_0;
  wire G3_n_spl_00;
  wire G3_n_spl_000;
  wire G3_n_spl_0000;
  wire G3_n_spl_0001;
  wire G3_n_spl_001;
  wire G3_n_spl_0010;
  wire G3_n_spl_01;
  wire G3_n_spl_010;
  wire G3_n_spl_011;
  wire G3_n_spl_1;
  wire G3_n_spl_10;
  wire G3_n_spl_100;
  wire G3_n_spl_101;
  wire G3_n_spl_11;
  wire G3_n_spl_110;
  wire G3_n_spl_111;
  wire G34_n_spl_;
  wire G34_n_spl_0;
  wire G34_n_spl_00;
  wire G34_n_spl_01;
  wire G34_n_spl_1;
  wire G34_n_spl_10;
  wire G32_n_spl_;
  wire G32_n_spl_0;
  wire G32_n_spl_00;
  wire G32_n_spl_01;
  wire G32_n_spl_1;
  wire G36_n_spl_;
  wire G36_n_spl_0;
  wire G36_n_spl_00;
  wire G36_n_spl_01;
  wire G36_n_spl_1;
  wire G10_p_spl_;
  wire G10_p_spl_0;
  wire G10_p_spl_00;
  wire G10_p_spl_000;
  wire G10_p_spl_001;
  wire G10_p_spl_01;
  wire G10_p_spl_010;
  wire G10_p_spl_011;
  wire G10_p_spl_1;
  wire G10_p_spl_10;
  wire G10_p_spl_100;
  wire G10_p_spl_101;
  wire G10_p_spl_11;
  wire G33_n_spl_;
  wire G33_n_spl_0;
  wire G33_n_spl_00;
  wire G33_n_spl_01;
  wire G33_n_spl_1;
  wire G14_p_spl_;
  wire G14_p_spl_0;
  wire G14_p_spl_00;
  wire G14_p_spl_000;
  wire G14_p_spl_001;
  wire G14_p_spl_01;
  wire G14_p_spl_010;
  wire G14_p_spl_011;
  wire G14_p_spl_1;
  wire G14_p_spl_10;
  wire G14_p_spl_100;
  wire G14_p_spl_101;
  wire G14_p_spl_11;
  wire G14_p_spl_110;
  wire G14_p_spl_111;
  wire G37_n_spl_;
  wire G37_n_spl_0;
  wire G37_n_spl_1;
  wire G31_n_spl_;
  wire G31_n_spl_0;
  wire G31_n_spl_00;
  wire G31_n_spl_01;
  wire G31_n_spl_1;
  wire G35_n_spl_;
  wire G35_n_spl_0;
  wire G35_n_spl_00;
  wire G35_n_spl_01;
  wire G35_n_spl_1;
  wire G35_n_spl_10;
  wire G30_n_spl_;
  wire G30_n_spl_0;
  wire G30_n_spl_00;
  wire G30_n_spl_01;
  wire G30_n_spl_1;
  wire G2_p_spl_;
  wire G2_p_spl_0;
  wire G2_p_spl_00;
  wire G2_p_spl_1;
  wire G1_p_spl_;
  wire G1_p_spl_0;
  wire G1_p_spl_00;
  wire G1_p_spl_000;
  wire G1_p_spl_01;
  wire G1_p_spl_1;
  wire G1_p_spl_10;
  wire G1_p_spl_11;
  wire G2_n_spl_;
  wire G2_n_spl_0;
  wire G2_n_spl_00;
  wire G2_n_spl_1;
  wire g73_p_spl_;
  wire g73_p_spl_0;
  wire G3_p_spl_;
  wire G3_p_spl_0;
  wire G3_p_spl_00;
  wire G3_p_spl_000;
  wire G3_p_spl_0000;
  wire G3_p_spl_0001;
  wire G3_p_spl_001;
  wire G3_p_spl_01;
  wire G3_p_spl_010;
  wire G3_p_spl_011;
  wire G3_p_spl_1;
  wire G3_p_spl_10;
  wire G3_p_spl_100;
  wire G3_p_spl_101;
  wire G3_p_spl_11;
  wire G3_p_spl_110;
  wire G3_p_spl_111;
  wire g73_n_spl_;
  wire g73_n_spl_0;
  wire g75_n_spl_;
  wire g75_p_spl_;
  wire g74_n_spl_;
  wire g76_n_spl_;
  wire g78_p_spl_;
  wire g78_n_spl_;
  wire g79_n_spl_;
  wire g79_n_spl_0;
  wire g79_n_spl_1;
  wire G36_p_spl_;
  wire G36_p_spl_0;
  wire G36_p_spl_1;
  wire G37_p_spl_;
  wire G37_p_spl_0;
  wire G34_p_spl_;
  wire G34_p_spl_0;
  wire G34_p_spl_00;
  wire G34_p_spl_1;
  wire G35_p_spl_;
  wire G35_p_spl_0;
  wire G35_p_spl_00;
  wire G35_p_spl_1;
  wire g87_p_spl_;
  wire g90_n_spl_;
  wire g87_n_spl_;
  wire g90_p_spl_;
  wire G32_p_spl_;
  wire G32_p_spl_0;
  wire G32_p_spl_00;
  wire G32_p_spl_1;
  wire G33_p_spl_;
  wire G33_p_spl_0;
  wire G33_p_spl_00;
  wire G33_p_spl_1;
  wire G30_p_spl_;
  wire G30_p_spl_0;
  wire G30_p_spl_00;
  wire G30_p_spl_1;
  wire G31_p_spl_;
  wire G31_p_spl_0;
  wire G31_p_spl_00;
  wire G31_p_spl_1;
  wire g96_n_spl_;
  wire g99_p_spl_;
  wire g96_p_spl_;
  wire g99_n_spl_;
  wire g102_p_spl_;
  wire g102_n_spl_;
  wire g106_n_spl_;
  wire g106_p_spl_;
  wire G14_n_spl_;
  wire G14_n_spl_0;
  wire G14_n_spl_00;
  wire G14_n_spl_000;
  wire G14_n_spl_001;
  wire G14_n_spl_01;
  wire G14_n_spl_010;
  wire G14_n_spl_011;
  wire G14_n_spl_1;
  wire G14_n_spl_10;
  wire G14_n_spl_100;
  wire G14_n_spl_101;
  wire G14_n_spl_11;
  wire G14_n_spl_110;
  wire G14_n_spl_111;
  wire g108_p_spl_;
  wire g111_n_spl_;
  wire g108_n_spl_;
  wire g111_p_spl_;
  wire g117_n_spl_;
  wire g117_p_spl_;
  wire g116_p_spl_;
  wire g119_n_spl_;
  wire g116_n_spl_;
  wire g119_p_spl_;
  wire g122_p_spl_;
  wire g122_n_spl_;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_00;
  wire G4_p_spl_000;
  wire G4_p_spl_0000;
  wire G4_p_spl_00000;
  wire G4_p_spl_00001;
  wire G4_p_spl_0001;
  wire G4_p_spl_00010;
  wire G4_p_spl_00011;
  wire G4_p_spl_001;
  wire G4_p_spl_0010;
  wire G4_p_spl_0011;
  wire G4_p_spl_01;
  wire G4_p_spl_010;
  wire G4_p_spl_0100;
  wire G4_p_spl_0101;
  wire G4_p_spl_011;
  wire G4_p_spl_0110;
  wire G4_p_spl_0111;
  wire G4_p_spl_1;
  wire G4_p_spl_10;
  wire G4_p_spl_100;
  wire G4_p_spl_1000;
  wire G4_p_spl_1001;
  wire G4_p_spl_101;
  wire G4_p_spl_1010;
  wire G4_p_spl_1011;
  wire G4_p_spl_11;
  wire G4_p_spl_110;
  wire G4_p_spl_1100;
  wire G4_p_spl_1101;
  wire G4_p_spl_111;
  wire G4_p_spl_1110;
  wire G4_p_spl_1111;
  wire G4_n_spl_;
  wire G4_n_spl_0;
  wire G4_n_spl_00;
  wire G4_n_spl_000;
  wire G4_n_spl_0000;
  wire G4_n_spl_00000;
  wire G4_n_spl_00001;
  wire G4_n_spl_0001;
  wire G4_n_spl_00010;
  wire G4_n_spl_00011;
  wire G4_n_spl_001;
  wire G4_n_spl_0010;
  wire G4_n_spl_0011;
  wire G4_n_spl_01;
  wire G4_n_spl_010;
  wire G4_n_spl_0100;
  wire G4_n_spl_0101;
  wire G4_n_spl_011;
  wire G4_n_spl_0110;
  wire G4_n_spl_0111;
  wire G4_n_spl_1;
  wire G4_n_spl_10;
  wire G4_n_spl_100;
  wire G4_n_spl_1000;
  wire G4_n_spl_1001;
  wire G4_n_spl_101;
  wire G4_n_spl_1010;
  wire G4_n_spl_1011;
  wire G4_n_spl_11;
  wire G4_n_spl_110;
  wire G4_n_spl_1100;
  wire G4_n_spl_1101;
  wire G4_n_spl_111;
  wire G4_n_spl_1110;
  wire G4_n_spl_1111;
  wire g126_n_spl_;
  wire g126_p_spl_;
  wire g129_p_spl_;
  wire g129_p_spl_0;
  wire g129_p_spl_00;
  wire g129_p_spl_000;
  wire g129_p_spl_001;
  wire g129_p_spl_01;
  wire g129_p_spl_1;
  wire g129_p_spl_10;
  wire g129_p_spl_11;
  wire g130_n_spl_;
  wire g130_n_spl_0;
  wire g130_n_spl_00;
  wire g130_n_spl_01;
  wire g130_n_spl_1;
  wire g130_n_spl_10;
  wire g130_n_spl_11;
  wire g129_n_spl_;
  wire g129_n_spl_0;
  wire g129_n_spl_00;
  wire g129_n_spl_000;
  wire g129_n_spl_001;
  wire g129_n_spl_01;
  wire g129_n_spl_1;
  wire g129_n_spl_10;
  wire g129_n_spl_11;
  wire g130_p_spl_;
  wire g130_p_spl_0;
  wire g130_p_spl_00;
  wire g130_p_spl_01;
  wire g130_p_spl_1;
  wire g130_p_spl_10;
  wire g130_p_spl_11;
  wire g131_p_spl_;
  wire g131_n_spl_;
  wire g133_n_spl_;
  wire g133_n_spl_0;
  wire g133_n_spl_1;
  wire g134_n_spl_;
  wire g134_n_spl_0;
  wire g133_p_spl_;
  wire g133_p_spl_0;
  wire g133_p_spl_1;
  wire g134_p_spl_;
  wire g134_p_spl_0;
  wire g137_n_spl_;
  wire g137_n_spl_0;
  wire g137_n_spl_00;
  wire g137_n_spl_000;
  wire g137_n_spl_01;
  wire g137_n_spl_1;
  wire g137_n_spl_10;
  wire g137_n_spl_11;
  wire g137_p_spl_;
  wire g137_p_spl_0;
  wire g137_p_spl_00;
  wire g137_p_spl_000;
  wire g137_p_spl_01;
  wire g137_p_spl_1;
  wire g137_p_spl_10;
  wire g137_p_spl_11;
  wire g138_p_spl_;
  wire g138_p_spl_0;
  wire g138_p_spl_00;
  wire g138_p_spl_01;
  wire g138_p_spl_1;
  wire g138_p_spl_10;
  wire g138_p_spl_11;
  wire g138_n_spl_;
  wire g138_n_spl_0;
  wire g138_n_spl_00;
  wire g138_n_spl_01;
  wire g138_n_spl_1;
  wire g138_n_spl_10;
  wire g138_n_spl_11;
  wire G39_p_spl_;
  wire G39_p_spl_0;
  wire G39_p_spl_00;
  wire G39_p_spl_000;
  wire G39_p_spl_01;
  wire G39_p_spl_1;
  wire G39_p_spl_10;
  wire G39_p_spl_11;
  wire G39_n_spl_;
  wire G39_n_spl_0;
  wire G39_n_spl_00;
  wire G39_n_spl_000;
  wire G39_n_spl_01;
  wire G39_n_spl_1;
  wire G39_n_spl_10;
  wire G39_n_spl_11;
  wire G5_p_spl_;
  wire G5_p_spl_0;
  wire G5_p_spl_00;
  wire G5_p_spl_01;
  wire G5_p_spl_1;
  wire G5_n_spl_;
  wire G5_n_spl_0;
  wire G5_n_spl_00;
  wire G5_n_spl_01;
  wire G5_n_spl_1;
  wire g146_n_spl_;
  wire g146_p_spl_;
  wire g147_n_spl_;
  wire g147_n_spl_0;
  wire g147_n_spl_00;
  wire g147_n_spl_000;
  wire g147_n_spl_01;
  wire g147_n_spl_1;
  wire g147_n_spl_10;
  wire g147_n_spl_11;
  wire g147_p_spl_;
  wire g147_p_spl_0;
  wire g147_p_spl_00;
  wire g147_p_spl_000;
  wire g147_p_spl_01;
  wire g147_p_spl_1;
  wire g147_p_spl_10;
  wire g147_p_spl_11;
  wire G6_n_spl_;
  wire G6_n_spl_0;
  wire G6_n_spl_00;
  wire G6_n_spl_01;
  wire G6_n_spl_1;
  wire G6_n_spl_10;
  wire G6_p_spl_;
  wire G6_p_spl_0;
  wire G6_p_spl_00;
  wire G6_p_spl_01;
  wire G6_p_spl_1;
  wire G6_p_spl_10;
  wire g149_p_spl_;
  wire g149_p_spl_0;
  wire g149_n_spl_;
  wire g149_n_spl_0;
  wire g148_p_spl_;
  wire g148_p_spl_0;
  wire g150_p_spl_;
  wire g150_p_spl_0;
  wire g150_p_spl_1;
  wire g148_n_spl_;
  wire g148_n_spl_0;
  wire g150_n_spl_;
  wire g150_n_spl_0;
  wire g150_n_spl_1;
  wire g153_p_spl_;
  wire g153_p_spl_0;
  wire g153_p_spl_00;
  wire g153_p_spl_01;
  wire g153_p_spl_1;
  wire g153_p_spl_10;
  wire g153_p_spl_11;
  wire g153_n_spl_;
  wire g153_n_spl_0;
  wire g153_n_spl_00;
  wire g153_n_spl_01;
  wire g153_n_spl_1;
  wire g153_n_spl_10;
  wire g153_n_spl_11;
  wire G41_n_spl_;
  wire G41_n_spl_0;
  wire G41_n_spl_00;
  wire G41_n_spl_01;
  wire G41_n_spl_1;
  wire G41_n_spl_10;
  wire G41_p_spl_;
  wire G41_p_spl_0;
  wire G41_p_spl_00;
  wire G41_p_spl_01;
  wire G41_p_spl_1;
  wire G41_p_spl_10;
  wire g151_n_spl_;
  wire g151_n_spl_0;
  wire g151_p_spl_;
  wire g151_p_spl_0;
  wire G25_n_spl_;
  wire G26_n_spl_;
  wire G26_n_spl_0;
  wire G25_p_spl_;
  wire G26_p_spl_;
  wire G26_p_spl_0;
  wire g161_p_spl_;
  wire g161_p_spl_0;
  wire g161_p_spl_1;
  wire g162_n_spl_;
  wire g162_n_spl_0;
  wire g162_n_spl_00;
  wire g162_n_spl_000;
  wire g162_n_spl_01;
  wire g162_n_spl_1;
  wire g162_n_spl_10;
  wire g162_n_spl_11;
  wire g161_n_spl_;
  wire g161_n_spl_0;
  wire g161_n_spl_1;
  wire g162_p_spl_;
  wire g162_p_spl_0;
  wire g162_p_spl_00;
  wire g162_p_spl_000;
  wire g162_p_spl_01;
  wire g162_p_spl_1;
  wire g162_p_spl_10;
  wire g162_p_spl_11;
  wire g145_p_spl_;
  wire g145_p_spl_0;
  wire g145_n_spl_;
  wire g145_n_spl_0;
  wire G23_n_spl_;
  wire G24_n_spl_;
  wire G24_n_spl_0;
  wire G24_n_spl_1;
  wire G23_p_spl_;
  wire G24_p_spl_;
  wire G24_p_spl_0;
  wire G24_p_spl_1;
  wire g165_n_spl_;
  wire g165_n_spl_0;
  wire g165_n_spl_00;
  wire g165_n_spl_01;
  wire g165_n_spl_1;
  wire g165_n_spl_10;
  wire g165_n_spl_11;
  wire g165_p_spl_;
  wire g165_p_spl_0;
  wire g165_p_spl_00;
  wire g165_p_spl_01;
  wire g165_p_spl_1;
  wire g165_p_spl_10;
  wire g165_p_spl_11;
  wire g167_n_spl_;
  wire g167_n_spl_0;
  wire g167_p_spl_;
  wire g167_p_spl_0;
  wire g169_n_spl_;
  wire g169_p_spl_;
  wire G40_n_spl_;
  wire G40_n_spl_0;
  wire G40_n_spl_00;
  wire G40_n_spl_01;
  wire G40_n_spl_1;
  wire G40_n_spl_10;
  wire G40_p_spl_;
  wire G40_p_spl_0;
  wire G40_p_spl_00;
  wire G40_p_spl_01;
  wire G40_p_spl_1;
  wire G40_p_spl_10;
  wire g186_p_spl_;
  wire g186_p_spl_0;
  wire g186_p_spl_1;
  wire g186_n_spl_;
  wire g186_n_spl_0;
  wire g186_n_spl_1;
  wire g177_p_spl_;
  wire g177_p_spl_0;
  wire g177_n_spl_;
  wire g177_n_spl_0;
  wire g190_n_spl_;
  wire g190_n_spl_0;
  wire g190_p_spl_;
  wire g190_p_spl_0;
  wire g196_n_spl_;
  wire g196_p_spl_;
  wire g212_p_spl_;
  wire g212_p_spl_0;
  wire g212_p_spl_1;
  wire g212_n_spl_;
  wire g212_n_spl_0;
  wire g212_n_spl_1;
  wire g202_p_spl_;
  wire g202_p_spl_0;
  wire g202_n_spl_;
  wire g202_n_spl_0;
  wire g216_n_spl_;
  wire g216_p_spl_;
  wire g223_n_spl_;
  wire g238_p_spl_;
  wire g238_p_spl_0;
  wire g238_p_spl_1;
  wire g238_n_spl_;
  wire g238_n_spl_0;
  wire g238_n_spl_1;
  wire g229_p_spl_;
  wire g229_p_spl_0;
  wire g229_n_spl_;
  wire g229_n_spl_0;
  wire g242_n_spl_;
  wire g242_n_spl_0;
  wire g242_p_spl_;
  wire g242_p_spl_0;
  wire g217_p_spl_;
  wire g217_p_spl_0;
  wire g217_p_spl_1;
  wire g243_p_spl_;
  wire g243_p_spl_0;
  wire g217_n_spl_;
  wire g217_n_spl_0;
  wire g217_n_spl_1;
  wire g243_n_spl_;
  wire g243_n_spl_0;
  wire g191_p_spl_;
  wire g191_p_spl_0;
  wire g244_p_spl_;
  wire g191_n_spl_;
  wire g191_n_spl_0;
  wire g244_n_spl_;
  wire g168_p_spl_;
  wire g168_p_spl_0;
  wire g245_p_spl_;
  wire g168_n_spl_;
  wire g168_n_spl_0;
  wire g245_n_spl_;
  wire g248_n_spl_;
  wire g248_n_spl_0;
  wire g248_n_spl_1;
  wire g248_p_spl_;
  wire g248_p_spl_0;
  wire g248_p_spl_1;
  wire g259_p_spl_;
  wire g259_p_spl_0;
  wire g259_p_spl_00;
  wire g259_p_spl_1;
  wire g259_n_spl_;
  wire g259_n_spl_0;
  wire g259_n_spl_00;
  wire g259_n_spl_1;
  wire g260_n_spl_;
  wire g260_n_spl_0;
  wire g260_n_spl_1;
  wire g260_p_spl_;
  wire g260_p_spl_0;
  wire g260_p_spl_1;
  wire g269_p_spl_;
  wire g269_n_spl_;
  wire g257_p_spl_;
  wire g257_p_spl_0;
  wire g257_n_spl_;
  wire g257_n_spl_0;
  wire g273_n_spl_;
  wire g273_n_spl_0;
  wire g273_p_spl_;
  wire g273_p_spl_0;
  wire g291_p_spl_;
  wire g291_n_spl_;
  wire g282_p_spl_;
  wire g282_p_spl_0;
  wire g282_n_spl_;
  wire g282_n_spl_0;
  wire g295_n_spl_;
  wire g295_n_spl_0;
  wire g295_p_spl_;
  wire g295_p_spl_0;
  wire G21_p_spl_;
  wire G21_p_spl_0;
  wire G21_p_spl_00;
  wire G21_p_spl_01;
  wire G21_p_spl_1;
  wire G21_p_spl_10;
  wire G21_p_spl_11;
  wire G21_n_spl_;
  wire G21_n_spl_0;
  wire G21_n_spl_00;
  wire G21_n_spl_01;
  wire G21_n_spl_1;
  wire G21_n_spl_10;
  wire G21_n_spl_11;
  wire G29_n_spl_;
  wire G29_p_spl_;
  wire g315_p_spl_;
  wire g315_n_spl_;
  wire g306_p_spl_;
  wire g306_p_spl_0;
  wire g306_n_spl_;
  wire g306_n_spl_0;
  wire g319_n_spl_;
  wire g319_p_spl_;
  wire g326_n_spl_;
  wire G22_p_spl_;
  wire G22_p_spl_0;
  wire G22_p_spl_00;
  wire G22_p_spl_01;
  wire G22_p_spl_1;
  wire G22_p_spl_10;
  wire G22_p_spl_11;
  wire G22_n_spl_;
  wire G22_n_spl_0;
  wire G22_n_spl_00;
  wire G22_n_spl_01;
  wire G22_n_spl_1;
  wire G22_n_spl_10;
  wire G22_n_spl_11;
  wire g341_p_spl_;
  wire g341_n_spl_;
  wire g332_p_spl_;
  wire g332_p_spl_0;
  wire g332_n_spl_;
  wire g332_n_spl_0;
  wire g345_n_spl_;
  wire g345_n_spl_0;
  wire g345_p_spl_;
  wire g345_p_spl_0;
  wire g320_p_spl_;
  wire g320_p_spl_0;
  wire g320_p_spl_1;
  wire g346_p_spl_;
  wire g346_p_spl_0;
  wire g320_n_spl_;
  wire g320_n_spl_0;
  wire g320_n_spl_1;
  wire g346_n_spl_;
  wire g346_n_spl_0;
  wire g296_p_spl_;
  wire g296_p_spl_0;
  wire g347_p_spl_;
  wire g296_n_spl_;
  wire g296_n_spl_0;
  wire g347_n_spl_;
  wire g274_p_spl_;
  wire g274_p_spl_0;
  wire g348_p_spl_;
  wire g274_n_spl_;
  wire g274_n_spl_0;
  wire g348_n_spl_;
  wire g246_p_spl_;
  wire g349_p_spl_;
  wire g349_p_spl_0;
  wire g349_p_spl_1;
  wire g356_n_spl_;
  wire g363_n_spl_;
  wire G27_p_spl_;
  wire G27_p_spl_0;
  wire g79_p_spl_;
  wire g79_p_spl_0;
  wire G27_n_spl_;
  wire G48_p_spl_;
  wire g365_p_spl_;
  wire g365_p_spl_0;
  wire g365_p_spl_1;
  wire G48_n_spl_;
  wire g365_n_spl_;
  wire g365_n_spl_0;
  wire g365_n_spl_1;
  wire g366_p_spl_;
  wire g366_p_spl_0;
  wire g366_p_spl_00;
  wire g366_p_spl_000;
  wire g366_p_spl_001;
  wire g366_p_spl_01;
  wire g366_p_spl_010;
  wire g366_p_spl_011;
  wire g366_p_spl_1;
  wire g366_p_spl_10;
  wire g366_p_spl_100;
  wire g366_p_spl_101;
  wire g366_p_spl_11;
  wire g366_n_spl_;
  wire g366_n_spl_0;
  wire g366_n_spl_00;
  wire g366_n_spl_000;
  wire g366_n_spl_001;
  wire g366_n_spl_01;
  wire g366_n_spl_010;
  wire g366_n_spl_011;
  wire g366_n_spl_1;
  wire g366_n_spl_10;
  wire g366_n_spl_100;
  wire g366_n_spl_101;
  wire g366_n_spl_11;
  wire g367_n_spl_;
  wire g367_p_spl_;
  wire g371_n_spl_;
  wire g371_p_spl_;
  wire G47_p_spl_;
  wire G47_p_spl_0;
  wire G47_p_spl_00;
  wire G47_p_spl_01;
  wire G47_p_spl_1;
  wire G47_p_spl_10;
  wire g374_p_spl_;
  wire g374_p_spl_0;
  wire g374_p_spl_1;
  wire G47_n_spl_;
  wire G47_n_spl_0;
  wire G47_n_spl_00;
  wire G47_n_spl_01;
  wire G47_n_spl_1;
  wire G47_n_spl_10;
  wire g374_n_spl_;
  wire g374_n_spl_0;
  wire g374_n_spl_1;
  wire g370_n_spl_;
  wire g370_n_spl_0;
  wire g370_n_spl_1;
  wire g370_p_spl_;
  wire g370_p_spl_0;
  wire g370_p_spl_1;
  wire g76_p_spl_;
  wire g377_n_spl_;
  wire g377_n_spl_0;
  wire g377_n_spl_00;
  wire g377_n_spl_01;
  wire g377_n_spl_1;
  wire g377_n_spl_10;
  wire g377_n_spl_11;
  wire g379_p_spl_;
  wire g379_p_spl_0;
  wire g379_p_spl_00;
  wire g379_p_spl_01;
  wire g379_p_spl_1;
  wire g379_p_spl_10;
  wire g382_p_spl_;
  wire g382_n_spl_;
  wire g377_p_spl_;
  wire g377_p_spl_0;
  wire g377_p_spl_00;
  wire g377_p_spl_01;
  wire g377_p_spl_1;
  wire g377_p_spl_10;
  wire g384_p_spl_;
  wire g384_p_spl_0;
  wire g384_p_spl_00;
  wire g384_p_spl_01;
  wire g384_p_spl_1;
  wire g384_p_spl_10;
  wire g384_n_spl_;
  wire g384_n_spl_0;
  wire g384_n_spl_00;
  wire g384_n_spl_01;
  wire g384_n_spl_1;
  wire g384_n_spl_10;
  wire g387_n_spl_;
  wire g387_n_spl_0;
  wire g387_p_spl_;
  wire g387_p_spl_0;
  wire g385_n_spl_;
  wire g385_n_spl_0;
  wire g385_n_spl_00;
  wire g385_n_spl_000;
  wire g385_n_spl_001;
  wire g385_n_spl_01;
  wire g385_n_spl_1;
  wire g385_n_spl_10;
  wire g385_n_spl_11;
  wire g385_p_spl_;
  wire g385_p_spl_0;
  wire g385_p_spl_00;
  wire g385_p_spl_000;
  wire g385_p_spl_001;
  wire g385_p_spl_01;
  wire g385_p_spl_1;
  wire g385_p_spl_10;
  wire g385_p_spl_11;
  wire g390_p_spl_;
  wire g390_p_spl_0;
  wire g390_p_spl_1;
  wire g390_n_spl_;
  wire g390_n_spl_0;
  wire g390_n_spl_1;
  wire g394_n_spl_;
  wire g394_n_spl_0;
  wire g394_n_spl_00;
  wire g394_n_spl_01;
  wire g394_n_spl_1;
  wire g394_p_spl_;
  wire g394_p_spl_0;
  wire g394_p_spl_00;
  wire g394_p_spl_01;
  wire g394_p_spl_1;
  wire g55_n_spl_;
  wire g393_p_spl_;
  wire g393_p_spl_0;
  wire g393_p_spl_00;
  wire g393_p_spl_000;
  wire g393_p_spl_001;
  wire g393_p_spl_01;
  wire g393_p_spl_010;
  wire g393_p_spl_011;
  wire g393_p_spl_1;
  wire g393_p_spl_10;
  wire g393_p_spl_100;
  wire g393_p_spl_101;
  wire g393_p_spl_11;
  wire g393_p_spl_110;
  wire g393_p_spl_111;
  wire g393_n_spl_;
  wire g393_n_spl_0;
  wire g393_n_spl_00;
  wire g393_n_spl_000;
  wire g393_n_spl_001;
  wire g393_n_spl_01;
  wire g393_n_spl_010;
  wire g393_n_spl_011;
  wire g393_n_spl_1;
  wire g393_n_spl_10;
  wire g393_n_spl_100;
  wire g393_n_spl_101;
  wire g393_n_spl_11;
  wire g393_n_spl_110;
  wire g393_n_spl_111;
  wire g404_n_spl_;
  wire g404_n_spl_0;
  wire g404_p_spl_;
  wire g404_p_spl_0;
  wire g403_n_spl_;
  wire g403_n_spl_0;
  wire g403_n_spl_1;
  wire g405_p_spl_;
  wire g403_p_spl_;
  wire g403_p_spl_0;
  wire g403_p_spl_1;
  wire g405_n_spl_;
  wire G45_p_spl_;
  wire g406_n_spl_;
  wire g406_n_spl_0;
  wire g406_n_spl_00;
  wire g406_n_spl_000;
  wire g406_n_spl_0000;
  wire g406_n_spl_001;
  wire g406_n_spl_01;
  wire g406_n_spl_010;
  wire g406_n_spl_011;
  wire g406_n_spl_1;
  wire g406_n_spl_10;
  wire g406_n_spl_100;
  wire g406_n_spl_101;
  wire g406_n_spl_11;
  wire g406_n_spl_110;
  wire g406_n_spl_111;
  wire G45_n_spl_;
  wire g406_p_spl_;
  wire g406_p_spl_0;
  wire g406_p_spl_00;
  wire g406_p_spl_000;
  wire g406_p_spl_0000;
  wire g406_p_spl_001;
  wire g406_p_spl_01;
  wire g406_p_spl_010;
  wire g406_p_spl_011;
  wire g406_p_spl_1;
  wire g406_p_spl_10;
  wire g406_p_spl_100;
  wire g406_p_spl_101;
  wire g406_p_spl_11;
  wire g406_p_spl_110;
  wire g406_p_spl_111;
  wire g408_p_spl_;
  wire g408_n_spl_;
  wire G44_p_spl_;
  wire G44_p_spl_0;
  wire g409_n_spl_;
  wire g409_n_spl_0;
  wire g409_n_spl_00;
  wire g409_n_spl_000;
  wire g409_n_spl_001;
  wire g409_n_spl_01;
  wire g409_n_spl_010;
  wire g409_n_spl_011;
  wire g409_n_spl_1;
  wire g409_n_spl_10;
  wire g409_n_spl_100;
  wire g409_n_spl_101;
  wire g409_n_spl_11;
  wire g409_n_spl_110;
  wire g409_n_spl_111;
  wire G44_n_spl_;
  wire G44_n_spl_0;
  wire g409_p_spl_;
  wire g409_p_spl_0;
  wire g409_p_spl_00;
  wire g409_p_spl_000;
  wire g409_p_spl_001;
  wire g409_p_spl_01;
  wire g409_p_spl_010;
  wire g409_p_spl_011;
  wire g409_p_spl_1;
  wire g409_p_spl_10;
  wire g409_p_spl_100;
  wire g409_p_spl_101;
  wire g409_p_spl_11;
  wire g409_p_spl_110;
  wire g409_p_spl_111;
  wire G42_p_spl_;
  wire G42_p_spl_0;
  wire G42_p_spl_1;
  wire g412_n_spl_;
  wire g412_n_spl_0;
  wire g412_n_spl_00;
  wire g412_n_spl_000;
  wire g412_n_spl_0000;
  wire g412_n_spl_0001;
  wire g412_n_spl_001;
  wire g412_n_spl_0010;
  wire g412_n_spl_01;
  wire g412_n_spl_010;
  wire g412_n_spl_011;
  wire g412_n_spl_1;
  wire g412_n_spl_10;
  wire g412_n_spl_100;
  wire g412_n_spl_101;
  wire g412_n_spl_11;
  wire g412_n_spl_110;
  wire g412_n_spl_111;
  wire G42_n_spl_;
  wire G42_n_spl_0;
  wire G42_n_spl_1;
  wire g412_p_spl_;
  wire g412_p_spl_0;
  wire g412_p_spl_00;
  wire g412_p_spl_000;
  wire g412_p_spl_0000;
  wire g412_p_spl_0001;
  wire g412_p_spl_001;
  wire g412_p_spl_0010;
  wire g412_p_spl_01;
  wire g412_p_spl_010;
  wire g412_p_spl_011;
  wire g412_p_spl_1;
  wire g412_p_spl_10;
  wire g412_p_spl_100;
  wire g412_p_spl_101;
  wire g412_p_spl_11;
  wire g412_p_spl_110;
  wire g412_p_spl_111;
  wire g414_n_spl_;
  wire g414_n_spl_0;
  wire g414_n_spl_00;
  wire g414_n_spl_000;
  wire g414_n_spl_0000;
  wire g414_n_spl_0001;
  wire g414_n_spl_001;
  wire g414_n_spl_01;
  wire g414_n_spl_010;
  wire g414_n_spl_011;
  wire g414_n_spl_1;
  wire g414_n_spl_10;
  wire g414_n_spl_100;
  wire g414_n_spl_101;
  wire g414_n_spl_11;
  wire g414_n_spl_110;
  wire g414_n_spl_111;
  wire g414_p_spl_;
  wire g414_p_spl_0;
  wire g414_p_spl_00;
  wire g414_p_spl_000;
  wire g414_p_spl_0000;
  wire g414_p_spl_0001;
  wire g414_p_spl_001;
  wire g414_p_spl_01;
  wire g414_p_spl_010;
  wire g414_p_spl_011;
  wire g414_p_spl_1;
  wire g414_p_spl_10;
  wire g414_p_spl_100;
  wire g414_p_spl_101;
  wire g414_p_spl_11;
  wire g414_p_spl_110;
  wire g414_p_spl_111;
  wire G43_p_spl_;
  wire G43_p_spl_0;
  wire G43_p_spl_1;
  wire G43_n_spl_;
  wire G43_n_spl_0;
  wire G43_n_spl_1;
  wire g416_p_spl_;
  wire g416_n_spl_;
  wire g423_n_spl_;
  wire g423_n_spl_0;
  wire g423_n_spl_00;
  wire g423_n_spl_000;
  wire g423_n_spl_001;
  wire g423_n_spl_01;
  wire g423_n_spl_010;
  wire g423_n_spl_011;
  wire g423_n_spl_1;
  wire g423_n_spl_10;
  wire g423_n_spl_11;
  wire g423_p_spl_;
  wire g423_p_spl_0;
  wire g423_p_spl_00;
  wire g423_p_spl_000;
  wire g423_p_spl_001;
  wire g423_p_spl_01;
  wire g423_p_spl_010;
  wire g423_p_spl_011;
  wire g423_p_spl_1;
  wire g423_p_spl_10;
  wire g423_p_spl_11;
  wire g425_n_spl_;
  wire g425_n_spl_0;
  wire g425_n_spl_00;
  wire g425_n_spl_000;
  wire g425_n_spl_001;
  wire g425_n_spl_01;
  wire g425_n_spl_010;
  wire g425_n_spl_011;
  wire g425_n_spl_1;
  wire g425_n_spl_10;
  wire g425_n_spl_100;
  wire g425_n_spl_101;
  wire g425_n_spl_11;
  wire g425_p_spl_;
  wire g425_p_spl_0;
  wire g425_p_spl_00;
  wire g425_p_spl_000;
  wire g425_p_spl_001;
  wire g425_p_spl_01;
  wire g425_p_spl_010;
  wire g425_p_spl_011;
  wire g425_p_spl_1;
  wire g425_p_spl_10;
  wire g425_p_spl_100;
  wire g425_p_spl_101;
  wire g425_p_spl_11;
  wire g432_n_spl_;
  wire g432_p_spl_;
  wire g430_n_spl_;
  wire g430_p_spl_;
  wire g438_n_spl_;
  wire g438_p_spl_;
  wire g440_n_spl_;
  wire g441_n_spl_;
  wire g440_p_spl_;
  wire g441_p_spl_;
  wire g439_p_spl_;
  wire g439_n_spl_;
  wire g453_n_spl_;
  wire g453_p_spl_;
  wire g452_p_spl_;
  wire g452_p_spl_0;
  wire g452_p_spl_1;
  wire g456_p_spl_;
  wire g456_p_spl_0;
  wire g456_p_spl_1;
  wire g452_n_spl_;
  wire g452_n_spl_0;
  wire g452_n_spl_1;
  wire g456_n_spl_;
  wire g456_n_spl_0;
  wire g456_n_spl_1;
  wire G20_p_spl_;
  wire G20_p_spl_0;
  wire G20_p_spl_00;
  wire G20_p_spl_1;
  wire G20_n_spl_;
  wire G20_n_spl_0;
  wire G20_n_spl_00;
  wire G20_n_spl_1;
  wire G18_p_spl_;
  wire G18_p_spl_0;
  wire G18_p_spl_1;
  wire G18_n_spl_;
  wire G18_n_spl_0;
  wire G18_n_spl_1;
  wire G19_p_spl_;
  wire G19_p_spl_0;
  wire G19_p_spl_00;
  wire G19_p_spl_1;
  wire G19_n_spl_;
  wire G19_n_spl_0;
  wire G19_n_spl_00;
  wire G19_n_spl_1;
  wire g480_n_spl_;
  wire g480_p_spl_;
  wire g500_p_spl_;
  wire g500_p_spl_0;
  wire g500_n_spl_;
  wire g500_n_spl_0;
  wire g379_n_spl_;
  wire g379_n_spl_0;
  wire g379_n_spl_00;
  wire g379_n_spl_01;
  wire g379_n_spl_1;
  wire g503_n_spl_;
  wire g503_p_spl_;
  wire g501_p_spl_;
  wire g504_p_spl_;
  wire g501_n_spl_;
  wire g504_n_spl_;
  wire g510_n_spl_;
  wire g510_p_spl_;
  wire g514_n_spl_;
  wire g514_p_spl_;
  wire g513_p_spl_;
  wire g513_p_spl_0;
  wire g513_p_spl_00;
  wire g513_p_spl_1;
  wire g517_p_spl_;
  wire g517_p_spl_0;
  wire g517_p_spl_00;
  wire g517_p_spl_1;
  wire g513_n_spl_;
  wire g513_n_spl_0;
  wire g513_n_spl_00;
  wire g513_n_spl_1;
  wire g517_n_spl_;
  wire g517_n_spl_0;
  wire g517_n_spl_00;
  wire g517_n_spl_1;
  wire g518_p_spl_;
  wire g519_p_spl_;
  wire g518_n_spl_;
  wire g519_n_spl_;
  wire g349_n_spl_;
  wire g520_n_spl_;
  wire g521_p_spl_;
  wire g521_p_spl_0;
  wire g520_p_spl_;
  wire g521_n_spl_;
  wire g521_n_spl_0;
  wire g528_p_spl_;
  wire g528_n_spl_;
  wire g530_n_spl_;
  wire g530_n_spl_0;
  wire g530_p_spl_;
  wire g530_p_spl_0;
  wire g527_n_spl_;
  wire g527_n_spl_0;
  wire g534_n_spl_;
  wire g534_n_spl_0;
  wire g534_n_spl_1;
  wire g527_p_spl_;
  wire g527_p_spl_0;
  wire g534_p_spl_;
  wire g534_p_spl_0;
  wire g534_p_spl_1;
  wire g552_n_spl_;
  wire g552_p_spl_;
  wire g555_p_spl_;
  wire g555_p_spl_0;
  wire g555_n_spl_;
  wire g555_n_spl_0;
  wire g569_n_spl_;
  wire g569_p_spl_;
  wire g579_n_spl_;
  wire g579_p_spl_;
  wire g594_n_spl_;
  wire g594_p_spl_;
  wire g376_p_spl_;
  wire g376_p_spl_0;
  wire g597_n_spl_;
  wire g597_n_spl_0;
  wire g597_n_spl_00;
  wire g597_n_spl_1;
  wire g376_n_spl_;
  wire g597_p_spl_;
  wire g597_p_spl_0;
  wire g597_p_spl_00;
  wire g597_p_spl_1;
  wire g600_n_spl_;
  wire g600_p_spl_;
  wire g601_n_spl_;
  wire g601_p_spl_;
  wire g603_n_spl_;
  wire g603_p_spl_;
  wire g605_p_spl_;
  wire g605_n_spl_;
  wire g598_n_spl_;
  wire g608_n_spl_;
  wire g598_p_spl_;
  wire g608_p_spl_;
  wire g613_n_spl_;
  wire g613_p_spl_;
  wire g617_p_spl_;
  wire g617_n_spl_;
  wire g616_n_spl_;
  wire g616_n_spl_0;
  wire g616_n_spl_1;
  wire g620_n_spl_;
  wire g620_n_spl_0;
  wire g620_n_spl_1;
  wire g616_p_spl_;
  wire g616_p_spl_0;
  wire g616_p_spl_1;
  wire g620_p_spl_;
  wire g620_p_spl_0;
  wire g620_p_spl_1;
  wire g628_n_spl_;
  wire g628_n_spl_0;
  wire g628_p_spl_;
  wire g628_p_spl_0;
  wire g653_n_spl_;
  wire g654_n_spl_;
  wire g653_p_spl_;
  wire g654_p_spl_;
  wire g649_p_spl_;
  wire g649_n_spl_;
  wire g685_p_spl_;
  wire g685_n_spl_;
  wire g706_n_spl_;
  wire g706_p_spl_;
  wire g705_n_spl_;
  wire g705_p_spl_;
  wire g723_p_spl_;
  wire g723_n_spl_;
  wire g726_p_spl_;
  wire g726_n_spl_;
  wire g724_p_spl_;
  wire g724_p_spl_0;
  wire g729_p_spl_;
  wire g724_n_spl_;
  wire g724_n_spl_0;
  wire g729_n_spl_;
  wire g730_n_spl_;
  wire g730_n_spl_0;
  wire g730_p_spl_;
  wire g730_p_spl_0;
  wire g733_p_spl_;
  wire g735_n_spl_;
  wire g733_n_spl_;
  wire g735_p_spl_;
  wire g738_n_spl_;
  wire g738_n_spl_0;
  wire g738_n_spl_1;
  wire g740_n_spl_;
  wire g740_n_spl_0;
  wire g738_p_spl_;
  wire g738_p_spl_0;
  wire g738_p_spl_1;
  wire g740_p_spl_;
  wire g740_p_spl_0;
  wire g732_p_spl_;
  wire g732_p_spl_0;
  wire g732_p_spl_1;
  wire g741_n_spl_;
  wire g741_n_spl_0;
  wire g732_n_spl_;
  wire g732_n_spl_0;
  wire g732_n_spl_1;
  wire g741_p_spl_;
  wire g741_p_spl_0;
  wire G17_p_spl_;
  wire G17_p_spl_0;
  wire G17_n_spl_;
  wire G17_n_spl_0;
  wire G16_n_spl_;
  wire G16_p_spl_;
  wire g779_n_spl_;
  wire g779_p_spl_;
  wire g782_p_spl_;
  wire g782_p_spl_0;
  wire g782_n_spl_;
  wire g782_n_spl_0;
  wire g818_p_spl_;
  wire g818_n_spl_;
  wire g626_p_spl_;
  wire g722_p_spl_;
  wire g626_n_spl_;
  wire g626_n_spl_0;
  wire g722_n_spl_;
  wire g722_n_spl_0;
  wire g778_p_spl_;
  wire g827_p_spl_;
  wire g778_n_spl_;
  wire g778_n_spl_0;
  wire g827_n_spl_;
  wire g827_n_spl_0;
  wire g509_p_spl_;
  wire g866_p_spl_;
  wire g509_n_spl_;
  wire g509_n_spl_0;
  wire g866_n_spl_;
  wire g866_n_spl_0;
  wire g451_p_spl_;
  wire g679_p_spl_;
  wire g451_n_spl_;
  wire g451_n_spl_0;
  wire g679_n_spl_;
  wire g679_n_spl_0;
  wire g869_n_spl_;
  wire g870_n_spl_;
  wire g868_n_spl_;
  wire g868_n_spl_0;
  wire g867_n_spl_;
  wire g874_n_spl_;
  wire g873_n_spl_;
  wire g879_p_spl_;
  wire g881_n_spl_;
  wire g879_n_spl_;
  wire g881_p_spl_;
  wire G50_n_spl_;
  wire g888_n_spl_;
  wire g888_n_spl_0;
  wire g888_n_spl_1;
  wire G50_p_spl_;
  wire g888_p_spl_;
  wire g888_p_spl_0;
  wire g888_p_spl_1;
  wire g886_p_spl_;
  wire g886_p_spl_0;
  wire g886_p_spl_1;
  wire g892_n_spl_;
  wire g886_n_spl_;
  wire g886_n_spl_0;
  wire g886_n_spl_1;
  wire g892_p_spl_;
  wire g884_n_spl_;
  wire g884_p_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  buf

  (
    G42_p,
    G42
  );


  not

  (
    G42_n,
    G42
  );


  buf

  (
    G43_p,
    G43
  );


  not

  (
    G43_n,
    G43
  );


  buf

  (
    G44_p,
    G44
  );


  not

  (
    G44_n,
    G44
  );


  buf

  (
    G45_p,
    G45
  );


  not

  (
    G45_n,
    G45
  );


  buf

  (
    G46_p,
    G46
  );


  not

  (
    G46_n,
    G46
  );


  buf

  (
    G47_p,
    G47
  );


  not

  (
    G47_n,
    G47
  );


  buf

  (
    G48_p,
    G48
  );


  not

  (
    G48_n,
    G48
  );


  buf

  (
    G49_p,
    G49
  );


  not

  (
    G49_n,
    G49
  );


  buf

  (
    G50_p,
    G50
  );


  not

  (
    G50_n,
    G50
  );


  and

  (
    g51_p,
    G7_n_spl_0000,
    G8_n_spl_000
  );


  or

  (
    g51_n,
    G7_p_spl_0000,
    G8_p_spl_000
  );


  and

  (
    g52_p,
    G9_n_spl_000,
    g51_p_spl_
  );


  or

  (
    g52_n,
    G9_p_spl_000,
    g51_n_spl_
  );


  and

  (
    g53_p,
    G10_n_spl_000,
    g52_p_spl_
  );


  and

  (
    g54_p,
    G12_n_spl_000,
    G13_n_spl_000
  );


  or

  (
    g54_n,
    G12_p_spl_000,
    G13_p_spl_000
  );


  and

  (
    g55_p,
    G11_p_spl_000,
    g54_n_spl_
  );


  or

  (
    g55_n,
    G11_n_spl_000,
    g54_p_spl_
  );


  and

  (
    g56_p,
    G1_n_spl_000,
    G3_n_spl_0000
  );


  or

  (
    g57_n,
    G11_p_spl_000,
    G34_n_spl_00
  );


  or

  (
    g58_n,
    G9_p_spl_000,
    G32_n_spl_00
  );


  and

  (
    g59_p,
    g57_n,
    g58_n
  );


  or

  (
    g60_n,
    G13_p_spl_000,
    G36_n_spl_00
  );


  or

  (
    g61_n,
    G10_p_spl_000,
    G33_n_spl_00
  );


  and

  (
    g62_p,
    g60_n,
    g61_n
  );


  and

  (
    g63_p,
    g59_p,
    g62_p
  );


  or

  (
    g64_n,
    G14_p_spl_000,
    G37_n_spl_0
  );


  or

  (
    g65_n,
    G8_p_spl_000,
    G31_n_spl_00
  );


  and

  (
    g66_p,
    g64_n,
    g65_n
  );


  or

  (
    g67_n,
    G12_p_spl_000,
    G35_n_spl_00
  );


  or

  (
    g68_n,
    G7_p_spl_0000,
    G30_n_spl_00
  );


  and

  (
    g69_p,
    g67_n,
    g68_n
  );


  and

  (
    g70_p,
    g66_p,
    g69_p
  );


  and

  (
    g71_p,
    g63_p,
    g70_p
  );


  or

  (
    g72_n,
    g56_p,
    g71_p
  );


  and

  (
    g73_p,
    G1_n_spl_000,
    G2_p_spl_00
  );


  or

  (
    g73_n,
    G1_p_spl_000,
    G2_n_spl_00
  );


  and

  (
    g74_p,
    G3_n_spl_0000,
    g73_p_spl_0
  );


  or

  (
    g74_n,
    G3_p_spl_0000,
    g73_n_spl_0
  );


  and

  (
    g75_p,
    G8_n_spl_000,
    G9_n_spl_000
  );


  or

  (
    g75_n,
    G8_p_spl_001,
    G9_p_spl_001
  );


  and

  (
    g76_p,
    G7_n_spl_0000,
    g75_n_spl_
  );


  or

  (
    g76_n,
    G7_p_spl_0001,
    g75_p_spl_
  );


  or

  (
    g77_n,
    g74_n_spl_,
    g76_n_spl_
  );


  and

  (
    g78_p,
    G1_n_spl_001,
    G2_n_spl_00
  );


  or

  (
    g78_n,
    G1_p_spl_000,
    G2_p_spl_00
  );


  and

  (
    g79_p,
    G3_n_spl_0001,
    g78_p_spl_
  );


  or

  (
    g79_n,
    G3_p_spl_0000,
    g78_n_spl_
  );


  and

  (
    g80_p,
    G35_n_spl_00,
    G36_n_spl_00
  );


  or

  (
    g81_n,
    G34_n_spl_00,
    g80_p
  );


  or

  (
    g82_n,
    g79_n_spl_0,
    g81_n
  );


  and

  (
    g83_p,
    g77_n,
    g82_n
  );


  and

  (
    g84_p,
    g72_n,
    g83_p
  );


  and

  (
    g85_p,
    G36_n_spl_01,
    G37_n_spl_0
  );


  or

  (
    g85_n,
    G36_p_spl_0,
    G37_p_spl_0
  );


  and

  (
    g86_p,
    G36_p_spl_0,
    G37_p_spl_0
  );


  or

  (
    g86_n,
    G36_n_spl_01,
    G37_n_spl_1
  );


  and

  (
    g87_p,
    g85_n,
    g86_n
  );


  or

  (
    g87_n,
    g85_p,
    g86_p
  );


  and

  (
    g88_p,
    G34_n_spl_01,
    G35_n_spl_01
  );


  or

  (
    g88_n,
    G34_p_spl_00,
    G35_p_spl_00
  );


  and

  (
    g89_p,
    G34_p_spl_00,
    G35_p_spl_00
  );


  or

  (
    g89_n,
    G34_n_spl_01,
    G35_n_spl_01
  );


  and

  (
    g90_p,
    g88_n,
    g89_n
  );


  or

  (
    g90_n,
    g88_p,
    g89_p
  );


  and

  (
    g91_p,
    g87_p_spl_,
    g90_n_spl_
  );


  or

  (
    g91_n,
    g87_n_spl_,
    g90_p_spl_
  );


  and

  (
    g92_p,
    g87_n_spl_,
    g90_p_spl_
  );


  or

  (
    g92_n,
    g87_p_spl_,
    g90_n_spl_
  );


  and

  (
    g93_p,
    g91_n,
    g92_n
  );


  or

  (
    g93_n,
    g91_p,
    g92_p
  );


  and

  (
    g94_p,
    G32_n_spl_00,
    G33_n_spl_00
  );


  or

  (
    g94_n,
    G32_p_spl_00,
    G33_p_spl_00
  );


  and

  (
    g95_p,
    G32_p_spl_00,
    G33_p_spl_00
  );


  or

  (
    g95_n,
    G32_n_spl_01,
    G33_n_spl_01
  );


  and

  (
    g96_p,
    g94_n,
    g95_n
  );


  or

  (
    g96_n,
    g94_p,
    g95_p
  );


  and

  (
    g97_p,
    G30_n_spl_00,
    G31_n_spl_00
  );


  or

  (
    g97_n,
    G30_p_spl_00,
    G31_p_spl_00
  );


  and

  (
    g98_p,
    G30_p_spl_00,
    G31_p_spl_00
  );


  or

  (
    g98_n,
    G30_n_spl_01,
    G31_n_spl_01
  );


  and

  (
    g99_p,
    g97_n,
    g98_n
  );


  or

  (
    g99_n,
    g97_p,
    g98_p
  );


  and

  (
    g100_p,
    g96_n_spl_,
    g99_p_spl_
  );


  or

  (
    g100_n,
    g96_p_spl_,
    g99_n_spl_
  );


  and

  (
    g101_p,
    g96_p_spl_,
    g99_n_spl_
  );


  or

  (
    g101_n,
    g96_n_spl_,
    g99_p_spl_
  );


  and

  (
    g102_p,
    g100_n,
    g101_n
  );


  or

  (
    g102_n,
    g100_p,
    g101_p
  );


  or

  (
    g103_n,
    g93_p,
    g102_p_spl_
  );


  or

  (
    g104_n,
    g93_n,
    g102_n_spl_
  );


  and

  (
    g105_p,
    g103_n,
    g104_n
  );


  and

  (
    g106_p,
    G11_n_spl_000,
    G12_n_spl_000
  );


  or

  (
    g106_n,
    G11_p_spl_001,
    G12_p_spl_001
  );


  and

  (
    g107_p,
    G11_p_spl_001,
    G12_p_spl_001
  );


  or

  (
    g107_n,
    G11_n_spl_001,
    G12_n_spl_001
  );


  and

  (
    g108_p,
    g106_n_spl_,
    g107_n
  );


  or

  (
    g108_n,
    g106_p_spl_,
    g107_p
  );


  and

  (
    g109_p,
    G13_n_spl_000,
    G14_n_spl_000
  );


  or

  (
    g109_n,
    G13_p_spl_001,
    G14_p_spl_000
  );


  and

  (
    g110_p,
    G13_p_spl_001,
    G14_p_spl_001
  );


  or

  (
    g110_n,
    G13_n_spl_001,
    G14_n_spl_000
  );


  and

  (
    g111_p,
    g109_n,
    g110_n
  );


  or

  (
    g111_n,
    g109_p,
    g110_p
  );


  and

  (
    g112_p,
    g108_p_spl_,
    g111_n_spl_
  );


  or

  (
    g112_n,
    g108_n_spl_,
    g111_p_spl_
  );


  and

  (
    g113_p,
    g108_n_spl_,
    g111_p_spl_
  );


  or

  (
    g113_n,
    g108_p_spl_,
    g111_n_spl_
  );


  and

  (
    g114_p,
    g112_n,
    g113_n
  );


  or

  (
    g114_n,
    g112_p,
    g113_p
  );


  and

  (
    g115_p,
    G7_p_spl_0001,
    G8_p_spl_001
  );


  or

  (
    g115_n,
    G7_n_spl_000,
    G8_n_spl_001
  );


  and

  (
    g116_p,
    g51_n_spl_,
    g115_n
  );


  or

  (
    g116_n,
    g51_p_spl_,
    g115_p
  );


  and

  (
    g117_p,
    G9_n_spl_001,
    G10_n_spl_000
  );


  or

  (
    g117_n,
    G9_p_spl_001,
    G10_p_spl_000
  );


  and

  (
    g118_p,
    G9_p_spl_010,
    G10_p_spl_001
  );


  or

  (
    g118_n,
    G9_n_spl_001,
    G10_n_spl_001
  );


  and

  (
    g119_p,
    g117_n_spl_,
    g118_n
  );


  or

  (
    g119_n,
    g117_p_spl_,
    g118_p
  );


  and

  (
    g120_p,
    g116_p_spl_,
    g119_n_spl_
  );


  or

  (
    g120_n,
    g116_n_spl_,
    g119_p_spl_
  );


  and

  (
    g121_p,
    g116_n_spl_,
    g119_p_spl_
  );


  or

  (
    g121_n,
    g116_p_spl_,
    g119_n_spl_
  );


  and

  (
    g122_p,
    g120_n,
    g121_n
  );


  or

  (
    g122_n,
    g120_p,
    g121_p
  );


  and

  (
    g123_p,
    g114_n,
    g122_p_spl_
  );


  and

  (
    g124_p,
    g114_p,
    g122_n_spl_
  );


  or

  (
    g125_n,
    g123_p,
    g124_p
  );


  and

  (
    g126_p,
    G1_p_spl_00,
    G2_p_spl_0
  );


  or

  (
    g126_n,
    G1_n_spl_001,
    G2_n_spl_0
  );


  and

  (
    g127_p,
    G1_p_spl_01,
    G3_p_spl_0001
  );


  or

  (
    g127_n,
    G1_n_spl_010,
    G3_n_spl_0001
  );


  and

  (
    g128_p,
    G4_p_spl_00000,
    g127_p
  );


  or

  (
    g128_n,
    G4_n_spl_00000,
    g127_n
  );


  and

  (
    g129_p,
    g126_n_spl_,
    g128_n
  );


  or

  (
    g129_n,
    g126_p_spl_,
    g128_p
  );


  and

  (
    g130_p,
    G3_p_spl_0001,
    g73_p_spl_0
  );


  or

  (
    g130_n,
    G3_n_spl_0010,
    g73_n_spl_0
  );


  and

  (
    g131_p,
    g129_p_spl_000,
    g130_n_spl_00
  );


  or

  (
    g131_n,
    g129_n_spl_000,
    g130_p_spl_00
  );


  and

  (
    g132_p,
    G1_n_spl_010,
    G4_p_spl_00000
  );


  or

  (
    g132_n,
    G1_p_spl_01,
    G4_n_spl_00000
  );


  and

  (
    g133_p,
    g131_p_spl_,
    g132_n
  );


  or

  (
    g133_n,
    g131_n_spl_,
    g132_p
  );


  and

  (
    g134_p,
    G3_p_spl_001,
    g129_n_spl_000
  );


  or

  (
    g134_n,
    G3_n_spl_0010,
    g129_p_spl_000
  );


  and

  (
    g135_p,
    g133_n_spl_0,
    g134_n_spl_0
  );


  or

  (
    g135_n,
    g133_p_spl_0,
    g134_p_spl_0
  );


  and

  (
    g136_p,
    G14_p_spl_001,
    g135_n
  );


  or

  (
    g136_n,
    G14_n_spl_001,
    g135_p
  );


  and

  (
    g137_p,
    G3_n_spl_001,
    G4_p_spl_00001
  );


  or

  (
    g137_n,
    G3_p_spl_001,
    G4_n_spl_00001
  );


  and

  (
    g138_p,
    G3_n_spl_010,
    g137_n_spl_000
  );


  or

  (
    g138_n,
    G3_p_spl_010,
    g137_p_spl_000
  );


  and

  (
    g139_p,
    G12_n_spl_001,
    g138_p_spl_00
  );


  or

  (
    g139_n,
    G12_p_spl_010,
    g138_n_spl_00
  );


  and

  (
    g140_p,
    G39_p_spl_000,
    g137_p_spl_000
  );


  or

  (
    g140_n,
    G39_n_spl_000,
    g137_n_spl_000
  );


  and

  (
    g141_p,
    g139_n,
    g140_n
  );


  or

  (
    g141_n,
    g139_p,
    g140_p
  );


  and

  (
    g142_p,
    g129_n_spl_001,
    g141_n
  );


  or

  (
    g142_n,
    g129_p_spl_001,
    g141_p
  );


  and

  (
    g143_p,
    G14_n_spl_001,
    g130_p_spl_00
  );


  or

  (
    g143_n,
    G14_p_spl_010,
    g130_n_spl_00
  );


  and

  (
    g144_p,
    g142_n,
    g143_n
  );


  or

  (
    g144_n,
    g142_p,
    g143_p
  );


  and

  (
    g145_p,
    g136_n,
    g144_p
  );


  or

  (
    g145_n,
    g136_p,
    g144_n
  );


  and

  (
    g146_p,
    G4_p_spl_00001,
    G5_p_spl_00
  );


  or

  (
    g146_n,
    G4_n_spl_00001,
    G5_n_spl_00
  );


  and

  (
    g147_p,
    g126_p_spl_,
    g146_n_spl_
  );


  or

  (
    g147_n,
    g126_n_spl_,
    g146_p_spl_
  );


  and

  (
    g148_p,
    G38_p,
    g147_n_spl_000
  );


  or

  (
    g148_n,
    G38_n,
    g147_p_spl_000
  );


  and

  (
    g149_p,
    G1_n_spl_01,
    G6_n_spl_00
  );


  or

  (
    g149_n,
    G1_p_spl_10,
    G6_p_spl_00
  );


  and

  (
    g150_p,
    G5_n_spl_00,
    g149_p_spl_0
  );


  or

  (
    g150_n,
    G5_p_spl_00,
    g149_n_spl_0
  );


  and

  (
    g151_p,
    g148_p_spl_0,
    g150_p_spl_0
  );


  or

  (
    g151_n,
    g148_n_spl_0,
    g150_n_spl_0
  );


  and

  (
    g152_p,
    G37_p_spl_,
    g150_n_spl_0
  );


  or

  (
    g152_n,
    G37_n_spl_1,
    g150_p_spl_0
  );


  and

  (
    g153_p,
    G4_n_spl_00010,
    G49_n
  );


  or

  (
    g153_n,
    G4_p_spl_00010,
    G49_p
  );


  and

  (
    g154_p,
    G35_p_spl_0,
    g153_p_spl_00
  );


  or

  (
    g154_n,
    G35_n_spl_10,
    g153_n_spl_00
  );


  and

  (
    g155_p,
    g152_n,
    g154_n
  );


  or

  (
    g155_n,
    g152_p,
    g154_p
  );


  and

  (
    g156_p,
    G4_n_spl_00010,
    G41_n_spl_00
  );


  or

  (
    g156_n,
    G4_p_spl_00010,
    G41_p_spl_00
  );


  and

  (
    g157_p,
    G4_p_spl_00011,
    G36_n_spl_1
  );


  or

  (
    g157_n,
    G4_n_spl_00011,
    G36_p_spl_1
  );


  and

  (
    g158_p,
    g156_n,
    g157_n
  );


  or

  (
    g158_n,
    g156_p,
    g157_p
  );


  and

  (
    g159_p,
    g155_p,
    g158_n
  );


  or

  (
    g159_n,
    g155_n,
    g158_p
  );


  and

  (
    g160_p,
    g147_n_spl_000,
    g159_n
  );


  or

  (
    g160_n,
    g147_p_spl_000,
    g159_p
  );


  and

  (
    g161_p,
    g151_n_spl_0,
    g160_n
  );


  or

  (
    g161_n,
    g151_p_spl_0,
    g160_p
  );


  and

  (
    g162_p,
    G25_n_spl_,
    G26_n_spl_0
  );


  or

  (
    g162_n,
    G25_p_spl_,
    G26_p_spl_0
  );


  and

  (
    g163_p,
    g161_p_spl_0,
    g162_n_spl_000
  );


  or

  (
    g163_n,
    g161_n_spl_0,
    g162_p_spl_000
  );


  and

  (
    g164_p,
    g145_p_spl_0,
    g163_n
  );


  or

  (
    g164_n,
    g145_n_spl_0,
    g163_p
  );


  and

  (
    g165_p,
    G23_n_spl_,
    G24_n_spl_0
  );


  or

  (
    g165_n,
    G23_p_spl_,
    G24_p_spl_0
  );


  and

  (
    g166_p,
    g145_n_spl_0,
    g161_p_spl_0
  );


  or

  (
    g166_n,
    g145_p_spl_0,
    g161_n_spl_0
  );


  and

  (
    g167_p,
    g165_n_spl_00,
    g166_p
  );


  or

  (
    g167_n,
    g165_p_spl_00,
    g166_n
  );


  and

  (
    g168_p,
    g164_n,
    g167_n_spl_0
  );


  or

  (
    g168_n,
    g164_p,
    g167_p_spl_0
  );


  and

  (
    g169_p,
    g130_n_spl_01,
    g134_n_spl_0
  );


  or

  (
    g169_n,
    g130_p_spl_01,
    g134_p_spl_0
  );


  and

  (
    g170_p,
    G13_n_spl_001,
    g169_n_spl_
  );


  or

  (
    g170_n,
    G13_p_spl_010,
    g169_p_spl_
  );


  and

  (
    g171_p,
    G11_n_spl_001,
    g138_p_spl_00
  );


  or

  (
    g171_n,
    G11_p_spl_010,
    g138_n_spl_00
  );


  and

  (
    g172_p,
    G14_p_spl_010,
    g137_p_spl_00
  );


  or

  (
    g172_n,
    G14_n_spl_010,
    g137_n_spl_00
  );


  and

  (
    g173_p,
    g171_n,
    g172_n
  );


  or

  (
    g173_n,
    g171_p,
    g172_p
  );


  and

  (
    g174_p,
    g129_n_spl_001,
    g173_n
  );


  or

  (
    g174_n,
    g129_p_spl_001,
    g173_p
  );


  and

  (
    g175_p,
    G13_p_spl_010,
    g133_p_spl_0
  );


  or

  (
    g175_n,
    G13_n_spl_010,
    g133_n_spl_0
  );


  and

  (
    g176_p,
    g174_n,
    g175_n
  );


  or

  (
    g176_n,
    g174_p,
    g175_p
  );


  and

  (
    g177_p,
    g170_n,
    g176_p
  );


  or

  (
    g177_n,
    g170_p,
    g176_n
  );


  and

  (
    g178_p,
    G36_p_spl_1,
    g150_n_spl_1
  );


  or

  (
    g178_n,
    G36_n_spl_1,
    g150_p_spl_1
  );


  and

  (
    g179_p,
    G34_p_spl_0,
    g153_p_spl_00
  );


  or

  (
    g179_n,
    G34_n_spl_10,
    g153_n_spl_00
  );


  and

  (
    g180_p,
    g178_n,
    g179_n
  );


  or

  (
    g180_n,
    g178_p,
    g179_p
  );


  and

  (
    g181_p,
    G4_n_spl_00011,
    G40_n_spl_00
  );


  or

  (
    g181_n,
    G4_p_spl_00011,
    G40_p_spl_00
  );


  and

  (
    g182_p,
    G4_p_spl_0010,
    G35_n_spl_10
  );


  or

  (
    g182_n,
    G4_n_spl_0010,
    G35_p_spl_1
  );


  and

  (
    g183_p,
    g181_n,
    g182_n
  );


  or

  (
    g183_n,
    g181_p,
    g182_p
  );


  and

  (
    g184_p,
    g180_p,
    g183_n
  );


  or

  (
    g184_n,
    g180_n,
    g183_p
  );


  and

  (
    g185_p,
    g147_n_spl_00,
    g184_n
  );


  or

  (
    g185_n,
    g147_p_spl_00,
    g184_p
  );


  and

  (
    g186_p,
    g151_n_spl_0,
    g185_n
  );


  or

  (
    g186_n,
    g151_p_spl_0,
    g185_p
  );


  and

  (
    g187_p,
    g162_n_spl_000,
    g186_p_spl_0
  );


  or

  (
    g187_n,
    g162_p_spl_000,
    g186_n_spl_0
  );


  and

  (
    g188_p,
    g177_p_spl_0,
    g187_n
  );


  or

  (
    g188_n,
    g177_n_spl_0,
    g187_p
  );


  and

  (
    g189_p,
    g165_n_spl_00,
    g177_n_spl_0
  );


  or

  (
    g189_n,
    g165_p_spl_00,
    g177_p_spl_0
  );


  and

  (
    g190_p,
    g186_p_spl_0,
    g189_p
  );


  or

  (
    g190_n,
    g186_n_spl_0,
    g189_n
  );


  and

  (
    g191_p,
    g188_n,
    g190_n_spl_0
  );


  or

  (
    g191_n,
    g188_p,
    g190_p_spl_0
  );


  and

  (
    g192_p,
    G11_p_spl_010,
    g133_n_spl_1
  );


  or

  (
    g192_n,
    G11_n_spl_010,
    g133_p_spl_1
  );


  and

  (
    g193_p,
    G11_n_spl_010,
    g130_n_spl_01
  );


  or

  (
    g193_n,
    G11_p_spl_011,
    g130_p_spl_01
  );


  and

  (
    g194_p,
    g192_n,
    g193_n
  );


  or

  (
    g194_n,
    g192_p,
    g193_p
  );


  and

  (
    g195_p,
    G12_n_spl_010,
    g137_p_spl_01
  );


  or

  (
    g195_n,
    G12_p_spl_010,
    g137_n_spl_01
  );


  and

  (
    g196_p,
    G13_n_spl_010,
    g106_p_spl_
  );


  or

  (
    g196_n,
    G13_p_spl_011,
    g106_n_spl_
  );


  and

  (
    g197_p,
    G3_p_spl_010,
    g196_n_spl_
  );


  or

  (
    g197_n,
    G3_n_spl_010,
    g196_p_spl_
  );


  and

  (
    g198_p,
    G9_n_spl_010,
    g138_p_spl_01
  );


  or

  (
    g198_n,
    G9_p_spl_010,
    g138_n_spl_01
  );


  and

  (
    g199_p,
    g197_n,
    g198_n
  );


  or

  (
    g199_n,
    g197_p,
    g198_p
  );


  and

  (
    g200_p,
    g195_n,
    g199_p
  );


  or

  (
    g200_n,
    g195_p,
    g199_n
  );


  and

  (
    g201_p,
    g129_n_spl_01,
    g200_n
  );


  or

  (
    g201_n,
    g129_p_spl_01,
    g200_p
  );


  and

  (
    g202_p,
    g194_n,
    g201_n
  );


  or

  (
    g202_n,
    g194_p,
    g201_p
  );


  and

  (
    g203_p,
    g148_p_spl_0,
    g149_p_spl_0
  );


  or

  (
    g203_n,
    g148_n_spl_0,
    g149_n_spl_0
  );


  and

  (
    g204_p,
    G4_p_spl_0010,
    G33_p_spl_0
  );


  or

  (
    g204_n,
    G4_n_spl_0010,
    G33_n_spl_01
  );


  and

  (
    g205_p,
    G4_n_spl_0011,
    G14_p_spl_011
  );


  or

  (
    g205_n,
    G4_p_spl_0011,
    G14_n_spl_010
  );


  and

  (
    g206_p,
    g204_n,
    g205_n
  );


  or

  (
    g206_n,
    g204_p,
    g205_p
  );


  and

  (
    g207_p,
    G34_p_spl_1,
    g149_n_spl_
  );


  or

  (
    g207_n,
    G34_n_spl_10,
    g149_p_spl_
  );


  and

  (
    g208_p,
    G32_p_spl_0,
    g153_p_spl_01
  );


  or

  (
    g208_n,
    G32_n_spl_01,
    g153_n_spl_01
  );


  and

  (
    g209_p,
    g207_n,
    g208_n
  );


  or

  (
    g209_n,
    g207_p,
    g208_p
  );


  and

  (
    g210_p,
    g206_p,
    g209_p
  );


  or

  (
    g210_n,
    g206_n,
    g209_n
  );


  and

  (
    g211_p,
    g147_n_spl_01,
    g210_n
  );


  or

  (
    g211_n,
    g147_p_spl_01,
    g210_p
  );


  and

  (
    g212_p,
    g203_n,
    g211_n
  );


  or

  (
    g212_n,
    g203_p,
    g211_p
  );


  and

  (
    g213_p,
    g162_n_spl_00,
    g212_p_spl_0
  );


  or

  (
    g213_n,
    g162_p_spl_00,
    g212_n_spl_0
  );


  and

  (
    g214_p,
    g202_p_spl_0,
    g213_n
  );


  or

  (
    g214_n,
    g202_n_spl_0,
    g213_p
  );


  and

  (
    g215_p,
    g165_n_spl_01,
    g202_n_spl_0
  );


  or

  (
    g215_n,
    g165_p_spl_01,
    g202_p_spl_0
  );


  and

  (
    g216_p,
    g212_p_spl_0,
    g215_p
  );


  or

  (
    g216_n,
    g212_n_spl_0,
    g215_n
  );


  and

  (
    g217_p,
    g214_n,
    g216_n_spl_
  );


  or

  (
    g217_n,
    g214_p,
    g216_p_spl_
  );


  and

  (
    g218_p,
    G12_p_spl_011,
    g133_n_spl_1
  );


  or

  (
    g218_n,
    G12_n_spl_010,
    g133_p_spl_1
  );


  and

  (
    g219_p,
    G12_n_spl_011,
    g130_n_spl_10
  );


  or

  (
    g219_n,
    G12_p_spl_011,
    g130_p_spl_10
  );


  and

  (
    g220_p,
    g218_n,
    g219_n
  );


  or

  (
    g220_n,
    g218_p,
    g219_p
  );


  and

  (
    g221_p,
    G13_p_spl_011,
    g137_p_spl_01
  );


  or

  (
    g221_n,
    G13_n_spl_011,
    g137_n_spl_01
  );


  and

  (
    g222_p,
    G12_p_spl_100,
    G13_p_spl_100
  );


  or

  (
    g222_n,
    G12_n_spl_011,
    G13_n_spl_011
  );


  and

  (
    g223_p,
    g54_n_spl_,
    g222_n
  );


  or

  (
    g223_n,
    g54_p_spl_,
    g222_p
  );


  and

  (
    g224_p,
    G3_p_spl_011,
    g223_p
  );


  or

  (
    g224_n,
    G3_n_spl_011,
    g223_n_spl_
  );


  and

  (
    g225_p,
    G10_p_spl_001,
    g138_p_spl_01
  );


  or

  (
    g225_n,
    G10_n_spl_001,
    g138_n_spl_01
  );


  and

  (
    g226_p,
    g224_n,
    g225_n
  );


  or

  (
    g226_n,
    g224_p,
    g225_p
  );


  and

  (
    g227_p,
    g221_n,
    g226_p
  );


  or

  (
    g227_n,
    g221_p,
    g226_n
  );


  and

  (
    g228_p,
    g129_n_spl_01,
    g227_n
  );


  or

  (
    g228_n,
    g129_p_spl_01,
    g227_p
  );


  and

  (
    g229_p,
    g220_n,
    g228_n
  );


  or

  (
    g229_n,
    g220_p,
    g228_p
  );


  and

  (
    g230_p,
    G35_p_spl_1,
    g150_n_spl_1
  );


  or

  (
    g230_n,
    G35_n_spl_1,
    g150_p_spl_1
  );


  and

  (
    g231_p,
    G33_p_spl_1,
    g153_p_spl_01
  );


  or

  (
    g231_n,
    G33_n_spl_1,
    g153_n_spl_01
  );


  and

  (
    g232_p,
    g230_n,
    g231_n
  );


  or

  (
    g232_n,
    g230_p,
    g231_p
  );


  and

  (
    g233_p,
    G4_n_spl_0011,
    G39_n_spl_000
  );


  or

  (
    g233_n,
    G4_p_spl_0011,
    G39_p_spl_000
  );


  and

  (
    g234_p,
    G4_p_spl_0100,
    G34_n_spl_1
  );


  or

  (
    g234_n,
    G4_n_spl_0100,
    G34_p_spl_1
  );


  and

  (
    g235_p,
    g233_n,
    g234_n
  );


  or

  (
    g235_n,
    g233_p,
    g234_p
  );


  and

  (
    g236_p,
    g232_p,
    g235_n
  );


  or

  (
    g236_n,
    g232_n,
    g235_p
  );


  and

  (
    g237_p,
    g147_n_spl_01,
    g236_n
  );


  or

  (
    g237_n,
    g147_p_spl_01,
    g236_p
  );


  and

  (
    g238_p,
    g151_n_spl_,
    g237_n
  );


  or

  (
    g238_n,
    g151_p_spl_,
    g237_p
  );


  and

  (
    g239_p,
    g162_n_spl_01,
    g238_p_spl_0
  );


  or

  (
    g239_n,
    g162_p_spl_01,
    g238_n_spl_0
  );


  and

  (
    g240_p,
    g229_p_spl_0,
    g239_n
  );


  or

  (
    g240_n,
    g229_n_spl_0,
    g239_p
  );


  and

  (
    g241_p,
    g165_n_spl_01,
    g229_n_spl_0
  );


  or

  (
    g241_n,
    g165_p_spl_01,
    g229_p_spl_0
  );


  and

  (
    g242_p,
    g238_p_spl_0,
    g241_p
  );


  or

  (
    g242_n,
    g238_n_spl_0,
    g241_n
  );


  and

  (
    g243_p,
    g240_n,
    g242_n_spl_0
  );


  or

  (
    g243_n,
    g240_p,
    g242_p_spl_0
  );


  and

  (
    g244_p,
    g217_p_spl_0,
    g243_p_spl_0
  );


  or

  (
    g244_n,
    g217_n_spl_0,
    g243_n_spl_0
  );


  and

  (
    g245_p,
    g191_p_spl_0,
    g244_p_spl_
  );


  or

  (
    g245_n,
    g191_n_spl_0,
    g244_n_spl_
  );


  and

  (
    g246_p,
    g168_p_spl_0,
    g245_p_spl_
  );


  or

  (
    g246_n,
    g168_n_spl_0,
    g245_n_spl_
  );


  and

  (
    g247_p,
    G1_n_spl_10,
    G3_p_spl_011
  );


  or

  (
    g247_n,
    G1_p_spl_10,
    G3_n_spl_011
  );


  and

  (
    g248_p,
    g131_p_spl_,
    g247_n
  );


  or

  (
    g248_n,
    g131_n_spl_,
    g247_p
  );


  and

  (
    g249_p,
    g134_n_spl_,
    g248_n_spl_0
  );


  or

  (
    g249_n,
    g134_p_spl_,
    g248_p_spl_0
  );


  and

  (
    g250_p,
    G10_p_spl_010,
    g249_n
  );


  or

  (
    g250_n,
    G10_n_spl_010,
    g249_p
  );


  and

  (
    g251_p,
    G8_n_spl_001,
    g138_p_spl_10
  );


  or

  (
    g251_n,
    G8_p_spl_010,
    g138_n_spl_10
  );


  and

  (
    g252_p,
    G11_n_spl_011,
    g137_p_spl_10
  );


  or

  (
    g252_n,
    G11_p_spl_011,
    g137_n_spl_10
  );


  and

  (
    g253_p,
    g251_n,
    g252_n
  );


  or

  (
    g253_n,
    g251_p,
    g252_p
  );


  and

  (
    g254_p,
    g129_n_spl_10,
    g253_n
  );


  or

  (
    g254_n,
    g129_p_spl_10,
    g253_p
  );


  and

  (
    g255_p,
    G10_n_spl_010,
    g130_p_spl_10
  );


  or

  (
    g255_n,
    G10_p_spl_010,
    g130_n_spl_10
  );


  and

  (
    g256_p,
    g254_n,
    g255_n
  );


  or

  (
    g256_n,
    g254_p,
    g255_p
  );


  and

  (
    g257_p,
    g250_n,
    g256_p
  );


  or

  (
    g257_n,
    g250_p,
    g256_n
  );


  and

  (
    g258_p,
    G5_n_spl_01,
    G6_n_spl_00
  );


  or

  (
    g258_n,
    G5_p_spl_01,
    G6_p_spl_00
  );


  and

  (
    g259_p,
    G1_n_spl_10,
    g258_n
  );


  or

  (
    g259_n,
    G1_p_spl_11,
    g258_p
  );


  and

  (
    g260_p,
    g148_p_spl_,
    g259_p_spl_00
  );


  or

  (
    g260_n,
    g148_n_spl_,
    g259_n_spl_00
  );


  and

  (
    g261_p,
    G33_p_spl_1,
    g259_n_spl_00
  );


  or

  (
    g261_n,
    G33_n_spl_1,
    g259_p_spl_00
  );


  and

  (
    g262_p,
    G31_p_spl_0,
    g153_p_spl_10
  );


  or

  (
    g262_n,
    G31_n_spl_01,
    g153_n_spl_10
  );


  and

  (
    g263_p,
    g261_n,
    g262_n
  );


  or

  (
    g263_n,
    g261_p,
    g262_p
  );


  and

  (
    g264_p,
    G4_n_spl_0100,
    G13_n_spl_100
  );


  or

  (
    g264_n,
    G4_p_spl_0100,
    G13_p_spl_100
  );


  and

  (
    g265_p,
    G4_p_spl_0101,
    G32_n_spl_1
  );


  or

  (
    g265_n,
    G4_n_spl_0101,
    G32_p_spl_1
  );


  and

  (
    g266_p,
    g264_n,
    g265_n
  );


  or

  (
    g266_n,
    g264_p,
    g265_p
  );


  and

  (
    g267_p,
    g263_p,
    g266_n
  );


  or

  (
    g267_n,
    g263_n,
    g266_p
  );


  and

  (
    g268_p,
    g147_n_spl_10,
    g267_n
  );


  or

  (
    g268_n,
    g147_p_spl_10,
    g267_p
  );


  and

  (
    g269_p,
    g260_n_spl_0,
    g268_n
  );


  or

  (
    g269_n,
    g260_p_spl_0,
    g268_p
  );


  and

  (
    g270_p,
    g162_n_spl_01,
    g269_p_spl_
  );


  or

  (
    g270_n,
    g162_p_spl_01,
    g269_n_spl_
  );


  and

  (
    g271_p,
    g257_p_spl_0,
    g270_n
  );


  or

  (
    g271_n,
    g257_n_spl_0,
    g270_p
  );


  and

  (
    g272_p,
    g165_n_spl_10,
    g257_n_spl_0
  );


  or

  (
    g272_n,
    g165_p_spl_10,
    g257_p_spl_0
  );


  and

  (
    g273_p,
    g269_p_spl_,
    g272_p
  );


  or

  (
    g273_n,
    g269_n_spl_,
    g272_n
  );


  and

  (
    g274_p,
    g271_n,
    g273_n_spl_0
  );


  or

  (
    g274_n,
    g271_p,
    g273_p_spl_0
  );


  and

  (
    g275_p,
    G9_n_spl_010,
    g169_n_spl_
  );


  or

  (
    g275_n,
    G9_p_spl_011,
    g169_p_spl_
  );


  and

  (
    g276_p,
    G7_p_spl_001,
    g138_p_spl_10
  );


  or

  (
    g276_n,
    G7_n_spl_001,
    g138_n_spl_10
  );


  and

  (
    g277_p,
    G10_p_spl_011,
    g137_p_spl_10
  );


  or

  (
    g277_n,
    G10_n_spl_011,
    g137_n_spl_10
  );


  and

  (
    g278_p,
    g276_n,
    g277_n
  );


  or

  (
    g278_n,
    g276_p,
    g277_p
  );


  and

  (
    g279_p,
    g129_n_spl_10,
    g278_n
  );


  or

  (
    g279_n,
    g129_p_spl_10,
    g278_p
  );


  and

  (
    g280_p,
    G9_p_spl_011,
    g248_p_spl_0
  );


  or

  (
    g280_n,
    G9_n_spl_011,
    g248_n_spl_0
  );


  and

  (
    g281_p,
    g279_n,
    g280_n
  );


  or

  (
    g281_n,
    g279_p,
    g280_p
  );


  and

  (
    g282_p,
    g275_n,
    g281_p
  );


  or

  (
    g282_n,
    g275_p,
    g281_n
  );


  and

  (
    g283_p,
    G32_p_spl_1,
    g259_n_spl_0
  );


  or

  (
    g283_n,
    G32_n_spl_1,
    g259_p_spl_0
  );


  and

  (
    g284_p,
    G30_p_spl_0,
    g153_p_spl_10
  );


  or

  (
    g284_n,
    G30_n_spl_01,
    g153_n_spl_10
  );


  and

  (
    g285_p,
    g283_n,
    g284_n
  );


  or

  (
    g285_n,
    g283_p,
    g284_p
  );


  and

  (
    g286_p,
    G4_n_spl_0101,
    G12_n_spl_100
  );


  or

  (
    g286_n,
    G4_p_spl_0101,
    G12_p_spl_100
  );


  and

  (
    g287_p,
    G4_p_spl_0110,
    G31_n_spl_1
  );


  or

  (
    g287_n,
    G4_n_spl_0110,
    G31_p_spl_1
  );


  and

  (
    g288_p,
    g286_n,
    g287_n
  );


  or

  (
    g288_n,
    g286_p,
    g287_p
  );


  and

  (
    g289_p,
    g285_p,
    g288_n
  );


  or

  (
    g289_n,
    g285_n,
    g288_p
  );


  and

  (
    g290_p,
    g147_n_spl_10,
    g289_n
  );


  or

  (
    g290_n,
    g147_p_spl_10,
    g289_p
  );


  and

  (
    g291_p,
    g260_n_spl_0,
    g290_n
  );


  or

  (
    g291_n,
    g260_p_spl_0,
    g290_p
  );


  and

  (
    g292_p,
    g162_n_spl_10,
    g291_p_spl_
  );


  or

  (
    g292_n,
    g162_p_spl_10,
    g291_n_spl_
  );


  and

  (
    g293_p,
    g282_p_spl_0,
    g292_n
  );


  or

  (
    g293_n,
    g282_n_spl_0,
    g292_p
  );


  and

  (
    g294_p,
    g165_n_spl_10,
    g282_n_spl_0
  );


  or

  (
    g294_n,
    g165_p_spl_10,
    g282_p_spl_0
  );


  and

  (
    g295_p,
    g291_p_spl_,
    g294_p
  );


  or

  (
    g295_n,
    g291_n_spl_,
    g294_n
  );


  and

  (
    g296_p,
    g293_n,
    g295_n_spl_0
  );


  or

  (
    g296_n,
    g293_p,
    g295_p_spl_0
  );


  and

  (
    g297_p,
    G7_p_spl_001,
    g248_n_spl_1
  );


  or

  (
    g297_n,
    G7_n_spl_001,
    g248_p_spl_1
  );


  and

  (
    g298_p,
    G7_n_spl_010,
    g130_n_spl_11
  );


  or

  (
    g298_n,
    G7_p_spl_010,
    g130_p_spl_11
  );


  and

  (
    g299_p,
    g297_n,
    g298_n
  );


  or

  (
    g299_n,
    g297_p,
    g298_p
  );


  and

  (
    g300_p,
    G8_n_spl_010,
    g137_p_spl_11
  );


  or

  (
    g300_n,
    G8_p_spl_010,
    g137_n_spl_11
  );


  and

  (
    g301_p,
    G3_p_spl_100,
    g52_n
  );


  or

  (
    g301_n,
    G3_n_spl_100,
    g52_p_spl_
  );


  and

  (
    g302_p,
    G21_p_spl_00,
    g138_p_spl_11
  );


  or

  (
    g302_n,
    G21_n_spl_00,
    g138_n_spl_11
  );


  and

  (
    g303_p,
    g301_n,
    g302_n
  );


  or

  (
    g303_n,
    g301_p,
    g302_p
  );


  and

  (
    g304_p,
    g300_n,
    g303_p
  );


  or

  (
    g304_n,
    g300_p,
    g303_n
  );


  and

  (
    g305_p,
    g129_n_spl_11,
    g304_n
  );


  or

  (
    g305_n,
    g129_p_spl_11,
    g304_p
  );


  and

  (
    g306_p,
    g299_n,
    g305_n
  );


  or

  (
    g306_n,
    g299_p,
    g305_p
  );


  and

  (
    g307_p,
    G30_p_spl_1,
    g259_n_spl_1
  );


  or

  (
    g307_n,
    G30_n_spl_1,
    g259_p_spl_1
  );


  and

  (
    g308_p,
    G28_p,
    g153_p_spl_11
  );


  or

  (
    g308_n,
    G28_n,
    g153_n_spl_11
  );


  and

  (
    g309_p,
    g307_n,
    g308_n
  );


  or

  (
    g309_n,
    g307_p,
    g308_p
  );


  and

  (
    g310_p,
    G4_n_spl_0110,
    G10_n_spl_011
  );


  or

  (
    g310_n,
    G4_p_spl_0110,
    G10_p_spl_011
  );


  and

  (
    g311_p,
    G4_p_spl_0111,
    G29_n_spl_
  );


  or

  (
    g311_n,
    G4_n_spl_0111,
    G29_p_spl_
  );


  and

  (
    g312_p,
    g310_n,
    g311_n
  );


  or

  (
    g312_n,
    g310_p,
    g311_p
  );


  and

  (
    g313_p,
    g309_p,
    g312_n
  );


  or

  (
    g313_n,
    g309_n,
    g312_p
  );


  and

  (
    g314_p,
    g147_n_spl_11,
    g313_n
  );


  or

  (
    g314_n,
    g147_p_spl_11,
    g313_p
  );


  and

  (
    g315_p,
    g260_n_spl_1,
    g314_n
  );


  or

  (
    g315_n,
    g260_p_spl_1,
    g314_p
  );


  and

  (
    g316_p,
    g162_n_spl_10,
    g315_p_spl_
  );


  or

  (
    g316_n,
    g162_p_spl_10,
    g315_n_spl_
  );


  and

  (
    g317_p,
    g306_p_spl_0,
    g316_n
  );


  or

  (
    g317_n,
    g306_n_spl_0,
    g316_p
  );


  and

  (
    g318_p,
    g165_n_spl_11,
    g306_n_spl_0
  );


  or

  (
    g318_n,
    g165_p_spl_11,
    g306_p_spl_0
  );


  and

  (
    g319_p,
    g315_p_spl_,
    g318_p
  );


  or

  (
    g319_n,
    g315_n_spl_,
    g318_n
  );


  and

  (
    g320_p,
    g317_n,
    g319_n_spl_
  );


  or

  (
    g320_n,
    g317_p,
    g319_p_spl_
  );


  and

  (
    g321_p,
    G8_p_spl_011,
    g248_n_spl_1
  );


  or

  (
    g321_n,
    G8_n_spl_010,
    g248_p_spl_1
  );


  and

  (
    g322_p,
    G8_n_spl_011,
    g130_n_spl_11
  );


  or

  (
    g322_n,
    G8_p_spl_011,
    g130_p_spl_11
  );


  and

  (
    g323_p,
    g321_n,
    g322_n
  );


  or

  (
    g323_n,
    g321_p,
    g322_p
  );


  and

  (
    g324_p,
    G9_n_spl_011,
    g137_p_spl_11
  );


  or

  (
    g324_n,
    G9_p_spl_100,
    g137_n_spl_11
  );


  and

  (
    g325_p,
    G8_p_spl_100,
    G9_p_spl_100
  );


  or

  (
    g325_n,
    G8_n_spl_011,
    G9_n_spl_100
  );


  and

  (
    g326_p,
    g75_n_spl_,
    g325_n
  );


  or

  (
    g326_n,
    g75_p_spl_,
    g325_p
  );


  and

  (
    g327_p,
    G3_p_spl_100,
    g326_p
  );


  or

  (
    g327_n,
    G3_n_spl_100,
    g326_n_spl_
  );


  and

  (
    g328_p,
    G22_p_spl_00,
    g138_p_spl_11
  );


  or

  (
    g328_n,
    G22_n_spl_00,
    g138_n_spl_11
  );


  and

  (
    g329_p,
    g327_n,
    g328_n
  );


  or

  (
    g329_n,
    g327_p,
    g328_p
  );


  and

  (
    g330_p,
    g324_n,
    g329_p
  );


  or

  (
    g330_n,
    g324_p,
    g329_n
  );


  and

  (
    g331_p,
    g129_n_spl_11,
    g330_n
  );


  or

  (
    g331_n,
    g129_p_spl_11,
    g330_p
  );


  and

  (
    g332_p,
    g323_n,
    g331_n
  );


  or

  (
    g332_n,
    g323_p,
    g331_p
  );


  and

  (
    g333_p,
    G31_p_spl_1,
    g259_n_spl_1
  );


  or

  (
    g333_n,
    G31_n_spl_1,
    g259_p_spl_1
  );


  and

  (
    g334_p,
    G29_p_spl_,
    g153_p_spl_11
  );


  or

  (
    g334_n,
    G29_n_spl_,
    g153_n_spl_11
  );


  and

  (
    g335_p,
    g333_n,
    g334_n
  );


  or

  (
    g335_n,
    g333_p,
    g334_p
  );


  and

  (
    g336_p,
    G4_n_spl_0111,
    G11_n_spl_011
  );


  or

  (
    g336_n,
    G4_p_spl_0111,
    G11_p_spl_100
  );


  and

  (
    g337_p,
    G4_p_spl_1000,
    G30_n_spl_1
  );


  or

  (
    g337_n,
    G4_n_spl_1000,
    G30_p_spl_1
  );


  and

  (
    g338_p,
    g336_n,
    g337_n
  );


  or

  (
    g338_n,
    g336_p,
    g337_p
  );


  and

  (
    g339_p,
    g335_p,
    g338_n
  );


  or

  (
    g339_n,
    g335_n,
    g338_p
  );


  and

  (
    g340_p,
    g147_n_spl_11,
    g339_n
  );


  or

  (
    g340_n,
    g147_p_spl_11,
    g339_p
  );


  and

  (
    g341_p,
    g260_n_spl_1,
    g340_n
  );


  or

  (
    g341_n,
    g260_p_spl_1,
    g340_p
  );


  and

  (
    g342_p,
    g162_n_spl_11,
    g341_p_spl_
  );


  or

  (
    g342_n,
    g162_p_spl_11,
    g341_n_spl_
  );


  and

  (
    g343_p,
    g332_p_spl_0,
    g342_n
  );


  or

  (
    g343_n,
    g332_n_spl_0,
    g342_p
  );


  and

  (
    g344_p,
    g165_n_spl_11,
    g332_n_spl_0
  );


  or

  (
    g344_n,
    g165_p_spl_11,
    g332_p_spl_0
  );


  and

  (
    g345_p,
    g341_p_spl_,
    g344_p
  );


  or

  (
    g345_n,
    g341_n_spl_,
    g344_n
  );


  and

  (
    g346_p,
    g343_n,
    g345_n_spl_0
  );


  or

  (
    g346_n,
    g343_p,
    g345_p_spl_0
  );


  and

  (
    g347_p,
    g320_p_spl_0,
    g346_p_spl_0
  );


  or

  (
    g347_n,
    g320_n_spl_0,
    g346_n_spl_0
  );


  and

  (
    g348_p,
    g296_p_spl_0,
    g347_p_spl_
  );


  or

  (
    g348_n,
    g296_n_spl_0,
    g347_n_spl_
  );


  and

  (
    g349_p,
    g274_p_spl_0,
    g348_p_spl_
  );


  or

  (
    g349_n,
    g274_n_spl_0,
    g348_n_spl_
  );


  and

  (
    g350_p,
    g246_p_spl_,
    g349_p_spl_0
  );


  and

  (
    g351_p,
    g190_p_spl_0,
    g244_p_spl_
  );


  or

  (
    g351_n,
    g190_n_spl_0,
    g244_n_spl_
  );


  and

  (
    g352_p,
    g217_p_spl_0,
    g242_p_spl_0
  );


  or

  (
    g352_n,
    g217_n_spl_0,
    g242_n_spl_0
  );


  and

  (
    g353_p,
    g351_n,
    g352_n
  );


  or

  (
    g353_n,
    g351_p,
    g352_p
  );


  and

  (
    g354_p,
    g167_p_spl_0,
    g245_p_spl_
  );


  or

  (
    g354_n,
    g167_n_spl_0,
    g245_n_spl_
  );


  and

  (
    g355_p,
    g216_n_spl_,
    g354_n
  );


  or

  (
    g355_n,
    g216_p_spl_,
    g354_p
  );


  and

  (
    g356_p,
    g353_p,
    g355_p
  );


  or

  (
    g356_n,
    g353_n,
    g355_n
  );


  and

  (
    g357_p,
    g349_p_spl_0,
    g356_n_spl_
  );


  and

  (
    g358_p,
    g295_p_spl_0,
    g347_p_spl_
  );


  or

  (
    g358_n,
    g295_n_spl_0,
    g347_n_spl_
  );


  and

  (
    g359_p,
    g320_p_spl_0,
    g345_p_spl_0
  );


  or

  (
    g359_n,
    g320_n_spl_0,
    g345_n_spl_0
  );


  and

  (
    g360_p,
    g358_n,
    g359_n
  );


  or

  (
    g360_n,
    g358_p,
    g359_p
  );


  and

  (
    g361_p,
    g273_p_spl_0,
    g348_p_spl_
  );


  or

  (
    g361_n,
    g273_n_spl_0,
    g348_n_spl_
  );


  and

  (
    g362_p,
    g319_n_spl_,
    g361_n
  );


  or

  (
    g362_n,
    g319_p_spl_,
    g361_p
  );


  and

  (
    g363_p,
    g360_p,
    g362_p
  );


  or

  (
    g363_n,
    g360_n,
    g362_n
  );


  or

  (
    g364_n,
    g357_p,
    g363_n_spl_
  );


  and

  (
    g365_p,
    G27_p_spl_0,
    g79_p_spl_0
  );


  or

  (
    g365_n,
    G27_n_spl_,
    g79_n_spl_0
  );


  and

  (
    g366_p,
    G48_p_spl_,
    g365_p_spl_0
  );


  or

  (
    g366_n,
    G48_n_spl_,
    g365_n_spl_0
  );


  and

  (
    g367_p,
    g177_n_spl_,
    g366_p_spl_000
  );


  or

  (
    g367_n,
    g177_p_spl_,
    g366_n_spl_000
  );


  and

  (
    g368_p,
    g191_n_spl_0,
    g367_n_spl_
  );


  or

  (
    g368_n,
    g191_p_spl_0,
    g367_p_spl_
  );


  and

  (
    g369_p,
    g191_p_spl_,
    g367_p_spl_
  );


  or

  (
    g369_n,
    g191_n_spl_,
    g367_n_spl_
  );


  and

  (
    g370_p,
    g368_n,
    g369_n
  );


  or

  (
    g370_n,
    g368_p,
    g369_p
  );


  and

  (
    g371_p,
    g145_n_spl_,
    g366_p_spl_000
  );


  or

  (
    g371_n,
    g145_p_spl_,
    g366_n_spl_000
  );


  and

  (
    g372_p,
    g168_n_spl_0,
    g371_n_spl_
  );


  or

  (
    g372_n,
    g168_p_spl_0,
    g371_p_spl_
  );


  and

  (
    g373_p,
    g168_p_spl_,
    g371_p_spl_
  );


  or

  (
    g373_n,
    g168_n_spl_,
    g371_n_spl_
  );


  and

  (
    g374_p,
    g372_n,
    g373_n
  );


  or

  (
    g374_n,
    g372_p,
    g373_p
  );


  and

  (
    g375_p,
    G47_p_spl_00,
    g374_p_spl_0
  );


  or

  (
    g375_n,
    G47_n_spl_00,
    g374_n_spl_0
  );


  and

  (
    g376_p,
    g370_n_spl_0,
    g375_p
  );


  or

  (
    g376_n,
    g370_p_spl_0,
    g375_n
  );


  and

  (
    g377_p,
    G5_p_spl_01,
    g79_p_spl_0
  );


  or

  (
    g377_n,
    G5_n_spl_01,
    g79_n_spl_1
  );


  and

  (
    g378_p,
    g76_p_spl_,
    g377_n_spl_00
  );


  and

  (
    g379_p,
    g356_n_spl_,
    g366_n_spl_001
  );


  or

  (
    g379_n,
    g356_p,
    g366_p_spl_001
  );


  and

  (
    g380_p,
    G1_n_spl_11,
    g379_p_spl_00
  );


  or

  (
    g381_n,
    g378_p,
    g380_p
  );


  and

  (
    g382_p,
    G2_n_spl_1,
    G3_n_spl_101
  );


  or

  (
    g382_n,
    G2_p_spl_1,
    G3_p_spl_101
  );


  and

  (
    g383_p,
    G6_p_spl_01,
    g382_p_spl_
  );


  or

  (
    g383_n,
    G6_n_spl_01,
    g382_n_spl_
  );


  and

  (
    g384_p,
    G1_n_spl_11,
    g383_n
  );


  or

  (
    g384_n,
    G1_p_spl_11,
    g383_p
  );


  and

  (
    g385_p,
    g377_p_spl_00,
    g384_p_spl_00
  );


  or

  (
    g385_n,
    g377_n_spl_00,
    g384_n_spl_00
  );


  and

  (
    g386_p,
    G47_n_spl_00,
    g374_p_spl_0
  );


  or

  (
    g386_n,
    G47_p_spl_00,
    g374_n_spl_0
  );


  and

  (
    g387_p,
    G47_p_spl_01,
    g374_n_spl_1
  );


  or

  (
    g387_n,
    G47_n_spl_01,
    g374_p_spl_1
  );


  and

  (
    g388_p,
    g386_n,
    g387_n_spl_0
  );


  or

  (
    g388_n,
    g386_p,
    g387_p_spl_0
  );


  and

  (
    g389_p,
    g385_n_spl_000,
    g388_p
  );


  or

  (
    g389_n,
    g385_p_spl_000,
    g388_n
  );


  and

  (
    g390_p,
    G4_p_spl_1000,
    g382_p_spl_
  );


  or

  (
    g390_n,
    G4_n_spl_1000,
    g382_n_spl_
  );


  and

  (
    g391_p,
    g374_p_spl_1,
    g390_p_spl_0
  );


  or

  (
    g391_n,
    g374_n_spl_1,
    g390_n_spl_0
  );


  and

  (
    g392_p,
    G3_p_spl_101,
    G23_n_spl_
  );


  or

  (
    g392_n,
    G3_n_spl_101,
    G23_p_spl_
  );


  and

  (
    g393_p,
    g73_p_spl_,
    g392_n
  );


  or

  (
    g393_n,
    g73_n_spl_,
    g392_p
  );


  and

  (
    g394_p,
    G4_n_spl_1001,
    g79_p_spl_
  );


  or

  (
    g394_n,
    G4_p_spl_1001,
    g79_n_spl_1
  );


  and

  (
    g395_p,
    G14_p_spl_011,
    g394_n_spl_00
  );


  or

  (
    g395_n,
    G14_n_spl_011,
    g394_p_spl_00
  );


  and

  (
    g396_p,
    G6_n_spl_01,
    g122_n_spl_
  );


  or

  (
    g396_n,
    G6_p_spl_01,
    g122_p_spl_
  );


  and

  (
    g397_p,
    G6_p_spl_10,
    g76_n_spl_
  );


  or

  (
    g397_n,
    G6_n_spl_10,
    g76_p_spl_
  );


  and

  (
    g398_p,
    g55_p,
    g397_n
  );


  or

  (
    g398_n,
    g55_n_spl_,
    g397_p
  );


  and

  (
    g399_p,
    g396_n,
    g398_p
  );


  or

  (
    g399_n,
    g396_p,
    g398_n
  );


  and

  (
    g400_p,
    g394_p_spl_00,
    g399_p
  );


  or

  (
    g400_n,
    g394_n_spl_00,
    g399_n
  );


  and

  (
    g401_p,
    g395_n,
    g400_n
  );


  or

  (
    g401_n,
    g395_p,
    g400_p
  );


  and

  (
    g402_p,
    g393_p_spl_000,
    g401_n
  );


  or

  (
    g402_n,
    g393_n_spl_000,
    g401_p
  );


  and

  (
    g403_p,
    G3_p_spl_110,
    G25_p_spl_
  );


  or

  (
    g403_n,
    G3_n_spl_110,
    G25_n_spl_
  );


  and

  (
    g404_p,
    G3_p_spl_110,
    G24_p_spl_0
  );


  or

  (
    g404_n,
    G3_n_spl_110,
    G24_n_spl_0
  );


  and

  (
    g405_p,
    G26_p_spl_0,
    g404_n_spl_0
  );


  or

  (
    g405_n,
    G26_n_spl_0,
    g404_p_spl_0
  );


  and

  (
    g406_p,
    g403_n_spl_0,
    g405_p_spl_
  );


  or

  (
    g406_n,
    g403_p_spl_0,
    g405_n_spl_
  );


  and

  (
    g407_p,
    G45_p_spl_,
    g406_n_spl_0000
  );


  or

  (
    g407_n,
    G45_n_spl_,
    g406_p_spl_0000
  );


  and

  (
    g408_p,
    G26_n_spl_,
    g404_n_spl_0
  );


  or

  (
    g408_n,
    G26_p_spl_,
    g404_p_spl_0
  );


  and

  (
    g409_p,
    g403_n_spl_0,
    g408_p_spl_
  );


  or

  (
    g409_n,
    g403_p_spl_0,
    g408_n_spl_
  );


  and

  (
    g410_p,
    G44_p_spl_0,
    g409_n_spl_000
  );


  or

  (
    g410_n,
    G44_n_spl_0,
    g409_p_spl_000
  );


  and

  (
    g411_p,
    g407_n,
    g410_n
  );


  or

  (
    g411_n,
    g407_p,
    g410_p
  );


  and

  (
    g412_p,
    g403_p_spl_1,
    g408_p_spl_
  );


  or

  (
    g412_n,
    g403_n_spl_1,
    g408_n_spl_
  );


  and

  (
    g413_p,
    G42_p_spl_0,
    g412_n_spl_0000
  );


  or

  (
    g413_n,
    G42_n_spl_0,
    g412_p_spl_0000
  );


  and

  (
    g414_p,
    g403_p_spl_1,
    g405_p_spl_
  );


  or

  (
    g414_n,
    g403_n_spl_1,
    g405_n_spl_
  );


  and

  (
    g415_p,
    G39_p_spl_00,
    g414_n_spl_0000
  );


  or

  (
    g415_n,
    G39_n_spl_00,
    g414_p_spl_0000
  );


  and

  (
    g416_p,
    g413_n,
    g415_n
  );


  or

  (
    g416_n,
    g413_p,
    g415_p
  );


  and

  (
    g417_p,
    G46_p,
    g412_n_spl_0000
  );


  or

  (
    g417_n,
    G46_n,
    g412_p_spl_0000
  );


  and

  (
    g418_p,
    G43_p_spl_0,
    g414_n_spl_0000
  );


  or

  (
    g418_n,
    G43_n_spl_0,
    g414_p_spl_0000
  );


  and

  (
    g419_p,
    g417_n,
    g418_n
  );


  or

  (
    g419_n,
    g417_p,
    g418_p
  );


  and

  (
    g420_p,
    g416_p_spl_,
    g419_p
  );


  or

  (
    g420_n,
    g416_n_spl_,
    g419_n
  );


  and

  (
    g421_p,
    g411_p,
    g420_p
  );


  or

  (
    g421_n,
    g411_n,
    g420_n
  );


  and

  (
    g422_p,
    G3_p_spl_111,
    g162_n_spl_11
  );


  or

  (
    g422_n,
    G3_n_spl_111,
    g162_p_spl_11
  );


  and

  (
    g423_p,
    g404_n_spl_,
    g422_n
  );


  or

  (
    g423_n,
    g404_p_spl_,
    g422_p
  );


  and

  (
    g424_p,
    G40_p_spl_00,
    g423_n_spl_000
  );


  or

  (
    g424_n,
    G40_n_spl_00,
    g423_p_spl_000
  );


  and

  (
    g425_p,
    G3_p_spl_111,
    g406_p_spl_0000
  );


  or

  (
    g425_n,
    G3_n_spl_111,
    g406_n_spl_0000
  );


  and

  (
    g426_p,
    G41_p_spl_00,
    g425_n_spl_000
  );


  or

  (
    g426_n,
    G41_n_spl_00,
    g425_p_spl_000
  );


  and

  (
    g427_p,
    G4_p_spl_1001,
    g426_n
  );


  or

  (
    g427_n,
    G4_n_spl_1001,
    g426_p
  );


  and

  (
    g428_p,
    g424_n,
    g427_p
  );


  or

  (
    g428_n,
    g424_p,
    g427_n
  );


  and

  (
    g429_p,
    g421_p,
    g428_p
  );


  or

  (
    g429_n,
    g421_n,
    g428_n
  );


  and

  (
    g430_p,
    G11_n_spl_100,
    g425_n_spl_000
  );


  or

  (
    g430_n,
    G11_p_spl_100,
    g425_p_spl_000
  );


  and

  (
    g431_p,
    G10_n_spl_100,
    g412_n_spl_0001
  );


  or

  (
    g431_n,
    G10_p_spl_100,
    g412_p_spl_0001
  );


  and

  (
    g432_p,
    G13_n_spl_100,
    g414_n_spl_0001
  );


  or

  (
    g432_n,
    G13_p_spl_101,
    g414_p_spl_0001
  );


  and

  (
    g433_p,
    g431_n,
    g432_n_spl_
  );


  or

  (
    g433_n,
    g431_p,
    g432_p_spl_
  );


  and

  (
    g434_p,
    g430_n_spl_,
    g433_p
  );


  or

  (
    g434_n,
    g430_p_spl_,
    g433_n
  );


  and

  (
    g435_p,
    G7_n_spl_010,
    g406_n_spl_000
  );


  or

  (
    g435_n,
    G7_p_spl_010,
    g406_p_spl_000
  );


  and

  (
    g436_p,
    G8_n_spl_100,
    g409_n_spl_000
  );


  or

  (
    g436_n,
    G8_p_spl_100,
    g409_p_spl_000
  );


  and

  (
    g437_p,
    g435_n,
    g436_n
  );


  or

  (
    g437_n,
    g435_p,
    g436_p
  );


  and

  (
    g438_p,
    G9_n_spl_100,
    g414_n_spl_0001
  );


  or

  (
    g438_n,
    G9_p_spl_101,
    g414_p_spl_0001
  );


  and

  (
    g439_p,
    G4_n_spl_1010,
    g438_n_spl_
  );


  or

  (
    g439_n,
    G4_p_spl_1010,
    g438_p_spl_
  );


  and

  (
    g440_p,
    G12_n_spl_100,
    g423_n_spl_000
  );


  or

  (
    g440_n,
    G12_p_spl_101,
    g423_p_spl_000
  );


  and

  (
    g441_p,
    G22_p_spl_00,
    g412_n_spl_0001
  );


  or

  (
    g441_n,
    G22_n_spl_00,
    g412_p_spl_0001
  );


  and

  (
    g442_p,
    g440_n_spl_,
    g441_n_spl_
  );


  or

  (
    g442_n,
    g440_p_spl_,
    g441_p_spl_
  );


  and

  (
    g443_p,
    g439_p_spl_,
    g442_p
  );


  or

  (
    g443_n,
    g439_n_spl_,
    g442_n
  );


  and

  (
    g444_p,
    g437_p,
    g443_p
  );


  or

  (
    g444_n,
    g437_n,
    g443_n
  );


  and

  (
    g445_p,
    g434_p,
    g444_p
  );


  or

  (
    g445_n,
    g434_n,
    g444_n
  );


  and

  (
    g446_p,
    g429_n,
    g445_n
  );


  or

  (
    g446_n,
    g429_p,
    g445_p
  );


  and

  (
    g447_p,
    g393_n_spl_000,
    g446_p
  );


  or

  (
    g447_n,
    g393_p_spl_000,
    g446_n
  );


  and

  (
    g448_p,
    g402_n,
    g447_n
  );


  or

  (
    g448_n,
    g402_p,
    g447_p
  );


  and

  (
    g449_p,
    g391_n,
    g448_n
  );


  or

  (
    g449_n,
    g391_p,
    g448_p
  );


  and

  (
    g450_p,
    g385_p_spl_000,
    g449_p
  );


  or

  (
    g450_n,
    g385_n_spl_000,
    g449_n
  );


  and

  (
    g451_p,
    g389_n,
    g450_n
  );


  or

  (
    g451_n,
    g389_p,
    g450_p
  );


  and

  (
    g452_p,
    G2_n_spl_1,
    G4_p_spl_1010
  );


  or

  (
    g452_n,
    G2_p_spl_1,
    G4_n_spl_1010
  );


  and

  (
    g453_p,
    g257_n_spl_,
    g366_p_spl_001
  );


  or

  (
    g453_n,
    g257_p_spl_,
    g366_n_spl_001
  );


  and

  (
    g454_p,
    g274_n_spl_0,
    g453_n_spl_
  );


  or

  (
    g454_n,
    g274_p_spl_0,
    g453_p_spl_
  );


  and

  (
    g455_p,
    g274_p_spl_,
    g453_p_spl_
  );


  or

  (
    g455_n,
    g274_n_spl_,
    g453_n_spl_
  );


  and

  (
    g456_p,
    g454_n,
    g455_n
  );


  or

  (
    g456_n,
    g454_p,
    g455_p
  );


  and

  (
    g457_p,
    g452_p_spl_0,
    g456_p_spl_0
  );


  or

  (
    g457_n,
    g452_n_spl_0,
    g456_n_spl_0
  );


  and

  (
    g458_p,
    G10_n_spl_100,
    g393_p_spl_001
  );


  or

  (
    g458_n,
    G10_p_spl_100,
    g393_n_spl_001
  );


  and

  (
    g459_p,
    g385_p_spl_001,
    g458_n
  );


  or

  (
    g459_n,
    g385_n_spl_001,
    g458_p
  );


  and

  (
    g460_p,
    G8_n_spl_100,
    g423_n_spl_001
  );


  or

  (
    g460_n,
    G8_p_spl_101,
    g423_p_spl_001
  );


  and

  (
    g461_p,
    g441_n_spl_,
    g460_n
  );


  or

  (
    g461_n,
    g441_p_spl_,
    g460_p
  );


  and

  (
    g462_p,
    G20_p_spl_00,
    g409_n_spl_001
  );


  or

  (
    g462_n,
    G20_n_spl_00,
    g409_p_spl_001
  );


  and

  (
    g463_p,
    G21_p_spl_00,
    g414_n_spl_001
  );


  or

  (
    g463_n,
    G21_n_spl_00,
    g414_p_spl_001
  );


  and

  (
    g464_p,
    g462_n,
    g463_n
  );


  or

  (
    g464_n,
    g462_p,
    g463_p
  );


  and

  (
    g465_p,
    g439_p_spl_,
    g464_p
  );


  or

  (
    g465_n,
    g439_n_spl_,
    g464_n
  );


  and

  (
    g466_p,
    g461_p,
    g465_p
  );


  or

  (
    g466_n,
    g461_n,
    g465_n
  );


  and

  (
    g467_p,
    G18_p_spl_0,
    g412_n_spl_0010
  );


  or

  (
    g467_n,
    G18_n_spl_0,
    g412_p_spl_0010
  );


  and

  (
    g468_p,
    G7_n_spl_011,
    g425_n_spl_001
  );


  or

  (
    g468_n,
    G7_p_spl_011,
    g425_p_spl_001
  );


  and

  (
    g469_p,
    G19_p_spl_00,
    g406_n_spl_001
  );


  or

  (
    g469_n,
    G19_n_spl_00,
    g406_p_spl_001
  );


  and

  (
    g470_p,
    g468_n,
    g469_n
  );


  or

  (
    g470_n,
    g468_p,
    g469_p
  );


  and

  (
    g471_p,
    g467_n,
    g470_p
  );


  or

  (
    g471_n,
    g467_p,
    g470_n
  );


  and

  (
    g472_p,
    g466_p,
    g471_p
  );


  or

  (
    g472_n,
    g466_n,
    g471_n
  );


  and

  (
    g473_p,
    G13_n_spl_101,
    g425_n_spl_001
  );


  or

  (
    g473_n,
    G13_p_spl_101,
    g425_p_spl_001
  );


  and

  (
    g474_p,
    g416_p_spl_,
    g440_n_spl_
  );


  or

  (
    g474_n,
    g416_n_spl_,
    g440_p_spl_
  );


  and

  (
    g475_p,
    g473_n,
    g474_p
  );


  or

  (
    g475_n,
    g473_p,
    g474_n
  );


  and

  (
    g476_p,
    G40_p_spl_01,
    g409_n_spl_001
  );


  or

  (
    g476_n,
    G40_n_spl_01,
    g409_p_spl_001
  );


  and

  (
    g477_p,
    G14_n_spl_011,
    g412_n_spl_0010
  );


  or

  (
    g477_n,
    G14_p_spl_100,
    g412_p_spl_0010
  );


  and

  (
    g478_p,
    g476_n,
    g477_n
  );


  or

  (
    g478_n,
    g476_p,
    g477_p
  );


  and

  (
    g479_p,
    G41_p_spl_01,
    g406_n_spl_001
  );


  or

  (
    g479_n,
    G41_n_spl_01,
    g406_p_spl_001
  );


  and

  (
    g480_p,
    G11_n_spl_100,
    g414_n_spl_001
  );


  or

  (
    g480_n,
    G11_p_spl_101,
    g414_p_spl_001
  );


  and

  (
    g481_p,
    g479_n,
    g480_n_spl_
  );


  or

  (
    g481_n,
    g479_p,
    g480_p_spl_
  );


  and

  (
    g482_p,
    g478_p,
    g481_p
  );


  or

  (
    g482_n,
    g478_n,
    g481_n
  );


  and

  (
    g483_p,
    G4_p_spl_1011,
    g482_p
  );


  or

  (
    g483_n,
    G4_n_spl_1011,
    g482_n
  );


  and

  (
    g484_p,
    g475_p,
    g483_p
  );


  or

  (
    g484_n,
    g475_n,
    g483_n
  );


  and

  (
    g485_p,
    g472_n,
    g484_n
  );


  or

  (
    g485_n,
    g472_p,
    g484_p
  );


  and

  (
    g486_p,
    g393_n_spl_001,
    g485_n
  );


  or

  (
    g486_n,
    g393_p_spl_001,
    g485_p
  );


  and

  (
    g487_p,
    g459_p,
    g486_n
  );


  or

  (
    g487_n,
    g459_n,
    g486_p
  );


  and

  (
    g488_p,
    g457_n,
    g487_p
  );


  or

  (
    g488_n,
    g457_p,
    g487_n
  );


  and

  (
    g489_p,
    g212_n_spl_1,
    g238_n_spl_1
  );


  or

  (
    g489_n,
    g212_p_spl_1,
    g238_p_spl_1
  );


  and

  (
    g490_p,
    g161_n_spl_1,
    g186_n_spl_1
  );


  or

  (
    g490_n,
    g161_p_spl_1,
    g186_p_spl_1
  );


  and

  (
    g491_p,
    g489_p,
    g490_p
  );


  or

  (
    g491_n,
    g489_n,
    g490_n
  );


  and

  (
    g492_p,
    G24_p_spl_1,
    g491_n
  );


  or

  (
    g492_n,
    G24_n_spl_1,
    g491_p
  );


  and

  (
    g493_p,
    g212_p_spl_1,
    g238_p_spl_1
  );


  or

  (
    g493_n,
    g212_n_spl_1,
    g238_n_spl_1
  );


  and

  (
    g494_p,
    g161_p_spl_1,
    g186_p_spl_1
  );


  or

  (
    g494_n,
    g161_n_spl_1,
    g186_n_spl_1
  );


  and

  (
    g495_p,
    g493_p,
    g494_p
  );


  or

  (
    g495_n,
    g493_n,
    g494_n
  );


  and

  (
    g496_p,
    G24_n_spl_1,
    g495_n
  );


  or

  (
    g496_n,
    G24_p_spl_1,
    g495_p
  );


  and

  (
    g497_p,
    g492_n,
    g496_n
  );


  or

  (
    g497_n,
    g492_p,
    g496_p
  );


  and

  (
    g498_p,
    g366_n_spl_010,
    g497_n
  );


  or

  (
    g498_n,
    g366_p_spl_010,
    g497_p
  );


  and

  (
    g499_p,
    g246_n,
    g366_p_spl_010
  );


  or

  (
    g499_n,
    g246_p_spl_,
    g366_n_spl_010
  );


  and

  (
    g500_p,
    g498_n,
    g499_n
  );


  or

  (
    g500_n,
    g498_p,
    g499_p
  );


  and

  (
    g501_p,
    G47_p_spl_01,
    g500_p_spl_0
  );


  or

  (
    g501_n,
    G47_n_spl_01,
    g500_n_spl_0
  );


  and

  (
    g502_p,
    g379_p_spl_00,
    g456_n_spl_0
  );


  or

  (
    g502_n,
    g379_n_spl_00,
    g456_p_spl_0
  );


  and

  (
    g503_p,
    g379_n_spl_00,
    g456_p_spl_1
  );


  or

  (
    g503_n,
    g379_p_spl_01,
    g456_n_spl_1
  );


  and

  (
    g504_p,
    g502_n,
    g503_n_spl_
  );


  or

  (
    g504_n,
    g502_p,
    g503_p_spl_
  );


  and

  (
    g505_p,
    g501_p_spl_,
    g504_p_spl_
  );


  or

  (
    g505_n,
    g501_n_spl_,
    g504_n_spl_
  );


  and

  (
    g506_p,
    g501_n_spl_,
    g504_n_spl_
  );


  or

  (
    g506_n,
    g501_p_spl_,
    g504_p_spl_
  );


  and

  (
    g507_p,
    g505_n,
    g506_n
  );


  or

  (
    g507_n,
    g505_p,
    g506_p
  );


  and

  (
    g508_p,
    g385_n_spl_001,
    g507_n
  );


  or

  (
    g508_n,
    g385_p_spl_001,
    g507_p
  );


  and

  (
    g509_p,
    g488_n,
    g508_n
  );


  or

  (
    g509_n,
    g488_p,
    g508_p
  );


  and

  (
    g510_p,
    g282_n_spl_,
    g366_p_spl_011
  );


  or

  (
    g510_n,
    g282_p_spl_,
    g366_n_spl_011
  );


  and

  (
    g511_p,
    g296_n_spl_0,
    g510_n_spl_
  );


  or

  (
    g511_n,
    g296_p_spl_0,
    g510_p_spl_
  );


  and

  (
    g512_p,
    g296_p_spl_,
    g510_p_spl_
  );


  or

  (
    g512_n,
    g296_n_spl_,
    g510_n_spl_
  );


  and

  (
    g513_p,
    g511_n,
    g512_n
  );


  or

  (
    g513_n,
    g511_p,
    g512_p
  );


  and

  (
    g514_p,
    g332_n_spl_,
    g365_p_spl_0
  );


  or

  (
    g514_n,
    g332_p_spl_,
    g365_n_spl_0
  );


  and

  (
    g515_p,
    g346_n_spl_0,
    g514_n_spl_
  );


  or

  (
    g515_n,
    g346_p_spl_0,
    g514_p_spl_
  );


  and

  (
    g516_p,
    g346_p_spl_,
    g514_p_spl_
  );


  or

  (
    g516_n,
    g346_n_spl_,
    g514_n_spl_
  );


  and

  (
    g517_p,
    g515_n,
    g516_n
  );


  or

  (
    g517_n,
    g515_p,
    g516_p
  );


  and

  (
    g518_p,
    g513_p_spl_00,
    g517_p_spl_00
  );


  or

  (
    g518_n,
    g513_n_spl_00,
    g517_n_spl_00
  );


  and

  (
    g519_p,
    g456_p_spl_1,
    g500_n_spl_0
  );


  or

  (
    g519_n,
    g456_n_spl_1,
    g500_p_spl_0
  );


  and

  (
    g520_p,
    g518_p_spl_,
    g519_p_spl_
  );


  or

  (
    g520_n,
    g518_n_spl_,
    g519_n_spl_
  );


  and

  (
    g521_p,
    g349_n_spl_,
    g500_n_spl_
  );


  or

  (
    g521_n,
    g349_p_spl_1,
    g500_p_spl_
  );


  and

  (
    g522_p,
    g520_n_spl_,
    g521_p_spl_0
  );


  or

  (
    g522_n,
    g520_p_spl_,
    g521_n_spl_0
  );


  and

  (
    g523_p,
    g520_p_spl_,
    g521_n_spl_0
  );


  or

  (
    g523_n,
    g520_n_spl_,
    g521_p_spl_0
  );


  and

  (
    g524_p,
    g522_n,
    g523_n
  );


  or

  (
    g524_n,
    g522_p,
    g523_p
  );


  and

  (
    g525_p,
    G47_p_spl_10,
    g524_n
  );


  or

  (
    g525_n,
    G47_n_spl_10,
    g524_p
  );


  and

  (
    g526_p,
    g349_n_spl_,
    g379_n_spl_01
  );


  or

  (
    g526_n,
    g349_p_spl_1,
    g379_p_spl_01
  );


  and

  (
    g527_p,
    g363_p,
    g526_n
  );


  or

  (
    g527_n,
    g363_n_spl_,
    g526_p
  );


  and

  (
    g528_p,
    g295_p_spl_,
    g366_n_spl_011
  );


  or

  (
    g528_n,
    g295_n_spl_,
    g366_p_spl_011
  );


  and

  (
    g529_p,
    g517_p_spl_00,
    g528_p_spl_
  );


  or

  (
    g529_n,
    g517_n_spl_00,
    g528_n_spl_
  );


  and

  (
    g530_p,
    g273_p_spl_,
    g366_n_spl_100
  );


  or

  (
    g530_n,
    g273_n_spl_,
    g366_p_spl_100
  );


  and

  (
    g531_p,
    g518_p_spl_,
    g530_n_spl_0
  );


  or

  (
    g531_n,
    g518_n_spl_,
    g530_p_spl_0
  );


  and

  (
    g532_p,
    g345_p_spl_,
    g365_n_spl_1
  );


  or

  (
    g532_n,
    g345_n_spl_,
    g365_p_spl_1
  );


  and

  (
    g533_p,
    g531_n,
    g532_n
  );


  or

  (
    g533_n,
    g531_p,
    g532_p
  );


  and

  (
    g534_p,
    g529_n,
    g533_p
  );


  or

  (
    g534_n,
    g529_p,
    g533_n
  );


  and

  (
    g535_p,
    g527_n_spl_0,
    g534_n_spl_0
  );


  or

  (
    g535_n,
    g527_p_spl_0,
    g534_p_spl_0
  );


  and

  (
    g536_p,
    g527_p_spl_0,
    g534_p_spl_0
  );


  or

  (
    g536_n,
    g527_n_spl_0,
    g534_n_spl_0
  );


  and

  (
    g537_p,
    g535_n,
    g536_n
  );


  or

  (
    g537_n,
    g535_p,
    g536_p
  );


  and

  (
    g538_p,
    g525_p,
    g537_n
  );


  and

  (
    g539_p,
    g525_n,
    g537_p
  );


  or

  (
    g540_n,
    g538_p,
    g539_p
  );


  and

  (
    g541_p,
    g74_n_spl_,
    g78_n_spl_
  );


  and

  (
    g542_p,
    g540_n,
    g541_p
  );


  and

  (
    g543_p,
    G10_n_spl_101,
    g326_n_spl_
  );


  or

  (
    g544_n,
    G7_p_spl_011,
    g543_p
  );


  or

  (
    g545_n,
    G7_n_spl_011,
    G9_n_spl_101
  );


  and

  (
    g546_p,
    g78_p_spl_,
    g545_n
  );


  and

  (
    g547_p,
    g544_n,
    g546_p
  );


  and

  (
    g548_p,
    G14_n_spl_100,
    g74_p
  );


  and

  (
    g549_p,
    g223_n_spl_,
    g548_p
  );


  or

  (
    g550_n,
    g547_p,
    g549_p
  );


  or

  (
    g551_n,
    g542_p,
    g550_n
  );


  and

  (
    g552_p,
    g202_n_spl_,
    g366_p_spl_100
  );


  or

  (
    g552_n,
    g202_p_spl_,
    g366_n_spl_100
  );


  and

  (
    g553_p,
    g217_n_spl_1,
    g552_n_spl_
  );


  or

  (
    g553_n,
    g217_p_spl_1,
    g552_p_spl_
  );


  and

  (
    g554_p,
    g217_p_spl_1,
    g552_p_spl_
  );


  or

  (
    g554_n,
    g217_n_spl_1,
    g552_n_spl_
  );


  and

  (
    g555_p,
    g553_n,
    g554_n
  );


  or

  (
    g555_n,
    g553_p,
    g554_p
  );


  and

  (
    g556_p,
    g390_p_spl_0,
    g555_p_spl_0
  );


  or

  (
    g556_n,
    g390_n_spl_0,
    g555_n_spl_0
  );


  and

  (
    g557_p,
    G11_p_spl_101,
    g394_n_spl_01
  );


  or

  (
    g557_n,
    G11_n_spl_10,
    g394_p_spl_01
  );


  and

  (
    g558_p,
    g393_p_spl_010,
    g557_n
  );


  or

  (
    g558_n,
    g393_n_spl_010,
    g557_p
  );


  and

  (
    g559_p,
    g385_p_spl_01,
    g558_n
  );


  or

  (
    g559_n,
    g385_n_spl_01,
    g558_p
  );


  and

  (
    g560_p,
    G41_p_spl_01,
    g409_n_spl_010
  );


  or

  (
    g560_n,
    G41_n_spl_01,
    g409_p_spl_010
  );


  and

  (
    g561_p,
    G42_p_spl_0,
    g406_n_spl_010
  );


  or

  (
    g561_n,
    G42_n_spl_0,
    g406_p_spl_010
  );


  and

  (
    g562_p,
    G4_p_spl_1011,
    g561_n
  );


  or

  (
    g562_n,
    G4_n_spl_1011,
    g561_p
  );


  and

  (
    g563_p,
    g560_n,
    g562_p
  );


  or

  (
    g563_n,
    g560_p,
    g562_n
  );


  and

  (
    g564_p,
    G13_n_spl_101,
    g423_n_spl_001
  );


  or

  (
    g564_n,
    G13_p_spl_110,
    g423_p_spl_001
  );


  and

  (
    g565_p,
    G14_n_spl_100,
    g425_n_spl_010
  );


  or

  (
    g565_n,
    G14_p_spl_100,
    g425_p_spl_010
  );


  and

  (
    g566_p,
    g564_n,
    g565_n
  );


  or

  (
    g566_n,
    g564_p,
    g565_p
  );


  and

  (
    g567_p,
    G39_n_spl_01,
    G43_n_spl_0
  );


  or

  (
    g567_n,
    G39_p_spl_01,
    G43_p_spl_0
  );


  and

  (
    g568_p,
    g412_n_spl_001,
    g567_n
  );


  or

  (
    g568_n,
    g412_p_spl_001,
    g567_p
  );


  and

  (
    g569_p,
    G12_p_spl_101,
    G40_n_spl_01
  );


  or

  (
    g569_n,
    G12_n_spl_101,
    G40_p_spl_01
  );


  and

  (
    g570_p,
    g414_n_spl_010,
    g569_n_spl_
  );


  or

  (
    g570_n,
    g414_p_spl_010,
    g569_p_spl_
  );


  and

  (
    g571_p,
    g568_n,
    g570_n
  );


  or

  (
    g571_n,
    g568_p,
    g570_p
  );


  and

  (
    g572_p,
    g566_p,
    g571_p
  );


  or

  (
    g572_n,
    g566_n,
    g571_n
  );


  and

  (
    g573_p,
    g563_p,
    g572_p
  );


  or

  (
    g573_n,
    g563_n,
    g572_n
  );


  and

  (
    g574_p,
    G8_n_spl_101,
    g425_n_spl_010
  );


  or

  (
    g574_n,
    G8_p_spl_101,
    g425_p_spl_010
  );


  and

  (
    g575_p,
    G7_n_spl_100,
    g412_n_spl_010
  );


  or

  (
    g575_n,
    G7_p_spl_100,
    g412_p_spl_010
  );


  and

  (
    g576_p,
    G10_n_spl_101,
    g414_n_spl_010
  );


  or

  (
    g576_n,
    G10_p_spl_101,
    g414_p_spl_010
  );


  and

  (
    g577_p,
    g575_n,
    g576_n
  );


  or

  (
    g577_n,
    g575_p,
    g576_p
  );


  and

  (
    g578_p,
    g574_n,
    g577_p
  );


  or

  (
    g578_n,
    g574_p,
    g577_n
  );


  and

  (
    g579_p,
    G9_n_spl_101,
    g423_n_spl_010
  );


  or

  (
    g579_n,
    G9_p_spl_101,
    g423_p_spl_010
  );


  and

  (
    g580_p,
    G20_p_spl_00,
    g406_n_spl_010
  );


  or

  (
    g580_n,
    G20_n_spl_00,
    g406_p_spl_010
  );


  and

  (
    g581_p,
    G21_p_spl_01,
    g409_n_spl_010
  );


  or

  (
    g581_n,
    G21_n_spl_01,
    g409_p_spl_010
  );


  and

  (
    g582_p,
    g580_n,
    g581_n
  );


  or

  (
    g582_n,
    g580_p,
    g581_p
  );


  and

  (
    g583_p,
    g579_n_spl_,
    g582_p
  );


  or

  (
    g583_n,
    g579_p_spl_,
    g582_n
  );


  and

  (
    g584_p,
    G19_p_spl_00,
    g412_n_spl_010
  );


  or

  (
    g584_n,
    G19_n_spl_00,
    g412_p_spl_010
  );


  and

  (
    g585_p,
    G22_p_spl_01,
    g414_n_spl_011
  );


  or

  (
    g585_n,
    G22_n_spl_01,
    g414_p_spl_011
  );


  and

  (
    g586_p,
    g584_n,
    g585_n
  );


  or

  (
    g586_n,
    g584_p,
    g585_p
  );


  and

  (
    g587_p,
    G4_n_spl_1100,
    g586_p
  );


  or

  (
    g587_n,
    G4_p_spl_1100,
    g586_n
  );


  and

  (
    g588_p,
    g583_p,
    g587_p
  );


  or

  (
    g588_n,
    g583_n,
    g587_n
  );


  and

  (
    g589_p,
    g578_p,
    g588_p
  );


  or

  (
    g589_n,
    g578_n,
    g588_n
  );


  and

  (
    g590_p,
    g573_n,
    g589_n
  );


  or

  (
    g590_n,
    g573_p,
    g589_p
  );


  and

  (
    g591_p,
    g393_n_spl_010,
    g590_n
  );


  or

  (
    g591_n,
    g393_p_spl_010,
    g590_p
  );


  and

  (
    g592_p,
    g559_p,
    g591_n
  );


  or

  (
    g592_n,
    g559_n,
    g591_p
  );


  and

  (
    g593_p,
    g556_n,
    g592_p
  );


  or

  (
    g593_n,
    g556_p,
    g592_n
  );


  and

  (
    g594_p,
    g229_n_spl_,
    g366_p_spl_101
  );


  or

  (
    g594_n,
    g229_p_spl_,
    g366_n_spl_101
  );


  and

  (
    g595_p,
    g243_n_spl_0,
    g594_n_spl_
  );


  or

  (
    g595_n,
    g243_p_spl_0,
    g594_p_spl_
  );


  and

  (
    g596_p,
    g243_p_spl_,
    g594_p_spl_
  );


  or

  (
    g596_n,
    g243_n_spl_,
    g594_n_spl_
  );


  and

  (
    g597_p,
    g595_n,
    g596_n
  );


  or

  (
    g597_n,
    g595_p,
    g596_p
  );


  and

  (
    g598_p,
    g376_p_spl_0,
    g597_n_spl_00
  );


  or

  (
    g598_n,
    g376_n_spl_,
    g597_p_spl_00
  );


  and

  (
    g599_p,
    g242_p_spl_,
    g366_n_spl_101
  );


  or

  (
    g599_n,
    g242_n_spl_,
    g366_p_spl_101
  );


  and

  (
    g600_p,
    g167_p_spl_,
    g366_n_spl_11
  );


  or

  (
    g600_n,
    g167_n_spl_,
    g366_p_spl_11
  );


  and

  (
    g601_p,
    g370_n_spl_0,
    g600_n_spl_
  );


  or

  (
    g601_n,
    g370_p_spl_0,
    g600_p_spl_
  );


  and

  (
    g602_p,
    g190_p_spl_,
    g366_n_spl_11
  );


  or

  (
    g602_n,
    g190_n_spl_,
    g366_p_spl_11
  );


  and

  (
    g603_p,
    g601_n_spl_,
    g602_n
  );


  or

  (
    g603_n,
    g601_p_spl_,
    g602_p
  );


  and

  (
    g604_p,
    g597_n_spl_00,
    g603_n_spl_
  );


  or

  (
    g604_n,
    g597_p_spl_00,
    g603_p_spl_
  );


  and

  (
    g605_p,
    g599_n,
    g604_n
  );


  or

  (
    g605_n,
    g599_p,
    g604_p
  );


  and

  (
    g606_p,
    g555_n_spl_0,
    g605_p_spl_
  );


  or

  (
    g606_n,
    g555_p_spl_0,
    g605_n_spl_
  );


  and

  (
    g607_p,
    g555_p_spl_,
    g605_n_spl_
  );


  or

  (
    g607_n,
    g555_n_spl_,
    g605_p_spl_
  );


  and

  (
    g608_p,
    g606_n,
    g607_n
  );


  or

  (
    g608_n,
    g606_p,
    g607_p
  );


  and

  (
    g609_p,
    g598_n_spl_,
    g608_n_spl_
  );


  or

  (
    g609_n,
    g598_p_spl_,
    g608_p_spl_
  );


  and

  (
    g610_p,
    g598_p_spl_,
    g608_p_spl_
  );


  or

  (
    g610_n,
    g598_n_spl_,
    g608_n_spl_
  );


  and

  (
    g611_p,
    g609_n,
    g610_n
  );


  or

  (
    g611_n,
    g609_p,
    g610_p
  );


  and

  (
    g612_p,
    g370_p_spl_1,
    g600_p_spl_
  );


  or

  (
    g612_n,
    g370_n_spl_1,
    g600_n_spl_
  );


  and

  (
    g613_p,
    g601_n_spl_,
    g612_n
  );


  or

  (
    g613_n,
    g601_p_spl_,
    g612_p
  );


  and

  (
    g614_p,
    g387_n_spl_0,
    g613_n_spl_
  );


  or

  (
    g614_n,
    g387_p_spl_0,
    g613_p_spl_
  );


  and

  (
    g615_p,
    g387_p_spl_,
    g613_p_spl_
  );


  or

  (
    g615_n,
    g387_n_spl_,
    g613_n_spl_
  );


  and

  (
    g616_p,
    g614_n,
    g615_n
  );


  or

  (
    g616_n,
    g614_p,
    g615_p
  );


  and

  (
    g617_p,
    g376_n_spl_,
    g603_n_spl_
  );


  or

  (
    g617_n,
    g376_p_spl_0,
    g603_p_spl_
  );


  and

  (
    g618_p,
    g597_p_spl_0,
    g617_p_spl_
  );


  or

  (
    g618_n,
    g597_n_spl_0,
    g617_n_spl_
  );


  and

  (
    g619_p,
    g597_n_spl_1,
    g617_n_spl_
  );


  or

  (
    g619_n,
    g597_p_spl_1,
    g617_p_spl_
  );


  and

  (
    g620_p,
    g618_n,
    g619_n
  );


  or

  (
    g620_n,
    g618_p,
    g619_p
  );


  and

  (
    g621_p,
    g616_n_spl_0,
    g620_n_spl_0
  );


  or

  (
    g621_n,
    g616_p_spl_0,
    g620_p_spl_0
  );


  and

  (
    g622_p,
    g379_p_spl_10,
    g621_n
  );


  or

  (
    g622_n,
    g379_n_spl_01,
    g621_p
  );


  and

  (
    g623_p,
    g377_n_spl_01,
    g622_n
  );


  or

  (
    g623_n,
    g377_p_spl_00,
    g622_p
  );


  and

  (
    g624_p,
    g384_p_spl_00,
    g623_n
  );


  or

  (
    g624_n,
    g384_n_spl_00,
    g623_p
  );


  and

  (
    g625_p,
    g611_n,
    g624_n
  );


  or

  (
    g625_n,
    g611_p,
    g624_p
  );


  and

  (
    g626_p,
    g593_n,
    g625_n
  );


  or

  (
    g626_n,
    g593_p,
    g625_p
  );


  and

  (
    g627_p,
    g379_p_spl_10,
    g616_p_spl_0
  );


  or

  (
    g627_n,
    g379_n_spl_1,
    g616_n_spl_0
  );


  and

  (
    g628_p,
    g379_n_spl_1,
    g616_n_spl_1
  );


  or

  (
    g628_n,
    g379_p_spl_1,
    g616_p_spl_1
  );


  and

  (
    g629_p,
    g627_n,
    g628_n_spl_0
  );


  or

  (
    g629_n,
    g627_p,
    g628_p_spl_0
  );


  and

  (
    g630_p,
    g377_n_spl_01,
    g629_p
  );


  or

  (
    g630_n,
    g377_p_spl_01,
    g629_n
  );


  and

  (
    g631_p,
    g384_n_spl_01,
    g616_n_spl_1
  );


  or

  (
    g631_n,
    g384_p_spl_01,
    g616_p_spl_1
  );


  and

  (
    g632_p,
    G39_p_spl_01,
    g423_n_spl_010
  );


  or

  (
    g632_n,
    G39_n_spl_01,
    g423_p_spl_010
  );


  and

  (
    g633_p,
    G40_p_spl_10,
    g425_n_spl_011
  );


  or

  (
    g633_n,
    G40_n_spl_10,
    g425_p_spl_011
  );


  and

  (
    g634_p,
    g632_n,
    g633_n
  );


  or

  (
    g634_n,
    g632_p,
    g633_p
  );


  and

  (
    g635_p,
    G43_p_spl_1,
    g409_n_spl_011
  );


  or

  (
    g635_n,
    G43_n_spl_1,
    g409_p_spl_011
  );


  and

  (
    g636_p,
    G44_p_spl_0,
    g406_n_spl_011
  );


  or

  (
    g636_n,
    G44_n_spl_0,
    g406_p_spl_011
  );


  and

  (
    g637_p,
    G4_p_spl_1100,
    g636_n
  );


  or

  (
    g637_n,
    G4_n_spl_1100,
    g636_p
  );


  and

  (
    g638_p,
    g635_n,
    g637_p
  );


  or

  (
    g638_n,
    g635_p,
    g637_n
  );


  and

  (
    g639_p,
    g634_p,
    g638_p
  );


  or

  (
    g639_n,
    g634_n,
    g638_n
  );


  and

  (
    g640_p,
    G41_n_spl_10,
    G45_n_spl_
  );


  or

  (
    g640_n,
    G41_p_spl_10,
    G45_p_spl_
  );


  and

  (
    g641_p,
    g412_n_spl_011,
    g640_n
  );


  or

  (
    g641_n,
    g412_p_spl_011,
    g640_p
  );


  and

  (
    g642_p,
    G14_p_spl_101,
    G42_n_spl_1
  );


  or

  (
    g642_n,
    G14_n_spl_101,
    G42_p_spl_1
  );


  and

  (
    g643_p,
    g414_n_spl_011,
    g642_n
  );


  or

  (
    g643_n,
    g414_p_spl_011,
    g642_p
  );


  and

  (
    g644_p,
    g641_n,
    g643_n
  );


  or

  (
    g644_n,
    g641_p,
    g643_p
  );


  and

  (
    g645_p,
    g639_p,
    g644_p
  );


  or

  (
    g645_n,
    g639_n,
    g644_n
  );


  and

  (
    g646_p,
    G12_n_spl_101,
    g414_n_spl_100
  );


  or

  (
    g646_n,
    G12_p_spl_110,
    g414_p_spl_100
  );


  and

  (
    g647_p,
    G10_n_spl_110,
    g425_n_spl_011
  );


  or

  (
    g647_n,
    G10_p_spl_101,
    g425_p_spl_011
  );


  and

  (
    g648_p,
    g646_n,
    g647_n
  );


  or

  (
    g648_n,
    g646_p,
    g647_p
  );


  and

  (
    g649_p,
    G4_n_spl_1101,
    g648_p
  );


  or

  (
    g649_n,
    G4_p_spl_1101,
    g648_n
  );


  and

  (
    g650_p,
    G22_p_spl_01,
    g406_n_spl_011
  );


  or

  (
    g650_n,
    G22_n_spl_01,
    g406_p_spl_011
  );


  and

  (
    g651_p,
    G7_n_spl_100,
    g409_n_spl_011
  );


  or

  (
    g651_n,
    G7_p_spl_100,
    g409_p_spl_011
  );


  and

  (
    g652_p,
    g650_n,
    g651_n
  );


  or

  (
    g652_n,
    g650_p,
    g651_p
  );


  and

  (
    g653_p,
    G8_n_spl_101,
    g414_n_spl_100
  );


  or

  (
    g653_n,
    G8_p_spl_110,
    g414_p_spl_100
  );


  and

  (
    g654_p,
    G11_n_spl_11,
    g423_n_spl_011
  );


  or

  (
    g654_n,
    G11_p_spl_11,
    g423_p_spl_011
  );


  and

  (
    g655_p,
    g653_n_spl_,
    g654_n_spl_
  );


  or

  (
    g655_n,
    g653_p_spl_,
    g654_p_spl_
  );


  and

  (
    g656_p,
    G9_p_spl_110,
    G21_n_spl_01
  );


  or

  (
    g656_n,
    G9_n_spl_110,
    G21_p_spl_01
  );


  and

  (
    g657_p,
    g412_n_spl_011,
    g656_n
  );


  or

  (
    g657_n,
    g412_p_spl_011,
    g656_p
  );


  and

  (
    g658_p,
    g655_p,
    g657_n
  );


  or

  (
    g658_n,
    g655_n,
    g657_p
  );


  and

  (
    g659_p,
    g652_p,
    g658_p
  );


  or

  (
    g659_n,
    g652_n,
    g658_n
  );


  and

  (
    g660_p,
    g649_p_spl_,
    g659_p
  );


  or

  (
    g660_n,
    g649_n_spl_,
    g659_n
  );


  and

  (
    g661_p,
    g645_n,
    g660_n
  );


  or

  (
    g661_n,
    g645_p,
    g660_p
  );


  and

  (
    g662_p,
    g393_n_spl_011,
    g661_n
  );


  or

  (
    g662_n,
    g393_p_spl_011,
    g661_p
  );


  and

  (
    g663_p,
    G6_n_spl_10,
    g102_p_spl_
  );


  or

  (
    g663_n,
    G6_p_spl_10,
    g102_n_spl_
  );


  and

  (
    g664_p,
    G7_n_spl_101,
    G8_p_spl_110
  );


  or

  (
    g664_n,
    G7_p_spl_101,
    G8_n_spl_110
  );


  and

  (
    g665_p,
    g117_n_spl_,
    g664_p
  );


  or

  (
    g665_n,
    g117_p_spl_,
    g664_n
  );


  and

  (
    g666_p,
    G6_p_spl_1,
    g665_p
  );


  or

  (
    g666_n,
    G6_n_spl_1,
    g665_n
  );


  and

  (
    g667_p,
    g663_n,
    g666_n
  );


  or

  (
    g667_n,
    g663_p,
    g666_p
  );


  and

  (
    g668_p,
    g196_p_spl_,
    g667_n
  );


  or

  (
    g668_n,
    g196_n_spl_,
    g667_p
  );


  and

  (
    g669_p,
    G14_n_spl_101,
    g668_p
  );


  or

  (
    g669_n,
    G14_p_spl_101,
    g668_n
  );


  and

  (
    g670_p,
    g394_p_spl_01,
    g669_p
  );


  or

  (
    g670_n,
    g394_n_spl_01,
    g669_n
  );


  and

  (
    g671_p,
    G13_p_spl_110,
    g394_n_spl_1
  );


  or

  (
    g671_n,
    G13_n_spl_110,
    g394_p_spl_1
  );


  and

  (
    g672_p,
    g670_n,
    g671_n
  );


  or

  (
    g672_n,
    g670_p,
    g671_p
  );


  and

  (
    g673_p,
    g393_p_spl_011,
    g672_p
  );


  or

  (
    g673_n,
    g393_n_spl_011,
    g672_n
  );


  and

  (
    g674_p,
    g370_p_spl_1,
    g390_p_spl_1
  );


  or

  (
    g674_n,
    g370_n_spl_1,
    g390_n_spl_1
  );


  and

  (
    g675_p,
    g385_p_spl_01,
    g674_n
  );


  or

  (
    g675_n,
    g385_n_spl_01,
    g674_p
  );


  and

  (
    g676_p,
    g673_n,
    g675_p
  );


  or

  (
    g676_n,
    g673_p,
    g675_n
  );


  and

  (
    g677_p,
    g662_n,
    g676_p
  );


  or

  (
    g677_n,
    g662_p,
    g676_n
  );


  and

  (
    g678_p,
    g631_n,
    g677_n
  );


  or

  (
    g678_n,
    g631_p,
    g677_p
  );


  and

  (
    g679_p,
    g630_n,
    g678_p
  );


  or

  (
    g679_n,
    g630_p,
    g678_n
  );


  and

  (
    g680_p,
    g620_p_spl_0,
    g628_n_spl_0
  );


  or

  (
    g680_n,
    g620_n_spl_0,
    g628_p_spl_0
  );


  and

  (
    g681_p,
    g620_n_spl_1,
    g628_p_spl_
  );


  or

  (
    g681_n,
    g620_p_spl_1,
    g628_n_spl_
  );


  and

  (
    g682_p,
    g680_n,
    g681_n
  );


  or

  (
    g682_n,
    g680_p,
    g681_p
  );


  and

  (
    g683_p,
    g377_n_spl_10,
    g682_n
  );


  or

  (
    g683_n,
    g377_p_spl_01,
    g682_p
  );


  and

  (
    g684_p,
    g384_n_spl_01,
    g620_n_spl_1
  );


  or

  (
    g684_n,
    g384_p_spl_01,
    g620_p_spl_1
  );


  and

  (
    g685_p,
    G4_p_spl_1101,
    g432_n_spl_
  );


  or

  (
    g685_n,
    G4_n_spl_1101,
    g432_p_spl_
  );


  and

  (
    g686_p,
    G43_p_spl_1,
    g406_n_spl_100
  );


  or

  (
    g686_n,
    G43_n_spl_1,
    g406_p_spl_100
  );


  and

  (
    g687_p,
    g685_p_spl_,
    g686_n
  );


  or

  (
    g687_n,
    g685_n_spl_,
    g686_p
  );


  and

  (
    g688_p,
    G14_n_spl_110,
    g423_n_spl_011
  );


  or

  (
    g688_n,
    G14_p_spl_110,
    g423_p_spl_011
  );


  and

  (
    g689_p,
    G41_p_spl_10,
    g414_n_spl_101
  );


  or

  (
    g689_n,
    G41_n_spl_10,
    g414_p_spl_101
  );


  and

  (
    g690_p,
    G42_p_spl_1,
    g409_n_spl_100
  );


  or

  (
    g690_n,
    G42_n_spl_1,
    g409_p_spl_100
  );


  and

  (
    g691_p,
    g689_n,
    g690_n
  );


  or

  (
    g691_n,
    g689_p,
    g690_p
  );


  and

  (
    g692_p,
    g688_n,
    g691_p
  );


  or

  (
    g692_n,
    g688_p,
    g691_n
  );


  and

  (
    g693_p,
    g687_p,
    g692_p
  );


  or

  (
    g693_n,
    g687_n,
    g692_n
  );


  and

  (
    g694_p,
    G39_p_spl_10,
    g425_n_spl_100
  );


  or

  (
    g694_n,
    G39_n_spl_10,
    g425_p_spl_100
  );


  and

  (
    g695_p,
    G40_n_spl_10,
    G44_n_spl_
  );


  or

  (
    g695_n,
    G40_p_spl_10,
    G44_p_spl_
  );


  and

  (
    g696_p,
    g412_n_spl_100,
    g695_n
  );


  or

  (
    g696_n,
    g412_p_spl_100,
    g695_p
  );


  and

  (
    g697_p,
    g694_n,
    g696_n
  );


  or

  (
    g697_n,
    g694_p,
    g696_p
  );


  and

  (
    g698_p,
    g693_p,
    g697_p
  );


  or

  (
    g698_n,
    g693_n,
    g697_n
  );


  and

  (
    g699_p,
    G21_p_spl_10,
    g406_n_spl_100
  );


  or

  (
    g699_n,
    G21_n_spl_10,
    g406_p_spl_100
  );


  and

  (
    g700_p,
    G22_p_spl_10,
    g409_n_spl_100
  );


  or

  (
    g700_n,
    G22_n_spl_10,
    g409_p_spl_100
  );


  and

  (
    g701_p,
    g699_n,
    g700_n
  );


  or

  (
    g701_n,
    g699_p,
    g700_p
  );


  and

  (
    g702_p,
    G9_n_spl_110,
    g425_n_spl_100
  );


  or

  (
    g702_n,
    G9_p_spl_110,
    g425_p_spl_100
  );


  and

  (
    g703_p,
    G4_n_spl_1110,
    g702_n
  );


  or

  (
    g703_n,
    G4_p_spl_1110,
    g702_p
  );


  and

  (
    g704_p,
    g701_p,
    g703_p
  );


  or

  (
    g704_n,
    g701_n,
    g703_n
  );


  and

  (
    g705_p,
    G10_n_spl_110,
    g423_n_spl_10
  );


  or

  (
    g705_n,
    G10_p_spl_11,
    g423_p_spl_10
  );


  and

  (
    g706_p,
    G8_p_spl_111,
    G20_n_spl_0
  );


  or

  (
    g706_n,
    G8_n_spl_110,
    G20_p_spl_0
  );


  and

  (
    g707_p,
    g412_n_spl_100,
    g706_n_spl_
  );


  or

  (
    g707_n,
    g412_p_spl_100,
    g706_p_spl_
  );


  and

  (
    g708_p,
    g705_n_spl_,
    g707_n
  );


  or

  (
    g708_n,
    g705_p_spl_,
    g707_p
  );


  and

  (
    g709_p,
    G7_n_spl_101,
    g414_n_spl_101
  );


  or

  (
    g709_n,
    G7_p_spl_101,
    g414_p_spl_101
  );


  and

  (
    g710_p,
    g480_n_spl_,
    g709_n
  );


  or

  (
    g710_n,
    g480_p_spl_,
    g709_p
  );


  and

  (
    g711_p,
    g708_p,
    g710_p
  );


  or

  (
    g711_n,
    g708_n,
    g710_n
  );


  and

  (
    g712_p,
    g704_p,
    g711_p
  );


  or

  (
    g712_n,
    g704_n,
    g711_n
  );


  and

  (
    g713_p,
    g698_n,
    g712_n
  );


  or

  (
    g713_n,
    g698_p,
    g712_p
  );


  and

  (
    g714_p,
    g393_n_spl_100,
    g713_n
  );


  or

  (
    g714_n,
    g393_p_spl_100,
    g713_p
  );


  and

  (
    g715_p,
    g390_p_spl_1,
    g597_p_spl_1
  );


  or

  (
    g715_n,
    g390_n_spl_1,
    g597_n_spl_1
  );


  and

  (
    g716_p,
    G12_p_spl_110,
    g394_n_spl_1
  );


  or

  (
    g716_n,
    G12_n_spl_11,
    g394_p_spl_1
  );


  and

  (
    g717_p,
    g393_p_spl_100,
    g716_n
  );


  or

  (
    g717_n,
    g393_n_spl_100,
    g716_p
  );


  and

  (
    g718_p,
    g385_p_spl_10,
    g717_n
  );


  or

  (
    g718_n,
    g385_n_spl_10,
    g717_p
  );


  and

  (
    g719_p,
    g715_n,
    g718_p
  );


  or

  (
    g719_n,
    g715_p,
    g718_n
  );


  and

  (
    g720_p,
    g714_n,
    g719_p
  );


  or

  (
    g720_n,
    g714_p,
    g719_n
  );


  and

  (
    g721_p,
    g684_n,
    g720_n
  );


  or

  (
    g721_n,
    g684_p,
    g720_p
  );


  and

  (
    g722_p,
    g683_n,
    g721_p
  );


  or

  (
    g722_n,
    g683_p,
    g721_n
  );


  and

  (
    g723_p,
    G47_p_spl_10,
    g519_p_spl_
  );


  or

  (
    g723_n,
    G47_n_spl_10,
    g519_n_spl_
  );


  and

  (
    g724_p,
    g513_p_spl_00,
    g723_p_spl_
  );


  or

  (
    g724_n,
    g513_n_spl_00,
    g723_n_spl_
  );


  and

  (
    g725_p,
    g513_p_spl_0,
    g530_n_spl_0
  );


  or

  (
    g725_n,
    g513_n_spl_0,
    g530_p_spl_0
  );


  and

  (
    g726_p,
    g528_n_spl_,
    g725_n
  );


  or

  (
    g726_n,
    g528_p_spl_,
    g725_p
  );


  and

  (
    g727_p,
    g517_p_spl_0,
    g726_p_spl_
  );


  or

  (
    g727_n,
    g517_n_spl_0,
    g726_n_spl_
  );


  and

  (
    g728_p,
    g517_n_spl_1,
    g726_n_spl_
  );


  or

  (
    g728_n,
    g517_p_spl_1,
    g726_p_spl_
  );


  and

  (
    g729_p,
    g727_n,
    g728_n
  );


  or

  (
    g729_n,
    g727_p,
    g728_p
  );


  and

  (
    g730_p,
    g724_p_spl_0,
    g729_p_spl_
  );


  or

  (
    g730_n,
    g724_n_spl_0,
    g729_n_spl_
  );


  and

  (
    g731_p,
    g724_n_spl_0,
    g729_n_spl_
  );


  or

  (
    g731_n,
    g724_p_spl_0,
    g729_p_spl_
  );


  and

  (
    g732_p,
    g730_n_spl_0,
    g731_n
  );


  or

  (
    g732_n,
    g730_p_spl_0,
    g731_p
  );


  and

  (
    g733_p,
    g503_n_spl_,
    g530_n_spl_
  );


  or

  (
    g733_n,
    g503_p_spl_,
    g530_p_spl_
  );


  and

  (
    g734_p,
    g513_n_spl_1,
    g723_n_spl_
  );


  or

  (
    g734_n,
    g513_p_spl_1,
    g723_p_spl_
  );


  and

  (
    g735_p,
    g724_n_spl_,
    g734_n
  );


  or

  (
    g735_n,
    g724_p_spl_,
    g734_p
  );


  and

  (
    g736_p,
    g733_p_spl_,
    g735_n_spl_
  );


  or

  (
    g736_n,
    g733_n_spl_,
    g735_p_spl_
  );


  and

  (
    g737_p,
    g733_n_spl_,
    g735_p_spl_
  );


  or

  (
    g737_n,
    g733_p_spl_,
    g735_n_spl_
  );


  and

  (
    g738_p,
    g736_n,
    g737_n
  );


  or

  (
    g738_n,
    g736_p,
    g737_p
  );


  and

  (
    g739_p,
    G47_p_spl_1,
    g527_n_spl_
  );


  or

  (
    g739_n,
    G47_n_spl_1,
    g527_p_spl_
  );


  and

  (
    g740_p,
    g521_p_spl_,
    g739_p
  );


  or

  (
    g740_n,
    g521_n_spl_,
    g739_n
  );


  and

  (
    g741_p,
    g738_n_spl_0,
    g740_n_spl_0
  );


  or

  (
    g741_n,
    g738_p_spl_0,
    g740_p_spl_0
  );


  and

  (
    g742_p,
    g732_p_spl_0,
    g741_n_spl_0
  );


  or

  (
    g742_n,
    g732_n_spl_0,
    g741_p_spl_0
  );


  and

  (
    g743_p,
    g732_n_spl_0,
    g741_p_spl_0
  );


  or

  (
    g743_n,
    g732_p_spl_0,
    g741_n_spl_0
  );


  and

  (
    g744_p,
    g742_n,
    g743_n
  );


  or

  (
    g744_n,
    g742_p,
    g743_p
  );


  and

  (
    g745_p,
    g377_n_spl_10,
    g744_n
  );


  or

  (
    g745_n,
    g377_p_spl_10,
    g744_p
  );


  and

  (
    g746_p,
    g452_p_spl_0,
    g517_p_spl_1
  );


  or

  (
    g746_n,
    g452_n_spl_0,
    g517_n_spl_1
  );


  and

  (
    g747_p,
    G8_n_spl_11,
    g393_p_spl_101
  );


  or

  (
    g747_n,
    G8_p_spl_111,
    g393_n_spl_101
  );


  and

  (
    g748_p,
    g385_p_spl_10,
    g747_n
  );


  or

  (
    g748_n,
    g385_n_spl_10,
    g747_p
  );


  and

  (
    g749_p,
    g430_n_spl_,
    g438_n_spl_
  );


  or

  (
    g749_n,
    g430_p_spl_,
    g438_p_spl_
  );


  and

  (
    g750_p,
    G39_p_spl_10,
    g406_n_spl_101
  );


  or

  (
    g750_n,
    G39_n_spl_10,
    g406_p_spl_101
  );


  and

  (
    g751_p,
    G14_n_spl_110,
    g409_n_spl_101
  );


  or

  (
    g751_n,
    G14_p_spl_110,
    g409_p_spl_101
  );


  and

  (
    g752_p,
    g750_n,
    g751_n
  );


  or

  (
    g752_n,
    g750_p,
    g751_p
  );


  and

  (
    g753_p,
    g705_n_spl_,
    g752_p
  );


  or

  (
    g753_n,
    g705_p_spl_,
    g752_n
  );


  and

  (
    g754_p,
    g412_n_spl_101,
    g569_n_spl_
  );


  or

  (
    g754_n,
    g412_p_spl_101,
    g569_p_spl_
  );


  and

  (
    g755_p,
    g685_p_spl_,
    g754_n
  );


  or

  (
    g755_n,
    g685_n_spl_,
    g754_p
  );


  and

  (
    g756_p,
    g753_p,
    g755_p
  );


  or

  (
    g756_n,
    g753_n,
    g755_n
  );


  and

  (
    g757_p,
    g749_p,
    g756_p
  );


  or

  (
    g757_n,
    g749_n,
    g756_n
  );


  and

  (
    g758_p,
    G21_p_spl_10,
    g425_n_spl_101
  );


  or

  (
    g758_n,
    G21_n_spl_10,
    g425_p_spl_101
  );


  and

  (
    g759_p,
    G17_p_spl_0,
    g406_n_spl_101
  );


  or

  (
    g759_n,
    G17_n_spl_0,
    g406_p_spl_101
  );


  and

  (
    g760_p,
    g758_n,
    g759_n
  );


  or

  (
    g760_n,
    g758_p,
    g759_p
  );


  and

  (
    g761_p,
    G22_p_spl_10,
    g423_n_spl_10
  );


  or

  (
    g761_n,
    G22_n_spl_10,
    g423_p_spl_10
  );


  and

  (
    g762_p,
    G4_n_spl_1110,
    g761_n
  );


  or

  (
    g762_n,
    G4_p_spl_1110,
    g761_p
  );


  and

  (
    g763_p,
    G18_p_spl_0,
    g409_n_spl_101
  );


  or

  (
    g763_n,
    G18_n_spl_0,
    g409_p_spl_101
  );


  and

  (
    g764_p,
    G16_n_spl_,
    G20_n_spl_1
  );


  or

  (
    g764_n,
    G16_p_spl_,
    G20_p_spl_1
  );


  and

  (
    g765_p,
    g412_n_spl_101,
    g764_n
  );


  or

  (
    g765_n,
    g412_p_spl_101,
    g764_p
  );


  and

  (
    g766_p,
    G7_p_spl_110,
    G19_n_spl_0
  );


  or

  (
    g766_n,
    G7_n_spl_110,
    G19_p_spl_0
  );


  and

  (
    g767_p,
    g414_n_spl_110,
    g766_n
  );


  or

  (
    g767_n,
    g414_p_spl_110,
    g766_p
  );


  and

  (
    g768_p,
    g765_n,
    g767_n
  );


  or

  (
    g768_n,
    g765_p,
    g767_p
  );


  and

  (
    g769_p,
    g763_n,
    g768_p
  );


  or

  (
    g769_n,
    g763_p,
    g768_n
  );


  and

  (
    g770_p,
    g762_p,
    g769_p
  );


  or

  (
    g770_n,
    g762_n,
    g769_n
  );


  and

  (
    g771_p,
    g760_p,
    g770_p
  );


  or

  (
    g771_n,
    g760_n,
    g770_n
  );


  and

  (
    g772_p,
    g757_n,
    g771_n
  );


  or

  (
    g772_n,
    g757_p,
    g771_p
  );


  and

  (
    g773_p,
    g393_n_spl_101,
    g772_n
  );


  or

  (
    g773_n,
    g393_p_spl_101,
    g772_p
  );


  and

  (
    g774_p,
    g748_p,
    g773_n
  );


  or

  (
    g774_n,
    g748_n,
    g773_p
  );


  and

  (
    g775_p,
    g746_n,
    g774_p
  );


  or

  (
    g775_n,
    g746_p,
    g774_n
  );


  and

  (
    g776_p,
    g384_n_spl_10,
    g732_n_spl_1
  );


  or

  (
    g776_n,
    g384_p_spl_10,
    g732_p_spl_1
  );


  and

  (
    g777_p,
    g775_n,
    g776_n
  );


  or

  (
    g777_n,
    g775_p,
    g776_p
  );


  and

  (
    g778_p,
    g745_n,
    g777_p
  );


  or

  (
    g778_n,
    g745_p,
    g777_n
  );


  and

  (
    g779_p,
    g306_n_spl_,
    g365_p_spl_1
  );


  or

  (
    g779_n,
    g306_p_spl_,
    g365_n_spl_1
  );


  and

  (
    g780_p,
    g320_n_spl_1,
    g779_n_spl_
  );


  or

  (
    g780_n,
    g320_p_spl_1,
    g779_p_spl_
  );


  and

  (
    g781_p,
    g320_p_spl_1,
    g779_p_spl_
  );


  or

  (
    g781_n,
    g320_n_spl_1,
    g779_n_spl_
  );


  and

  (
    g782_p,
    g780_n,
    g781_n
  );


  or

  (
    g782_n,
    g780_p,
    g781_p
  );


  and

  (
    g783_p,
    g452_p_spl_1,
    g782_p_spl_0
  );


  or

  (
    g783_n,
    g452_n_spl_1,
    g782_n_spl_0
  );


  and

  (
    g784_p,
    G11_p_spl_11,
    G39_n_spl_11
  );


  or

  (
    g784_n,
    G11_n_spl_11,
    G39_p_spl_11
  );


  and

  (
    g785_p,
    g412_n_spl_110,
    g784_n
  );


  or

  (
    g785_n,
    g412_p_spl_110,
    g784_p
  );


  and

  (
    g786_p,
    G5_p_spl_1,
    g579_n_spl_
  );


  or

  (
    g786_n,
    G5_n_spl_1,
    g579_p_spl_
  );


  and

  (
    g787_p,
    g649_p_spl_,
    g786_p
  );


  or

  (
    g787_n,
    g649_n_spl_,
    g786_n
  );


  and

  (
    g788_p,
    G14_n_spl_111,
    g406_n_spl_110
  );


  or

  (
    g788_n,
    G14_p_spl_111,
    g406_p_spl_110
  );


  and

  (
    g789_p,
    G13_n_spl_110,
    g409_n_spl_110
  );


  or

  (
    g789_n,
    G13_p_spl_111,
    g409_p_spl_110
  );


  and

  (
    g790_p,
    g788_n,
    g789_n
  );


  or

  (
    g790_n,
    g788_p,
    g789_p
  );


  and

  (
    g791_p,
    g653_n_spl_,
    g790_p
  );


  or

  (
    g791_n,
    g653_p_spl_,
    g790_n
  );


  and

  (
    g792_p,
    g787_p,
    g791_p
  );


  or

  (
    g792_n,
    g787_n,
    g791_n
  );


  and

  (
    g793_p,
    g785_n,
    g792_p
  );


  or

  (
    g793_n,
    g785_p,
    g792_n
  );


  and

  (
    g794_p,
    G5_n_spl_1,
    G7_n_spl_110
  );


  or

  (
    g794_n,
    G5_p_spl_1,
    G7_p_spl_110
  );


  and

  (
    g795_p,
    G17_p_spl_0,
    g409_n_spl_110
  );


  or

  (
    g795_n,
    G17_n_spl_0,
    g409_p_spl_110
  );


  and

  (
    g796_p,
    G15_n,
    G19_n_spl_1
  );


  or

  (
    g796_n,
    G15_p,
    G19_p_spl_1
  );


  and

  (
    g797_p,
    g412_n_spl_110,
    g796_n
  );


  or

  (
    g797_n,
    g412_p_spl_110,
    g796_p
  );


  and

  (
    g798_p,
    G18_n_spl_1,
    G22_n_spl_11
  );


  or

  (
    g798_n,
    G18_p_spl_1,
    G22_p_spl_11
  );


  and

  (
    g799_p,
    g414_n_spl_110,
    g798_n
  );


  or

  (
    g799_n,
    g414_p_spl_110,
    g798_p
  );


  and

  (
    g800_p,
    g797_n,
    g799_n
  );


  or

  (
    g800_n,
    g797_p,
    g799_p
  );


  and

  (
    g801_p,
    g795_n,
    g800_p
  );


  or

  (
    g801_n,
    g795_p,
    g800_n
  );


  and

  (
    g802_p,
    G21_p_spl_11,
    g423_n_spl_11
  );


  or

  (
    g802_n,
    G21_n_spl_11,
    g423_p_spl_11
  );


  and

  (
    g803_p,
    g146_p_spl_,
    g802_n
  );


  or

  (
    g803_n,
    g146_n_spl_,
    g802_p
  );


  and

  (
    g804_p,
    G20_p_spl_1,
    g425_n_spl_101
  );


  or

  (
    g804_n,
    G20_n_spl_1,
    g425_p_spl_101
  );


  and

  (
    g805_p,
    G16_p_spl_,
    g406_n_spl_110
  );


  or

  (
    g805_n,
    G16_n_spl_,
    g406_p_spl_110
  );


  and

  (
    g806_p,
    g804_n,
    g805_n
  );


  or

  (
    g806_n,
    g804_p,
    g805_p
  );


  and

  (
    g807_p,
    g803_p,
    g806_p
  );


  or

  (
    g807_n,
    g803_n,
    g806_n
  );


  and

  (
    g808_p,
    g801_p,
    g807_p
  );


  or

  (
    g808_n,
    g801_n,
    g807_n
  );


  and

  (
    g809_p,
    g794_n,
    g808_n
  );


  or

  (
    g809_n,
    g794_p,
    g808_p
  );


  and

  (
    g810_p,
    g793_n,
    g809_p
  );


  or

  (
    g810_n,
    g793_p,
    g809_n
  );


  and

  (
    g811_p,
    g393_n_spl_110,
    g810_n
  );


  or

  (
    g811_n,
    g393_p_spl_110,
    g810_p
  );


  and

  (
    g812_p,
    G7_n_spl_111,
    g393_p_spl_110
  );


  or

  (
    g812_n,
    G7_p_spl_111,
    g393_n_spl_110
  );


  and

  (
    g813_p,
    g385_p_spl_11,
    g812_n
  );


  or

  (
    g813_n,
    g385_n_spl_11,
    g812_p
  );


  and

  (
    g814_p,
    g811_n,
    g813_p
  );


  or

  (
    g814_n,
    g811_p,
    g813_n
  );


  and

  (
    g815_p,
    g783_n,
    g814_p
  );


  or

  (
    g815_n,
    g783_p,
    g814_n
  );


  and

  (
    g816_p,
    g534_p_spl_1,
    g782_n_spl_0
  );


  or

  (
    g816_n,
    g534_n_spl_1,
    g782_p_spl_0
  );


  and

  (
    g817_p,
    g534_n_spl_1,
    g782_p_spl_
  );


  or

  (
    g817_n,
    g534_p_spl_1,
    g782_n_spl_
  );


  and

  (
    g818_p,
    g816_n,
    g817_n
  );


  or

  (
    g818_n,
    g816_p,
    g817_p
  );


  and

  (
    g819_p,
    g730_n_spl_0,
    g818_p_spl_
  );


  or

  (
    g819_n,
    g730_p_spl_0,
    g818_n_spl_
  );


  and

  (
    g820_p,
    g730_p_spl_,
    g818_n_spl_
  );


  or

  (
    g820_n,
    g730_n_spl_,
    g818_p_spl_
  );


  and

  (
    g821_p,
    g819_n,
    g820_n
  );


  or

  (
    g821_n,
    g819_p,
    g820_p
  );


  and

  (
    g822_p,
    g732_n_spl_1,
    g738_n_spl_0
  );


  or

  (
    g822_n,
    g732_p_spl_1,
    g738_p_spl_0
  );


  and

  (
    g823_p,
    g740_p_spl_0,
    g822_n
  );


  or

  (
    g823_n,
    g740_n_spl_0,
    g822_p
  );


  and

  (
    g824_p,
    g377_n_spl_11,
    g823_n
  );


  or

  (
    g824_n,
    g377_p_spl_10,
    g823_p
  );


  and

  (
    g825_p,
    g384_p_spl_10,
    g824_n
  );


  or

  (
    g825_n,
    g384_n_spl_10,
    g824_p
  );


  and

  (
    g826_p,
    g821_n,
    g825_n
  );


  or

  (
    g826_n,
    g821_p,
    g825_p
  );


  and

  (
    g827_p,
    g815_n,
    g826_n
  );


  or

  (
    g827_n,
    g815_p,
    g826_p
  );


  and

  (
    g828_p,
    g452_p_spl_1,
    g513_p_spl_1
  );


  or

  (
    g828_n,
    g452_n_spl_1,
    g513_n_spl_1
  );


  and

  (
    g829_p,
    G9_n_spl_11,
    g393_p_spl_111
  );


  or

  (
    g829_n,
    G9_p_spl_11,
    g393_n_spl_111
  );


  and

  (
    g830_p,
    g385_p_spl_11,
    g829_n
  );


  or

  (
    g830_n,
    g385_n_spl_11,
    g829_p
  );


  and

  (
    g831_p,
    G13_p_spl_111,
    G41_n_spl_1
  );


  or

  (
    g831_n,
    G13_n_spl_11,
    G41_p_spl_1
  );


  and

  (
    g832_p,
    g412_n_spl_111,
    g831_n
  );


  or

  (
    g832_n,
    g412_p_spl_111,
    g831_p
  );


  and

  (
    g833_p,
    G10_p_spl_11,
    G14_p_spl_111
  );


  or

  (
    g833_n,
    G10_n_spl_11,
    G14_n_spl_111
  );


  and

  (
    g834_p,
    g414_n_spl_111,
    g833_n
  );


  or

  (
    g834_n,
    g414_p_spl_111,
    g833_p
  );


  and

  (
    g835_p,
    g832_n,
    g834_n
  );


  or

  (
    g835_n,
    g832_p,
    g834_p
  );


  and

  (
    g836_p,
    g654_n_spl_,
    g835_p
  );


  or

  (
    g836_n,
    g654_p_spl_,
    g835_n
  );


  and

  (
    g837_p,
    G39_p_spl_11,
    g409_n_spl_111
  );


  or

  (
    g837_n,
    G39_n_spl_11,
    g409_p_spl_111
  );


  and

  (
    g838_p,
    G4_p_spl_1111,
    g837_n
  );


  or

  (
    g838_n,
    G4_n_spl_1111,
    g837_p
  );


  and

  (
    g839_p,
    G40_p_spl_1,
    g406_n_spl_111
  );


  or

  (
    g839_n,
    G40_n_spl_1,
    g406_p_spl_111
  );


  and

  (
    g840_p,
    G12_n_spl_11,
    g425_n_spl_11
  );


  or

  (
    g840_n,
    G12_p_spl_11,
    g425_p_spl_11
  );


  and

  (
    g841_p,
    g839_n,
    g840_n
  );


  or

  (
    g841_n,
    g839_p,
    g840_p
  );


  and

  (
    g842_p,
    g838_p,
    g841_p
  );


  or

  (
    g842_n,
    g838_n,
    g841_n
  );


  and

  (
    g843_p,
    g836_p,
    g842_p
  );


  or

  (
    g843_n,
    g836_n,
    g842_n
  );


  and

  (
    g844_p,
    G22_p_spl_11,
    g425_n_spl_11
  );


  or

  (
    g844_n,
    G22_n_spl_11,
    g425_p_spl_11
  );


  and

  (
    g845_p,
    G17_n_spl_,
    G21_n_spl_11
  );


  or

  (
    g845_n,
    G17_p_spl_,
    G21_p_spl_11
  );


  and

  (
    g846_p,
    g412_n_spl_111,
    g845_n
  );


  or

  (
    g846_n,
    g412_p_spl_111,
    g845_p
  );


  and

  (
    g847_p,
    g414_n_spl_111,
    g706_n_spl_
  );


  or

  (
    g847_n,
    g414_p_spl_111,
    g706_p_spl_
  );


  and

  (
    g848_p,
    g846_n,
    g847_n
  );


  or

  (
    g848_n,
    g846_p,
    g847_p
  );


  and

  (
    g849_p,
    g844_n,
    g848_p
  );


  or

  (
    g849_n,
    g844_p,
    g848_n
  );


  and

  (
    g850_p,
    G7_n_spl_111,
    g423_n_spl_11
  );


  or

  (
    g850_n,
    G7_p_spl_111,
    g423_p_spl_11
  );


  and

  (
    g851_p,
    G4_n_spl_1111,
    g850_n
  );


  or

  (
    g851_n,
    G4_p_spl_1111,
    g850_p
  );


  and

  (
    g852_p,
    G19_p_spl_1,
    g409_n_spl_111
  );


  or

  (
    g852_n,
    G19_n_spl_1,
    g409_p_spl_111
  );


  and

  (
    g853_p,
    G18_p_spl_1,
    g406_n_spl_111
  );


  or

  (
    g853_n,
    G18_n_spl_1,
    g406_p_spl_111
  );


  and

  (
    g854_p,
    g852_n,
    g853_n
  );


  or

  (
    g854_n,
    g852_p,
    g853_p
  );


  and

  (
    g855_p,
    g851_p,
    g854_p
  );


  or

  (
    g855_n,
    g851_n,
    g854_n
  );


  and

  (
    g856_p,
    g849_p,
    g855_p
  );


  or

  (
    g856_n,
    g849_n,
    g855_n
  );


  and

  (
    g857_p,
    g843_n,
    g856_n
  );


  or

  (
    g857_n,
    g843_p,
    g856_p
  );


  and

  (
    g858_p,
    g393_n_spl_111,
    g857_n
  );


  or

  (
    g858_n,
    g393_p_spl_111,
    g857_p
  );


  and

  (
    g859_p,
    g830_p,
    g858_n
  );


  or

  (
    g859_n,
    g830_n,
    g858_p
  );


  and

  (
    g860_p,
    g828_n,
    g859_p
  );


  or

  (
    g860_n,
    g828_p,
    g859_n
  );


  and

  (
    g861_p,
    g738_p_spl_1,
    g740_p_spl_
  );


  or

  (
    g861_n,
    g738_n_spl_1,
    g740_n_spl_
  );


  and

  (
    g862_p,
    g384_n_spl_1,
    g738_n_spl_1
  );


  or

  (
    g862_n,
    g384_p_spl_1,
    g738_p_spl_1
  );


  and

  (
    g863_p,
    g377_n_spl_11,
    g741_n_spl_
  );


  or

  (
    g863_n,
    g377_p_spl_1,
    g741_p_spl_
  );


  and

  (
    g864_p,
    g862_n,
    g863_n
  );


  or

  (
    g864_n,
    g862_p,
    g863_p
  );


  and

  (
    g865_p,
    g861_n,
    g864_n
  );


  or

  (
    g865_n,
    g861_p,
    g864_p
  );


  and

  (
    g866_p,
    g860_n,
    g865_n
  );


  or

  (
    g866_n,
    g860_p,
    g865_p
  );


  and

  (
    g867_p,
    g626_p_spl_,
    g722_p_spl_
  );


  or

  (
    g867_n,
    g626_n_spl_0,
    g722_n_spl_0
  );


  and

  (
    g868_p,
    g778_p_spl_,
    g827_p_spl_
  );


  or

  (
    g868_n,
    g778_n_spl_0,
    g827_n_spl_0
  );


  and

  (
    g869_p,
    g509_p_spl_,
    g866_p_spl_
  );


  or

  (
    g869_n,
    g509_n_spl_0,
    g866_n_spl_0
  );


  and

  (
    g870_p,
    g451_p_spl_,
    g679_p_spl_
  );


  or

  (
    g870_n,
    g451_n_spl_0,
    g679_n_spl_0
  );


  or

  (
    g871_n,
    g869_n_spl_,
    g870_n_spl_
  );


  or

  (
    g872_n,
    g868_n_spl_0,
    g871_n
  );


  or

  (
    g873_n,
    g867_n_spl_,
    g872_n
  );


  and

  (
    g874_p,
    G27_p_spl_0,
    G48_p_spl_
  );


  or

  (
    g874_n,
    G27_n_spl_,
    G48_n_spl_
  );


  or

  (
    g875_n,
    g868_n_spl_0,
    g874_n_spl_
  );


  and

  (
    g876_p,
    G27_p_spl_,
    g875_n
  );


  and

  (
    g877_p,
    g873_n_spl_,
    g876_p
  );


  and

  (
    g878_p,
    g451_n_spl_0,
    g679_n_spl_0
  );


  or

  (
    g878_n,
    g451_p_spl_,
    g679_p_spl_
  );


  and

  (
    g879_p,
    g870_n_spl_,
    g878_n
  );


  or

  (
    g879_n,
    g870_p,
    g878_p
  );


  and

  (
    g880_p,
    g626_n_spl_0,
    g722_n_spl_0
  );


  or

  (
    g880_n,
    g626_p_spl_,
    g722_p_spl_
  );


  and

  (
    g881_p,
    g867_n_spl_,
    g880_n
  );


  or

  (
    g881_n,
    g867_p,
    g880_p
  );


  and

  (
    g882_p,
    g879_p_spl_,
    g881_n_spl_
  );


  or

  (
    g882_n,
    g879_n_spl_,
    g881_p_spl_
  );


  and

  (
    g883_p,
    g879_n_spl_,
    g881_p_spl_
  );


  or

  (
    g883_n,
    g879_p_spl_,
    g881_n_spl_
  );


  and

  (
    g884_p,
    g882_n,
    g883_n
  );


  or

  (
    g884_n,
    g882_p,
    g883_p
  );


  and

  (
    g885_p,
    g509_n_spl_0,
    g866_n_spl_0
  );


  or

  (
    g885_n,
    g509_p_spl_,
    g866_p_spl_
  );


  and

  (
    g886_p,
    g869_n_spl_,
    g885_n
  );


  or

  (
    g886_n,
    g869_p,
    g885_p
  );


  and

  (
    g887_p,
    g778_n_spl_0,
    g827_n_spl_0
  );


  or

  (
    g887_n,
    g778_p_spl_,
    g827_p_spl_
  );


  and

  (
    g888_p,
    g868_n_spl_,
    g887_n
  );


  or

  (
    g888_n,
    g868_p,
    g887_p
  );


  and

  (
    g889_p,
    G50_n_spl_,
    g888_n_spl_0
  );


  or

  (
    g889_n,
    G50_p_spl_,
    g888_p_spl_0
  );


  and

  (
    g890_p,
    G50_p_spl_,
    g888_p_spl_0
  );


  or

  (
    g890_n,
    G50_n_spl_,
    g888_n_spl_0
  );


  and

  (
    g891_p,
    g874_n_spl_,
    g890_n
  );


  or

  (
    g891_n,
    g874_p,
    g890_p
  );


  and

  (
    g892_p,
    g889_n,
    g891_p
  );


  or

  (
    g892_n,
    g889_p,
    g891_n
  );


  and

  (
    g893_p,
    g886_p_spl_0,
    g892_n_spl_
  );


  or

  (
    g893_n,
    g886_n_spl_0,
    g892_p_spl_
  );


  and

  (
    g894_p,
    g886_n_spl_0,
    g892_p_spl_
  );


  or

  (
    g894_n,
    g886_p_spl_0,
    g892_n_spl_
  );


  and

  (
    g895_p,
    g893_n,
    g894_n
  );


  or

  (
    g895_n,
    g893_p,
    g894_p
  );


  and

  (
    g896_p,
    g884_n_spl_,
    g895_p
  );


  and

  (
    g897_p,
    g884_p_spl_,
    g895_n
  );


  or

  (
    g898_n,
    g896_p,
    g897_p
  );


  and

  (
    g899_p,
    g886_n_spl_1,
    g888_n_spl_1
  );


  or

  (
    g899_n,
    g886_p_spl_1,
    g888_p_spl_1
  );


  and

  (
    g900_p,
    g886_p_spl_1,
    g888_p_spl_1
  );


  or

  (
    g900_n,
    g886_n_spl_1,
    g888_n_spl_1
  );


  and

  (
    g901_p,
    g899_n,
    g900_n
  );


  or

  (
    g901_n,
    g899_p,
    g900_p
  );


  or

  (
    g902_n,
    g884_p_spl_,
    g901_p
  );


  or

  (
    g903_n,
    g884_n_spl_,
    g901_n
  );


  and

  (
    g904_p,
    g902_n,
    g903_n
  );


  buf

  (
    G3519,
    g53_p
  );


  buf

  (
    G3520,
    g55_n_spl_
  );


  buf

  (
    G3521,
    g84_p
  );


  buf

  (
    G3522,
    g105_p
  );


  buf

  (
    G3523,
    g125_n
  );


  buf

  (
    G3524,
    g350_p
  );


  buf

  (
    G3525,
    g364_n
  );


  buf

  (
    G3526,
    g376_p_spl_
  );


  buf

  (
    G3527,
    g381_n
  );


  buf

  (
    G3528,
    g451_n_spl_
  );


  buf

  (
    G3529,
    g509_n_spl_
  );


  buf

  (
    G3530,
    g551_n
  );


  buf

  (
    G3531,
    g626_n_spl_
  );


  buf

  (
    G3532,
    g679_n_spl_
  );


  buf

  (
    G3533,
    g722_n_spl_
  );


  buf

  (
    G3534,
    g778_n_spl_
  );


  buf

  (
    G3535,
    g827_n_spl_
  );


  buf

  (
    G3536,
    g866_n_spl_
  );


  buf

  (
    G3537,
    g873_n_spl_
  );


  not

  (
    G3538,
    g877_p
  );


  buf

  (
    G3539,
    g898_n
  );


  buf

  (
    G3540,
    g904_p
  );


  buf

  (
    G7_n_spl_,
    G7_n
  );


  buf

  (
    G7_n_spl_0,
    G7_n_spl_
  );


  buf

  (
    G7_n_spl_00,
    G7_n_spl_0
  );


  buf

  (
    G7_n_spl_000,
    G7_n_spl_00
  );


  buf

  (
    G7_n_spl_0000,
    G7_n_spl_000
  );


  buf

  (
    G7_n_spl_001,
    G7_n_spl_00
  );


  buf

  (
    G7_n_spl_01,
    G7_n_spl_0
  );


  buf

  (
    G7_n_spl_010,
    G7_n_spl_01
  );


  buf

  (
    G7_n_spl_011,
    G7_n_spl_01
  );


  buf

  (
    G7_n_spl_1,
    G7_n_spl_
  );


  buf

  (
    G7_n_spl_10,
    G7_n_spl_1
  );


  buf

  (
    G7_n_spl_100,
    G7_n_spl_10
  );


  buf

  (
    G7_n_spl_101,
    G7_n_spl_10
  );


  buf

  (
    G7_n_spl_11,
    G7_n_spl_1
  );


  buf

  (
    G7_n_spl_110,
    G7_n_spl_11
  );


  buf

  (
    G7_n_spl_111,
    G7_n_spl_11
  );


  buf

  (
    G8_n_spl_,
    G8_n
  );


  buf

  (
    G8_n_spl_0,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_00,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_000,
    G8_n_spl_00
  );


  buf

  (
    G8_n_spl_001,
    G8_n_spl_00
  );


  buf

  (
    G8_n_spl_01,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_010,
    G8_n_spl_01
  );


  buf

  (
    G8_n_spl_011,
    G8_n_spl_01
  );


  buf

  (
    G8_n_spl_1,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_10,
    G8_n_spl_1
  );


  buf

  (
    G8_n_spl_100,
    G8_n_spl_10
  );


  buf

  (
    G8_n_spl_101,
    G8_n_spl_10
  );


  buf

  (
    G8_n_spl_11,
    G8_n_spl_1
  );


  buf

  (
    G8_n_spl_110,
    G8_n_spl_11
  );


  buf

  (
    G7_p_spl_,
    G7_p
  );


  buf

  (
    G7_p_spl_0,
    G7_p_spl_
  );


  buf

  (
    G7_p_spl_00,
    G7_p_spl_0
  );


  buf

  (
    G7_p_spl_000,
    G7_p_spl_00
  );


  buf

  (
    G7_p_spl_0000,
    G7_p_spl_000
  );


  buf

  (
    G7_p_spl_0001,
    G7_p_spl_000
  );


  buf

  (
    G7_p_spl_001,
    G7_p_spl_00
  );


  buf

  (
    G7_p_spl_01,
    G7_p_spl_0
  );


  buf

  (
    G7_p_spl_010,
    G7_p_spl_01
  );


  buf

  (
    G7_p_spl_011,
    G7_p_spl_01
  );


  buf

  (
    G7_p_spl_1,
    G7_p_spl_
  );


  buf

  (
    G7_p_spl_10,
    G7_p_spl_1
  );


  buf

  (
    G7_p_spl_100,
    G7_p_spl_10
  );


  buf

  (
    G7_p_spl_101,
    G7_p_spl_10
  );


  buf

  (
    G7_p_spl_11,
    G7_p_spl_1
  );


  buf

  (
    G7_p_spl_110,
    G7_p_spl_11
  );


  buf

  (
    G7_p_spl_111,
    G7_p_spl_11
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_00,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_000,
    G8_p_spl_00
  );


  buf

  (
    G8_p_spl_001,
    G8_p_spl_00
  );


  buf

  (
    G8_p_spl_01,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_010,
    G8_p_spl_01
  );


  buf

  (
    G8_p_spl_011,
    G8_p_spl_01
  );


  buf

  (
    G8_p_spl_1,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_10,
    G8_p_spl_1
  );


  buf

  (
    G8_p_spl_100,
    G8_p_spl_10
  );


  buf

  (
    G8_p_spl_101,
    G8_p_spl_10
  );


  buf

  (
    G8_p_spl_11,
    G8_p_spl_1
  );


  buf

  (
    G8_p_spl_110,
    G8_p_spl_11
  );


  buf

  (
    G8_p_spl_111,
    G8_p_spl_11
  );


  buf

  (
    G9_n_spl_,
    G9_n
  );


  buf

  (
    G9_n_spl_0,
    G9_n_spl_
  );


  buf

  (
    G9_n_spl_00,
    G9_n_spl_0
  );


  buf

  (
    G9_n_spl_000,
    G9_n_spl_00
  );


  buf

  (
    G9_n_spl_001,
    G9_n_spl_00
  );


  buf

  (
    G9_n_spl_01,
    G9_n_spl_0
  );


  buf

  (
    G9_n_spl_010,
    G9_n_spl_01
  );


  buf

  (
    G9_n_spl_011,
    G9_n_spl_01
  );


  buf

  (
    G9_n_spl_1,
    G9_n_spl_
  );


  buf

  (
    G9_n_spl_10,
    G9_n_spl_1
  );


  buf

  (
    G9_n_spl_100,
    G9_n_spl_10
  );


  buf

  (
    G9_n_spl_101,
    G9_n_spl_10
  );


  buf

  (
    G9_n_spl_11,
    G9_n_spl_1
  );


  buf

  (
    G9_n_spl_110,
    G9_n_spl_11
  );


  buf

  (
    g51_p_spl_,
    g51_p
  );


  buf

  (
    G9_p_spl_,
    G9_p
  );


  buf

  (
    G9_p_spl_0,
    G9_p_spl_
  );


  buf

  (
    G9_p_spl_00,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_000,
    G9_p_spl_00
  );


  buf

  (
    G9_p_spl_001,
    G9_p_spl_00
  );


  buf

  (
    G9_p_spl_01,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_010,
    G9_p_spl_01
  );


  buf

  (
    G9_p_spl_011,
    G9_p_spl_01
  );


  buf

  (
    G9_p_spl_1,
    G9_p_spl_
  );


  buf

  (
    G9_p_spl_10,
    G9_p_spl_1
  );


  buf

  (
    G9_p_spl_100,
    G9_p_spl_10
  );


  buf

  (
    G9_p_spl_101,
    G9_p_spl_10
  );


  buf

  (
    G9_p_spl_11,
    G9_p_spl_1
  );


  buf

  (
    G9_p_spl_110,
    G9_p_spl_11
  );


  buf

  (
    g51_n_spl_,
    g51_n
  );


  buf

  (
    G10_n_spl_,
    G10_n
  );


  buf

  (
    G10_n_spl_0,
    G10_n_spl_
  );


  buf

  (
    G10_n_spl_00,
    G10_n_spl_0
  );


  buf

  (
    G10_n_spl_000,
    G10_n_spl_00
  );


  buf

  (
    G10_n_spl_001,
    G10_n_spl_00
  );


  buf

  (
    G10_n_spl_01,
    G10_n_spl_0
  );


  buf

  (
    G10_n_spl_010,
    G10_n_spl_01
  );


  buf

  (
    G10_n_spl_011,
    G10_n_spl_01
  );


  buf

  (
    G10_n_spl_1,
    G10_n_spl_
  );


  buf

  (
    G10_n_spl_10,
    G10_n_spl_1
  );


  buf

  (
    G10_n_spl_100,
    G10_n_spl_10
  );


  buf

  (
    G10_n_spl_101,
    G10_n_spl_10
  );


  buf

  (
    G10_n_spl_11,
    G10_n_spl_1
  );


  buf

  (
    G10_n_spl_110,
    G10_n_spl_11
  );


  buf

  (
    g52_p_spl_,
    g52_p
  );


  buf

  (
    G12_n_spl_,
    G12_n
  );


  buf

  (
    G12_n_spl_0,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_00,
    G12_n_spl_0
  );


  buf

  (
    G12_n_spl_000,
    G12_n_spl_00
  );


  buf

  (
    G12_n_spl_001,
    G12_n_spl_00
  );


  buf

  (
    G12_n_spl_01,
    G12_n_spl_0
  );


  buf

  (
    G12_n_spl_010,
    G12_n_spl_01
  );


  buf

  (
    G12_n_spl_011,
    G12_n_spl_01
  );


  buf

  (
    G12_n_spl_1,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_10,
    G12_n_spl_1
  );


  buf

  (
    G12_n_spl_100,
    G12_n_spl_10
  );


  buf

  (
    G12_n_spl_101,
    G12_n_spl_10
  );


  buf

  (
    G12_n_spl_11,
    G12_n_spl_1
  );


  buf

  (
    G13_n_spl_,
    G13_n
  );


  buf

  (
    G13_n_spl_0,
    G13_n_spl_
  );


  buf

  (
    G13_n_spl_00,
    G13_n_spl_0
  );


  buf

  (
    G13_n_spl_000,
    G13_n_spl_00
  );


  buf

  (
    G13_n_spl_001,
    G13_n_spl_00
  );


  buf

  (
    G13_n_spl_01,
    G13_n_spl_0
  );


  buf

  (
    G13_n_spl_010,
    G13_n_spl_01
  );


  buf

  (
    G13_n_spl_011,
    G13_n_spl_01
  );


  buf

  (
    G13_n_spl_1,
    G13_n_spl_
  );


  buf

  (
    G13_n_spl_10,
    G13_n_spl_1
  );


  buf

  (
    G13_n_spl_100,
    G13_n_spl_10
  );


  buf

  (
    G13_n_spl_101,
    G13_n_spl_10
  );


  buf

  (
    G13_n_spl_11,
    G13_n_spl_1
  );


  buf

  (
    G13_n_spl_110,
    G13_n_spl_11
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_00,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_000,
    G12_p_spl_00
  );


  buf

  (
    G12_p_spl_001,
    G12_p_spl_00
  );


  buf

  (
    G12_p_spl_01,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_010,
    G12_p_spl_01
  );


  buf

  (
    G12_p_spl_011,
    G12_p_spl_01
  );


  buf

  (
    G12_p_spl_1,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_10,
    G12_p_spl_1
  );


  buf

  (
    G12_p_spl_100,
    G12_p_spl_10
  );


  buf

  (
    G12_p_spl_101,
    G12_p_spl_10
  );


  buf

  (
    G12_p_spl_11,
    G12_p_spl_1
  );


  buf

  (
    G12_p_spl_110,
    G12_p_spl_11
  );


  buf

  (
    G13_p_spl_,
    G13_p
  );


  buf

  (
    G13_p_spl_0,
    G13_p_spl_
  );


  buf

  (
    G13_p_spl_00,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_000,
    G13_p_spl_00
  );


  buf

  (
    G13_p_spl_001,
    G13_p_spl_00
  );


  buf

  (
    G13_p_spl_01,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_010,
    G13_p_spl_01
  );


  buf

  (
    G13_p_spl_011,
    G13_p_spl_01
  );


  buf

  (
    G13_p_spl_1,
    G13_p_spl_
  );


  buf

  (
    G13_p_spl_10,
    G13_p_spl_1
  );


  buf

  (
    G13_p_spl_100,
    G13_p_spl_10
  );


  buf

  (
    G13_p_spl_101,
    G13_p_spl_10
  );


  buf

  (
    G13_p_spl_11,
    G13_p_spl_1
  );


  buf

  (
    G13_p_spl_110,
    G13_p_spl_11
  );


  buf

  (
    G13_p_spl_111,
    G13_p_spl_11
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    G11_p_spl_0,
    G11_p_spl_
  );


  buf

  (
    G11_p_spl_00,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_000,
    G11_p_spl_00
  );


  buf

  (
    G11_p_spl_001,
    G11_p_spl_00
  );


  buf

  (
    G11_p_spl_01,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_010,
    G11_p_spl_01
  );


  buf

  (
    G11_p_spl_011,
    G11_p_spl_01
  );


  buf

  (
    G11_p_spl_1,
    G11_p_spl_
  );


  buf

  (
    G11_p_spl_10,
    G11_p_spl_1
  );


  buf

  (
    G11_p_spl_100,
    G11_p_spl_10
  );


  buf

  (
    G11_p_spl_101,
    G11_p_spl_10
  );


  buf

  (
    G11_p_spl_11,
    G11_p_spl_1
  );


  buf

  (
    g54_n_spl_,
    g54_n
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    G11_n_spl_0,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_00,
    G11_n_spl_0
  );


  buf

  (
    G11_n_spl_000,
    G11_n_spl_00
  );


  buf

  (
    G11_n_spl_001,
    G11_n_spl_00
  );


  buf

  (
    G11_n_spl_01,
    G11_n_spl_0
  );


  buf

  (
    G11_n_spl_010,
    G11_n_spl_01
  );


  buf

  (
    G11_n_spl_011,
    G11_n_spl_01
  );


  buf

  (
    G11_n_spl_1,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_10,
    G11_n_spl_1
  );


  buf

  (
    G11_n_spl_100,
    G11_n_spl_10
  );


  buf

  (
    G11_n_spl_11,
    G11_n_spl_1
  );


  buf

  (
    g54_p_spl_,
    g54_p
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    G1_n_spl_00,
    G1_n_spl_0
  );


  buf

  (
    G1_n_spl_000,
    G1_n_spl_00
  );


  buf

  (
    G1_n_spl_001,
    G1_n_spl_00
  );


  buf

  (
    G1_n_spl_01,
    G1_n_spl_0
  );


  buf

  (
    G1_n_spl_010,
    G1_n_spl_01
  );


  buf

  (
    G1_n_spl_1,
    G1_n_spl_
  );


  buf

  (
    G1_n_spl_10,
    G1_n_spl_1
  );


  buf

  (
    G1_n_spl_11,
    G1_n_spl_1
  );


  buf

  (
    G3_n_spl_,
    G3_n
  );


  buf

  (
    G3_n_spl_0,
    G3_n_spl_
  );


  buf

  (
    G3_n_spl_00,
    G3_n_spl_0
  );


  buf

  (
    G3_n_spl_000,
    G3_n_spl_00
  );


  buf

  (
    G3_n_spl_0000,
    G3_n_spl_000
  );


  buf

  (
    G3_n_spl_0001,
    G3_n_spl_000
  );


  buf

  (
    G3_n_spl_001,
    G3_n_spl_00
  );


  buf

  (
    G3_n_spl_0010,
    G3_n_spl_001
  );


  buf

  (
    G3_n_spl_01,
    G3_n_spl_0
  );


  buf

  (
    G3_n_spl_010,
    G3_n_spl_01
  );


  buf

  (
    G3_n_spl_011,
    G3_n_spl_01
  );


  buf

  (
    G3_n_spl_1,
    G3_n_spl_
  );


  buf

  (
    G3_n_spl_10,
    G3_n_spl_1
  );


  buf

  (
    G3_n_spl_100,
    G3_n_spl_10
  );


  buf

  (
    G3_n_spl_101,
    G3_n_spl_10
  );


  buf

  (
    G3_n_spl_11,
    G3_n_spl_1
  );


  buf

  (
    G3_n_spl_110,
    G3_n_spl_11
  );


  buf

  (
    G3_n_spl_111,
    G3_n_spl_11
  );


  buf

  (
    G34_n_spl_,
    G34_n
  );


  buf

  (
    G34_n_spl_0,
    G34_n_spl_
  );


  buf

  (
    G34_n_spl_00,
    G34_n_spl_0
  );


  buf

  (
    G34_n_spl_01,
    G34_n_spl_0
  );


  buf

  (
    G34_n_spl_1,
    G34_n_spl_
  );


  buf

  (
    G34_n_spl_10,
    G34_n_spl_1
  );


  buf

  (
    G32_n_spl_,
    G32_n
  );


  buf

  (
    G32_n_spl_0,
    G32_n_spl_
  );


  buf

  (
    G32_n_spl_00,
    G32_n_spl_0
  );


  buf

  (
    G32_n_spl_01,
    G32_n_spl_0
  );


  buf

  (
    G32_n_spl_1,
    G32_n_spl_
  );


  buf

  (
    G36_n_spl_,
    G36_n
  );


  buf

  (
    G36_n_spl_0,
    G36_n_spl_
  );


  buf

  (
    G36_n_spl_00,
    G36_n_spl_0
  );


  buf

  (
    G36_n_spl_01,
    G36_n_spl_0
  );


  buf

  (
    G36_n_spl_1,
    G36_n_spl_
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


  buf

  (
    G10_p_spl_0,
    G10_p_spl_
  );


  buf

  (
    G10_p_spl_00,
    G10_p_spl_0
  );


  buf

  (
    G10_p_spl_000,
    G10_p_spl_00
  );


  buf

  (
    G10_p_spl_001,
    G10_p_spl_00
  );


  buf

  (
    G10_p_spl_01,
    G10_p_spl_0
  );


  buf

  (
    G10_p_spl_010,
    G10_p_spl_01
  );


  buf

  (
    G10_p_spl_011,
    G10_p_spl_01
  );


  buf

  (
    G10_p_spl_1,
    G10_p_spl_
  );


  buf

  (
    G10_p_spl_10,
    G10_p_spl_1
  );


  buf

  (
    G10_p_spl_100,
    G10_p_spl_10
  );


  buf

  (
    G10_p_spl_101,
    G10_p_spl_10
  );


  buf

  (
    G10_p_spl_11,
    G10_p_spl_1
  );


  buf

  (
    G33_n_spl_,
    G33_n
  );


  buf

  (
    G33_n_spl_0,
    G33_n_spl_
  );


  buf

  (
    G33_n_spl_00,
    G33_n_spl_0
  );


  buf

  (
    G33_n_spl_01,
    G33_n_spl_0
  );


  buf

  (
    G33_n_spl_1,
    G33_n_spl_
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G14_p_spl_0,
    G14_p_spl_
  );


  buf

  (
    G14_p_spl_00,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_000,
    G14_p_spl_00
  );


  buf

  (
    G14_p_spl_001,
    G14_p_spl_00
  );


  buf

  (
    G14_p_spl_01,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_010,
    G14_p_spl_01
  );


  buf

  (
    G14_p_spl_011,
    G14_p_spl_01
  );


  buf

  (
    G14_p_spl_1,
    G14_p_spl_
  );


  buf

  (
    G14_p_spl_10,
    G14_p_spl_1
  );


  buf

  (
    G14_p_spl_100,
    G14_p_spl_10
  );


  buf

  (
    G14_p_spl_101,
    G14_p_spl_10
  );


  buf

  (
    G14_p_spl_11,
    G14_p_spl_1
  );


  buf

  (
    G14_p_spl_110,
    G14_p_spl_11
  );


  buf

  (
    G14_p_spl_111,
    G14_p_spl_11
  );


  buf

  (
    G37_n_spl_,
    G37_n
  );


  buf

  (
    G37_n_spl_0,
    G37_n_spl_
  );


  buf

  (
    G37_n_spl_1,
    G37_n_spl_
  );


  buf

  (
    G31_n_spl_,
    G31_n
  );


  buf

  (
    G31_n_spl_0,
    G31_n_spl_
  );


  buf

  (
    G31_n_spl_00,
    G31_n_spl_0
  );


  buf

  (
    G31_n_spl_01,
    G31_n_spl_0
  );


  buf

  (
    G31_n_spl_1,
    G31_n_spl_
  );


  buf

  (
    G35_n_spl_,
    G35_n
  );


  buf

  (
    G35_n_spl_0,
    G35_n_spl_
  );


  buf

  (
    G35_n_spl_00,
    G35_n_spl_0
  );


  buf

  (
    G35_n_spl_01,
    G35_n_spl_0
  );


  buf

  (
    G35_n_spl_1,
    G35_n_spl_
  );


  buf

  (
    G35_n_spl_10,
    G35_n_spl_1
  );


  buf

  (
    G30_n_spl_,
    G30_n
  );


  buf

  (
    G30_n_spl_0,
    G30_n_spl_
  );


  buf

  (
    G30_n_spl_00,
    G30_n_spl_0
  );


  buf

  (
    G30_n_spl_01,
    G30_n_spl_0
  );


  buf

  (
    G30_n_spl_1,
    G30_n_spl_
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G2_p_spl_0,
    G2_p_spl_
  );


  buf

  (
    G2_p_spl_00,
    G2_p_spl_0
  );


  buf

  (
    G2_p_spl_1,
    G2_p_spl_
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G1_p_spl_0,
    G1_p_spl_
  );


  buf

  (
    G1_p_spl_00,
    G1_p_spl_0
  );


  buf

  (
    G1_p_spl_000,
    G1_p_spl_00
  );


  buf

  (
    G1_p_spl_01,
    G1_p_spl_0
  );


  buf

  (
    G1_p_spl_1,
    G1_p_spl_
  );


  buf

  (
    G1_p_spl_10,
    G1_p_spl_1
  );


  buf

  (
    G1_p_spl_11,
    G1_p_spl_1
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G2_n_spl_0,
    G2_n_spl_
  );


  buf

  (
    G2_n_spl_00,
    G2_n_spl_0
  );


  buf

  (
    G2_n_spl_1,
    G2_n_spl_
  );


  buf

  (
    g73_p_spl_,
    g73_p
  );


  buf

  (
    g73_p_spl_0,
    g73_p_spl_
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G3_p_spl_0,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_00,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_000,
    G3_p_spl_00
  );


  buf

  (
    G3_p_spl_0000,
    G3_p_spl_000
  );


  buf

  (
    G3_p_spl_0001,
    G3_p_spl_000
  );


  buf

  (
    G3_p_spl_001,
    G3_p_spl_00
  );


  buf

  (
    G3_p_spl_01,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_010,
    G3_p_spl_01
  );


  buf

  (
    G3_p_spl_011,
    G3_p_spl_01
  );


  buf

  (
    G3_p_spl_1,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_10,
    G3_p_spl_1
  );


  buf

  (
    G3_p_spl_100,
    G3_p_spl_10
  );


  buf

  (
    G3_p_spl_101,
    G3_p_spl_10
  );


  buf

  (
    G3_p_spl_11,
    G3_p_spl_1
  );


  buf

  (
    G3_p_spl_110,
    G3_p_spl_11
  );


  buf

  (
    G3_p_spl_111,
    G3_p_spl_11
  );


  buf

  (
    g73_n_spl_,
    g73_n
  );


  buf

  (
    g73_n_spl_0,
    g73_n_spl_
  );


  buf

  (
    g75_n_spl_,
    g75_n
  );


  buf

  (
    g75_p_spl_,
    g75_p
  );


  buf

  (
    g74_n_spl_,
    g74_n
  );


  buf

  (
    g76_n_spl_,
    g76_n
  );


  buf

  (
    g78_p_spl_,
    g78_p
  );


  buf

  (
    g78_n_spl_,
    g78_n
  );


  buf

  (
    g79_n_spl_,
    g79_n
  );


  buf

  (
    g79_n_spl_0,
    g79_n_spl_
  );


  buf

  (
    g79_n_spl_1,
    g79_n_spl_
  );


  buf

  (
    G36_p_spl_,
    G36_p
  );


  buf

  (
    G36_p_spl_0,
    G36_p_spl_
  );


  buf

  (
    G36_p_spl_1,
    G36_p_spl_
  );


  buf

  (
    G37_p_spl_,
    G37_p
  );


  buf

  (
    G37_p_spl_0,
    G37_p_spl_
  );


  buf

  (
    G34_p_spl_,
    G34_p
  );


  buf

  (
    G34_p_spl_0,
    G34_p_spl_
  );


  buf

  (
    G34_p_spl_00,
    G34_p_spl_0
  );


  buf

  (
    G34_p_spl_1,
    G34_p_spl_
  );


  buf

  (
    G35_p_spl_,
    G35_p
  );


  buf

  (
    G35_p_spl_0,
    G35_p_spl_
  );


  buf

  (
    G35_p_spl_00,
    G35_p_spl_0
  );


  buf

  (
    G35_p_spl_1,
    G35_p_spl_
  );


  buf

  (
    g87_p_spl_,
    g87_p
  );


  buf

  (
    g90_n_spl_,
    g90_n
  );


  buf

  (
    g87_n_spl_,
    g87_n
  );


  buf

  (
    g90_p_spl_,
    g90_p
  );


  buf

  (
    G32_p_spl_,
    G32_p
  );


  buf

  (
    G32_p_spl_0,
    G32_p_spl_
  );


  buf

  (
    G32_p_spl_00,
    G32_p_spl_0
  );


  buf

  (
    G32_p_spl_1,
    G32_p_spl_
  );


  buf

  (
    G33_p_spl_,
    G33_p
  );


  buf

  (
    G33_p_spl_0,
    G33_p_spl_
  );


  buf

  (
    G33_p_spl_00,
    G33_p_spl_0
  );


  buf

  (
    G33_p_spl_1,
    G33_p_spl_
  );


  buf

  (
    G30_p_spl_,
    G30_p
  );


  buf

  (
    G30_p_spl_0,
    G30_p_spl_
  );


  buf

  (
    G30_p_spl_00,
    G30_p_spl_0
  );


  buf

  (
    G30_p_spl_1,
    G30_p_spl_
  );


  buf

  (
    G31_p_spl_,
    G31_p
  );


  buf

  (
    G31_p_spl_0,
    G31_p_spl_
  );


  buf

  (
    G31_p_spl_00,
    G31_p_spl_0
  );


  buf

  (
    G31_p_spl_1,
    G31_p_spl_
  );


  buf

  (
    g96_n_spl_,
    g96_n
  );


  buf

  (
    g99_p_spl_,
    g99_p
  );


  buf

  (
    g96_p_spl_,
    g96_p
  );


  buf

  (
    g99_n_spl_,
    g99_n
  );


  buf

  (
    g102_p_spl_,
    g102_p
  );


  buf

  (
    g102_n_spl_,
    g102_n
  );


  buf

  (
    g106_n_spl_,
    g106_n
  );


  buf

  (
    g106_p_spl_,
    g106_p
  );


  buf

  (
    G14_n_spl_,
    G14_n
  );


  buf

  (
    G14_n_spl_0,
    G14_n_spl_
  );


  buf

  (
    G14_n_spl_00,
    G14_n_spl_0
  );


  buf

  (
    G14_n_spl_000,
    G14_n_spl_00
  );


  buf

  (
    G14_n_spl_001,
    G14_n_spl_00
  );


  buf

  (
    G14_n_spl_01,
    G14_n_spl_0
  );


  buf

  (
    G14_n_spl_010,
    G14_n_spl_01
  );


  buf

  (
    G14_n_spl_011,
    G14_n_spl_01
  );


  buf

  (
    G14_n_spl_1,
    G14_n_spl_
  );


  buf

  (
    G14_n_spl_10,
    G14_n_spl_1
  );


  buf

  (
    G14_n_spl_100,
    G14_n_spl_10
  );


  buf

  (
    G14_n_spl_101,
    G14_n_spl_10
  );


  buf

  (
    G14_n_spl_11,
    G14_n_spl_1
  );


  buf

  (
    G14_n_spl_110,
    G14_n_spl_11
  );


  buf

  (
    G14_n_spl_111,
    G14_n_spl_11
  );


  buf

  (
    g108_p_spl_,
    g108_p
  );


  buf

  (
    g111_n_spl_,
    g111_n
  );


  buf

  (
    g108_n_spl_,
    g108_n
  );


  buf

  (
    g111_p_spl_,
    g111_p
  );


  buf

  (
    g117_n_spl_,
    g117_n
  );


  buf

  (
    g117_p_spl_,
    g117_p
  );


  buf

  (
    g116_p_spl_,
    g116_p
  );


  buf

  (
    g119_n_spl_,
    g119_n
  );


  buf

  (
    g116_n_spl_,
    g116_n
  );


  buf

  (
    g119_p_spl_,
    g119_p
  );


  buf

  (
    g122_p_spl_,
    g122_p
  );


  buf

  (
    g122_n_spl_,
    g122_n
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_00,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_000,
    G4_p_spl_00
  );


  buf

  (
    G4_p_spl_0000,
    G4_p_spl_000
  );


  buf

  (
    G4_p_spl_00000,
    G4_p_spl_0000
  );


  buf

  (
    G4_p_spl_00001,
    G4_p_spl_0000
  );


  buf

  (
    G4_p_spl_0001,
    G4_p_spl_000
  );


  buf

  (
    G4_p_spl_00010,
    G4_p_spl_0001
  );


  buf

  (
    G4_p_spl_00011,
    G4_p_spl_0001
  );


  buf

  (
    G4_p_spl_001,
    G4_p_spl_00
  );


  buf

  (
    G4_p_spl_0010,
    G4_p_spl_001
  );


  buf

  (
    G4_p_spl_0011,
    G4_p_spl_001
  );


  buf

  (
    G4_p_spl_01,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_010,
    G4_p_spl_01
  );


  buf

  (
    G4_p_spl_0100,
    G4_p_spl_010
  );


  buf

  (
    G4_p_spl_0101,
    G4_p_spl_010
  );


  buf

  (
    G4_p_spl_011,
    G4_p_spl_01
  );


  buf

  (
    G4_p_spl_0110,
    G4_p_spl_011
  );


  buf

  (
    G4_p_spl_0111,
    G4_p_spl_011
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_10,
    G4_p_spl_1
  );


  buf

  (
    G4_p_spl_100,
    G4_p_spl_10
  );


  buf

  (
    G4_p_spl_1000,
    G4_p_spl_100
  );


  buf

  (
    G4_p_spl_1001,
    G4_p_spl_100
  );


  buf

  (
    G4_p_spl_101,
    G4_p_spl_10
  );


  buf

  (
    G4_p_spl_1010,
    G4_p_spl_101
  );


  buf

  (
    G4_p_spl_1011,
    G4_p_spl_101
  );


  buf

  (
    G4_p_spl_11,
    G4_p_spl_1
  );


  buf

  (
    G4_p_spl_110,
    G4_p_spl_11
  );


  buf

  (
    G4_p_spl_1100,
    G4_p_spl_110
  );


  buf

  (
    G4_p_spl_1101,
    G4_p_spl_110
  );


  buf

  (
    G4_p_spl_111,
    G4_p_spl_11
  );


  buf

  (
    G4_p_spl_1110,
    G4_p_spl_111
  );


  buf

  (
    G4_p_spl_1111,
    G4_p_spl_111
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    G4_n_spl_0,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_00,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_000,
    G4_n_spl_00
  );


  buf

  (
    G4_n_spl_0000,
    G4_n_spl_000
  );


  buf

  (
    G4_n_spl_00000,
    G4_n_spl_0000
  );


  buf

  (
    G4_n_spl_00001,
    G4_n_spl_0000
  );


  buf

  (
    G4_n_spl_0001,
    G4_n_spl_000
  );


  buf

  (
    G4_n_spl_00010,
    G4_n_spl_0001
  );


  buf

  (
    G4_n_spl_00011,
    G4_n_spl_0001
  );


  buf

  (
    G4_n_spl_001,
    G4_n_spl_00
  );


  buf

  (
    G4_n_spl_0010,
    G4_n_spl_001
  );


  buf

  (
    G4_n_spl_0011,
    G4_n_spl_001
  );


  buf

  (
    G4_n_spl_01,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_010,
    G4_n_spl_01
  );


  buf

  (
    G4_n_spl_0100,
    G4_n_spl_010
  );


  buf

  (
    G4_n_spl_0101,
    G4_n_spl_010
  );


  buf

  (
    G4_n_spl_011,
    G4_n_spl_01
  );


  buf

  (
    G4_n_spl_0110,
    G4_n_spl_011
  );


  buf

  (
    G4_n_spl_0111,
    G4_n_spl_011
  );


  buf

  (
    G4_n_spl_1,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_10,
    G4_n_spl_1
  );


  buf

  (
    G4_n_spl_100,
    G4_n_spl_10
  );


  buf

  (
    G4_n_spl_1000,
    G4_n_spl_100
  );


  buf

  (
    G4_n_spl_1001,
    G4_n_spl_100
  );


  buf

  (
    G4_n_spl_101,
    G4_n_spl_10
  );


  buf

  (
    G4_n_spl_1010,
    G4_n_spl_101
  );


  buf

  (
    G4_n_spl_1011,
    G4_n_spl_101
  );


  buf

  (
    G4_n_spl_11,
    G4_n_spl_1
  );


  buf

  (
    G4_n_spl_110,
    G4_n_spl_11
  );


  buf

  (
    G4_n_spl_1100,
    G4_n_spl_110
  );


  buf

  (
    G4_n_spl_1101,
    G4_n_spl_110
  );


  buf

  (
    G4_n_spl_111,
    G4_n_spl_11
  );


  buf

  (
    G4_n_spl_1110,
    G4_n_spl_111
  );


  buf

  (
    G4_n_spl_1111,
    G4_n_spl_111
  );


  buf

  (
    g126_n_spl_,
    g126_n
  );


  buf

  (
    g126_p_spl_,
    g126_p
  );


  buf

  (
    g129_p_spl_,
    g129_p
  );


  buf

  (
    g129_p_spl_0,
    g129_p_spl_
  );


  buf

  (
    g129_p_spl_00,
    g129_p_spl_0
  );


  buf

  (
    g129_p_spl_000,
    g129_p_spl_00
  );


  buf

  (
    g129_p_spl_001,
    g129_p_spl_00
  );


  buf

  (
    g129_p_spl_01,
    g129_p_spl_0
  );


  buf

  (
    g129_p_spl_1,
    g129_p_spl_
  );


  buf

  (
    g129_p_spl_10,
    g129_p_spl_1
  );


  buf

  (
    g129_p_spl_11,
    g129_p_spl_1
  );


  buf

  (
    g130_n_spl_,
    g130_n
  );


  buf

  (
    g130_n_spl_0,
    g130_n_spl_
  );


  buf

  (
    g130_n_spl_00,
    g130_n_spl_0
  );


  buf

  (
    g130_n_spl_01,
    g130_n_spl_0
  );


  buf

  (
    g130_n_spl_1,
    g130_n_spl_
  );


  buf

  (
    g130_n_spl_10,
    g130_n_spl_1
  );


  buf

  (
    g130_n_spl_11,
    g130_n_spl_1
  );


  buf

  (
    g129_n_spl_,
    g129_n
  );


  buf

  (
    g129_n_spl_0,
    g129_n_spl_
  );


  buf

  (
    g129_n_spl_00,
    g129_n_spl_0
  );


  buf

  (
    g129_n_spl_000,
    g129_n_spl_00
  );


  buf

  (
    g129_n_spl_001,
    g129_n_spl_00
  );


  buf

  (
    g129_n_spl_01,
    g129_n_spl_0
  );


  buf

  (
    g129_n_spl_1,
    g129_n_spl_
  );


  buf

  (
    g129_n_spl_10,
    g129_n_spl_1
  );


  buf

  (
    g129_n_spl_11,
    g129_n_spl_1
  );


  buf

  (
    g130_p_spl_,
    g130_p
  );


  buf

  (
    g130_p_spl_0,
    g130_p_spl_
  );


  buf

  (
    g130_p_spl_00,
    g130_p_spl_0
  );


  buf

  (
    g130_p_spl_01,
    g130_p_spl_0
  );


  buf

  (
    g130_p_spl_1,
    g130_p_spl_
  );


  buf

  (
    g130_p_spl_10,
    g130_p_spl_1
  );


  buf

  (
    g130_p_spl_11,
    g130_p_spl_1
  );


  buf

  (
    g131_p_spl_,
    g131_p
  );


  buf

  (
    g131_n_spl_,
    g131_n
  );


  buf

  (
    g133_n_spl_,
    g133_n
  );


  buf

  (
    g133_n_spl_0,
    g133_n_spl_
  );


  buf

  (
    g133_n_spl_1,
    g133_n_spl_
  );


  buf

  (
    g134_n_spl_,
    g134_n
  );


  buf

  (
    g134_n_spl_0,
    g134_n_spl_
  );


  buf

  (
    g133_p_spl_,
    g133_p
  );


  buf

  (
    g133_p_spl_0,
    g133_p_spl_
  );


  buf

  (
    g133_p_spl_1,
    g133_p_spl_
  );


  buf

  (
    g134_p_spl_,
    g134_p
  );


  buf

  (
    g134_p_spl_0,
    g134_p_spl_
  );


  buf

  (
    g137_n_spl_,
    g137_n
  );


  buf

  (
    g137_n_spl_0,
    g137_n_spl_
  );


  buf

  (
    g137_n_spl_00,
    g137_n_spl_0
  );


  buf

  (
    g137_n_spl_000,
    g137_n_spl_00
  );


  buf

  (
    g137_n_spl_01,
    g137_n_spl_0
  );


  buf

  (
    g137_n_spl_1,
    g137_n_spl_
  );


  buf

  (
    g137_n_spl_10,
    g137_n_spl_1
  );


  buf

  (
    g137_n_spl_11,
    g137_n_spl_1
  );


  buf

  (
    g137_p_spl_,
    g137_p
  );


  buf

  (
    g137_p_spl_0,
    g137_p_spl_
  );


  buf

  (
    g137_p_spl_00,
    g137_p_spl_0
  );


  buf

  (
    g137_p_spl_000,
    g137_p_spl_00
  );


  buf

  (
    g137_p_spl_01,
    g137_p_spl_0
  );


  buf

  (
    g137_p_spl_1,
    g137_p_spl_
  );


  buf

  (
    g137_p_spl_10,
    g137_p_spl_1
  );


  buf

  (
    g137_p_spl_11,
    g137_p_spl_1
  );


  buf

  (
    g138_p_spl_,
    g138_p
  );


  buf

  (
    g138_p_spl_0,
    g138_p_spl_
  );


  buf

  (
    g138_p_spl_00,
    g138_p_spl_0
  );


  buf

  (
    g138_p_spl_01,
    g138_p_spl_0
  );


  buf

  (
    g138_p_spl_1,
    g138_p_spl_
  );


  buf

  (
    g138_p_spl_10,
    g138_p_spl_1
  );


  buf

  (
    g138_p_spl_11,
    g138_p_spl_1
  );


  buf

  (
    g138_n_spl_,
    g138_n
  );


  buf

  (
    g138_n_spl_0,
    g138_n_spl_
  );


  buf

  (
    g138_n_spl_00,
    g138_n_spl_0
  );


  buf

  (
    g138_n_spl_01,
    g138_n_spl_0
  );


  buf

  (
    g138_n_spl_1,
    g138_n_spl_
  );


  buf

  (
    g138_n_spl_10,
    g138_n_spl_1
  );


  buf

  (
    g138_n_spl_11,
    g138_n_spl_1
  );


  buf

  (
    G39_p_spl_,
    G39_p
  );


  buf

  (
    G39_p_spl_0,
    G39_p_spl_
  );


  buf

  (
    G39_p_spl_00,
    G39_p_spl_0
  );


  buf

  (
    G39_p_spl_000,
    G39_p_spl_00
  );


  buf

  (
    G39_p_spl_01,
    G39_p_spl_0
  );


  buf

  (
    G39_p_spl_1,
    G39_p_spl_
  );


  buf

  (
    G39_p_spl_10,
    G39_p_spl_1
  );


  buf

  (
    G39_p_spl_11,
    G39_p_spl_1
  );


  buf

  (
    G39_n_spl_,
    G39_n
  );


  buf

  (
    G39_n_spl_0,
    G39_n_spl_
  );


  buf

  (
    G39_n_spl_00,
    G39_n_spl_0
  );


  buf

  (
    G39_n_spl_000,
    G39_n_spl_00
  );


  buf

  (
    G39_n_spl_01,
    G39_n_spl_0
  );


  buf

  (
    G39_n_spl_1,
    G39_n_spl_
  );


  buf

  (
    G39_n_spl_10,
    G39_n_spl_1
  );


  buf

  (
    G39_n_spl_11,
    G39_n_spl_1
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G5_p_spl_0,
    G5_p_spl_
  );


  buf

  (
    G5_p_spl_00,
    G5_p_spl_0
  );


  buf

  (
    G5_p_spl_01,
    G5_p_spl_0
  );


  buf

  (
    G5_p_spl_1,
    G5_p_spl_
  );


  buf

  (
    G5_n_spl_,
    G5_n
  );


  buf

  (
    G5_n_spl_0,
    G5_n_spl_
  );


  buf

  (
    G5_n_spl_00,
    G5_n_spl_0
  );


  buf

  (
    G5_n_spl_01,
    G5_n_spl_0
  );


  buf

  (
    G5_n_spl_1,
    G5_n_spl_
  );


  buf

  (
    g146_n_spl_,
    g146_n
  );


  buf

  (
    g146_p_spl_,
    g146_p
  );


  buf

  (
    g147_n_spl_,
    g147_n
  );


  buf

  (
    g147_n_spl_0,
    g147_n_spl_
  );


  buf

  (
    g147_n_spl_00,
    g147_n_spl_0
  );


  buf

  (
    g147_n_spl_000,
    g147_n_spl_00
  );


  buf

  (
    g147_n_spl_01,
    g147_n_spl_0
  );


  buf

  (
    g147_n_spl_1,
    g147_n_spl_
  );


  buf

  (
    g147_n_spl_10,
    g147_n_spl_1
  );


  buf

  (
    g147_n_spl_11,
    g147_n_spl_1
  );


  buf

  (
    g147_p_spl_,
    g147_p
  );


  buf

  (
    g147_p_spl_0,
    g147_p_spl_
  );


  buf

  (
    g147_p_spl_00,
    g147_p_spl_0
  );


  buf

  (
    g147_p_spl_000,
    g147_p_spl_00
  );


  buf

  (
    g147_p_spl_01,
    g147_p_spl_0
  );


  buf

  (
    g147_p_spl_1,
    g147_p_spl_
  );


  buf

  (
    g147_p_spl_10,
    g147_p_spl_1
  );


  buf

  (
    g147_p_spl_11,
    g147_p_spl_1
  );


  buf

  (
    G6_n_spl_,
    G6_n
  );


  buf

  (
    G6_n_spl_0,
    G6_n_spl_
  );


  buf

  (
    G6_n_spl_00,
    G6_n_spl_0
  );


  buf

  (
    G6_n_spl_01,
    G6_n_spl_0
  );


  buf

  (
    G6_n_spl_1,
    G6_n_spl_
  );


  buf

  (
    G6_n_spl_10,
    G6_n_spl_1
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G6_p_spl_0,
    G6_p_spl_
  );


  buf

  (
    G6_p_spl_00,
    G6_p_spl_0
  );


  buf

  (
    G6_p_spl_01,
    G6_p_spl_0
  );


  buf

  (
    G6_p_spl_1,
    G6_p_spl_
  );


  buf

  (
    G6_p_spl_10,
    G6_p_spl_1
  );


  buf

  (
    g149_p_spl_,
    g149_p
  );


  buf

  (
    g149_p_spl_0,
    g149_p_spl_
  );


  buf

  (
    g149_n_spl_,
    g149_n
  );


  buf

  (
    g149_n_spl_0,
    g149_n_spl_
  );


  buf

  (
    g148_p_spl_,
    g148_p
  );


  buf

  (
    g148_p_spl_0,
    g148_p_spl_
  );


  buf

  (
    g150_p_spl_,
    g150_p
  );


  buf

  (
    g150_p_spl_0,
    g150_p_spl_
  );


  buf

  (
    g150_p_spl_1,
    g150_p_spl_
  );


  buf

  (
    g148_n_spl_,
    g148_n
  );


  buf

  (
    g148_n_spl_0,
    g148_n_spl_
  );


  buf

  (
    g150_n_spl_,
    g150_n
  );


  buf

  (
    g150_n_spl_0,
    g150_n_spl_
  );


  buf

  (
    g150_n_spl_1,
    g150_n_spl_
  );


  buf

  (
    g153_p_spl_,
    g153_p
  );


  buf

  (
    g153_p_spl_0,
    g153_p_spl_
  );


  buf

  (
    g153_p_spl_00,
    g153_p_spl_0
  );


  buf

  (
    g153_p_spl_01,
    g153_p_spl_0
  );


  buf

  (
    g153_p_spl_1,
    g153_p_spl_
  );


  buf

  (
    g153_p_spl_10,
    g153_p_spl_1
  );


  buf

  (
    g153_p_spl_11,
    g153_p_spl_1
  );


  buf

  (
    g153_n_spl_,
    g153_n
  );


  buf

  (
    g153_n_spl_0,
    g153_n_spl_
  );


  buf

  (
    g153_n_spl_00,
    g153_n_spl_0
  );


  buf

  (
    g153_n_spl_01,
    g153_n_spl_0
  );


  buf

  (
    g153_n_spl_1,
    g153_n_spl_
  );


  buf

  (
    g153_n_spl_10,
    g153_n_spl_1
  );


  buf

  (
    g153_n_spl_11,
    g153_n_spl_1
  );


  buf

  (
    G41_n_spl_,
    G41_n
  );


  buf

  (
    G41_n_spl_0,
    G41_n_spl_
  );


  buf

  (
    G41_n_spl_00,
    G41_n_spl_0
  );


  buf

  (
    G41_n_spl_01,
    G41_n_spl_0
  );


  buf

  (
    G41_n_spl_1,
    G41_n_spl_
  );


  buf

  (
    G41_n_spl_10,
    G41_n_spl_1
  );


  buf

  (
    G41_p_spl_,
    G41_p
  );


  buf

  (
    G41_p_spl_0,
    G41_p_spl_
  );


  buf

  (
    G41_p_spl_00,
    G41_p_spl_0
  );


  buf

  (
    G41_p_spl_01,
    G41_p_spl_0
  );


  buf

  (
    G41_p_spl_1,
    G41_p_spl_
  );


  buf

  (
    G41_p_spl_10,
    G41_p_spl_1
  );


  buf

  (
    g151_n_spl_,
    g151_n
  );


  buf

  (
    g151_n_spl_0,
    g151_n_spl_
  );


  buf

  (
    g151_p_spl_,
    g151_p
  );


  buf

  (
    g151_p_spl_0,
    g151_p_spl_
  );


  buf

  (
    G25_n_spl_,
    G25_n
  );


  buf

  (
    G26_n_spl_,
    G26_n
  );


  buf

  (
    G26_n_spl_0,
    G26_n_spl_
  );


  buf

  (
    G25_p_spl_,
    G25_p
  );


  buf

  (
    G26_p_spl_,
    G26_p
  );


  buf

  (
    G26_p_spl_0,
    G26_p_spl_
  );


  buf

  (
    g161_p_spl_,
    g161_p
  );


  buf

  (
    g161_p_spl_0,
    g161_p_spl_
  );


  buf

  (
    g161_p_spl_1,
    g161_p_spl_
  );


  buf

  (
    g162_n_spl_,
    g162_n
  );


  buf

  (
    g162_n_spl_0,
    g162_n_spl_
  );


  buf

  (
    g162_n_spl_00,
    g162_n_spl_0
  );


  buf

  (
    g162_n_spl_000,
    g162_n_spl_00
  );


  buf

  (
    g162_n_spl_01,
    g162_n_spl_0
  );


  buf

  (
    g162_n_spl_1,
    g162_n_spl_
  );


  buf

  (
    g162_n_spl_10,
    g162_n_spl_1
  );


  buf

  (
    g162_n_spl_11,
    g162_n_spl_1
  );


  buf

  (
    g161_n_spl_,
    g161_n
  );


  buf

  (
    g161_n_spl_0,
    g161_n_spl_
  );


  buf

  (
    g161_n_spl_1,
    g161_n_spl_
  );


  buf

  (
    g162_p_spl_,
    g162_p
  );


  buf

  (
    g162_p_spl_0,
    g162_p_spl_
  );


  buf

  (
    g162_p_spl_00,
    g162_p_spl_0
  );


  buf

  (
    g162_p_spl_000,
    g162_p_spl_00
  );


  buf

  (
    g162_p_spl_01,
    g162_p_spl_0
  );


  buf

  (
    g162_p_spl_1,
    g162_p_spl_
  );


  buf

  (
    g162_p_spl_10,
    g162_p_spl_1
  );


  buf

  (
    g162_p_spl_11,
    g162_p_spl_1
  );


  buf

  (
    g145_p_spl_,
    g145_p
  );


  buf

  (
    g145_p_spl_0,
    g145_p_spl_
  );


  buf

  (
    g145_n_spl_,
    g145_n
  );


  buf

  (
    g145_n_spl_0,
    g145_n_spl_
  );


  buf

  (
    G23_n_spl_,
    G23_n
  );


  buf

  (
    G24_n_spl_,
    G24_n
  );


  buf

  (
    G24_n_spl_0,
    G24_n_spl_
  );


  buf

  (
    G24_n_spl_1,
    G24_n_spl_
  );


  buf

  (
    G23_p_spl_,
    G23_p
  );


  buf

  (
    G24_p_spl_,
    G24_p
  );


  buf

  (
    G24_p_spl_0,
    G24_p_spl_
  );


  buf

  (
    G24_p_spl_1,
    G24_p_spl_
  );


  buf

  (
    g165_n_spl_,
    g165_n
  );


  buf

  (
    g165_n_spl_0,
    g165_n_spl_
  );


  buf

  (
    g165_n_spl_00,
    g165_n_spl_0
  );


  buf

  (
    g165_n_spl_01,
    g165_n_spl_0
  );


  buf

  (
    g165_n_spl_1,
    g165_n_spl_
  );


  buf

  (
    g165_n_spl_10,
    g165_n_spl_1
  );


  buf

  (
    g165_n_spl_11,
    g165_n_spl_1
  );


  buf

  (
    g165_p_spl_,
    g165_p
  );


  buf

  (
    g165_p_spl_0,
    g165_p_spl_
  );


  buf

  (
    g165_p_spl_00,
    g165_p_spl_0
  );


  buf

  (
    g165_p_spl_01,
    g165_p_spl_0
  );


  buf

  (
    g165_p_spl_1,
    g165_p_spl_
  );


  buf

  (
    g165_p_spl_10,
    g165_p_spl_1
  );


  buf

  (
    g165_p_spl_11,
    g165_p_spl_1
  );


  buf

  (
    g167_n_spl_,
    g167_n
  );


  buf

  (
    g167_n_spl_0,
    g167_n_spl_
  );


  buf

  (
    g167_p_spl_,
    g167_p
  );


  buf

  (
    g167_p_spl_0,
    g167_p_spl_
  );


  buf

  (
    g169_n_spl_,
    g169_n
  );


  buf

  (
    g169_p_spl_,
    g169_p
  );


  buf

  (
    G40_n_spl_,
    G40_n
  );


  buf

  (
    G40_n_spl_0,
    G40_n_spl_
  );


  buf

  (
    G40_n_spl_00,
    G40_n_spl_0
  );


  buf

  (
    G40_n_spl_01,
    G40_n_spl_0
  );


  buf

  (
    G40_n_spl_1,
    G40_n_spl_
  );


  buf

  (
    G40_n_spl_10,
    G40_n_spl_1
  );


  buf

  (
    G40_p_spl_,
    G40_p
  );


  buf

  (
    G40_p_spl_0,
    G40_p_spl_
  );


  buf

  (
    G40_p_spl_00,
    G40_p_spl_0
  );


  buf

  (
    G40_p_spl_01,
    G40_p_spl_0
  );


  buf

  (
    G40_p_spl_1,
    G40_p_spl_
  );


  buf

  (
    G40_p_spl_10,
    G40_p_spl_1
  );


  buf

  (
    g186_p_spl_,
    g186_p
  );


  buf

  (
    g186_p_spl_0,
    g186_p_spl_
  );


  buf

  (
    g186_p_spl_1,
    g186_p_spl_
  );


  buf

  (
    g186_n_spl_,
    g186_n
  );


  buf

  (
    g186_n_spl_0,
    g186_n_spl_
  );


  buf

  (
    g186_n_spl_1,
    g186_n_spl_
  );


  buf

  (
    g177_p_spl_,
    g177_p
  );


  buf

  (
    g177_p_spl_0,
    g177_p_spl_
  );


  buf

  (
    g177_n_spl_,
    g177_n
  );


  buf

  (
    g177_n_spl_0,
    g177_n_spl_
  );


  buf

  (
    g190_n_spl_,
    g190_n
  );


  buf

  (
    g190_n_spl_0,
    g190_n_spl_
  );


  buf

  (
    g190_p_spl_,
    g190_p
  );


  buf

  (
    g190_p_spl_0,
    g190_p_spl_
  );


  buf

  (
    g196_n_spl_,
    g196_n
  );


  buf

  (
    g196_p_spl_,
    g196_p
  );


  buf

  (
    g212_p_spl_,
    g212_p
  );


  buf

  (
    g212_p_spl_0,
    g212_p_spl_
  );


  buf

  (
    g212_p_spl_1,
    g212_p_spl_
  );


  buf

  (
    g212_n_spl_,
    g212_n
  );


  buf

  (
    g212_n_spl_0,
    g212_n_spl_
  );


  buf

  (
    g212_n_spl_1,
    g212_n_spl_
  );


  buf

  (
    g202_p_spl_,
    g202_p
  );


  buf

  (
    g202_p_spl_0,
    g202_p_spl_
  );


  buf

  (
    g202_n_spl_,
    g202_n
  );


  buf

  (
    g202_n_spl_0,
    g202_n_spl_
  );


  buf

  (
    g216_n_spl_,
    g216_n
  );


  buf

  (
    g216_p_spl_,
    g216_p
  );


  buf

  (
    g223_n_spl_,
    g223_n
  );


  buf

  (
    g238_p_spl_,
    g238_p
  );


  buf

  (
    g238_p_spl_0,
    g238_p_spl_
  );


  buf

  (
    g238_p_spl_1,
    g238_p_spl_
  );


  buf

  (
    g238_n_spl_,
    g238_n
  );


  buf

  (
    g238_n_spl_0,
    g238_n_spl_
  );


  buf

  (
    g238_n_spl_1,
    g238_n_spl_
  );


  buf

  (
    g229_p_spl_,
    g229_p
  );


  buf

  (
    g229_p_spl_0,
    g229_p_spl_
  );


  buf

  (
    g229_n_spl_,
    g229_n
  );


  buf

  (
    g229_n_spl_0,
    g229_n_spl_
  );


  buf

  (
    g242_n_spl_,
    g242_n
  );


  buf

  (
    g242_n_spl_0,
    g242_n_spl_
  );


  buf

  (
    g242_p_spl_,
    g242_p
  );


  buf

  (
    g242_p_spl_0,
    g242_p_spl_
  );


  buf

  (
    g217_p_spl_,
    g217_p
  );


  buf

  (
    g217_p_spl_0,
    g217_p_spl_
  );


  buf

  (
    g217_p_spl_1,
    g217_p_spl_
  );


  buf

  (
    g243_p_spl_,
    g243_p
  );


  buf

  (
    g243_p_spl_0,
    g243_p_spl_
  );


  buf

  (
    g217_n_spl_,
    g217_n
  );


  buf

  (
    g217_n_spl_0,
    g217_n_spl_
  );


  buf

  (
    g217_n_spl_1,
    g217_n_spl_
  );


  buf

  (
    g243_n_spl_,
    g243_n
  );


  buf

  (
    g243_n_spl_0,
    g243_n_spl_
  );


  buf

  (
    g191_p_spl_,
    g191_p
  );


  buf

  (
    g191_p_spl_0,
    g191_p_spl_
  );


  buf

  (
    g244_p_spl_,
    g244_p
  );


  buf

  (
    g191_n_spl_,
    g191_n
  );


  buf

  (
    g191_n_spl_0,
    g191_n_spl_
  );


  buf

  (
    g244_n_spl_,
    g244_n
  );


  buf

  (
    g168_p_spl_,
    g168_p
  );


  buf

  (
    g168_p_spl_0,
    g168_p_spl_
  );


  buf

  (
    g245_p_spl_,
    g245_p
  );


  buf

  (
    g168_n_spl_,
    g168_n
  );


  buf

  (
    g168_n_spl_0,
    g168_n_spl_
  );


  buf

  (
    g245_n_spl_,
    g245_n
  );


  buf

  (
    g248_n_spl_,
    g248_n
  );


  buf

  (
    g248_n_spl_0,
    g248_n_spl_
  );


  buf

  (
    g248_n_spl_1,
    g248_n_spl_
  );


  buf

  (
    g248_p_spl_,
    g248_p
  );


  buf

  (
    g248_p_spl_0,
    g248_p_spl_
  );


  buf

  (
    g248_p_spl_1,
    g248_p_spl_
  );


  buf

  (
    g259_p_spl_,
    g259_p
  );


  buf

  (
    g259_p_spl_0,
    g259_p_spl_
  );


  buf

  (
    g259_p_spl_00,
    g259_p_spl_0
  );


  buf

  (
    g259_p_spl_1,
    g259_p_spl_
  );


  buf

  (
    g259_n_spl_,
    g259_n
  );


  buf

  (
    g259_n_spl_0,
    g259_n_spl_
  );


  buf

  (
    g259_n_spl_00,
    g259_n_spl_0
  );


  buf

  (
    g259_n_spl_1,
    g259_n_spl_
  );


  buf

  (
    g260_n_spl_,
    g260_n
  );


  buf

  (
    g260_n_spl_0,
    g260_n_spl_
  );


  buf

  (
    g260_n_spl_1,
    g260_n_spl_
  );


  buf

  (
    g260_p_spl_,
    g260_p
  );


  buf

  (
    g260_p_spl_0,
    g260_p_spl_
  );


  buf

  (
    g260_p_spl_1,
    g260_p_spl_
  );


  buf

  (
    g269_p_spl_,
    g269_p
  );


  buf

  (
    g269_n_spl_,
    g269_n
  );


  buf

  (
    g257_p_spl_,
    g257_p
  );


  buf

  (
    g257_p_spl_0,
    g257_p_spl_
  );


  buf

  (
    g257_n_spl_,
    g257_n
  );


  buf

  (
    g257_n_spl_0,
    g257_n_spl_
  );


  buf

  (
    g273_n_spl_,
    g273_n
  );


  buf

  (
    g273_n_spl_0,
    g273_n_spl_
  );


  buf

  (
    g273_p_spl_,
    g273_p
  );


  buf

  (
    g273_p_spl_0,
    g273_p_spl_
  );


  buf

  (
    g291_p_spl_,
    g291_p
  );


  buf

  (
    g291_n_spl_,
    g291_n
  );


  buf

  (
    g282_p_spl_,
    g282_p
  );


  buf

  (
    g282_p_spl_0,
    g282_p_spl_
  );


  buf

  (
    g282_n_spl_,
    g282_n
  );


  buf

  (
    g282_n_spl_0,
    g282_n_spl_
  );


  buf

  (
    g295_n_spl_,
    g295_n
  );


  buf

  (
    g295_n_spl_0,
    g295_n_spl_
  );


  buf

  (
    g295_p_spl_,
    g295_p
  );


  buf

  (
    g295_p_spl_0,
    g295_p_spl_
  );


  buf

  (
    G21_p_spl_,
    G21_p
  );


  buf

  (
    G21_p_spl_0,
    G21_p_spl_
  );


  buf

  (
    G21_p_spl_00,
    G21_p_spl_0
  );


  buf

  (
    G21_p_spl_01,
    G21_p_spl_0
  );


  buf

  (
    G21_p_spl_1,
    G21_p_spl_
  );


  buf

  (
    G21_p_spl_10,
    G21_p_spl_1
  );


  buf

  (
    G21_p_spl_11,
    G21_p_spl_1
  );


  buf

  (
    G21_n_spl_,
    G21_n
  );


  buf

  (
    G21_n_spl_0,
    G21_n_spl_
  );


  buf

  (
    G21_n_spl_00,
    G21_n_spl_0
  );


  buf

  (
    G21_n_spl_01,
    G21_n_spl_0
  );


  buf

  (
    G21_n_spl_1,
    G21_n_spl_
  );


  buf

  (
    G21_n_spl_10,
    G21_n_spl_1
  );


  buf

  (
    G21_n_spl_11,
    G21_n_spl_1
  );


  buf

  (
    G29_n_spl_,
    G29_n
  );


  buf

  (
    G29_p_spl_,
    G29_p
  );


  buf

  (
    g315_p_spl_,
    g315_p
  );


  buf

  (
    g315_n_spl_,
    g315_n
  );


  buf

  (
    g306_p_spl_,
    g306_p
  );


  buf

  (
    g306_p_spl_0,
    g306_p_spl_
  );


  buf

  (
    g306_n_spl_,
    g306_n
  );


  buf

  (
    g306_n_spl_0,
    g306_n_spl_
  );


  buf

  (
    g319_n_spl_,
    g319_n
  );


  buf

  (
    g319_p_spl_,
    g319_p
  );


  buf

  (
    g326_n_spl_,
    g326_n
  );


  buf

  (
    G22_p_spl_,
    G22_p
  );


  buf

  (
    G22_p_spl_0,
    G22_p_spl_
  );


  buf

  (
    G22_p_spl_00,
    G22_p_spl_0
  );


  buf

  (
    G22_p_spl_01,
    G22_p_spl_0
  );


  buf

  (
    G22_p_spl_1,
    G22_p_spl_
  );


  buf

  (
    G22_p_spl_10,
    G22_p_spl_1
  );


  buf

  (
    G22_p_spl_11,
    G22_p_spl_1
  );


  buf

  (
    G22_n_spl_,
    G22_n
  );


  buf

  (
    G22_n_spl_0,
    G22_n_spl_
  );


  buf

  (
    G22_n_spl_00,
    G22_n_spl_0
  );


  buf

  (
    G22_n_spl_01,
    G22_n_spl_0
  );


  buf

  (
    G22_n_spl_1,
    G22_n_spl_
  );


  buf

  (
    G22_n_spl_10,
    G22_n_spl_1
  );


  buf

  (
    G22_n_spl_11,
    G22_n_spl_1
  );


  buf

  (
    g341_p_spl_,
    g341_p
  );


  buf

  (
    g341_n_spl_,
    g341_n
  );


  buf

  (
    g332_p_spl_,
    g332_p
  );


  buf

  (
    g332_p_spl_0,
    g332_p_spl_
  );


  buf

  (
    g332_n_spl_,
    g332_n
  );


  buf

  (
    g332_n_spl_0,
    g332_n_spl_
  );


  buf

  (
    g345_n_spl_,
    g345_n
  );


  buf

  (
    g345_n_spl_0,
    g345_n_spl_
  );


  buf

  (
    g345_p_spl_,
    g345_p
  );


  buf

  (
    g345_p_spl_0,
    g345_p_spl_
  );


  buf

  (
    g320_p_spl_,
    g320_p
  );


  buf

  (
    g320_p_spl_0,
    g320_p_spl_
  );


  buf

  (
    g320_p_spl_1,
    g320_p_spl_
  );


  buf

  (
    g346_p_spl_,
    g346_p
  );


  buf

  (
    g346_p_spl_0,
    g346_p_spl_
  );


  buf

  (
    g320_n_spl_,
    g320_n
  );


  buf

  (
    g320_n_spl_0,
    g320_n_spl_
  );


  buf

  (
    g320_n_spl_1,
    g320_n_spl_
  );


  buf

  (
    g346_n_spl_,
    g346_n
  );


  buf

  (
    g346_n_spl_0,
    g346_n_spl_
  );


  buf

  (
    g296_p_spl_,
    g296_p
  );


  buf

  (
    g296_p_spl_0,
    g296_p_spl_
  );


  buf

  (
    g347_p_spl_,
    g347_p
  );


  buf

  (
    g296_n_spl_,
    g296_n
  );


  buf

  (
    g296_n_spl_0,
    g296_n_spl_
  );


  buf

  (
    g347_n_spl_,
    g347_n
  );


  buf

  (
    g274_p_spl_,
    g274_p
  );


  buf

  (
    g274_p_spl_0,
    g274_p_spl_
  );


  buf

  (
    g348_p_spl_,
    g348_p
  );


  buf

  (
    g274_n_spl_,
    g274_n
  );


  buf

  (
    g274_n_spl_0,
    g274_n_spl_
  );


  buf

  (
    g348_n_spl_,
    g348_n
  );


  buf

  (
    g246_p_spl_,
    g246_p
  );


  buf

  (
    g349_p_spl_,
    g349_p
  );


  buf

  (
    g349_p_spl_0,
    g349_p_spl_
  );


  buf

  (
    g349_p_spl_1,
    g349_p_spl_
  );


  buf

  (
    g356_n_spl_,
    g356_n
  );


  buf

  (
    g363_n_spl_,
    g363_n
  );


  buf

  (
    G27_p_spl_,
    G27_p
  );


  buf

  (
    G27_p_spl_0,
    G27_p_spl_
  );


  buf

  (
    g79_p_spl_,
    g79_p
  );


  buf

  (
    g79_p_spl_0,
    g79_p_spl_
  );


  buf

  (
    G27_n_spl_,
    G27_n
  );


  buf

  (
    G48_p_spl_,
    G48_p
  );


  buf

  (
    g365_p_spl_,
    g365_p
  );


  buf

  (
    g365_p_spl_0,
    g365_p_spl_
  );


  buf

  (
    g365_p_spl_1,
    g365_p_spl_
  );


  buf

  (
    G48_n_spl_,
    G48_n
  );


  buf

  (
    g365_n_spl_,
    g365_n
  );


  buf

  (
    g365_n_spl_0,
    g365_n_spl_
  );


  buf

  (
    g365_n_spl_1,
    g365_n_spl_
  );


  buf

  (
    g366_p_spl_,
    g366_p
  );


  buf

  (
    g366_p_spl_0,
    g366_p_spl_
  );


  buf

  (
    g366_p_spl_00,
    g366_p_spl_0
  );


  buf

  (
    g366_p_spl_000,
    g366_p_spl_00
  );


  buf

  (
    g366_p_spl_001,
    g366_p_spl_00
  );


  buf

  (
    g366_p_spl_01,
    g366_p_spl_0
  );


  buf

  (
    g366_p_spl_010,
    g366_p_spl_01
  );


  buf

  (
    g366_p_spl_011,
    g366_p_spl_01
  );


  buf

  (
    g366_p_spl_1,
    g366_p_spl_
  );


  buf

  (
    g366_p_spl_10,
    g366_p_spl_1
  );


  buf

  (
    g366_p_spl_100,
    g366_p_spl_10
  );


  buf

  (
    g366_p_spl_101,
    g366_p_spl_10
  );


  buf

  (
    g366_p_spl_11,
    g366_p_spl_1
  );


  buf

  (
    g366_n_spl_,
    g366_n
  );


  buf

  (
    g366_n_spl_0,
    g366_n_spl_
  );


  buf

  (
    g366_n_spl_00,
    g366_n_spl_0
  );


  buf

  (
    g366_n_spl_000,
    g366_n_spl_00
  );


  buf

  (
    g366_n_spl_001,
    g366_n_spl_00
  );


  buf

  (
    g366_n_spl_01,
    g366_n_spl_0
  );


  buf

  (
    g366_n_spl_010,
    g366_n_spl_01
  );


  buf

  (
    g366_n_spl_011,
    g366_n_spl_01
  );


  buf

  (
    g366_n_spl_1,
    g366_n_spl_
  );


  buf

  (
    g366_n_spl_10,
    g366_n_spl_1
  );


  buf

  (
    g366_n_spl_100,
    g366_n_spl_10
  );


  buf

  (
    g366_n_spl_101,
    g366_n_spl_10
  );


  buf

  (
    g366_n_spl_11,
    g366_n_spl_1
  );


  buf

  (
    g367_n_spl_,
    g367_n
  );


  buf

  (
    g367_p_spl_,
    g367_p
  );


  buf

  (
    g371_n_spl_,
    g371_n
  );


  buf

  (
    g371_p_spl_,
    g371_p
  );


  buf

  (
    G47_p_spl_,
    G47_p
  );


  buf

  (
    G47_p_spl_0,
    G47_p_spl_
  );


  buf

  (
    G47_p_spl_00,
    G47_p_spl_0
  );


  buf

  (
    G47_p_spl_01,
    G47_p_spl_0
  );


  buf

  (
    G47_p_spl_1,
    G47_p_spl_
  );


  buf

  (
    G47_p_spl_10,
    G47_p_spl_1
  );


  buf

  (
    g374_p_spl_,
    g374_p
  );


  buf

  (
    g374_p_spl_0,
    g374_p_spl_
  );


  buf

  (
    g374_p_spl_1,
    g374_p_spl_
  );


  buf

  (
    G47_n_spl_,
    G47_n
  );


  buf

  (
    G47_n_spl_0,
    G47_n_spl_
  );


  buf

  (
    G47_n_spl_00,
    G47_n_spl_0
  );


  buf

  (
    G47_n_spl_01,
    G47_n_spl_0
  );


  buf

  (
    G47_n_spl_1,
    G47_n_spl_
  );


  buf

  (
    G47_n_spl_10,
    G47_n_spl_1
  );


  buf

  (
    g374_n_spl_,
    g374_n
  );


  buf

  (
    g374_n_spl_0,
    g374_n_spl_
  );


  buf

  (
    g374_n_spl_1,
    g374_n_spl_
  );


  buf

  (
    g370_n_spl_,
    g370_n
  );


  buf

  (
    g370_n_spl_0,
    g370_n_spl_
  );


  buf

  (
    g370_n_spl_1,
    g370_n_spl_
  );


  buf

  (
    g370_p_spl_,
    g370_p
  );


  buf

  (
    g370_p_spl_0,
    g370_p_spl_
  );


  buf

  (
    g370_p_spl_1,
    g370_p_spl_
  );


  buf

  (
    g76_p_spl_,
    g76_p
  );


  buf

  (
    g377_n_spl_,
    g377_n
  );


  buf

  (
    g377_n_spl_0,
    g377_n_spl_
  );


  buf

  (
    g377_n_spl_00,
    g377_n_spl_0
  );


  buf

  (
    g377_n_spl_01,
    g377_n_spl_0
  );


  buf

  (
    g377_n_spl_1,
    g377_n_spl_
  );


  buf

  (
    g377_n_spl_10,
    g377_n_spl_1
  );


  buf

  (
    g377_n_spl_11,
    g377_n_spl_1
  );


  buf

  (
    g379_p_spl_,
    g379_p
  );


  buf

  (
    g379_p_spl_0,
    g379_p_spl_
  );


  buf

  (
    g379_p_spl_00,
    g379_p_spl_0
  );


  buf

  (
    g379_p_spl_01,
    g379_p_spl_0
  );


  buf

  (
    g379_p_spl_1,
    g379_p_spl_
  );


  buf

  (
    g379_p_spl_10,
    g379_p_spl_1
  );


  buf

  (
    g382_p_spl_,
    g382_p
  );


  buf

  (
    g382_n_spl_,
    g382_n
  );


  buf

  (
    g377_p_spl_,
    g377_p
  );


  buf

  (
    g377_p_spl_0,
    g377_p_spl_
  );


  buf

  (
    g377_p_spl_00,
    g377_p_spl_0
  );


  buf

  (
    g377_p_spl_01,
    g377_p_spl_0
  );


  buf

  (
    g377_p_spl_1,
    g377_p_spl_
  );


  buf

  (
    g377_p_spl_10,
    g377_p_spl_1
  );


  buf

  (
    g384_p_spl_,
    g384_p
  );


  buf

  (
    g384_p_spl_0,
    g384_p_spl_
  );


  buf

  (
    g384_p_spl_00,
    g384_p_spl_0
  );


  buf

  (
    g384_p_spl_01,
    g384_p_spl_0
  );


  buf

  (
    g384_p_spl_1,
    g384_p_spl_
  );


  buf

  (
    g384_p_spl_10,
    g384_p_spl_1
  );


  buf

  (
    g384_n_spl_,
    g384_n
  );


  buf

  (
    g384_n_spl_0,
    g384_n_spl_
  );


  buf

  (
    g384_n_spl_00,
    g384_n_spl_0
  );


  buf

  (
    g384_n_spl_01,
    g384_n_spl_0
  );


  buf

  (
    g384_n_spl_1,
    g384_n_spl_
  );


  buf

  (
    g384_n_spl_10,
    g384_n_spl_1
  );


  buf

  (
    g387_n_spl_,
    g387_n
  );


  buf

  (
    g387_n_spl_0,
    g387_n_spl_
  );


  buf

  (
    g387_p_spl_,
    g387_p
  );


  buf

  (
    g387_p_spl_0,
    g387_p_spl_
  );


  buf

  (
    g385_n_spl_,
    g385_n
  );


  buf

  (
    g385_n_spl_0,
    g385_n_spl_
  );


  buf

  (
    g385_n_spl_00,
    g385_n_spl_0
  );


  buf

  (
    g385_n_spl_000,
    g385_n_spl_00
  );


  buf

  (
    g385_n_spl_001,
    g385_n_spl_00
  );


  buf

  (
    g385_n_spl_01,
    g385_n_spl_0
  );


  buf

  (
    g385_n_spl_1,
    g385_n_spl_
  );


  buf

  (
    g385_n_spl_10,
    g385_n_spl_1
  );


  buf

  (
    g385_n_spl_11,
    g385_n_spl_1
  );


  buf

  (
    g385_p_spl_,
    g385_p
  );


  buf

  (
    g385_p_spl_0,
    g385_p_spl_
  );


  buf

  (
    g385_p_spl_00,
    g385_p_spl_0
  );


  buf

  (
    g385_p_spl_000,
    g385_p_spl_00
  );


  buf

  (
    g385_p_spl_001,
    g385_p_spl_00
  );


  buf

  (
    g385_p_spl_01,
    g385_p_spl_0
  );


  buf

  (
    g385_p_spl_1,
    g385_p_spl_
  );


  buf

  (
    g385_p_spl_10,
    g385_p_spl_1
  );


  buf

  (
    g385_p_spl_11,
    g385_p_spl_1
  );


  buf

  (
    g390_p_spl_,
    g390_p
  );


  buf

  (
    g390_p_spl_0,
    g390_p_spl_
  );


  buf

  (
    g390_p_spl_1,
    g390_p_spl_
  );


  buf

  (
    g390_n_spl_,
    g390_n
  );


  buf

  (
    g390_n_spl_0,
    g390_n_spl_
  );


  buf

  (
    g390_n_spl_1,
    g390_n_spl_
  );


  buf

  (
    g394_n_spl_,
    g394_n
  );


  buf

  (
    g394_n_spl_0,
    g394_n_spl_
  );


  buf

  (
    g394_n_spl_00,
    g394_n_spl_0
  );


  buf

  (
    g394_n_spl_01,
    g394_n_spl_0
  );


  buf

  (
    g394_n_spl_1,
    g394_n_spl_
  );


  buf

  (
    g394_p_spl_,
    g394_p
  );


  buf

  (
    g394_p_spl_0,
    g394_p_spl_
  );


  buf

  (
    g394_p_spl_00,
    g394_p_spl_0
  );


  buf

  (
    g394_p_spl_01,
    g394_p_spl_0
  );


  buf

  (
    g394_p_spl_1,
    g394_p_spl_
  );


  buf

  (
    g55_n_spl_,
    g55_n
  );


  buf

  (
    g393_p_spl_,
    g393_p
  );


  buf

  (
    g393_p_spl_0,
    g393_p_spl_
  );


  buf

  (
    g393_p_spl_00,
    g393_p_spl_0
  );


  buf

  (
    g393_p_spl_000,
    g393_p_spl_00
  );


  buf

  (
    g393_p_spl_001,
    g393_p_spl_00
  );


  buf

  (
    g393_p_spl_01,
    g393_p_spl_0
  );


  buf

  (
    g393_p_spl_010,
    g393_p_spl_01
  );


  buf

  (
    g393_p_spl_011,
    g393_p_spl_01
  );


  buf

  (
    g393_p_spl_1,
    g393_p_spl_
  );


  buf

  (
    g393_p_spl_10,
    g393_p_spl_1
  );


  buf

  (
    g393_p_spl_100,
    g393_p_spl_10
  );


  buf

  (
    g393_p_spl_101,
    g393_p_spl_10
  );


  buf

  (
    g393_p_spl_11,
    g393_p_spl_1
  );


  buf

  (
    g393_p_spl_110,
    g393_p_spl_11
  );


  buf

  (
    g393_p_spl_111,
    g393_p_spl_11
  );


  buf

  (
    g393_n_spl_,
    g393_n
  );


  buf

  (
    g393_n_spl_0,
    g393_n_spl_
  );


  buf

  (
    g393_n_spl_00,
    g393_n_spl_0
  );


  buf

  (
    g393_n_spl_000,
    g393_n_spl_00
  );


  buf

  (
    g393_n_spl_001,
    g393_n_spl_00
  );


  buf

  (
    g393_n_spl_01,
    g393_n_spl_0
  );


  buf

  (
    g393_n_spl_010,
    g393_n_spl_01
  );


  buf

  (
    g393_n_spl_011,
    g393_n_spl_01
  );


  buf

  (
    g393_n_spl_1,
    g393_n_spl_
  );


  buf

  (
    g393_n_spl_10,
    g393_n_spl_1
  );


  buf

  (
    g393_n_spl_100,
    g393_n_spl_10
  );


  buf

  (
    g393_n_spl_101,
    g393_n_spl_10
  );


  buf

  (
    g393_n_spl_11,
    g393_n_spl_1
  );


  buf

  (
    g393_n_spl_110,
    g393_n_spl_11
  );


  buf

  (
    g393_n_spl_111,
    g393_n_spl_11
  );


  buf

  (
    g404_n_spl_,
    g404_n
  );


  buf

  (
    g404_n_spl_0,
    g404_n_spl_
  );


  buf

  (
    g404_p_spl_,
    g404_p
  );


  buf

  (
    g404_p_spl_0,
    g404_p_spl_
  );


  buf

  (
    g403_n_spl_,
    g403_n
  );


  buf

  (
    g403_n_spl_0,
    g403_n_spl_
  );


  buf

  (
    g403_n_spl_1,
    g403_n_spl_
  );


  buf

  (
    g405_p_spl_,
    g405_p
  );


  buf

  (
    g403_p_spl_,
    g403_p
  );


  buf

  (
    g403_p_spl_0,
    g403_p_spl_
  );


  buf

  (
    g403_p_spl_1,
    g403_p_spl_
  );


  buf

  (
    g405_n_spl_,
    g405_n
  );


  buf

  (
    G45_p_spl_,
    G45_p
  );


  buf

  (
    g406_n_spl_,
    g406_n
  );


  buf

  (
    g406_n_spl_0,
    g406_n_spl_
  );


  buf

  (
    g406_n_spl_00,
    g406_n_spl_0
  );


  buf

  (
    g406_n_spl_000,
    g406_n_spl_00
  );


  buf

  (
    g406_n_spl_0000,
    g406_n_spl_000
  );


  buf

  (
    g406_n_spl_001,
    g406_n_spl_00
  );


  buf

  (
    g406_n_spl_01,
    g406_n_spl_0
  );


  buf

  (
    g406_n_spl_010,
    g406_n_spl_01
  );


  buf

  (
    g406_n_spl_011,
    g406_n_spl_01
  );


  buf

  (
    g406_n_spl_1,
    g406_n_spl_
  );


  buf

  (
    g406_n_spl_10,
    g406_n_spl_1
  );


  buf

  (
    g406_n_spl_100,
    g406_n_spl_10
  );


  buf

  (
    g406_n_spl_101,
    g406_n_spl_10
  );


  buf

  (
    g406_n_spl_11,
    g406_n_spl_1
  );


  buf

  (
    g406_n_spl_110,
    g406_n_spl_11
  );


  buf

  (
    g406_n_spl_111,
    g406_n_spl_11
  );


  buf

  (
    G45_n_spl_,
    G45_n
  );


  buf

  (
    g406_p_spl_,
    g406_p
  );


  buf

  (
    g406_p_spl_0,
    g406_p_spl_
  );


  buf

  (
    g406_p_spl_00,
    g406_p_spl_0
  );


  buf

  (
    g406_p_spl_000,
    g406_p_spl_00
  );


  buf

  (
    g406_p_spl_0000,
    g406_p_spl_000
  );


  buf

  (
    g406_p_spl_001,
    g406_p_spl_00
  );


  buf

  (
    g406_p_spl_01,
    g406_p_spl_0
  );


  buf

  (
    g406_p_spl_010,
    g406_p_spl_01
  );


  buf

  (
    g406_p_spl_011,
    g406_p_spl_01
  );


  buf

  (
    g406_p_spl_1,
    g406_p_spl_
  );


  buf

  (
    g406_p_spl_10,
    g406_p_spl_1
  );


  buf

  (
    g406_p_spl_100,
    g406_p_spl_10
  );


  buf

  (
    g406_p_spl_101,
    g406_p_spl_10
  );


  buf

  (
    g406_p_spl_11,
    g406_p_spl_1
  );


  buf

  (
    g406_p_spl_110,
    g406_p_spl_11
  );


  buf

  (
    g406_p_spl_111,
    g406_p_spl_11
  );


  buf

  (
    g408_p_spl_,
    g408_p
  );


  buf

  (
    g408_n_spl_,
    g408_n
  );


  buf

  (
    G44_p_spl_,
    G44_p
  );


  buf

  (
    G44_p_spl_0,
    G44_p_spl_
  );


  buf

  (
    g409_n_spl_,
    g409_n
  );


  buf

  (
    g409_n_spl_0,
    g409_n_spl_
  );


  buf

  (
    g409_n_spl_00,
    g409_n_spl_0
  );


  buf

  (
    g409_n_spl_000,
    g409_n_spl_00
  );


  buf

  (
    g409_n_spl_001,
    g409_n_spl_00
  );


  buf

  (
    g409_n_spl_01,
    g409_n_spl_0
  );


  buf

  (
    g409_n_spl_010,
    g409_n_spl_01
  );


  buf

  (
    g409_n_spl_011,
    g409_n_spl_01
  );


  buf

  (
    g409_n_spl_1,
    g409_n_spl_
  );


  buf

  (
    g409_n_spl_10,
    g409_n_spl_1
  );


  buf

  (
    g409_n_spl_100,
    g409_n_spl_10
  );


  buf

  (
    g409_n_spl_101,
    g409_n_spl_10
  );


  buf

  (
    g409_n_spl_11,
    g409_n_spl_1
  );


  buf

  (
    g409_n_spl_110,
    g409_n_spl_11
  );


  buf

  (
    g409_n_spl_111,
    g409_n_spl_11
  );


  buf

  (
    G44_n_spl_,
    G44_n
  );


  buf

  (
    G44_n_spl_0,
    G44_n_spl_
  );


  buf

  (
    g409_p_spl_,
    g409_p
  );


  buf

  (
    g409_p_spl_0,
    g409_p_spl_
  );


  buf

  (
    g409_p_spl_00,
    g409_p_spl_0
  );


  buf

  (
    g409_p_spl_000,
    g409_p_spl_00
  );


  buf

  (
    g409_p_spl_001,
    g409_p_spl_00
  );


  buf

  (
    g409_p_spl_01,
    g409_p_spl_0
  );


  buf

  (
    g409_p_spl_010,
    g409_p_spl_01
  );


  buf

  (
    g409_p_spl_011,
    g409_p_spl_01
  );


  buf

  (
    g409_p_spl_1,
    g409_p_spl_
  );


  buf

  (
    g409_p_spl_10,
    g409_p_spl_1
  );


  buf

  (
    g409_p_spl_100,
    g409_p_spl_10
  );


  buf

  (
    g409_p_spl_101,
    g409_p_spl_10
  );


  buf

  (
    g409_p_spl_11,
    g409_p_spl_1
  );


  buf

  (
    g409_p_spl_110,
    g409_p_spl_11
  );


  buf

  (
    g409_p_spl_111,
    g409_p_spl_11
  );


  buf

  (
    G42_p_spl_,
    G42_p
  );


  buf

  (
    G42_p_spl_0,
    G42_p_spl_
  );


  buf

  (
    G42_p_spl_1,
    G42_p_spl_
  );


  buf

  (
    g412_n_spl_,
    g412_n
  );


  buf

  (
    g412_n_spl_0,
    g412_n_spl_
  );


  buf

  (
    g412_n_spl_00,
    g412_n_spl_0
  );


  buf

  (
    g412_n_spl_000,
    g412_n_spl_00
  );


  buf

  (
    g412_n_spl_0000,
    g412_n_spl_000
  );


  buf

  (
    g412_n_spl_0001,
    g412_n_spl_000
  );


  buf

  (
    g412_n_spl_001,
    g412_n_spl_00
  );


  buf

  (
    g412_n_spl_0010,
    g412_n_spl_001
  );


  buf

  (
    g412_n_spl_01,
    g412_n_spl_0
  );


  buf

  (
    g412_n_spl_010,
    g412_n_spl_01
  );


  buf

  (
    g412_n_spl_011,
    g412_n_spl_01
  );


  buf

  (
    g412_n_spl_1,
    g412_n_spl_
  );


  buf

  (
    g412_n_spl_10,
    g412_n_spl_1
  );


  buf

  (
    g412_n_spl_100,
    g412_n_spl_10
  );


  buf

  (
    g412_n_spl_101,
    g412_n_spl_10
  );


  buf

  (
    g412_n_spl_11,
    g412_n_spl_1
  );


  buf

  (
    g412_n_spl_110,
    g412_n_spl_11
  );


  buf

  (
    g412_n_spl_111,
    g412_n_spl_11
  );


  buf

  (
    G42_n_spl_,
    G42_n
  );


  buf

  (
    G42_n_spl_0,
    G42_n_spl_
  );


  buf

  (
    G42_n_spl_1,
    G42_n_spl_
  );


  buf

  (
    g412_p_spl_,
    g412_p
  );


  buf

  (
    g412_p_spl_0,
    g412_p_spl_
  );


  buf

  (
    g412_p_spl_00,
    g412_p_spl_0
  );


  buf

  (
    g412_p_spl_000,
    g412_p_spl_00
  );


  buf

  (
    g412_p_spl_0000,
    g412_p_spl_000
  );


  buf

  (
    g412_p_spl_0001,
    g412_p_spl_000
  );


  buf

  (
    g412_p_spl_001,
    g412_p_spl_00
  );


  buf

  (
    g412_p_spl_0010,
    g412_p_spl_001
  );


  buf

  (
    g412_p_spl_01,
    g412_p_spl_0
  );


  buf

  (
    g412_p_spl_010,
    g412_p_spl_01
  );


  buf

  (
    g412_p_spl_011,
    g412_p_spl_01
  );


  buf

  (
    g412_p_spl_1,
    g412_p_spl_
  );


  buf

  (
    g412_p_spl_10,
    g412_p_spl_1
  );


  buf

  (
    g412_p_spl_100,
    g412_p_spl_10
  );


  buf

  (
    g412_p_spl_101,
    g412_p_spl_10
  );


  buf

  (
    g412_p_spl_11,
    g412_p_spl_1
  );


  buf

  (
    g412_p_spl_110,
    g412_p_spl_11
  );


  buf

  (
    g412_p_spl_111,
    g412_p_spl_11
  );


  buf

  (
    g414_n_spl_,
    g414_n
  );


  buf

  (
    g414_n_spl_0,
    g414_n_spl_
  );


  buf

  (
    g414_n_spl_00,
    g414_n_spl_0
  );


  buf

  (
    g414_n_spl_000,
    g414_n_spl_00
  );


  buf

  (
    g414_n_spl_0000,
    g414_n_spl_000
  );


  buf

  (
    g414_n_spl_0001,
    g414_n_spl_000
  );


  buf

  (
    g414_n_spl_001,
    g414_n_spl_00
  );


  buf

  (
    g414_n_spl_01,
    g414_n_spl_0
  );


  buf

  (
    g414_n_spl_010,
    g414_n_spl_01
  );


  buf

  (
    g414_n_spl_011,
    g414_n_spl_01
  );


  buf

  (
    g414_n_spl_1,
    g414_n_spl_
  );


  buf

  (
    g414_n_spl_10,
    g414_n_spl_1
  );


  buf

  (
    g414_n_spl_100,
    g414_n_spl_10
  );


  buf

  (
    g414_n_spl_101,
    g414_n_spl_10
  );


  buf

  (
    g414_n_spl_11,
    g414_n_spl_1
  );


  buf

  (
    g414_n_spl_110,
    g414_n_spl_11
  );


  buf

  (
    g414_n_spl_111,
    g414_n_spl_11
  );


  buf

  (
    g414_p_spl_,
    g414_p
  );


  buf

  (
    g414_p_spl_0,
    g414_p_spl_
  );


  buf

  (
    g414_p_spl_00,
    g414_p_spl_0
  );


  buf

  (
    g414_p_spl_000,
    g414_p_spl_00
  );


  buf

  (
    g414_p_spl_0000,
    g414_p_spl_000
  );


  buf

  (
    g414_p_spl_0001,
    g414_p_spl_000
  );


  buf

  (
    g414_p_spl_001,
    g414_p_spl_00
  );


  buf

  (
    g414_p_spl_01,
    g414_p_spl_0
  );


  buf

  (
    g414_p_spl_010,
    g414_p_spl_01
  );


  buf

  (
    g414_p_spl_011,
    g414_p_spl_01
  );


  buf

  (
    g414_p_spl_1,
    g414_p_spl_
  );


  buf

  (
    g414_p_spl_10,
    g414_p_spl_1
  );


  buf

  (
    g414_p_spl_100,
    g414_p_spl_10
  );


  buf

  (
    g414_p_spl_101,
    g414_p_spl_10
  );


  buf

  (
    g414_p_spl_11,
    g414_p_spl_1
  );


  buf

  (
    g414_p_spl_110,
    g414_p_spl_11
  );


  buf

  (
    g414_p_spl_111,
    g414_p_spl_11
  );


  buf

  (
    G43_p_spl_,
    G43_p
  );


  buf

  (
    G43_p_spl_0,
    G43_p_spl_
  );


  buf

  (
    G43_p_spl_1,
    G43_p_spl_
  );


  buf

  (
    G43_n_spl_,
    G43_n
  );


  buf

  (
    G43_n_spl_0,
    G43_n_spl_
  );


  buf

  (
    G43_n_spl_1,
    G43_n_spl_
  );


  buf

  (
    g416_p_spl_,
    g416_p
  );


  buf

  (
    g416_n_spl_,
    g416_n
  );


  buf

  (
    g423_n_spl_,
    g423_n
  );


  buf

  (
    g423_n_spl_0,
    g423_n_spl_
  );


  buf

  (
    g423_n_spl_00,
    g423_n_spl_0
  );


  buf

  (
    g423_n_spl_000,
    g423_n_spl_00
  );


  buf

  (
    g423_n_spl_001,
    g423_n_spl_00
  );


  buf

  (
    g423_n_spl_01,
    g423_n_spl_0
  );


  buf

  (
    g423_n_spl_010,
    g423_n_spl_01
  );


  buf

  (
    g423_n_spl_011,
    g423_n_spl_01
  );


  buf

  (
    g423_n_spl_1,
    g423_n_spl_
  );


  buf

  (
    g423_n_spl_10,
    g423_n_spl_1
  );


  buf

  (
    g423_n_spl_11,
    g423_n_spl_1
  );


  buf

  (
    g423_p_spl_,
    g423_p
  );


  buf

  (
    g423_p_spl_0,
    g423_p_spl_
  );


  buf

  (
    g423_p_spl_00,
    g423_p_spl_0
  );


  buf

  (
    g423_p_spl_000,
    g423_p_spl_00
  );


  buf

  (
    g423_p_spl_001,
    g423_p_spl_00
  );


  buf

  (
    g423_p_spl_01,
    g423_p_spl_0
  );


  buf

  (
    g423_p_spl_010,
    g423_p_spl_01
  );


  buf

  (
    g423_p_spl_011,
    g423_p_spl_01
  );


  buf

  (
    g423_p_spl_1,
    g423_p_spl_
  );


  buf

  (
    g423_p_spl_10,
    g423_p_spl_1
  );


  buf

  (
    g423_p_spl_11,
    g423_p_spl_1
  );


  buf

  (
    g425_n_spl_,
    g425_n
  );


  buf

  (
    g425_n_spl_0,
    g425_n_spl_
  );


  buf

  (
    g425_n_spl_00,
    g425_n_spl_0
  );


  buf

  (
    g425_n_spl_000,
    g425_n_spl_00
  );


  buf

  (
    g425_n_spl_001,
    g425_n_spl_00
  );


  buf

  (
    g425_n_spl_01,
    g425_n_spl_0
  );


  buf

  (
    g425_n_spl_010,
    g425_n_spl_01
  );


  buf

  (
    g425_n_spl_011,
    g425_n_spl_01
  );


  buf

  (
    g425_n_spl_1,
    g425_n_spl_
  );


  buf

  (
    g425_n_spl_10,
    g425_n_spl_1
  );


  buf

  (
    g425_n_spl_100,
    g425_n_spl_10
  );


  buf

  (
    g425_n_spl_101,
    g425_n_spl_10
  );


  buf

  (
    g425_n_spl_11,
    g425_n_spl_1
  );


  buf

  (
    g425_p_spl_,
    g425_p
  );


  buf

  (
    g425_p_spl_0,
    g425_p_spl_
  );


  buf

  (
    g425_p_spl_00,
    g425_p_spl_0
  );


  buf

  (
    g425_p_spl_000,
    g425_p_spl_00
  );


  buf

  (
    g425_p_spl_001,
    g425_p_spl_00
  );


  buf

  (
    g425_p_spl_01,
    g425_p_spl_0
  );


  buf

  (
    g425_p_spl_010,
    g425_p_spl_01
  );


  buf

  (
    g425_p_spl_011,
    g425_p_spl_01
  );


  buf

  (
    g425_p_spl_1,
    g425_p_spl_
  );


  buf

  (
    g425_p_spl_10,
    g425_p_spl_1
  );


  buf

  (
    g425_p_spl_100,
    g425_p_spl_10
  );


  buf

  (
    g425_p_spl_101,
    g425_p_spl_10
  );


  buf

  (
    g425_p_spl_11,
    g425_p_spl_1
  );


  buf

  (
    g432_n_spl_,
    g432_n
  );


  buf

  (
    g432_p_spl_,
    g432_p
  );


  buf

  (
    g430_n_spl_,
    g430_n
  );


  buf

  (
    g430_p_spl_,
    g430_p
  );


  buf

  (
    g438_n_spl_,
    g438_n
  );


  buf

  (
    g438_p_spl_,
    g438_p
  );


  buf

  (
    g440_n_spl_,
    g440_n
  );


  buf

  (
    g441_n_spl_,
    g441_n
  );


  buf

  (
    g440_p_spl_,
    g440_p
  );


  buf

  (
    g441_p_spl_,
    g441_p
  );


  buf

  (
    g439_p_spl_,
    g439_p
  );


  buf

  (
    g439_n_spl_,
    g439_n
  );


  buf

  (
    g453_n_spl_,
    g453_n
  );


  buf

  (
    g453_p_spl_,
    g453_p
  );


  buf

  (
    g452_p_spl_,
    g452_p
  );


  buf

  (
    g452_p_spl_0,
    g452_p_spl_
  );


  buf

  (
    g452_p_spl_1,
    g452_p_spl_
  );


  buf

  (
    g456_p_spl_,
    g456_p
  );


  buf

  (
    g456_p_spl_0,
    g456_p_spl_
  );


  buf

  (
    g456_p_spl_1,
    g456_p_spl_
  );


  buf

  (
    g452_n_spl_,
    g452_n
  );


  buf

  (
    g452_n_spl_0,
    g452_n_spl_
  );


  buf

  (
    g452_n_spl_1,
    g452_n_spl_
  );


  buf

  (
    g456_n_spl_,
    g456_n
  );


  buf

  (
    g456_n_spl_0,
    g456_n_spl_
  );


  buf

  (
    g456_n_spl_1,
    g456_n_spl_
  );


  buf

  (
    G20_p_spl_,
    G20_p
  );


  buf

  (
    G20_p_spl_0,
    G20_p_spl_
  );


  buf

  (
    G20_p_spl_00,
    G20_p_spl_0
  );


  buf

  (
    G20_p_spl_1,
    G20_p_spl_
  );


  buf

  (
    G20_n_spl_,
    G20_n
  );


  buf

  (
    G20_n_spl_0,
    G20_n_spl_
  );


  buf

  (
    G20_n_spl_00,
    G20_n_spl_0
  );


  buf

  (
    G20_n_spl_1,
    G20_n_spl_
  );


  buf

  (
    G18_p_spl_,
    G18_p
  );


  buf

  (
    G18_p_spl_0,
    G18_p_spl_
  );


  buf

  (
    G18_p_spl_1,
    G18_p_spl_
  );


  buf

  (
    G18_n_spl_,
    G18_n
  );


  buf

  (
    G18_n_spl_0,
    G18_n_spl_
  );


  buf

  (
    G18_n_spl_1,
    G18_n_spl_
  );


  buf

  (
    G19_p_spl_,
    G19_p
  );


  buf

  (
    G19_p_spl_0,
    G19_p_spl_
  );


  buf

  (
    G19_p_spl_00,
    G19_p_spl_0
  );


  buf

  (
    G19_p_spl_1,
    G19_p_spl_
  );


  buf

  (
    G19_n_spl_,
    G19_n
  );


  buf

  (
    G19_n_spl_0,
    G19_n_spl_
  );


  buf

  (
    G19_n_spl_00,
    G19_n_spl_0
  );


  buf

  (
    G19_n_spl_1,
    G19_n_spl_
  );


  buf

  (
    g480_n_spl_,
    g480_n
  );


  buf

  (
    g480_p_spl_,
    g480_p
  );


  buf

  (
    g500_p_spl_,
    g500_p
  );


  buf

  (
    g500_p_spl_0,
    g500_p_spl_
  );


  buf

  (
    g500_n_spl_,
    g500_n
  );


  buf

  (
    g500_n_spl_0,
    g500_n_spl_
  );


  buf

  (
    g379_n_spl_,
    g379_n
  );


  buf

  (
    g379_n_spl_0,
    g379_n_spl_
  );


  buf

  (
    g379_n_spl_00,
    g379_n_spl_0
  );


  buf

  (
    g379_n_spl_01,
    g379_n_spl_0
  );


  buf

  (
    g379_n_spl_1,
    g379_n_spl_
  );


  buf

  (
    g503_n_spl_,
    g503_n
  );


  buf

  (
    g503_p_spl_,
    g503_p
  );


  buf

  (
    g501_p_spl_,
    g501_p
  );


  buf

  (
    g504_p_spl_,
    g504_p
  );


  buf

  (
    g501_n_spl_,
    g501_n
  );


  buf

  (
    g504_n_spl_,
    g504_n
  );


  buf

  (
    g510_n_spl_,
    g510_n
  );


  buf

  (
    g510_p_spl_,
    g510_p
  );


  buf

  (
    g514_n_spl_,
    g514_n
  );


  buf

  (
    g514_p_spl_,
    g514_p
  );


  buf

  (
    g513_p_spl_,
    g513_p
  );


  buf

  (
    g513_p_spl_0,
    g513_p_spl_
  );


  buf

  (
    g513_p_spl_00,
    g513_p_spl_0
  );


  buf

  (
    g513_p_spl_1,
    g513_p_spl_
  );


  buf

  (
    g517_p_spl_,
    g517_p
  );


  buf

  (
    g517_p_spl_0,
    g517_p_spl_
  );


  buf

  (
    g517_p_spl_00,
    g517_p_spl_0
  );


  buf

  (
    g517_p_spl_1,
    g517_p_spl_
  );


  buf

  (
    g513_n_spl_,
    g513_n
  );


  buf

  (
    g513_n_spl_0,
    g513_n_spl_
  );


  buf

  (
    g513_n_spl_00,
    g513_n_spl_0
  );


  buf

  (
    g513_n_spl_1,
    g513_n_spl_
  );


  buf

  (
    g517_n_spl_,
    g517_n
  );


  buf

  (
    g517_n_spl_0,
    g517_n_spl_
  );


  buf

  (
    g517_n_spl_00,
    g517_n_spl_0
  );


  buf

  (
    g517_n_spl_1,
    g517_n_spl_
  );


  buf

  (
    g518_p_spl_,
    g518_p
  );


  buf

  (
    g519_p_spl_,
    g519_p
  );


  buf

  (
    g518_n_spl_,
    g518_n
  );


  buf

  (
    g519_n_spl_,
    g519_n
  );


  buf

  (
    g349_n_spl_,
    g349_n
  );


  buf

  (
    g520_n_spl_,
    g520_n
  );


  buf

  (
    g521_p_spl_,
    g521_p
  );


  buf

  (
    g521_p_spl_0,
    g521_p_spl_
  );


  buf

  (
    g520_p_spl_,
    g520_p
  );


  buf

  (
    g521_n_spl_,
    g521_n
  );


  buf

  (
    g521_n_spl_0,
    g521_n_spl_
  );


  buf

  (
    g528_p_spl_,
    g528_p
  );


  buf

  (
    g528_n_spl_,
    g528_n
  );


  buf

  (
    g530_n_spl_,
    g530_n
  );


  buf

  (
    g530_n_spl_0,
    g530_n_spl_
  );


  buf

  (
    g530_p_spl_,
    g530_p
  );


  buf

  (
    g530_p_spl_0,
    g530_p_spl_
  );


  buf

  (
    g527_n_spl_,
    g527_n
  );


  buf

  (
    g527_n_spl_0,
    g527_n_spl_
  );


  buf

  (
    g534_n_spl_,
    g534_n
  );


  buf

  (
    g534_n_spl_0,
    g534_n_spl_
  );


  buf

  (
    g534_n_spl_1,
    g534_n_spl_
  );


  buf

  (
    g527_p_spl_,
    g527_p
  );


  buf

  (
    g527_p_spl_0,
    g527_p_spl_
  );


  buf

  (
    g534_p_spl_,
    g534_p
  );


  buf

  (
    g534_p_spl_0,
    g534_p_spl_
  );


  buf

  (
    g534_p_spl_1,
    g534_p_spl_
  );


  buf

  (
    g552_n_spl_,
    g552_n
  );


  buf

  (
    g552_p_spl_,
    g552_p
  );


  buf

  (
    g555_p_spl_,
    g555_p
  );


  buf

  (
    g555_p_spl_0,
    g555_p_spl_
  );


  buf

  (
    g555_n_spl_,
    g555_n
  );


  buf

  (
    g555_n_spl_0,
    g555_n_spl_
  );


  buf

  (
    g569_n_spl_,
    g569_n
  );


  buf

  (
    g569_p_spl_,
    g569_p
  );


  buf

  (
    g579_n_spl_,
    g579_n
  );


  buf

  (
    g579_p_spl_,
    g579_p
  );


  buf

  (
    g594_n_spl_,
    g594_n
  );


  buf

  (
    g594_p_spl_,
    g594_p
  );


  buf

  (
    g376_p_spl_,
    g376_p
  );


  buf

  (
    g376_p_spl_0,
    g376_p_spl_
  );


  buf

  (
    g597_n_spl_,
    g597_n
  );


  buf

  (
    g597_n_spl_0,
    g597_n_spl_
  );


  buf

  (
    g597_n_spl_00,
    g597_n_spl_0
  );


  buf

  (
    g597_n_spl_1,
    g597_n_spl_
  );


  buf

  (
    g376_n_spl_,
    g376_n
  );


  buf

  (
    g597_p_spl_,
    g597_p
  );


  buf

  (
    g597_p_spl_0,
    g597_p_spl_
  );


  buf

  (
    g597_p_spl_00,
    g597_p_spl_0
  );


  buf

  (
    g597_p_spl_1,
    g597_p_spl_
  );


  buf

  (
    g600_n_spl_,
    g600_n
  );


  buf

  (
    g600_p_spl_,
    g600_p
  );


  buf

  (
    g601_n_spl_,
    g601_n
  );


  buf

  (
    g601_p_spl_,
    g601_p
  );


  buf

  (
    g603_n_spl_,
    g603_n
  );


  buf

  (
    g603_p_spl_,
    g603_p
  );


  buf

  (
    g605_p_spl_,
    g605_p
  );


  buf

  (
    g605_n_spl_,
    g605_n
  );


  buf

  (
    g598_n_spl_,
    g598_n
  );


  buf

  (
    g608_n_spl_,
    g608_n
  );


  buf

  (
    g598_p_spl_,
    g598_p
  );


  buf

  (
    g608_p_spl_,
    g608_p
  );


  buf

  (
    g613_n_spl_,
    g613_n
  );


  buf

  (
    g613_p_spl_,
    g613_p
  );


  buf

  (
    g617_p_spl_,
    g617_p
  );


  buf

  (
    g617_n_spl_,
    g617_n
  );


  buf

  (
    g616_n_spl_,
    g616_n
  );


  buf

  (
    g616_n_spl_0,
    g616_n_spl_
  );


  buf

  (
    g616_n_spl_1,
    g616_n_spl_
  );


  buf

  (
    g620_n_spl_,
    g620_n
  );


  buf

  (
    g620_n_spl_0,
    g620_n_spl_
  );


  buf

  (
    g620_n_spl_1,
    g620_n_spl_
  );


  buf

  (
    g616_p_spl_,
    g616_p
  );


  buf

  (
    g616_p_spl_0,
    g616_p_spl_
  );


  buf

  (
    g616_p_spl_1,
    g616_p_spl_
  );


  buf

  (
    g620_p_spl_,
    g620_p
  );


  buf

  (
    g620_p_spl_0,
    g620_p_spl_
  );


  buf

  (
    g620_p_spl_1,
    g620_p_spl_
  );


  buf

  (
    g628_n_spl_,
    g628_n
  );


  buf

  (
    g628_n_spl_0,
    g628_n_spl_
  );


  buf

  (
    g628_p_spl_,
    g628_p
  );


  buf

  (
    g628_p_spl_0,
    g628_p_spl_
  );


  buf

  (
    g653_n_spl_,
    g653_n
  );


  buf

  (
    g654_n_spl_,
    g654_n
  );


  buf

  (
    g653_p_spl_,
    g653_p
  );


  buf

  (
    g654_p_spl_,
    g654_p
  );


  buf

  (
    g649_p_spl_,
    g649_p
  );


  buf

  (
    g649_n_spl_,
    g649_n
  );


  buf

  (
    g685_p_spl_,
    g685_p
  );


  buf

  (
    g685_n_spl_,
    g685_n
  );


  buf

  (
    g706_n_spl_,
    g706_n
  );


  buf

  (
    g706_p_spl_,
    g706_p
  );


  buf

  (
    g705_n_spl_,
    g705_n
  );


  buf

  (
    g705_p_spl_,
    g705_p
  );


  buf

  (
    g723_p_spl_,
    g723_p
  );


  buf

  (
    g723_n_spl_,
    g723_n
  );


  buf

  (
    g726_p_spl_,
    g726_p
  );


  buf

  (
    g726_n_spl_,
    g726_n
  );


  buf

  (
    g724_p_spl_,
    g724_p
  );


  buf

  (
    g724_p_spl_0,
    g724_p_spl_
  );


  buf

  (
    g729_p_spl_,
    g729_p
  );


  buf

  (
    g724_n_spl_,
    g724_n
  );


  buf

  (
    g724_n_spl_0,
    g724_n_spl_
  );


  buf

  (
    g729_n_spl_,
    g729_n
  );


  buf

  (
    g730_n_spl_,
    g730_n
  );


  buf

  (
    g730_n_spl_0,
    g730_n_spl_
  );


  buf

  (
    g730_p_spl_,
    g730_p
  );


  buf

  (
    g730_p_spl_0,
    g730_p_spl_
  );


  buf

  (
    g733_p_spl_,
    g733_p
  );


  buf

  (
    g735_n_spl_,
    g735_n
  );


  buf

  (
    g733_n_spl_,
    g733_n
  );


  buf

  (
    g735_p_spl_,
    g735_p
  );


  buf

  (
    g738_n_spl_,
    g738_n
  );


  buf

  (
    g738_n_spl_0,
    g738_n_spl_
  );


  buf

  (
    g738_n_spl_1,
    g738_n_spl_
  );


  buf

  (
    g740_n_spl_,
    g740_n
  );


  buf

  (
    g740_n_spl_0,
    g740_n_spl_
  );


  buf

  (
    g738_p_spl_,
    g738_p
  );


  buf

  (
    g738_p_spl_0,
    g738_p_spl_
  );


  buf

  (
    g738_p_spl_1,
    g738_p_spl_
  );


  buf

  (
    g740_p_spl_,
    g740_p
  );


  buf

  (
    g740_p_spl_0,
    g740_p_spl_
  );


  buf

  (
    g732_p_spl_,
    g732_p
  );


  buf

  (
    g732_p_spl_0,
    g732_p_spl_
  );


  buf

  (
    g732_p_spl_1,
    g732_p_spl_
  );


  buf

  (
    g741_n_spl_,
    g741_n
  );


  buf

  (
    g741_n_spl_0,
    g741_n_spl_
  );


  buf

  (
    g732_n_spl_,
    g732_n
  );


  buf

  (
    g732_n_spl_0,
    g732_n_spl_
  );


  buf

  (
    g732_n_spl_1,
    g732_n_spl_
  );


  buf

  (
    g741_p_spl_,
    g741_p
  );


  buf

  (
    g741_p_spl_0,
    g741_p_spl_
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    G17_p_spl_0,
    G17_p_spl_
  );


  buf

  (
    G17_n_spl_,
    G17_n
  );


  buf

  (
    G17_n_spl_0,
    G17_n_spl_
  );


  buf

  (
    G16_n_spl_,
    G16_n
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    g779_n_spl_,
    g779_n
  );


  buf

  (
    g779_p_spl_,
    g779_p
  );


  buf

  (
    g782_p_spl_,
    g782_p
  );


  buf

  (
    g782_p_spl_0,
    g782_p_spl_
  );


  buf

  (
    g782_n_spl_,
    g782_n
  );


  buf

  (
    g782_n_spl_0,
    g782_n_spl_
  );


  buf

  (
    g818_p_spl_,
    g818_p
  );


  buf

  (
    g818_n_spl_,
    g818_n
  );


  buf

  (
    g626_p_spl_,
    g626_p
  );


  buf

  (
    g722_p_spl_,
    g722_p
  );


  buf

  (
    g626_n_spl_,
    g626_n
  );


  buf

  (
    g626_n_spl_0,
    g626_n_spl_
  );


  buf

  (
    g722_n_spl_,
    g722_n
  );


  buf

  (
    g722_n_spl_0,
    g722_n_spl_
  );


  buf

  (
    g778_p_spl_,
    g778_p
  );


  buf

  (
    g827_p_spl_,
    g827_p
  );


  buf

  (
    g778_n_spl_,
    g778_n
  );


  buf

  (
    g778_n_spl_0,
    g778_n_spl_
  );


  buf

  (
    g827_n_spl_,
    g827_n
  );


  buf

  (
    g827_n_spl_0,
    g827_n_spl_
  );


  buf

  (
    g509_p_spl_,
    g509_p
  );


  buf

  (
    g866_p_spl_,
    g866_p
  );


  buf

  (
    g509_n_spl_,
    g509_n
  );


  buf

  (
    g509_n_spl_0,
    g509_n_spl_
  );


  buf

  (
    g866_n_spl_,
    g866_n
  );


  buf

  (
    g866_n_spl_0,
    g866_n_spl_
  );


  buf

  (
    g451_p_spl_,
    g451_p
  );


  buf

  (
    g679_p_spl_,
    g679_p
  );


  buf

  (
    g451_n_spl_,
    g451_n
  );


  buf

  (
    g451_n_spl_0,
    g451_n_spl_
  );


  buf

  (
    g679_n_spl_,
    g679_n
  );


  buf

  (
    g679_n_spl_0,
    g679_n_spl_
  );


  buf

  (
    g869_n_spl_,
    g869_n
  );


  buf

  (
    g870_n_spl_,
    g870_n
  );


  buf

  (
    g868_n_spl_,
    g868_n
  );


  buf

  (
    g868_n_spl_0,
    g868_n_spl_
  );


  buf

  (
    g867_n_spl_,
    g867_n
  );


  buf

  (
    g874_n_spl_,
    g874_n
  );


  buf

  (
    g873_n_spl_,
    g873_n
  );


  buf

  (
    g879_p_spl_,
    g879_p
  );


  buf

  (
    g881_n_spl_,
    g881_n
  );


  buf

  (
    g879_n_spl_,
    g879_n
  );


  buf

  (
    g881_p_spl_,
    g881_p
  );


  buf

  (
    G50_n_spl_,
    G50_n
  );


  buf

  (
    g888_n_spl_,
    g888_n
  );


  buf

  (
    g888_n_spl_0,
    g888_n_spl_
  );


  buf

  (
    g888_n_spl_1,
    g888_n_spl_
  );


  buf

  (
    G50_p_spl_,
    G50_p
  );


  buf

  (
    g888_p_spl_,
    g888_p
  );


  buf

  (
    g888_p_spl_0,
    g888_p_spl_
  );


  buf

  (
    g888_p_spl_1,
    g888_p_spl_
  );


  buf

  (
    g886_p_spl_,
    g886_p
  );


  buf

  (
    g886_p_spl_0,
    g886_p_spl_
  );


  buf

  (
    g886_p_spl_1,
    g886_p_spl_
  );


  buf

  (
    g892_n_spl_,
    g892_n
  );


  buf

  (
    g886_n_spl_,
    g886_n
  );


  buf

  (
    g886_n_spl_0,
    g886_n_spl_
  );


  buf

  (
    g886_n_spl_1,
    g886_n_spl_
  );


  buf

  (
    g892_p_spl_,
    g892_p
  );


  buf

  (
    g884_n_spl_,
    g884_n
  );


  buf

  (
    g884_p_spl_,
    g884_p
  );


endmodule
