
module mymod
(
  enable,
  reset,
  input_f[0],
  input_f[1],
  input_f[2],
  input_f[3],
  input_f[4],
  input_f[5],
  input_f[6],
  input_f[7],
  input_w[0],
  input_w[1],
  input_w[2],
  input_w[3],
  input_w[4],
  input_w[5],
  input_w[6],
  input_w[7],
  psum_reg[0],
  psum_reg[1],
  psum_reg[2],
  psum_reg[3],
  psum_reg[4],
  psum_reg[5],
  psum_reg[6],
  psum_reg[7],
  output_f[0],
  output_f[1],
  output_f[2],
  output_f[3],
  output_f[4],
  output_f[5],
  output_f[6],
  output_f[7],
  psum_next[0],
  psum_next[1],
  psum_next[2],
  psum_next[3],
  psum_next[4],
  psum_next[5],
  psum_next[6],
  psum_next[7]
);

  input enable;input reset;input input_f[0];input input_f[1];input input_f[2];input input_f[3];input input_f[4];input input_f[5];input input_f[6];input input_f[7];input input_w[0];input input_w[1];input input_w[2];input input_w[3];input input_w[4];input input_w[5];input input_w[6];input input_w[7];input psum_reg[0];input psum_reg[1];input psum_reg[2];input psum_reg[3];input psum_reg[4];input psum_reg[5];input psum_reg[6];input psum_reg[7];
  output output_f[0];output output_f[1];output output_f[2];output output_f[3];output output_f[4];output output_f[5];output output_f[6];output output_f[7];output psum_next[0];output psum_next[1];output psum_next[2];output psum_next[3];output psum_next[4];output psum_next[5];output psum_next[6];output psum_next[7];
  wire enable_p;
  wire enable_n;
  wire reset_p;
  wire reset_n;
  wire input_f[0]_p;
  wire input_f[0]_n;
  wire input_f[1]_p;
  wire input_f[1]_n;
  wire input_f[2]_p;
  wire input_f[2]_n;
  wire input_f[3]_p;
  wire input_f[3]_n;
  wire input_f[4]_p;
  wire input_f[4]_n;
  wire input_f[5]_p;
  wire input_f[5]_n;
  wire input_f[6]_p;
  wire input_f[6]_n;
  wire input_f[7]_p;
  wire input_f[7]_n;
  wire input_w[0]_p;
  wire input_w[0]_n;
  wire input_w[1]_p;
  wire input_w[1]_n;
  wire input_w[2]_p;
  wire input_w[2]_n;
  wire input_w[3]_p;
  wire input_w[3]_n;
  wire input_w[4]_p;
  wire input_w[4]_n;
  wire input_w[5]_p;
  wire input_w[5]_n;
  wire input_w[6]_p;
  wire input_w[6]_n;
  wire input_w[7]_p;
  wire input_w[7]_n;
  wire psum_reg[0]_p;
  wire psum_reg[0]_n;
  wire psum_reg[1]_p;
  wire psum_reg[1]_n;
  wire psum_reg[2]_p;
  wire psum_reg[2]_n;
  wire psum_reg[3]_p;
  wire psum_reg[3]_n;
  wire psum_reg[4]_p;
  wire psum_reg[4]_n;
  wire psum_reg[5]_p;
  wire psum_reg[5]_n;
  wire psum_reg[6]_p;
  wire psum_reg[6]_n;
  wire psum_reg[7]_p;
  wire psum_reg[7]_n;
  wire g27_p;
  wire g27_n;
  wire g28_p;
  wire g28_n;
  wire g29_p;
  wire g29_n;
  wire g30_p;
  wire g30_n;
  wire g31_p;
  wire g31_n;
  wire g32_p;
  wire g32_n;
  wire g33_p;
  wire g33_n;
  wire g34_p;
  wire g34_n;
  wire g35_p;
  wire g35_n;
  wire g36_p;
  wire g36_n;
  wire g37_p;
  wire g37_n;
  wire g38_p;
  wire g38_n;
  wire g39_p;
  wire g39_n;
  wire g40_p;
  wire g40_n;
  wire g41_p;
  wire g41_n;
  wire g42_p;
  wire g42_n;
  wire g43_p;
  wire g43_n;
  wire g44_p;
  wire g44_n;
  wire g45_p;
  wire g45_n;
  wire g46_p;
  wire g46_n;
  wire g47_p;
  wire g47_n;
  wire g48_p;
  wire g48_n;
  wire g49_p;
  wire g49_n;
  wire g50_p;
  wire g50_n;
  wire g51_p;
  wire g51_n;
  wire g52_p;
  wire g52_n;
  wire g53_p;
  wire g53_n;
  wire g54_p;
  wire g54_n;
  wire g55_p;
  wire g55_n;
  wire g56_p;
  wire g56_n;
  wire g57_p;
  wire g57_n;
  wire g58_p;
  wire g58_n;
  wire g59_p;
  wire g59_n;
  wire g60_p;
  wire g60_n;
  wire g61_p;
  wire g61_n;
  wire g62_p;
  wire g62_n;
  wire g63_p;
  wire g63_n;
  wire g64_p;
  wire g64_n;
  wire g65_p;
  wire g65_n;
  wire g66_p;
  wire g66_n;
  wire g67_p;
  wire g67_n;
  wire g68_p;
  wire g68_n;
  wire g69_p;
  wire g69_n;
  wire g70_p;
  wire g70_n;
  wire g71_p;
  wire g71_n;
  wire g72_p;
  wire g72_n;
  wire g73_p;
  wire g73_n;
  wire g74_p;
  wire g74_n;
  wire g75_p;
  wire g75_n;
  wire g76_p;
  wire g76_n;
  wire g77_p;
  wire g77_n;
  wire g78_p;
  wire g78_n;
  wire g79_p;
  wire g79_n;
  wire g80_p;
  wire g80_n;
  wire g81_p;
  wire g81_n;
  wire g82_p;
  wire g82_n;
  wire g83_p;
  wire g83_n;
  wire g84_p;
  wire g84_n;
  wire g85_p;
  wire g85_n;
  wire g86_p;
  wire g86_n;
  wire g87_p;
  wire g87_n;
  wire g88_p;
  wire g88_n;
  wire g89_p;
  wire g89_n;
  wire g90_p;
  wire g90_n;
  wire g91_p;
  wire g91_n;
  wire g92_p;
  wire g92_n;
  wire g93_p;
  wire g93_n;
  wire g94_p;
  wire g94_n;
  wire g95_p;
  wire g95_n;
  wire g96_p;
  wire g96_n;
  wire g97_p;
  wire g97_n;
  wire g98_p;
  wire g98_n;
  wire g99_p;
  wire g99_n;
  wire g100_p;
  wire g100_n;
  wire g101_p;
  wire g101_n;
  wire g102_p;
  wire g102_n;
  wire g103_p;
  wire g103_n;
  wire g104_p;
  wire g104_n;
  wire g105_p;
  wire g105_n;
  wire g106_p;
  wire g106_n;
  wire g107_p;
  wire g107_n;
  wire g108_p;
  wire g108_n;
  wire g109_p;
  wire g109_n;
  wire g110_p;
  wire g110_n;
  wire g111_p;
  wire g111_n;
  wire g112_p;
  wire g112_n;
  wire g113_p;
  wire g113_n;
  wire g114_p;
  wire g114_n;
  wire g115_p;
  wire g115_n;
  wire g116_p;
  wire g116_n;
  wire g117_p;
  wire g117_n;
  wire g118_p;
  wire g118_n;
  wire g119_p;
  wire g119_n;
  wire g120_p;
  wire g120_n;
  wire g121_p;
  wire g121_n;
  wire g122_p;
  wire g122_n;
  wire g123_p;
  wire g123_n;
  wire g124_p;
  wire g124_n;
  wire g125_p;
  wire g125_n;
  wire g126_p;
  wire g126_n;
  wire g127_p;
  wire g127_n;
  wire g128_p;
  wire g128_n;
  wire g129_p;
  wire g129_n;
  wire g130_p;
  wire g130_n;
  wire g131_p;
  wire g131_n;
  wire g132_p;
  wire g132_n;
  wire g133_p;
  wire g133_n;
  wire g134_p;
  wire g134_n;
  wire g135_p;
  wire g135_n;
  wire g136_p;
  wire g136_n;
  wire g137_p;
  wire g137_n;
  wire g138_p;
  wire g138_n;
  wire g139_p;
  wire g139_n;
  wire g140_p;
  wire g140_n;
  wire g141_p;
  wire g141_n;
  wire g142_p;
  wire g142_n;
  wire g143_p;
  wire g143_n;
  wire g144_p;
  wire g144_n;
  wire g145_p;
  wire g145_n;
  wire g146_p;
  wire g146_n;
  wire g147_p;
  wire g147_n;
  wire g148_p;
  wire g148_n;
  wire g149_p;
  wire g149_n;
  wire g150_p;
  wire g150_n;
  wire g151_p;
  wire g151_n;
  wire g152_p;
  wire g152_n;
  wire g153_p;
  wire g153_n;
  wire g154_p;
  wire g154_n;
  wire g155_p;
  wire g155_n;
  wire g156_p;
  wire g156_n;
  wire g157_p;
  wire g157_n;
  wire g158_p;
  wire g158_n;
  wire g159_p;
  wire g159_n;
  wire g160_p;
  wire g160_n;
  wire g161_p;
  wire g161_n;
  wire g162_p;
  wire g162_n;
  wire g163_p;
  wire g163_n;
  wire g164_p;
  wire g164_n;
  wire g165_p;
  wire g165_n;
  wire g166_p;
  wire g166_n;
  wire g167_p;
  wire g167_n;
  wire g168_p;
  wire g168_n;
  wire g169_p;
  wire g169_n;
  wire g170_p;
  wire g170_n;
  wire g171_p;
  wire g171_n;
  wire g172_p;
  wire g172_n;
  wire g173_p;
  wire g173_n;
  wire g174_p;
  wire g174_n;
  wire g175_p;
  wire g175_n;
  wire g176_p;
  wire g176_n;
  wire g177_p;
  wire g177_n;
  wire g178_p;
  wire g178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire reset_n_spl_;
  wire reset_n_spl_0;
  wire reset_n_spl_00;
  wire reset_n_spl_01;
  wire reset_n_spl_1;
  wire reset_n_spl_10;
  wire reset_n_spl_11;
  wire reset_p_spl_;
  wire reset_p_spl_0;
  wire reset_p_spl_00;
  wire reset_p_spl_01;
  wire reset_p_spl_1;
  wire reset_p_spl_10;
  wire reset_p_spl_11;
  wire enable_n_spl_;
  wire enable_n_spl_0;
  wire enable_n_spl_00;
  wire enable_n_spl_01;
  wire enable_n_spl_1;
  wire enable_n_spl_10;
  wire enable_n_spl_11;
  wire g27_p_spl_;
  wire g27_p_spl_0;
  wire input_f[7]_p_spl_;
  wire input_f[7]_p_spl_0;
  wire input_f[7]_p_spl_00;
  wire input_f[7]_p_spl_01;
  wire input_f[7]_p_spl_1;
  wire input_f[7]_p_spl_10;
  wire input_f[7]_p_spl_11;
  wire input_w[0]_p_spl_;
  wire input_w[0]_p_spl_0;
  wire input_w[0]_p_spl_00;
  wire input_w[0]_p_spl_000;
  wire input_w[0]_p_spl_01;
  wire input_w[0]_p_spl_1;
  wire input_w[0]_p_spl_10;
  wire input_w[0]_p_spl_11;
  wire input_f[7]_n_spl_;
  wire input_f[7]_n_spl_0;
  wire input_f[7]_n_spl_00;
  wire input_f[7]_n_spl_01;
  wire input_f[7]_n_spl_1;
  wire input_f[7]_n_spl_10;
  wire input_f[7]_n_spl_11;
  wire input_w[0]_n_spl_;
  wire input_w[0]_n_spl_0;
  wire input_w[0]_n_spl_00;
  wire input_w[0]_n_spl_000;
  wire input_w[0]_n_spl_01;
  wire input_w[0]_n_spl_1;
  wire input_w[0]_n_spl_10;
  wire input_w[0]_n_spl_11;
  wire input_w[1]_p_spl_;
  wire input_w[1]_p_spl_0;
  wire input_w[1]_p_spl_00;
  wire input_w[1]_p_spl_000;
  wire input_w[1]_p_spl_01;
  wire input_w[1]_p_spl_1;
  wire input_w[1]_p_spl_10;
  wire input_w[1]_p_spl_11;
  wire g29_p_spl_;
  wire g29_p_spl_0;
  wire input_w[1]_n_spl_;
  wire input_w[1]_n_spl_0;
  wire input_w[1]_n_spl_00;
  wire input_w[1]_n_spl_000;
  wire input_w[1]_n_spl_01;
  wire input_w[1]_n_spl_1;
  wire input_w[1]_n_spl_10;
  wire input_w[1]_n_spl_11;
  wire g29_n_spl_;
  wire g29_n_spl_0;
  wire input_w[2]_p_spl_;
  wire input_w[2]_p_spl_0;
  wire input_w[2]_p_spl_00;
  wire input_w[2]_p_spl_000;
  wire input_w[2]_p_spl_01;
  wire input_w[2]_p_spl_1;
  wire input_w[2]_p_spl_10;
  wire input_w[2]_p_spl_11;
  wire g30_p_spl_;
  wire g30_p_spl_0;
  wire input_w[2]_n_spl_;
  wire input_w[2]_n_spl_0;
  wire input_w[2]_n_spl_00;
  wire input_w[2]_n_spl_000;
  wire input_w[2]_n_spl_01;
  wire input_w[2]_n_spl_1;
  wire input_w[2]_n_spl_10;
  wire input_w[2]_n_spl_11;
  wire g30_n_spl_;
  wire g30_n_spl_0;
  wire g32_n_spl_;
  wire g34_n_spl_;
  wire g34_n_spl_0;
  wire g32_p_spl_;
  wire g34_p_spl_;
  wire g34_p_spl_0;
  wire g31_n_spl_;
  wire g31_n_spl_0;
  wire g31_n_spl_00;
  wire g31_n_spl_01;
  wire g31_n_spl_1;
  wire g35_n_spl_;
  wire g35_n_spl_0;
  wire g31_p_spl_;
  wire g31_p_spl_0;
  wire g31_p_spl_00;
  wire g31_p_spl_01;
  wire g31_p_spl_1;
  wire g35_p_spl_;
  wire g35_p_spl_0;
  wire input_f[5]_p_spl_;
  wire input_f[5]_p_spl_0;
  wire input_f[5]_p_spl_00;
  wire input_f[5]_p_spl_01;
  wire input_f[5]_p_spl_1;
  wire input_f[5]_p_spl_10;
  wire input_f[5]_p_spl_11;
  wire input_w[5]_p_spl_;
  wire input_w[5]_p_spl_0;
  wire input_w[5]_p_spl_00;
  wire input_w[5]_p_spl_01;
  wire input_w[5]_p_spl_1;
  wire input_w[5]_p_spl_10;
  wire input_w[5]_p_spl_11;
  wire input_f[5]_n_spl_;
  wire input_f[5]_n_spl_0;
  wire input_f[5]_n_spl_00;
  wire input_f[5]_n_spl_01;
  wire input_f[5]_n_spl_1;
  wire input_f[5]_n_spl_10;
  wire input_f[5]_n_spl_11;
  wire input_w[5]_n_spl_;
  wire input_w[5]_n_spl_0;
  wire input_w[5]_n_spl_00;
  wire input_w[5]_n_spl_01;
  wire input_w[5]_n_spl_1;
  wire input_w[5]_n_spl_10;
  wire input_w[5]_n_spl_11;
  wire input_w[3]_p_spl_;
  wire input_w[3]_p_spl_0;
  wire input_w[3]_p_spl_00;
  wire input_w[3]_p_spl_000;
  wire input_w[3]_p_spl_01;
  wire input_w[3]_p_spl_1;
  wire input_w[3]_p_spl_10;
  wire input_w[3]_p_spl_11;
  wire input_w[3]_n_spl_;
  wire input_w[3]_n_spl_0;
  wire input_w[3]_n_spl_00;
  wire input_w[3]_n_spl_000;
  wire input_w[3]_n_spl_01;
  wire input_w[3]_n_spl_1;
  wire input_w[3]_n_spl_10;
  wire input_w[3]_n_spl_11;
  wire input_f[6]_p_spl_;
  wire input_f[6]_p_spl_0;
  wire input_f[6]_p_spl_00;
  wire input_f[6]_p_spl_01;
  wire input_f[6]_p_spl_1;
  wire input_f[6]_p_spl_10;
  wire input_f[6]_p_spl_11;
  wire input_w[4]_p_spl_;
  wire input_w[4]_p_spl_0;
  wire input_w[4]_p_spl_00;
  wire input_w[4]_p_spl_000;
  wire input_w[4]_p_spl_01;
  wire input_w[4]_p_spl_1;
  wire input_w[4]_p_spl_10;
  wire input_w[4]_p_spl_11;
  wire input_f[6]_n_spl_;
  wire input_f[6]_n_spl_0;
  wire input_f[6]_n_spl_00;
  wire input_f[6]_n_spl_01;
  wire input_f[6]_n_spl_1;
  wire input_f[6]_n_spl_10;
  wire input_f[6]_n_spl_11;
  wire input_w[4]_n_spl_;
  wire input_w[4]_n_spl_0;
  wire input_w[4]_n_spl_00;
  wire input_w[4]_n_spl_000;
  wire input_w[4]_n_spl_01;
  wire input_w[4]_n_spl_1;
  wire input_w[4]_n_spl_10;
  wire input_w[4]_n_spl_11;
  wire g38_p_spl_;
  wire g38_p_spl_0;
  wire g39_p_spl_;
  wire g39_p_spl_0;
  wire g38_n_spl_;
  wire g38_n_spl_0;
  wire g39_n_spl_;
  wire g39_n_spl_0;
  wire g40_n_spl_;
  wire g40_p_spl_;
  wire g37_p_spl_;
  wire g42_p_spl_;
  wire g37_n_spl_;
  wire g42_n_spl_;
  wire g43_n_spl_;
  wire g43_p_spl_;
  wire g36_p_spl_;
  wire g36_p_spl_0;
  wire g36_p_spl_00;
  wire g36_p_spl_01;
  wire g36_p_spl_1;
  wire g45_p_spl_;
  wire g36_n_spl_;
  wire g36_n_spl_0;
  wire g36_n_spl_00;
  wire g36_n_spl_01;
  wire g36_n_spl_1;
  wire g45_n_spl_;
  wire g46_n_spl_;
  wire g46_p_spl_;
  wire g49_n_spl_;
  wire g49_n_spl_0;
  wire g49_p_spl_;
  wire g49_p_spl_0;
  wire g51_p_spl_;
  wire g51_p_spl_0;
  wire g51_p_spl_1;
  wire g52_p_spl_;
  wire g51_n_spl_;
  wire g51_n_spl_0;
  wire g51_n_spl_1;
  wire g52_n_spl_;
  wire g53_n_spl_;
  wire g53_p_spl_;
  wire g55_p_spl_;
  wire g55_n_spl_;
  wire g56_n_spl_;
  wire g56_p_spl_;
  wire g47_n_spl_;
  wire g58_p_spl_;
  wire g47_p_spl_;
  wire g58_n_spl_;
  wire input_f[4]_p_spl_;
  wire input_f[4]_p_spl_0;
  wire input_f[4]_p_spl_00;
  wire input_f[4]_p_spl_01;
  wire input_f[4]_p_spl_1;
  wire input_f[4]_p_spl_10;
  wire input_f[4]_p_spl_11;
  wire input_w[6]_p_spl_;
  wire input_w[6]_p_spl_0;
  wire input_w[6]_p_spl_00;
  wire input_w[6]_p_spl_01;
  wire input_w[6]_p_spl_1;
  wire input_w[6]_p_spl_10;
  wire input_w[6]_p_spl_11;
  wire input_f[4]_n_spl_;
  wire input_f[4]_n_spl_0;
  wire input_f[4]_n_spl_00;
  wire input_f[4]_n_spl_01;
  wire input_f[4]_n_spl_1;
  wire input_f[4]_n_spl_10;
  wire input_f[4]_n_spl_11;
  wire input_w[6]_n_spl_;
  wire input_w[6]_n_spl_0;
  wire input_w[6]_n_spl_00;
  wire input_w[6]_n_spl_01;
  wire input_w[6]_n_spl_1;
  wire input_w[6]_n_spl_10;
  wire input_w[6]_n_spl_11;
  wire input_f[3]_n_spl_;
  wire input_f[3]_n_spl_0;
  wire input_f[3]_n_spl_00;
  wire input_f[3]_n_spl_01;
  wire input_f[3]_n_spl_1;
  wire input_f[3]_n_spl_10;
  wire input_f[3]_n_spl_11;
  wire input_w[7]_p_spl_;
  wire input_w[7]_p_spl_0;
  wire input_w[7]_p_spl_00;
  wire input_w[7]_p_spl_000;
  wire input_w[7]_p_spl_001;
  wire input_w[7]_p_spl_01;
  wire input_w[7]_p_spl_1;
  wire input_w[7]_p_spl_10;
  wire input_w[7]_p_spl_11;
  wire input_f[3]_p_spl_;
  wire input_f[3]_p_spl_0;
  wire input_f[3]_p_spl_00;
  wire input_f[3]_p_spl_01;
  wire input_f[3]_p_spl_1;
  wire input_f[3]_p_spl_10;
  wire input_f[3]_p_spl_11;
  wire input_w[7]_n_spl_;
  wire input_w[7]_n_spl_0;
  wire input_w[7]_n_spl_00;
  wire input_w[7]_n_spl_000;
  wire input_w[7]_n_spl_001;
  wire input_w[7]_n_spl_01;
  wire input_w[7]_n_spl_1;
  wire input_w[7]_n_spl_10;
  wire input_w[7]_n_spl_11;
  wire g60_p_spl_;
  wire g61_p_spl_;
  wire g60_n_spl_;
  wire g61_n_spl_;
  wire g64_p_spl_;
  wire g65_p_spl_;
  wire g64_n_spl_;
  wire g65_n_spl_;
  wire g66_n_spl_;
  wire g66_n_spl_0;
  wire g66_p_spl_;
  wire g66_p_spl_0;
  wire g63_n_spl_;
  wire g68_p_spl_;
  wire g63_p_spl_;
  wire g68_n_spl_;
  wire g69_n_spl_;
  wire g69_p_spl_;
  wire g62_p_spl_;
  wire g62_p_spl_0;
  wire g71_p_spl_;
  wire g62_n_spl_;
  wire g62_n_spl_0;
  wire g71_n_spl_;
  wire g72_n_spl_;
  wire g72_p_spl_;
  wire g59_n_spl_;
  wire g59_p_spl_;
  wire g74_p_spl_;
  wire g76_p_spl_;
  wire g74_n_spl_;
  wire g76_n_spl_;
  wire g77_n_spl_;
  wire g77_p_spl_;
  wire g80_p_spl_;
  wire g81_p_spl_;
  wire g80_n_spl_;
  wire g81_n_spl_;
  wire g82_n_spl_;
  wire g82_n_spl_0;
  wire g82_p_spl_;
  wire g82_p_spl_0;
  wire g79_n_spl_;
  wire g84_p_spl_;
  wire g79_p_spl_;
  wire g84_n_spl_;
  wire g85_n_spl_;
  wire g85_p_spl_;
  wire g87_p_spl_;
  wire g87_n_spl_;
  wire g88_n_spl_;
  wire g88_p_spl_;
  wire g92_p_spl_;
  wire g92_n_spl_;
  wire g93_n_spl_;
  wire g93_p_spl_;
  wire g95_p_spl_;
  wire g95_p_spl_0;
  wire g95_p_spl_1;
  wire g95_n_spl_;
  wire g95_n_spl_0;
  wire g95_n_spl_1;
  wire g91_n_spl_;
  wire g98_n_spl_;
  wire g91_p_spl_;
  wire g98_p_spl_;
  wire g99_n_spl_;
  wire g99_p_spl_;
  wire g90_p_spl_;
  wire g101_p_spl_;
  wire g90_n_spl_;
  wire g101_n_spl_;
  wire g102_n_spl_;
  wire g102_p_spl_;
  wire g78_n_spl_;
  wire g104_p_spl_;
  wire g78_p_spl_;
  wire g104_n_spl_;
  wire g105_n_spl_;
  wire g105_p_spl_;
  wire g106_n_spl_;
  wire g108_p_spl_;
  wire g106_p_spl_;
  wire g108_n_spl_;
  wire g109_n_spl_;
  wire g109_p_spl_;
  wire g113_n_spl_;
  wire g113_n_spl_0;
  wire g113_p_spl_;
  wire g113_p_spl_0;
  wire g117_p_spl_;
  wire g118_n_spl_;
  wire g117_n_spl_;
  wire g118_p_spl_;
  wire g119_n_spl_;
  wire g119_p_spl_;
  wire g116_n_spl_;
  wire g116_n_spl_0;
  wire g116_n_spl_1;
  wire g121_n_spl_;
  wire g116_p_spl_;
  wire g116_p_spl_0;
  wire g116_p_spl_1;
  wire g121_p_spl_;
  wire g122_n_spl_;
  wire g122_p_spl_;
  wire g124_p_spl_;
  wire g124_n_spl_;
  wire g125_n_spl_;
  wire g125_p_spl_;
  wire g115_p_spl_;
  wire g115_p_spl_0;
  wire g115_p_spl_1;
  wire g127_p_spl_;
  wire g115_n_spl_;
  wire g115_n_spl_0;
  wire g115_n_spl_1;
  wire g127_n_spl_;
  wire g128_n_spl_;
  wire g128_p_spl_;
  wire g112_n_spl_;
  wire g130_p_spl_;
  wire g112_p_spl_;
  wire g130_n_spl_;
  wire g131_n_spl_;
  wire g131_p_spl_;
  wire g111_n_spl_;
  wire g133_p_spl_;
  wire g111_p_spl_;
  wire g133_n_spl_;
  wire g134_n_spl_;
  wire g134_p_spl_;
  wire g110_n_spl_;
  wire g136_p_spl_;
  wire g110_p_spl_;
  wire g136_n_spl_;
  wire g139_p_spl_;
  wire g139_p_spl_0;
  wire g139_p_spl_1;
  wire g139_n_spl_;
  wire g139_n_spl_0;
  wire g139_n_spl_1;
  wire g140_n_spl_;
  wire g140_p_spl_;
  wire g138_p_spl_;
  wire g144_p_spl_;
  wire g138_n_spl_;
  wire g144_n_spl_;
  wire g145_n_spl_;
  wire g145_p_spl_;
  wire g148_n_spl_;
  wire g148_n_spl_0;
  wire g148_p_spl_;
  wire g148_p_spl_0;
  wire g147_p_spl_;
  wire g153_p_spl_;
  wire g147_n_spl_;
  wire g153_n_spl_;
  wire g154_n_spl_;
  wire g154_p_spl_;
  wire g155_n_spl_;
  wire g157_p_spl_;
  wire g155_p_spl_;
  wire g157_n_spl_;
  wire input_f[2]_n_spl_;
  wire input_f[2]_n_spl_0;
  wire input_f[2]_n_spl_00;
  wire input_f[2]_n_spl_01;
  wire input_f[2]_n_spl_1;
  wire input_f[2]_n_spl_10;
  wire input_f[2]_n_spl_11;
  wire input_f[2]_p_spl_;
  wire input_f[2]_p_spl_0;
  wire input_f[2]_p_spl_00;
  wire input_f[2]_p_spl_01;
  wire input_f[2]_p_spl_1;
  wire input_f[2]_p_spl_10;
  wire input_f[2]_p_spl_11;
  wire g159_p_spl_;
  wire g160_p_spl_;
  wire g159_n_spl_;
  wire g160_n_spl_;
  wire g162_n_spl_;
  wire g164_p_spl_;
  wire g162_p_spl_;
  wire g164_n_spl_;
  wire g165_n_spl_;
  wire g165_p_spl_;
  wire g161_p_spl_;
  wire g161_p_spl_0;
  wire g167_p_spl_;
  wire g161_n_spl_;
  wire g161_n_spl_0;
  wire g167_n_spl_;
  wire g168_n_spl_;
  wire g168_p_spl_;
  wire g158_n_spl_;
  wire g158_p_spl_;
  wire g170_p_spl_;
  wire g172_p_spl_;
  wire g170_n_spl_;
  wire g172_n_spl_;
  wire g173_n_spl_;
  wire g173_p_spl_;
  wire g174_n_spl_;
  wire g176_p_spl_;
  wire g174_p_spl_;
  wire g176_n_spl_;
  wire g177_n_spl_;
  wire g177_p_spl_;
  wire g178_n_spl_;
  wire g180_p_spl_;
  wire g178_p_spl_;
  wire g180_n_spl_;
  wire g181_n_spl_;
  wire g181_p_spl_;
  wire g182_n_spl_;
  wire g184_p_spl_;
  wire g182_p_spl_;
  wire g184_n_spl_;
  wire g186_n_spl_;
  wire g186_p_spl_;
  wire g187_p_spl_;
  wire g187_p_spl_0;
  wire g189_p_spl_;
  wire g187_n_spl_;
  wire g187_n_spl_0;
  wire g189_n_spl_;
  wire g190_n_spl_;
  wire g190_p_spl_;
  wire g192_p_spl_;
  wire g192_n_spl_;
  wire g191_n_spl_;
  wire g195_n_spl_;
  wire g191_p_spl_;
  wire g195_p_spl_;
  wire g198_p_spl_;
  wire g198_n_spl_;
  wire g199_n_spl_;
  wire g199_p_spl_;
  wire g197_p_spl_;
  wire g201_p_spl_;
  wire g197_n_spl_;
  wire g201_n_spl_;
  wire g202_n_spl_;
  wire g202_p_spl_;
  wire g196_n_spl_;
  wire g196_p_spl_;
  wire g204_p_spl_;
  wire g206_p_spl_;
  wire g204_n_spl_;
  wire g206_n_spl_;
  wire g207_n_spl_;
  wire g207_p_spl_;
  wire g208_n_spl_;
  wire g210_p_spl_;
  wire g208_p_spl_;
  wire g210_n_spl_;
  wire input_f[1]_n_spl_;
  wire input_f[1]_n_spl_0;
  wire input_f[1]_n_spl_00;
  wire input_f[1]_n_spl_01;
  wire input_f[1]_n_spl_1;
  wire input_f[1]_n_spl_10;
  wire input_f[1]_n_spl_11;
  wire input_f[1]_p_spl_;
  wire input_f[1]_p_spl_0;
  wire input_f[1]_p_spl_00;
  wire input_f[1]_p_spl_01;
  wire input_f[1]_p_spl_1;
  wire input_f[1]_p_spl_10;
  wire input_f[1]_p_spl_11;
  wire g212_p_spl_;
  wire g212_p_spl_0;
  wire g213_p_spl_;
  wire g212_n_spl_;
  wire g212_n_spl_0;
  wire g213_n_spl_;
  wire g215_n_spl_;
  wire g217_p_spl_;
  wire g215_p_spl_;
  wire g217_n_spl_;
  wire g218_n_spl_;
  wire g218_p_spl_;
  wire g214_p_spl_;
  wire g214_p_spl_0;
  wire g220_p_spl_;
  wire g214_n_spl_;
  wire g214_n_spl_0;
  wire g220_n_spl_;
  wire g221_n_spl_;
  wire g221_p_spl_;
  wire g211_n_spl_;
  wire g211_p_spl_;
  wire g223_p_spl_;
  wire g225_p_spl_;
  wire g223_n_spl_;
  wire g225_n_spl_;
  wire g226_n_spl_;
  wire g226_p_spl_;
  wire g227_n_spl_;
  wire g229_p_spl_;
  wire g227_p_spl_;
  wire g229_n_spl_;
  wire g230_n_spl_;
  wire g230_p_spl_;
  wire g231_n_spl_;
  wire g233_p_spl_;
  wire g231_p_spl_;
  wire g233_n_spl_;
  wire g234_n_spl_;
  wire g234_p_spl_;
  wire g235_n_spl_;
  wire g237_p_spl_;
  wire g235_p_spl_;
  wire g237_n_spl_;
  wire g238_n_spl_;
  wire g238_p_spl_;
  wire g241_p_spl_;
  wire g241_p_spl_0;
  wire g241_n_spl_;
  wire g241_n_spl_0;
  wire g242_n_spl_;
  wire g242_p_spl_;
  wire g243_p_spl_;
  wire g243_p_spl_0;
  wire g247_p_spl_;
  wire g243_n_spl_;
  wire g243_n_spl_0;
  wire g247_n_spl_;
  wire g248_n_spl_;
  wire g248_p_spl_;
  wire g249_n_spl_;
  wire g251_p_spl_;
  wire g249_p_spl_;
  wire g251_n_spl_;
  wire g252_n_spl_;
  wire g252_p_spl_;
  wire g256_n_spl_;
  wire g256_p_spl_;
  wire g255_p_spl_;
  wire g255_p_spl_0;
  wire g260_p_spl_;
  wire g255_n_spl_;
  wire g255_n_spl_0;
  wire g260_n_spl_;
  wire g261_n_spl_;
  wire g261_p_spl_;
  wire g254_p_spl_;
  wire g263_p_spl_;
  wire g254_n_spl_;
  wire g263_n_spl_;
  wire g264_n_spl_;
  wire g264_p_spl_;
  wire g265_n_spl_;
  wire g267_p_spl_;
  wire g265_p_spl_;
  wire g267_n_spl_;
  wire g269_p_spl_;
  wire g269_p_spl_0;
  wire g269_n_spl_;
  wire g269_n_spl_0;
  wire input_f[0]_n_spl_;
  wire input_f[0]_n_spl_0;
  wire input_f[0]_n_spl_00;
  wire input_f[0]_n_spl_01;
  wire input_f[0]_n_spl_1;
  wire input_f[0]_n_spl_10;
  wire input_f[0]_n_spl_11;
  wire input_f[0]_p_spl_;
  wire input_f[0]_p_spl_0;
  wire input_f[0]_p_spl_00;
  wire input_f[0]_p_spl_01;
  wire input_f[0]_p_spl_1;
  wire input_f[0]_p_spl_10;
  wire input_f[0]_p_spl_11;
  wire g270_n_spl_;
  wire g270_p_spl_;
  wire g271_p_spl_;
  wire g275_p_spl_;
  wire g271_n_spl_;
  wire g275_n_spl_;
  wire g276_n_spl_;
  wire g276_p_spl_;
  wire g278_n_spl_;
  wire g280_p_spl_;
  wire g278_p_spl_;
  wire g280_n_spl_;
  wire g281_n_spl_;
  wire g281_p_spl_;
  wire g277_n_spl_;
  wire g283_p_spl_;
  wire g277_p_spl_;
  wire g283_n_spl_;
  wire g284_n_spl_;
  wire g284_p_spl_;
  wire g268_n_spl_;
  wire g268_p_spl_;
  wire g286_p_spl_;
  wire g288_p_spl_;
  wire g286_n_spl_;
  wire g288_n_spl_;
  wire g289_n_spl_;
  wire g289_p_spl_;
  wire g290_n_spl_;
  wire g292_p_spl_;
  wire g290_p_spl_;
  wire g292_n_spl_;
  wire g293_n_spl_;
  wire g293_p_spl_;
  wire g294_n_spl_;
  wire g296_p_spl_;
  wire g294_p_spl_;
  wire g296_n_spl_;
  wire g297_n_spl_;
  wire g297_p_spl_;
  wire g298_n_spl_;
  wire g300_p_spl_;
  wire g298_p_spl_;
  wire g300_n_spl_;
  wire g301_n_spl_;
  wire g301_p_spl_;
  wire g304_p_spl_;
  wire g304_n_spl_;
  wire g305_n_spl_;
  wire g305_p_spl_;
  wire g306_p_spl_;
  wire g308_p_spl_;
  wire g306_n_spl_;
  wire g308_n_spl_;
  wire g309_n_spl_;
  wire g309_p_spl_;
  wire g310_n_spl_;
  wire g312_p_spl_;
  wire g310_p_spl_;
  wire g312_n_spl_;
  wire g314_p_spl_;
  wire g314_p_spl_0;
  wire g314_n_spl_;
  wire g314_n_spl_0;
  wire g315_n_spl_;
  wire g315_p_spl_;
  wire g319_p_spl_;
  wire g319_n_spl_;
  wire g320_n_spl_;
  wire g320_p_spl_;
  wire g313_n_spl_;
  wire g313_p_spl_;
  wire g322_p_spl_;
  wire g324_p_spl_;
  wire g322_n_spl_;
  wire g324_n_spl_;
  wire g325_n_spl_;
  wire g325_p_spl_;
  wire g326_n_spl_;
  wire g328_p_spl_;
  wire g326_p_spl_;
  wire g328_n_spl_;
  wire g329_n_spl_;
  wire g329_p_spl_;
  wire g332_n_spl_;
  wire g334_p_spl_;
  wire g332_p_spl_;
  wire g334_n_spl_;
  wire g335_n_spl_;
  wire g335_n_spl_0;
  wire g335_p_spl_;
  wire g335_p_spl_0;
  wire g331_p_spl_;
  wire g337_p_spl_;
  wire g331_n_spl_;
  wire g337_n_spl_;
  wire g338_n_spl_;
  wire g338_p_spl_;
  wire g339_n_spl_;
  wire g341_p_spl_;
  wire g339_p_spl_;
  wire g341_n_spl_;
  wire g342_n_spl_;
  wire g342_p_spl_;
  wire g344_p_spl_;
  wire g344_n_spl_;
  wire g345_n_spl_;
  wire g345_p_spl_;
  wire g346_n_spl_;
  wire g348_p_spl_;
  wire g346_p_spl_;
  wire g348_n_spl_;
  wire g350_p_spl_;
  wire g351_p_spl_;
  wire g351_p_spl_0;
  wire g350_n_spl_;
  wire g351_n_spl_;
  wire g351_n_spl_0;
  wire g352_n_spl_;
  wire g352_p_spl_;
  wire g353_p_spl_;
  wire g355_p_spl_;
  wire g353_n_spl_;
  wire g355_n_spl_;
  wire g356_n_spl_;
  wire g356_p_spl_;
  wire g357_n_spl_;
  wire g359_p_spl_;
  wire g357_p_spl_;
  wire g359_n_spl_;
  wire g362_p_spl_;
  wire g362_p_spl_0;
  wire g362_n_spl_;
  wire g362_n_spl_0;
  wire g363_n_spl_;
  wire g363_p_spl_;
  wire g361_p_spl_;
  wire g365_p_spl_;
  wire g361_n_spl_;
  wire g365_n_spl_;
  wire g366_n_spl_;
  wire g366_p_spl_;
  wire g360_n_spl_;
  wire g360_p_spl_;
  wire g368_p_spl_;
  wire g370_p_spl_;
  wire g368_n_spl_;
  wire g370_n_spl_;
  wire g371_n_spl_;
  wire g371_p_spl_;
  wire g372_n_spl_;
  wire g374_p_spl_;
  wire g372_p_spl_;
  wire g374_n_spl_;
  wire g376_n_spl_;
  wire g377_p_spl_;
  wire g376_p_spl_;
  wire g377_n_spl_;
  wire g378_n_spl_;
  wire g378_n_spl_0;
  wire g378_p_spl_;
  wire g378_p_spl_0;
  wire g375_n_spl_;
  wire g375_p_spl_;
  wire g380_p_spl_;
  wire g382_p_spl_;
  wire g380_n_spl_;
  wire g382_n_spl_;
  wire g383_n_spl_;
  wire g383_p_spl_;
  wire g384_n_spl_;
  wire g386_p_spl_;
  wire g384_p_spl_;
  wire g386_n_spl_;
  wire g387_n_spl_;
  wire g387_p_spl_;
  wire g389_p_spl_;
  wire g389_n_spl_;
  wire g390_n_spl_;
  wire g390_p_spl_;
  wire g391_n_spl_;
  wire g393_p_spl_;
  wire g391_p_spl_;
  wire g393_n_spl_;
  wire g395_p_spl_;
  wire g395_p_spl_0;
  wire g395_n_spl_;
  wire g395_n_spl_0;
  wire g396_n_spl_;
  wire g396_p_spl_;
  wire g397_p_spl_;
  wire g401_p_spl_;
  wire g397_n_spl_;
  wire g401_n_spl_;
  wire g402_n_spl_;
  wire g402_p_spl_;
  wire g403_n_spl_;
  wire g405_p_spl_;
  wire g403_p_spl_;
  wire g405_n_spl_;
  wire g407_p_spl_;
  wire g407_p_spl_0;
  wire g407_n_spl_;
  wire g407_n_spl_0;
  wire g408_n_spl_;
  wire g408_n_spl_0;
  wire g408_p_spl_;
  wire g408_p_spl_0;
  wire g406_n_spl_;
  wire g406_p_spl_;
  wire g412_p_spl_;
  wire g414_p_spl_;
  wire g412_n_spl_;
  wire g414_n_spl_;
  wire g415_n_spl_;
  wire g415_p_spl_;
  wire g416_n_spl_;
  wire g418_p_spl_;
  wire g416_p_spl_;
  wire g418_n_spl_;
  wire g419_n_spl_;
  wire g419_p_spl_;
  wire g421_p_spl_;
  wire g421_n_spl_;
  wire g422_n_spl_;
  wire g422_p_spl_;
  wire g423_n_spl_;
  wire g425_p_spl_;
  wire g423_p_spl_;
  wire g425_n_spl_;
  wire g426_p_spl_;
  wire g426_p_spl_0;
  wire g428_p_spl_;
  wire g426_n_spl_;
  wire g426_n_spl_0;
  wire g428_n_spl_;
  wire g430_p_spl_;
  wire g430_p_spl_0;
  wire g430_n_spl_;
  wire g430_n_spl_0;
  wire g431_n_spl_;
  wire g431_p_spl_;
  wire g432_p_spl_;
  wire g434_p_spl_;
  wire g432_n_spl_;
  wire g434_n_spl_;
  wire g435_n_spl_;
  wire g435_p_spl_;
  wire g436_n_spl_;
  wire g438_p_spl_;
  wire g436_p_spl_;
  wire g438_n_spl_;
  wire g439_n_spl_;
  wire g439_p_spl_;
  wire g441_p_spl_;
  wire g441_n_spl_;
  wire g442_n_spl_;
  wire g442_p_spl_;
  wire g443_n_spl_;
  wire g445_p_spl_;
  wire g443_p_spl_;
  wire g445_n_spl_;
  wire g446_p_spl_;
  wire g446_p_spl_0;
  wire g448_p_spl_;
  wire g446_n_spl_;
  wire g446_n_spl_0;
  wire g448_n_spl_;
  wire g449_p_spl_;
  wire g449_p_spl_0;
  wire g451_p_spl_;
  wire g449_n_spl_;
  wire g449_n_spl_0;
  wire g451_n_spl_;
  wire g453_p_spl_;
  wire g453_n_spl_;
  wire g454_p_spl_;
  wire g454_p_spl_0;
  wire g456_p_spl_;
  wire g454_n_spl_;
  wire g454_n_spl_0;
  wire g456_n_spl_;
  wire g457_p_spl_;
  wire g457_p_spl_0;
  wire g459_p_spl_;
  wire g457_n_spl_;
  wire g457_n_spl_0;
  wire g459_n_spl_;
  wire g460_p_spl_;
  wire g460_p_spl_0;
  wire g462_p_spl_;
  wire g460_n_spl_;
  wire g460_n_spl_0;
  wire g462_n_spl_;
  wire g463_p_spl_;
  wire g463_p_spl_0;
  wire g465_p_spl_;
  wire g463_n_spl_;
  wire g463_n_spl_0;
  wire g465_n_spl_;
  wire g452_n_spl_;
  wire g452_p_spl_;
  wire g466_p_spl_;
  wire g466_p_spl_0;
  wire g468_p_spl_;
  wire g466_n_spl_;
  wire g466_n_spl_0;
  wire g468_n_spl_;
  wire g469_n_spl_;
  wire g469_p_spl_;
  wire g429_n_spl_;
  wire g429_p_spl_;
  wire g470_n_spl_;
  wire g472_p_spl_;
  wire g470_p_spl_;
  wire g472_n_spl_;
  wire g473_n_spl_;
  wire g473_p_spl_;
  wire g394_n_spl_;
  wire g394_p_spl_;
  wire g474_n_spl_;
  wire g476_p_spl_;
  wire g474_p_spl_;
  wire g476_n_spl_;
  wire g477_n_spl_;
  wire g477_p_spl_;
  wire g349_n_spl_;
  wire g349_p_spl_;
  wire g478_n_spl_;
  wire g480_p_spl_;
  wire g478_p_spl_;
  wire g480_n_spl_;
  wire g481_n_spl_;
  wire g481_p_spl_;
  wire g303_p_spl_;
  wire g482_n_spl_;
  wire g303_n_spl_;
  wire g482_p_spl_;
  wire g483_n_spl_;
  wire g483_p_spl_;
  wire g240_p_spl_;
  wire g484_n_spl_;
  wire g240_n_spl_;
  wire g484_p_spl_;
  wire g485_n_spl_;
  wire g485_p_spl_;
  wire g185_n_spl_;
  wire g185_p_spl_;
  wire g486_n_spl_;
  wire g488_p_spl_;
  wire g486_p_spl_;
  wire g488_n_spl_;
  wire g489_n_spl_;
  wire g489_p_spl_;
  wire g137_n_spl_;
  wire g137_p_spl_;
  wire g490_n_spl_;
  wire g492_p_spl_;
  wire g490_p_spl_;
  wire g492_n_spl_;
  wire g493_n_spl_;
  wire g493_p_spl_;
  wire g498_p_spl_;
  wire g498_n_spl_;
  wire g499_n_spl_;
  wire g499_n_spl_0;
  wire g499_p_spl_;
  wire g499_p_spl_0;
  wire g501_n_spl_;
  wire g501_p_spl_;
  wire g502_n_spl_;
  wire g502_p_spl_;
  wire g504_n_spl_;
  wire g505_n_spl_;
  wire g504_p_spl_;
  wire g505_p_spl_;
  wire g506_n_spl_;
  wire g506_p_spl_;
  wire g496_n_spl_;
  wire g508_p_spl_;
  wire g496_p_spl_;
  wire g508_n_spl_;
  wire g509_n_spl_;
  wire g509_p_spl_;
  wire g495_n_spl_;
  wire g511_p_spl_;
  wire g495_p_spl_;
  wire g511_n_spl_;
  wire g512_n_spl_;
  wire g512_p_spl_;
  wire g494_n_spl_;
  wire g514_p_spl_;
  wire g494_p_spl_;
  wire g514_n_spl_;
  wire g516_p_spl_;
  wire g516_n_spl_;
  wire g515_n_spl_;
  wire g515_p_spl_;
  wire g533_n_spl_;
  wire g535_n_spl_;
  wire g533_p_spl_;
  wire g535_p_spl_;
  wire g531_n_spl_;
  wire g531_p_spl_;
  wire g529_n_spl_;
  wire g529_p_spl_;
  wire g540_n_spl_;
  wire g542_n_spl_;
  wire g540_p_spl_;
  wire g542_p_spl_;
  wire g525_n_spl_;
  wire g525_p_spl_;
  wire g523_n_spl_;
  wire g523_n_spl_0;
  wire g523_n_spl_1;
  wire g523_p_spl_;
  wire g523_p_spl_0;
  wire g523_p_spl_1;
  wire g554_n_spl_;
  wire g554_n_spl_0;
  wire g554_n_spl_00;
  wire g554_n_spl_01;
  wire g554_n_spl_1;
  wire g554_n_spl_10;
  wire g554_p_spl_;
  wire g554_p_spl_0;
  wire g554_p_spl_00;
  wire g554_p_spl_01;
  wire g554_p_spl_1;
  wire g554_p_spl_10;
  wire g547_n_spl_;
  wire g547_n_spl_0;
  wire g547_n_spl_00;
  wire g547_n_spl_01;
  wire g547_n_spl_1;
  wire g547_n_spl_10;
  wire g547_p_spl_;
  wire g547_p_spl_0;
  wire g547_p_spl_00;
  wire g547_p_spl_01;
  wire g547_p_spl_1;
  wire g547_p_spl_10;
  wire g558_n_spl_;
  wire g559_p_spl_;
  wire g558_p_spl_;
  wire g559_n_spl_;
  wire g559_n_spl_0;
  wire g564_n_spl_;
  wire g565_p_spl_;
  wire g564_p_spl_;
  wire g565_n_spl_;
  wire g565_n_spl_0;
  wire g570_n_spl_;
  wire g571_p_spl_;
  wire g570_p_spl_;
  wire g571_n_spl_;
  wire g571_n_spl_0;
  wire g572_n_spl_;
  wire g572_p_spl_;
  wire g578_n_spl_;
  wire g579_p_spl_;
  wire g578_p_spl_;
  wire g579_n_spl_;
  wire g579_n_spl_0;
  wire g585_n_spl_;
  wire g586_p_spl_;
  wire g585_p_spl_;
  wire g586_n_spl_;
  wire g586_n_spl_0;
  wire g589_p_spl_;
  wire g595_n_spl_;
  wire g589_n_spl_;
  wire g589_n_spl_0;
  wire g595_p_spl_;
  wire g598_n_spl_;
  wire g598_n_spl_0;
  wire g600_n_spl_;
  wire g597_n_spl_;
  wire g601_p_spl_;
  wire g601_p_spl_0;
  wire g597_p_spl_;
  wire g601_n_spl_;
  wire g596_n_spl_;
  wire g596_p_spl_;
  wire g588_n_spl_;
  wire g603_n_spl_;
  wire g588_p_spl_;
  wire g603_p_spl_;
  wire g587_n_spl_;
  wire g587_p_spl_;
  wire g581_n_spl_;
  wire g605_n_spl_;
  wire g581_p_spl_;
  wire g605_p_spl_;
  wire g580_n_spl_;
  wire g580_p_spl_;
  wire g574_n_spl_;
  wire g607_p_spl_;
  wire g608_p_spl_;
  wire g566_n_spl_;
  wire g566_p_spl_;
  wire g609_p_spl_;
  wire g611_n_spl_;
  wire g612_p_spl_;
  wire g560_n_spl_;
  wire g560_p_spl_;
  wire g613_p_spl_;
  wire g615_n_spl_;
  wire g616_p_spl_;
  wire g27_n_spl_;
  wire g617_p_spl_;
  wire g617_p_spl_0;
  wire g618_n_spl_;
  wire g618_p_spl_;
  wire g621_p_spl_;
  wire g622_p_spl_;
  wire g617_n_spl_;
  wire g622_n_spl_;
  wire g620_p_spl_;
  wire g620_p_spl_0;
  wire g620_p_spl_00;
  wire g620_p_spl_01;
  wire g620_p_spl_1;
  wire g620_p_spl_10;
  wire g620_p_spl_11;
  wire g626_n_spl_;
  wire g630_p_spl_;
  wire g630_p_spl_0;
  wire g630_p_spl_00;
  wire g630_p_spl_01;
  wire g630_p_spl_1;
  wire g630_p_spl_10;
  wire g628_n_spl_;
  wire g628_n_spl_0;
  wire g628_n_spl_00;
  wire g628_n_spl_01;
  wire g628_n_spl_1;
  wire g628_n_spl_10;
  wire g628_n_spl_11;
  wire g636_n_spl_;
  wire g645_n_spl_;
  wire g654_n_spl_;
  wire g663_n_spl_;
  wire g670_n_spl_;
  wire g677_n_spl_;
  wire g684_n_spl_;

  buf

  (
    enable_p,
    enable
  );


  not

  (
    enable_n,
    enable
  );


  buf

  (
    reset_p,
    reset
  );


  not

  (
    reset_n,
    reset
  );


  buf

  (
    input_f[0]_p,
    input_f[0]
  );


  not

  (
    input_f[0]_n,
    input_f[0]
  );


  buf

  (
    input_f[1]_p,
    input_f[1]
  );


  not

  (
    input_f[1]_n,
    input_f[1]
  );


  buf

  (
    input_f[2]_p,
    input_f[2]
  );


  not

  (
    input_f[2]_n,
    input_f[2]
  );


  buf

  (
    input_f[3]_p,
    input_f[3]
  );


  not

  (
    input_f[3]_n,
    input_f[3]
  );


  buf

  (
    input_f[4]_p,
    input_f[4]
  );


  not

  (
    input_f[4]_n,
    input_f[4]
  );


  buf

  (
    input_f[5]_p,
    input_f[5]
  );


  not

  (
    input_f[5]_n,
    input_f[5]
  );


  buf

  (
    input_f[6]_p,
    input_f[6]
  );


  not

  (
    input_f[6]_n,
    input_f[6]
  );


  buf

  (
    input_f[7]_p,
    input_f[7]
  );


  not

  (
    input_f[7]_n,
    input_f[7]
  );


  buf

  (
    input_w[0]_p,
    input_w[0]
  );


  not

  (
    input_w[0]_n,
    input_w[0]
  );


  buf

  (
    input_w[1]_p,
    input_w[1]
  );


  not

  (
    input_w[1]_n,
    input_w[1]
  );


  buf

  (
    input_w[2]_p,
    input_w[2]
  );


  not

  (
    input_w[2]_n,
    input_w[2]
  );


  buf

  (
    input_w[3]_p,
    input_w[3]
  );


  not

  (
    input_w[3]_n,
    input_w[3]
  );


  buf

  (
    input_w[4]_p,
    input_w[4]
  );


  not

  (
    input_w[4]_n,
    input_w[4]
  );


  buf

  (
    input_w[5]_p,
    input_w[5]
  );


  not

  (
    input_w[5]_n,
    input_w[5]
  );


  buf

  (
    input_w[6]_p,
    input_w[6]
  );


  not

  (
    input_w[6]_n,
    input_w[6]
  );


  buf

  (
    input_w[7]_p,
    input_w[7]
  );


  not

  (
    input_w[7]_n,
    input_w[7]
  );


  buf

  (
    psum_reg[0]_p,
    psum_reg[0]
  );


  not

  (
    psum_reg[0]_n,
    psum_reg[0]
  );


  buf

  (
    psum_reg[1]_p,
    psum_reg[1]
  );


  not

  (
    psum_reg[1]_n,
    psum_reg[1]
  );


  buf

  (
    psum_reg[2]_p,
    psum_reg[2]
  );


  not

  (
    psum_reg[2]_n,
    psum_reg[2]
  );


  buf

  (
    psum_reg[3]_p,
    psum_reg[3]
  );


  not

  (
    psum_reg[3]_n,
    psum_reg[3]
  );


  buf

  (
    psum_reg[4]_p,
    psum_reg[4]
  );


  not

  (
    psum_reg[4]_n,
    psum_reg[4]
  );


  buf

  (
    psum_reg[5]_p,
    psum_reg[5]
  );


  not

  (
    psum_reg[5]_n,
    psum_reg[5]
  );


  buf

  (
    psum_reg[6]_p,
    psum_reg[6]
  );


  not

  (
    psum_reg[6]_n,
    psum_reg[6]
  );


  buf

  (
    psum_reg[7]_p,
    psum_reg[7]
  );


  not

  (
    psum_reg[7]_n,
    psum_reg[7]
  );


  and

  (
    g27_p,
    reset_n_spl_00,
    psum_reg[7]_p
  );


  or

  (
    g27_n,
    reset_p_spl_00,
    psum_reg[7]_n
  );


  and

  (
    g28_p,
    enable_n_spl_00,
    g27_p_spl_0
  );


  and

  (
    g29_p,
    input_f[7]_p_spl_00,
    input_w[0]_p_spl_000
  );


  or

  (
    g29_n,
    input_f[7]_n_spl_00,
    input_w[0]_n_spl_000
  );


  and

  (
    g30_p,
    input_w[1]_p_spl_000,
    g29_p_spl_0
  );


  or

  (
    g30_n,
    input_w[1]_n_spl_000,
    g29_n_spl_0
  );


  and

  (
    g31_p,
    input_w[2]_p_spl_000,
    g30_p_spl_0
  );


  or

  (
    g31_n,
    input_w[2]_n_spl_000,
    g30_n_spl_0
  );


  and

  (
    g32_p,
    input_f[7]_p_spl_00,
    input_w[2]_p_spl_000
  );


  or

  (
    g32_n,
    input_f[7]_n_spl_00,
    input_w[2]_n_spl_000
  );


  and

  (
    g33_p,
    input_w[0]_n_spl_000,
    input_w[1]_n_spl_000
  );


  or

  (
    g33_n,
    input_w[0]_p_spl_000,
    input_w[1]_p_spl_000
  );


  and

  (
    g34_p,
    input_f[7]_p_spl_01,
    g33_n
  );


  or

  (
    g34_n,
    input_f[7]_n_spl_01,
    g33_p
  );


  and

  (
    g35_p,
    g32_n_spl_,
    g34_n_spl_0
  );


  or

  (
    g35_n,
    g32_p_spl_,
    g34_p_spl_0
  );


  and

  (
    g36_p,
    g31_n_spl_00,
    g35_n_spl_0
  );


  or

  (
    g36_n,
    g31_p_spl_00,
    g35_p_spl_0
  );


  and

  (
    g37_p,
    input_f[5]_p_spl_00,
    input_w[5]_p_spl_00
  );


  or

  (
    g37_n,
    input_f[5]_n_spl_00,
    input_w[5]_n_spl_00
  );


  and

  (
    g38_p,
    input_f[7]_p_spl_01,
    input_w[3]_p_spl_000
  );


  or

  (
    g38_n,
    input_f[7]_n_spl_01,
    input_w[3]_n_spl_000
  );


  and

  (
    g39_p,
    input_f[6]_p_spl_00,
    input_w[4]_p_spl_000
  );


  or

  (
    g39_n,
    input_f[6]_n_spl_00,
    input_w[4]_n_spl_000
  );


  and

  (
    g40_p,
    g38_p_spl_0,
    g39_p_spl_0
  );


  or

  (
    g40_n,
    g38_n_spl_0,
    g39_n_spl_0
  );


  and

  (
    g41_p,
    g38_n_spl_0,
    g39_n_spl_0
  );


  or

  (
    g41_n,
    g38_p_spl_0,
    g39_p_spl_0
  );


  and

  (
    g42_p,
    g40_n_spl_,
    g41_n
  );


  or

  (
    g42_n,
    g40_p_spl_,
    g41_p
  );


  and

  (
    g43_p,
    g37_p_spl_,
    g42_p_spl_
  );


  or

  (
    g43_n,
    g37_n_spl_,
    g42_n_spl_
  );


  and

  (
    g44_p,
    g37_n_spl_,
    g42_n_spl_
  );


  or

  (
    g44_n,
    g37_p_spl_,
    g42_p_spl_
  );


  and

  (
    g45_p,
    g43_n_spl_,
    g44_n
  );


  or

  (
    g45_n,
    g43_p_spl_,
    g44_p
  );


  and

  (
    g46_p,
    g36_p_spl_00,
    g45_p_spl_
  );


  or

  (
    g46_n,
    g36_n_spl_00,
    g45_n_spl_
  );


  and

  (
    g47_p,
    g31_n_spl_00,
    g46_n_spl_
  );


  or

  (
    g47_n,
    g31_p_spl_00,
    g46_p_spl_
  );


  and

  (
    g48_p,
    input_w[3]_n_spl_000,
    input_w[4]_n_spl_000
  );


  or

  (
    g48_n,
    input_w[3]_p_spl_000,
    input_w[4]_p_spl_000
  );


  and

  (
    g49_p,
    input_w[4]_p_spl_00,
    g38_p_spl_
  );


  or

  (
    g49_n,
    input_w[4]_n_spl_00,
    g38_n_spl_
  );


  and

  (
    g50_p,
    input_f[7]_p_spl_10,
    g49_n_spl_0
  );


  or

  (
    g50_n,
    input_f[7]_n_spl_10,
    g49_p_spl_0
  );


  and

  (
    g51_p,
    g48_n,
    g50_p
  );


  or

  (
    g51_n,
    g48_p,
    g50_n
  );


  and

  (
    g52_p,
    input_f[6]_p_spl_00,
    input_w[5]_p_spl_00
  );


  or

  (
    g52_n,
    input_f[6]_n_spl_00,
    input_w[5]_n_spl_00
  );


  and

  (
    g53_p,
    g51_p_spl_0,
    g52_p_spl_
  );


  or

  (
    g53_n,
    g51_n_spl_0,
    g52_n_spl_
  );


  and

  (
    g54_p,
    g51_n_spl_0,
    g52_n_spl_
  );


  or

  (
    g54_n,
    g51_p_spl_0,
    g52_p_spl_
  );


  and

  (
    g55_p,
    g53_n_spl_,
    g54_n
  );


  or

  (
    g55_n,
    g53_p_spl_,
    g54_p
  );


  and

  (
    g56_p,
    g36_p_spl_00,
    g55_p_spl_
  );


  or

  (
    g56_n,
    g36_n_spl_00,
    g55_n_spl_
  );


  and

  (
    g57_p,
    g36_n_spl_01,
    g55_n_spl_
  );


  or

  (
    g57_n,
    g36_p_spl_01,
    g55_p_spl_
  );


  and

  (
    g58_p,
    g56_n_spl_,
    g57_n
  );


  or

  (
    g58_n,
    g56_p_spl_,
    g57_p
  );


  and

  (
    g59_p,
    g47_n_spl_,
    g58_p_spl_
  );


  or

  (
    g59_n,
    g47_p_spl_,
    g58_n_spl_
  );


  and

  (
    g60_p,
    input_f[4]_p_spl_00,
    input_w[6]_p_spl_00
  );


  or

  (
    g60_n,
    input_f[4]_n_spl_00,
    input_w[6]_n_spl_00
  );


  and

  (
    g61_p,
    input_f[3]_n_spl_00,
    input_w[7]_p_spl_000
  );


  or

  (
    g61_n,
    input_f[3]_p_spl_00,
    input_w[7]_n_spl_000
  );


  and

  (
    g62_p,
    g60_p_spl_,
    g61_p_spl_
  );


  or

  (
    g62_n,
    g60_n_spl_,
    g61_n_spl_
  );


  and

  (
    g63_p,
    g40_n_spl_,
    g43_n_spl_
  );


  or

  (
    g63_n,
    g40_p_spl_,
    g43_p_spl_
  );


  and

  (
    g64_p,
    input_f[5]_p_spl_00,
    input_w[6]_p_spl_00
  );


  or

  (
    g64_n,
    input_f[5]_n_spl_00,
    input_w[6]_n_spl_00
  );


  and

  (
    g65_p,
    input_f[4]_n_spl_00,
    input_w[7]_p_spl_000
  );


  or

  (
    g65_n,
    input_f[4]_p_spl_00,
    input_w[7]_n_spl_000
  );


  and

  (
    g66_p,
    g64_p_spl_,
    g65_p_spl_
  );


  or

  (
    g66_n,
    g64_n_spl_,
    g65_n_spl_
  );


  and

  (
    g67_p,
    g64_n_spl_,
    g65_n_spl_
  );


  or

  (
    g67_n,
    g64_p_spl_,
    g65_p_spl_
  );


  and

  (
    g68_p,
    g66_n_spl_0,
    g67_n
  );


  or

  (
    g68_n,
    g66_p_spl_0,
    g67_p
  );


  and

  (
    g69_p,
    g63_n_spl_,
    g68_p_spl_
  );


  or

  (
    g69_n,
    g63_p_spl_,
    g68_n_spl_
  );


  and

  (
    g70_p,
    g63_p_spl_,
    g68_n_spl_
  );


  or

  (
    g70_n,
    g63_n_spl_,
    g68_p_spl_
  );


  and

  (
    g71_p,
    g69_n_spl_,
    g70_n
  );


  or

  (
    g71_n,
    g69_p_spl_,
    g70_p
  );


  and

  (
    g72_p,
    g62_p_spl_0,
    g71_p_spl_
  );


  or

  (
    g72_n,
    g62_n_spl_0,
    g71_n_spl_
  );


  and

  (
    g73_p,
    g62_n_spl_0,
    g71_n_spl_
  );


  or

  (
    g73_n,
    g62_p_spl_0,
    g71_p_spl_
  );


  and

  (
    g74_p,
    g72_n_spl_,
    g73_n
  );


  or

  (
    g74_n,
    g72_p_spl_,
    g73_p
  );


  and

  (
    g75_p,
    g47_p_spl_,
    g58_n_spl_
  );


  or

  (
    g75_n,
    g47_n_spl_,
    g58_p_spl_
  );


  and

  (
    g76_p,
    g59_n_spl_,
    g75_n
  );


  or

  (
    g76_n,
    g59_p_spl_,
    g75_p
  );


  and

  (
    g77_p,
    g74_p_spl_,
    g76_p_spl_
  );


  or

  (
    g77_n,
    g74_n_spl_,
    g76_n_spl_
  );


  and

  (
    g78_p,
    g59_n_spl_,
    g77_n_spl_
  );


  or

  (
    g78_n,
    g59_p_spl_,
    g77_p_spl_
  );


  and

  (
    g79_p,
    g49_n_spl_0,
    g53_n_spl_
  );


  or

  (
    g79_n,
    g49_p_spl_0,
    g53_p_spl_
  );


  and

  (
    g80_p,
    input_f[6]_p_spl_01,
    input_w[6]_p_spl_01
  );


  or

  (
    g80_n,
    input_f[6]_n_spl_01,
    input_w[6]_n_spl_01
  );


  and

  (
    g81_p,
    input_f[5]_n_spl_01,
    input_w[7]_p_spl_001
  );


  or

  (
    g81_n,
    input_f[5]_p_spl_01,
    input_w[7]_n_spl_001
  );


  and

  (
    g82_p,
    g80_p_spl_,
    g81_p_spl_
  );


  or

  (
    g82_n,
    g80_n_spl_,
    g81_n_spl_
  );


  and

  (
    g83_p,
    g80_n_spl_,
    g81_n_spl_
  );


  or

  (
    g83_n,
    g80_p_spl_,
    g81_p_spl_
  );


  and

  (
    g84_p,
    g82_n_spl_0,
    g83_n
  );


  or

  (
    g84_n,
    g82_p_spl_0,
    g83_p
  );


  and

  (
    g85_p,
    g79_n_spl_,
    g84_p_spl_
  );


  or

  (
    g85_n,
    g79_p_spl_,
    g84_n_spl_
  );


  and

  (
    g86_p,
    g79_p_spl_,
    g84_n_spl_
  );


  or

  (
    g86_n,
    g79_n_spl_,
    g84_p_spl_
  );


  and

  (
    g87_p,
    g85_n_spl_,
    g86_n
  );


  or

  (
    g87_n,
    g85_p_spl_,
    g86_p
  );


  and

  (
    g88_p,
    g66_p_spl_0,
    g87_p_spl_
  );


  or

  (
    g88_n,
    g66_n_spl_0,
    g87_n_spl_
  );


  and

  (
    g89_p,
    g66_n_spl_,
    g87_n_spl_
  );


  or

  (
    g89_n,
    g66_p_spl_,
    g87_p_spl_
  );


  and

  (
    g90_p,
    g88_n_spl_,
    g89_n
  );


  or

  (
    g90_n,
    g88_p_spl_,
    g89_p
  );


  and

  (
    g91_p,
    g31_n_spl_01,
    g56_n_spl_
  );


  or

  (
    g91_n,
    g31_p_spl_01,
    g56_p_spl_
  );


  and

  (
    g92_p,
    input_f[7]_p_spl_10,
    input_w[5]_p_spl_01
  );


  or

  (
    g92_n,
    input_f[7]_n_spl_10,
    input_w[5]_n_spl_01
  );


  and

  (
    g93_p,
    g51_p_spl_1,
    g92_p_spl_
  );


  or

  (
    g93_n,
    g51_n_spl_1,
    g92_n_spl_
  );


  and

  (
    g94_p,
    g51_n_spl_1,
    g92_n_spl_
  );


  or

  (
    g94_n,
    g51_p_spl_1,
    g92_p_spl_
  );


  and

  (
    g95_p,
    g93_n_spl_,
    g94_n
  );


  or

  (
    g95_n,
    g93_p_spl_,
    g94_p
  );


  and

  (
    g96_p,
    g36_n_spl_01,
    g95_p_spl_0
  );


  or

  (
    g96_n,
    g36_p_spl_01,
    g95_n_spl_0
  );


  and

  (
    g97_p,
    g36_p_spl_1,
    g95_n_spl_0
  );


  or

  (
    g97_n,
    g36_n_spl_1,
    g95_p_spl_0
  );


  and

  (
    g98_p,
    g96_n,
    g97_n
  );


  or

  (
    g98_n,
    g96_p,
    g97_p
  );


  and

  (
    g99_p,
    g91_n_spl_,
    g98_n_spl_
  );


  or

  (
    g99_n,
    g91_p_spl_,
    g98_p_spl_
  );


  and

  (
    g100_p,
    g91_p_spl_,
    g98_p_spl_
  );


  or

  (
    g100_n,
    g91_n_spl_,
    g98_n_spl_
  );


  and

  (
    g101_p,
    g99_n_spl_,
    g100_n
  );


  or

  (
    g101_n,
    g99_p_spl_,
    g100_p
  );


  and

  (
    g102_p,
    g90_p_spl_,
    g101_p_spl_
  );


  or

  (
    g102_n,
    g90_n_spl_,
    g101_n_spl_
  );


  and

  (
    g103_p,
    g90_n_spl_,
    g101_n_spl_
  );


  or

  (
    g103_n,
    g90_p_spl_,
    g101_p_spl_
  );


  and

  (
    g104_p,
    g102_n_spl_,
    g103_n
  );


  or

  (
    g104_n,
    g102_p_spl_,
    g103_p
  );


  and

  (
    g105_p,
    g78_n_spl_,
    g104_p_spl_
  );


  or

  (
    g105_n,
    g78_p_spl_,
    g104_n_spl_
  );


  and

  (
    g106_p,
    g69_n_spl_,
    g72_n_spl_
  );


  or

  (
    g106_n,
    g69_p_spl_,
    g72_p_spl_
  );


  and

  (
    g107_p,
    g78_p_spl_,
    g104_n_spl_
  );


  or

  (
    g107_n,
    g78_n_spl_,
    g104_p_spl_
  );


  and

  (
    g108_p,
    g105_n_spl_,
    g107_n
  );


  or

  (
    g108_n,
    g105_p_spl_,
    g107_p
  );


  and

  (
    g109_p,
    g106_n_spl_,
    g108_p_spl_
  );


  or

  (
    g109_n,
    g106_p_spl_,
    g108_n_spl_
  );


  and

  (
    g110_p,
    g105_n_spl_,
    g109_n_spl_
  );


  or

  (
    g110_n,
    g105_p_spl_,
    g109_p_spl_
  );


  and

  (
    g111_p,
    g85_n_spl_,
    g88_n_spl_
  );


  or

  (
    g111_n,
    g85_p_spl_,
    g88_p_spl_
  );


  and

  (
    g112_p,
    g99_n_spl_,
    g102_n_spl_
  );


  or

  (
    g112_n,
    g99_p_spl_,
    g102_p_spl_
  );


  and

  (
    g113_p,
    g31_p_spl_01,
    g95_p_spl_1
  );


  or

  (
    g113_n,
    g31_n_spl_01,
    g95_n_spl_1
  );


  and

  (
    g114_p,
    g35_p_spl_0,
    g95_n_spl_1
  );


  or

  (
    g114_n,
    g35_n_spl_0,
    g95_p_spl_1
  );


  and

  (
    g115_p,
    g113_n_spl_0,
    g114_n
  );


  or

  (
    g115_n,
    g113_p_spl_0,
    g114_p
  );


  and

  (
    g116_p,
    g49_n_spl_,
    g93_n_spl_
  );


  or

  (
    g116_n,
    g49_p_spl_,
    g93_p_spl_
  );


  and

  (
    g117_p,
    input_f[7]_p_spl_11,
    input_w[6]_p_spl_01
  );


  or

  (
    g117_n,
    input_f[7]_n_spl_11,
    input_w[6]_n_spl_01
  );


  and

  (
    g118_p,
    input_f[6]_n_spl_01,
    input_w[7]_p_spl_001
  );


  or

  (
    g118_n,
    input_f[6]_p_spl_01,
    input_w[7]_n_spl_001
  );


  and

  (
    g119_p,
    g117_p_spl_,
    g118_n_spl_
  );


  or

  (
    g119_n,
    g117_n_spl_,
    g118_p_spl_
  );


  and

  (
    g120_p,
    g117_n_spl_,
    g118_p_spl_
  );


  or

  (
    g120_n,
    g117_p_spl_,
    g118_n_spl_
  );


  and

  (
    g121_p,
    g119_n_spl_,
    g120_n
  );


  or

  (
    g121_n,
    g119_p_spl_,
    g120_p
  );


  and

  (
    g122_p,
    g116_n_spl_0,
    g121_n_spl_
  );


  or

  (
    g122_n,
    g116_p_spl_0,
    g121_p_spl_
  );


  and

  (
    g123_p,
    g116_p_spl_0,
    g121_p_spl_
  );


  or

  (
    g123_n,
    g116_n_spl_0,
    g121_n_spl_
  );


  and

  (
    g124_p,
    g122_n_spl_,
    g123_n
  );


  or

  (
    g124_n,
    g122_p_spl_,
    g123_p
  );


  and

  (
    g125_p,
    g82_p_spl_0,
    g124_p_spl_
  );


  or

  (
    g125_n,
    g82_n_spl_0,
    g124_n_spl_
  );


  and

  (
    g126_p,
    g82_n_spl_,
    g124_n_spl_
  );


  or

  (
    g126_n,
    g82_p_spl_,
    g124_p_spl_
  );


  and

  (
    g127_p,
    g125_n_spl_,
    g126_n
  );


  or

  (
    g127_n,
    g125_p_spl_,
    g126_p
  );


  and

  (
    g128_p,
    g115_p_spl_0,
    g127_p_spl_
  );


  or

  (
    g128_n,
    g115_n_spl_0,
    g127_n_spl_
  );


  and

  (
    g129_p,
    g115_n_spl_0,
    g127_n_spl_
  );


  or

  (
    g129_n,
    g115_p_spl_0,
    g127_p_spl_
  );


  and

  (
    g130_p,
    g128_n_spl_,
    g129_n
  );


  or

  (
    g130_n,
    g128_p_spl_,
    g129_p
  );


  and

  (
    g131_p,
    g112_n_spl_,
    g130_p_spl_
  );


  or

  (
    g131_n,
    g112_p_spl_,
    g130_n_spl_
  );


  and

  (
    g132_p,
    g112_p_spl_,
    g130_n_spl_
  );


  or

  (
    g132_n,
    g112_n_spl_,
    g130_p_spl_
  );


  and

  (
    g133_p,
    g131_n_spl_,
    g132_n
  );


  or

  (
    g133_n,
    g131_p_spl_,
    g132_p
  );


  and

  (
    g134_p,
    g111_n_spl_,
    g133_p_spl_
  );


  or

  (
    g134_n,
    g111_p_spl_,
    g133_n_spl_
  );


  and

  (
    g135_p,
    g111_p_spl_,
    g133_n_spl_
  );


  or

  (
    g135_n,
    g111_n_spl_,
    g133_p_spl_
  );


  and

  (
    g136_p,
    g134_n_spl_,
    g135_n
  );


  or

  (
    g136_n,
    g134_p_spl_,
    g135_p
  );


  and

  (
    g137_p,
    g110_n_spl_,
    g136_p_spl_
  );


  or

  (
    g137_n,
    g110_p_spl_,
    g136_n_spl_
  );


  and

  (
    g138_p,
    input_f[4]_p_spl_01,
    input_w[5]_p_spl_01
  );


  or

  (
    g138_n,
    input_f[4]_n_spl_01,
    input_w[5]_n_spl_01
  );


  and

  (
    g139_p,
    input_f[5]_p_spl_01,
    input_w[3]_p_spl_00
  );


  or

  (
    g139_n,
    input_f[5]_n_spl_01,
    input_w[3]_n_spl_00
  );


  and

  (
    g140_p,
    g39_p_spl_,
    g139_p_spl_0
  );


  or

  (
    g140_n,
    g39_n_spl_,
    g139_n_spl_0
  );


  and

  (
    g141_p,
    input_f[6]_p_spl_10,
    input_w[3]_p_spl_01
  );


  or

  (
    g141_n,
    input_f[6]_n_spl_10,
    input_w[3]_n_spl_01
  );


  and

  (
    g142_p,
    input_f[5]_p_spl_10,
    input_w[4]_p_spl_01
  );


  or

  (
    g142_n,
    input_f[5]_n_spl_10,
    input_w[4]_n_spl_01
  );


  and

  (
    g143_p,
    g141_n,
    g142_n
  );


  or

  (
    g143_n,
    g141_p,
    g142_p
  );


  and

  (
    g144_p,
    g140_n_spl_,
    g143_n
  );


  or

  (
    g144_n,
    g140_p_spl_,
    g143_p
  );


  and

  (
    g145_p,
    g138_p_spl_,
    g144_p_spl_
  );


  or

  (
    g145_n,
    g138_n_spl_,
    g144_n_spl_
  );


  and

  (
    g146_p,
    g138_n_spl_,
    g144_n_spl_
  );


  or

  (
    g146_n,
    g138_p_spl_,
    g144_p_spl_
  );


  and

  (
    g147_p,
    g145_n_spl_,
    g146_n
  );


  or

  (
    g147_n,
    g145_p_spl_,
    g146_p
  );


  and

  (
    g148_p,
    input_f[6]_p_spl_10,
    input_w[2]_p_spl_00
  );


  or

  (
    g148_n,
    input_f[6]_n_spl_10,
    input_w[2]_n_spl_00
  );


  and

  (
    g149_p,
    g32_p_spl_,
    g148_n_spl_0
  );


  or

  (
    g149_n,
    g32_n_spl_,
    g148_p_spl_0
  );


  and

  (
    g150_p,
    g34_p_spl_0,
    g149_p
  );


  or

  (
    g150_n,
    g34_n_spl_0,
    g149_n
  );


  and

  (
    g151_p,
    g35_n_spl_,
    g150_n
  );


  or

  (
    g151_n,
    g35_p_spl_,
    g150_p
  );


  and

  (
    g152_p,
    g30_n_spl_0,
    g151_n
  );


  or

  (
    g152_n,
    g30_p_spl_0,
    g151_p
  );


  and

  (
    g153_p,
    g31_n_spl_1,
    g152_n
  );


  or

  (
    g153_n,
    g31_p_spl_1,
    g152_p
  );


  and

  (
    g154_p,
    g147_p_spl_,
    g153_p_spl_
  );


  or

  (
    g154_n,
    g147_n_spl_,
    g153_n_spl_
  );


  and

  (
    g155_p,
    g31_n_spl_1,
    g154_n_spl_
  );


  or

  (
    g155_n,
    g31_p_spl_1,
    g154_p_spl_
  );


  and

  (
    g156_p,
    g36_n_spl_1,
    g45_n_spl_
  );


  or

  (
    g156_n,
    g36_p_spl_1,
    g45_p_spl_
  );


  and

  (
    g157_p,
    g46_n_spl_,
    g156_n
  );


  or

  (
    g157_n,
    g46_p_spl_,
    g156_p
  );


  and

  (
    g158_p,
    g155_n_spl_,
    g157_p_spl_
  );


  or

  (
    g158_n,
    g155_p_spl_,
    g157_n_spl_
  );


  and

  (
    g159_p,
    input_f[3]_p_spl_00,
    input_w[6]_p_spl_10
  );


  or

  (
    g159_n,
    input_f[3]_n_spl_00,
    input_w[6]_n_spl_10
  );


  and

  (
    g160_p,
    input_f[2]_n_spl_00,
    input_w[7]_p_spl_01
  );


  or

  (
    g160_n,
    input_f[2]_p_spl_00,
    input_w[7]_n_spl_01
  );


  and

  (
    g161_p,
    g159_p_spl_,
    g160_p_spl_
  );


  or

  (
    g161_n,
    g159_n_spl_,
    g160_n_spl_
  );


  and

  (
    g162_p,
    g140_n_spl_,
    g145_n_spl_
  );


  or

  (
    g162_n,
    g140_p_spl_,
    g145_p_spl_
  );


  and

  (
    g163_p,
    g60_n_spl_,
    g61_n_spl_
  );


  or

  (
    g163_n,
    g60_p_spl_,
    g61_p_spl_
  );


  and

  (
    g164_p,
    g62_n_spl_,
    g163_n
  );


  or

  (
    g164_n,
    g62_p_spl_,
    g163_p
  );


  and

  (
    g165_p,
    g162_n_spl_,
    g164_p_spl_
  );


  or

  (
    g165_n,
    g162_p_spl_,
    g164_n_spl_
  );


  and

  (
    g166_p,
    g162_p_spl_,
    g164_n_spl_
  );


  or

  (
    g166_n,
    g162_n_spl_,
    g164_p_spl_
  );


  and

  (
    g167_p,
    g165_n_spl_,
    g166_n
  );


  or

  (
    g167_n,
    g165_p_spl_,
    g166_p
  );


  and

  (
    g168_p,
    g161_p_spl_0,
    g167_p_spl_
  );


  or

  (
    g168_n,
    g161_n_spl_0,
    g167_n_spl_
  );


  and

  (
    g169_p,
    g161_n_spl_0,
    g167_n_spl_
  );


  or

  (
    g169_n,
    g161_p_spl_0,
    g167_p_spl_
  );


  and

  (
    g170_p,
    g168_n_spl_,
    g169_n
  );


  or

  (
    g170_n,
    g168_p_spl_,
    g169_p
  );


  and

  (
    g171_p,
    g155_p_spl_,
    g157_n_spl_
  );


  or

  (
    g171_n,
    g155_n_spl_,
    g157_p_spl_
  );


  and

  (
    g172_p,
    g158_n_spl_,
    g171_n
  );


  or

  (
    g172_n,
    g158_p_spl_,
    g171_p
  );


  and

  (
    g173_p,
    g170_p_spl_,
    g172_p_spl_
  );


  or

  (
    g173_n,
    g170_n_spl_,
    g172_n_spl_
  );


  and

  (
    g174_p,
    g158_n_spl_,
    g173_n_spl_
  );


  or

  (
    g174_n,
    g158_p_spl_,
    g173_p_spl_
  );


  and

  (
    g175_p,
    g74_n_spl_,
    g76_n_spl_
  );


  or

  (
    g175_n,
    g74_p_spl_,
    g76_p_spl_
  );


  and

  (
    g176_p,
    g77_n_spl_,
    g175_n
  );


  or

  (
    g176_n,
    g77_p_spl_,
    g175_p
  );


  and

  (
    g177_p,
    g174_n_spl_,
    g176_p_spl_
  );


  or

  (
    g177_n,
    g174_p_spl_,
    g176_n_spl_
  );


  and

  (
    g178_p,
    g165_n_spl_,
    g168_n_spl_
  );


  or

  (
    g178_n,
    g165_p_spl_,
    g168_p_spl_
  );


  and

  (
    g179_p,
    g174_p_spl_,
    g176_n_spl_
  );


  or

  (
    g179_n,
    g174_n_spl_,
    g176_p_spl_
  );


  and

  (
    g180_p,
    g177_n_spl_,
    g179_n
  );


  or

  (
    g180_n,
    g177_p_spl_,
    g179_p
  );


  and

  (
    g181_p,
    g178_n_spl_,
    g180_p_spl_
  );


  or

  (
    g181_n,
    g178_p_spl_,
    g180_n_spl_
  );


  and

  (
    g182_p,
    g177_n_spl_,
    g181_n_spl_
  );


  or

  (
    g182_n,
    g177_p_spl_,
    g181_p_spl_
  );


  and

  (
    g183_p,
    g106_p_spl_,
    g108_n_spl_
  );


  or

  (
    g183_n,
    g106_n_spl_,
    g108_p_spl_
  );


  and

  (
    g184_p,
    g109_n_spl_,
    g183_n
  );


  or

  (
    g184_n,
    g109_p_spl_,
    g183_p
  );


  and

  (
    g185_p,
    g182_n_spl_,
    g184_p_spl_
  );


  or

  (
    g185_n,
    g182_p_spl_,
    g184_n_spl_
  );


  and

  (
    g186_p,
    input_w[7]_p_spl_01,
    g29_p_spl_0
  );


  or

  (
    g186_n,
    input_w[7]_n_spl_01,
    g29_n_spl_0
  );


  and

  (
    g187_p,
    input_f[6]_p_spl_11,
    input_w[1]_p_spl_00
  );


  or

  (
    g187_n,
    input_f[6]_n_spl_11,
    input_w[1]_n_spl_00
  );


  and

  (
    g188_p,
    input_w[7]_n_spl_10,
    g29_n_spl_
  );


  or

  (
    g188_n,
    input_w[7]_p_spl_10,
    g29_p_spl_
  );


  and

  (
    g189_p,
    g186_n_spl_,
    g188_n
  );


  or

  (
    g189_n,
    g186_p_spl_,
    g188_p
  );


  and

  (
    g190_p,
    g187_p_spl_0,
    g189_p_spl_
  );


  or

  (
    g190_n,
    g187_n_spl_0,
    g189_n_spl_
  );


  and

  (
    g191_p,
    g186_n_spl_,
    g190_n_spl_
  );


  or

  (
    g191_n,
    g186_p_spl_,
    g190_p_spl_
  );


  and

  (
    g192_p,
    g30_n_spl_,
    g34_p_spl_
  );


  or

  (
    g192_n,
    g30_p_spl_,
    g34_n_spl_
  );


  and

  (
    g193_p,
    g148_n_spl_0,
    g192_p_spl_
  );


  or

  (
    g193_n,
    g148_p_spl_0,
    g192_n_spl_
  );


  and

  (
    g194_p,
    g148_p_spl_,
    g192_n_spl_
  );


  or

  (
    g194_n,
    g148_n_spl_,
    g192_p_spl_
  );


  and

  (
    g195_p,
    g193_n,
    g194_n
  );


  or

  (
    g195_n,
    g193_p,
    g194_p
  );


  and

  (
    g196_p,
    g191_n_spl_,
    g195_n_spl_
  );


  or

  (
    g196_n,
    g191_p_spl_,
    g195_p_spl_
  );


  and

  (
    g197_p,
    input_f[3]_p_spl_01,
    input_w[5]_p_spl_10
  );


  or

  (
    g197_n,
    input_f[3]_n_spl_01,
    input_w[5]_n_spl_10
  );


  and

  (
    g198_p,
    input_f[4]_p_spl_01,
    input_w[4]_p_spl_01
  );


  or

  (
    g198_n,
    input_f[4]_n_spl_01,
    input_w[4]_n_spl_01
  );


  and

  (
    g199_p,
    g139_p_spl_0,
    g198_p_spl_
  );


  or

  (
    g199_n,
    g139_n_spl_0,
    g198_n_spl_
  );


  and

  (
    g200_p,
    g139_n_spl_1,
    g198_n_spl_
  );


  or

  (
    g200_n,
    g139_p_spl_1,
    g198_p_spl_
  );


  and

  (
    g201_p,
    g199_n_spl_,
    g200_n
  );


  or

  (
    g201_n,
    g199_p_spl_,
    g200_p
  );


  and

  (
    g202_p,
    g197_p_spl_,
    g201_p_spl_
  );


  or

  (
    g202_n,
    g197_n_spl_,
    g201_n_spl_
  );


  and

  (
    g203_p,
    g197_n_spl_,
    g201_n_spl_
  );


  or

  (
    g203_n,
    g197_p_spl_,
    g201_p_spl_
  );


  and

  (
    g204_p,
    g202_n_spl_,
    g203_n
  );


  or

  (
    g204_n,
    g202_p_spl_,
    g203_p
  );


  and

  (
    g205_p,
    g191_p_spl_,
    g195_p_spl_
  );


  or

  (
    g205_n,
    g191_n_spl_,
    g195_n_spl_
  );


  and

  (
    g206_p,
    g196_n_spl_,
    g205_n
  );


  or

  (
    g206_n,
    g196_p_spl_,
    g205_p
  );


  and

  (
    g207_p,
    g204_p_spl_,
    g206_p_spl_
  );


  or

  (
    g207_n,
    g204_n_spl_,
    g206_n_spl_
  );


  and

  (
    g208_p,
    g196_n_spl_,
    g207_n_spl_
  );


  or

  (
    g208_n,
    g196_p_spl_,
    g207_p_spl_
  );


  and

  (
    g209_p,
    g147_n_spl_,
    g153_n_spl_
  );


  or

  (
    g209_n,
    g147_p_spl_,
    g153_p_spl_
  );


  and

  (
    g210_p,
    g154_n_spl_,
    g209_n
  );


  or

  (
    g210_n,
    g154_p_spl_,
    g209_p
  );


  and

  (
    g211_p,
    g208_n_spl_,
    g210_p_spl_
  );


  or

  (
    g211_n,
    g208_p_spl_,
    g210_n_spl_
  );


  and

  (
    g212_p,
    input_f[2]_p_spl_00,
    input_w[6]_p_spl_10
  );


  or

  (
    g212_n,
    input_f[2]_n_spl_00,
    input_w[6]_n_spl_10
  );


  and

  (
    g213_p,
    input_f[1]_n_spl_00,
    input_w[7]_p_spl_10
  );


  or

  (
    g213_n,
    input_f[1]_p_spl_00,
    input_w[7]_n_spl_10
  );


  and

  (
    g214_p,
    g212_p_spl_0,
    g213_p_spl_
  );


  or

  (
    g214_n,
    g212_n_spl_0,
    g213_n_spl_
  );


  and

  (
    g215_p,
    g199_n_spl_,
    g202_n_spl_
  );


  or

  (
    g215_n,
    g199_p_spl_,
    g202_p_spl_
  );


  and

  (
    g216_p,
    g159_n_spl_,
    g160_n_spl_
  );


  or

  (
    g216_n,
    g159_p_spl_,
    g160_p_spl_
  );


  and

  (
    g217_p,
    g161_n_spl_,
    g216_n
  );


  or

  (
    g217_n,
    g161_p_spl_,
    g216_p
  );


  and

  (
    g218_p,
    g215_n_spl_,
    g217_p_spl_
  );


  or

  (
    g218_n,
    g215_p_spl_,
    g217_n_spl_
  );


  and

  (
    g219_p,
    g215_p_spl_,
    g217_n_spl_
  );


  or

  (
    g219_n,
    g215_n_spl_,
    g217_p_spl_
  );


  and

  (
    g220_p,
    g218_n_spl_,
    g219_n
  );


  or

  (
    g220_n,
    g218_p_spl_,
    g219_p
  );


  and

  (
    g221_p,
    g214_p_spl_0,
    g220_p_spl_
  );


  or

  (
    g221_n,
    g214_n_spl_0,
    g220_n_spl_
  );


  and

  (
    g222_p,
    g214_n_spl_0,
    g220_n_spl_
  );


  or

  (
    g222_n,
    g214_p_spl_0,
    g220_p_spl_
  );


  and

  (
    g223_p,
    g221_n_spl_,
    g222_n
  );


  or

  (
    g223_n,
    g221_p_spl_,
    g222_p
  );


  and

  (
    g224_p,
    g208_p_spl_,
    g210_n_spl_
  );


  or

  (
    g224_n,
    g208_n_spl_,
    g210_p_spl_
  );


  and

  (
    g225_p,
    g211_n_spl_,
    g224_n
  );


  or

  (
    g225_n,
    g211_p_spl_,
    g224_p
  );


  and

  (
    g226_p,
    g223_p_spl_,
    g225_p_spl_
  );


  or

  (
    g226_n,
    g223_n_spl_,
    g225_n_spl_
  );


  and

  (
    g227_p,
    g211_n_spl_,
    g226_n_spl_
  );


  or

  (
    g227_n,
    g211_p_spl_,
    g226_p_spl_
  );


  and

  (
    g228_p,
    g170_n_spl_,
    g172_n_spl_
  );


  or

  (
    g228_n,
    g170_p_spl_,
    g172_p_spl_
  );


  and

  (
    g229_p,
    g173_n_spl_,
    g228_n
  );


  or

  (
    g229_n,
    g173_p_spl_,
    g228_p
  );


  and

  (
    g230_p,
    g227_n_spl_,
    g229_p_spl_
  );


  or

  (
    g230_n,
    g227_p_spl_,
    g229_n_spl_
  );


  and

  (
    g231_p,
    g218_n_spl_,
    g221_n_spl_
  );


  or

  (
    g231_n,
    g218_p_spl_,
    g221_p_spl_
  );


  and

  (
    g232_p,
    g227_p_spl_,
    g229_n_spl_
  );


  or

  (
    g232_n,
    g227_n_spl_,
    g229_p_spl_
  );


  and

  (
    g233_p,
    g230_n_spl_,
    g232_n
  );


  or

  (
    g233_n,
    g230_p_spl_,
    g232_p
  );


  and

  (
    g234_p,
    g231_n_spl_,
    g233_p_spl_
  );


  or

  (
    g234_n,
    g231_p_spl_,
    g233_n_spl_
  );


  and

  (
    g235_p,
    g230_n_spl_,
    g234_n_spl_
  );


  or

  (
    g235_n,
    g230_p_spl_,
    g234_p_spl_
  );


  and

  (
    g236_p,
    g178_p_spl_,
    g180_n_spl_
  );


  or

  (
    g236_n,
    g178_n_spl_,
    g180_p_spl_
  );


  and

  (
    g237_p,
    g181_n_spl_,
    g236_n
  );


  or

  (
    g237_n,
    g181_p_spl_,
    g236_p
  );


  and

  (
    g238_p,
    g235_n_spl_,
    g237_p_spl_
  );


  or

  (
    g238_n,
    g235_p_spl_,
    g237_n_spl_
  );


  and

  (
    g239_p,
    g235_p_spl_,
    g237_n_spl_
  );


  or

  (
    g239_n,
    g235_n_spl_,
    g237_p_spl_
  );


  and

  (
    g240_p,
    g238_n_spl_,
    g239_n
  );


  or

  (
    g240_n,
    g238_p_spl_,
    g239_p
  );


  and

  (
    g241_p,
    input_f[5]_p_spl_10,
    input_w[0]_p_spl_00
  );


  or

  (
    g241_n,
    input_f[5]_n_spl_10,
    input_w[0]_n_spl_00
  );


  and

  (
    g242_p,
    g187_p_spl_0,
    g241_p_spl_0
  );


  or

  (
    g242_n,
    g187_n_spl_0,
    g241_n_spl_0
  );


  and

  (
    g243_p,
    input_f[4]_p_spl_10,
    input_w[2]_p_spl_01
  );


  or

  (
    g243_n,
    input_f[4]_n_spl_10,
    input_w[2]_n_spl_01
  );


  and

  (
    g244_p,
    input_f[6]_p_spl_11,
    input_w[0]_p_spl_01
  );


  or

  (
    g244_n,
    input_f[6]_n_spl_11,
    input_w[0]_n_spl_01
  );


  and

  (
    g245_p,
    input_f[5]_p_spl_11,
    input_w[1]_p_spl_01
  );


  or

  (
    g245_n,
    input_f[5]_n_spl_11,
    input_w[1]_n_spl_01
  );


  and

  (
    g246_p,
    g244_n,
    g245_n
  );


  or

  (
    g246_n,
    g244_p,
    g245_p
  );


  and

  (
    g247_p,
    g242_n_spl_,
    g246_n
  );


  or

  (
    g247_n,
    g242_p_spl_,
    g246_p
  );


  and

  (
    g248_p,
    g243_p_spl_0,
    g247_p_spl_
  );


  or

  (
    g248_n,
    g243_n_spl_0,
    g247_n_spl_
  );


  and

  (
    g249_p,
    g242_n_spl_,
    g248_n_spl_
  );


  or

  (
    g249_n,
    g242_p_spl_,
    g248_p_spl_
  );


  and

  (
    g250_p,
    g187_n_spl_,
    g189_n_spl_
  );


  or

  (
    g250_n,
    g187_p_spl_,
    g189_p_spl_
  );


  and

  (
    g251_p,
    g190_n_spl_,
    g250_n
  );


  or

  (
    g251_n,
    g190_p_spl_,
    g250_p
  );


  and

  (
    g252_p,
    g249_n_spl_,
    g251_p_spl_
  );


  or

  (
    g252_n,
    g249_p_spl_,
    g251_n_spl_
  );


  and

  (
    g253_p,
    g249_p_spl_,
    g251_n_spl_
  );


  or

  (
    g253_n,
    g249_n_spl_,
    g251_p_spl_
  );


  and

  (
    g254_p,
    g252_n_spl_,
    g253_n
  );


  or

  (
    g254_n,
    g252_p_spl_,
    g253_p
  );


  and

  (
    g255_p,
    input_f[3]_p_spl_01,
    input_w[4]_p_spl_10
  );


  or

  (
    g255_n,
    input_f[3]_n_spl_01,
    input_w[4]_n_spl_10
  );


  and

  (
    g256_p,
    g139_p_spl_1,
    g243_p_spl_0
  );


  or

  (
    g256_n,
    g139_n_spl_1,
    g243_n_spl_0
  );


  and

  (
    g257_p,
    input_f[4]_p_spl_10,
    input_w[3]_p_spl_01
  );


  or

  (
    g257_n,
    input_f[4]_n_spl_10,
    input_w[3]_n_spl_01
  );


  and

  (
    g258_p,
    input_f[5]_p_spl_11,
    input_w[2]_p_spl_01
  );


  or

  (
    g258_n,
    input_f[5]_n_spl_11,
    input_w[2]_n_spl_01
  );


  and

  (
    g259_p,
    g257_n,
    g258_n
  );


  or

  (
    g259_n,
    g257_p,
    g258_p
  );


  and

  (
    g260_p,
    g256_n_spl_,
    g259_n
  );


  or

  (
    g260_n,
    g256_p_spl_,
    g259_p
  );


  and

  (
    g261_p,
    g255_p_spl_0,
    g260_p_spl_
  );


  or

  (
    g261_n,
    g255_n_spl_0,
    g260_n_spl_
  );


  and

  (
    g262_p,
    g255_n_spl_0,
    g260_n_spl_
  );


  or

  (
    g262_n,
    g255_p_spl_0,
    g260_p_spl_
  );


  and

  (
    g263_p,
    g261_n_spl_,
    g262_n
  );


  or

  (
    g263_n,
    g261_p_spl_,
    g262_p
  );


  and

  (
    g264_p,
    g254_p_spl_,
    g263_p_spl_
  );


  or

  (
    g264_n,
    g254_n_spl_,
    g263_n_spl_
  );


  and

  (
    g265_p,
    g252_n_spl_,
    g264_n_spl_
  );


  or

  (
    g265_n,
    g252_p_spl_,
    g264_p_spl_
  );


  and

  (
    g266_p,
    g204_n_spl_,
    g206_n_spl_
  );


  or

  (
    g266_n,
    g204_p_spl_,
    g206_p_spl_
  );


  and

  (
    g267_p,
    g207_n_spl_,
    g266_n
  );


  or

  (
    g267_n,
    g207_p_spl_,
    g266_p
  );


  and

  (
    g268_p,
    g265_n_spl_,
    g267_p_spl_
  );


  or

  (
    g268_n,
    g265_p_spl_,
    g267_n_spl_
  );


  and

  (
    g269_p,
    input_f[1]_p_spl_00,
    input_w[5]_p_spl_10
  );


  or

  (
    g269_n,
    input_f[1]_n_spl_00,
    input_w[5]_n_spl_10
  );


  and

  (
    g270_p,
    g212_p_spl_0,
    g269_p_spl_0
  );


  or

  (
    g270_n,
    g212_n_spl_0,
    g269_n_spl_0
  );


  and

  (
    g271_p,
    input_f[0]_n_spl_00,
    input_w[7]_p_spl_11
  );


  or

  (
    g271_n,
    input_f[0]_p_spl_00,
    input_w[7]_n_spl_11
  );


  and

  (
    g272_p,
    input_f[2]_p_spl_01,
    input_w[5]_p_spl_11
  );


  or

  (
    g272_n,
    input_f[2]_n_spl_01,
    input_w[5]_n_spl_11
  );


  and

  (
    g273_p,
    input_f[1]_p_spl_01,
    input_w[6]_p_spl_11
  );


  or

  (
    g273_n,
    input_f[1]_n_spl_01,
    input_w[6]_n_spl_11
  );


  and

  (
    g274_p,
    g272_n,
    g273_n
  );


  or

  (
    g274_n,
    g272_p,
    g273_p
  );


  and

  (
    g275_p,
    g270_n_spl_,
    g274_n
  );


  or

  (
    g275_n,
    g270_p_spl_,
    g274_p
  );


  and

  (
    g276_p,
    g271_p_spl_,
    g275_p_spl_
  );


  or

  (
    g276_n,
    g271_n_spl_,
    g275_n_spl_
  );


  and

  (
    g277_p,
    g270_n_spl_,
    g276_n_spl_
  );


  or

  (
    g277_n,
    g270_p_spl_,
    g276_p_spl_
  );


  and

  (
    g278_p,
    g256_n_spl_,
    g261_n_spl_
  );


  or

  (
    g278_n,
    g256_p_spl_,
    g261_p_spl_
  );


  and

  (
    g279_p,
    g212_n_spl_,
    g213_n_spl_
  );


  or

  (
    g279_n,
    g212_p_spl_,
    g213_p_spl_
  );


  and

  (
    g280_p,
    g214_n_spl_,
    g279_n
  );


  or

  (
    g280_n,
    g214_p_spl_,
    g279_p
  );


  and

  (
    g281_p,
    g278_n_spl_,
    g280_p_spl_
  );


  or

  (
    g281_n,
    g278_p_spl_,
    g280_n_spl_
  );


  and

  (
    g282_p,
    g278_p_spl_,
    g280_n_spl_
  );


  or

  (
    g282_n,
    g278_n_spl_,
    g280_p_spl_
  );


  and

  (
    g283_p,
    g281_n_spl_,
    g282_n
  );


  or

  (
    g283_n,
    g281_p_spl_,
    g282_p
  );


  and

  (
    g284_p,
    g277_n_spl_,
    g283_p_spl_
  );


  or

  (
    g284_n,
    g277_p_spl_,
    g283_n_spl_
  );


  and

  (
    g285_p,
    g277_p_spl_,
    g283_n_spl_
  );


  or

  (
    g285_n,
    g277_n_spl_,
    g283_p_spl_
  );


  and

  (
    g286_p,
    g284_n_spl_,
    g285_n
  );


  or

  (
    g286_n,
    g284_p_spl_,
    g285_p
  );


  and

  (
    g287_p,
    g265_p_spl_,
    g267_n_spl_
  );


  or

  (
    g287_n,
    g265_n_spl_,
    g267_p_spl_
  );


  and

  (
    g288_p,
    g268_n_spl_,
    g287_n
  );


  or

  (
    g288_n,
    g268_p_spl_,
    g287_p
  );


  and

  (
    g289_p,
    g286_p_spl_,
    g288_p_spl_
  );


  or

  (
    g289_n,
    g286_n_spl_,
    g288_n_spl_
  );


  and

  (
    g290_p,
    g268_n_spl_,
    g289_n_spl_
  );


  or

  (
    g290_n,
    g268_p_spl_,
    g289_p_spl_
  );


  and

  (
    g291_p,
    g223_n_spl_,
    g225_n_spl_
  );


  or

  (
    g291_n,
    g223_p_spl_,
    g225_p_spl_
  );


  and

  (
    g292_p,
    g226_n_spl_,
    g291_n
  );


  or

  (
    g292_n,
    g226_p_spl_,
    g291_p
  );


  and

  (
    g293_p,
    g290_n_spl_,
    g292_p_spl_
  );


  or

  (
    g293_n,
    g290_p_spl_,
    g292_n_spl_
  );


  and

  (
    g294_p,
    g281_n_spl_,
    g284_n_spl_
  );


  or

  (
    g294_n,
    g281_p_spl_,
    g284_p_spl_
  );


  and

  (
    g295_p,
    g290_p_spl_,
    g292_n_spl_
  );


  or

  (
    g295_n,
    g290_n_spl_,
    g292_p_spl_
  );


  and

  (
    g296_p,
    g293_n_spl_,
    g295_n
  );


  or

  (
    g296_n,
    g293_p_spl_,
    g295_p
  );


  and

  (
    g297_p,
    g294_n_spl_,
    g296_p_spl_
  );


  or

  (
    g297_n,
    g294_p_spl_,
    g296_n_spl_
  );


  and

  (
    g298_p,
    g293_n_spl_,
    g297_n_spl_
  );


  or

  (
    g298_n,
    g293_p_spl_,
    g297_p_spl_
  );


  and

  (
    g299_p,
    g231_p_spl_,
    g233_n_spl_
  );


  or

  (
    g299_n,
    g231_n_spl_,
    g233_p_spl_
  );


  and

  (
    g300_p,
    g234_n_spl_,
    g299_n
  );


  or

  (
    g300_n,
    g234_p_spl_,
    g299_p
  );


  and

  (
    g301_p,
    g298_n_spl_,
    g300_p_spl_
  );


  or

  (
    g301_n,
    g298_p_spl_,
    g300_n_spl_
  );


  and

  (
    g302_p,
    g298_p_spl_,
    g300_n_spl_
  );


  or

  (
    g302_n,
    g298_n_spl_,
    g300_p_spl_
  );


  and

  (
    g303_p,
    g301_n_spl_,
    g302_n
  );


  or

  (
    g303_n,
    g301_p_spl_,
    g302_p
  );


  and

  (
    g304_p,
    input_f[4]_p_spl_11,
    input_w[1]_p_spl_01
  );


  or

  (
    g304_n,
    input_f[4]_n_spl_11,
    input_w[1]_n_spl_01
  );


  and

  (
    g305_p,
    g241_p_spl_0,
    g304_p_spl_
  );


  or

  (
    g305_n,
    g241_n_spl_0,
    g304_n_spl_
  );


  and

  (
    g306_p,
    input_f[3]_p_spl_10,
    input_w[2]_p_spl_10
  );


  or

  (
    g306_n,
    input_f[3]_n_spl_10,
    input_w[2]_n_spl_10
  );


  and

  (
    g307_p,
    g241_n_spl_,
    g304_n_spl_
  );


  or

  (
    g307_n,
    g241_p_spl_,
    g304_p_spl_
  );


  and

  (
    g308_p,
    g305_n_spl_,
    g307_n
  );


  or

  (
    g308_n,
    g305_p_spl_,
    g307_p
  );


  and

  (
    g309_p,
    g306_p_spl_,
    g308_p_spl_
  );


  or

  (
    g309_n,
    g306_n_spl_,
    g308_n_spl_
  );


  and

  (
    g310_p,
    g305_n_spl_,
    g309_n_spl_
  );


  or

  (
    g310_n,
    g305_p_spl_,
    g309_p_spl_
  );


  and

  (
    g311_p,
    g243_n_spl_,
    g247_n_spl_
  );


  or

  (
    g311_n,
    g243_p_spl_,
    g247_p_spl_
  );


  and

  (
    g312_p,
    g248_n_spl_,
    g311_n
  );


  or

  (
    g312_n,
    g248_p_spl_,
    g311_p
  );


  and

  (
    g313_p,
    g310_n_spl_,
    g312_p_spl_
  );


  or

  (
    g313_n,
    g310_p_spl_,
    g312_n_spl_
  );


  and

  (
    g314_p,
    input_f[2]_p_spl_01,
    input_w[3]_p_spl_10
  );


  or

  (
    g314_n,
    input_f[2]_n_spl_01,
    input_w[3]_n_spl_10
  );


  and

  (
    g315_p,
    g255_p_spl_,
    g314_p_spl_0
  );


  or

  (
    g315_n,
    g255_n_spl_,
    g314_n_spl_0
  );


  and

  (
    g316_p,
    input_f[3]_p_spl_10,
    input_w[3]_p_spl_10
  );


  or

  (
    g316_n,
    input_f[3]_n_spl_10,
    input_w[3]_n_spl_10
  );


  and

  (
    g317_p,
    input_f[2]_p_spl_10,
    input_w[4]_p_spl_10
  );


  or

  (
    g317_n,
    input_f[2]_n_spl_10,
    input_w[4]_n_spl_10
  );


  and

  (
    g318_p,
    g316_n,
    g317_n
  );


  or

  (
    g318_n,
    g316_p,
    g317_p
  );


  and

  (
    g319_p,
    g315_n_spl_,
    g318_n
  );


  or

  (
    g319_n,
    g315_p_spl_,
    g318_p
  );


  and

  (
    g320_p,
    g269_p_spl_0,
    g319_p_spl_
  );


  or

  (
    g320_n,
    g269_n_spl_0,
    g319_n_spl_
  );


  and

  (
    g321_p,
    g269_n_spl_,
    g319_n_spl_
  );


  or

  (
    g321_n,
    g269_p_spl_,
    g319_p_spl_
  );


  and

  (
    g322_p,
    g320_n_spl_,
    g321_n
  );


  or

  (
    g322_n,
    g320_p_spl_,
    g321_p
  );


  and

  (
    g323_p,
    g310_p_spl_,
    g312_n_spl_
  );


  or

  (
    g323_n,
    g310_n_spl_,
    g312_p_spl_
  );


  and

  (
    g324_p,
    g313_n_spl_,
    g323_n
  );


  or

  (
    g324_n,
    g313_p_spl_,
    g323_p
  );


  and

  (
    g325_p,
    g322_p_spl_,
    g324_p_spl_
  );


  or

  (
    g325_n,
    g322_n_spl_,
    g324_n_spl_
  );


  and

  (
    g326_p,
    g313_n_spl_,
    g325_n_spl_
  );


  or

  (
    g326_n,
    g313_p_spl_,
    g325_p_spl_
  );


  and

  (
    g327_p,
    g254_n_spl_,
    g263_n_spl_
  );


  or

  (
    g327_n,
    g254_p_spl_,
    g263_p_spl_
  );


  and

  (
    g328_p,
    g264_n_spl_,
    g327_n
  );


  or

  (
    g328_n,
    g264_p_spl_,
    g327_p
  );


  and

  (
    g329_p,
    g326_n_spl_,
    g328_p_spl_
  );


  or

  (
    g329_n,
    g326_p_spl_,
    g328_n_spl_
  );


  and

  (
    g330_p,
    g326_p_spl_,
    g328_n_spl_
  );


  or

  (
    g330_n,
    g326_n_spl_,
    g328_p_spl_
  );


  and

  (
    g331_p,
    g329_n_spl_,
    g330_n
  );


  or

  (
    g331_n,
    g329_p_spl_,
    g330_p
  );


  and

  (
    g332_p,
    g315_n_spl_,
    g320_n_spl_
  );


  or

  (
    g332_n,
    g315_p_spl_,
    g320_p_spl_
  );


  and

  (
    g333_p,
    g271_n_spl_,
    g275_n_spl_
  );


  or

  (
    g333_n,
    g271_p_spl_,
    g275_p_spl_
  );


  and

  (
    g334_p,
    g276_n_spl_,
    g333_n
  );


  or

  (
    g334_n,
    g276_p_spl_,
    g333_p
  );


  and

  (
    g335_p,
    g332_n_spl_,
    g334_p_spl_
  );


  or

  (
    g335_n,
    g332_p_spl_,
    g334_n_spl_
  );


  and

  (
    g336_p,
    g332_p_spl_,
    g334_n_spl_
  );


  or

  (
    g336_n,
    g332_n_spl_,
    g334_p_spl_
  );


  and

  (
    g337_p,
    g335_n_spl_0,
    g336_n
  );


  or

  (
    g337_n,
    g335_p_spl_0,
    g336_p
  );


  and

  (
    g338_p,
    g331_p_spl_,
    g337_p_spl_
  );


  or

  (
    g338_n,
    g331_n_spl_,
    g337_n_spl_
  );


  and

  (
    g339_p,
    g329_n_spl_,
    g338_n_spl_
  );


  or

  (
    g339_n,
    g329_p_spl_,
    g338_p_spl_
  );


  and

  (
    g340_p,
    g286_n_spl_,
    g288_n_spl_
  );


  or

  (
    g340_n,
    g286_p_spl_,
    g288_p_spl_
  );


  and

  (
    g341_p,
    g289_n_spl_,
    g340_n
  );


  or

  (
    g341_n,
    g289_p_spl_,
    g340_p
  );


  and

  (
    g342_p,
    g339_n_spl_,
    g341_p_spl_
  );


  or

  (
    g342_n,
    g339_p_spl_,
    g341_n_spl_
  );


  and

  (
    g343_p,
    g339_p_spl_,
    g341_n_spl_
  );


  or

  (
    g343_n,
    g339_n_spl_,
    g341_p_spl_
  );


  and

  (
    g344_p,
    g342_n_spl_,
    g343_n
  );


  or

  (
    g344_n,
    g342_p_spl_,
    g343_p
  );


  and

  (
    g345_p,
    g335_p_spl_0,
    g344_p_spl_
  );


  or

  (
    g345_n,
    g335_n_spl_0,
    g344_n_spl_
  );


  and

  (
    g346_p,
    g342_n_spl_,
    g345_n_spl_
  );


  or

  (
    g346_n,
    g342_p_spl_,
    g345_p_spl_
  );


  and

  (
    g347_p,
    g294_p_spl_,
    g296_n_spl_
  );


  or

  (
    g347_n,
    g294_n_spl_,
    g296_p_spl_
  );


  and

  (
    g348_p,
    g297_n_spl_,
    g347_n
  );


  or

  (
    g348_n,
    g297_p_spl_,
    g347_p
  );


  and

  (
    g349_p,
    g346_n_spl_,
    g348_p_spl_
  );


  or

  (
    g349_n,
    g346_p_spl_,
    g348_n_spl_
  );


  and

  (
    g350_p,
    input_f[4]_p_spl_11,
    input_w[0]_p_spl_01
  );


  or

  (
    g350_n,
    input_f[4]_n_spl_11,
    input_w[0]_n_spl_01
  );


  and

  (
    g351_p,
    input_f[3]_p_spl_11,
    input_w[1]_p_spl_10
  );


  or

  (
    g351_n,
    input_f[3]_n_spl_11,
    input_w[1]_n_spl_10
  );


  and

  (
    g352_p,
    g350_p_spl_,
    g351_p_spl_0
  );


  or

  (
    g352_n,
    g350_n_spl_,
    g351_n_spl_0
  );


  and

  (
    g353_p,
    input_f[2]_p_spl_10,
    input_w[2]_p_spl_10
  );


  or

  (
    g353_n,
    input_f[2]_n_spl_10,
    input_w[2]_n_spl_10
  );


  and

  (
    g354_p,
    g350_n_spl_,
    g351_n_spl_0
  );


  or

  (
    g354_n,
    g350_p_spl_,
    g351_p_spl_0
  );


  and

  (
    g355_p,
    g352_n_spl_,
    g354_n
  );


  or

  (
    g355_n,
    g352_p_spl_,
    g354_p
  );


  and

  (
    g356_p,
    g353_p_spl_,
    g355_p_spl_
  );


  or

  (
    g356_n,
    g353_n_spl_,
    g355_n_spl_
  );


  and

  (
    g357_p,
    g352_n_spl_,
    g356_n_spl_
  );


  or

  (
    g357_n,
    g352_p_spl_,
    g356_p_spl_
  );


  and

  (
    g358_p,
    g306_n_spl_,
    g308_n_spl_
  );


  or

  (
    g358_n,
    g306_p_spl_,
    g308_p_spl_
  );


  and

  (
    g359_p,
    g309_n_spl_,
    g358_n
  );


  or

  (
    g359_n,
    g309_p_spl_,
    g358_p
  );


  and

  (
    g360_p,
    g357_n_spl_,
    g359_p_spl_
  );


  or

  (
    g360_n,
    g357_p_spl_,
    g359_n_spl_
  );


  and

  (
    g361_p,
    input_f[0]_p_spl_00,
    input_w[5]_p_spl_11
  );


  or

  (
    g361_n,
    input_f[0]_n_spl_00,
    input_w[5]_n_spl_11
  );


  and

  (
    g362_p,
    input_f[1]_p_spl_01,
    input_w[4]_p_spl_11
  );


  or

  (
    g362_n,
    input_f[1]_n_spl_01,
    input_w[4]_n_spl_11
  );


  and

  (
    g363_p,
    g314_p_spl_0,
    g362_p_spl_0
  );


  or

  (
    g363_n,
    g314_n_spl_0,
    g362_n_spl_0
  );


  and

  (
    g364_p,
    g314_n_spl_,
    g362_n_spl_0
  );


  or

  (
    g364_n,
    g314_p_spl_,
    g362_p_spl_0
  );


  and

  (
    g365_p,
    g363_n_spl_,
    g364_n
  );


  or

  (
    g365_n,
    g363_p_spl_,
    g364_p
  );


  and

  (
    g366_p,
    g361_p_spl_,
    g365_p_spl_
  );


  or

  (
    g366_n,
    g361_n_spl_,
    g365_n_spl_
  );


  and

  (
    g367_p,
    g361_n_spl_,
    g365_n_spl_
  );


  or

  (
    g367_n,
    g361_p_spl_,
    g365_p_spl_
  );


  and

  (
    g368_p,
    g366_n_spl_,
    g367_n
  );


  or

  (
    g368_n,
    g366_p_spl_,
    g367_p
  );


  and

  (
    g369_p,
    g357_p_spl_,
    g359_n_spl_
  );


  or

  (
    g369_n,
    g357_n_spl_,
    g359_p_spl_
  );


  and

  (
    g370_p,
    g360_n_spl_,
    g369_n
  );


  or

  (
    g370_n,
    g360_p_spl_,
    g369_p
  );


  and

  (
    g371_p,
    g368_p_spl_,
    g370_p_spl_
  );


  or

  (
    g371_n,
    g368_n_spl_,
    g370_n_spl_
  );


  and

  (
    g372_p,
    g360_n_spl_,
    g371_n_spl_
  );


  or

  (
    g372_n,
    g360_p_spl_,
    g371_p_spl_
  );


  and

  (
    g373_p,
    g322_n_spl_,
    g324_n_spl_
  );


  or

  (
    g373_n,
    g322_p_spl_,
    g324_p_spl_
  );


  and

  (
    g374_p,
    g325_n_spl_,
    g373_n
  );


  or

  (
    g374_n,
    g325_p_spl_,
    g373_p
  );


  and

  (
    g375_p,
    g372_n_spl_,
    g374_p_spl_
  );


  or

  (
    g375_n,
    g372_p_spl_,
    g374_n_spl_
  );


  and

  (
    g376_p,
    g363_n_spl_,
    g366_n_spl_
  );


  or

  (
    g376_n,
    g363_p_spl_,
    g366_p_spl_
  );


  and

  (
    g377_p,
    input_f[0]_p_spl_01,
    input_w[6]_p_spl_11
  );


  or

  (
    g377_n,
    input_f[0]_n_spl_01,
    input_w[6]_n_spl_11
  );


  and

  (
    g378_p,
    g376_n_spl_,
    g377_p_spl_
  );


  or

  (
    g378_n,
    g376_p_spl_,
    g377_n_spl_
  );


  and

  (
    g379_p,
    g376_p_spl_,
    g377_n_spl_
  );


  or

  (
    g379_n,
    g376_n_spl_,
    g377_p_spl_
  );


  and

  (
    g380_p,
    g378_n_spl_0,
    g379_n
  );


  or

  (
    g380_n,
    g378_p_spl_0,
    g379_p
  );


  and

  (
    g381_p,
    g372_p_spl_,
    g374_n_spl_
  );


  or

  (
    g381_n,
    g372_n_spl_,
    g374_p_spl_
  );


  and

  (
    g382_p,
    g375_n_spl_,
    g381_n
  );


  or

  (
    g382_n,
    g375_p_spl_,
    g381_p
  );


  and

  (
    g383_p,
    g380_p_spl_,
    g382_p_spl_
  );


  or

  (
    g383_n,
    g380_n_spl_,
    g382_n_spl_
  );


  and

  (
    g384_p,
    g375_n_spl_,
    g383_n_spl_
  );


  or

  (
    g384_n,
    g375_p_spl_,
    g383_p_spl_
  );


  and

  (
    g385_p,
    g331_n_spl_,
    g337_n_spl_
  );


  or

  (
    g385_n,
    g331_p_spl_,
    g337_p_spl_
  );


  and

  (
    g386_p,
    g338_n_spl_,
    g385_n
  );


  or

  (
    g386_n,
    g338_p_spl_,
    g385_p
  );


  and

  (
    g387_p,
    g384_n_spl_,
    g386_p_spl_
  );


  or

  (
    g387_n,
    g384_p_spl_,
    g386_n_spl_
  );


  and

  (
    g388_p,
    g384_p_spl_,
    g386_n_spl_
  );


  or

  (
    g388_n,
    g384_n_spl_,
    g386_p_spl_
  );


  and

  (
    g389_p,
    g387_n_spl_,
    g388_n
  );


  or

  (
    g389_n,
    g387_p_spl_,
    g388_p
  );


  and

  (
    g390_p,
    g378_p_spl_0,
    g389_p_spl_
  );


  or

  (
    g390_n,
    g378_n_spl_0,
    g389_n_spl_
  );


  and

  (
    g391_p,
    g387_n_spl_,
    g390_n_spl_
  );


  or

  (
    g391_n,
    g387_p_spl_,
    g390_p_spl_
  );


  and

  (
    g392_p,
    g335_n_spl_,
    g344_n_spl_
  );


  or

  (
    g392_n,
    g335_p_spl_,
    g344_p_spl_
  );


  and

  (
    g393_p,
    g345_n_spl_,
    g392_n
  );


  or

  (
    g393_n,
    g345_p_spl_,
    g392_p
  );


  and

  (
    g394_p,
    g391_n_spl_,
    g393_p_spl_
  );


  or

  (
    g394_n,
    g391_p_spl_,
    g393_n_spl_
  );


  and

  (
    g395_p,
    input_f[2]_p_spl_11,
    input_w[0]_p_spl_10
  );


  or

  (
    g395_n,
    input_f[2]_n_spl_11,
    input_w[0]_n_spl_10
  );


  and

  (
    g396_p,
    g351_p_spl_,
    g395_p_spl_0
  );


  or

  (
    g396_n,
    g351_n_spl_,
    g395_n_spl_0
  );


  and

  (
    g397_p,
    input_f[1]_p_spl_10,
    input_w[2]_p_spl_11
  );


  or

  (
    g397_n,
    input_f[1]_n_spl_10,
    input_w[2]_n_spl_11
  );


  and

  (
    g398_p,
    input_f[3]_p_spl_11,
    input_w[0]_p_spl_10
  );


  or

  (
    g398_n,
    input_f[3]_n_spl_11,
    input_w[0]_n_spl_10
  );


  and

  (
    g399_p,
    input_f[2]_p_spl_11,
    input_w[1]_p_spl_10
  );


  or

  (
    g399_n,
    input_f[2]_n_spl_11,
    input_w[1]_n_spl_10
  );


  and

  (
    g400_p,
    g398_n,
    g399_n
  );


  or

  (
    g400_n,
    g398_p,
    g399_p
  );


  and

  (
    g401_p,
    g396_n_spl_,
    g400_n
  );


  or

  (
    g401_n,
    g396_p_spl_,
    g400_p
  );


  and

  (
    g402_p,
    g397_p_spl_,
    g401_p_spl_
  );


  or

  (
    g402_n,
    g397_n_spl_,
    g401_n_spl_
  );


  and

  (
    g403_p,
    g396_n_spl_,
    g402_n_spl_
  );


  or

  (
    g403_n,
    g396_p_spl_,
    g402_p_spl_
  );


  and

  (
    g404_p,
    g353_n_spl_,
    g355_n_spl_
  );


  or

  (
    g404_n,
    g353_p_spl_,
    g355_p_spl_
  );


  and

  (
    g405_p,
    g356_n_spl_,
    g404_n
  );


  or

  (
    g405_n,
    g356_p_spl_,
    g404_p
  );


  and

  (
    g406_p,
    g403_n_spl_,
    g405_p_spl_
  );


  or

  (
    g406_n,
    g403_p_spl_,
    g405_n_spl_
  );


  and

  (
    g407_p,
    input_f[0]_p_spl_01,
    input_w[3]_p_spl_11
  );


  or

  (
    g407_n,
    input_f[0]_n_spl_01,
    input_w[3]_n_spl_11
  );


  and

  (
    g408_p,
    g362_p_spl_,
    g407_p_spl_0
  );


  or

  (
    g408_n,
    g362_n_spl_,
    g407_n_spl_0
  );


  and

  (
    g409_p,
    input_f[1]_p_spl_10,
    input_w[3]_p_spl_11
  );


  or

  (
    g409_n,
    input_f[1]_n_spl_10,
    input_w[3]_n_spl_11
  );


  and

  (
    g410_p,
    input_f[0]_p_spl_10,
    input_w[4]_p_spl_11
  );


  or

  (
    g410_n,
    input_f[0]_n_spl_10,
    input_w[4]_n_spl_11
  );


  and

  (
    g411_p,
    g409_n,
    g410_n
  );


  or

  (
    g411_n,
    g409_p,
    g410_p
  );


  and

  (
    g412_p,
    g408_n_spl_0,
    g411_n
  );


  or

  (
    g412_n,
    g408_p_spl_0,
    g411_p
  );


  and

  (
    g413_p,
    g403_p_spl_,
    g405_n_spl_
  );


  or

  (
    g413_n,
    g403_n_spl_,
    g405_p_spl_
  );


  and

  (
    g414_p,
    g406_n_spl_,
    g413_n
  );


  or

  (
    g414_n,
    g406_p_spl_,
    g413_p
  );


  and

  (
    g415_p,
    g412_p_spl_,
    g414_p_spl_
  );


  or

  (
    g415_n,
    g412_n_spl_,
    g414_n_spl_
  );


  and

  (
    g416_p,
    g406_n_spl_,
    g415_n_spl_
  );


  or

  (
    g416_n,
    g406_p_spl_,
    g415_p_spl_
  );


  and

  (
    g417_p,
    g368_n_spl_,
    g370_n_spl_
  );


  or

  (
    g417_n,
    g368_p_spl_,
    g370_p_spl_
  );


  and

  (
    g418_p,
    g371_n_spl_,
    g417_n
  );


  or

  (
    g418_n,
    g371_p_spl_,
    g417_p
  );


  and

  (
    g419_p,
    g416_n_spl_,
    g418_p_spl_
  );


  or

  (
    g419_n,
    g416_p_spl_,
    g418_n_spl_
  );


  and

  (
    g420_p,
    g416_p_spl_,
    g418_n_spl_
  );


  or

  (
    g420_n,
    g416_n_spl_,
    g418_p_spl_
  );


  and

  (
    g421_p,
    g419_n_spl_,
    g420_n
  );


  or

  (
    g421_n,
    g419_p_spl_,
    g420_p
  );


  and

  (
    g422_p,
    g408_p_spl_0,
    g421_p_spl_
  );


  or

  (
    g422_n,
    g408_n_spl_0,
    g421_n_spl_
  );


  and

  (
    g423_p,
    g419_n_spl_,
    g422_n_spl_
  );


  or

  (
    g423_n,
    g419_p_spl_,
    g422_p_spl_
  );


  and

  (
    g424_p,
    g380_n_spl_,
    g382_n_spl_
  );


  or

  (
    g424_n,
    g380_p_spl_,
    g382_p_spl_
  );


  and

  (
    g425_p,
    g383_n_spl_,
    g424_n
  );


  or

  (
    g425_n,
    g383_p_spl_,
    g424_p
  );


  and

  (
    g426_p,
    g423_n_spl_,
    g425_p_spl_
  );


  or

  (
    g426_n,
    g423_p_spl_,
    g425_n_spl_
  );


  and

  (
    g427_p,
    g378_n_spl_,
    g389_n_spl_
  );


  or

  (
    g427_n,
    g378_p_spl_,
    g389_p_spl_
  );


  and

  (
    g428_p,
    g390_n_spl_,
    g427_n
  );


  or

  (
    g428_n,
    g390_p_spl_,
    g427_p
  );


  and

  (
    g429_p,
    g426_p_spl_0,
    g428_p_spl_
  );


  or

  (
    g429_n,
    g426_n_spl_0,
    g428_n_spl_
  );


  and

  (
    g430_p,
    input_f[1]_p_spl_11,
    input_w[1]_p_spl_11
  );


  or

  (
    g430_n,
    input_f[1]_n_spl_11,
    input_w[1]_n_spl_11
  );


  and

  (
    g431_p,
    g395_p_spl_0,
    g430_p_spl_0
  );


  or

  (
    g431_n,
    g395_n_spl_0,
    g430_n_spl_0
  );


  and

  (
    g432_p,
    input_f[0]_p_spl_10,
    input_w[2]_p_spl_11
  );


  or

  (
    g432_n,
    input_f[0]_n_spl_10,
    input_w[2]_n_spl_11
  );


  and

  (
    g433_p,
    g395_n_spl_,
    g430_n_spl_0
  );


  or

  (
    g433_n,
    g395_p_spl_,
    g430_p_spl_0
  );


  and

  (
    g434_p,
    g431_n_spl_,
    g433_n
  );


  or

  (
    g434_n,
    g431_p_spl_,
    g433_p
  );


  and

  (
    g435_p,
    g432_p_spl_,
    g434_p_spl_
  );


  or

  (
    g435_n,
    g432_n_spl_,
    g434_n_spl_
  );


  and

  (
    g436_p,
    g431_n_spl_,
    g435_n_spl_
  );


  or

  (
    g436_n,
    g431_p_spl_,
    g435_p_spl_
  );


  and

  (
    g437_p,
    g397_n_spl_,
    g401_n_spl_
  );


  or

  (
    g437_n,
    g397_p_spl_,
    g401_p_spl_
  );


  and

  (
    g438_p,
    g402_n_spl_,
    g437_n
  );


  or

  (
    g438_n,
    g402_p_spl_,
    g437_p
  );


  and

  (
    g439_p,
    g436_n_spl_,
    g438_p_spl_
  );


  or

  (
    g439_n,
    g436_p_spl_,
    g438_n_spl_
  );


  and

  (
    g440_p,
    g436_p_spl_,
    g438_n_spl_
  );


  or

  (
    g440_n,
    g436_n_spl_,
    g438_p_spl_
  );


  and

  (
    g441_p,
    g439_n_spl_,
    g440_n
  );


  or

  (
    g441_n,
    g439_p_spl_,
    g440_p
  );


  and

  (
    g442_p,
    g407_p_spl_0,
    g441_p_spl_
  );


  or

  (
    g442_n,
    g407_n_spl_0,
    g441_n_spl_
  );


  and

  (
    g443_p,
    g439_n_spl_,
    g442_n_spl_
  );


  or

  (
    g443_n,
    g439_p_spl_,
    g442_p_spl_
  );


  and

  (
    g444_p,
    g412_n_spl_,
    g414_n_spl_
  );


  or

  (
    g444_n,
    g412_p_spl_,
    g414_p_spl_
  );


  and

  (
    g445_p,
    g415_n_spl_,
    g444_n
  );


  or

  (
    g445_n,
    g415_p_spl_,
    g444_p
  );


  and

  (
    g446_p,
    g443_n_spl_,
    g445_p_spl_
  );


  or

  (
    g446_n,
    g443_p_spl_,
    g445_n_spl_
  );


  and

  (
    g447_p,
    g408_n_spl_,
    g421_n_spl_
  );


  or

  (
    g447_n,
    g408_p_spl_,
    g421_p_spl_
  );


  and

  (
    g448_p,
    g422_n_spl_,
    g447_n
  );


  or

  (
    g448_n,
    g422_p_spl_,
    g447_p
  );


  and

  (
    g449_p,
    g446_p_spl_0,
    g448_p_spl_
  );


  or

  (
    g449_n,
    g446_n_spl_0,
    g448_n_spl_
  );


  and

  (
    g450_p,
    g423_p_spl_,
    g425_n_spl_
  );


  or

  (
    g450_n,
    g423_n_spl_,
    g425_p_spl_
  );


  and

  (
    g451_p,
    g426_n_spl_0,
    g450_n
  );


  or

  (
    g451_n,
    g426_p_spl_0,
    g450_p
  );


  and

  (
    g452_p,
    g449_p_spl_0,
    g451_p_spl_
  );


  or

  (
    g452_n,
    g449_n_spl_0,
    g451_n_spl_
  );


  and

  (
    g453_p,
    input_f[0]_p_spl_11,
    input_w[0]_p_spl_11
  );


  or

  (
    g453_n,
    input_f[0]_n_spl_11,
    input_w[0]_n_spl_11
  );


  and

  (
    g454_p,
    g430_p_spl_,
    g453_p_spl_
  );


  or

  (
    g454_n,
    g430_n_spl_,
    g453_n_spl_
  );


  and

  (
    g455_p,
    g432_n_spl_,
    g434_n_spl_
  );


  or

  (
    g455_n,
    g432_p_spl_,
    g434_p_spl_
  );


  and

  (
    g456_p,
    g435_n_spl_,
    g455_n
  );


  or

  (
    g456_n,
    g435_p_spl_,
    g455_p
  );


  and

  (
    g457_p,
    g454_p_spl_0,
    g456_p_spl_
  );


  or

  (
    g457_n,
    g454_n_spl_0,
    g456_n_spl_
  );


  and

  (
    g458_p,
    g407_n_spl_,
    g441_n_spl_
  );


  or

  (
    g458_n,
    g407_p_spl_,
    g441_p_spl_
  );


  and

  (
    g459_p,
    g442_n_spl_,
    g458_n
  );


  or

  (
    g459_n,
    g442_p_spl_,
    g458_p
  );


  and

  (
    g460_p,
    g457_p_spl_0,
    g459_p_spl_
  );


  or

  (
    g460_n,
    g457_n_spl_0,
    g459_n_spl_
  );


  and

  (
    g461_p,
    g443_p_spl_,
    g445_n_spl_
  );


  or

  (
    g461_n,
    g443_n_spl_,
    g445_p_spl_
  );


  and

  (
    g462_p,
    g446_n_spl_0,
    g461_n
  );


  or

  (
    g462_n,
    g446_p_spl_0,
    g461_p
  );


  and

  (
    g463_p,
    g460_p_spl_0,
    g462_p_spl_
  );


  or

  (
    g463_n,
    g460_n_spl_0,
    g462_n_spl_
  );


  and

  (
    g464_p,
    g446_n_spl_,
    g448_n_spl_
  );


  or

  (
    g464_n,
    g446_p_spl_,
    g448_p_spl_
  );


  and

  (
    g465_p,
    g449_n_spl_0,
    g464_n
  );


  or

  (
    g465_n,
    g449_p_spl_0,
    g464_p
  );


  and

  (
    g466_p,
    g463_p_spl_0,
    g465_p_spl_
  );


  or

  (
    g466_n,
    g463_n_spl_0,
    g465_n_spl_
  );


  and

  (
    g467_p,
    g449_n_spl_,
    g451_n_spl_
  );


  or

  (
    g467_n,
    g449_p_spl_,
    g451_p_spl_
  );


  and

  (
    g468_p,
    g452_n_spl_,
    g467_n
  );


  or

  (
    g468_n,
    g452_p_spl_,
    g467_p
  );


  and

  (
    g469_p,
    g466_p_spl_0,
    g468_p_spl_
  );


  or

  (
    g469_n,
    g466_n_spl_0,
    g468_n_spl_
  );


  and

  (
    g470_p,
    g452_n_spl_,
    g469_n_spl_
  );


  or

  (
    g470_n,
    g452_p_spl_,
    g469_p_spl_
  );


  and

  (
    g471_p,
    g426_n_spl_,
    g428_n_spl_
  );


  or

  (
    g471_n,
    g426_p_spl_,
    g428_p_spl_
  );


  and

  (
    g472_p,
    g429_n_spl_,
    g471_n
  );


  or

  (
    g472_n,
    g429_p_spl_,
    g471_p
  );


  and

  (
    g473_p,
    g470_n_spl_,
    g472_p_spl_
  );


  or

  (
    g473_n,
    g470_p_spl_,
    g472_n_spl_
  );


  and

  (
    g474_p,
    g429_n_spl_,
    g473_n_spl_
  );


  or

  (
    g474_n,
    g429_p_spl_,
    g473_p_spl_
  );


  and

  (
    g475_p,
    g391_p_spl_,
    g393_n_spl_
  );


  or

  (
    g475_n,
    g391_n_spl_,
    g393_p_spl_
  );


  and

  (
    g476_p,
    g394_n_spl_,
    g475_n
  );


  or

  (
    g476_n,
    g394_p_spl_,
    g475_p
  );


  and

  (
    g477_p,
    g474_n_spl_,
    g476_p_spl_
  );


  or

  (
    g477_n,
    g474_p_spl_,
    g476_n_spl_
  );


  and

  (
    g478_p,
    g394_n_spl_,
    g477_n_spl_
  );


  or

  (
    g478_n,
    g394_p_spl_,
    g477_p_spl_
  );


  and

  (
    g479_p,
    g346_p_spl_,
    g348_n_spl_
  );


  or

  (
    g479_n,
    g346_n_spl_,
    g348_p_spl_
  );


  and

  (
    g480_p,
    g349_n_spl_,
    g479_n
  );


  or

  (
    g480_n,
    g349_p_spl_,
    g479_p
  );


  and

  (
    g481_p,
    g478_n_spl_,
    g480_p_spl_
  );


  or

  (
    g481_n,
    g478_p_spl_,
    g480_n_spl_
  );


  and

  (
    g482_p,
    g349_n_spl_,
    g481_n_spl_
  );


  or

  (
    g482_n,
    g349_p_spl_,
    g481_p_spl_
  );


  and

  (
    g483_p,
    g303_p_spl_,
    g482_n_spl_
  );


  or

  (
    g483_n,
    g303_n_spl_,
    g482_p_spl_
  );


  and

  (
    g484_p,
    g301_n_spl_,
    g483_n_spl_
  );


  or

  (
    g484_n,
    g301_p_spl_,
    g483_p_spl_
  );


  and

  (
    g485_p,
    g240_p_spl_,
    g484_n_spl_
  );


  or

  (
    g485_n,
    g240_n_spl_,
    g484_p_spl_
  );


  and

  (
    g486_p,
    g238_n_spl_,
    g485_n_spl_
  );


  or

  (
    g486_n,
    g238_p_spl_,
    g485_p_spl_
  );


  and

  (
    g487_p,
    g182_p_spl_,
    g184_n_spl_
  );


  or

  (
    g487_n,
    g182_n_spl_,
    g184_p_spl_
  );


  and

  (
    g488_p,
    g185_n_spl_,
    g487_n
  );


  or

  (
    g488_n,
    g185_p_spl_,
    g487_p
  );


  and

  (
    g489_p,
    g486_n_spl_,
    g488_p_spl_
  );


  or

  (
    g489_n,
    g486_p_spl_,
    g488_n_spl_
  );


  and

  (
    g490_p,
    g185_n_spl_,
    g489_n_spl_
  );


  or

  (
    g490_n,
    g185_p_spl_,
    g489_p_spl_
  );


  and

  (
    g491_p,
    g110_p_spl_,
    g136_n_spl_
  );


  or

  (
    g491_n,
    g110_n_spl_,
    g136_p_spl_
  );


  and

  (
    g492_p,
    g137_n_spl_,
    g491_n
  );


  or

  (
    g492_n,
    g137_p_spl_,
    g491_p
  );


  and

  (
    g493_p,
    g490_n_spl_,
    g492_p_spl_
  );


  or

  (
    g493_n,
    g490_p_spl_,
    g492_n_spl_
  );


  and

  (
    g494_p,
    g137_n_spl_,
    g493_n_spl_
  );


  or

  (
    g494_n,
    g137_p_spl_,
    g493_p_spl_
  );


  and

  (
    g495_p,
    g131_n_spl_,
    g134_n_spl_
  );


  or

  (
    g495_n,
    g131_p_spl_,
    g134_p_spl_
  );


  and

  (
    g496_p,
    g122_n_spl_,
    g125_n_spl_
  );


  or

  (
    g496_n,
    g122_p_spl_,
    g125_p_spl_
  );


  and

  (
    g497_p,
    input_f[7]_n_spl_11,
    input_w[7]_p_spl_11
  );


  or

  (
    g497_n,
    input_f[7]_p_spl_11,
    input_w[7]_n_spl_11
  );


  and

  (
    g498_p,
    g119_n_spl_,
    g497_n
  );


  or

  (
    g498_n,
    g119_p_spl_,
    g497_p
  );


  and

  (
    g499_p,
    g116_p_spl_1,
    g498_p_spl_
  );


  or

  (
    g499_n,
    g116_n_spl_1,
    g498_n_spl_
  );


  and

  (
    g500_p,
    g116_n_spl_1,
    g498_n_spl_
  );


  or

  (
    g500_n,
    g116_p_spl_1,
    g498_p_spl_
  );


  and

  (
    g501_p,
    g499_n_spl_0,
    g500_n
  );


  or

  (
    g501_n,
    g499_p_spl_0,
    g500_p
  );


  and

  (
    g502_p,
    g115_p_spl_1,
    g501_n_spl_
  );


  or

  (
    g502_n,
    g115_n_spl_1,
    g501_p_spl_
  );


  and

  (
    g503_p,
    g115_n_spl_1,
    g501_p_spl_
  );


  or

  (
    g503_n,
    g115_p_spl_1,
    g501_n_spl_
  );


  and

  (
    g504_p,
    g502_n_spl_,
    g503_n
  );


  or

  (
    g504_n,
    g502_p_spl_,
    g503_p
  );


  and

  (
    g505_p,
    g113_n_spl_0,
    g128_n_spl_
  );


  or

  (
    g505_n,
    g113_p_spl_0,
    g128_p_spl_
  );


  and

  (
    g506_p,
    g504_n_spl_,
    g505_n_spl_
  );


  or

  (
    g506_n,
    g504_p_spl_,
    g505_p_spl_
  );


  and

  (
    g507_p,
    g504_p_spl_,
    g505_p_spl_
  );


  or

  (
    g507_n,
    g504_n_spl_,
    g505_n_spl_
  );


  and

  (
    g508_p,
    g506_n_spl_,
    g507_n
  );


  or

  (
    g508_n,
    g506_p_spl_,
    g507_p
  );


  and

  (
    g509_p,
    g496_n_spl_,
    g508_p_spl_
  );


  or

  (
    g509_n,
    g496_p_spl_,
    g508_n_spl_
  );


  and

  (
    g510_p,
    g496_p_spl_,
    g508_n_spl_
  );


  or

  (
    g510_n,
    g496_n_spl_,
    g508_p_spl_
  );


  and

  (
    g511_p,
    g509_n_spl_,
    g510_n
  );


  or

  (
    g511_n,
    g509_p_spl_,
    g510_p
  );


  and

  (
    g512_p,
    g495_n_spl_,
    g511_p_spl_
  );


  or

  (
    g512_n,
    g495_p_spl_,
    g511_n_spl_
  );


  and

  (
    g513_p,
    g495_p_spl_,
    g511_n_spl_
  );


  or

  (
    g513_n,
    g495_n_spl_,
    g511_p_spl_
  );


  and

  (
    g514_p,
    g512_n_spl_,
    g513_n
  );


  or

  (
    g514_n,
    g512_p_spl_,
    g513_p
  );


  and

  (
    g515_p,
    g494_n_spl_,
    g514_p_spl_
  );


  or

  (
    g515_n,
    g494_p_spl_,
    g514_n_spl_
  );


  and

  (
    g516_p,
    g113_n_spl_,
    g502_n_spl_
  );


  or

  (
    g516_n,
    g113_p_spl_,
    g502_p_spl_
  );


  and

  (
    g517_p,
    g499_p_spl_0,
    g516_p_spl_
  );


  or

  (
    g517_n,
    g499_n_spl_0,
    g516_n_spl_
  );


  and

  (
    g518_p,
    g499_n_spl_,
    g516_n_spl_
  );


  or

  (
    g518_n,
    g499_p_spl_,
    g516_p_spl_
  );


  and

  (
    g519_p,
    g506_n_spl_,
    g509_n_spl_
  );


  or

  (
    g519_n,
    g506_p_spl_,
    g509_p_spl_
  );


  and

  (
    g520_p,
    g518_n,
    g519_n
  );


  or

  (
    g520_n,
    g518_p,
    g519_p
  );


  and

  (
    g521_p,
    g517_n,
    g520_n
  );


  or

  (
    g521_n,
    g517_p,
    g520_p
  );


  and

  (
    g522_p,
    g512_n_spl_,
    g521_p
  );


  or

  (
    g522_n,
    g512_p_spl_,
    g521_n
  );


  and

  (
    g523_p,
    g515_n_spl_,
    g522_p
  );


  or

  (
    g523_n,
    g515_p_spl_,
    g522_n
  );


  and

  (
    g524_p,
    g490_p_spl_,
    g492_n_spl_
  );


  or

  (
    g524_n,
    g490_n_spl_,
    g492_p_spl_
  );


  and

  (
    g525_p,
    g493_n_spl_,
    g524_n
  );


  or

  (
    g525_n,
    g493_p_spl_,
    g524_p
  );


  and

  (
    g526_p,
    g494_p_spl_,
    g514_n_spl_
  );


  or

  (
    g526_n,
    g494_n_spl_,
    g514_p_spl_
  );


  and

  (
    g527_p,
    g515_n_spl_,
    g526_n
  );


  or

  (
    g527_n,
    g515_p_spl_,
    g526_p
  );


  and

  (
    g528_p,
    g486_p_spl_,
    g488_n_spl_
  );


  or

  (
    g528_n,
    g486_n_spl_,
    g488_p_spl_
  );


  and

  (
    g529_p,
    g489_n_spl_,
    g528_n
  );


  or

  (
    g529_n,
    g489_p_spl_,
    g528_p
  );


  and

  (
    g530_p,
    g303_n_spl_,
    g482_p_spl_
  );


  or

  (
    g530_n,
    g303_p_spl_,
    g482_n_spl_
  );


  and

  (
    g531_p,
    g483_n_spl_,
    g530_n
  );


  or

  (
    g531_n,
    g483_p_spl_,
    g530_p
  );


  and

  (
    g532_p,
    g470_p_spl_,
    g472_n_spl_
  );


  or

  (
    g532_n,
    g470_n_spl_,
    g472_p_spl_
  );


  and

  (
    g533_p,
    g473_n_spl_,
    g532_n
  );


  or

  (
    g533_n,
    g473_p_spl_,
    g532_p
  );


  and

  (
    g534_p,
    g474_p_spl_,
    g476_n_spl_
  );


  or

  (
    g534_n,
    g474_n_spl_,
    g476_p_spl_
  );


  and

  (
    g535_p,
    g477_n_spl_,
    g534_n
  );


  or

  (
    g535_n,
    g477_p_spl_,
    g534_p
  );


  and

  (
    g536_p,
    g533_n_spl_,
    g535_n_spl_
  );


  or

  (
    g536_n,
    g533_p_spl_,
    g535_p_spl_
  );


  and

  (
    g537_p,
    g531_n_spl_,
    g536_p
  );


  or

  (
    g537_n,
    g531_p_spl_,
    g536_n
  );


  and

  (
    g538_p,
    g529_n_spl_,
    g537_p
  );


  or

  (
    g538_n,
    g529_p_spl_,
    g537_n
  );


  and

  (
    g539_p,
    g240_n_spl_,
    g484_p_spl_
  );


  or

  (
    g539_n,
    g240_p_spl_,
    g484_n_spl_
  );


  and

  (
    g540_p,
    g485_n_spl_,
    g539_n
  );


  or

  (
    g540_n,
    g485_p_spl_,
    g539_p
  );


  and

  (
    g541_p,
    g478_p_spl_,
    g480_n_spl_
  );


  or

  (
    g541_n,
    g478_n_spl_,
    g480_p_spl_
  );


  and

  (
    g542_p,
    g481_n_spl_,
    g541_n
  );


  or

  (
    g542_n,
    g481_p_spl_,
    g541_p
  );


  and

  (
    g543_p,
    g540_n_spl_,
    g542_n_spl_
  );


  or

  (
    g543_n,
    g540_p_spl_,
    g542_p_spl_
  );


  and

  (
    g544_p,
    g538_p,
    g543_p
  );


  or

  (
    g544_n,
    g538_n,
    g543_n
  );


  and

  (
    g545_p,
    g527_n,
    g544_p
  );


  or

  (
    g545_n,
    g527_p,
    g544_n
  );


  and

  (
    g546_p,
    g525_n_spl_,
    g545_p
  );


  or

  (
    g546_n,
    g525_p_spl_,
    g545_n
  );


  and

  (
    g547_p,
    g523_n_spl_0,
    g546_n
  );


  or

  (
    g547_n,
    g523_p_spl_0,
    g546_p
  );


  and

  (
    g548_p,
    g533_p_spl_,
    g535_p_spl_
  );


  or

  (
    g548_n,
    g533_n_spl_,
    g535_n_spl_
  );


  and

  (
    g549_p,
    g531_p_spl_,
    g548_p
  );


  or

  (
    g549_n,
    g531_n_spl_,
    g548_n
  );


  and

  (
    g550_p,
    g540_p_spl_,
    g549_p
  );


  or

  (
    g550_n,
    g540_n_spl_,
    g549_n
  );


  and

  (
    g551_p,
    g529_p_spl_,
    g550_p
  );


  or

  (
    g551_n,
    g529_n_spl_,
    g550_n
  );


  and

  (
    g552_p,
    g542_p_spl_,
    g551_p
  );


  or

  (
    g552_n,
    g542_n_spl_,
    g551_n
  );


  and

  (
    g553_p,
    g525_p_spl_,
    g552_p
  );


  or

  (
    g553_n,
    g525_n_spl_,
    g552_n
  );


  and

  (
    g554_p,
    g523_p_spl_0,
    g553_n
  );


  or

  (
    g554_n,
    g523_n_spl_0,
    g553_p
  );


  and

  (
    g555_p,
    g466_n_spl_0,
    g468_n_spl_
  );


  or

  (
    g555_n,
    g466_p_spl_0,
    g468_p_spl_
  );


  and

  (
    g556_p,
    g554_n_spl_00,
    g555_n
  );


  or

  (
    g556_n,
    g554_p_spl_00,
    g555_p
  );


  and

  (
    g557_p,
    g469_n_spl_,
    g556_p
  );


  or

  (
    g557_n,
    g469_p_spl_,
    g556_n
  );


  and

  (
    g558_p,
    g547_n_spl_00,
    g557_n
  );


  or

  (
    g558_n,
    g547_p_spl_00,
    g557_p
  );


  and

  (
    g559_p,
    reset_n_spl_00,
    psum_reg[6]_p
  );


  or

  (
    g559_n,
    reset_p_spl_00,
    psum_reg[6]_n
  );


  and

  (
    g560_p,
    g558_n_spl_,
    g559_p_spl_
  );


  or

  (
    g560_n,
    g558_p_spl_,
    g559_n_spl_0
  );


  and

  (
    g561_p,
    g463_n_spl_0,
    g465_n_spl_
  );


  or

  (
    g561_n,
    g463_p_spl_0,
    g465_p_spl_
  );


  and

  (
    g562_p,
    g554_n_spl_00,
    g561_n
  );


  or

  (
    g562_n,
    g554_p_spl_00,
    g561_p
  );


  and

  (
    g563_p,
    g466_n_spl_,
    g562_p
  );


  or

  (
    g563_n,
    g466_p_spl_,
    g562_n
  );


  and

  (
    g564_p,
    g547_n_spl_00,
    g563_n
  );


  or

  (
    g564_n,
    g547_p_spl_00,
    g563_p
  );


  and

  (
    g565_p,
    reset_n_spl_01,
    psum_reg[5]_p
  );


  or

  (
    g565_n,
    reset_p_spl_01,
    psum_reg[5]_n
  );


  and

  (
    g566_p,
    g564_n_spl_,
    g565_p_spl_
  );


  or

  (
    g566_n,
    g564_p_spl_,
    g565_n_spl_0
  );


  and

  (
    g567_p,
    g460_n_spl_0,
    g462_n_spl_
  );


  or

  (
    g567_n,
    g460_p_spl_0,
    g462_p_spl_
  );


  and

  (
    g568_p,
    g554_n_spl_01,
    g567_n
  );


  or

  (
    g568_n,
    g554_p_spl_01,
    g567_p
  );


  and

  (
    g569_p,
    g463_n_spl_,
    g568_p
  );


  or

  (
    g569_n,
    g463_p_spl_,
    g568_n
  );


  and

  (
    g570_p,
    g547_n_spl_01,
    g569_n
  );


  or

  (
    g570_n,
    g547_p_spl_01,
    g569_p
  );


  and

  (
    g571_p,
    reset_n_spl_01,
    psum_reg[4]_p
  );


  or

  (
    g571_n,
    reset_p_spl_01,
    psum_reg[4]_n
  );


  and

  (
    g572_p,
    g570_n_spl_,
    g571_p_spl_
  );


  or

  (
    g572_n,
    g570_p_spl_,
    g571_n_spl_0
  );


  and

  (
    g573_p,
    g570_p_spl_,
    g571_n_spl_0
  );


  or

  (
    g573_n,
    g570_n_spl_,
    g571_p_spl_
  );


  and

  (
    g574_p,
    g572_n_spl_,
    g573_n
  );


  or

  (
    g574_n,
    g572_p_spl_,
    g573_p
  );


  and

  (
    g575_p,
    g457_n_spl_0,
    g459_n_spl_
  );


  or

  (
    g575_n,
    g457_p_spl_0,
    g459_p_spl_
  );


  and

  (
    g576_p,
    g554_n_spl_01,
    g575_n
  );


  or

  (
    g576_n,
    g554_p_spl_01,
    g575_p
  );


  and

  (
    g577_p,
    g460_n_spl_,
    g576_p
  );


  or

  (
    g577_n,
    g460_p_spl_,
    g576_n
  );


  and

  (
    g578_p,
    g547_n_spl_01,
    g577_n
  );


  or

  (
    g578_n,
    g547_p_spl_01,
    g577_p
  );


  and

  (
    g579_p,
    reset_n_spl_10,
    psum_reg[3]_p
  );


  or

  (
    g579_n,
    reset_p_spl_10,
    psum_reg[3]_n
  );


  and

  (
    g580_p,
    g578_n_spl_,
    g579_p_spl_
  );


  or

  (
    g580_n,
    g578_p_spl_,
    g579_n_spl_0
  );


  and

  (
    g581_p,
    g578_p_spl_,
    g579_n_spl_0
  );


  or

  (
    g581_n,
    g578_n_spl_,
    g579_p_spl_
  );


  and

  (
    g582_p,
    g454_n_spl_0,
    g456_n_spl_
  );


  or

  (
    g582_n,
    g454_p_spl_0,
    g456_p_spl_
  );


  and

  (
    g583_p,
    g554_n_spl_10,
    g582_n
  );


  or

  (
    g583_n,
    g554_p_spl_10,
    g582_p
  );


  and

  (
    g584_p,
    g457_n_spl_,
    g583_p
  );


  or

  (
    g584_n,
    g457_p_spl_,
    g583_n
  );


  and

  (
    g585_p,
    g547_n_spl_10,
    g584_n
  );


  or

  (
    g585_n,
    g547_p_spl_10,
    g584_p
  );


  and

  (
    g586_p,
    reset_n_spl_10,
    psum_reg[2]_p
  );


  or

  (
    g586_n,
    reset_p_spl_10,
    psum_reg[2]_n
  );


  and

  (
    g587_p,
    g585_n_spl_,
    g586_p_spl_
  );


  or

  (
    g587_n,
    g585_p_spl_,
    g586_n_spl_0
  );


  and

  (
    g588_p,
    g585_p_spl_,
    g586_n_spl_0
  );


  or

  (
    g588_n,
    g585_n_spl_,
    g586_p_spl_
  );


  and

  (
    g589_p,
    reset_n_spl_11,
    psum_reg[1]_p
  );


  or

  (
    g589_n,
    reset_p_spl_11,
    psum_reg[1]_n
  );


  and

  (
    g590_p,
    input_f[1]_p_spl_11,
    input_w[0]_p_spl_11
  );


  or

  (
    g590_n,
    input_f[1]_n_spl_11,
    input_w[0]_n_spl_11
  );


  and

  (
    g591_p,
    input_f[0]_p_spl_11,
    input_w[1]_p_spl_11
  );


  or

  (
    g591_n,
    input_f[0]_n_spl_11,
    input_w[1]_n_spl_11
  );


  and

  (
    g592_p,
    g590_n,
    g591_n
  );


  or

  (
    g592_n,
    g590_p,
    g591_p
  );


  and

  (
    g593_p,
    g554_n_spl_10,
    g592_n
  );


  or

  (
    g593_n,
    g554_p_spl_10,
    g592_p
  );


  and

  (
    g594_p,
    g454_n_spl_,
    g593_p
  );


  or

  (
    g594_n,
    g454_p_spl_,
    g593_n
  );


  and

  (
    g595_p,
    g547_n_spl_10,
    g594_n
  );


  or

  (
    g595_n,
    g547_p_spl_10,
    g594_p
  );


  and

  (
    g596_p,
    g589_p_spl_,
    g595_n_spl_
  );


  or

  (
    g596_n,
    g589_n_spl_0,
    g595_p_spl_
  );


  and

  (
    g597_p,
    g589_n_spl_0,
    g595_p_spl_
  );


  or

  (
    g597_n,
    g589_p_spl_,
    g595_n_spl_
  );


  and

  (
    g598_p,
    reset_n_spl_11,
    psum_reg[0]_p
  );


  or

  (
    g598_n,
    reset_p_spl_11,
    psum_reg[0]_n
  );


  and

  (
    g599_p,
    g453_n_spl_,
    g547_n_spl_1
  );


  or

  (
    g599_n,
    g453_p_spl_,
    g547_p_spl_1
  );


  and

  (
    g600_p,
    g554_n_spl_1,
    g599_n
  );


  or

  (
    g600_n,
    g554_p_spl_1,
    g599_p
  );


  and

  (
    g601_p,
    g598_p,
    g600_p
  );


  or

  (
    g601_n,
    g598_n_spl_0,
    g600_n_spl_
  );


  and

  (
    g602_p,
    g597_n_spl_,
    g601_p_spl_0
  );


  or

  (
    g602_n,
    g597_p_spl_,
    g601_n_spl_
  );


  and

  (
    g603_p,
    g596_n_spl_,
    g602_n
  );


  or

  (
    g603_n,
    g596_p_spl_,
    g602_p
  );


  and

  (
    g604_p,
    g588_n_spl_,
    g603_n_spl_
  );


  or

  (
    g604_n,
    g588_p_spl_,
    g603_p_spl_
  );


  and

  (
    g605_p,
    g587_n_spl_,
    g604_n
  );


  or

  (
    g605_n,
    g587_p_spl_,
    g604_p
  );


  and

  (
    g606_p,
    g581_n_spl_,
    g605_n_spl_
  );


  or

  (
    g606_n,
    g581_p_spl_,
    g605_p_spl_
  );


  and

  (
    g607_p,
    g580_n_spl_,
    g606_n
  );


  or

  (
    g607_n,
    g580_p_spl_,
    g606_p
  );


  and

  (
    g608_p,
    g574_p,
    g607_n
  );


  or

  (
    g608_n,
    g574_n_spl_,
    g607_p_spl_
  );


  and

  (
    g609_p,
    g572_n_spl_,
    g608_n
  );


  or

  (
    g609_n,
    g572_p_spl_,
    g608_p_spl_
  );


  and

  (
    g610_p,
    g564_p_spl_,
    g565_n_spl_0
  );


  or

  (
    g610_n,
    g564_n_spl_,
    g565_p_spl_
  );


  and

  (
    g611_p,
    g566_n_spl_,
    g610_n
  );


  or

  (
    g611_n,
    g566_p_spl_,
    g610_p
  );


  and

  (
    g612_p,
    g609_n,
    g611_p
  );


  or

  (
    g612_n,
    g609_p_spl_,
    g611_n_spl_
  );


  and

  (
    g613_p,
    g566_n_spl_,
    g612_n
  );


  or

  (
    g613_n,
    g566_p_spl_,
    g612_p_spl_
  );


  and

  (
    g614_p,
    g558_p_spl_,
    g559_n_spl_0
  );


  or

  (
    g614_n,
    g558_n_spl_,
    g559_p_spl_
  );


  and

  (
    g615_p,
    g560_n_spl_,
    g614_n
  );


  or

  (
    g615_n,
    g560_p_spl_,
    g614_p
  );


  and

  (
    g616_p,
    g613_n,
    g615_p
  );


  or

  (
    g616_n,
    g613_p_spl_,
    g615_n_spl_
  );


  and

  (
    g617_p,
    g560_n_spl_,
    g616_n
  );


  or

  (
    g617_n,
    g560_p_spl_,
    g616_p_spl_
  );


  and

  (
    g618_p,
    g27_n_spl_,
    g523_n_spl_1
  );


  or

  (
    g618_n,
    g27_p_spl_0,
    g523_p_spl_1
  );


  or

  (
    g619_n,
    g617_p_spl_0,
    g618_n_spl_
  );


  and

  (
    g620_p,
    enable_p,
    g619_n
  );


  and

  (
    g621_p,
    g27_p_spl_,
    g523_p_spl_1
  );


  or

  (
    g621_n,
    g27_n_spl_,
    g523_n_spl_1
  );


  and

  (
    g622_p,
    g618_n_spl_,
    g621_n
  );


  or

  (
    g622_n,
    g618_p_spl_,
    g621_p_spl_
  );


  and

  (
    g623_p,
    g617_p_spl_0,
    g622_p_spl_
  );


  or

  (
    g623_n,
    g617_n_spl_,
    g622_n_spl_
  );


  and

  (
    g624_p,
    g617_n_spl_,
    g622_n_spl_
  );


  or

  (
    g624_n,
    g617_p_spl_,
    g622_p_spl_
  );


  and

  (
    g625_p,
    g623_n,
    g624_n
  );


  or

  (
    g625_n,
    g623_p,
    g624_p
  );


  or

  (
    g626_n,
    g621_p_spl_,
    g625_n
  );


  and

  (
    g627_p,
    g620_p_spl_00,
    g626_n_spl_
  );


  or

  (
    g628_n,
    g28_p,
    g627_p
  );


  or

  (
    g629_n,
    g618_p_spl_,
    g625_p
  );


  and

  (
    g630_p,
    g626_n_spl_,
    g629_n
  );


  and

  (
    g631_p,
    g598_n_spl_0,
    g600_n_spl_
  );


  or

  (
    g632_n,
    g601_p_spl_0,
    g631_p
  );


  or

  (
    g633_n,
    g630_p_spl_00,
    g632_n
  );


  and

  (
    g634_p,
    g620_p_spl_00,
    g633_n
  );


  and

  (
    g635_p,
    enable_n_spl_00,
    g598_n_spl_
  );


  or

  (
    g636_n,
    g634_p,
    g635_p
  );


  or

  (
    g637_n,
    g628_n_spl_00,
    g636_n_spl_
  );


  and

  (
    g638_p,
    g596_n_spl_,
    g597_n_spl_
  );


  or

  (
    g638_n,
    g596_p_spl_,
    g597_p_spl_
  );


  and

  (
    g639_p,
    g601_p_spl_,
    g638_p
  );


  and

  (
    g640_p,
    g601_n_spl_,
    g638_n
  );


  or

  (
    g641_n,
    g639_p,
    g640_p
  );


  or

  (
    g642_n,
    g630_p_spl_00,
    g641_n
  );


  and

  (
    g643_p,
    g620_p_spl_01,
    g642_n
  );


  and

  (
    g644_p,
    enable_n_spl_01,
    g589_n_spl_
  );


  or

  (
    g645_n,
    g643_p,
    g644_p
  );


  or

  (
    g646_n,
    g628_n_spl_00,
    g645_n_spl_
  );


  and

  (
    g647_p,
    g587_n_spl_,
    g588_n_spl_
  );


  or

  (
    g647_n,
    g587_p_spl_,
    g588_p_spl_
  );


  or

  (
    g648_n,
    g603_n_spl_,
    g647_n
  );


  or

  (
    g649_n,
    g603_p_spl_,
    g647_p
  );


  and

  (
    g650_p,
    g648_n,
    g649_n
  );


  or

  (
    g651_n,
    g630_p_spl_01,
    g650_p
  );


  and

  (
    g652_p,
    g620_p_spl_01,
    g651_n
  );


  and

  (
    g653_p,
    enable_n_spl_01,
    g586_n_spl_
  );


  or

  (
    g654_n,
    g652_p,
    g653_p
  );


  or

  (
    g655_n,
    g628_n_spl_01,
    g654_n_spl_
  );


  and

  (
    g656_p,
    g580_n_spl_,
    g581_n_spl_
  );


  or

  (
    g656_n,
    g580_p_spl_,
    g581_p_spl_
  );


  or

  (
    g657_n,
    g605_n_spl_,
    g656_n
  );


  or

  (
    g658_n,
    g605_p_spl_,
    g656_p
  );


  and

  (
    g659_p,
    g657_n,
    g658_n
  );


  or

  (
    g660_n,
    g630_p_spl_01,
    g659_p
  );


  and

  (
    g661_p,
    g620_p_spl_10,
    g660_n
  );


  and

  (
    g662_p,
    enable_n_spl_10,
    g579_n_spl_
  );


  or

  (
    g663_n,
    g661_p,
    g662_p
  );


  or

  (
    g664_n,
    g628_n_spl_01,
    g663_n_spl_
  );


  and

  (
    g665_p,
    g574_n_spl_,
    g607_p_spl_
  );


  or

  (
    g666_n,
    g608_p_spl_,
    g665_p
  );


  or

  (
    g667_n,
    g630_p_spl_10,
    g666_n
  );


  and

  (
    g668_p,
    g620_p_spl_10,
    g667_n
  );


  and

  (
    g669_p,
    enable_n_spl_10,
    g571_n_spl_
  );


  or

  (
    g670_n,
    g668_p,
    g669_p
  );


  or

  (
    g671_n,
    g628_n_spl_10,
    g670_n_spl_
  );


  and

  (
    g672_p,
    enable_n_spl_11,
    g565_n_spl_
  );


  and

  (
    g673_p,
    g609_p_spl_,
    g611_n_spl_
  );


  or

  (
    g674_n,
    g630_p_spl_10,
    g673_p
  );


  or

  (
    g675_n,
    g612_p_spl_,
    g674_n
  );


  and

  (
    g676_p,
    g620_p_spl_11,
    g675_n
  );


  or

  (
    g677_n,
    g672_p,
    g676_p
  );


  or

  (
    g678_n,
    g628_n_spl_10,
    g677_n_spl_
  );


  and

  (
    g679_p,
    enable_n_spl_11,
    g559_n_spl_
  );


  and

  (
    g680_p,
    g613_p_spl_,
    g615_n_spl_
  );


  or

  (
    g681_n,
    g630_p_spl_1,
    g680_p
  );


  or

  (
    g682_n,
    g616_p_spl_,
    g681_n
  );


  and

  (
    g683_p,
    g620_p_spl_11,
    g682_n
  );


  or

  (
    g684_n,
    g679_p,
    g683_p
  );


  or

  (
    g685_n,
    g628_n_spl_11,
    g684_n_spl_
  );


  not

  (
    output_f[0],
    g637_n
  );


  not

  (
    output_f[1],
    g646_n
  );


  not

  (
    output_f[2],
    g655_n
  );


  not

  (
    output_f[3],
    g664_n
  );


  not

  (
    output_f[4],
    g671_n
  );


  not

  (
    output_f[5],
    g678_n
  );


  not

  (
    output_f[6],
    g685_n
  );


  buf

  (
    output_f[7],
    1'b0
  );


  not

  (
    psum_next[0],
    g636_n_spl_
  );


  not

  (
    psum_next[1],
    g645_n_spl_
  );


  not

  (
    psum_next[2],
    g654_n_spl_
  );


  not

  (
    psum_next[3],
    g663_n_spl_
  );


  not

  (
    psum_next[4],
    g670_n_spl_
  );


  not

  (
    psum_next[5],
    g677_n_spl_
  );


  not

  (
    psum_next[6],
    g684_n_spl_
  );


  buf

  (
    psum_next[7],
    g628_n_spl_11
  );


  buf

  (
    reset_n_spl_,
    reset_n
  );


  buf

  (
    reset_n_spl_0,
    reset_n_spl_
  );


  buf

  (
    reset_n_spl_00,
    reset_n_spl_0
  );


  buf

  (
    reset_n_spl_01,
    reset_n_spl_0
  );


  buf

  (
    reset_n_spl_1,
    reset_n_spl_
  );


  buf

  (
    reset_n_spl_10,
    reset_n_spl_1
  );


  buf

  (
    reset_n_spl_11,
    reset_n_spl_1
  );


  buf

  (
    reset_p_spl_,
    reset_p
  );


  buf

  (
    reset_p_spl_0,
    reset_p_spl_
  );


  buf

  (
    reset_p_spl_00,
    reset_p_spl_0
  );


  buf

  (
    reset_p_spl_01,
    reset_p_spl_0
  );


  buf

  (
    reset_p_spl_1,
    reset_p_spl_
  );


  buf

  (
    reset_p_spl_10,
    reset_p_spl_1
  );


  buf

  (
    reset_p_spl_11,
    reset_p_spl_1
  );


  buf

  (
    enable_n_spl_,
    enable_n
  );


  buf

  (
    enable_n_spl_0,
    enable_n_spl_
  );


  buf

  (
    enable_n_spl_00,
    enable_n_spl_0
  );


  buf

  (
    enable_n_spl_01,
    enable_n_spl_0
  );


  buf

  (
    enable_n_spl_1,
    enable_n_spl_
  );


  buf

  (
    enable_n_spl_10,
    enable_n_spl_1
  );


  buf

  (
    enable_n_spl_11,
    enable_n_spl_1
  );


  buf

  (
    g27_p_spl_,
    g27_p
  );


  buf

  (
    g27_p_spl_0,
    g27_p_spl_
  );


  buf

  (
    input_f[7]_p_spl_,
    input_f[7]_p
  );


  buf

  (
    input_f[7]_p_spl_0,
    input_f[7]_p_spl_
  );


  buf

  (
    input_f[7]_p_spl_00,
    input_f[7]_p_spl_0
  );


  buf

  (
    input_f[7]_p_spl_01,
    input_f[7]_p_spl_0
  );


  buf

  (
    input_f[7]_p_spl_1,
    input_f[7]_p_spl_
  );


  buf

  (
    input_f[7]_p_spl_10,
    input_f[7]_p_spl_1
  );


  buf

  (
    input_f[7]_p_spl_11,
    input_f[7]_p_spl_1
  );


  buf

  (
    input_w[0]_p_spl_,
    input_w[0]_p
  );


  buf

  (
    input_w[0]_p_spl_0,
    input_w[0]_p_spl_
  );


  buf

  (
    input_w[0]_p_spl_00,
    input_w[0]_p_spl_0
  );


  buf

  (
    input_w[0]_p_spl_000,
    input_w[0]_p_spl_00
  );


  buf

  (
    input_w[0]_p_spl_01,
    input_w[0]_p_spl_0
  );


  buf

  (
    input_w[0]_p_spl_1,
    input_w[0]_p_spl_
  );


  buf

  (
    input_w[0]_p_spl_10,
    input_w[0]_p_spl_1
  );


  buf

  (
    input_w[0]_p_spl_11,
    input_w[0]_p_spl_1
  );


  buf

  (
    input_f[7]_n_spl_,
    input_f[7]_n
  );


  buf

  (
    input_f[7]_n_spl_0,
    input_f[7]_n_spl_
  );


  buf

  (
    input_f[7]_n_spl_00,
    input_f[7]_n_spl_0
  );


  buf

  (
    input_f[7]_n_spl_01,
    input_f[7]_n_spl_0
  );


  buf

  (
    input_f[7]_n_spl_1,
    input_f[7]_n_spl_
  );


  buf

  (
    input_f[7]_n_spl_10,
    input_f[7]_n_spl_1
  );


  buf

  (
    input_f[7]_n_spl_11,
    input_f[7]_n_spl_1
  );


  buf

  (
    input_w[0]_n_spl_,
    input_w[0]_n
  );


  buf

  (
    input_w[0]_n_spl_0,
    input_w[0]_n_spl_
  );


  buf

  (
    input_w[0]_n_spl_00,
    input_w[0]_n_spl_0
  );


  buf

  (
    input_w[0]_n_spl_000,
    input_w[0]_n_spl_00
  );


  buf

  (
    input_w[0]_n_spl_01,
    input_w[0]_n_spl_0
  );


  buf

  (
    input_w[0]_n_spl_1,
    input_w[0]_n_spl_
  );


  buf

  (
    input_w[0]_n_spl_10,
    input_w[0]_n_spl_1
  );


  buf

  (
    input_w[0]_n_spl_11,
    input_w[0]_n_spl_1
  );


  buf

  (
    input_w[1]_p_spl_,
    input_w[1]_p
  );


  buf

  (
    input_w[1]_p_spl_0,
    input_w[1]_p_spl_
  );


  buf

  (
    input_w[1]_p_spl_00,
    input_w[1]_p_spl_0
  );


  buf

  (
    input_w[1]_p_spl_000,
    input_w[1]_p_spl_00
  );


  buf

  (
    input_w[1]_p_spl_01,
    input_w[1]_p_spl_0
  );


  buf

  (
    input_w[1]_p_spl_1,
    input_w[1]_p_spl_
  );


  buf

  (
    input_w[1]_p_spl_10,
    input_w[1]_p_spl_1
  );


  buf

  (
    input_w[1]_p_spl_11,
    input_w[1]_p_spl_1
  );


  buf

  (
    g29_p_spl_,
    g29_p
  );


  buf

  (
    g29_p_spl_0,
    g29_p_spl_
  );


  buf

  (
    input_w[1]_n_spl_,
    input_w[1]_n
  );


  buf

  (
    input_w[1]_n_spl_0,
    input_w[1]_n_spl_
  );


  buf

  (
    input_w[1]_n_spl_00,
    input_w[1]_n_spl_0
  );


  buf

  (
    input_w[1]_n_spl_000,
    input_w[1]_n_spl_00
  );


  buf

  (
    input_w[1]_n_spl_01,
    input_w[1]_n_spl_0
  );


  buf

  (
    input_w[1]_n_spl_1,
    input_w[1]_n_spl_
  );


  buf

  (
    input_w[1]_n_spl_10,
    input_w[1]_n_spl_1
  );


  buf

  (
    input_w[1]_n_spl_11,
    input_w[1]_n_spl_1
  );


  buf

  (
    g29_n_spl_,
    g29_n
  );


  buf

  (
    g29_n_spl_0,
    g29_n_spl_
  );


  buf

  (
    input_w[2]_p_spl_,
    input_w[2]_p
  );


  buf

  (
    input_w[2]_p_spl_0,
    input_w[2]_p_spl_
  );


  buf

  (
    input_w[2]_p_spl_00,
    input_w[2]_p_spl_0
  );


  buf

  (
    input_w[2]_p_spl_000,
    input_w[2]_p_spl_00
  );


  buf

  (
    input_w[2]_p_spl_01,
    input_w[2]_p_spl_0
  );


  buf

  (
    input_w[2]_p_spl_1,
    input_w[2]_p_spl_
  );


  buf

  (
    input_w[2]_p_spl_10,
    input_w[2]_p_spl_1
  );


  buf

  (
    input_w[2]_p_spl_11,
    input_w[2]_p_spl_1
  );


  buf

  (
    g30_p_spl_,
    g30_p
  );


  buf

  (
    g30_p_spl_0,
    g30_p_spl_
  );


  buf

  (
    input_w[2]_n_spl_,
    input_w[2]_n
  );


  buf

  (
    input_w[2]_n_spl_0,
    input_w[2]_n_spl_
  );


  buf

  (
    input_w[2]_n_spl_00,
    input_w[2]_n_spl_0
  );


  buf

  (
    input_w[2]_n_spl_000,
    input_w[2]_n_spl_00
  );


  buf

  (
    input_w[2]_n_spl_01,
    input_w[2]_n_spl_0
  );


  buf

  (
    input_w[2]_n_spl_1,
    input_w[2]_n_spl_
  );


  buf

  (
    input_w[2]_n_spl_10,
    input_w[2]_n_spl_1
  );


  buf

  (
    input_w[2]_n_spl_11,
    input_w[2]_n_spl_1
  );


  buf

  (
    g30_n_spl_,
    g30_n
  );


  buf

  (
    g30_n_spl_0,
    g30_n_spl_
  );


  buf

  (
    g32_n_spl_,
    g32_n
  );


  buf

  (
    g34_n_spl_,
    g34_n
  );


  buf

  (
    g34_n_spl_0,
    g34_n_spl_
  );


  buf

  (
    g32_p_spl_,
    g32_p
  );


  buf

  (
    g34_p_spl_,
    g34_p
  );


  buf

  (
    g34_p_spl_0,
    g34_p_spl_
  );


  buf

  (
    g31_n_spl_,
    g31_n
  );


  buf

  (
    g31_n_spl_0,
    g31_n_spl_
  );


  buf

  (
    g31_n_spl_00,
    g31_n_spl_0
  );


  buf

  (
    g31_n_spl_01,
    g31_n_spl_0
  );


  buf

  (
    g31_n_spl_1,
    g31_n_spl_
  );


  buf

  (
    g35_n_spl_,
    g35_n
  );


  buf

  (
    g35_n_spl_0,
    g35_n_spl_
  );


  buf

  (
    g31_p_spl_,
    g31_p
  );


  buf

  (
    g31_p_spl_0,
    g31_p_spl_
  );


  buf

  (
    g31_p_spl_00,
    g31_p_spl_0
  );


  buf

  (
    g31_p_spl_01,
    g31_p_spl_0
  );


  buf

  (
    g31_p_spl_1,
    g31_p_spl_
  );


  buf

  (
    g35_p_spl_,
    g35_p
  );


  buf

  (
    g35_p_spl_0,
    g35_p_spl_
  );


  buf

  (
    input_f[5]_p_spl_,
    input_f[5]_p
  );


  buf

  (
    input_f[5]_p_spl_0,
    input_f[5]_p_spl_
  );


  buf

  (
    input_f[5]_p_spl_00,
    input_f[5]_p_spl_0
  );


  buf

  (
    input_f[5]_p_spl_01,
    input_f[5]_p_spl_0
  );


  buf

  (
    input_f[5]_p_spl_1,
    input_f[5]_p_spl_
  );


  buf

  (
    input_f[5]_p_spl_10,
    input_f[5]_p_spl_1
  );


  buf

  (
    input_f[5]_p_spl_11,
    input_f[5]_p_spl_1
  );


  buf

  (
    input_w[5]_p_spl_,
    input_w[5]_p
  );


  buf

  (
    input_w[5]_p_spl_0,
    input_w[5]_p_spl_
  );


  buf

  (
    input_w[5]_p_spl_00,
    input_w[5]_p_spl_0
  );


  buf

  (
    input_w[5]_p_spl_01,
    input_w[5]_p_spl_0
  );


  buf

  (
    input_w[5]_p_spl_1,
    input_w[5]_p_spl_
  );


  buf

  (
    input_w[5]_p_spl_10,
    input_w[5]_p_spl_1
  );


  buf

  (
    input_w[5]_p_spl_11,
    input_w[5]_p_spl_1
  );


  buf

  (
    input_f[5]_n_spl_,
    input_f[5]_n
  );


  buf

  (
    input_f[5]_n_spl_0,
    input_f[5]_n_spl_
  );


  buf

  (
    input_f[5]_n_spl_00,
    input_f[5]_n_spl_0
  );


  buf

  (
    input_f[5]_n_spl_01,
    input_f[5]_n_spl_0
  );


  buf

  (
    input_f[5]_n_spl_1,
    input_f[5]_n_spl_
  );


  buf

  (
    input_f[5]_n_spl_10,
    input_f[5]_n_spl_1
  );


  buf

  (
    input_f[5]_n_spl_11,
    input_f[5]_n_spl_1
  );


  buf

  (
    input_w[5]_n_spl_,
    input_w[5]_n
  );


  buf

  (
    input_w[5]_n_spl_0,
    input_w[5]_n_spl_
  );


  buf

  (
    input_w[5]_n_spl_00,
    input_w[5]_n_spl_0
  );


  buf

  (
    input_w[5]_n_spl_01,
    input_w[5]_n_spl_0
  );


  buf

  (
    input_w[5]_n_spl_1,
    input_w[5]_n_spl_
  );


  buf

  (
    input_w[5]_n_spl_10,
    input_w[5]_n_spl_1
  );


  buf

  (
    input_w[5]_n_spl_11,
    input_w[5]_n_spl_1
  );


  buf

  (
    input_w[3]_p_spl_,
    input_w[3]_p
  );


  buf

  (
    input_w[3]_p_spl_0,
    input_w[3]_p_spl_
  );


  buf

  (
    input_w[3]_p_spl_00,
    input_w[3]_p_spl_0
  );


  buf

  (
    input_w[3]_p_spl_000,
    input_w[3]_p_spl_00
  );


  buf

  (
    input_w[3]_p_spl_01,
    input_w[3]_p_spl_0
  );


  buf

  (
    input_w[3]_p_spl_1,
    input_w[3]_p_spl_
  );


  buf

  (
    input_w[3]_p_spl_10,
    input_w[3]_p_spl_1
  );


  buf

  (
    input_w[3]_p_spl_11,
    input_w[3]_p_spl_1
  );


  buf

  (
    input_w[3]_n_spl_,
    input_w[3]_n
  );


  buf

  (
    input_w[3]_n_spl_0,
    input_w[3]_n_spl_
  );


  buf

  (
    input_w[3]_n_spl_00,
    input_w[3]_n_spl_0
  );


  buf

  (
    input_w[3]_n_spl_000,
    input_w[3]_n_spl_00
  );


  buf

  (
    input_w[3]_n_spl_01,
    input_w[3]_n_spl_0
  );


  buf

  (
    input_w[3]_n_spl_1,
    input_w[3]_n_spl_
  );


  buf

  (
    input_w[3]_n_spl_10,
    input_w[3]_n_spl_1
  );


  buf

  (
    input_w[3]_n_spl_11,
    input_w[3]_n_spl_1
  );


  buf

  (
    input_f[6]_p_spl_,
    input_f[6]_p
  );


  buf

  (
    input_f[6]_p_spl_0,
    input_f[6]_p_spl_
  );


  buf

  (
    input_f[6]_p_spl_00,
    input_f[6]_p_spl_0
  );


  buf

  (
    input_f[6]_p_spl_01,
    input_f[6]_p_spl_0
  );


  buf

  (
    input_f[6]_p_spl_1,
    input_f[6]_p_spl_
  );


  buf

  (
    input_f[6]_p_spl_10,
    input_f[6]_p_spl_1
  );


  buf

  (
    input_f[6]_p_spl_11,
    input_f[6]_p_spl_1
  );


  buf

  (
    input_w[4]_p_spl_,
    input_w[4]_p
  );


  buf

  (
    input_w[4]_p_spl_0,
    input_w[4]_p_spl_
  );


  buf

  (
    input_w[4]_p_spl_00,
    input_w[4]_p_spl_0
  );


  buf

  (
    input_w[4]_p_spl_000,
    input_w[4]_p_spl_00
  );


  buf

  (
    input_w[4]_p_spl_01,
    input_w[4]_p_spl_0
  );


  buf

  (
    input_w[4]_p_spl_1,
    input_w[4]_p_spl_
  );


  buf

  (
    input_w[4]_p_spl_10,
    input_w[4]_p_spl_1
  );


  buf

  (
    input_w[4]_p_spl_11,
    input_w[4]_p_spl_1
  );


  buf

  (
    input_f[6]_n_spl_,
    input_f[6]_n
  );


  buf

  (
    input_f[6]_n_spl_0,
    input_f[6]_n_spl_
  );


  buf

  (
    input_f[6]_n_spl_00,
    input_f[6]_n_spl_0
  );


  buf

  (
    input_f[6]_n_spl_01,
    input_f[6]_n_spl_0
  );


  buf

  (
    input_f[6]_n_spl_1,
    input_f[6]_n_spl_
  );


  buf

  (
    input_f[6]_n_spl_10,
    input_f[6]_n_spl_1
  );


  buf

  (
    input_f[6]_n_spl_11,
    input_f[6]_n_spl_1
  );


  buf

  (
    input_w[4]_n_spl_,
    input_w[4]_n
  );


  buf

  (
    input_w[4]_n_spl_0,
    input_w[4]_n_spl_
  );


  buf

  (
    input_w[4]_n_spl_00,
    input_w[4]_n_spl_0
  );


  buf

  (
    input_w[4]_n_spl_000,
    input_w[4]_n_spl_00
  );


  buf

  (
    input_w[4]_n_spl_01,
    input_w[4]_n_spl_0
  );


  buf

  (
    input_w[4]_n_spl_1,
    input_w[4]_n_spl_
  );


  buf

  (
    input_w[4]_n_spl_10,
    input_w[4]_n_spl_1
  );


  buf

  (
    input_w[4]_n_spl_11,
    input_w[4]_n_spl_1
  );


  buf

  (
    g38_p_spl_,
    g38_p
  );


  buf

  (
    g38_p_spl_0,
    g38_p_spl_
  );


  buf

  (
    g39_p_spl_,
    g39_p
  );


  buf

  (
    g39_p_spl_0,
    g39_p_spl_
  );


  buf

  (
    g38_n_spl_,
    g38_n
  );


  buf

  (
    g38_n_spl_0,
    g38_n_spl_
  );


  buf

  (
    g39_n_spl_,
    g39_n
  );


  buf

  (
    g39_n_spl_0,
    g39_n_spl_
  );


  buf

  (
    g40_n_spl_,
    g40_n
  );


  buf

  (
    g40_p_spl_,
    g40_p
  );


  buf

  (
    g37_p_spl_,
    g37_p
  );


  buf

  (
    g42_p_spl_,
    g42_p
  );


  buf

  (
    g37_n_spl_,
    g37_n
  );


  buf

  (
    g42_n_spl_,
    g42_n
  );


  buf

  (
    g43_n_spl_,
    g43_n
  );


  buf

  (
    g43_p_spl_,
    g43_p
  );


  buf

  (
    g36_p_spl_,
    g36_p
  );


  buf

  (
    g36_p_spl_0,
    g36_p_spl_
  );


  buf

  (
    g36_p_spl_00,
    g36_p_spl_0
  );


  buf

  (
    g36_p_spl_01,
    g36_p_spl_0
  );


  buf

  (
    g36_p_spl_1,
    g36_p_spl_
  );


  buf

  (
    g45_p_spl_,
    g45_p
  );


  buf

  (
    g36_n_spl_,
    g36_n
  );


  buf

  (
    g36_n_spl_0,
    g36_n_spl_
  );


  buf

  (
    g36_n_spl_00,
    g36_n_spl_0
  );


  buf

  (
    g36_n_spl_01,
    g36_n_spl_0
  );


  buf

  (
    g36_n_spl_1,
    g36_n_spl_
  );


  buf

  (
    g45_n_spl_,
    g45_n
  );


  buf

  (
    g46_n_spl_,
    g46_n
  );


  buf

  (
    g46_p_spl_,
    g46_p
  );


  buf

  (
    g49_n_spl_,
    g49_n
  );


  buf

  (
    g49_n_spl_0,
    g49_n_spl_
  );


  buf

  (
    g49_p_spl_,
    g49_p
  );


  buf

  (
    g49_p_spl_0,
    g49_p_spl_
  );


  buf

  (
    g51_p_spl_,
    g51_p
  );


  buf

  (
    g51_p_spl_0,
    g51_p_spl_
  );


  buf

  (
    g51_p_spl_1,
    g51_p_spl_
  );


  buf

  (
    g52_p_spl_,
    g52_p
  );


  buf

  (
    g51_n_spl_,
    g51_n
  );


  buf

  (
    g51_n_spl_0,
    g51_n_spl_
  );


  buf

  (
    g51_n_spl_1,
    g51_n_spl_
  );


  buf

  (
    g52_n_spl_,
    g52_n
  );


  buf

  (
    g53_n_spl_,
    g53_n
  );


  buf

  (
    g53_p_spl_,
    g53_p
  );


  buf

  (
    g55_p_spl_,
    g55_p
  );


  buf

  (
    g55_n_spl_,
    g55_n
  );


  buf

  (
    g56_n_spl_,
    g56_n
  );


  buf

  (
    g56_p_spl_,
    g56_p
  );


  buf

  (
    g47_n_spl_,
    g47_n
  );


  buf

  (
    g58_p_spl_,
    g58_p
  );


  buf

  (
    g47_p_spl_,
    g47_p
  );


  buf

  (
    g58_n_spl_,
    g58_n
  );


  buf

  (
    input_f[4]_p_spl_,
    input_f[4]_p
  );


  buf

  (
    input_f[4]_p_spl_0,
    input_f[4]_p_spl_
  );


  buf

  (
    input_f[4]_p_spl_00,
    input_f[4]_p_spl_0
  );


  buf

  (
    input_f[4]_p_spl_01,
    input_f[4]_p_spl_0
  );


  buf

  (
    input_f[4]_p_spl_1,
    input_f[4]_p_spl_
  );


  buf

  (
    input_f[4]_p_spl_10,
    input_f[4]_p_spl_1
  );


  buf

  (
    input_f[4]_p_spl_11,
    input_f[4]_p_spl_1
  );


  buf

  (
    input_w[6]_p_spl_,
    input_w[6]_p
  );


  buf

  (
    input_w[6]_p_spl_0,
    input_w[6]_p_spl_
  );


  buf

  (
    input_w[6]_p_spl_00,
    input_w[6]_p_spl_0
  );


  buf

  (
    input_w[6]_p_spl_01,
    input_w[6]_p_spl_0
  );


  buf

  (
    input_w[6]_p_spl_1,
    input_w[6]_p_spl_
  );


  buf

  (
    input_w[6]_p_spl_10,
    input_w[6]_p_spl_1
  );


  buf

  (
    input_w[6]_p_spl_11,
    input_w[6]_p_spl_1
  );


  buf

  (
    input_f[4]_n_spl_,
    input_f[4]_n
  );


  buf

  (
    input_f[4]_n_spl_0,
    input_f[4]_n_spl_
  );


  buf

  (
    input_f[4]_n_spl_00,
    input_f[4]_n_spl_0
  );


  buf

  (
    input_f[4]_n_spl_01,
    input_f[4]_n_spl_0
  );


  buf

  (
    input_f[4]_n_spl_1,
    input_f[4]_n_spl_
  );


  buf

  (
    input_f[4]_n_spl_10,
    input_f[4]_n_spl_1
  );


  buf

  (
    input_f[4]_n_spl_11,
    input_f[4]_n_spl_1
  );


  buf

  (
    input_w[6]_n_spl_,
    input_w[6]_n
  );


  buf

  (
    input_w[6]_n_spl_0,
    input_w[6]_n_spl_
  );


  buf

  (
    input_w[6]_n_spl_00,
    input_w[6]_n_spl_0
  );


  buf

  (
    input_w[6]_n_spl_01,
    input_w[6]_n_spl_0
  );


  buf

  (
    input_w[6]_n_spl_1,
    input_w[6]_n_spl_
  );


  buf

  (
    input_w[6]_n_spl_10,
    input_w[6]_n_spl_1
  );


  buf

  (
    input_w[6]_n_spl_11,
    input_w[6]_n_spl_1
  );


  buf

  (
    input_f[3]_n_spl_,
    input_f[3]_n
  );


  buf

  (
    input_f[3]_n_spl_0,
    input_f[3]_n_spl_
  );


  buf

  (
    input_f[3]_n_spl_00,
    input_f[3]_n_spl_0
  );


  buf

  (
    input_f[3]_n_spl_01,
    input_f[3]_n_spl_0
  );


  buf

  (
    input_f[3]_n_spl_1,
    input_f[3]_n_spl_
  );


  buf

  (
    input_f[3]_n_spl_10,
    input_f[3]_n_spl_1
  );


  buf

  (
    input_f[3]_n_spl_11,
    input_f[3]_n_spl_1
  );


  buf

  (
    input_w[7]_p_spl_,
    input_w[7]_p
  );


  buf

  (
    input_w[7]_p_spl_0,
    input_w[7]_p_spl_
  );


  buf

  (
    input_w[7]_p_spl_00,
    input_w[7]_p_spl_0
  );


  buf

  (
    input_w[7]_p_spl_000,
    input_w[7]_p_spl_00
  );


  buf

  (
    input_w[7]_p_spl_001,
    input_w[7]_p_spl_00
  );


  buf

  (
    input_w[7]_p_spl_01,
    input_w[7]_p_spl_0
  );


  buf

  (
    input_w[7]_p_spl_1,
    input_w[7]_p_spl_
  );


  buf

  (
    input_w[7]_p_spl_10,
    input_w[7]_p_spl_1
  );


  buf

  (
    input_w[7]_p_spl_11,
    input_w[7]_p_spl_1
  );


  buf

  (
    input_f[3]_p_spl_,
    input_f[3]_p
  );


  buf

  (
    input_f[3]_p_spl_0,
    input_f[3]_p_spl_
  );


  buf

  (
    input_f[3]_p_spl_00,
    input_f[3]_p_spl_0
  );


  buf

  (
    input_f[3]_p_spl_01,
    input_f[3]_p_spl_0
  );


  buf

  (
    input_f[3]_p_spl_1,
    input_f[3]_p_spl_
  );


  buf

  (
    input_f[3]_p_spl_10,
    input_f[3]_p_spl_1
  );


  buf

  (
    input_f[3]_p_spl_11,
    input_f[3]_p_spl_1
  );


  buf

  (
    input_w[7]_n_spl_,
    input_w[7]_n
  );


  buf

  (
    input_w[7]_n_spl_0,
    input_w[7]_n_spl_
  );


  buf

  (
    input_w[7]_n_spl_00,
    input_w[7]_n_spl_0
  );


  buf

  (
    input_w[7]_n_spl_000,
    input_w[7]_n_spl_00
  );


  buf

  (
    input_w[7]_n_spl_001,
    input_w[7]_n_spl_00
  );


  buf

  (
    input_w[7]_n_spl_01,
    input_w[7]_n_spl_0
  );


  buf

  (
    input_w[7]_n_spl_1,
    input_w[7]_n_spl_
  );


  buf

  (
    input_w[7]_n_spl_10,
    input_w[7]_n_spl_1
  );


  buf

  (
    input_w[7]_n_spl_11,
    input_w[7]_n_spl_1
  );


  buf

  (
    g60_p_spl_,
    g60_p
  );


  buf

  (
    g61_p_spl_,
    g61_p
  );


  buf

  (
    g60_n_spl_,
    g60_n
  );


  buf

  (
    g61_n_spl_,
    g61_n
  );


  buf

  (
    g64_p_spl_,
    g64_p
  );


  buf

  (
    g65_p_spl_,
    g65_p
  );


  buf

  (
    g64_n_spl_,
    g64_n
  );


  buf

  (
    g65_n_spl_,
    g65_n
  );


  buf

  (
    g66_n_spl_,
    g66_n
  );


  buf

  (
    g66_n_spl_0,
    g66_n_spl_
  );


  buf

  (
    g66_p_spl_,
    g66_p
  );


  buf

  (
    g66_p_spl_0,
    g66_p_spl_
  );


  buf

  (
    g63_n_spl_,
    g63_n
  );


  buf

  (
    g68_p_spl_,
    g68_p
  );


  buf

  (
    g63_p_spl_,
    g63_p
  );


  buf

  (
    g68_n_spl_,
    g68_n
  );


  buf

  (
    g69_n_spl_,
    g69_n
  );


  buf

  (
    g69_p_spl_,
    g69_p
  );


  buf

  (
    g62_p_spl_,
    g62_p
  );


  buf

  (
    g62_p_spl_0,
    g62_p_spl_
  );


  buf

  (
    g71_p_spl_,
    g71_p
  );


  buf

  (
    g62_n_spl_,
    g62_n
  );


  buf

  (
    g62_n_spl_0,
    g62_n_spl_
  );


  buf

  (
    g71_n_spl_,
    g71_n
  );


  buf

  (
    g72_n_spl_,
    g72_n
  );


  buf

  (
    g72_p_spl_,
    g72_p
  );


  buf

  (
    g59_n_spl_,
    g59_n
  );


  buf

  (
    g59_p_spl_,
    g59_p
  );


  buf

  (
    g74_p_spl_,
    g74_p
  );


  buf

  (
    g76_p_spl_,
    g76_p
  );


  buf

  (
    g74_n_spl_,
    g74_n
  );


  buf

  (
    g76_n_spl_,
    g76_n
  );


  buf

  (
    g77_n_spl_,
    g77_n
  );


  buf

  (
    g77_p_spl_,
    g77_p
  );


  buf

  (
    g80_p_spl_,
    g80_p
  );


  buf

  (
    g81_p_spl_,
    g81_p
  );


  buf

  (
    g80_n_spl_,
    g80_n
  );


  buf

  (
    g81_n_spl_,
    g81_n
  );


  buf

  (
    g82_n_spl_,
    g82_n
  );


  buf

  (
    g82_n_spl_0,
    g82_n_spl_
  );


  buf

  (
    g82_p_spl_,
    g82_p
  );


  buf

  (
    g82_p_spl_0,
    g82_p_spl_
  );


  buf

  (
    g79_n_spl_,
    g79_n
  );


  buf

  (
    g84_p_spl_,
    g84_p
  );


  buf

  (
    g79_p_spl_,
    g79_p
  );


  buf

  (
    g84_n_spl_,
    g84_n
  );


  buf

  (
    g85_n_spl_,
    g85_n
  );


  buf

  (
    g85_p_spl_,
    g85_p
  );


  buf

  (
    g87_p_spl_,
    g87_p
  );


  buf

  (
    g87_n_spl_,
    g87_n
  );


  buf

  (
    g88_n_spl_,
    g88_n
  );


  buf

  (
    g88_p_spl_,
    g88_p
  );


  buf

  (
    g92_p_spl_,
    g92_p
  );


  buf

  (
    g92_n_spl_,
    g92_n
  );


  buf

  (
    g93_n_spl_,
    g93_n
  );


  buf

  (
    g93_p_spl_,
    g93_p
  );


  buf

  (
    g95_p_spl_,
    g95_p
  );


  buf

  (
    g95_p_spl_0,
    g95_p_spl_
  );


  buf

  (
    g95_p_spl_1,
    g95_p_spl_
  );


  buf

  (
    g95_n_spl_,
    g95_n
  );


  buf

  (
    g95_n_spl_0,
    g95_n_spl_
  );


  buf

  (
    g95_n_spl_1,
    g95_n_spl_
  );


  buf

  (
    g91_n_spl_,
    g91_n
  );


  buf

  (
    g98_n_spl_,
    g98_n
  );


  buf

  (
    g91_p_spl_,
    g91_p
  );


  buf

  (
    g98_p_spl_,
    g98_p
  );


  buf

  (
    g99_n_spl_,
    g99_n
  );


  buf

  (
    g99_p_spl_,
    g99_p
  );


  buf

  (
    g90_p_spl_,
    g90_p
  );


  buf

  (
    g101_p_spl_,
    g101_p
  );


  buf

  (
    g90_n_spl_,
    g90_n
  );


  buf

  (
    g101_n_spl_,
    g101_n
  );


  buf

  (
    g102_n_spl_,
    g102_n
  );


  buf

  (
    g102_p_spl_,
    g102_p
  );


  buf

  (
    g78_n_spl_,
    g78_n
  );


  buf

  (
    g104_p_spl_,
    g104_p
  );


  buf

  (
    g78_p_spl_,
    g78_p
  );


  buf

  (
    g104_n_spl_,
    g104_n
  );


  buf

  (
    g105_n_spl_,
    g105_n
  );


  buf

  (
    g105_p_spl_,
    g105_p
  );


  buf

  (
    g106_n_spl_,
    g106_n
  );


  buf

  (
    g108_p_spl_,
    g108_p
  );


  buf

  (
    g106_p_spl_,
    g106_p
  );


  buf

  (
    g108_n_spl_,
    g108_n
  );


  buf

  (
    g109_n_spl_,
    g109_n
  );


  buf

  (
    g109_p_spl_,
    g109_p
  );


  buf

  (
    g113_n_spl_,
    g113_n
  );


  buf

  (
    g113_n_spl_0,
    g113_n_spl_
  );


  buf

  (
    g113_p_spl_,
    g113_p
  );


  buf

  (
    g113_p_spl_0,
    g113_p_spl_
  );


  buf

  (
    g117_p_spl_,
    g117_p
  );


  buf

  (
    g118_n_spl_,
    g118_n
  );


  buf

  (
    g117_n_spl_,
    g117_n
  );


  buf

  (
    g118_p_spl_,
    g118_p
  );


  buf

  (
    g119_n_spl_,
    g119_n
  );


  buf

  (
    g119_p_spl_,
    g119_p
  );


  buf

  (
    g116_n_spl_,
    g116_n
  );


  buf

  (
    g116_n_spl_0,
    g116_n_spl_
  );


  buf

  (
    g116_n_spl_1,
    g116_n_spl_
  );


  buf

  (
    g121_n_spl_,
    g121_n
  );


  buf

  (
    g116_p_spl_,
    g116_p
  );


  buf

  (
    g116_p_spl_0,
    g116_p_spl_
  );


  buf

  (
    g116_p_spl_1,
    g116_p_spl_
  );


  buf

  (
    g121_p_spl_,
    g121_p
  );


  buf

  (
    g122_n_spl_,
    g122_n
  );


  buf

  (
    g122_p_spl_,
    g122_p
  );


  buf

  (
    g124_p_spl_,
    g124_p
  );


  buf

  (
    g124_n_spl_,
    g124_n
  );


  buf

  (
    g125_n_spl_,
    g125_n
  );


  buf

  (
    g125_p_spl_,
    g125_p
  );


  buf

  (
    g115_p_spl_,
    g115_p
  );


  buf

  (
    g115_p_spl_0,
    g115_p_spl_
  );


  buf

  (
    g115_p_spl_1,
    g115_p_spl_
  );


  buf

  (
    g127_p_spl_,
    g127_p
  );


  buf

  (
    g115_n_spl_,
    g115_n
  );


  buf

  (
    g115_n_spl_0,
    g115_n_spl_
  );


  buf

  (
    g115_n_spl_1,
    g115_n_spl_
  );


  buf

  (
    g127_n_spl_,
    g127_n
  );


  buf

  (
    g128_n_spl_,
    g128_n
  );


  buf

  (
    g128_p_spl_,
    g128_p
  );


  buf

  (
    g112_n_spl_,
    g112_n
  );


  buf

  (
    g130_p_spl_,
    g130_p
  );


  buf

  (
    g112_p_spl_,
    g112_p
  );


  buf

  (
    g130_n_spl_,
    g130_n
  );


  buf

  (
    g131_n_spl_,
    g131_n
  );


  buf

  (
    g131_p_spl_,
    g131_p
  );


  buf

  (
    g111_n_spl_,
    g111_n
  );


  buf

  (
    g133_p_spl_,
    g133_p
  );


  buf

  (
    g111_p_spl_,
    g111_p
  );


  buf

  (
    g133_n_spl_,
    g133_n
  );


  buf

  (
    g134_n_spl_,
    g134_n
  );


  buf

  (
    g134_p_spl_,
    g134_p
  );


  buf

  (
    g110_n_spl_,
    g110_n
  );


  buf

  (
    g136_p_spl_,
    g136_p
  );


  buf

  (
    g110_p_spl_,
    g110_p
  );


  buf

  (
    g136_n_spl_,
    g136_n
  );


  buf

  (
    g139_p_spl_,
    g139_p
  );


  buf

  (
    g139_p_spl_0,
    g139_p_spl_
  );


  buf

  (
    g139_p_spl_1,
    g139_p_spl_
  );


  buf

  (
    g139_n_spl_,
    g139_n
  );


  buf

  (
    g139_n_spl_0,
    g139_n_spl_
  );


  buf

  (
    g139_n_spl_1,
    g139_n_spl_
  );


  buf

  (
    g140_n_spl_,
    g140_n
  );


  buf

  (
    g140_p_spl_,
    g140_p
  );


  buf

  (
    g138_p_spl_,
    g138_p
  );


  buf

  (
    g144_p_spl_,
    g144_p
  );


  buf

  (
    g138_n_spl_,
    g138_n
  );


  buf

  (
    g144_n_spl_,
    g144_n
  );


  buf

  (
    g145_n_spl_,
    g145_n
  );


  buf

  (
    g145_p_spl_,
    g145_p
  );


  buf

  (
    g148_n_spl_,
    g148_n
  );


  buf

  (
    g148_n_spl_0,
    g148_n_spl_
  );


  buf

  (
    g148_p_spl_,
    g148_p
  );


  buf

  (
    g148_p_spl_0,
    g148_p_spl_
  );


  buf

  (
    g147_p_spl_,
    g147_p
  );


  buf

  (
    g153_p_spl_,
    g153_p
  );


  buf

  (
    g147_n_spl_,
    g147_n
  );


  buf

  (
    g153_n_spl_,
    g153_n
  );


  buf

  (
    g154_n_spl_,
    g154_n
  );


  buf

  (
    g154_p_spl_,
    g154_p
  );


  buf

  (
    g155_n_spl_,
    g155_n
  );


  buf

  (
    g157_p_spl_,
    g157_p
  );


  buf

  (
    g155_p_spl_,
    g155_p
  );


  buf

  (
    g157_n_spl_,
    g157_n
  );


  buf

  (
    input_f[2]_n_spl_,
    input_f[2]_n
  );


  buf

  (
    input_f[2]_n_spl_0,
    input_f[2]_n_spl_
  );


  buf

  (
    input_f[2]_n_spl_00,
    input_f[2]_n_spl_0
  );


  buf

  (
    input_f[2]_n_spl_01,
    input_f[2]_n_spl_0
  );


  buf

  (
    input_f[2]_n_spl_1,
    input_f[2]_n_spl_
  );


  buf

  (
    input_f[2]_n_spl_10,
    input_f[2]_n_spl_1
  );


  buf

  (
    input_f[2]_n_spl_11,
    input_f[2]_n_spl_1
  );


  buf

  (
    input_f[2]_p_spl_,
    input_f[2]_p
  );


  buf

  (
    input_f[2]_p_spl_0,
    input_f[2]_p_spl_
  );


  buf

  (
    input_f[2]_p_spl_00,
    input_f[2]_p_spl_0
  );


  buf

  (
    input_f[2]_p_spl_01,
    input_f[2]_p_spl_0
  );


  buf

  (
    input_f[2]_p_spl_1,
    input_f[2]_p_spl_
  );


  buf

  (
    input_f[2]_p_spl_10,
    input_f[2]_p_spl_1
  );


  buf

  (
    input_f[2]_p_spl_11,
    input_f[2]_p_spl_1
  );


  buf

  (
    g159_p_spl_,
    g159_p
  );


  buf

  (
    g160_p_spl_,
    g160_p
  );


  buf

  (
    g159_n_spl_,
    g159_n
  );


  buf

  (
    g160_n_spl_,
    g160_n
  );


  buf

  (
    g162_n_spl_,
    g162_n
  );


  buf

  (
    g164_p_spl_,
    g164_p
  );


  buf

  (
    g162_p_spl_,
    g162_p
  );


  buf

  (
    g164_n_spl_,
    g164_n
  );


  buf

  (
    g165_n_spl_,
    g165_n
  );


  buf

  (
    g165_p_spl_,
    g165_p
  );


  buf

  (
    g161_p_spl_,
    g161_p
  );


  buf

  (
    g161_p_spl_0,
    g161_p_spl_
  );


  buf

  (
    g167_p_spl_,
    g167_p
  );


  buf

  (
    g161_n_spl_,
    g161_n
  );


  buf

  (
    g161_n_spl_0,
    g161_n_spl_
  );


  buf

  (
    g167_n_spl_,
    g167_n
  );


  buf

  (
    g168_n_spl_,
    g168_n
  );


  buf

  (
    g168_p_spl_,
    g168_p
  );


  buf

  (
    g158_n_spl_,
    g158_n
  );


  buf

  (
    g158_p_spl_,
    g158_p
  );


  buf

  (
    g170_p_spl_,
    g170_p
  );


  buf

  (
    g172_p_spl_,
    g172_p
  );


  buf

  (
    g170_n_spl_,
    g170_n
  );


  buf

  (
    g172_n_spl_,
    g172_n
  );


  buf

  (
    g173_n_spl_,
    g173_n
  );


  buf

  (
    g173_p_spl_,
    g173_p
  );


  buf

  (
    g174_n_spl_,
    g174_n
  );


  buf

  (
    g176_p_spl_,
    g176_p
  );


  buf

  (
    g174_p_spl_,
    g174_p
  );


  buf

  (
    g176_n_spl_,
    g176_n
  );


  buf

  (
    g177_n_spl_,
    g177_n
  );


  buf

  (
    g177_p_spl_,
    g177_p
  );


  buf

  (
    g178_n_spl_,
    g178_n
  );


  buf

  (
    g180_p_spl_,
    g180_p
  );


  buf

  (
    g178_p_spl_,
    g178_p
  );


  buf

  (
    g180_n_spl_,
    g180_n
  );


  buf

  (
    g181_n_spl_,
    g181_n
  );


  buf

  (
    g181_p_spl_,
    g181_p
  );


  buf

  (
    g182_n_spl_,
    g182_n
  );


  buf

  (
    g184_p_spl_,
    g184_p
  );


  buf

  (
    g182_p_spl_,
    g182_p
  );


  buf

  (
    g184_n_spl_,
    g184_n
  );


  buf

  (
    g186_n_spl_,
    g186_n
  );


  buf

  (
    g186_p_spl_,
    g186_p
  );


  buf

  (
    g187_p_spl_,
    g187_p
  );


  buf

  (
    g187_p_spl_0,
    g187_p_spl_
  );


  buf

  (
    g189_p_spl_,
    g189_p
  );


  buf

  (
    g187_n_spl_,
    g187_n
  );


  buf

  (
    g187_n_spl_0,
    g187_n_spl_
  );


  buf

  (
    g189_n_spl_,
    g189_n
  );


  buf

  (
    g190_n_spl_,
    g190_n
  );


  buf

  (
    g190_p_spl_,
    g190_p
  );


  buf

  (
    g192_p_spl_,
    g192_p
  );


  buf

  (
    g192_n_spl_,
    g192_n
  );


  buf

  (
    g191_n_spl_,
    g191_n
  );


  buf

  (
    g195_n_spl_,
    g195_n
  );


  buf

  (
    g191_p_spl_,
    g191_p
  );


  buf

  (
    g195_p_spl_,
    g195_p
  );


  buf

  (
    g198_p_spl_,
    g198_p
  );


  buf

  (
    g198_n_spl_,
    g198_n
  );


  buf

  (
    g199_n_spl_,
    g199_n
  );


  buf

  (
    g199_p_spl_,
    g199_p
  );


  buf

  (
    g197_p_spl_,
    g197_p
  );


  buf

  (
    g201_p_spl_,
    g201_p
  );


  buf

  (
    g197_n_spl_,
    g197_n
  );


  buf

  (
    g201_n_spl_,
    g201_n
  );


  buf

  (
    g202_n_spl_,
    g202_n
  );


  buf

  (
    g202_p_spl_,
    g202_p
  );


  buf

  (
    g196_n_spl_,
    g196_n
  );


  buf

  (
    g196_p_spl_,
    g196_p
  );


  buf

  (
    g204_p_spl_,
    g204_p
  );


  buf

  (
    g206_p_spl_,
    g206_p
  );


  buf

  (
    g204_n_spl_,
    g204_n
  );


  buf

  (
    g206_n_spl_,
    g206_n
  );


  buf

  (
    g207_n_spl_,
    g207_n
  );


  buf

  (
    g207_p_spl_,
    g207_p
  );


  buf

  (
    g208_n_spl_,
    g208_n
  );


  buf

  (
    g210_p_spl_,
    g210_p
  );


  buf

  (
    g208_p_spl_,
    g208_p
  );


  buf

  (
    g210_n_spl_,
    g210_n
  );


  buf

  (
    input_f[1]_n_spl_,
    input_f[1]_n
  );


  buf

  (
    input_f[1]_n_spl_0,
    input_f[1]_n_spl_
  );


  buf

  (
    input_f[1]_n_spl_00,
    input_f[1]_n_spl_0
  );


  buf

  (
    input_f[1]_n_spl_01,
    input_f[1]_n_spl_0
  );


  buf

  (
    input_f[1]_n_spl_1,
    input_f[1]_n_spl_
  );


  buf

  (
    input_f[1]_n_spl_10,
    input_f[1]_n_spl_1
  );


  buf

  (
    input_f[1]_n_spl_11,
    input_f[1]_n_spl_1
  );


  buf

  (
    input_f[1]_p_spl_,
    input_f[1]_p
  );


  buf

  (
    input_f[1]_p_spl_0,
    input_f[1]_p_spl_
  );


  buf

  (
    input_f[1]_p_spl_00,
    input_f[1]_p_spl_0
  );


  buf

  (
    input_f[1]_p_spl_01,
    input_f[1]_p_spl_0
  );


  buf

  (
    input_f[1]_p_spl_1,
    input_f[1]_p_spl_
  );


  buf

  (
    input_f[1]_p_spl_10,
    input_f[1]_p_spl_1
  );


  buf

  (
    input_f[1]_p_spl_11,
    input_f[1]_p_spl_1
  );


  buf

  (
    g212_p_spl_,
    g212_p
  );


  buf

  (
    g212_p_spl_0,
    g212_p_spl_
  );


  buf

  (
    g213_p_spl_,
    g213_p
  );


  buf

  (
    g212_n_spl_,
    g212_n
  );


  buf

  (
    g212_n_spl_0,
    g212_n_spl_
  );


  buf

  (
    g213_n_spl_,
    g213_n
  );


  buf

  (
    g215_n_spl_,
    g215_n
  );


  buf

  (
    g217_p_spl_,
    g217_p
  );


  buf

  (
    g215_p_spl_,
    g215_p
  );


  buf

  (
    g217_n_spl_,
    g217_n
  );


  buf

  (
    g218_n_spl_,
    g218_n
  );


  buf

  (
    g218_p_spl_,
    g218_p
  );


  buf

  (
    g214_p_spl_,
    g214_p
  );


  buf

  (
    g214_p_spl_0,
    g214_p_spl_
  );


  buf

  (
    g220_p_spl_,
    g220_p
  );


  buf

  (
    g214_n_spl_,
    g214_n
  );


  buf

  (
    g214_n_spl_0,
    g214_n_spl_
  );


  buf

  (
    g220_n_spl_,
    g220_n
  );


  buf

  (
    g221_n_spl_,
    g221_n
  );


  buf

  (
    g221_p_spl_,
    g221_p
  );


  buf

  (
    g211_n_spl_,
    g211_n
  );


  buf

  (
    g211_p_spl_,
    g211_p
  );


  buf

  (
    g223_p_spl_,
    g223_p
  );


  buf

  (
    g225_p_spl_,
    g225_p
  );


  buf

  (
    g223_n_spl_,
    g223_n
  );


  buf

  (
    g225_n_spl_,
    g225_n
  );


  buf

  (
    g226_n_spl_,
    g226_n
  );


  buf

  (
    g226_p_spl_,
    g226_p
  );


  buf

  (
    g227_n_spl_,
    g227_n
  );


  buf

  (
    g229_p_spl_,
    g229_p
  );


  buf

  (
    g227_p_spl_,
    g227_p
  );


  buf

  (
    g229_n_spl_,
    g229_n
  );


  buf

  (
    g230_n_spl_,
    g230_n
  );


  buf

  (
    g230_p_spl_,
    g230_p
  );


  buf

  (
    g231_n_spl_,
    g231_n
  );


  buf

  (
    g233_p_spl_,
    g233_p
  );


  buf

  (
    g231_p_spl_,
    g231_p
  );


  buf

  (
    g233_n_spl_,
    g233_n
  );


  buf

  (
    g234_n_spl_,
    g234_n
  );


  buf

  (
    g234_p_spl_,
    g234_p
  );


  buf

  (
    g235_n_spl_,
    g235_n
  );


  buf

  (
    g237_p_spl_,
    g237_p
  );


  buf

  (
    g235_p_spl_,
    g235_p
  );


  buf

  (
    g237_n_spl_,
    g237_n
  );


  buf

  (
    g238_n_spl_,
    g238_n
  );


  buf

  (
    g238_p_spl_,
    g238_p
  );


  buf

  (
    g241_p_spl_,
    g241_p
  );


  buf

  (
    g241_p_spl_0,
    g241_p_spl_
  );


  buf

  (
    g241_n_spl_,
    g241_n
  );


  buf

  (
    g241_n_spl_0,
    g241_n_spl_
  );


  buf

  (
    g242_n_spl_,
    g242_n
  );


  buf

  (
    g242_p_spl_,
    g242_p
  );


  buf

  (
    g243_p_spl_,
    g243_p
  );


  buf

  (
    g243_p_spl_0,
    g243_p_spl_
  );


  buf

  (
    g247_p_spl_,
    g247_p
  );


  buf

  (
    g243_n_spl_,
    g243_n
  );


  buf

  (
    g243_n_spl_0,
    g243_n_spl_
  );


  buf

  (
    g247_n_spl_,
    g247_n
  );


  buf

  (
    g248_n_spl_,
    g248_n
  );


  buf

  (
    g248_p_spl_,
    g248_p
  );


  buf

  (
    g249_n_spl_,
    g249_n
  );


  buf

  (
    g251_p_spl_,
    g251_p
  );


  buf

  (
    g249_p_spl_,
    g249_p
  );


  buf

  (
    g251_n_spl_,
    g251_n
  );


  buf

  (
    g252_n_spl_,
    g252_n
  );


  buf

  (
    g252_p_spl_,
    g252_p
  );


  buf

  (
    g256_n_spl_,
    g256_n
  );


  buf

  (
    g256_p_spl_,
    g256_p
  );


  buf

  (
    g255_p_spl_,
    g255_p
  );


  buf

  (
    g255_p_spl_0,
    g255_p_spl_
  );


  buf

  (
    g260_p_spl_,
    g260_p
  );


  buf

  (
    g255_n_spl_,
    g255_n
  );


  buf

  (
    g255_n_spl_0,
    g255_n_spl_
  );


  buf

  (
    g260_n_spl_,
    g260_n
  );


  buf

  (
    g261_n_spl_,
    g261_n
  );


  buf

  (
    g261_p_spl_,
    g261_p
  );


  buf

  (
    g254_p_spl_,
    g254_p
  );


  buf

  (
    g263_p_spl_,
    g263_p
  );


  buf

  (
    g254_n_spl_,
    g254_n
  );


  buf

  (
    g263_n_spl_,
    g263_n
  );


  buf

  (
    g264_n_spl_,
    g264_n
  );


  buf

  (
    g264_p_spl_,
    g264_p
  );


  buf

  (
    g265_n_spl_,
    g265_n
  );


  buf

  (
    g267_p_spl_,
    g267_p
  );


  buf

  (
    g265_p_spl_,
    g265_p
  );


  buf

  (
    g267_n_spl_,
    g267_n
  );


  buf

  (
    g269_p_spl_,
    g269_p
  );


  buf

  (
    g269_p_spl_0,
    g269_p_spl_
  );


  buf

  (
    g269_n_spl_,
    g269_n
  );


  buf

  (
    g269_n_spl_0,
    g269_n_spl_
  );


  buf

  (
    input_f[0]_n_spl_,
    input_f[0]_n
  );


  buf

  (
    input_f[0]_n_spl_0,
    input_f[0]_n_spl_
  );


  buf

  (
    input_f[0]_n_spl_00,
    input_f[0]_n_spl_0
  );


  buf

  (
    input_f[0]_n_spl_01,
    input_f[0]_n_spl_0
  );


  buf

  (
    input_f[0]_n_spl_1,
    input_f[0]_n_spl_
  );


  buf

  (
    input_f[0]_n_spl_10,
    input_f[0]_n_spl_1
  );


  buf

  (
    input_f[0]_n_spl_11,
    input_f[0]_n_spl_1
  );


  buf

  (
    input_f[0]_p_spl_,
    input_f[0]_p
  );


  buf

  (
    input_f[0]_p_spl_0,
    input_f[0]_p_spl_
  );


  buf

  (
    input_f[0]_p_spl_00,
    input_f[0]_p_spl_0
  );


  buf

  (
    input_f[0]_p_spl_01,
    input_f[0]_p_spl_0
  );


  buf

  (
    input_f[0]_p_spl_1,
    input_f[0]_p_spl_
  );


  buf

  (
    input_f[0]_p_spl_10,
    input_f[0]_p_spl_1
  );


  buf

  (
    input_f[0]_p_spl_11,
    input_f[0]_p_spl_1
  );


  buf

  (
    g270_n_spl_,
    g270_n
  );


  buf

  (
    g270_p_spl_,
    g270_p
  );


  buf

  (
    g271_p_spl_,
    g271_p
  );


  buf

  (
    g275_p_spl_,
    g275_p
  );


  buf

  (
    g271_n_spl_,
    g271_n
  );


  buf

  (
    g275_n_spl_,
    g275_n
  );


  buf

  (
    g276_n_spl_,
    g276_n
  );


  buf

  (
    g276_p_spl_,
    g276_p
  );


  buf

  (
    g278_n_spl_,
    g278_n
  );


  buf

  (
    g280_p_spl_,
    g280_p
  );


  buf

  (
    g278_p_spl_,
    g278_p
  );


  buf

  (
    g280_n_spl_,
    g280_n
  );


  buf

  (
    g281_n_spl_,
    g281_n
  );


  buf

  (
    g281_p_spl_,
    g281_p
  );


  buf

  (
    g277_n_spl_,
    g277_n
  );


  buf

  (
    g283_p_spl_,
    g283_p
  );


  buf

  (
    g277_p_spl_,
    g277_p
  );


  buf

  (
    g283_n_spl_,
    g283_n
  );


  buf

  (
    g284_n_spl_,
    g284_n
  );


  buf

  (
    g284_p_spl_,
    g284_p
  );


  buf

  (
    g268_n_spl_,
    g268_n
  );


  buf

  (
    g268_p_spl_,
    g268_p
  );


  buf

  (
    g286_p_spl_,
    g286_p
  );


  buf

  (
    g288_p_spl_,
    g288_p
  );


  buf

  (
    g286_n_spl_,
    g286_n
  );


  buf

  (
    g288_n_spl_,
    g288_n
  );


  buf

  (
    g289_n_spl_,
    g289_n
  );


  buf

  (
    g289_p_spl_,
    g289_p
  );


  buf

  (
    g290_n_spl_,
    g290_n
  );


  buf

  (
    g292_p_spl_,
    g292_p
  );


  buf

  (
    g290_p_spl_,
    g290_p
  );


  buf

  (
    g292_n_spl_,
    g292_n
  );


  buf

  (
    g293_n_spl_,
    g293_n
  );


  buf

  (
    g293_p_spl_,
    g293_p
  );


  buf

  (
    g294_n_spl_,
    g294_n
  );


  buf

  (
    g296_p_spl_,
    g296_p
  );


  buf

  (
    g294_p_spl_,
    g294_p
  );


  buf

  (
    g296_n_spl_,
    g296_n
  );


  buf

  (
    g297_n_spl_,
    g297_n
  );


  buf

  (
    g297_p_spl_,
    g297_p
  );


  buf

  (
    g298_n_spl_,
    g298_n
  );


  buf

  (
    g300_p_spl_,
    g300_p
  );


  buf

  (
    g298_p_spl_,
    g298_p
  );


  buf

  (
    g300_n_spl_,
    g300_n
  );


  buf

  (
    g301_n_spl_,
    g301_n
  );


  buf

  (
    g301_p_spl_,
    g301_p
  );


  buf

  (
    g304_p_spl_,
    g304_p
  );


  buf

  (
    g304_n_spl_,
    g304_n
  );


  buf

  (
    g305_n_spl_,
    g305_n
  );


  buf

  (
    g305_p_spl_,
    g305_p
  );


  buf

  (
    g306_p_spl_,
    g306_p
  );


  buf

  (
    g308_p_spl_,
    g308_p
  );


  buf

  (
    g306_n_spl_,
    g306_n
  );


  buf

  (
    g308_n_spl_,
    g308_n
  );


  buf

  (
    g309_n_spl_,
    g309_n
  );


  buf

  (
    g309_p_spl_,
    g309_p
  );


  buf

  (
    g310_n_spl_,
    g310_n
  );


  buf

  (
    g312_p_spl_,
    g312_p
  );


  buf

  (
    g310_p_spl_,
    g310_p
  );


  buf

  (
    g312_n_spl_,
    g312_n
  );


  buf

  (
    g314_p_spl_,
    g314_p
  );


  buf

  (
    g314_p_spl_0,
    g314_p_spl_
  );


  buf

  (
    g314_n_spl_,
    g314_n
  );


  buf

  (
    g314_n_spl_0,
    g314_n_spl_
  );


  buf

  (
    g315_n_spl_,
    g315_n
  );


  buf

  (
    g315_p_spl_,
    g315_p
  );


  buf

  (
    g319_p_spl_,
    g319_p
  );


  buf

  (
    g319_n_spl_,
    g319_n
  );


  buf

  (
    g320_n_spl_,
    g320_n
  );


  buf

  (
    g320_p_spl_,
    g320_p
  );


  buf

  (
    g313_n_spl_,
    g313_n
  );


  buf

  (
    g313_p_spl_,
    g313_p
  );


  buf

  (
    g322_p_spl_,
    g322_p
  );


  buf

  (
    g324_p_spl_,
    g324_p
  );


  buf

  (
    g322_n_spl_,
    g322_n
  );


  buf

  (
    g324_n_spl_,
    g324_n
  );


  buf

  (
    g325_n_spl_,
    g325_n
  );


  buf

  (
    g325_p_spl_,
    g325_p
  );


  buf

  (
    g326_n_spl_,
    g326_n
  );


  buf

  (
    g328_p_spl_,
    g328_p
  );


  buf

  (
    g326_p_spl_,
    g326_p
  );


  buf

  (
    g328_n_spl_,
    g328_n
  );


  buf

  (
    g329_n_spl_,
    g329_n
  );


  buf

  (
    g329_p_spl_,
    g329_p
  );


  buf

  (
    g332_n_spl_,
    g332_n
  );


  buf

  (
    g334_p_spl_,
    g334_p
  );


  buf

  (
    g332_p_spl_,
    g332_p
  );


  buf

  (
    g334_n_spl_,
    g334_n
  );


  buf

  (
    g335_n_spl_,
    g335_n
  );


  buf

  (
    g335_n_spl_0,
    g335_n_spl_
  );


  buf

  (
    g335_p_spl_,
    g335_p
  );


  buf

  (
    g335_p_spl_0,
    g335_p_spl_
  );


  buf

  (
    g331_p_spl_,
    g331_p
  );


  buf

  (
    g337_p_spl_,
    g337_p
  );


  buf

  (
    g331_n_spl_,
    g331_n
  );


  buf

  (
    g337_n_spl_,
    g337_n
  );


  buf

  (
    g338_n_spl_,
    g338_n
  );


  buf

  (
    g338_p_spl_,
    g338_p
  );


  buf

  (
    g339_n_spl_,
    g339_n
  );


  buf

  (
    g341_p_spl_,
    g341_p
  );


  buf

  (
    g339_p_spl_,
    g339_p
  );


  buf

  (
    g341_n_spl_,
    g341_n
  );


  buf

  (
    g342_n_spl_,
    g342_n
  );


  buf

  (
    g342_p_spl_,
    g342_p
  );


  buf

  (
    g344_p_spl_,
    g344_p
  );


  buf

  (
    g344_n_spl_,
    g344_n
  );


  buf

  (
    g345_n_spl_,
    g345_n
  );


  buf

  (
    g345_p_spl_,
    g345_p
  );


  buf

  (
    g346_n_spl_,
    g346_n
  );


  buf

  (
    g348_p_spl_,
    g348_p
  );


  buf

  (
    g346_p_spl_,
    g346_p
  );


  buf

  (
    g348_n_spl_,
    g348_n
  );


  buf

  (
    g350_p_spl_,
    g350_p
  );


  buf

  (
    g351_p_spl_,
    g351_p
  );


  buf

  (
    g351_p_spl_0,
    g351_p_spl_
  );


  buf

  (
    g350_n_spl_,
    g350_n
  );


  buf

  (
    g351_n_spl_,
    g351_n
  );


  buf

  (
    g351_n_spl_0,
    g351_n_spl_
  );


  buf

  (
    g352_n_spl_,
    g352_n
  );


  buf

  (
    g352_p_spl_,
    g352_p
  );


  buf

  (
    g353_p_spl_,
    g353_p
  );


  buf

  (
    g355_p_spl_,
    g355_p
  );


  buf

  (
    g353_n_spl_,
    g353_n
  );


  buf

  (
    g355_n_spl_,
    g355_n
  );


  buf

  (
    g356_n_spl_,
    g356_n
  );


  buf

  (
    g356_p_spl_,
    g356_p
  );


  buf

  (
    g357_n_spl_,
    g357_n
  );


  buf

  (
    g359_p_spl_,
    g359_p
  );


  buf

  (
    g357_p_spl_,
    g357_p
  );


  buf

  (
    g359_n_spl_,
    g359_n
  );


  buf

  (
    g362_p_spl_,
    g362_p
  );


  buf

  (
    g362_p_spl_0,
    g362_p_spl_
  );


  buf

  (
    g362_n_spl_,
    g362_n
  );


  buf

  (
    g362_n_spl_0,
    g362_n_spl_
  );


  buf

  (
    g363_n_spl_,
    g363_n
  );


  buf

  (
    g363_p_spl_,
    g363_p
  );


  buf

  (
    g361_p_spl_,
    g361_p
  );


  buf

  (
    g365_p_spl_,
    g365_p
  );


  buf

  (
    g361_n_spl_,
    g361_n
  );


  buf

  (
    g365_n_spl_,
    g365_n
  );


  buf

  (
    g366_n_spl_,
    g366_n
  );


  buf

  (
    g366_p_spl_,
    g366_p
  );


  buf

  (
    g360_n_spl_,
    g360_n
  );


  buf

  (
    g360_p_spl_,
    g360_p
  );


  buf

  (
    g368_p_spl_,
    g368_p
  );


  buf

  (
    g370_p_spl_,
    g370_p
  );


  buf

  (
    g368_n_spl_,
    g368_n
  );


  buf

  (
    g370_n_spl_,
    g370_n
  );


  buf

  (
    g371_n_spl_,
    g371_n
  );


  buf

  (
    g371_p_spl_,
    g371_p
  );


  buf

  (
    g372_n_spl_,
    g372_n
  );


  buf

  (
    g374_p_spl_,
    g374_p
  );


  buf

  (
    g372_p_spl_,
    g372_p
  );


  buf

  (
    g374_n_spl_,
    g374_n
  );


  buf

  (
    g376_n_spl_,
    g376_n
  );


  buf

  (
    g377_p_spl_,
    g377_p
  );


  buf

  (
    g376_p_spl_,
    g376_p
  );


  buf

  (
    g377_n_spl_,
    g377_n
  );


  buf

  (
    g378_n_spl_,
    g378_n
  );


  buf

  (
    g378_n_spl_0,
    g378_n_spl_
  );


  buf

  (
    g378_p_spl_,
    g378_p
  );


  buf

  (
    g378_p_spl_0,
    g378_p_spl_
  );


  buf

  (
    g375_n_spl_,
    g375_n
  );


  buf

  (
    g375_p_spl_,
    g375_p
  );


  buf

  (
    g380_p_spl_,
    g380_p
  );


  buf

  (
    g382_p_spl_,
    g382_p
  );


  buf

  (
    g380_n_spl_,
    g380_n
  );


  buf

  (
    g382_n_spl_,
    g382_n
  );


  buf

  (
    g383_n_spl_,
    g383_n
  );


  buf

  (
    g383_p_spl_,
    g383_p
  );


  buf

  (
    g384_n_spl_,
    g384_n
  );


  buf

  (
    g386_p_spl_,
    g386_p
  );


  buf

  (
    g384_p_spl_,
    g384_p
  );


  buf

  (
    g386_n_spl_,
    g386_n
  );


  buf

  (
    g387_n_spl_,
    g387_n
  );


  buf

  (
    g387_p_spl_,
    g387_p
  );


  buf

  (
    g389_p_spl_,
    g389_p
  );


  buf

  (
    g389_n_spl_,
    g389_n
  );


  buf

  (
    g390_n_spl_,
    g390_n
  );


  buf

  (
    g390_p_spl_,
    g390_p
  );


  buf

  (
    g391_n_spl_,
    g391_n
  );


  buf

  (
    g393_p_spl_,
    g393_p
  );


  buf

  (
    g391_p_spl_,
    g391_p
  );


  buf

  (
    g393_n_spl_,
    g393_n
  );


  buf

  (
    g395_p_spl_,
    g395_p
  );


  buf

  (
    g395_p_spl_0,
    g395_p_spl_
  );


  buf

  (
    g395_n_spl_,
    g395_n
  );


  buf

  (
    g395_n_spl_0,
    g395_n_spl_
  );


  buf

  (
    g396_n_spl_,
    g396_n
  );


  buf

  (
    g396_p_spl_,
    g396_p
  );


  buf

  (
    g397_p_spl_,
    g397_p
  );


  buf

  (
    g401_p_spl_,
    g401_p
  );


  buf

  (
    g397_n_spl_,
    g397_n
  );


  buf

  (
    g401_n_spl_,
    g401_n
  );


  buf

  (
    g402_n_spl_,
    g402_n
  );


  buf

  (
    g402_p_spl_,
    g402_p
  );


  buf

  (
    g403_n_spl_,
    g403_n
  );


  buf

  (
    g405_p_spl_,
    g405_p
  );


  buf

  (
    g403_p_spl_,
    g403_p
  );


  buf

  (
    g405_n_spl_,
    g405_n
  );


  buf

  (
    g407_p_spl_,
    g407_p
  );


  buf

  (
    g407_p_spl_0,
    g407_p_spl_
  );


  buf

  (
    g407_n_spl_,
    g407_n
  );


  buf

  (
    g407_n_spl_0,
    g407_n_spl_
  );


  buf

  (
    g408_n_spl_,
    g408_n
  );


  buf

  (
    g408_n_spl_0,
    g408_n_spl_
  );


  buf

  (
    g408_p_spl_,
    g408_p
  );


  buf

  (
    g408_p_spl_0,
    g408_p_spl_
  );


  buf

  (
    g406_n_spl_,
    g406_n
  );


  buf

  (
    g406_p_spl_,
    g406_p
  );


  buf

  (
    g412_p_spl_,
    g412_p
  );


  buf

  (
    g414_p_spl_,
    g414_p
  );


  buf

  (
    g412_n_spl_,
    g412_n
  );


  buf

  (
    g414_n_spl_,
    g414_n
  );


  buf

  (
    g415_n_spl_,
    g415_n
  );


  buf

  (
    g415_p_spl_,
    g415_p
  );


  buf

  (
    g416_n_spl_,
    g416_n
  );


  buf

  (
    g418_p_spl_,
    g418_p
  );


  buf

  (
    g416_p_spl_,
    g416_p
  );


  buf

  (
    g418_n_spl_,
    g418_n
  );


  buf

  (
    g419_n_spl_,
    g419_n
  );


  buf

  (
    g419_p_spl_,
    g419_p
  );


  buf

  (
    g421_p_spl_,
    g421_p
  );


  buf

  (
    g421_n_spl_,
    g421_n
  );


  buf

  (
    g422_n_spl_,
    g422_n
  );


  buf

  (
    g422_p_spl_,
    g422_p
  );


  buf

  (
    g423_n_spl_,
    g423_n
  );


  buf

  (
    g425_p_spl_,
    g425_p
  );


  buf

  (
    g423_p_spl_,
    g423_p
  );


  buf

  (
    g425_n_spl_,
    g425_n
  );


  buf

  (
    g426_p_spl_,
    g426_p
  );


  buf

  (
    g426_p_spl_0,
    g426_p_spl_
  );


  buf

  (
    g428_p_spl_,
    g428_p
  );


  buf

  (
    g426_n_spl_,
    g426_n
  );


  buf

  (
    g426_n_spl_0,
    g426_n_spl_
  );


  buf

  (
    g428_n_spl_,
    g428_n
  );


  buf

  (
    g430_p_spl_,
    g430_p
  );


  buf

  (
    g430_p_spl_0,
    g430_p_spl_
  );


  buf

  (
    g430_n_spl_,
    g430_n
  );


  buf

  (
    g430_n_spl_0,
    g430_n_spl_
  );


  buf

  (
    g431_n_spl_,
    g431_n
  );


  buf

  (
    g431_p_spl_,
    g431_p
  );


  buf

  (
    g432_p_spl_,
    g432_p
  );


  buf

  (
    g434_p_spl_,
    g434_p
  );


  buf

  (
    g432_n_spl_,
    g432_n
  );


  buf

  (
    g434_n_spl_,
    g434_n
  );


  buf

  (
    g435_n_spl_,
    g435_n
  );


  buf

  (
    g435_p_spl_,
    g435_p
  );


  buf

  (
    g436_n_spl_,
    g436_n
  );


  buf

  (
    g438_p_spl_,
    g438_p
  );


  buf

  (
    g436_p_spl_,
    g436_p
  );


  buf

  (
    g438_n_spl_,
    g438_n
  );


  buf

  (
    g439_n_spl_,
    g439_n
  );


  buf

  (
    g439_p_spl_,
    g439_p
  );


  buf

  (
    g441_p_spl_,
    g441_p
  );


  buf

  (
    g441_n_spl_,
    g441_n
  );


  buf

  (
    g442_n_spl_,
    g442_n
  );


  buf

  (
    g442_p_spl_,
    g442_p
  );


  buf

  (
    g443_n_spl_,
    g443_n
  );


  buf

  (
    g445_p_spl_,
    g445_p
  );


  buf

  (
    g443_p_spl_,
    g443_p
  );


  buf

  (
    g445_n_spl_,
    g445_n
  );


  buf

  (
    g446_p_spl_,
    g446_p
  );


  buf

  (
    g446_p_spl_0,
    g446_p_spl_
  );


  buf

  (
    g448_p_spl_,
    g448_p
  );


  buf

  (
    g446_n_spl_,
    g446_n
  );


  buf

  (
    g446_n_spl_0,
    g446_n_spl_
  );


  buf

  (
    g448_n_spl_,
    g448_n
  );


  buf

  (
    g449_p_spl_,
    g449_p
  );


  buf

  (
    g449_p_spl_0,
    g449_p_spl_
  );


  buf

  (
    g451_p_spl_,
    g451_p
  );


  buf

  (
    g449_n_spl_,
    g449_n
  );


  buf

  (
    g449_n_spl_0,
    g449_n_spl_
  );


  buf

  (
    g451_n_spl_,
    g451_n
  );


  buf

  (
    g453_p_spl_,
    g453_p
  );


  buf

  (
    g453_n_spl_,
    g453_n
  );


  buf

  (
    g454_p_spl_,
    g454_p
  );


  buf

  (
    g454_p_spl_0,
    g454_p_spl_
  );


  buf

  (
    g456_p_spl_,
    g456_p
  );


  buf

  (
    g454_n_spl_,
    g454_n
  );


  buf

  (
    g454_n_spl_0,
    g454_n_spl_
  );


  buf

  (
    g456_n_spl_,
    g456_n
  );


  buf

  (
    g457_p_spl_,
    g457_p
  );


  buf

  (
    g457_p_spl_0,
    g457_p_spl_
  );


  buf

  (
    g459_p_spl_,
    g459_p
  );


  buf

  (
    g457_n_spl_,
    g457_n
  );


  buf

  (
    g457_n_spl_0,
    g457_n_spl_
  );


  buf

  (
    g459_n_spl_,
    g459_n
  );


  buf

  (
    g460_p_spl_,
    g460_p
  );


  buf

  (
    g460_p_spl_0,
    g460_p_spl_
  );


  buf

  (
    g462_p_spl_,
    g462_p
  );


  buf

  (
    g460_n_spl_,
    g460_n
  );


  buf

  (
    g460_n_spl_0,
    g460_n_spl_
  );


  buf

  (
    g462_n_spl_,
    g462_n
  );


  buf

  (
    g463_p_spl_,
    g463_p
  );


  buf

  (
    g463_p_spl_0,
    g463_p_spl_
  );


  buf

  (
    g465_p_spl_,
    g465_p
  );


  buf

  (
    g463_n_spl_,
    g463_n
  );


  buf

  (
    g463_n_spl_0,
    g463_n_spl_
  );


  buf

  (
    g465_n_spl_,
    g465_n
  );


  buf

  (
    g452_n_spl_,
    g452_n
  );


  buf

  (
    g452_p_spl_,
    g452_p
  );


  buf

  (
    g466_p_spl_,
    g466_p
  );


  buf

  (
    g466_p_spl_0,
    g466_p_spl_
  );


  buf

  (
    g468_p_spl_,
    g468_p
  );


  buf

  (
    g466_n_spl_,
    g466_n
  );


  buf

  (
    g466_n_spl_0,
    g466_n_spl_
  );


  buf

  (
    g468_n_spl_,
    g468_n
  );


  buf

  (
    g469_n_spl_,
    g469_n
  );


  buf

  (
    g469_p_spl_,
    g469_p
  );


  buf

  (
    g429_n_spl_,
    g429_n
  );


  buf

  (
    g429_p_spl_,
    g429_p
  );


  buf

  (
    g470_n_spl_,
    g470_n
  );


  buf

  (
    g472_p_spl_,
    g472_p
  );


  buf

  (
    g470_p_spl_,
    g470_p
  );


  buf

  (
    g472_n_spl_,
    g472_n
  );


  buf

  (
    g473_n_spl_,
    g473_n
  );


  buf

  (
    g473_p_spl_,
    g473_p
  );


  buf

  (
    g394_n_spl_,
    g394_n
  );


  buf

  (
    g394_p_spl_,
    g394_p
  );


  buf

  (
    g474_n_spl_,
    g474_n
  );


  buf

  (
    g476_p_spl_,
    g476_p
  );


  buf

  (
    g474_p_spl_,
    g474_p
  );


  buf

  (
    g476_n_spl_,
    g476_n
  );


  buf

  (
    g477_n_spl_,
    g477_n
  );


  buf

  (
    g477_p_spl_,
    g477_p
  );


  buf

  (
    g349_n_spl_,
    g349_n
  );


  buf

  (
    g349_p_spl_,
    g349_p
  );


  buf

  (
    g478_n_spl_,
    g478_n
  );


  buf

  (
    g480_p_spl_,
    g480_p
  );


  buf

  (
    g478_p_spl_,
    g478_p
  );


  buf

  (
    g480_n_spl_,
    g480_n
  );


  buf

  (
    g481_n_spl_,
    g481_n
  );


  buf

  (
    g481_p_spl_,
    g481_p
  );


  buf

  (
    g303_p_spl_,
    g303_p
  );


  buf

  (
    g482_n_spl_,
    g482_n
  );


  buf

  (
    g303_n_spl_,
    g303_n
  );


  buf

  (
    g482_p_spl_,
    g482_p
  );


  buf

  (
    g483_n_spl_,
    g483_n
  );


  buf

  (
    g483_p_spl_,
    g483_p
  );


  buf

  (
    g240_p_spl_,
    g240_p
  );


  buf

  (
    g484_n_spl_,
    g484_n
  );


  buf

  (
    g240_n_spl_,
    g240_n
  );


  buf

  (
    g484_p_spl_,
    g484_p
  );


  buf

  (
    g485_n_spl_,
    g485_n
  );


  buf

  (
    g485_p_spl_,
    g485_p
  );


  buf

  (
    g185_n_spl_,
    g185_n
  );


  buf

  (
    g185_p_spl_,
    g185_p
  );


  buf

  (
    g486_n_spl_,
    g486_n
  );


  buf

  (
    g488_p_spl_,
    g488_p
  );


  buf

  (
    g486_p_spl_,
    g486_p
  );


  buf

  (
    g488_n_spl_,
    g488_n
  );


  buf

  (
    g489_n_spl_,
    g489_n
  );


  buf

  (
    g489_p_spl_,
    g489_p
  );


  buf

  (
    g137_n_spl_,
    g137_n
  );


  buf

  (
    g137_p_spl_,
    g137_p
  );


  buf

  (
    g490_n_spl_,
    g490_n
  );


  buf

  (
    g492_p_spl_,
    g492_p
  );


  buf

  (
    g490_p_spl_,
    g490_p
  );


  buf

  (
    g492_n_spl_,
    g492_n
  );


  buf

  (
    g493_n_spl_,
    g493_n
  );


  buf

  (
    g493_p_spl_,
    g493_p
  );


  buf

  (
    g498_p_spl_,
    g498_p
  );


  buf

  (
    g498_n_spl_,
    g498_n
  );


  buf

  (
    g499_n_spl_,
    g499_n
  );


  buf

  (
    g499_n_spl_0,
    g499_n_spl_
  );


  buf

  (
    g499_p_spl_,
    g499_p
  );


  buf

  (
    g499_p_spl_0,
    g499_p_spl_
  );


  buf

  (
    g501_n_spl_,
    g501_n
  );


  buf

  (
    g501_p_spl_,
    g501_p
  );


  buf

  (
    g502_n_spl_,
    g502_n
  );


  buf

  (
    g502_p_spl_,
    g502_p
  );


  buf

  (
    g504_n_spl_,
    g504_n
  );


  buf

  (
    g505_n_spl_,
    g505_n
  );


  buf

  (
    g504_p_spl_,
    g504_p
  );


  buf

  (
    g505_p_spl_,
    g505_p
  );


  buf

  (
    g506_n_spl_,
    g506_n
  );


  buf

  (
    g506_p_spl_,
    g506_p
  );


  buf

  (
    g496_n_spl_,
    g496_n
  );


  buf

  (
    g508_p_spl_,
    g508_p
  );


  buf

  (
    g496_p_spl_,
    g496_p
  );


  buf

  (
    g508_n_spl_,
    g508_n
  );


  buf

  (
    g509_n_spl_,
    g509_n
  );


  buf

  (
    g509_p_spl_,
    g509_p
  );


  buf

  (
    g495_n_spl_,
    g495_n
  );


  buf

  (
    g511_p_spl_,
    g511_p
  );


  buf

  (
    g495_p_spl_,
    g495_p
  );


  buf

  (
    g511_n_spl_,
    g511_n
  );


  buf

  (
    g512_n_spl_,
    g512_n
  );


  buf

  (
    g512_p_spl_,
    g512_p
  );


  buf

  (
    g494_n_spl_,
    g494_n
  );


  buf

  (
    g514_p_spl_,
    g514_p
  );


  buf

  (
    g494_p_spl_,
    g494_p
  );


  buf

  (
    g514_n_spl_,
    g514_n
  );


  buf

  (
    g516_p_spl_,
    g516_p
  );


  buf

  (
    g516_n_spl_,
    g516_n
  );


  buf

  (
    g515_n_spl_,
    g515_n
  );


  buf

  (
    g515_p_spl_,
    g515_p
  );


  buf

  (
    g533_n_spl_,
    g533_n
  );


  buf

  (
    g535_n_spl_,
    g535_n
  );


  buf

  (
    g533_p_spl_,
    g533_p
  );


  buf

  (
    g535_p_spl_,
    g535_p
  );


  buf

  (
    g531_n_spl_,
    g531_n
  );


  buf

  (
    g531_p_spl_,
    g531_p
  );


  buf

  (
    g529_n_spl_,
    g529_n
  );


  buf

  (
    g529_p_spl_,
    g529_p
  );


  buf

  (
    g540_n_spl_,
    g540_n
  );


  buf

  (
    g542_n_spl_,
    g542_n
  );


  buf

  (
    g540_p_spl_,
    g540_p
  );


  buf

  (
    g542_p_spl_,
    g542_p
  );


  buf

  (
    g525_n_spl_,
    g525_n
  );


  buf

  (
    g525_p_spl_,
    g525_p
  );


  buf

  (
    g523_n_spl_,
    g523_n
  );


  buf

  (
    g523_n_spl_0,
    g523_n_spl_
  );


  buf

  (
    g523_n_spl_1,
    g523_n_spl_
  );


  buf

  (
    g523_p_spl_,
    g523_p
  );


  buf

  (
    g523_p_spl_0,
    g523_p_spl_
  );


  buf

  (
    g523_p_spl_1,
    g523_p_spl_
  );


  buf

  (
    g554_n_spl_,
    g554_n
  );


  buf

  (
    g554_n_spl_0,
    g554_n_spl_
  );


  buf

  (
    g554_n_spl_00,
    g554_n_spl_0
  );


  buf

  (
    g554_n_spl_01,
    g554_n_spl_0
  );


  buf

  (
    g554_n_spl_1,
    g554_n_spl_
  );


  buf

  (
    g554_n_spl_10,
    g554_n_spl_1
  );


  buf

  (
    g554_p_spl_,
    g554_p
  );


  buf

  (
    g554_p_spl_0,
    g554_p_spl_
  );


  buf

  (
    g554_p_spl_00,
    g554_p_spl_0
  );


  buf

  (
    g554_p_spl_01,
    g554_p_spl_0
  );


  buf

  (
    g554_p_spl_1,
    g554_p_spl_
  );


  buf

  (
    g554_p_spl_10,
    g554_p_spl_1
  );


  buf

  (
    g547_n_spl_,
    g547_n
  );


  buf

  (
    g547_n_spl_0,
    g547_n_spl_
  );


  buf

  (
    g547_n_spl_00,
    g547_n_spl_0
  );


  buf

  (
    g547_n_spl_01,
    g547_n_spl_0
  );


  buf

  (
    g547_n_spl_1,
    g547_n_spl_
  );


  buf

  (
    g547_n_spl_10,
    g547_n_spl_1
  );


  buf

  (
    g547_p_spl_,
    g547_p
  );


  buf

  (
    g547_p_spl_0,
    g547_p_spl_
  );


  buf

  (
    g547_p_spl_00,
    g547_p_spl_0
  );


  buf

  (
    g547_p_spl_01,
    g547_p_spl_0
  );


  buf

  (
    g547_p_spl_1,
    g547_p_spl_
  );


  buf

  (
    g547_p_spl_10,
    g547_p_spl_1
  );


  buf

  (
    g558_n_spl_,
    g558_n
  );


  buf

  (
    g559_p_spl_,
    g559_p
  );


  buf

  (
    g558_p_spl_,
    g558_p
  );


  buf

  (
    g559_n_spl_,
    g559_n
  );


  buf

  (
    g559_n_spl_0,
    g559_n_spl_
  );


  buf

  (
    g564_n_spl_,
    g564_n
  );


  buf

  (
    g565_p_spl_,
    g565_p
  );


  buf

  (
    g564_p_spl_,
    g564_p
  );


  buf

  (
    g565_n_spl_,
    g565_n
  );


  buf

  (
    g565_n_spl_0,
    g565_n_spl_
  );


  buf

  (
    g570_n_spl_,
    g570_n
  );


  buf

  (
    g571_p_spl_,
    g571_p
  );


  buf

  (
    g570_p_spl_,
    g570_p
  );


  buf

  (
    g571_n_spl_,
    g571_n
  );


  buf

  (
    g571_n_spl_0,
    g571_n_spl_
  );


  buf

  (
    g572_n_spl_,
    g572_n
  );


  buf

  (
    g572_p_spl_,
    g572_p
  );


  buf

  (
    g578_n_spl_,
    g578_n
  );


  buf

  (
    g579_p_spl_,
    g579_p
  );


  buf

  (
    g578_p_spl_,
    g578_p
  );


  buf

  (
    g579_n_spl_,
    g579_n
  );


  buf

  (
    g579_n_spl_0,
    g579_n_spl_
  );


  buf

  (
    g585_n_spl_,
    g585_n
  );


  buf

  (
    g586_p_spl_,
    g586_p
  );


  buf

  (
    g585_p_spl_,
    g585_p
  );


  buf

  (
    g586_n_spl_,
    g586_n
  );


  buf

  (
    g586_n_spl_0,
    g586_n_spl_
  );


  buf

  (
    g589_p_spl_,
    g589_p
  );


  buf

  (
    g595_n_spl_,
    g595_n
  );


  buf

  (
    g589_n_spl_,
    g589_n
  );


  buf

  (
    g589_n_spl_0,
    g589_n_spl_
  );


  buf

  (
    g595_p_spl_,
    g595_p
  );


  buf

  (
    g598_n_spl_,
    g598_n
  );


  buf

  (
    g598_n_spl_0,
    g598_n_spl_
  );


  buf

  (
    g600_n_spl_,
    g600_n
  );


  buf

  (
    g597_n_spl_,
    g597_n
  );


  buf

  (
    g601_p_spl_,
    g601_p
  );


  buf

  (
    g601_p_spl_0,
    g601_p_spl_
  );


  buf

  (
    g597_p_spl_,
    g597_p
  );


  buf

  (
    g601_n_spl_,
    g601_n
  );


  buf

  (
    g596_n_spl_,
    g596_n
  );


  buf

  (
    g596_p_spl_,
    g596_p
  );


  buf

  (
    g588_n_spl_,
    g588_n
  );


  buf

  (
    g603_n_spl_,
    g603_n
  );


  buf

  (
    g588_p_spl_,
    g588_p
  );


  buf

  (
    g603_p_spl_,
    g603_p
  );


  buf

  (
    g587_n_spl_,
    g587_n
  );


  buf

  (
    g587_p_spl_,
    g587_p
  );


  buf

  (
    g581_n_spl_,
    g581_n
  );


  buf

  (
    g605_n_spl_,
    g605_n
  );


  buf

  (
    g581_p_spl_,
    g581_p
  );


  buf

  (
    g605_p_spl_,
    g605_p
  );


  buf

  (
    g580_n_spl_,
    g580_n
  );


  buf

  (
    g580_p_spl_,
    g580_p
  );


  buf

  (
    g574_n_spl_,
    g574_n
  );


  buf

  (
    g607_p_spl_,
    g607_p
  );


  buf

  (
    g608_p_spl_,
    g608_p
  );


  buf

  (
    g566_n_spl_,
    g566_n
  );


  buf

  (
    g566_p_spl_,
    g566_p
  );


  buf

  (
    g609_p_spl_,
    g609_p
  );


  buf

  (
    g611_n_spl_,
    g611_n
  );


  buf

  (
    g612_p_spl_,
    g612_p
  );


  buf

  (
    g560_n_spl_,
    g560_n
  );


  buf

  (
    g560_p_spl_,
    g560_p
  );


  buf

  (
    g613_p_spl_,
    g613_p
  );


  buf

  (
    g615_n_spl_,
    g615_n
  );


  buf

  (
    g616_p_spl_,
    g616_p
  );


  buf

  (
    g27_n_spl_,
    g27_n
  );


  buf

  (
    g617_p_spl_,
    g617_p
  );


  buf

  (
    g617_p_spl_0,
    g617_p_spl_
  );


  buf

  (
    g618_n_spl_,
    g618_n
  );


  buf

  (
    g618_p_spl_,
    g618_p
  );


  buf

  (
    g621_p_spl_,
    g621_p
  );


  buf

  (
    g622_p_spl_,
    g622_p
  );


  buf

  (
    g617_n_spl_,
    g617_n
  );


  buf

  (
    g622_n_spl_,
    g622_n
  );


  buf

  (
    g620_p_spl_,
    g620_p
  );


  buf

  (
    g620_p_spl_0,
    g620_p_spl_
  );


  buf

  (
    g620_p_spl_00,
    g620_p_spl_0
  );


  buf

  (
    g620_p_spl_01,
    g620_p_spl_0
  );


  buf

  (
    g620_p_spl_1,
    g620_p_spl_
  );


  buf

  (
    g620_p_spl_10,
    g620_p_spl_1
  );


  buf

  (
    g620_p_spl_11,
    g620_p_spl_1
  );


  buf

  (
    g626_n_spl_,
    g626_n
  );


  buf

  (
    g630_p_spl_,
    g630_p
  );


  buf

  (
    g630_p_spl_0,
    g630_p_spl_
  );


  buf

  (
    g630_p_spl_00,
    g630_p_spl_0
  );


  buf

  (
    g630_p_spl_01,
    g630_p_spl_0
  );


  buf

  (
    g630_p_spl_1,
    g630_p_spl_
  );


  buf

  (
    g630_p_spl_10,
    g630_p_spl_1
  );


  buf

  (
    g628_n_spl_,
    g628_n
  );


  buf

  (
    g628_n_spl_0,
    g628_n_spl_
  );


  buf

  (
    g628_n_spl_00,
    g628_n_spl_0
  );


  buf

  (
    g628_n_spl_01,
    g628_n_spl_0
  );


  buf

  (
    g628_n_spl_1,
    g628_n_spl_
  );


  buf

  (
    g628_n_spl_10,
    g628_n_spl_1
  );


  buf

  (
    g628_n_spl_11,
    g628_n_spl_1
  );


  buf

  (
    g636_n_spl_,
    g636_n
  );


  buf

  (
    g645_n_spl_,
    g645_n
  );


  buf

  (
    g654_n_spl_,
    g654_n
  );


  buf

  (
    g663_n_spl_,
    g663_n
  );


  buf

  (
    g670_n_spl_,
    g670_n
  );


  buf

  (
    g677_n_spl_,
    g677_n
  );


  buf

  (
    g684_n_spl_,
    g684_n
  );


endmodule
