// Benchmark "mymod" written by ABC on Sun Oct 29 19:31:54 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58,
    G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70, G71, G72,
    G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86,
    G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G109, G110, G111, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G124,
    G125, G126, G127, G128, G129, G130, G131, G132, G133, G134, G135, G136,
    G137, G138, G139, G140, G141, G142, G143, G144, G145, G146, G147, G148,
    G149, G150, G151, G152, G153, G154, G155, G156, G157,
    G2531, G2532, G2533, G2534, G2535, G2536, G2537, G2538, G2539, G2540,
    G2541, G2542, G2543, G2544, G2545, G2546, G2547, G2548, G2549, G2550,
    G2551, G2552, G2553, G2554, G2555, G2556, G2557, G2558, G2559, G2560,
    G2561, G2562, G2563, G2564, G2565, G2566, G2567, G2568, G2569, G2570,
    G2571, G2572, G2573, G2574, G2575, G2576, G2577, G2578, G2579, G2580,
    G2581, G2582, G2583, G2584, G2585, G2586, G2587, G2588, G2589, G2590,
    G2591, G2592, G2593, G2594  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70,
    G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98,
    G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G110,
    G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G133, G134,
    G135, G136, G137, G138, G139, G140, G141, G142, G143, G144, G145, G146,
    G147, G148, G149, G150, G151, G152, G153, G154, G155, G156, G157;
  output G2531, G2532, G2533, G2534, G2535, G2536, G2537, G2538, G2539, G2540,
    G2541, G2542, G2543, G2544, G2545, G2546, G2547, G2548, G2549, G2550,
    G2551, G2552, G2553, G2554, G2555, G2556, G2557, G2558, G2559, G2560,
    G2561, G2562, G2563, G2564, G2565, G2566, G2567, G2568, G2569, G2570,
    G2571, G2572, G2573, G2574, G2575, G2576, G2577, G2578, G2579, G2580,
    G2581, G2582, G2583, G2584, G2585, G2586, G2587, G2588, G2589, G2590,
    G2591, G2592, G2593, G2594;
  reg n1416_lo, n1419_lo, n1422_lo, n1425_lo, n1428_lo, n1431_lo, n1434_lo,
    n1437_lo, n1440_lo, n1443_lo, n1446_lo, n1449_lo, n1452_lo, n1455_lo,
    n1458_lo, n1464_lo, n1467_lo, n1470_lo, n1476_lo, n1479_lo, n1482_lo,
    n1488_lo, n1491_lo, n1494_lo, n1497_lo, n1500_lo, n1512_lo, n1515_lo,
    n1518_lo, n1521_lo, n1524_lo, n1527_lo, n1530_lo, n1533_lo, n1536_lo,
    n1539_lo, n1542_lo, n1545_lo, n1548_lo, n1551_lo, n1554_lo, n1560_lo,
    n1563_lo, n1566_lo, n1572_lo, n1575_lo, n1578_lo, n1584_lo, n1587_lo,
    n1590_lo, n1596_lo, n1599_lo, n1602_lo, n1608_lo, n1611_lo, n1614_lo,
    n1620_lo, n1623_lo, n1626_lo, n1632_lo, n1635_lo, n1638_lo, n1644_lo,
    n1647_lo, n1650_lo, n1656_lo, n1659_lo, n1662_lo, n1668_lo, n1671_lo,
    n1674_lo, n1677_lo, n1680_lo, n1683_lo, n1686_lo, n1692_lo, n1695_lo,
    n1698_lo, n1704_lo, n1707_lo, n1710_lo, n1716_lo, n1719_lo, n1722_lo,
    n1728_lo, n1731_lo, n1734_lo, n1740_lo, n1743_lo, n1746_lo, n1749_lo,
    n1752_lo, n1755_lo, n1758_lo, n1761_lo, n1764_lo, n1776_lo, n1779_lo,
    n1788_lo, n1791_lo, n1794_lo, n1797_lo, n1800_lo, n1812_lo, n1824_lo,
    n1836_lo, n1848_lo, n1860_lo, n1872_lo, n1884_lo, n1896_lo, n1899_lo,
    n1908_lo, n1911_lo, n1920_lo, n1923_lo, n1926_lo, n1929_lo, n1932_lo,
    n1944_lo, n1956_lo, n1968_lo, n1980_lo, n1992_lo, n2004_lo, n2016_lo,
    n2019_lo, n2028_lo, n2031_lo, n2040_lo, n2043_lo, n2046_lo, n2049_lo,
    n2052_lo, n2064_lo, n2076_lo, n2088_lo, n2100_lo, n2112_lo, n2124_lo,
    n2136_lo, n2148_lo, n2151_lo, n2160_lo, n2163_lo, n2172_lo, n2175_lo,
    n2178_lo, n2181_lo, n2184_lo, n2196_lo, n2208_lo, n2220_lo, n2232_lo,
    n2244_lo, n2256_lo, n2268_lo, n2280_lo, n2283_lo, n2292_lo, n2295_lo,
    n2298_lo, n2301_lo, n2304_lo, n2316_lo, n2319_lo, n2322_lo, n2325_lo,
    n2328_lo, n2331_lo, n2340_lo, n2343_lo, n2376_lo, n2379_lo, n2388_lo,
    n2400_lo, n2412_lo, n2415_lo, n2424_lo, n2436_lo, n2439_lo, n2442_lo,
    n2445_lo, n2448_lo, n2451_lo, n2460_lo, n2463_lo, n2496_lo, n2499_lo,
    n2508_lo, n2520_lo, n2532_lo, n2535_lo, n2544_lo, n2556_lo, n2559_lo,
    n2562_lo, n2565_lo, n2568_lo, n2571_lo, n2580_lo, n2583_lo, n2616_lo,
    n2619_lo, n2628_lo, n2640_lo, n2652_lo, n2655_lo, n2664_lo, n2676_lo,
    n2679_lo, n2682_lo, n2685_lo, n2688_lo, n2691_lo, n2700_lo, n2703_lo,
    n2736_lo, n2739_lo, n2748_lo, n2760_lo, n2772_lo, n2775_lo, n2784_lo,
    n2787_lo, n2790_lo, n2793_lo, n2796_lo, n2799_lo, n2802_lo, n2805_lo,
    n2808_lo, n2820_lo, n2823_lo, n2826_lo, n2832_lo, n2835_lo, n2838_lo,
    n2841_lo, n2844_lo, n2856_lo, n2859_lo, n2862_lo, n2865_lo, n2868_lo,
    n2871_lo, n2874_lo, n2877_lo, n2880_lo, n2883_lo, n2886_lo, n2889_lo,
    n2892_lo, n2895_lo, n2898_lo, n2901_lo, n2904_lo, n2907_lo, n2916_lo,
    n2928_lo, n2940_lo, n2952_lo, n2955_lo, n2964_lo, n2976_lo, n2988_lo,
    n2991_lo, n3000_lo, n3003_lo, n3012_lo, n3015_lo, n3024_lo, n3027_lo,
    n3036_lo, n3039_lo, n3048_lo, n3051_lo, n3054_lo, n3057_lo, n3060_lo,
    n3072_lo, n3081_lo, n3084_lo, n3087_lo, n3093_lo, n3096_lo, n3105_lo,
    n3108_lo, n3117_lo, n3120_lo, n3123_lo, n3126_lo, n3129_lo, n3132_lo,
    n3135_lo, n3138_lo, n3141_lo, n3168_lo, n3171_lo, n3174_lo, n3177_lo,
    n3180_lo, n3183_lo, n3192_lo, n3195_lo, n3204_lo, n3207_lo, n3216_lo,
    n3219_lo, n3228_lo, n3231_lo, n3240_lo, n3243_lo, n3252_lo, n3255_lo,
    n3258_lo, n3264_lo, n3267_lo, n3270_lo, n3276_lo, n3279_lo, n3282_lo,
    n3288_lo, n3291_lo, n3294_lo, n4537_o2, n4538_o2, n4710_o2, n4711_o2,
    n1211_inv, n1214_inv, n1217_inv, n1220_inv, n4927_o2, n4928_o2,
    n1229_inv, n1232_inv, n1235_inv, n5178_o2, n5179_o2, n5477_o2,
    n5478_o2, n5479_o2, n5222_o2, n5223_o2, n5553_o2, n5554_o2, G491_o2,
    n2922_lo_buf_o2, n2946_lo_buf_o2, n2970_lo_buf_o2, n2982_lo_buf_o2,
    n3066_lo_buf_o2, n3078_lo_buf_o2, n3102_lo_buf_o2, n3114_lo_buf_o2,
    G1321_o2, G1033_o2, G1030_o2, G1072_o2, n1304_inv, n1307_inv,
    n2958_lo_buf_o2, n2994_lo_buf_o2, n3006_lo_buf_o2, n3030_lo_buf_o2,
    n3042_lo_buf_o2, n3090_lo_buf_o2, n1328_inv, n1331_inv, n1334_inv,
    n1337_inv, n1340_inv, n1343_inv, n1346_inv, n1349_inv, G1036_o2,
    G1062_o2, G1067_o2, G1014_o2, n1364_inv, n1367_inv, n3018_lo_buf_o2,
    G766_o2, n1376_inv, n1379_inv, n1382_inv, n1385_inv, n1388_inv,
    n1391_inv, G1017_o2, G1008_o2, n1400_inv, n1403_inv, n2910_lo_buf_o2,
    n1409_inv, G2138_o2, G2147_o2, n1418_inv, G1137_o2, G1329_o2, G374_o2,
    G386_o2, G663_o2, G674_o2, G578_o2, G575_o2, G2505_o2, n1448_inv,
    G987_o2, G984_o2, G1862_o2, G1859_o2, G1260_o2, G1865_o2, G2073_o2,
    G1402_o2, G2048_o2, G2276_o2, n1481_inv, G2141_o2, G2008_o2, G2011_o2,
    G2150_o2, G2026_o2, G2029_o2, G2023_o2, G2041_o2, G2017_o2, G2020_o2,
    G2035_o2, G2038_o2, G2228_o2, G2231_o2, G2234_o2, G2237_o2, G1904_o2,
    G1907_o2, G1928_o2, G1931_o2, G1893_o2, G1896_o2, G1899_o2, G1937_o2,
    G1940_o2, G1943_o2, G1336_o2, G1996_o2, G1999_o2, G2002_o2, G2005_o2,
    G2014_o2, G2032_o2, G1076_o2, G1002_o2, G998_o2, G1890_o2, G1934_o2,
    G1044_o2, G1039_o2, n1770_lo_buf_o2, G342_o2, G354_o2, G1193_o2,
    n3234_lo_buf_o2, n3246_lo_buf_o2, G783_o2, G786_o2, G792_o2, G795_o2,
    G815_o2, G818_o2, G824_o2, G827_o2, G789_o2, G798_o2, G801_o2, G807_o2,
    G812_o2, G821_o2, G804_o2, G780_o2, G1231_o2, G1572_o2, G1377_o2,
    G1253_o2, G1359_o2, G1258_o2, G1367_o2, G1358_o2, G1366_o2, G2057_o2,
    G2117_o2, G2118_o2, G1254_o2, G1259_o2, G2058_o2, G405_o2, G417_o2,
    G1269_o2, G1275_o2, G1287_o2, G1266_o2, G1272_o2, G1278_o2, G1281_o2,
    G1284_o2, G1290_o2, G1293_o2, G1299_o2, G1305_o2, G1296_o2, G1302_o2,
    G1308_o2, G1311_o2, G811_o2, G810_o2, G1728_o2, G2512_o2, G1114_o2,
    G1113_o2, G1992_o2, G1991_o2, G1426_o2, G1966_o2, G2211_o2, G1509_o2,
    G2153_o2, G2329_o2, G1540_o2, G2167_o2, G2191_o2, G1234_o2, G1132_o2,
    G1129_o2, G2088_o2, G2106_o2, G1314_o2, G636_o2, G647_o2,
    n3186_lo_buf_o2, n3198_lo_buf_o2, n3210_lo_buf_o2, n3222_lo_buf_o2,
    G1225_o2, G1342_o2, G1222_o2, G1228_o2, G1348_o2, G1345_o2, G1351_o2,
    G2242_o2, G2260_o2, G1374_o2, G1537_o2, G301_o2, G313_o2, G2365_o2,
    G2255_o2, G2253_o2, G2395_o2, G2272_o2, G2270_o2, G2245_o2, G2262_o2,
    G2249_o2, G2247_o2, G2266_o2, G2264_o2, G2403_o2, G2401_o2, G2410_o2,
    G2408_o2, G2306_o2, G2305_o2, G2314_o2, G2313_o2, G2303_o2, G2302_o2,
    G2301_o2, G2311_o2, G2310_o2, G2309_o2, G2404_o2, G2411_o2, G2420_o2,
    G2419_o2, G2433_o2, G2432_o2, G402_o2, G403_o2, G1053_o2, G1049_o2,
    n2003_inv, G1364_o2, G1079_o2, G1478_o2, G707_o2, G718_o2, G2417_o2,
    G2414_o2, G2431_o2, G2428_o2, G1653_o2, G2213_o2, G2221_o2, G2250_o2,
    G2267_o2, G1365_o2, G1368_o2, G1371_o2, G2218_o2, G2225_o2,
    n1503_lo_buf_o2, n1863_lo_buf_o2, n1887_lo_buf_o2, n1983_lo_buf_o2,
    n2007_lo_buf_o2, n2115_lo_buf_o2, n2139_lo_buf_o2, n2247_lo_buf_o2,
    n2271_lo_buf_o2, n2919_lo_buf_o2, n2943_lo_buf_o2, n2967_lo_buf_o2,
    n2979_lo_buf_o2, n3063_lo_buf_o2, n3075_lo_buf_o2, n3099_lo_buf_o2,
    n3111_lo_buf_o2, G878_o2, G875_o2, G661_o2, G660_o2, G879_o2, G876_o2,
    G1320_o2, G941_o2, G732_o2, G942_o2, G1493_o2, G1498_o2, G877_o2,
    G874_o2, n1806_lo_buf_o2, n1878_lo_buf_o2, n1938_lo_buf_o2,
    n1998_lo_buf_o2, n2058_lo_buf_o2, n2130_lo_buf_o2, n2190_lo_buf_o2,
    n2262_lo_buf_o2, n2310_lo_buf_o2, n2406_lo_buf_o2, n2430_lo_buf_o2,
    n2526_lo_buf_o2, n2550_lo_buf_o2, n2646_lo_buf_o2, n2670_lo_buf_o2,
    n2766_lo_buf_o2, G603_o2, G614_o2, G1026_o2, G1021_o2, G940_o2,
    G1636_o2, G1684_o2, n2352_lo_buf_o2, n2364_lo_buf_o2, n2472_lo_buf_o2,
    n2484_lo_buf_o2, n2592_lo_buf_o2, n2604_lo_buf_o2, n2712_lo_buf_o2,
    n2724_lo_buf_o2, n3150_lo_buf_o2, n3162_lo_buf_o2;
  wire new_n1576_, new_n1578_, new_n1580_, new_n1582_, new_n1584_,
    new_n1586_, new_n1588_, new_n1590_, new_n1592_, new_n1594_, new_n1596_,
    new_n1598_, new_n1600_, new_n1602_, new_n1604_, new_n1606_, new_n1608_,
    new_n1610_, new_n1612_, new_n1614_, new_n1616_, new_n1618_, new_n1620_,
    new_n1622_, new_n1624_, new_n1626_, new_n1628_, new_n1630_, new_n1632_,
    new_n1634_, new_n1636_, new_n1638_, new_n1640_, new_n1642_, new_n1644_,
    new_n1646_, new_n1648_, new_n1650_, new_n1652_, new_n1654_, new_n1656_,
    new_n1658_, new_n1660_, new_n1662_, new_n1664_, new_n1666_, new_n1668_,
    new_n1670_, new_n1672_, new_n1674_, new_n1676_, new_n1678_, new_n1680_,
    new_n1682_, new_n1684_, new_n1686_, new_n1688_, new_n1690_, new_n1692_,
    new_n1694_, new_n1696_, new_n1698_, new_n1700_, new_n1702_, new_n1704_,
    new_n1706_, new_n1708_, new_n1710_, new_n1712_, new_n1714_, new_n1716_,
    new_n1718_, new_n1720_, new_n1722_, new_n1724_, new_n1726_, new_n1728_,
    new_n1730_, new_n1732_, new_n1734_, new_n1736_, new_n1738_, new_n1740_,
    new_n1742_, new_n1744_, new_n1746_, new_n1748_, new_n1750_, new_n1752_,
    new_n1754_, new_n1756_, new_n1758_, new_n1760_, new_n1762_, new_n1764_,
    new_n1766_, new_n1768_, new_n1770_, new_n1772_, new_n1774_, new_n1776_,
    new_n1778_, new_n1780_, new_n1782_, new_n1784_, new_n1786_, new_n1788_,
    new_n1790_, new_n1792_, new_n1794_, new_n1796_, new_n1798_, new_n1800_,
    new_n1802_, new_n1804_, new_n1806_, new_n1808_, new_n1810_, new_n1812_,
    new_n1814_, new_n1816_, new_n1818_, new_n1820_, new_n1822_, new_n1824_,
    new_n1826_, new_n1828_, new_n1830_, new_n1832_, new_n1834_, new_n1836_,
    new_n1838_, new_n1840_, new_n1842_, new_n1844_, new_n1846_, new_n1848_,
    new_n1850_, new_n1852_, new_n1854_, new_n1856_, new_n1858_, new_n1860_,
    new_n1862_, new_n1864_, new_n1866_, new_n1868_, new_n1870_, new_n1872_,
    new_n1874_, new_n1876_, new_n1878_, new_n1880_, new_n1882_, new_n1884_,
    new_n1886_, new_n1888_, new_n1890_, new_n1892_, new_n1894_, new_n1896_,
    new_n1898_, new_n1900_, new_n1902_, new_n1905_, new_n1906_, new_n1908_,
    new_n1910_, new_n1912_, new_n1914_, new_n1916_, new_n1918_, new_n1920_,
    new_n1922_, new_n1924_, new_n1926_, new_n1928_, new_n1930_, new_n1932_,
    new_n1934_, new_n1936_, new_n1939_, new_n1940_, new_n1942_, new_n1944_,
    new_n1946_, new_n1949_, new_n1950_, new_n1952_, new_n1954_, new_n1956_,
    new_n1958_, new_n1960_, new_n1962_, new_n1965_, new_n1966_, new_n1968_,
    new_n1970_, new_n1971_, new_n1972_, new_n1974_, new_n1976_, new_n1978_,
    new_n1980_, new_n1982_, new_n1984_, new_n1986_, new_n1988_, new_n1990_,
    new_n1992_, new_n1994_, new_n1996_, new_n1998_, new_n2000_, new_n2002_,
    new_n2004_, new_n2006_, new_n2008_, new_n2010_, new_n2012_, new_n2014_,
    new_n2016_, new_n2018_, new_n2020_, new_n2022_, new_n2024_, new_n2026_,
    new_n2028_, new_n2030_, new_n2033_, new_n2034_, new_n2036_, new_n2038_,
    new_n2039_, new_n2040_, new_n2042_, new_n2044_, new_n2046_, new_n2048_,
    new_n2050_, new_n2052_, new_n2054_, new_n2056_, new_n2058_, new_n2060_,
    new_n2062_, new_n2064_, new_n2066_, new_n2068_, new_n2071_, new_n2072_,
    new_n2074_, new_n2076_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2084_, new_n2086_, new_n2088_, new_n2090_, new_n2093_, new_n2094_,
    new_n2096_, new_n2098_, new_n2100_, new_n2102_, new_n2104_, new_n2106_,
    new_n2108_, new_n2110_, new_n2112_, new_n2114_, new_n2116_, new_n2118_,
    new_n2120_, new_n2122_, new_n2125_, new_n2126_, new_n2128_, new_n2130_,
    new_n2132_, new_n2134_, new_n2136_, new_n2138_, new_n2140_, new_n2142_,
    new_n2144_, new_n2146_, new_n2148_, new_n2150_, new_n2152_, new_n2155_,
    new_n2156_, new_n2158_, new_n2160_, new_n2162_, new_n2164_, new_n2166_,
    new_n2168_, new_n2170_, new_n2172_, new_n2174_, new_n2176_, new_n2178_,
    new_n2180_, new_n2182_, new_n2184_, new_n2187_, new_n2188_, new_n2190_,
    new_n2192_, new_n2194_, new_n2196_, new_n2198_, new_n2200_, new_n2202_,
    new_n2204_, new_n2206_, new_n2208_, new_n2210_, new_n2212_, new_n2214_,
    new_n2216_, new_n2218_, new_n2220_, new_n2222_, new_n2225_, new_n2226_,
    new_n2228_, new_n2230_, new_n2232_, new_n2234_, new_n2236_, new_n2238_,
    new_n2240_, new_n2242_, new_n2244_, new_n2246_, new_n2248_, new_n2250_,
    new_n2252_, new_n2255_, new_n2256_, new_n2258_, new_n2260_, new_n2262_,
    new_n2264_, new_n2266_, new_n2268_, new_n2270_, new_n2272_, new_n2274_,
    new_n2276_, new_n2278_, new_n2280_, new_n2282_, new_n2285_, new_n2286_,
    new_n2288_, new_n2290_, new_n2292_, new_n2294_, new_n2296_, new_n2298_,
    new_n2300_, new_n2302_, new_n2304_, new_n2306_, new_n2308_, new_n2310_,
    new_n2312_, new_n2315_, new_n2316_, new_n2318_, new_n2320_, new_n2322_,
    new_n2324_, new_n2326_, new_n2328_, new_n2330_, new_n2332_, new_n2334_,
    new_n2336_, new_n2338_, new_n2340_, new_n2342_, new_n2343_, new_n2344_,
    new_n2346_, new_n2348_, new_n2351_, new_n2352_, new_n2353_, new_n2354_,
    new_n2356_, new_n2358_, new_n2359_, new_n2360_, new_n2362_, new_n2364_,
    new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2372_,
    new_n2374_, new_n2376_, new_n2377_, new_n2378_, new_n2380_, new_n2382_,
    new_n2384_, new_n2385_, new_n2386_, new_n2388_, new_n2390_, new_n2392_,
    new_n2393_, new_n2394_, new_n2396_, new_n2398_, new_n2401_, new_n2402_,
    new_n2404_, new_n2406_, new_n2408_, new_n2410_, new_n2412_, new_n2414_,
    new_n2415_, new_n2416_, new_n2418_, new_n2420_, new_n2422_, new_n2424_,
    new_n2426_, new_n2428_, new_n2430_, new_n2431_, new_n2432_, new_n2434_,
    new_n2435_, new_n2436_, new_n2438_, new_n2439_, new_n2440_, new_n2442_,
    new_n2444_, new_n2447_, new_n2448_, new_n2450_, new_n2453_, new_n2454_,
    new_n2456_, new_n2457_, new_n2459_, new_n2460_, new_n2463_, new_n2464_,
    new_n2467_, new_n2468_, new_n2470_, new_n2472_, new_n2474_, new_n2475_,
    new_n2476_, new_n2478_, new_n2480_, new_n2482_, new_n2483_, new_n2484_,
    new_n2486_, new_n2488_, new_n2490_, new_n2491_, new_n2492_, new_n2494_,
    new_n2496_, new_n2498_, new_n2500_, new_n2502_, new_n2504_, new_n2506_,
    new_n2508_, new_n2510_, new_n2512_, new_n2514_, new_n2516_, new_n2518_,
    new_n2520_, new_n2521_, new_n2522_, new_n2524_, new_n2526_, new_n2527_,
    new_n2528_, new_n2530_, new_n2532_, new_n2533_, new_n2534_, new_n2536_,
    new_n2538_, new_n2539_, new_n2541_, new_n2543_, new_n2545_, new_n2547_,
    new_n2548_, new_n2550_, new_n2552_, new_n2554_, new_n2557_, new_n2558_,
    new_n2559_, new_n2560_, new_n2562_, new_n2564_, new_n2566_, new_n2567_,
    new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2580_, new_n2582_,
    new_n2584_, new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_,
    new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_,
    new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2604_, new_n2606_, new_n2608_, new_n2610_, new_n2612_,
    new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_,
    new_n2620_, new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_,
    new_n2626_, new_n2628_, new_n2630_, new_n2632_, new_n2634_, new_n2636_,
    new_n2638_, new_n2640_, new_n2642_, new_n2644_, new_n2646_, new_n2648_,
    new_n2650_, new_n2652_, new_n2654_, new_n2655_, new_n2657_, new_n2658_,
    new_n2660_, new_n2662_, new_n2664_, new_n2666_, new_n2668_, new_n2670_,
    new_n2672_, new_n2673_, new_n2674_, new_n2676_, new_n2678_, new_n2679_,
    new_n2680_, new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_,
    new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_,
    new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_,
    new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_,
    new_n2713_, new_n2714_, new_n2715_, new_n2717_, new_n2718_, new_n2721_,
    new_n2722_, new_n2725_, new_n2726_, new_n2728_, new_n2730_, new_n2731_,
    new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_,
    new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2744_,
    new_n2746_, new_n2748_, new_n2750_, new_n2752_, new_n2754_, new_n2755_,
    new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_,
    new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_,
    new_n2768_, new_n2769_, new_n2771_, new_n2773_, new_n2775_, new_n2777_,
    new_n2779_, new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_,
    new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_,
    new_n2792_, new_n2794_, new_n2796_, new_n2798_, new_n2799_, new_n2800_,
    new_n2803_, new_n2805_, new_n2806_, new_n2808_, new_n2810_, new_n2811_,
    new_n2813_, new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_,
    new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_,
    new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_,
    new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_,
    new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_,
    new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_,
    new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_,
    new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_,
    new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_,
    new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_,
    new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_,
    new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2885_, new_n2887_,
    new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_,
    new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_,
    new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_,
    new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_,
    new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_,
    new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_,
    new_n2924_, new_n2925_, new_n2926_, new_n2928_, new_n2929_, new_n2930_,
    new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_,
    new_n2939_, new_n2940_, new_n2943_, new_n2944_, new_n2947_, new_n2948_,
    new_n2949_, new_n2951_, new_n2953_, new_n2954_, new_n2955_, new_n2956_,
    new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2962_, new_n2964_,
    new_n2965_, new_n2966_, new_n2968_, new_n2970_, new_n2971_, new_n2972_,
    new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_,
    new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_,
    new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_,
    new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_,
    new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_,
    new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_,
    new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_,
    new_n3015_, new_n3017_, new_n3019_, new_n3021_, new_n3023_, new_n3025_,
    new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_,
    new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_,
    new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_,
    new_n3046_, new_n3048_, new_n3050_, new_n3052_, new_n3054_, new_n3056_,
    new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_,
    new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_,
    new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_,
    new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_,
    new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3086_, new_n3088_,
    new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_,
    new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_,
    new_n3101_, new_n3102_, new_n3104_, new_n3106_, new_n3107_, new_n3108_,
    new_n3109_, new_n3110_, new_n3111_, new_n3113_, new_n3115_, new_n3117_,
    new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_,
    new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_,
    new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_,
    new_n3136_, new_n3137_, new_n3138_, new_n3140_, new_n3142_, new_n3143_,
    new_n3144_, new_n3145_, new_n3146_, new_n3148_, new_n3150_, new_n3152_,
    new_n3154_, new_n3156_, new_n3158_, new_n3160_, new_n3162_, new_n3163_,
    new_n3164_, new_n3166_, new_n3168_, new_n3170_, new_n3171_, new_n3172_,
    new_n3173_, new_n3174_, new_n3176_, new_n3178_, new_n3180_, new_n3181_,
    new_n3182_, new_n3184_, new_n3185_, new_n3186_, new_n3188_, new_n3189_,
    new_n3190_, new_n3192_, new_n3193_, new_n3194_, new_n3196_, new_n3198_,
    new_n3200_, new_n3202_, new_n3204_, new_n3206_, new_n3208_, new_n3210_,
    new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3216_, new_n3218_,
    new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3227_,
    new_n3228_, new_n3231_, new_n3232_, new_n3235_, new_n3236_, new_n3239_,
    new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_,
    new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_,
    new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_,
    new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_,
    new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_,
    new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_,
    new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_,
    new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_,
    new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_,
    new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_,
    new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_,
    new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_,
    new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_,
    new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_,
    new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_,
    new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_,
    new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_,
    new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_,
    new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_,
    new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_,
    new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_,
    new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_,
    new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_,
    new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_,
    new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_,
    new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_,
    new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_,
    new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_,
    new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_,
    new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_,
    new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_,
    new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_,
    new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_,
    new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_,
    new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_,
    new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_,
    new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_,
    new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_,
    new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_,
    new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_,
    new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_,
    new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_,
    new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_,
    new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_,
    new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_,
    new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_,
    new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_,
    new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_,
    new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_,
    new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_,
    new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_,
    new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_,
    new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_,
    new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_,
    new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_,
    new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_,
    new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_,
    new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_,
    new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_,
    new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_,
    new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_,
    new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_,
    new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_,
    new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_,
    new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_,
    new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_,
    new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_,
    new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_,
    new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_,
    new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_,
    new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_,
    new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_,
    new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_,
    new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_,
    new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_,
    new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_,
    new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_,
    new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_,
    new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_,
    new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_,
    new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_,
    new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_,
    new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_,
    new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_,
    new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_,
    new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_,
    new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_,
    new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_,
    new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_,
    new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_,
    new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_,
    new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_,
    new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_,
    new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_,
    new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_,
    new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_,
    new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_,
    new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_,
    new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_,
    new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_,
    new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_,
    new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_,
    new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_,
    new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_,
    new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_,
    new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_,
    new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_,
    new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_,
    new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_,
    new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_,
    new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_,
    new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_,
    new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_,
    new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_,
    new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_,
    new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_,
    new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_,
    new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_,
    new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_,
    new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_,
    new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_,
    new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_,
    new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_,
    new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_,
    new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_,
    new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_,
    new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_,
    new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_,
    new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_,
    new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_,
    new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_,
    new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_,
    new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_,
    new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_,
    new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_,
    new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_,
    new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_,
    new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_,
    new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_,
    new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_,
    new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_,
    new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_,
    new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_,
    new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_,
    new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_,
    new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_,
    new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_,
    new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_,
    new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_,
    new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_,
    new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_,
    new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_,
    new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n5047_, new_n5048_,
    new_n5049_, new_n5050_, new_n5051_, new_n5052_, new_n5053_, new_n5054_,
    new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_, new_n5060_,
    new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_, new_n5066_,
    new_n5067_, new_n5068_, new_n5069_, new_n5070_, new_n5071_, new_n5072_,
    new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_, new_n5078_,
    new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_, new_n5084_,
    new_n5085_, new_n5086_, new_n5087_, new_n5088_, new_n5089_, new_n5090_,
    new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_, new_n5096_,
    new_n5097_, new_n5098_, new_n5099_, new_n5100_, new_n5101_, new_n5102_,
    new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_, new_n5108_,
    new_n5109_, new_n5110_, new_n5111_, new_n5112_, new_n5113_, new_n5114_,
    new_n5115_, new_n5116_, new_n5117_, new_n5118_, new_n5119_, new_n5120_,
    new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_, new_n5126_,
    new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_, new_n5132_,
    new_n5133_, new_n5134_, new_n5135_, new_n5136_, new_n5137_, new_n5138_,
    new_n5139_, new_n5140_, new_n5141_, new_n5142_, new_n5143_, new_n5144_,
    new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_, new_n5150_,
    new_n5151_, new_n5152_, new_n5153_, new_n5154_, new_n5155_, new_n5156_,
    new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5161_, new_n5162_,
    new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5167_, new_n5168_,
    new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5173_, new_n5174_,
    new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5179_, new_n5180_,
    new_n5181_, new_n5182_, new_n5183_, new_n5184_, new_n5185_, new_n5186_,
    new_n5187_, new_n5188_, new_n5189_, new_n5190_, new_n5191_, new_n5192_,
    new_n5193_, new_n5194_, new_n5195_, new_n5196_, new_n5197_, new_n5198_,
    new_n5199_, new_n5200_, new_n5201_, new_n5202_, new_n5203_, new_n5204_,
    new_n5205_, new_n5206_, new_n5207_, new_n5208_, new_n5209_, new_n5210_,
    new_n5211_, new_n5212_, new_n5213_, new_n5214_, new_n5215_, new_n5216_,
    new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_, new_n5222_,
    new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_, new_n5228_,
    new_n5229_, new_n5230_, new_n5231_, new_n5232_, new_n5233_, new_n5234_,
    new_n5235_, new_n5236_, new_n5237_, new_n5238_, new_n5239_, new_n5240_,
    new_n5241_, new_n5242_, new_n5243_, new_n5244_, new_n5245_, new_n5246_,
    new_n5247_, new_n5248_, new_n5249_, new_n5250_, new_n5251_, new_n5252_,
    new_n5253_, new_n5254_, new_n5255_, new_n5256_, new_n5257_, new_n5258_,
    new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5263_, new_n5264_,
    new_n5265_, new_n5266_, new_n5267_, new_n5268_, new_n5269_, new_n5270_,
    new_n5271_, new_n5272_, new_n5273_, new_n5274_, new_n5275_, new_n5276_,
    new_n5277_, new_n5278_, new_n5279_, new_n5280_, new_n5281_, new_n5282_,
    new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_, new_n5288_,
    new_n5289_, new_n5290_, new_n5291_, new_n5292_, new_n5293_, new_n5294_,
    new_n5295_, new_n5296_, new_n5297_, new_n5298_, new_n5299_, new_n5300_,
    new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_, new_n5306_,
    new_n5307_, new_n5308_, new_n5309_, new_n5310_, new_n5311_, new_n5312_,
    new_n5313_, new_n5314_, new_n5315_, new_n5316_, new_n5317_, new_n5318_,
    new_n5319_, new_n5320_, new_n5321_, new_n5322_, new_n5323_, new_n5324_,
    new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_, new_n5330_,
    new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_, new_n5336_,
    new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_, new_n5342_,
    new_n5343_, new_n5344_, new_n5345_, new_n5346_, new_n5347_, new_n5348_,
    new_n5349_, new_n5350_, new_n5351_, new_n5352_, new_n5353_, new_n5354_,
    new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_, new_n5360_,
    new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_, new_n5366_,
    new_n5367_, new_n5368_, new_n5369_, new_n5370_, new_n5371_, new_n5372_,
    new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_, new_n5378_,
    new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_, new_n5384_,
    new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_, new_n5390_,
    new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_, new_n5396_,
    new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_, new_n5402_,
    new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_, new_n5408_,
    new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_, new_n5414_,
    new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_, new_n5420_,
    new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_, new_n5426_,
    new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_, new_n5432_,
    new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_, new_n5438_,
    new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_, new_n5444_,
    new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_, new_n5450_,
    new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_, new_n5456_,
    new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_, new_n5462_,
    new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_, new_n5468_,
    new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_, new_n5474_,
    new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5479_, new_n5480_,
    new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_,
    new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5492_,
    new_n5493_, new_n5494_, new_n5495_, new_n5496_, new_n5497_, new_n5498_,
    new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_, new_n5504_,
    new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_, new_n5510_,
    new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_, new_n5516_,
    new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_, new_n5522_,
    new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_, new_n5528_,
    new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_, new_n5534_,
    new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_, new_n5540_,
    new_n5541_, new_n5542_, new_n5543_, new_n5544_, new_n5545_, new_n5546_,
    new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_, new_n5552_,
    new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_, new_n5558_,
    new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_, new_n5564_,
    new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_, new_n5570_,
    new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_, new_n5576_,
    new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_, new_n5582_,
    new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_, new_n5588_,
    new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_, new_n5594_,
    new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_, new_n5600_,
    new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_, new_n5606_,
    new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_, new_n5612_,
    new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_, new_n5618_,
    new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_, new_n5624_,
    new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_, new_n5630_,
    new_n5631_, new_n5632_, new_n5633_, new_n5634_, new_n5635_, new_n5636_,
    new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_, new_n5642_,
    new_n5643_, new_n5644_, new_n5645_, new_n5646_, new_n5647_, new_n5648_,
    new_n5649_, new_n5650_, new_n5651_, new_n5652_, new_n5653_, new_n5654_,
    new_n5655_, new_n5656_, new_n5657_, new_n5658_, new_n5659_, new_n5660_,
    new_n5661_, new_n5662_, new_n5663_, new_n5664_, new_n5665_, new_n5666_,
    new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_, new_n5672_,
    new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_, new_n5678_,
    new_n5679_, new_n5680_, new_n5681_, new_n5682_, new_n5683_, new_n5684_,
    new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_, new_n5690_,
    new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_, new_n5696_,
    new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_, new_n5702_,
    new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_, new_n5708_,
    new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_, new_n5714_,
    new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_, new_n5720_,
    new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_, new_n5726_,
    new_n5727_, new_n5728_, new_n5729_, new_n5730_, new_n5731_, new_n5732_,
    new_n5733_, new_n5734_, new_n5735_, new_n5736_, new_n5737_, new_n5738_,
    new_n5739_, new_n5740_, new_n5741_, new_n5742_, new_n5743_, new_n5744_,
    new_n5745_, new_n5746_, new_n5747_, new_n5748_, new_n5749_, new_n5750_,
    new_n5751_, new_n5752_, new_n5753_, new_n5754_, new_n5755_, new_n5756_,
    new_n5757_, new_n5758_, new_n5759_, new_n5760_, new_n5761_, new_n5762_,
    new_n5763_, new_n5764_, new_n5765_, new_n5766_, new_n5767_, new_n5768_,
    new_n5769_, new_n5770_, new_n5771_, new_n5772_, new_n5773_, new_n5774_,
    new_n5775_, new_n5776_, new_n5777_, new_n5778_, new_n5779_, new_n5780_,
    new_n5781_, new_n5782_, new_n5783_, new_n5784_, new_n5785_, new_n5786_,
    new_n5787_, new_n5788_, new_n5789_, new_n5790_, n1416_li, n1419_li,
    n1422_li, n1425_li, n1428_li, n1431_li, n1434_li, n1437_li, n1440_li,
    n1443_li, n1446_li, n1449_li, n1452_li, n1455_li, n1458_li, n1464_li,
    n1467_li, n1470_li, n1476_li, n1479_li, n1482_li, n1488_li, n1491_li,
    n1494_li, n1497_li, n1500_li, n1512_li, n1515_li, n1518_li, n1521_li,
    n1524_li, n1527_li, n1530_li, n1533_li, n1536_li, n1539_li, n1542_li,
    n1545_li, n1548_li, n1551_li, n1554_li, n1560_li, n1563_li, n1566_li,
    n1572_li, n1575_li, n1578_li, n1584_li, n1587_li, n1590_li, n1596_li,
    n1599_li, n1602_li, n1608_li, n1611_li, n1614_li, n1620_li, n1623_li,
    n1626_li, n1632_li, n1635_li, n1638_li, n1644_li, n1647_li, n1650_li,
    n1656_li, n1659_li, n1662_li, n1668_li, n1671_li, n1674_li, n1677_li,
    n1680_li, n1683_li, n1686_li, n1692_li, n1695_li, n1698_li, n1704_li,
    n1707_li, n1710_li, n1716_li, n1719_li, n1722_li, n1728_li, n1731_li,
    n1734_li, n1740_li, n1743_li, n1746_li, n1749_li, n1752_li, n1755_li,
    n1758_li, n1761_li, n1764_li, n1776_li, n1779_li, n1788_li, n1791_li,
    n1794_li, n1797_li, n1800_li, n1812_li, n1824_li, n1836_li, n1848_li,
    n1860_li, n1872_li, n1884_li, n1896_li, n1899_li, n1908_li, n1911_li,
    n1920_li, n1923_li, n1926_li, n1929_li, n1932_li, n1944_li, n1956_li,
    n1968_li, n1980_li, n1992_li, n2004_li, n2016_li, n2019_li, n2028_li,
    n2031_li, n2040_li, n2043_li, n2046_li, n2049_li, n2052_li, n2064_li,
    n2076_li, n2088_li, n2100_li, n2112_li, n2124_li, n2136_li, n2148_li,
    n2151_li, n2160_li, n2163_li, n2172_li, n2175_li, n2178_li, n2181_li,
    n2184_li, n2196_li, n2208_li, n2220_li, n2232_li, n2244_li, n2256_li,
    n2268_li, n2280_li, n2283_li, n2292_li, n2295_li, n2298_li, n2301_li,
    n2304_li, n2316_li, n2319_li, n2322_li, n2325_li, n2328_li, n2331_li,
    n2340_li, n2343_li, n2376_li, n2379_li, n2388_li, n2400_li, n2412_li,
    n2415_li, n2424_li, n2436_li, n2439_li, n2442_li, n2445_li, n2448_li,
    n2451_li, n2460_li, n2463_li, n2496_li, n2499_li, n2508_li, n2520_li,
    n2532_li, n2535_li, n2544_li, n2556_li, n2559_li, n2562_li, n2565_li,
    n2568_li, n2571_li, n2580_li, n2583_li, n2616_li, n2619_li, n2628_li,
    n2640_li, n2652_li, n2655_li, n2664_li, n2676_li, n2679_li, n2682_li,
    n2685_li, n2688_li, n2691_li, n2700_li, n2703_li, n2736_li, n2739_li,
    n2748_li, n2760_li, n2772_li, n2775_li, n2784_li, n2787_li, n2790_li,
    n2793_li, n2796_li, n2799_li, n2802_li, n2805_li, n2808_li, n2820_li,
    n2823_li, n2826_li, n2832_li, n2835_li, n2838_li, n2841_li, n2844_li,
    n2856_li, n2859_li, n2862_li, n2865_li, n2868_li, n2871_li, n2874_li,
    n2877_li, n2880_li, n2883_li, n2886_li, n2889_li, n2892_li, n2895_li,
    n2898_li, n2901_li, n2904_li, n2907_li, n2916_li, n2928_li, n2940_li,
    n2952_li, n2955_li, n2964_li, n2976_li, n2988_li, n2991_li, n3000_li,
    n3003_li, n3012_li, n3015_li, n3024_li, n3027_li, n3036_li, n3039_li,
    n3048_li, n3051_li, n3054_li, n3057_li, n3060_li, n3072_li, n3081_li,
    n3084_li, n3087_li, n3093_li, n3096_li, n3105_li, n3108_li, n3117_li,
    n3120_li, n3123_li, n3126_li, n3129_li, n3132_li, n3135_li, n3138_li,
    n3141_li, n3168_li, n3171_li, n3174_li, n3177_li, n3180_li, n3183_li,
    n3192_li, n3195_li, n3204_li, n3207_li, n3216_li, n3219_li, n3228_li,
    n3231_li, n3240_li, n3243_li, n3252_li, n3255_li, n3258_li, n3264_li,
    n3267_li, n3270_li, n3276_li, n3279_li, n3282_li, n3288_li, n3291_li,
    n3294_li, n4537_i2, n4538_i2, n4710_i2, n4711_i2, n4803_i2, n4804_i2,
    n4843_i2, n4844_i2, n4927_i2, n4928_i2, n4945_i2, n4946_i2, n5009_i2,
    n5178_i2, n5179_i2, n5477_i2, n5478_i2, n5479_i2, n5222_i2, n5223_i2,
    n5553_i2, n5554_i2, G491_i2, n2922_lo_buf_i2, n2946_lo_buf_i2,
    n2970_lo_buf_i2, n2982_lo_buf_i2, n3066_lo_buf_i2, n3078_lo_buf_i2,
    n3102_lo_buf_i2, n3114_lo_buf_i2, G1321_i2, G1033_i2, G1030_i2,
    G1072_i2, G1159_i2, G1152_i2, n2958_lo_buf_i2, n2994_lo_buf_i2,
    n3006_lo_buf_i2, n3030_lo_buf_i2, n3042_lo_buf_i2, n3090_lo_buf_i2,
    G370_i2, G447_i2, G455_i2, G459_i2, G497_i2, G503_i2, G511_i2, G515_i2,
    G1036_i2, G1062_i2, G1067_i2, G1014_i2, G1171_i2, G1166_i2,
    n3018_lo_buf_i2, G766_i2, G451_i2, G463_i2, G467_i2, G475_i2, G479_i2,
    G507_i2, G1017_i2, G1008_i2, G1176_i2, G1144_i2, n2910_lo_buf_i2,
    G471_i2, G2138_i2, G2147_i2, G1148_i2, G1137_i2, G1329_i2, G374_i2,
    G386_i2, G663_i2, G674_i2, G578_i2, G575_i2, G2505_i2, G2508_i2,
    G987_i2, G984_i2, G1862_i2, G1859_i2, G1260_i2, G1865_i2, G2073_i2,
    G1402_i2, G2048_i2, G2276_i2, G366_i2, G2141_i2, G2008_i2, G2011_i2,
    G2150_i2, G2026_i2, G2029_i2, G2023_i2, G2041_i2, G2017_i2, G2020_i2,
    G2035_i2, G2038_i2, G2228_i2, G2231_i2, G2234_i2, G2237_i2, G1904_i2,
    G1907_i2, G1928_i2, G1931_i2, G1893_i2, G1896_i2, G1899_i2, G1937_i2,
    G1940_i2, G1943_i2, G1336_i2, G1996_i2, G1999_i2, G2002_i2, G2005_i2,
    G2014_i2, G2032_i2, G1076_i2, G1002_i2, G998_i2, G1890_i2, G1934_i2,
    G1044_i2, G1039_i2, n1770_lo_buf_i2, G342_i2, G354_i2, G1193_i2,
    n3234_lo_buf_i2, n3246_lo_buf_i2, G783_i2, G786_i2, G792_i2, G795_i2,
    G815_i2, G818_i2, G824_i2, G827_i2, G789_i2, G798_i2, G801_i2, G807_i2,
    G812_i2, G821_i2, G804_i2, G780_i2, G1231_i2, G1572_i2, G1377_i2,
    G1253_i2, G1359_i2, G1258_i2, G1367_i2, G1358_i2, G1366_i2, G2057_i2,
    G2117_i2, G2118_i2, G1254_i2, G1259_i2, G2058_i2, G405_i2, G417_i2,
    G1269_i2, G1275_i2, G1287_i2, G1266_i2, G1272_i2, G1278_i2, G1281_i2,
    G1284_i2, G1290_i2, G1293_i2, G1299_i2, G1305_i2, G1296_i2, G1302_i2,
    G1308_i2, G1311_i2, G811_i2, G810_i2, G1728_i2, G2512_i2, G1114_i2,
    G1113_i2, G1992_i2, G1991_i2, G1426_i2, G1966_i2, G2211_i2, G1509_i2,
    G2153_i2, G2329_i2, G1540_i2, G2167_i2, G2191_i2, G1234_i2, G1132_i2,
    G1129_i2, G2088_i2, G2106_i2, G1314_i2, G636_i2, G647_i2,
    n3186_lo_buf_i2, n3198_lo_buf_i2, n3210_lo_buf_i2, n3222_lo_buf_i2,
    G1225_i2, G1342_i2, G1222_i2, G1228_i2, G1348_i2, G1345_i2, G1351_i2,
    G2242_i2, G2260_i2, G1374_i2, G1537_i2, G301_i2, G313_i2, G2365_i2,
    G2255_i2, G2253_i2, G2395_i2, G2272_i2, G2270_i2, G2245_i2, G2262_i2,
    G2249_i2, G2247_i2, G2266_i2, G2264_i2, G2403_i2, G2401_i2, G2410_i2,
    G2408_i2, G2306_i2, G2305_i2, G2314_i2, G2313_i2, G2303_i2, G2302_i2,
    G2301_i2, G2311_i2, G2310_i2, G2309_i2, G2404_i2, G2411_i2, G2420_i2,
    G2419_i2, G2433_i2, G2432_i2, G402_i2, G403_i2, G1053_i2, G1049_i2,
    G1058_i2, G1364_i2, G1079_i2, G1478_i2, G707_i2, G718_i2, G2417_i2,
    G2414_i2, G2431_i2, G2428_i2, G1653_i2, G2213_i2, G2221_i2, G2250_i2,
    G2267_i2, G1365_i2, G1368_i2, G1371_i2, G2218_i2, G2225_i2,
    n1503_lo_buf_i2, n1863_lo_buf_i2, n1887_lo_buf_i2, n1983_lo_buf_i2,
    n2007_lo_buf_i2, n2115_lo_buf_i2, n2139_lo_buf_i2, n2247_lo_buf_i2,
    n2271_lo_buf_i2, n2919_lo_buf_i2, n2943_lo_buf_i2, n2967_lo_buf_i2,
    n2979_lo_buf_i2, n3063_lo_buf_i2, n3075_lo_buf_i2, n3099_lo_buf_i2,
    n3111_lo_buf_i2, G878_i2, G875_i2, G661_i2, G660_i2, G879_i2, G876_i2,
    G1320_i2, G941_i2, G732_i2, G942_i2, G1493_i2, G1498_i2, G877_i2,
    G874_i2, n1806_lo_buf_i2, n1878_lo_buf_i2, n1938_lo_buf_i2,
    n1998_lo_buf_i2, n2058_lo_buf_i2, n2130_lo_buf_i2, n2190_lo_buf_i2,
    n2262_lo_buf_i2, n2310_lo_buf_i2, n2406_lo_buf_i2, n2430_lo_buf_i2,
    n2526_lo_buf_i2, n2550_lo_buf_i2, n2646_lo_buf_i2, n2670_lo_buf_i2,
    n2766_lo_buf_i2, G603_i2, G614_i2, G1026_i2, G1021_i2, G940_i2,
    G1636_i2, G1684_i2, n2352_lo_buf_i2, n2364_lo_buf_i2, n2472_lo_buf_i2,
    n2484_lo_buf_i2, n2592_lo_buf_i2, n2604_lo_buf_i2, n2712_lo_buf_i2,
    n2724_lo_buf_i2, n3150_lo_buf_i2, n3162_lo_buf_i2;
  assign new_n1576_ = G1;
  assign new_n1578_ = G2;
  assign new_n1580_ = G3;
  assign new_n1582_ = G4;
  assign new_n1584_ = G5;
  assign new_n1586_ = G6;
  assign new_n1588_ = G7;
  assign new_n1590_ = G8;
  assign new_n1592_ = G9;
  assign new_n1594_ = G10;
  assign new_n1596_ = G11;
  assign new_n1598_ = G12;
  assign new_n1600_ = G13;
  assign new_n1602_ = G14;
  assign new_n1604_ = G15;
  assign new_n1606_ = G16;
  assign new_n1608_ = G17;
  assign new_n1610_ = G18;
  assign new_n1612_ = G19;
  assign new_n1614_ = G20;
  assign new_n1616_ = G21;
  assign new_n1618_ = G22;
  assign new_n1620_ = G23;
  assign new_n1622_ = G24;
  assign new_n1624_ = G25;
  assign new_n1626_ = G26;
  assign new_n1628_ = G27;
  assign new_n1630_ = G28;
  assign new_n1632_ = G29;
  assign new_n1634_ = G30;
  assign new_n1636_ = G31;
  assign new_n1638_ = G32;
  assign new_n1640_ = G33;
  assign new_n1642_ = G34;
  assign new_n1644_ = G35;
  assign new_n1646_ = G36;
  assign new_n1648_ = G37;
  assign new_n1650_ = G38;
  assign new_n1652_ = G39;
  assign new_n1654_ = G40;
  assign new_n1656_ = G41;
  assign new_n1658_ = G42;
  assign new_n1660_ = G43;
  assign new_n1662_ = G44;
  assign new_n1664_ = G45;
  assign new_n1666_ = G46;
  assign new_n1668_ = G47;
  assign new_n1670_ = G48;
  assign new_n1672_ = G49;
  assign new_n1674_ = G50;
  assign new_n1676_ = G51;
  assign new_n1678_ = G52;
  assign new_n1680_ = G53;
  assign new_n1682_ = G54;
  assign new_n1684_ = G55;
  assign new_n1686_ = G56;
  assign new_n1688_ = G57;
  assign new_n1690_ = G58;
  assign new_n1692_ = G59;
  assign new_n1694_ = G60;
  assign new_n1696_ = G61;
  assign new_n1698_ = G62;
  assign new_n1700_ = G63;
  assign new_n1702_ = G64;
  assign new_n1704_ = G65;
  assign new_n1706_ = G66;
  assign new_n1708_ = G67;
  assign new_n1710_ = G68;
  assign new_n1712_ = G69;
  assign new_n1714_ = G70;
  assign new_n1716_ = G71;
  assign new_n1718_ = G72;
  assign new_n1720_ = G73;
  assign new_n1722_ = G74;
  assign new_n1724_ = G75;
  assign new_n1726_ = G76;
  assign new_n1728_ = G77;
  assign new_n1730_ = G78;
  assign new_n1732_ = G79;
  assign new_n1734_ = G80;
  assign new_n1736_ = G81;
  assign new_n1738_ = G82;
  assign new_n1740_ = G83;
  assign new_n1742_ = G84;
  assign new_n1744_ = G85;
  assign new_n1746_ = G86;
  assign new_n1748_ = G87;
  assign new_n1750_ = G88;
  assign new_n1752_ = G89;
  assign new_n1754_ = G90;
  assign new_n1756_ = G91;
  assign new_n1758_ = G92;
  assign new_n1760_ = G93;
  assign new_n1762_ = G94;
  assign new_n1764_ = G95;
  assign new_n1766_ = G96;
  assign new_n1768_ = G97;
  assign new_n1770_ = G98;
  assign new_n1772_ = G99;
  assign new_n1774_ = G100;
  assign new_n1776_ = G101;
  assign new_n1778_ = G102;
  assign new_n1780_ = G103;
  assign new_n1782_ = G104;
  assign new_n1784_ = G105;
  assign new_n1786_ = G106;
  assign new_n1788_ = G107;
  assign new_n1790_ = G108;
  assign new_n1792_ = G109;
  assign new_n1794_ = G110;
  assign new_n1796_ = G111;
  assign new_n1798_ = G112;
  assign new_n1800_ = G113;
  assign new_n1802_ = G114;
  assign new_n1804_ = G115;
  assign new_n1806_ = G116;
  assign new_n1808_ = G117;
  assign new_n1810_ = G118;
  assign new_n1812_ = G119;
  assign new_n1814_ = G120;
  assign new_n1816_ = G121;
  assign new_n1818_ = G122;
  assign new_n1820_ = G123;
  assign new_n1822_ = G124;
  assign new_n1824_ = G125;
  assign new_n1826_ = G126;
  assign new_n1828_ = G127;
  assign new_n1830_ = G128;
  assign new_n1832_ = G129;
  assign new_n1834_ = G130;
  assign new_n1836_ = G131;
  assign new_n1838_ = G132;
  assign new_n1840_ = G133;
  assign new_n1842_ = G134;
  assign new_n1844_ = G135;
  assign new_n1846_ = G136;
  assign new_n1848_ = G137;
  assign new_n1850_ = G138;
  assign new_n1852_ = G139;
  assign new_n1854_ = G140;
  assign new_n1856_ = G141;
  assign new_n1858_ = G142;
  assign new_n1860_ = G143;
  assign new_n1862_ = G144;
  assign new_n1864_ = G145;
  assign new_n1866_ = G146;
  assign new_n1868_ = G147;
  assign new_n1870_ = G148;
  assign new_n1872_ = G149;
  assign new_n1874_ = G150;
  assign new_n1876_ = G151;
  assign new_n1878_ = G152;
  assign new_n1880_ = G153;
  assign new_n1882_ = G154;
  assign new_n1884_ = G155;
  assign new_n1886_ = G156;
  assign new_n1888_ = G157;
  assign new_n1890_ = n1416_lo;
  assign new_n1892_ = n1419_lo;
  assign new_n1894_ = n1422_lo;
  assign new_n1896_ = n1425_lo;
  assign new_n1898_ = n1428_lo;
  assign new_n1900_ = n1431_lo;
  assign new_n1902_ = n1434_lo;
  assign new_n1905_ = ~n1437_lo;
  assign new_n1906_ = n1440_lo;
  assign new_n1908_ = n1443_lo;
  assign new_n1910_ = n1446_lo;
  assign new_n1912_ = n1449_lo;
  assign new_n1914_ = n1452_lo;
  assign new_n1916_ = n1455_lo;
  assign new_n1918_ = n1458_lo;
  assign new_n1920_ = n1464_lo;
  assign new_n1922_ = n1467_lo;
  assign new_n1924_ = n1470_lo;
  assign new_n1926_ = n1476_lo;
  assign new_n1928_ = n1479_lo;
  assign new_n1930_ = n1482_lo;
  assign new_n1932_ = n1488_lo;
  assign new_n1934_ = n1491_lo;
  assign new_n1936_ = n1494_lo;
  assign new_n1939_ = ~n1497_lo;
  assign new_n1940_ = n1500_lo;
  assign new_n1942_ = n1512_lo;
  assign new_n1944_ = n1515_lo;
  assign new_n1946_ = n1518_lo;
  assign new_n1949_ = ~n1521_lo;
  assign new_n1950_ = n1524_lo;
  assign new_n1952_ = n1527_lo;
  assign new_n1954_ = n1530_lo;
  assign new_n1956_ = n1533_lo;
  assign new_n1958_ = n1536_lo;
  assign new_n1960_ = n1539_lo;
  assign new_n1962_ = n1542_lo;
  assign new_n1965_ = ~n1545_lo;
  assign new_n1966_ = n1548_lo;
  assign new_n1968_ = n1551_lo;
  assign new_n1970_ = n1554_lo;
  assign new_n1971_ = ~n1554_lo;
  assign new_n1972_ = n1560_lo;
  assign new_n1974_ = n1563_lo;
  assign new_n1976_ = n1566_lo;
  assign new_n1978_ = n1572_lo;
  assign new_n1980_ = n1575_lo;
  assign new_n1982_ = n1578_lo;
  assign new_n1984_ = n1584_lo;
  assign new_n1986_ = n1587_lo;
  assign new_n1988_ = n1590_lo;
  assign new_n1990_ = n1596_lo;
  assign new_n1992_ = n1599_lo;
  assign new_n1994_ = n1602_lo;
  assign new_n1996_ = n1608_lo;
  assign new_n1998_ = n1611_lo;
  assign new_n2000_ = n1614_lo;
  assign new_n2002_ = n1620_lo;
  assign new_n2004_ = n1623_lo;
  assign new_n2006_ = n1626_lo;
  assign new_n2008_ = n1632_lo;
  assign new_n2010_ = n1635_lo;
  assign new_n2012_ = n1638_lo;
  assign new_n2014_ = n1644_lo;
  assign new_n2016_ = n1647_lo;
  assign new_n2018_ = n1650_lo;
  assign new_n2020_ = n1656_lo;
  assign new_n2022_ = n1659_lo;
  assign new_n2024_ = n1662_lo;
  assign new_n2026_ = n1668_lo;
  assign new_n2028_ = n1671_lo;
  assign new_n2030_ = n1674_lo;
  assign new_n2033_ = ~n1677_lo;
  assign new_n2034_ = n1680_lo;
  assign new_n2036_ = n1683_lo;
  assign new_n2038_ = n1686_lo;
  assign new_n2039_ = ~n1686_lo;
  assign new_n2040_ = n1692_lo;
  assign new_n2042_ = n1695_lo;
  assign new_n2044_ = n1698_lo;
  assign new_n2046_ = n1704_lo;
  assign new_n2048_ = n1707_lo;
  assign new_n2050_ = n1710_lo;
  assign new_n2052_ = n1716_lo;
  assign new_n2054_ = n1719_lo;
  assign new_n2056_ = n1722_lo;
  assign new_n2058_ = n1728_lo;
  assign new_n2060_ = n1731_lo;
  assign new_n2062_ = n1734_lo;
  assign new_n2064_ = n1740_lo;
  assign new_n2066_ = n1743_lo;
  assign new_n2068_ = n1746_lo;
  assign new_n2071_ = ~n1749_lo;
  assign new_n2072_ = n1752_lo;
  assign new_n2074_ = n1755_lo;
  assign new_n2076_ = n1758_lo;
  assign new_n2079_ = ~n1761_lo;
  assign new_n2080_ = n1764_lo;
  assign new_n2081_ = ~n1764_lo;
  assign new_n2082_ = n1776_lo;
  assign new_n2084_ = n1779_lo;
  assign new_n2086_ = n1788_lo;
  assign new_n2088_ = n1791_lo;
  assign new_n2090_ = n1794_lo;
  assign new_n2093_ = ~n1797_lo;
  assign new_n2094_ = n1800_lo;
  assign new_n2096_ = n1812_lo;
  assign new_n2098_ = n1824_lo;
  assign new_n2100_ = n1836_lo;
  assign new_n2102_ = n1848_lo;
  assign new_n2104_ = n1860_lo;
  assign new_n2106_ = n1872_lo;
  assign new_n2108_ = n1884_lo;
  assign new_n2110_ = n1896_lo;
  assign new_n2112_ = n1899_lo;
  assign new_n2114_ = n1908_lo;
  assign new_n2116_ = n1911_lo;
  assign new_n2118_ = n1920_lo;
  assign new_n2120_ = n1923_lo;
  assign new_n2122_ = n1926_lo;
  assign new_n2125_ = ~n1929_lo;
  assign new_n2126_ = n1932_lo;
  assign new_n2128_ = n1944_lo;
  assign new_n2130_ = n1956_lo;
  assign new_n2132_ = n1968_lo;
  assign new_n2134_ = n1980_lo;
  assign new_n2136_ = n1992_lo;
  assign new_n2138_ = n2004_lo;
  assign new_n2140_ = n2016_lo;
  assign new_n2142_ = n2019_lo;
  assign new_n2144_ = n2028_lo;
  assign new_n2146_ = n2031_lo;
  assign new_n2148_ = n2040_lo;
  assign new_n2150_ = n2043_lo;
  assign new_n2152_ = n2046_lo;
  assign new_n2155_ = ~n2049_lo;
  assign new_n2156_ = n2052_lo;
  assign new_n2158_ = n2064_lo;
  assign new_n2160_ = n2076_lo;
  assign new_n2162_ = n2088_lo;
  assign new_n2164_ = n2100_lo;
  assign new_n2166_ = n2112_lo;
  assign new_n2168_ = n2124_lo;
  assign new_n2170_ = n2136_lo;
  assign new_n2172_ = n2148_lo;
  assign new_n2174_ = n2151_lo;
  assign new_n2176_ = n2160_lo;
  assign new_n2178_ = n2163_lo;
  assign new_n2180_ = n2172_lo;
  assign new_n2182_ = n2175_lo;
  assign new_n2184_ = n2178_lo;
  assign new_n2187_ = ~n2181_lo;
  assign new_n2188_ = n2184_lo;
  assign new_n2190_ = n2196_lo;
  assign new_n2192_ = n2208_lo;
  assign new_n2194_ = n2220_lo;
  assign new_n2196_ = n2232_lo;
  assign new_n2198_ = n2244_lo;
  assign new_n2200_ = n2256_lo;
  assign new_n2202_ = n2268_lo;
  assign new_n2204_ = n2280_lo;
  assign new_n2206_ = n2283_lo;
  assign new_n2208_ = n2292_lo;
  assign new_n2210_ = n2295_lo;
  assign new_n2212_ = n2298_lo;
  assign new_n2214_ = n2301_lo;
  assign new_n2216_ = n2304_lo;
  assign new_n2218_ = n2316_lo;
  assign new_n2220_ = n2319_lo;
  assign new_n2222_ = n2322_lo;
  assign new_n2225_ = ~n2325_lo;
  assign new_n2226_ = n2328_lo;
  assign new_n2228_ = n2331_lo;
  assign new_n2230_ = n2340_lo;
  assign new_n2232_ = n2343_lo;
  assign new_n2234_ = n2376_lo;
  assign new_n2236_ = n2379_lo;
  assign new_n2238_ = n2388_lo;
  assign new_n2240_ = n2400_lo;
  assign new_n2242_ = n2412_lo;
  assign new_n2244_ = n2415_lo;
  assign new_n2246_ = n2424_lo;
  assign new_n2248_ = n2436_lo;
  assign new_n2250_ = n2439_lo;
  assign new_n2252_ = n2442_lo;
  assign new_n2255_ = ~n2445_lo;
  assign new_n2256_ = n2448_lo;
  assign new_n2258_ = n2451_lo;
  assign new_n2260_ = n2460_lo;
  assign new_n2262_ = n2463_lo;
  assign new_n2264_ = n2496_lo;
  assign new_n2266_ = n2499_lo;
  assign new_n2268_ = n2508_lo;
  assign new_n2270_ = n2520_lo;
  assign new_n2272_ = n2532_lo;
  assign new_n2274_ = n2535_lo;
  assign new_n2276_ = n2544_lo;
  assign new_n2278_ = n2556_lo;
  assign new_n2280_ = n2559_lo;
  assign new_n2282_ = n2562_lo;
  assign new_n2285_ = ~n2565_lo;
  assign new_n2286_ = n2568_lo;
  assign new_n2288_ = n2571_lo;
  assign new_n2290_ = n2580_lo;
  assign new_n2292_ = n2583_lo;
  assign new_n2294_ = n2616_lo;
  assign new_n2296_ = n2619_lo;
  assign new_n2298_ = n2628_lo;
  assign new_n2300_ = n2640_lo;
  assign new_n2302_ = n2652_lo;
  assign new_n2304_ = n2655_lo;
  assign new_n2306_ = n2664_lo;
  assign new_n2308_ = n2676_lo;
  assign new_n2310_ = n2679_lo;
  assign new_n2312_ = n2682_lo;
  assign new_n2315_ = ~n2685_lo;
  assign new_n2316_ = n2688_lo;
  assign new_n2318_ = n2691_lo;
  assign new_n2320_ = n2700_lo;
  assign new_n2322_ = n2703_lo;
  assign new_n2324_ = n2736_lo;
  assign new_n2326_ = n2739_lo;
  assign new_n2328_ = n2748_lo;
  assign new_n2330_ = n2760_lo;
  assign new_n2332_ = n2772_lo;
  assign new_n2334_ = n2775_lo;
  assign new_n2336_ = n2784_lo;
  assign new_n2338_ = n2787_lo;
  assign new_n2340_ = n2790_lo;
  assign new_n2342_ = n2793_lo;
  assign new_n2343_ = ~n2793_lo;
  assign new_n2344_ = n2796_lo;
  assign new_n2346_ = n2799_lo;
  assign new_n2348_ = n2802_lo;
  assign new_n2351_ = ~n2805_lo;
  assign new_n2352_ = n2808_lo;
  assign new_n2353_ = ~n2808_lo;
  assign new_n2354_ = n2820_lo;
  assign new_n2356_ = n2823_lo;
  assign new_n2358_ = n2826_lo;
  assign new_n2359_ = ~n2826_lo;
  assign new_n2360_ = n2832_lo;
  assign new_n2362_ = n2835_lo;
  assign new_n2364_ = n2838_lo;
  assign new_n2366_ = n2841_lo;
  assign new_n2367_ = ~n2841_lo;
  assign new_n2368_ = n2844_lo;
  assign new_n2369_ = ~n2844_lo;
  assign new_n2370_ = n2856_lo;
  assign new_n2372_ = n2859_lo;
  assign new_n2374_ = n2862_lo;
  assign new_n2376_ = n2865_lo;
  assign new_n2377_ = ~n2865_lo;
  assign new_n2378_ = n2868_lo;
  assign new_n2380_ = n2871_lo;
  assign new_n2382_ = n2874_lo;
  assign new_n2384_ = n2877_lo;
  assign new_n2385_ = ~n2877_lo;
  assign new_n2386_ = n2880_lo;
  assign new_n2388_ = n2883_lo;
  assign new_n2390_ = n2886_lo;
  assign new_n2392_ = n2889_lo;
  assign new_n2393_ = ~n2889_lo;
  assign new_n2394_ = n2892_lo;
  assign new_n2396_ = n2895_lo;
  assign new_n2398_ = n2898_lo;
  assign new_n2401_ = ~n2901_lo;
  assign new_n2402_ = n2904_lo;
  assign new_n2404_ = n2907_lo;
  assign new_n2406_ = n2916_lo;
  assign new_n2408_ = n2928_lo;
  assign new_n2410_ = n2940_lo;
  assign new_n2412_ = n2952_lo;
  assign new_n2414_ = n2955_lo;
  assign new_n2415_ = ~n2955_lo;
  assign new_n2416_ = n2964_lo;
  assign new_n2418_ = n2976_lo;
  assign new_n2420_ = n2988_lo;
  assign new_n2422_ = n2991_lo;
  assign new_n2424_ = n3000_lo;
  assign new_n2426_ = n3003_lo;
  assign new_n2428_ = n3012_lo;
  assign new_n2430_ = n3015_lo;
  assign new_n2431_ = ~n3015_lo;
  assign new_n2432_ = n3024_lo;
  assign new_n2434_ = n3027_lo;
  assign new_n2435_ = ~n3027_lo;
  assign new_n2436_ = n3036_lo;
  assign new_n2438_ = n3039_lo;
  assign new_n2439_ = ~n3039_lo;
  assign new_n2440_ = n3048_lo;
  assign new_n2442_ = n3051_lo;
  assign new_n2444_ = n3054_lo;
  assign new_n2447_ = ~n3057_lo;
  assign new_n2448_ = n3060_lo;
  assign new_n2450_ = n3072_lo;
  assign new_n2453_ = ~n3081_lo;
  assign new_n2454_ = n3084_lo;
  assign new_n2456_ = n3087_lo;
  assign new_n2457_ = ~n3087_lo;
  assign new_n2459_ = ~n3093_lo;
  assign new_n2460_ = n3096_lo;
  assign new_n2463_ = ~n3105_lo;
  assign new_n2464_ = n3108_lo;
  assign new_n2467_ = ~n3117_lo;
  assign new_n2468_ = n3120_lo;
  assign new_n2470_ = n3123_lo;
  assign new_n2472_ = n3126_lo;
  assign new_n2474_ = n3129_lo;
  assign new_n2475_ = ~n3129_lo;
  assign new_n2476_ = n3132_lo;
  assign new_n2478_ = n3135_lo;
  assign new_n2480_ = n3138_lo;
  assign new_n2482_ = n3141_lo;
  assign new_n2483_ = ~n3141_lo;
  assign new_n2484_ = n3168_lo;
  assign new_n2486_ = n3171_lo;
  assign new_n2488_ = n3174_lo;
  assign new_n2490_ = n3177_lo;
  assign new_n2491_ = ~n3177_lo;
  assign new_n2492_ = n3180_lo;
  assign new_n2494_ = n3183_lo;
  assign new_n2496_ = n3192_lo;
  assign new_n2498_ = n3195_lo;
  assign new_n2500_ = n3204_lo;
  assign new_n2502_ = n3207_lo;
  assign new_n2504_ = n3216_lo;
  assign new_n2506_ = n3219_lo;
  assign new_n2508_ = n3228_lo;
  assign new_n2510_ = n3231_lo;
  assign new_n2512_ = n3240_lo;
  assign new_n2514_ = n3243_lo;
  assign new_n2516_ = n3252_lo;
  assign new_n2518_ = n3255_lo;
  assign new_n2520_ = n3258_lo;
  assign new_n2521_ = ~n3258_lo;
  assign new_n2522_ = n3264_lo;
  assign new_n2524_ = n3267_lo;
  assign new_n2526_ = n3270_lo;
  assign new_n2527_ = ~n3270_lo;
  assign new_n2528_ = n3276_lo;
  assign new_n2530_ = n3279_lo;
  assign new_n2532_ = n3282_lo;
  assign new_n2533_ = ~n3282_lo;
  assign new_n2534_ = n3288_lo;
  assign new_n2536_ = n3291_lo;
  assign new_n2538_ = n3294_lo;
  assign new_n2539_ = ~n3294_lo;
  assign new_n2541_ = ~n4537_o2;
  assign new_n2543_ = ~n4538_o2;
  assign new_n2545_ = ~n4710_o2;
  assign new_n2547_ = ~n4711_o2;
  assign new_n2548_ = n1211_inv;
  assign new_n2550_ = n1214_inv;
  assign new_n2552_ = n1217_inv;
  assign new_n2554_ = n1220_inv;
  assign new_n2557_ = ~n4927_o2;
  assign new_n2558_ = n4928_o2;
  assign new_n2559_ = ~n4928_o2;
  assign new_n2560_ = n1229_inv;
  assign new_n2562_ = n1232_inv;
  assign new_n2564_ = n1235_inv;
  assign new_n2566_ = n5178_o2;
  assign new_n2567_ = ~n5178_o2;
  assign new_n2568_ = n5179_o2;
  assign new_n2569_ = ~n5179_o2;
  assign new_n2570_ = n5477_o2;
  assign new_n2571_ = ~n5477_o2;
  assign new_n2573_ = ~n5478_o2;
  assign new_n2574_ = n5479_o2;
  assign new_n2575_ = ~n5479_o2;
  assign new_n2576_ = n5222_o2;
  assign new_n2577_ = ~n5222_o2;
  assign new_n2578_ = n5223_o2;
  assign new_n2580_ = n5553_o2;
  assign new_n2582_ = n5554_o2;
  assign new_n2584_ = G491_o2;
  assign new_n2586_ = n2922_lo_buf_o2;
  assign new_n2587_ = ~n2922_lo_buf_o2;
  assign new_n2588_ = n2946_lo_buf_o2;
  assign new_n2589_ = ~n2946_lo_buf_o2;
  assign new_n2590_ = n2970_lo_buf_o2;
  assign new_n2591_ = ~n2970_lo_buf_o2;
  assign new_n2592_ = n2982_lo_buf_o2;
  assign new_n2593_ = ~n2982_lo_buf_o2;
  assign new_n2594_ = n3066_lo_buf_o2;
  assign new_n2595_ = ~n3066_lo_buf_o2;
  assign new_n2596_ = n3078_lo_buf_o2;
  assign new_n2597_ = ~n3078_lo_buf_o2;
  assign new_n2598_ = n3102_lo_buf_o2;
  assign new_n2599_ = ~n3102_lo_buf_o2;
  assign new_n2600_ = n3114_lo_buf_o2;
  assign new_n2601_ = ~n3114_lo_buf_o2;
  assign new_n2602_ = G1321_o2;
  assign new_n2603_ = ~G1321_o2;
  assign new_n2604_ = G1033_o2;
  assign new_n2606_ = G1030_o2;
  assign new_n2608_ = G1072_o2;
  assign new_n2610_ = n1304_inv;
  assign new_n2612_ = n1307_inv;
  assign new_n2614_ = n2958_lo_buf_o2;
  assign new_n2615_ = ~n2958_lo_buf_o2;
  assign new_n2616_ = n2994_lo_buf_o2;
  assign new_n2617_ = ~n2994_lo_buf_o2;
  assign new_n2618_ = n3006_lo_buf_o2;
  assign new_n2619_ = ~n3006_lo_buf_o2;
  assign new_n2620_ = n3030_lo_buf_o2;
  assign new_n2621_ = ~n3030_lo_buf_o2;
  assign new_n2622_ = n3042_lo_buf_o2;
  assign new_n2623_ = ~n3042_lo_buf_o2;
  assign new_n2624_ = n3090_lo_buf_o2;
  assign new_n2625_ = ~n3090_lo_buf_o2;
  assign new_n2626_ = n1328_inv;
  assign new_n2628_ = n1331_inv;
  assign new_n2630_ = n1334_inv;
  assign new_n2632_ = n1337_inv;
  assign new_n2634_ = n1340_inv;
  assign new_n2636_ = n1343_inv;
  assign new_n2638_ = n1346_inv;
  assign new_n2640_ = n1349_inv;
  assign new_n2642_ = G1036_o2;
  assign new_n2644_ = G1062_o2;
  assign new_n2646_ = G1067_o2;
  assign new_n2648_ = G1014_o2;
  assign new_n2650_ = n1364_inv;
  assign new_n2652_ = n1367_inv;
  assign new_n2654_ = n3018_lo_buf_o2;
  assign new_n2655_ = ~n3018_lo_buf_o2;
  assign new_n2657_ = ~G766_o2;
  assign new_n2658_ = n1376_inv;
  assign new_n2660_ = n1379_inv;
  assign new_n2662_ = n1382_inv;
  assign new_n2664_ = n1385_inv;
  assign new_n2666_ = n1388_inv;
  assign new_n2668_ = n1391_inv;
  assign new_n2670_ = G1017_o2;
  assign new_n2672_ = G1008_o2;
  assign new_n2673_ = ~G1008_o2;
  assign new_n2674_ = n1400_inv;
  assign new_n2676_ = n1403_inv;
  assign new_n2678_ = n2910_lo_buf_o2;
  assign new_n2679_ = ~n2910_lo_buf_o2;
  assign new_n2680_ = n1409_inv;
  assign new_n2682_ = G2138_o2;
  assign new_n2683_ = ~G2138_o2;
  assign new_n2684_ = G2147_o2;
  assign new_n2685_ = ~G2147_o2;
  assign new_n2686_ = n1418_inv;
  assign new_n2688_ = G1137_o2;
  assign new_n2689_ = ~G1137_o2;
  assign new_n2690_ = G1329_o2;
  assign new_n2691_ = ~G1329_o2;
  assign new_n2692_ = G374_o2;
  assign new_n2693_ = ~G374_o2;
  assign new_n2694_ = G386_o2;
  assign new_n2695_ = ~G386_o2;
  assign new_n2696_ = G663_o2;
  assign new_n2697_ = ~G663_o2;
  assign new_n2698_ = G674_o2;
  assign new_n2699_ = ~G674_o2;
  assign new_n2700_ = G578_o2;
  assign new_n2701_ = ~G578_o2;
  assign new_n2702_ = G575_o2;
  assign new_n2703_ = ~G575_o2;
  assign new_n2705_ = ~G2505_o2;
  assign new_n2706_ = n1448_inv;
  assign new_n2707_ = ~n1448_inv;
  assign new_n2708_ = G987_o2;
  assign new_n2709_ = ~G987_o2;
  assign new_n2710_ = G984_o2;
  assign new_n2711_ = ~G984_o2;
  assign new_n2712_ = G1862_o2;
  assign new_n2713_ = ~G1862_o2;
  assign new_n2714_ = G1859_o2;
  assign new_n2715_ = ~G1859_o2;
  assign new_n2717_ = ~G1260_o2;
  assign new_n2718_ = G1865_o2;
  assign new_n2721_ = ~G2073_o2;
  assign new_n2722_ = G1402_o2;
  assign new_n2725_ = ~G2048_o2;
  assign new_n2726_ = G2276_o2;
  assign new_n2728_ = n1481_inv;
  assign new_n2730_ = G2141_o2;
  assign new_n2731_ = ~G2141_o2;
  assign new_n2732_ = G2008_o2;
  assign new_n2733_ = ~G2008_o2;
  assign new_n2734_ = G2011_o2;
  assign new_n2735_ = ~G2011_o2;
  assign new_n2736_ = G2150_o2;
  assign new_n2737_ = ~G2150_o2;
  assign new_n2738_ = G2026_o2;
  assign new_n2739_ = ~G2026_o2;
  assign new_n2740_ = G2029_o2;
  assign new_n2741_ = ~G2029_o2;
  assign new_n2742_ = G2023_o2;
  assign new_n2744_ = G2041_o2;
  assign new_n2746_ = G2017_o2;
  assign new_n2748_ = G2020_o2;
  assign new_n2750_ = G2035_o2;
  assign new_n2752_ = G2038_o2;
  assign new_n2754_ = G2228_o2;
  assign new_n2755_ = ~G2228_o2;
  assign new_n2756_ = G2231_o2;
  assign new_n2757_ = ~G2231_o2;
  assign new_n2758_ = G2234_o2;
  assign new_n2759_ = ~G2234_o2;
  assign new_n2760_ = G2237_o2;
  assign new_n2761_ = ~G2237_o2;
  assign new_n2762_ = G1904_o2;
  assign new_n2763_ = ~G1904_o2;
  assign new_n2764_ = G1907_o2;
  assign new_n2765_ = ~G1907_o2;
  assign new_n2766_ = G1928_o2;
  assign new_n2767_ = ~G1928_o2;
  assign new_n2768_ = G1931_o2;
  assign new_n2769_ = ~G1931_o2;
  assign new_n2771_ = ~G1893_o2;
  assign new_n2773_ = ~G1896_o2;
  assign new_n2775_ = ~G1899_o2;
  assign new_n2777_ = ~G1937_o2;
  assign new_n2779_ = ~G1940_o2;
  assign new_n2781_ = ~G1943_o2;
  assign new_n2782_ = G1336_o2;
  assign new_n2783_ = ~G1336_o2;
  assign new_n2784_ = G1996_o2;
  assign new_n2785_ = ~G1996_o2;
  assign new_n2786_ = G1999_o2;
  assign new_n2787_ = ~G1999_o2;
  assign new_n2788_ = G2002_o2;
  assign new_n2789_ = ~G2002_o2;
  assign new_n2790_ = G2005_o2;
  assign new_n2791_ = ~G2005_o2;
  assign new_n2792_ = G2014_o2;
  assign new_n2794_ = G2032_o2;
  assign new_n2796_ = G1076_o2;
  assign new_n2798_ = G1002_o2;
  assign new_n2799_ = ~G1002_o2;
  assign new_n2800_ = G998_o2;
  assign new_n2803_ = ~G1890_o2;
  assign new_n2805_ = ~G1934_o2;
  assign new_n2806_ = G1044_o2;
  assign new_n2808_ = G1039_o2;
  assign new_n2810_ = n1770_lo_buf_o2;
  assign new_n2811_ = ~n1770_lo_buf_o2;
  assign new_n2813_ = ~G342_o2;
  assign new_n2815_ = ~G354_o2;
  assign new_n2816_ = G1193_o2;
  assign new_n2817_ = ~G1193_o2;
  assign new_n2818_ = n3234_lo_buf_o2;
  assign new_n2819_ = ~n3234_lo_buf_o2;
  assign new_n2820_ = n3246_lo_buf_o2;
  assign new_n2821_ = ~n3246_lo_buf_o2;
  assign new_n2822_ = G783_o2;
  assign new_n2823_ = ~G783_o2;
  assign new_n2824_ = G786_o2;
  assign new_n2825_ = ~G786_o2;
  assign new_n2826_ = G792_o2;
  assign new_n2827_ = ~G792_o2;
  assign new_n2828_ = G795_o2;
  assign new_n2829_ = ~G795_o2;
  assign new_n2830_ = G815_o2;
  assign new_n2831_ = ~G815_o2;
  assign new_n2832_ = G818_o2;
  assign new_n2833_ = ~G818_o2;
  assign new_n2834_ = G824_o2;
  assign new_n2835_ = ~G824_o2;
  assign new_n2836_ = G827_o2;
  assign new_n2837_ = ~G827_o2;
  assign new_n2838_ = G789_o2;
  assign new_n2839_ = ~G789_o2;
  assign new_n2840_ = G798_o2;
  assign new_n2841_ = ~G798_o2;
  assign new_n2842_ = G801_o2;
  assign new_n2843_ = ~G801_o2;
  assign new_n2844_ = G807_o2;
  assign new_n2845_ = ~G807_o2;
  assign new_n2846_ = G812_o2;
  assign new_n2847_ = ~G812_o2;
  assign new_n2848_ = G821_o2;
  assign new_n2849_ = ~G821_o2;
  assign new_n2850_ = G804_o2;
  assign new_n2851_ = ~G804_o2;
  assign new_n2852_ = G780_o2;
  assign new_n2853_ = ~G780_o2;
  assign new_n2854_ = G1231_o2;
  assign new_n2855_ = ~G1231_o2;
  assign new_n2856_ = G1572_o2;
  assign new_n2857_ = ~G1572_o2;
  assign new_n2858_ = G1377_o2;
  assign new_n2859_ = ~G1377_o2;
  assign new_n2860_ = G1253_o2;
  assign new_n2861_ = ~G1253_o2;
  assign new_n2862_ = G1359_o2;
  assign new_n2863_ = ~G1359_o2;
  assign new_n2864_ = G1258_o2;
  assign new_n2865_ = ~G1258_o2;
  assign new_n2866_ = G1367_o2;
  assign new_n2867_ = ~G1367_o2;
  assign new_n2868_ = G1358_o2;
  assign new_n2869_ = ~G1358_o2;
  assign new_n2870_ = G1366_o2;
  assign new_n2871_ = ~G1366_o2;
  assign new_n2872_ = G2057_o2;
  assign new_n2873_ = ~G2057_o2;
  assign new_n2874_ = G2117_o2;
  assign new_n2875_ = ~G2117_o2;
  assign new_n2876_ = G2118_o2;
  assign new_n2877_ = ~G2118_o2;
  assign new_n2878_ = G1254_o2;
  assign new_n2879_ = ~G1254_o2;
  assign new_n2880_ = G1259_o2;
  assign new_n2881_ = ~G1259_o2;
  assign new_n2882_ = G2058_o2;
  assign new_n2883_ = ~G2058_o2;
  assign new_n2885_ = ~G405_o2;
  assign new_n2887_ = ~G417_o2;
  assign new_n2888_ = G1269_o2;
  assign new_n2889_ = ~G1269_o2;
  assign new_n2890_ = G1275_o2;
  assign new_n2891_ = ~G1275_o2;
  assign new_n2892_ = G1287_o2;
  assign new_n2893_ = ~G1287_o2;
  assign new_n2894_ = G1266_o2;
  assign new_n2895_ = ~G1266_o2;
  assign new_n2896_ = G1272_o2;
  assign new_n2897_ = ~G1272_o2;
  assign new_n2898_ = G1278_o2;
  assign new_n2899_ = ~G1278_o2;
  assign new_n2900_ = G1281_o2;
  assign new_n2901_ = ~G1281_o2;
  assign new_n2902_ = G1284_o2;
  assign new_n2903_ = ~G1284_o2;
  assign new_n2904_ = G1290_o2;
  assign new_n2905_ = ~G1290_o2;
  assign new_n2906_ = G1293_o2;
  assign new_n2907_ = ~G1293_o2;
  assign new_n2908_ = G1299_o2;
  assign new_n2909_ = ~G1299_o2;
  assign new_n2910_ = G1305_o2;
  assign new_n2911_ = ~G1305_o2;
  assign new_n2912_ = G1296_o2;
  assign new_n2913_ = ~G1296_o2;
  assign new_n2914_ = G1302_o2;
  assign new_n2915_ = ~G1302_o2;
  assign new_n2916_ = G1308_o2;
  assign new_n2917_ = ~G1308_o2;
  assign new_n2918_ = G1311_o2;
  assign new_n2919_ = ~G1311_o2;
  assign new_n2920_ = G811_o2;
  assign new_n2921_ = ~G811_o2;
  assign new_n2922_ = G810_o2;
  assign new_n2923_ = ~G810_o2;
  assign new_n2924_ = G1728_o2;
  assign new_n2925_ = ~G1728_o2;
  assign new_n2926_ = G2512_o2;
  assign new_n2928_ = G1114_o2;
  assign new_n2929_ = ~G1114_o2;
  assign new_n2930_ = G1113_o2;
  assign new_n2931_ = ~G1113_o2;
  assign new_n2932_ = G1992_o2;
  assign new_n2933_ = ~G1992_o2;
  assign new_n2934_ = G1991_o2;
  assign new_n2935_ = ~G1991_o2;
  assign new_n2936_ = G1426_o2;
  assign new_n2939_ = ~G1966_o2;
  assign new_n2940_ = G2211_o2;
  assign new_n2943_ = ~G1509_o2;
  assign new_n2944_ = G2153_o2;
  assign new_n2947_ = ~G2329_o2;
  assign new_n2948_ = G1540_o2;
  assign new_n2949_ = ~G1540_o2;
  assign new_n2951_ = ~G2167_o2;
  assign new_n2953_ = ~G2191_o2;
  assign new_n2954_ = G1234_o2;
  assign new_n2955_ = ~G1234_o2;
  assign new_n2956_ = G1132_o2;
  assign new_n2957_ = ~G1132_o2;
  assign new_n2958_ = G1129_o2;
  assign new_n2959_ = ~G1129_o2;
  assign new_n2960_ = G2088_o2;
  assign new_n2962_ = G2106_o2;
  assign new_n2964_ = G1314_o2;
  assign new_n2965_ = ~G1314_o2;
  assign new_n2966_ = G636_o2;
  assign new_n2968_ = G647_o2;
  assign new_n2970_ = n3186_lo_buf_o2;
  assign new_n2971_ = ~n3186_lo_buf_o2;
  assign new_n2972_ = n3198_lo_buf_o2;
  assign new_n2973_ = ~n3198_lo_buf_o2;
  assign new_n2974_ = n3210_lo_buf_o2;
  assign new_n2975_ = ~n3210_lo_buf_o2;
  assign new_n2976_ = n3222_lo_buf_o2;
  assign new_n2977_ = ~n3222_lo_buf_o2;
  assign new_n2978_ = G1225_o2;
  assign new_n2979_ = ~G1225_o2;
  assign new_n2980_ = G1342_o2;
  assign new_n2981_ = ~G1342_o2;
  assign new_n2982_ = G1222_o2;
  assign new_n2983_ = ~G1222_o2;
  assign new_n2984_ = G1228_o2;
  assign new_n2985_ = ~G1228_o2;
  assign new_n2986_ = G1348_o2;
  assign new_n2987_ = ~G1348_o2;
  assign new_n2988_ = G1345_o2;
  assign new_n2989_ = ~G1345_o2;
  assign new_n2990_ = G1351_o2;
  assign new_n2991_ = ~G1351_o2;
  assign new_n2992_ = G2242_o2;
  assign new_n2993_ = ~G2242_o2;
  assign new_n2994_ = G2260_o2;
  assign new_n2995_ = ~G2260_o2;
  assign new_n2996_ = G1374_o2;
  assign new_n2997_ = ~G1374_o2;
  assign new_n2998_ = G1537_o2;
  assign new_n2999_ = ~G1537_o2;
  assign new_n3000_ = G301_o2;
  assign new_n3001_ = ~G301_o2;
  assign new_n3002_ = G313_o2;
  assign new_n3003_ = ~G313_o2;
  assign new_n3004_ = G2365_o2;
  assign new_n3005_ = ~G2365_o2;
  assign new_n3006_ = G2255_o2;
  assign new_n3007_ = ~G2255_o2;
  assign new_n3008_ = G2253_o2;
  assign new_n3009_ = ~G2253_o2;
  assign new_n3010_ = G2395_o2;
  assign new_n3011_ = ~G2395_o2;
  assign new_n3012_ = G2272_o2;
  assign new_n3013_ = ~G2272_o2;
  assign new_n3014_ = G2270_o2;
  assign new_n3015_ = ~G2270_o2;
  assign new_n3017_ = ~G2245_o2;
  assign new_n3019_ = ~G2262_o2;
  assign new_n3021_ = ~G2249_o2;
  assign new_n3023_ = ~G2247_o2;
  assign new_n3025_ = ~G2266_o2;
  assign new_n3027_ = ~G2264_o2;
  assign new_n3028_ = G2403_o2;
  assign new_n3029_ = ~G2403_o2;
  assign new_n3030_ = G2401_o2;
  assign new_n3031_ = ~G2401_o2;
  assign new_n3032_ = G2410_o2;
  assign new_n3033_ = ~G2410_o2;
  assign new_n3034_ = G2408_o2;
  assign new_n3035_ = ~G2408_o2;
  assign new_n3036_ = G2306_o2;
  assign new_n3037_ = ~G2306_o2;
  assign new_n3038_ = G2305_o2;
  assign new_n3039_ = ~G2305_o2;
  assign new_n3040_ = G2314_o2;
  assign new_n3041_ = ~G2314_o2;
  assign new_n3042_ = G2313_o2;
  assign new_n3043_ = ~G2313_o2;
  assign new_n3044_ = G2303_o2;
  assign new_n3046_ = G2302_o2;
  assign new_n3048_ = G2301_o2;
  assign new_n3050_ = G2311_o2;
  assign new_n3052_ = G2310_o2;
  assign new_n3054_ = G2309_o2;
  assign new_n3056_ = G2404_o2;
  assign new_n3057_ = ~G2404_o2;
  assign new_n3058_ = G2411_o2;
  assign new_n3059_ = ~G2411_o2;
  assign new_n3060_ = G2420_o2;
  assign new_n3061_ = ~G2420_o2;
  assign new_n3062_ = G2419_o2;
  assign new_n3063_ = ~G2419_o2;
  assign new_n3064_ = G2433_o2;
  assign new_n3065_ = ~G2433_o2;
  assign new_n3066_ = G2432_o2;
  assign new_n3067_ = ~G2432_o2;
  assign new_n3068_ = G402_o2;
  assign new_n3069_ = ~G402_o2;
  assign new_n3070_ = G403_o2;
  assign new_n3071_ = ~G403_o2;
  assign new_n3072_ = G1053_o2;
  assign new_n3073_ = ~G1053_o2;
  assign new_n3074_ = G1049_o2;
  assign new_n3075_ = ~G1049_o2;
  assign new_n3076_ = n2003_inv;
  assign new_n3077_ = ~n2003_inv;
  assign new_n3078_ = G1364_o2;
  assign new_n3079_ = ~G1364_o2;
  assign new_n3080_ = G1079_o2;
  assign new_n3081_ = ~G1079_o2;
  assign new_n3082_ = G1478_o2;
  assign new_n3083_ = ~G1478_o2;
  assign new_n3084_ = G707_o2;
  assign new_n3086_ = G718_o2;
  assign new_n3088_ = G2417_o2;
  assign new_n3089_ = ~G2417_o2;
  assign new_n3090_ = G2414_o2;
  assign new_n3091_ = ~G2414_o2;
  assign new_n3092_ = G2431_o2;
  assign new_n3093_ = ~G2431_o2;
  assign new_n3094_ = G2428_o2;
  assign new_n3095_ = ~G2428_o2;
  assign new_n3096_ = G1653_o2;
  assign new_n3097_ = ~G1653_o2;
  assign new_n3098_ = G2213_o2;
  assign new_n3099_ = ~G2213_o2;
  assign new_n3100_ = G2221_o2;
  assign new_n3101_ = ~G2221_o2;
  assign new_n3102_ = G2250_o2;
  assign new_n3104_ = G2267_o2;
  assign new_n3106_ = G1365_o2;
  assign new_n3107_ = ~G1365_o2;
  assign new_n3108_ = G1368_o2;
  assign new_n3109_ = ~G1368_o2;
  assign new_n3110_ = G1371_o2;
  assign new_n3111_ = ~G1371_o2;
  assign new_n3113_ = ~G2218_o2;
  assign new_n3115_ = ~G2225_o2;
  assign new_n3117_ = ~n1503_lo_buf_o2;
  assign new_n3118_ = n1863_lo_buf_o2;
  assign new_n3119_ = ~n1863_lo_buf_o2;
  assign new_n3120_ = n1887_lo_buf_o2;
  assign new_n3121_ = ~n1887_lo_buf_o2;
  assign new_n3122_ = n1983_lo_buf_o2;
  assign new_n3123_ = ~n1983_lo_buf_o2;
  assign new_n3124_ = n2007_lo_buf_o2;
  assign new_n3125_ = ~n2007_lo_buf_o2;
  assign new_n3126_ = n2115_lo_buf_o2;
  assign new_n3127_ = ~n2115_lo_buf_o2;
  assign new_n3128_ = n2139_lo_buf_o2;
  assign new_n3129_ = ~n2139_lo_buf_o2;
  assign new_n3130_ = n2247_lo_buf_o2;
  assign new_n3131_ = ~n2247_lo_buf_o2;
  assign new_n3132_ = n2271_lo_buf_o2;
  assign new_n3133_ = ~n2271_lo_buf_o2;
  assign new_n3134_ = n2919_lo_buf_o2;
  assign new_n3135_ = ~n2919_lo_buf_o2;
  assign new_n3136_ = n2943_lo_buf_o2;
  assign new_n3137_ = ~n2943_lo_buf_o2;
  assign new_n3138_ = n2967_lo_buf_o2;
  assign new_n3140_ = n2979_lo_buf_o2;
  assign new_n3142_ = n3063_lo_buf_o2;
  assign new_n3143_ = ~n3063_lo_buf_o2;
  assign new_n3144_ = n3075_lo_buf_o2;
  assign new_n3145_ = ~n3075_lo_buf_o2;
  assign new_n3146_ = n3099_lo_buf_o2;
  assign new_n3148_ = n3111_lo_buf_o2;
  assign new_n3150_ = G878_o2;
  assign new_n3152_ = G875_o2;
  assign new_n3154_ = G661_o2;
  assign new_n3156_ = G660_o2;
  assign new_n3158_ = G879_o2;
  assign new_n3160_ = G876_o2;
  assign new_n3162_ = G1320_o2;
  assign new_n3163_ = ~G1320_o2;
  assign new_n3164_ = G941_o2;
  assign new_n3166_ = G732_o2;
  assign new_n3168_ = G942_o2;
  assign new_n3170_ = G1493_o2;
  assign new_n3171_ = ~G1493_o2;
  assign new_n3172_ = G1498_o2;
  assign new_n3173_ = ~G1498_o2;
  assign new_n3174_ = G877_o2;
  assign new_n3176_ = G874_o2;
  assign new_n3178_ = n1806_lo_buf_o2;
  assign new_n3180_ = n1878_lo_buf_o2;
  assign new_n3181_ = ~n1878_lo_buf_o2;
  assign new_n3182_ = n1938_lo_buf_o2;
  assign new_n3184_ = n1998_lo_buf_o2;
  assign new_n3185_ = ~n1998_lo_buf_o2;
  assign new_n3186_ = n2058_lo_buf_o2;
  assign new_n3188_ = n2130_lo_buf_o2;
  assign new_n3189_ = ~n2130_lo_buf_o2;
  assign new_n3190_ = n2190_lo_buf_o2;
  assign new_n3192_ = n2262_lo_buf_o2;
  assign new_n3193_ = ~n2262_lo_buf_o2;
  assign new_n3194_ = n2310_lo_buf_o2;
  assign new_n3196_ = n2406_lo_buf_o2;
  assign new_n3198_ = n2430_lo_buf_o2;
  assign new_n3200_ = n2526_lo_buf_o2;
  assign new_n3202_ = n2550_lo_buf_o2;
  assign new_n3204_ = n2646_lo_buf_o2;
  assign new_n3206_ = n2670_lo_buf_o2;
  assign new_n3208_ = n2766_lo_buf_o2;
  assign new_n3210_ = G603_o2;
  assign new_n3211_ = ~G603_o2;
  assign new_n3212_ = G614_o2;
  assign new_n3213_ = ~G614_o2;
  assign new_n3214_ = G1026_o2;
  assign new_n3216_ = G1021_o2;
  assign new_n3218_ = G940_o2;
  assign new_n3220_ = G1636_o2;
  assign new_n3221_ = ~G1636_o2;
  assign new_n3222_ = G1684_o2;
  assign new_n3223_ = ~G1684_o2;
  assign new_n3224_ = n2352_lo_buf_o2;
  assign new_n3227_ = ~n2364_lo_buf_o2;
  assign new_n3228_ = n2472_lo_buf_o2;
  assign new_n3231_ = ~n2484_lo_buf_o2;
  assign new_n3232_ = n2592_lo_buf_o2;
  assign new_n3235_ = ~n2604_lo_buf_o2;
  assign new_n3236_ = n2712_lo_buf_o2;
  assign new_n3239_ = ~n2724_lo_buf_o2;
  assign new_n3240_ = n3150_lo_buf_o2;
  assign new_n3241_ = ~n3150_lo_buf_o2;
  assign new_n3242_ = n3162_lo_buf_o2;
  assign new_n3243_ = ~n3162_lo_buf_o2;
  assign new_n3244_ = new_n2467_ | new_n2463_;
  assign new_n3245_ = new_n3244_ | new_n2459_;
  assign new_n3246_ = new_n3245_ | new_n2453_;
  assign new_n3247_ = new_n1965_ | new_n1905_;
  assign new_n3248_ = new_n3247_ | new_n5047_;
  assign new_n3249_ = new_n5049_ & new_n2214_;
  assign new_n3250_ = new_n5047_ | new_n1939_;
  assign new_n3251_ = new_n5052_ | new_n2367_;
  assign new_n3252_ = new_n5052_ | new_n2491_;
  assign new_n3253_ = new_n5053_ | new_n5054_;
  assign new_n3254_ = new_n3253_ | new_n5055_;
  assign new_n3255_ = new_n3254_ | new_n5056_;
  assign new_n3256_ = new_n5057_ | new_n5058_;
  assign new_n3257_ = new_n3256_ | new_n5059_;
  assign new_n3258_ = new_n3257_ | new_n5060_;
  assign new_n3259_ = new_n5061_ | new_n5062_;
  assign new_n3260_ = new_n5061_ & new_n2490_;
  assign new_n3261_ = new_n5062_ & new_n2366_;
  assign new_n3262_ = new_n3261_ | new_n3260_;
  assign new_n3263_ = new_n2566_ & new_n5064_;
  assign new_n3264_ = new_n3263_ | new_n5066_;
  assign new_n3265_ = new_n2376_ | new_n2351_;
  assign new_n3266_ = new_n5067_ | new_n2071_;
  assign new_n3267_ = new_n3266_ | new_n5069_;
  assign new_n3268_ = new_n1912_ & new_n1896_;
  assign new_n3269_ = new_n5067_ | new_n5069_;
  assign new_n3270_ = new_n3269_ | new_n3268_;
  assign new_n3271_ = new_n2559_ | new_n5073_;
  assign new_n3272_ = new_n5075_ | new_n5078_;
  assign new_n3273_ = new_n3272_ & new_n3271_;
  assign new_n3274_ = new_n5080_ | new_n5073_;
  assign new_n3275_ = new_n5081_ | new_n5078_;
  assign new_n3276_ = new_n3275_ & new_n3274_;
  assign new_n3277_ = new_n2602_ & new_n5066_;
  assign new_n3278_ = new_n2558_ & new_n5064_;
  assign new_n3279_ = new_n3278_ | new_n3277_;
  assign new_n3280_ = new_n2567_ | new_n5072_;
  assign new_n3281_ = new_n2603_ | new_n5077_;
  assign new_n3282_ = new_n3281_ & new_n3280_;
  assign new_n3283_ = new_n2574_ | new_n2482_;
  assign new_n3284_ = new_n5082_ & new_n2483_;
  assign new_n3285_ = new_n5082_ & new_n2575_;
  assign new_n3286_ = new_n3285_ | new_n3284_;
  assign new_n3287_ = new_n5083_ | new_n2474_;
  assign new_n3288_ = new_n5084_ & new_n2475_;
  assign new_n3289_ = new_n5084_ & new_n2570_;
  assign new_n3290_ = new_n3289_ | new_n3288_;
  assign new_n3291_ = new_n3290_ | new_n3286_;
  assign new_n3292_ = new_n2943_ | new_n2717_;
  assign new_n3293_ = new_n2936_ | new_n2722_;
  assign new_n3294_ = new_n3293_ & new_n3292_;
  assign new_n3295_ = new_n3294_ & new_n1956_;
  assign new_n3296_ = new_n2922_ & new_n2701_;
  assign new_n3297_ = new_n2923_ | new_n2700_;
  assign new_n3298_ = new_n2920_ & new_n2703_;
  assign new_n3299_ = new_n2921_ | new_n2702_;
  assign new_n3300_ = new_n3299_ & new_n3297_;
  assign new_n3301_ = new_n3298_ | new_n3296_;
  assign new_n3302_ = new_n2881_ & new_n2867_;
  assign new_n3303_ = new_n2880_ | new_n2866_;
  assign new_n3304_ = new_n2871_ & new_n2865_;
  assign new_n3305_ = new_n2870_ | new_n2864_;
  assign new_n3306_ = new_n3304_ & new_n3302_;
  assign new_n3307_ = new_n3305_ | new_n3303_;
  assign new_n3308_ = new_n3307_ | new_n3300_;
  assign new_n3309_ = new_n3306_ | new_n3301_;
  assign new_n3310_ = new_n3309_ & new_n3308_;
  assign new_n3311_ = new_n2931_ & new_n2708_;
  assign new_n3312_ = new_n2930_ | new_n2709_;
  assign new_n3313_ = new_n2929_ & new_n2710_;
  assign new_n3314_ = new_n2928_ | new_n2711_;
  assign new_n3315_ = new_n3314_ & new_n3312_;
  assign new_n3316_ = new_n3313_ | new_n3311_;
  assign new_n3317_ = new_n2879_ & new_n2863_;
  assign new_n3318_ = new_n2878_ | new_n2862_;
  assign new_n3319_ = new_n2869_ & new_n2861_;
  assign new_n3320_ = new_n2868_ | new_n2860_;
  assign new_n3321_ = new_n3319_ & new_n3317_;
  assign new_n3322_ = new_n3320_ | new_n3318_;
  assign new_n3323_ = new_n3322_ | new_n3315_;
  assign new_n3324_ = new_n3321_ | new_n3316_;
  assign new_n3325_ = new_n3324_ & new_n3323_;
  assign new_n3326_ = new_n2906_ & new_n2845_;
  assign new_n3327_ = new_n2907_ & new_n2844_;
  assign new_n3328_ = new_n3327_ | new_n3326_;
  assign new_n3329_ = new_n2904_ & new_n2851_;
  assign new_n3330_ = new_n2905_ & new_n2850_;
  assign new_n3331_ = new_n3330_ | new_n3329_;
  assign new_n3332_ = new_n2892_ & new_n2843_;
  assign new_n3333_ = new_n2893_ & new_n2842_;
  assign new_n3334_ = new_n3333_ | new_n3332_;
  assign new_n3335_ = new_n2902_ & new_n2841_;
  assign new_n3336_ = new_n2903_ & new_n2840_;
  assign new_n3337_ = new_n3336_ | new_n3335_;
  assign new_n3338_ = new_n2900_ & new_n2829_;
  assign new_n3339_ = new_n2901_ & new_n2828_;
  assign new_n3340_ = new_n3339_ | new_n3338_;
  assign new_n3341_ = new_n3331_ | new_n3328_;
  assign new_n3342_ = new_n3341_ | new_n3334_;
  assign new_n3343_ = new_n3342_ | new_n3337_;
  assign new_n3344_ = new_n3343_ | new_n3340_;
  assign new_n3345_ = new_n2898_ & new_n2827_;
  assign new_n3346_ = new_n2899_ & new_n2826_;
  assign new_n3347_ = new_n3346_ | new_n3345_;
  assign new_n3348_ = new_n2890_ & new_n2839_;
  assign new_n3349_ = new_n2891_ & new_n2838_;
  assign new_n3350_ = new_n3349_ | new_n3348_;
  assign new_n3351_ = new_n2896_ & new_n2825_;
  assign new_n3352_ = new_n2897_ & new_n2824_;
  assign new_n3353_ = new_n3352_ | new_n3351_;
  assign new_n3354_ = new_n2888_ & new_n2823_;
  assign new_n3355_ = new_n2889_ & new_n2822_;
  assign new_n3356_ = new_n3355_ | new_n3354_;
  assign new_n3357_ = new_n2894_ & new_n2853_;
  assign new_n3358_ = new_n2895_ & new_n2852_;
  assign new_n3359_ = new_n3358_ | new_n3357_;
  assign new_n3360_ = new_n3350_ | new_n3347_;
  assign new_n3361_ = new_n3360_ | new_n3353_;
  assign new_n3362_ = new_n3361_ | new_n3356_;
  assign new_n3363_ = new_n3362_ | new_n3359_;
  assign new_n3364_ = new_n3363_ | new_n3344_;
  assign new_n3365_ = new_n2657_ | new_n2033_;
  assign new_n3366_ = new_n2584_ | new_n5083_;
  assign new_n3367_ = new_n3366_ & new_n3365_;
  assign new_n3368_ = new_n2918_ & new_n2837_;
  assign new_n3369_ = new_n2919_ & new_n2836_;
  assign new_n3370_ = new_n3369_ | new_n3368_;
  assign new_n3371_ = new_n3370_ | new_n3367_;
  assign new_n3372_ = new_n2916_ & new_n2835_;
  assign new_n3373_ = new_n2917_ & new_n2834_;
  assign new_n3374_ = new_n3373_ | new_n3372_;
  assign new_n3375_ = new_n2910_ & new_n2849_;
  assign new_n3376_ = new_n2911_ & new_n2848_;
  assign new_n3377_ = new_n3376_ | new_n3375_;
  assign new_n3378_ = new_n2914_ & new_n2833_;
  assign new_n3379_ = new_n2915_ & new_n2832_;
  assign new_n3380_ = new_n3379_ | new_n3378_;
  assign new_n3381_ = new_n2908_ & new_n2831_;
  assign new_n3382_ = new_n2909_ & new_n2830_;
  assign new_n3383_ = new_n3382_ | new_n3381_;
  assign new_n3384_ = new_n2912_ & new_n2847_;
  assign new_n3385_ = new_n2913_ & new_n2846_;
  assign new_n3386_ = new_n3385_ | new_n3384_;
  assign new_n3387_ = new_n3377_ | new_n3374_;
  assign new_n3388_ = new_n3387_ | new_n3380_;
  assign new_n3389_ = new_n3388_ | new_n3383_;
  assign new_n3390_ = new_n3389_ | new_n3386_;
  assign new_n3391_ = new_n3390_ | new_n3371_;
  assign new_n3392_ = new_n5074_ | new_n5085_;
  assign new_n3393_ = new_n5079_ | new_n5085_;
  assign new_n3394_ = new_n3393_ & new_n3392_;
  assign new_n3395_ = new_n3391_ | new_n3364_;
  assign new_n3396_ = new_n3395_ | new_n3394_;
  assign new_n3397_ = new_n5086_ & new_n5087_;
  assign new_n3398_ = new_n5088_ | new_n5089_;
  assign new_n3399_ = new_n5088_ & new_n5089_;
  assign new_n3400_ = new_n5086_ | new_n5087_;
  assign new_n3401_ = new_n3400_ & new_n3398_;
  assign new_n3402_ = new_n3399_ | new_n3397_;
  assign new_n3403_ = new_n3402_ & new_n2569_;
  assign new_n3404_ = new_n3401_ & new_n5091_;
  assign new_n3405_ = new_n3404_ | new_n3403_;
  assign new_n3406_ = new_n3405_ & new_n5065_;
  assign new_n3407_ = new_n5091_ & new_n5063_;
  assign new_n3408_ = new_n3407_ | new_n3406_;
  assign new_n3409_ = new_n2944_ | new_n2718_;
  assign new_n3410_ = new_n2939_ | new_n2725_;
  assign new_n3411_ = new_n3410_ & new_n3409_;
  assign new_n3412_ = new_n3411_ & new_n5092_;
  assign new_n3413_ = new_n5090_ | new_n5074_;
  assign new_n3414_ = new_n2935_ & new_n2712_;
  assign new_n3415_ = new_n2934_ | new_n2713_;
  assign new_n3416_ = new_n2933_ & new_n2714_;
  assign new_n3417_ = new_n2932_ | new_n2715_;
  assign new_n3418_ = new_n3417_ & new_n3415_;
  assign new_n3419_ = new_n3416_ | new_n3414_;
  assign new_n3420_ = new_n2883_ & new_n2876_;
  assign new_n3421_ = new_n2882_ | new_n2877_;
  assign new_n3422_ = new_n2875_ & new_n2873_;
  assign new_n3423_ = new_n2874_ | new_n2872_;
  assign new_n3424_ = new_n3422_ & new_n3420_;
  assign new_n3425_ = new_n3423_ | new_n3421_;
  assign new_n3426_ = new_n3425_ | new_n3418_;
  assign new_n3427_ = new_n3424_ | new_n3419_;
  assign new_n3428_ = new_n3427_ & new_n3426_;
  assign new_n3429_ = new_n3428_ | new_n5079_;
  assign new_n3430_ = new_n3429_ & new_n3413_;
  assign new_n3431_ = new_n2947_ | new_n2721_;
  assign new_n3432_ = new_n2940_ | new_n2726_;
  assign new_n3433_ = new_n3432_ & new_n3431_;
  assign new_n3434_ = new_n3433_ & new_n5092_;
  assign new_n3435_ = new_n5093_ & new_n2707_;
  assign new_n3436_ = new_n5093_ & new_n2705_;
  assign new_n3437_ = new_n3436_ | new_n3435_;
  assign new_n3438_ = new_n5094_ | new_n5095_;
  assign new_n3439_ = new_n3438_ | new_n5096_;
  assign new_n3440_ = new_n5097_ | new_n5098_;
  assign new_n3441_ = new_n3440_ | new_n5099_;
  assign new_n3442_ = new_n3441_ | new_n3439_;
  assign new_n3443_ = new_n3442_ | new_n5070_;
  assign new_n3444_ = new_n5100_ & new_n2359_;
  assign new_n3445_ = new_n5102_ | new_n2358_;
  assign new_n3446_ = new_n3174_ | new_n3150_;
  assign new_n3447_ = new_n3446_ | new_n3158_;
  assign new_n3448_ = new_n3447_ | new_n3154_;
  assign new_n3449_ = new_n3176_ | new_n3152_;
  assign new_n3450_ = new_n3449_ | new_n3160_;
  assign new_n3451_ = new_n3450_ | new_n3156_;
  assign new_n3452_ = new_n3218_ | new_n3164_;
  assign new_n3453_ = new_n3452_ | new_n3168_;
  assign new_n3454_ = new_n3453_ | new_n3166_;
  assign new_n3455_ = new_n3190_ & new_n5104_;
  assign new_n3456_ = new_n3455_ & new_n5105_;
  assign new_n3457_ = new_n3178_ & new_n5106_;
  assign new_n3458_ = new_n3457_ & new_n5105_;
  assign new_n3459_ = new_n3182_ & new_n5104_;
  assign new_n3460_ = new_n3459_ & new_n5107_;
  assign new_n3461_ = new_n3186_ & new_n5106_;
  assign new_n3462_ = new_n3461_ & new_n5107_;
  assign new_n3463_ = new_n3458_ | new_n3456_;
  assign new_n3464_ = new_n3463_ | new_n3460_;
  assign new_n3465_ = new_n3464_ | new_n3462_;
  assign new_n3466_ = new_n3206_ & new_n5110_;
  assign new_n3467_ = new_n3466_ & new_n5117_;
  assign new_n3468_ = new_n3194_ & new_n5124_;
  assign new_n3469_ = new_n3468_ & new_n5117_;
  assign new_n3470_ = new_n3202_ & new_n5110_;
  assign new_n3471_ = new_n3470_ & new_n5131_;
  assign new_n3472_ = new_n3198_ & new_n5124_;
  assign new_n3473_ = new_n3472_ & new_n5131_;
  assign new_n3474_ = new_n3469_ | new_n3467_;
  assign new_n3475_ = new_n3474_ | new_n3471_;
  assign new_n3476_ = new_n3475_ | new_n3473_;
  assign new_n3477_ = new_n3208_ & new_n5111_;
  assign new_n3478_ = new_n3477_ & new_n5118_;
  assign new_n3479_ = new_n3196_ & new_n5125_;
  assign new_n3480_ = new_n3479_ & new_n5118_;
  assign new_n3481_ = new_n3204_ & new_n5111_;
  assign new_n3482_ = new_n3481_ & new_n5132_;
  assign new_n3483_ = new_n3200_ & new_n5125_;
  assign new_n3484_ = new_n3483_ & new_n5132_;
  assign new_n3485_ = new_n3480_ | new_n3478_;
  assign new_n3486_ = new_n3485_ | new_n3482_;
  assign new_n3487_ = new_n3486_ | new_n3484_;
  assign new_n3488_ = new_n5139_ & new_n3192_;
  assign new_n3489_ = new_n5147_ | new_n3193_;
  assign new_n3490_ = new_n3488_ & new_n5153_;
  assign new_n3491_ = new_n3489_ | new_n5161_;
  assign new_n3492_ = new_n3180_ & new_n5167_;
  assign new_n3493_ = new_n3181_ | new_n5175_;
  assign new_n3494_ = new_n3492_ & new_n5153_;
  assign new_n3495_ = new_n3493_ | new_n5161_;
  assign new_n3496_ = new_n5139_ & new_n3184_;
  assign new_n3497_ = new_n5147_ | new_n3185_;
  assign new_n3498_ = new_n3496_ & new_n5181_;
  assign new_n3499_ = new_n3497_ | new_n5189_;
  assign new_n3500_ = new_n3188_ & new_n5167_;
  assign new_n3501_ = new_n3189_ | new_n5175_;
  assign new_n3502_ = new_n3500_ & new_n5181_;
  assign new_n3503_ = new_n3501_ | new_n5189_;
  assign new_n3504_ = new_n3495_ & new_n3491_;
  assign new_n3505_ = new_n3494_ | new_n3490_;
  assign new_n3506_ = new_n3504_ & new_n3499_;
  assign new_n3507_ = new_n3505_ | new_n3498_;
  assign new_n3508_ = new_n3506_ & new_n3503_;
  assign new_n3509_ = new_n3507_ | new_n3502_;
  assign new_n3510_ = new_n5140_ & new_n3130_;
  assign new_n3511_ = new_n5148_ | new_n3131_;
  assign new_n3512_ = new_n3510_ & new_n5154_;
  assign new_n3513_ = new_n3511_ | new_n5162_;
  assign new_n3514_ = new_n3118_ & new_n5168_;
  assign new_n3515_ = new_n3119_ | new_n5176_;
  assign new_n3516_ = new_n3514_ & new_n5154_;
  assign new_n3517_ = new_n3515_ | new_n5162_;
  assign new_n3518_ = new_n5140_ & new_n3122_;
  assign new_n3519_ = new_n5148_ | new_n3123_;
  assign new_n3520_ = new_n3518_ & new_n5182_;
  assign new_n3521_ = new_n3519_ | new_n5190_;
  assign new_n3522_ = new_n3126_ & new_n5168_;
  assign new_n3523_ = new_n3127_ | new_n5176_;
  assign new_n3524_ = new_n3522_ & new_n5182_;
  assign new_n3525_ = new_n3523_ | new_n5190_;
  assign new_n3526_ = new_n3517_ & new_n3513_;
  assign new_n3527_ = new_n3516_ | new_n3512_;
  assign new_n3528_ = new_n3526_ & new_n3521_;
  assign new_n3529_ = new_n3527_ | new_n3520_;
  assign new_n3530_ = new_n3528_ & new_n3525_;
  assign new_n3531_ = new_n3529_ | new_n3524_;
  assign new_n3532_ = new_n5141_ & new_n3132_;
  assign new_n3533_ = new_n5149_ | new_n3133_;
  assign new_n3534_ = new_n3532_ & new_n5155_;
  assign new_n3535_ = new_n3533_ | new_n5163_;
  assign new_n3536_ = new_n3120_ & new_n5169_;
  assign new_n3537_ = new_n3121_ | new_n5177_;
  assign new_n3538_ = new_n3536_ & new_n5155_;
  assign new_n3539_ = new_n3537_ | new_n5163_;
  assign new_n3540_ = new_n5141_ & new_n3124_;
  assign new_n3541_ = new_n5149_ | new_n3125_;
  assign new_n3542_ = new_n3540_ & new_n5183_;
  assign new_n3543_ = new_n3541_ | new_n5191_;
  assign new_n3544_ = new_n3128_ & new_n5169_;
  assign new_n3545_ = new_n3129_ | new_n5177_;
  assign new_n3546_ = new_n3544_ & new_n5183_;
  assign new_n3547_ = new_n3545_ | new_n5191_;
  assign new_n3548_ = new_n3539_ & new_n3535_;
  assign new_n3549_ = new_n3538_ | new_n3534_;
  assign new_n3550_ = new_n3548_ & new_n3543_;
  assign new_n3551_ = new_n3549_ | new_n3542_;
  assign new_n3552_ = new_n3550_ & new_n3547_;
  assign new_n3553_ = new_n3551_ | new_n3546_;
  assign new_n3554_ = new_n5195_ & new_n5202_;
  assign new_n3555_ = new_n5206_ | new_n5214_;
  assign new_n3556_ = new_n5206_ & new_n5216_;
  assign new_n3557_ = new_n5195_ | new_n5218_;
  assign new_n3558_ = new_n3557_ & new_n3555_;
  assign new_n3559_ = new_n3556_ | new_n3554_;
  assign new_n3560_ = new_n5223_ & new_n5202_;
  assign new_n3561_ = new_n5233_ | new_n5214_;
  assign new_n3562_ = new_n5233_ & new_n5216_;
  assign new_n3563_ = new_n5223_ | new_n5218_;
  assign new_n3564_ = new_n3563_ & new_n3561_;
  assign new_n3565_ = new_n3562_ | new_n3560_;
  assign new_n3566_ = new_n2775_ & new_n2742_;
  assign new_n3567_ = new_n3048_ | new_n3017_;
  assign new_n3568_ = new_n2773_ & new_n2748_;
  assign new_n3569_ = new_n3568_ & new_n5241_;
  assign new_n3570_ = new_n3046_ | new_n3023_;
  assign new_n3571_ = new_n2771_ & new_n2746_;
  assign new_n3572_ = new_n5244_ & new_n5241_;
  assign new_n3573_ = new_n3572_ & new_n3571_;
  assign new_n3574_ = new_n3044_ | new_n3021_;
  assign new_n3575_ = new_n2803_ & new_n2792_;
  assign new_n3576_ = new_n5245_ & new_n5242_;
  assign new_n3577_ = new_n3576_ & new_n3575_;
  assign new_n3578_ = new_n3577_ & new_n5244_;
  assign new_n3579_ = new_n3569_ | new_n3566_;
  assign new_n3580_ = new_n3579_ | new_n3573_;
  assign new_n3581_ = new_n3580_ | new_n3578_;
  assign new_n3582_ = new_n2765_ & new_n2734_;
  assign new_n3583_ = new_n2764_ | new_n2735_;
  assign new_n3584_ = new_n3039_ & new_n3008_;
  assign new_n3585_ = new_n3038_ | new_n3009_;
  assign new_n3586_ = new_n2763_ & new_n2732_;
  assign new_n3587_ = new_n2762_ | new_n2733_;
  assign new_n3588_ = new_n3586_ & new_n5248_;
  assign new_n3589_ = new_n3587_ | new_n5252_;
  assign new_n3590_ = new_n3037_ & new_n3006_;
  assign new_n3591_ = new_n3036_ | new_n3007_;
  assign new_n3592_ = new_n2787_ & new_n2756_;
  assign new_n3593_ = new_n2786_ | new_n2757_;
  assign new_n3594_ = new_n5255_ & new_n5248_;
  assign new_n3595_ = new_n5258_ | new_n5252_;
  assign new_n3596_ = new_n3594_ & new_n3592_;
  assign new_n3597_ = new_n3595_ | new_n3593_;
  assign new_n3598_ = new_n3063_ & new_n3030_;
  assign new_n3599_ = new_n3062_ | new_n3031_;
  assign new_n3600_ = new_n2785_ & new_n2754_;
  assign new_n3601_ = new_n2784_ | new_n2755_;
  assign new_n3602_ = new_n5261_ & new_n5247_;
  assign new_n3603_ = new_n5263_ | new_n5251_;
  assign new_n3604_ = new_n3602_ & new_n3600_;
  assign new_n3605_ = new_n3603_ | new_n3601_;
  assign new_n3606_ = new_n3604_ & new_n5255_;
  assign new_n3607_ = new_n3605_ | new_n5258_;
  assign new_n3608_ = new_n3061_ & new_n3028_;
  assign new_n3609_ = new_n3060_ | new_n3029_;
  assign new_n3610_ = new_n5264_ & new_n2731_;
  assign new_n3611_ = new_n5265_ | new_n2730_;
  assign new_n3612_ = new_n5266_ & new_n5261_;
  assign new_n3613_ = new_n5267_ | new_n5263_;
  assign new_n3614_ = new_n3612_ & new_n5249_;
  assign new_n3615_ = new_n3613_ | new_n5253_;
  assign new_n3616_ = new_n3614_ & new_n3610_;
  assign new_n3617_ = new_n3615_ | new_n3611_;
  assign new_n3618_ = new_n3616_ & new_n5256_;
  assign new_n3619_ = new_n3617_ | new_n5259_;
  assign new_n3620_ = new_n3589_ & new_n3583_;
  assign new_n3621_ = new_n3588_ | new_n3582_;
  assign new_n3622_ = new_n3620_ & new_n3597_;
  assign new_n3623_ = new_n3621_ | new_n3596_;
  assign new_n3624_ = new_n3622_ & new_n3607_;
  assign new_n3625_ = new_n3623_ | new_n3606_;
  assign new_n3626_ = new_n3624_ & new_n3619_;
  assign new_n3627_ = new_n3625_ | new_n3618_;
  assign new_n3628_ = new_n3056_ & new_n3005_;
  assign new_n3629_ = new_n3057_ | new_n3004_;
  assign new_n3630_ = new_n3629_ & new_n5256_;
  assign new_n3631_ = new_n3628_ | new_n5259_;
  assign new_n3632_ = new_n3630_ & new_n5260_;
  assign new_n3633_ = new_n3631_ | new_n5262_;
  assign new_n3634_ = new_n3632_ & new_n5249_;
  assign new_n3635_ = new_n3633_ | new_n5253_;
  assign new_n3636_ = new_n3634_ & new_n5266_;
  assign new_n3637_ = new_n3635_ | new_n5267_;
  assign new_n3638_ = new_n5269_ & new_n2683_;
  assign new_n3639_ = new_n5271_ | new_n2682_;
  assign new_n3640_ = new_n5272_ & new_n2993_;
  assign new_n3641_ = new_n5273_ | new_n2992_;
  assign new_n3642_ = new_n5272_ & new_n3088_;
  assign new_n3643_ = new_n5273_ | new_n3089_;
  assign new_n3644_ = new_n3642_ & new_n3099_;
  assign new_n3645_ = new_n3643_ | new_n3098_;
  assign new_n3646_ = new_n3641_ & new_n3639_;
  assign new_n3647_ = new_n3640_ | new_n3638_;
  assign new_n3648_ = new_n3646_ & new_n3645_;
  assign new_n3649_ = new_n3647_ | new_n3644_;
  assign new_n3650_ = new_n3649_ & new_n3636_;
  assign new_n3651_ = new_n3648_ | new_n3637_;
  assign new_n3652_ = new_n3651_ & new_n3626_;
  assign new_n3653_ = new_n3650_ | new_n3627_;
  assign new_n3654_ = new_n3652_ & new_n5274_;
  assign new_n3655_ = new_n3102_ & new_n2960_;
  assign new_n3656_ = new_n3113_ & new_n2951_;
  assign new_n3657_ = new_n3656_ | new_n3655_;
  assign new_n3658_ = new_n3657_ & new_n5243_;
  assign new_n3659_ = new_n3658_ & new_n5245_;
  assign new_n3660_ = new_n3659_ & new_n5242_;
  assign new_n3661_ = new_n3660_ | new_n5274_;
  assign new_n3662_ = new_n3661_ & new_n3653_;
  assign new_n3663_ = new_n3662_ | new_n3654_;
  assign new_n3664_ = new_n2781_ & new_n2744_;
  assign new_n3665_ = new_n3054_ | new_n3019_;
  assign new_n3666_ = new_n2779_ & new_n2752_;
  assign new_n3667_ = new_n3666_ & new_n5276_;
  assign new_n3668_ = new_n3052_ | new_n3027_;
  assign new_n3669_ = new_n2777_ & new_n2750_;
  assign new_n3670_ = new_n5279_ & new_n5276_;
  assign new_n3671_ = new_n3670_ & new_n3669_;
  assign new_n3672_ = new_n3050_ | new_n3025_;
  assign new_n3673_ = new_n2805_ & new_n2794_;
  assign new_n3674_ = new_n5280_ & new_n5277_;
  assign new_n3675_ = new_n3674_ & new_n3673_;
  assign new_n3676_ = new_n3675_ & new_n5279_;
  assign new_n3677_ = new_n3667_ | new_n3664_;
  assign new_n3678_ = new_n3677_ | new_n3671_;
  assign new_n3679_ = new_n3678_ | new_n3676_;
  assign new_n3680_ = new_n2769_ & new_n2740_;
  assign new_n3681_ = new_n2768_ | new_n2741_;
  assign new_n3682_ = new_n3043_ & new_n3014_;
  assign new_n3683_ = new_n3042_ | new_n3015_;
  assign new_n3684_ = new_n2767_ & new_n2738_;
  assign new_n3685_ = new_n2766_ | new_n2739_;
  assign new_n3686_ = new_n3684_ & new_n5283_;
  assign new_n3687_ = new_n3685_ | new_n5287_;
  assign new_n3688_ = new_n3041_ & new_n3012_;
  assign new_n3689_ = new_n3040_ | new_n3013_;
  assign new_n3690_ = new_n2791_ & new_n2760_;
  assign new_n3691_ = new_n2790_ | new_n2761_;
  assign new_n3692_ = new_n5290_ & new_n5283_;
  assign new_n3693_ = new_n5293_ | new_n5287_;
  assign new_n3694_ = new_n3692_ & new_n3690_;
  assign new_n3695_ = new_n3693_ | new_n3691_;
  assign new_n3696_ = new_n3067_ & new_n3034_;
  assign new_n3697_ = new_n3066_ | new_n3035_;
  assign new_n3698_ = new_n2789_ & new_n2758_;
  assign new_n3699_ = new_n2788_ | new_n2759_;
  assign new_n3700_ = new_n5296_ & new_n5282_;
  assign new_n3701_ = new_n5298_ | new_n5286_;
  assign new_n3702_ = new_n3700_ & new_n3698_;
  assign new_n3703_ = new_n3701_ | new_n3699_;
  assign new_n3704_ = new_n3702_ & new_n5290_;
  assign new_n3705_ = new_n3703_ | new_n5293_;
  assign new_n3706_ = new_n3065_ & new_n3032_;
  assign new_n3707_ = new_n3064_ | new_n3033_;
  assign new_n3708_ = new_n5264_ & new_n2737_;
  assign new_n3709_ = new_n5265_ | new_n2736_;
  assign new_n3710_ = new_n5299_ & new_n5296_;
  assign new_n3711_ = new_n5300_ | new_n5298_;
  assign new_n3712_ = new_n3710_ & new_n5284_;
  assign new_n3713_ = new_n3711_ | new_n5288_;
  assign new_n3714_ = new_n3712_ & new_n3708_;
  assign new_n3715_ = new_n3713_ | new_n3709_;
  assign new_n3716_ = new_n3714_ & new_n5291_;
  assign new_n3717_ = new_n3715_ | new_n5294_;
  assign new_n3718_ = new_n3687_ & new_n3681_;
  assign new_n3719_ = new_n3686_ | new_n3680_;
  assign new_n3720_ = new_n3718_ & new_n3695_;
  assign new_n3721_ = new_n3719_ | new_n3694_;
  assign new_n3722_ = new_n3720_ & new_n3705_;
  assign new_n3723_ = new_n3721_ | new_n3704_;
  assign new_n3724_ = new_n3722_ & new_n3717_;
  assign new_n3725_ = new_n3723_ | new_n3716_;
  assign new_n3726_ = new_n3058_ & new_n3011_;
  assign new_n3727_ = new_n3059_ | new_n3010_;
  assign new_n3728_ = new_n3727_ & new_n5291_;
  assign new_n3729_ = new_n3726_ | new_n5294_;
  assign new_n3730_ = new_n3728_ & new_n5295_;
  assign new_n3731_ = new_n3729_ | new_n5297_;
  assign new_n3732_ = new_n3730_ & new_n5284_;
  assign new_n3733_ = new_n3731_ | new_n5288_;
  assign new_n3734_ = new_n3732_ & new_n5299_;
  assign new_n3735_ = new_n3733_ | new_n5300_;
  assign new_n3736_ = new_n5269_ & new_n2685_;
  assign new_n3737_ = new_n5271_ | new_n2684_;
  assign new_n3738_ = new_n5301_ & new_n2995_;
  assign new_n3739_ = new_n5302_ | new_n2994_;
  assign new_n3740_ = new_n5301_ & new_n3092_;
  assign new_n3741_ = new_n5302_ | new_n3093_;
  assign new_n3742_ = new_n3740_ & new_n3101_;
  assign new_n3743_ = new_n3741_ | new_n3100_;
  assign new_n3744_ = new_n3739_ & new_n3737_;
  assign new_n3745_ = new_n3738_ | new_n3736_;
  assign new_n3746_ = new_n3744_ & new_n3743_;
  assign new_n3747_ = new_n3745_ | new_n3742_;
  assign new_n3748_ = new_n3747_ & new_n3734_;
  assign new_n3749_ = new_n3746_ | new_n3735_;
  assign new_n3750_ = new_n3749_ & new_n3724_;
  assign new_n3751_ = new_n3748_ | new_n3725_;
  assign new_n3752_ = new_n3750_ & new_n5303_;
  assign new_n3753_ = new_n3104_ & new_n2962_;
  assign new_n3754_ = new_n3115_ & new_n2953_;
  assign new_n3755_ = new_n3754_ | new_n3753_;
  assign new_n3756_ = new_n3755_ & new_n5278_;
  assign new_n3757_ = new_n3756_ & new_n5280_;
  assign new_n3758_ = new_n3757_ & new_n5277_;
  assign new_n3759_ = new_n3758_ | new_n5303_;
  assign new_n3760_ = new_n3759_ & new_n3751_;
  assign new_n3761_ = new_n3760_ | new_n3752_;
  assign new_n3762_ = new_n2654_ & new_n2619_;
  assign new_n3763_ = new_n2655_ & new_n2618_;
  assign new_n3764_ = new_n3763_ | new_n3762_;
  assign new_n3765_ = new_n2622_ & new_n2621_;
  assign new_n3766_ = new_n2623_ & new_n2620_;
  assign new_n3767_ = new_n3766_ | new_n3765_;
  assign new_n3768_ = new_n5304_ & new_n5305_;
  assign new_n3769_ = new_n5306_ | new_n5307_;
  assign new_n3770_ = new_n5306_ & new_n5307_;
  assign new_n3771_ = new_n5304_ | new_n5305_;
  assign new_n3772_ = new_n3771_ & new_n3769_;
  assign new_n3773_ = new_n3770_ | new_n3768_;
  assign new_n3774_ = new_n5308_ & new_n5309_;
  assign new_n3775_ = new_n5310_ | new_n5311_;
  assign new_n3776_ = new_n5310_ & new_n5311_;
  assign new_n3777_ = new_n5308_ | new_n5309_;
  assign new_n3778_ = new_n3777_ & new_n3775_;
  assign new_n3779_ = new_n3776_ | new_n3774_;
  assign new_n3780_ = new_n5312_ & new_n5313_;
  assign new_n3781_ = new_n5314_ | new_n5315_;
  assign new_n3782_ = new_n5314_ & new_n5315_;
  assign new_n3783_ = new_n5312_ | new_n5313_;
  assign new_n3784_ = new_n3783_ & new_n3781_;
  assign new_n3785_ = new_n3782_ | new_n3780_;
  assign new_n3786_ = new_n5316_ & new_n5317_;
  assign new_n3787_ = new_n5318_ | new_n5319_;
  assign new_n3788_ = new_n5318_ & new_n5319_;
  assign new_n3789_ = new_n5316_ | new_n5317_;
  assign new_n3790_ = new_n3789_ & new_n3787_;
  assign new_n3791_ = new_n3788_ | new_n3786_;
  assign new_n3792_ = new_n3790_ & new_n3785_;
  assign new_n3793_ = new_n3791_ & new_n3784_;
  assign new_n3794_ = new_n3793_ | new_n3792_;
  assign new_n3795_ = new_n5321_ & new_n5323_;
  assign new_n3796_ = new_n5324_ | new_n5326_;
  assign new_n3797_ = new_n5324_ & new_n5326_;
  assign new_n3798_ = new_n5321_ | new_n5323_;
  assign new_n3799_ = new_n3798_ & new_n3796_;
  assign new_n3800_ = new_n3797_ | new_n3795_;
  assign new_n3801_ = new_n5328_ & new_n5329_;
  assign new_n3802_ = new_n5331_ | new_n5333_;
  assign new_n3803_ = new_n5331_ & new_n5333_;
  assign new_n3804_ = new_n5328_ | new_n5329_;
  assign new_n3805_ = new_n3804_ & new_n3802_;
  assign new_n3806_ = new_n3803_ | new_n3801_;
  assign new_n3807_ = new_n3806_ | new_n3799_;
  assign new_n3808_ = new_n3805_ | new_n3800_;
  assign new_n3809_ = new_n3808_ & new_n3807_;
  assign new_n3810_ = new_n3778_ & new_n5335_;
  assign new_n3811_ = new_n5337_ & new_n3772_;
  assign new_n3812_ = new_n3811_ | new_n3810_;
  assign new_n3813_ = new_n5338_ & new_n5339_;
  assign new_n3814_ = new_n5340_ | new_n5341_;
  assign new_n3815_ = new_n5340_ & new_n5341_;
  assign new_n3816_ = new_n5338_ | new_n5339_;
  assign new_n3817_ = new_n3816_ & new_n3814_;
  assign new_n3818_ = new_n3815_ | new_n3813_;
  assign new_n3819_ = new_n5342_ & new_n5343_;
  assign new_n3820_ = new_n5344_ | new_n5345_;
  assign new_n3821_ = new_n5344_ & new_n5345_;
  assign new_n3822_ = new_n5342_ | new_n5343_;
  assign new_n3823_ = new_n3822_ & new_n3820_;
  assign new_n3824_ = new_n3821_ | new_n3819_;
  assign new_n3825_ = new_n3069_ & new_n2820_;
  assign new_n3826_ = new_n3068_ | new_n2821_;
  assign new_n3827_ = new_n3071_ & new_n2818_;
  assign new_n3828_ = new_n3070_ | new_n2819_;
  assign new_n3829_ = new_n3828_ & new_n3826_;
  assign new_n3830_ = new_n3827_ | new_n3825_;
  assign new_n3831_ = new_n5346_ | new_n5347_;
  assign new_n3832_ = new_n3831_ | new_n5348_;
  assign new_n3833_ = new_n5346_ | new_n5349_;
  assign new_n3834_ = new_n3833_ | new_n5350_;
  assign new_n3835_ = new_n3834_ & new_n3832_;
  assign new_n3836_ = new_n5351_ | new_n5349_;
  assign new_n3837_ = new_n3836_ | new_n5348_;
  assign new_n3838_ = new_n5351_ | new_n5347_;
  assign new_n3839_ = new_n3838_ | new_n5350_;
  assign new_n3840_ = new_n3839_ & new_n3837_;
  assign new_n3841_ = new_n3840_ & new_n3835_;
  assign new_n3842_ = new_n5352_ & new_n5353_;
  assign new_n3843_ = new_n5354_ | new_n5355_;
  assign new_n3844_ = new_n5354_ & new_n5355_;
  assign new_n3845_ = new_n5352_ | new_n5353_;
  assign new_n3846_ = new_n3845_ & new_n3843_;
  assign new_n3847_ = new_n3844_ | new_n3842_;
  assign new_n3848_ = new_n5356_ & new_n5357_;
  assign new_n3849_ = new_n5358_ | new_n5359_;
  assign new_n3850_ = new_n5358_ & new_n5359_;
  assign new_n3851_ = new_n5356_ | new_n5357_;
  assign new_n3852_ = new_n3851_ & new_n3849_;
  assign new_n3853_ = new_n3850_ | new_n3848_;
  assign new_n3854_ = new_n3078_ & new_n2955_;
  assign new_n3855_ = new_n3079_ | new_n2954_;
  assign new_n3856_ = new_n3106_ & new_n2855_;
  assign new_n3857_ = new_n3107_ | new_n2854_;
  assign new_n3858_ = new_n3857_ & new_n3855_;
  assign new_n3859_ = new_n3856_ | new_n3854_;
  assign new_n3860_ = new_n5360_ & new_n5361_;
  assign new_n3861_ = new_n3860_ & new_n5362_;
  assign new_n3862_ = new_n5360_ & new_n5363_;
  assign new_n3863_ = new_n3862_ & new_n5364_;
  assign new_n3864_ = new_n3863_ | new_n3861_;
  assign new_n3865_ = new_n5365_ & new_n5363_;
  assign new_n3866_ = new_n3865_ & new_n5362_;
  assign new_n3867_ = new_n5365_ & new_n5361_;
  assign new_n3868_ = new_n3867_ & new_n5364_;
  assign new_n3869_ = new_n3868_ | new_n3866_;
  assign new_n3870_ = new_n3869_ | new_n3864_;
  assign new_n3871_ = new_n5366_ & new_n5367_;
  assign new_n3872_ = new_n5368_ | new_n5369_;
  assign new_n3873_ = new_n5368_ & new_n5369_;
  assign new_n3874_ = new_n5366_ | new_n5367_;
  assign new_n3875_ = new_n3874_ & new_n3872_;
  assign new_n3876_ = new_n3873_ | new_n3871_;
  assign new_n3877_ = new_n5370_ & new_n5371_;
  assign new_n3878_ = new_n5372_ | new_n5373_;
  assign new_n3879_ = new_n5372_ & new_n5373_;
  assign new_n3880_ = new_n5370_ | new_n5371_;
  assign new_n3881_ = new_n3880_ & new_n3878_;
  assign new_n3882_ = new_n3879_ | new_n3877_;
  assign new_n3883_ = new_n3083_ & new_n2949_;
  assign new_n3884_ = new_n3082_ | new_n2948_;
  assign new_n3885_ = new_n3096_ & new_n2858_;
  assign new_n3886_ = new_n3097_ | new_n2859_;
  assign new_n3887_ = new_n3886_ & new_n3884_;
  assign new_n3888_ = new_n3885_ | new_n3883_;
  assign new_n3889_ = new_n5374_ | new_n5375_;
  assign new_n3890_ = new_n3889_ | new_n5376_;
  assign new_n3891_ = new_n5374_ | new_n5377_;
  assign new_n3892_ = new_n3891_ | new_n5378_;
  assign new_n3893_ = new_n3892_ & new_n3890_;
  assign new_n3894_ = new_n5379_ | new_n5377_;
  assign new_n3895_ = new_n3894_ | new_n5376_;
  assign new_n3896_ = new_n5379_ | new_n5375_;
  assign new_n3897_ = new_n3896_ | new_n5378_;
  assign new_n3898_ = new_n3897_ & new_n3895_;
  assign new_n3899_ = new_n3898_ & new_n3893_;
  assign new_n3900_ = new_n5196_ & new_n5380_;
  assign new_n3901_ = new_n5207_ & new_n5381_;
  assign new_n3902_ = new_n3901_ | new_n3900_;
  assign new_n3903_ = new_n5196_ | new_n5383_;
  assign new_n3904_ = new_n3903_ | new_n5388_;
  assign new_n3905_ = new_n5198_ | new_n5401_;
  assign new_n3906_ = new_n3905_ | new_n5388_;
  assign new_n3907_ = new_n5224_ & new_n5380_;
  assign new_n3908_ = new_n5234_ & new_n5381_;
  assign new_n3909_ = new_n3908_ | new_n3907_;
  assign new_n3910_ = new_n5224_ | new_n5383_;
  assign new_n3911_ = new_n3910_ | new_n5389_;
  assign new_n3912_ = new_n5226_ | new_n5401_;
  assign new_n3913_ = new_n3912_ | new_n5389_;
  assign new_n3914_ = new_n5198_ | new_n5405_;
  assign new_n3915_ = new_n2817_ & new_n2810_;
  assign new_n3916_ = new_n2816_ | new_n2811_;
  assign new_n3917_ = new_n3915_ & new_n3163_;
  assign new_n3918_ = new_n3916_ | new_n3162_;
  assign new_n3919_ = new_n5409_ | new_n3914_;
  assign new_n3920_ = new_n5226_ | new_n5405_;
  assign new_n3921_ = new_n3920_ | new_n5409_;
  assign new_n3922_ = new_n5207_ & new_n5411_;
  assign new_n3923_ = new_n3922_ & new_n5414_;
  assign new_n3924_ = new_n5209_ & new_n5419_;
  assign new_n3925_ = new_n3924_ & new_n5414_;
  assign new_n3926_ = new_n5234_ & new_n5411_;
  assign new_n3927_ = new_n3926_ & new_n5415_;
  assign new_n3928_ = new_n5236_ & new_n5419_;
  assign new_n3929_ = new_n3928_ & new_n5415_;
  assign new_n3930_ = new_n5209_ | new_n5421_;
  assign new_n3931_ = new_n5197_ | new_n5424_;
  assign new_n3932_ = new_n3931_ & new_n3930_;
  assign new_n3933_ = new_n3932_ | new_n5391_;
  assign new_n3934_ = new_n5208_ | new_n5427_;
  assign new_n3935_ = new_n5200_ | new_n5430_;
  assign new_n3936_ = new_n3935_ & new_n3934_;
  assign new_n3937_ = new_n3936_ | new_n5391_;
  assign new_n3938_ = new_n5236_ | new_n5421_;
  assign new_n3939_ = new_n5225_ | new_n5424_;
  assign new_n3940_ = new_n3939_ & new_n3938_;
  assign new_n3941_ = new_n3940_ | new_n5392_;
  assign new_n3942_ = new_n5235_ | new_n5427_;
  assign new_n3943_ = new_n5228_ | new_n5430_;
  assign new_n3944_ = new_n3943_ & new_n3942_;
  assign new_n3945_ = new_n3944_ | new_n5392_;
  assign new_n3946_ = new_n5434_ | new_n5437_;
  assign new_n3947_ = new_n3946_ | new_n5395_;
  assign new_n3948_ = new_n5441_ | new_n5437_;
  assign new_n3949_ = new_n3948_ | new_n5395_;
  assign new_n3950_ = new_n5434_ | new_n5444_;
  assign new_n3951_ = new_n3950_ | new_n5396_;
  assign new_n3952_ = new_n5441_ | new_n5444_;
  assign new_n3953_ = new_n3952_ | new_n5396_;
  assign new_n3954_ = new_n5447_ & new_n5448_;
  assign new_n3955_ = new_n3954_ & new_n5417_;
  assign new_n3956_ = new_n5450_ & new_n5448_;
  assign new_n3957_ = new_n3956_ & new_n5417_;
  assign new_n3958_ = new_n5452_ | new_n5453_;
  assign new_n3959_ = new_n3958_ | new_n5410_;
  assign new_n3960_ = new_n5456_ | new_n5438_;
  assign new_n3961_ = new_n5456_ | new_n5461_;
  assign new_n3962_ = new_n3961_ & new_n3960_;
  assign new_n3963_ = new_n3962_ | new_n5398_;
  assign new_n3964_ = new_n5464_ | new_n5438_;
  assign new_n3965_ = new_n5464_ | new_n5461_;
  assign new_n3966_ = new_n3965_ & new_n3964_;
  assign new_n3967_ = new_n3966_ | new_n5398_;
  assign new_n3968_ = new_n5457_ | new_n5445_;
  assign new_n3969_ = new_n5457_ | new_n5468_;
  assign new_n3970_ = new_n3969_ & new_n3968_;
  assign new_n3971_ = new_n3970_ | new_n5399_;
  assign new_n3972_ = new_n5465_ | new_n5445_;
  assign new_n3973_ = new_n5465_ | new_n5468_;
  assign new_n3974_ = new_n3973_ & new_n3972_;
  assign new_n3975_ = new_n3974_ | new_n5399_;
  assign new_n3976_ = new_n5211_ & new_n5469_;
  assign new_n3977_ = new_n3976_ & new_n5418_;
  assign new_n3978_ = new_n5238_ & new_n5469_;
  assign new_n3979_ = new_n3978_ & new_n5418_;
  assign new_n3980_ = new_n5113_ & new_n2326_;
  assign new_n3981_ = new_n3980_ & new_n5120_;
  assign new_n3982_ = new_n5127_ & new_n2236_;
  assign new_n3983_ = new_n3982_ & new_n5120_;
  assign new_n3984_ = new_n5113_ & new_n2296_;
  assign new_n3985_ = new_n3984_ & new_n5134_;
  assign new_n3986_ = new_n5127_ & new_n2266_;
  assign new_n3987_ = new_n3986_ & new_n5134_;
  assign new_n3988_ = new_n3983_ | new_n3981_;
  assign new_n3989_ = new_n3988_ | new_n3985_;
  assign new_n3990_ = new_n3989_ | new_n3987_;
  assign new_n3991_ = new_n5143_ & new_n2178_;
  assign new_n3992_ = new_n3991_ & new_n5157_;
  assign new_n3993_ = new_n5171_ & new_n2084_;
  assign new_n3994_ = new_n3993_ & new_n5157_;
  assign new_n3995_ = new_n5143_ & new_n2116_;
  assign new_n3996_ = new_n3995_ & new_n5185_;
  assign new_n3997_ = new_n5171_ & new_n2146_;
  assign new_n3998_ = new_n3997_ & new_n5185_;
  assign new_n3999_ = new_n3994_ | new_n3992_;
  assign new_n4000_ = new_n3999_ | new_n3996_;
  assign new_n4001_ = new_n4000_ | new_n3998_;
  assign new_n4002_ = new_n5144_ & new_n2206_;
  assign new_n4003_ = new_n4002_ & new_n5158_;
  assign new_n4004_ = new_n5172_ & new_n2112_;
  assign new_n4005_ = new_n4004_ & new_n5158_;
  assign new_n4006_ = new_n5144_ & new_n2142_;
  assign new_n4007_ = new_n4006_ & new_n5186_;
  assign new_n4008_ = new_n5172_ & new_n2174_;
  assign new_n4009_ = new_n4008_ & new_n5186_;
  assign new_n4010_ = new_n4005_ | new_n4003_;
  assign new_n4011_ = new_n4010_ | new_n4007_;
  assign new_n4012_ = new_n4011_ | new_n4009_;
  assign new_n4013_ = new_n5471_ | new_n5453_;
  assign new_n4014_ = new_n4013_ | new_n5410_;
  assign new_n4015_ = new_n5476_ & new_n3236_;
  assign new_n4016_ = new_n4015_ & new_n5485_;
  assign new_n4017_ = new_n5493_ & new_n3224_;
  assign new_n4018_ = new_n4017_ & new_n5485_;
  assign new_n4019_ = new_n5476_ & new_n3232_;
  assign new_n4020_ = new_n4019_ & new_n5498_;
  assign new_n4021_ = new_n5493_ & new_n3228_;
  assign new_n4022_ = new_n4021_ & new_n5498_;
  assign new_n4023_ = new_n4018_ | new_n4016_;
  assign new_n4024_ = new_n4023_ | new_n4020_;
  assign new_n4025_ = new_n4024_ | new_n4022_;
  assign new_n4026_ = new_n5494_ | new_n3239_;
  assign new_n4027_ = new_n4026_ | new_n5499_;
  assign new_n4028_ = new_n5477_ | new_n3227_;
  assign new_n4029_ = new_n4028_ | new_n5499_;
  assign new_n4030_ = new_n5494_ | new_n3235_;
  assign new_n4031_ = new_n4030_ | new_n5486_;
  assign new_n4032_ = new_n5477_ | new_n3231_;
  assign new_n4033_ = new_n4032_ | new_n5486_;
  assign new_n4034_ = new_n4029_ & new_n4027_;
  assign new_n4035_ = new_n4034_ & new_n4031_;
  assign new_n4036_ = new_n4035_ & new_n4033_;
  assign new_n4037_ = new_n5501_ & new_n5502_;
  assign new_n4038_ = new_n5503_ | new_n5504_;
  assign new_n4039_ = new_n5503_ & new_n5504_;
  assign new_n4040_ = new_n5501_ | new_n5502_;
  assign new_n4041_ = new_n4040_ & new_n4038_;
  assign new_n4042_ = new_n4039_ | new_n4037_;
  assign new_n4043_ = new_n5505_ & new_n5506_;
  assign new_n4044_ = new_n5507_ | new_n5508_;
  assign new_n4045_ = new_n5507_ & new_n5508_;
  assign new_n4046_ = new_n5505_ | new_n5506_;
  assign new_n4047_ = new_n4046_ & new_n4044_;
  assign new_n4048_ = new_n4045_ | new_n4043_;
  assign new_n4049_ = new_n2616_ & new_n2593_;
  assign new_n4050_ = new_n2617_ & new_n2592_;
  assign new_n4051_ = new_n4050_ | new_n4049_;
  assign new_n4052_ = new_n5509_ | new_n5510_;
  assign new_n4053_ = new_n4052_ | new_n5512_;
  assign new_n4054_ = new_n5514_ & new_n5510_;
  assign new_n4055_ = new_n4054_ & new_n5512_;
  assign new_n4056_ = new_n5516_ & new_n5517_;
  assign new_n4057_ = new_n5518_ | new_n5520_;
  assign new_n4058_ = new_n5518_ & new_n5520_;
  assign new_n4059_ = new_n5516_ | new_n5517_;
  assign new_n4060_ = new_n4059_ & new_n4057_;
  assign new_n4061_ = new_n4058_ | new_n4056_;
  assign new_n4062_ = new_n5521_ & new_n5522_;
  assign new_n4063_ = new_n5523_ | new_n5524_;
  assign new_n4064_ = new_n5523_ & new_n5524_;
  assign new_n4065_ = new_n5521_ | new_n5522_;
  assign new_n4066_ = new_n4065_ & new_n4063_;
  assign new_n4067_ = new_n4064_ | new_n4062_;
  assign new_n4068_ = new_n5525_ & new_n2599_;
  assign new_n4069_ = new_n2601_ & new_n5526_;
  assign new_n4070_ = new_n4069_ | new_n4068_;
  assign new_n4071_ = new_n5527_ | new_n5528_;
  assign new_n4072_ = new_n4071_ | new_n5530_;
  assign new_n4073_ = new_n5532_ & new_n5528_;
  assign new_n4074_ = new_n4073_ & new_n5530_;
  assign new_n4075_ = new_n5509_ & new_n5533_;
  assign new_n4076_ = new_n4075_ & new_n5513_;
  assign new_n4077_ = new_n5527_ & new_n5534_;
  assign new_n4078_ = new_n4077_ & new_n5531_;
  assign new_n4079_ = new_n5535_ & new_n5536_;
  assign new_n4080_ = new_n5537_ | new_n5538_;
  assign new_n4081_ = new_n5537_ & new_n5538_;
  assign new_n4082_ = new_n5535_ | new_n5536_;
  assign new_n4083_ = new_n4082_ & new_n4080_;
  assign new_n4084_ = new_n4081_ | new_n4079_;
  assign new_n4085_ = new_n5268_ & new_n2688_;
  assign new_n4086_ = new_n5270_ & new_n2689_;
  assign new_n4087_ = new_n4086_ | new_n4085_;
  assign new_n4088_ = new_n5539_ | new_n5541_;
  assign new_n4089_ = new_n4088_ | new_n5544_;
  assign new_n4090_ = new_n5546_ & new_n5541_;
  assign new_n4091_ = new_n4090_ & new_n5544_;
  assign new_n4092_ = new_n5539_ & new_n5547_;
  assign new_n4093_ = new_n4092_ & new_n5545_;
  assign new_n4094_ = new_n5514_ | new_n5533_;
  assign new_n4095_ = new_n4094_ | new_n5513_;
  assign new_n4096_ = new_n5532_ | new_n5534_;
  assign new_n4097_ = new_n4096_ | new_n5531_;
  assign new_n4098_ = new_n5546_ | new_n5547_;
  assign new_n4099_ = new_n4098_ | new_n5545_;
  assign new_n4100_ = new_n5551_ & new_n1918_;
  assign new_n4101_ = new_n5102_ & new_n5559_;
  assign new_n4102_ = new_n4101_ | new_n4100_;
  assign new_n4103_ = new_n5551_ & new_n1924_;
  assign new_n4104_ = new_n5564_ & new_n5559_;
  assign new_n4105_ = new_n4104_ | new_n4103_;
  assign new_n4106_ = new_n5550_ & new_n1930_;
  assign new_n4107_ = new_n2604_ & new_n5558_;
  assign new_n4108_ = new_n4107_ | new_n4106_;
  assign new_n4109_ = new_n1976_ & new_n5552_;
  assign new_n4110_ = new_n5566_ & new_n5560_;
  assign new_n4111_ = new_n4110_ | new_n4109_;
  assign new_n4112_ = new_n1982_ & new_n5552_;
  assign new_n4113_ = new_n2648_ & new_n5560_;
  assign new_n4114_ = new_n4113_ | new_n4112_;
  assign new_n4115_ = new_n1988_ & new_n5554_;
  assign new_n4116_ = new_n5567_ & new_n5562_;
  assign new_n4117_ = new_n4116_ | new_n4115_;
  assign new_n4118_ = new_n1994_ & new_n5554_;
  assign new_n4119_ = new_n5568_ & new_n5562_;
  assign new_n4120_ = new_n4119_ | new_n4118_;
  assign new_n4121_ = new_n2000_ & new_n5555_;
  assign new_n4122_ = new_n2606_ & new_n5563_;
  assign new_n4123_ = new_n4122_ | new_n4121_;
  assign new_n4124_ = new_n2006_ & new_n5555_;
  assign new_n4125_ = new_n2642_ & new_n5563_;
  assign new_n4126_ = new_n4125_ | new_n4124_;
  assign new_n4127_ = new_n5572_ & new_n2012_;
  assign new_n4128_ = new_n2644_ & new_n5579_;
  assign new_n4129_ = new_n4128_ | new_n4127_;
  assign new_n4130_ = new_n5572_ & new_n2018_;
  assign new_n4131_ = new_n2608_ & new_n5579_;
  assign new_n4132_ = new_n4131_ | new_n4130_;
  assign new_n4133_ = new_n5571_ & new_n2024_;
  assign new_n4134_ = new_n5583_ & new_n5580_;
  assign new_n4135_ = new_n4134_ | new_n4133_;
  assign new_n4136_ = new_n2044_ & new_n5573_;
  assign new_n4137_ = new_n2646_ & new_n5580_;
  assign new_n4138_ = new_n4137_ | new_n4136_;
  assign new_n4139_ = new_n2050_ & new_n5573_;
  assign new_n4140_ = new_n2796_ & new_n5582_;
  assign new_n4141_ = new_n4140_ | new_n4139_;
  assign new_n4142_ = new_n2056_ & new_n5575_;
  assign new_n4143_ = new_n5327_ & new_n5582_;
  assign new_n4144_ = new_n4143_ | new_n4142_;
  assign new_n4145_ = new_n2062_ & new_n5575_;
  assign new_n4146_ = new_n5322_ & new_n5581_;
  assign new_n4147_ = new_n4146_ | new_n4145_;
  assign new_n4148_ = new_n5566_ | new_n5103_;
  assign new_n4149_ = new_n2799_ | new_n5100_;
  assign new_n4150_ = new_n4149_ & new_n4148_;
  assign new_n4151_ = new_n5584_ & new_n5585_;
  assign new_n4152_ = new_n5586_ | new_n2408_;
  assign new_n4153_ = new_n5587_ | new_n5589_;
  assign new_n4154_ = new_n4153_ | new_n2081_;
  assign new_n4155_ = new_n5200_ & new_n5590_;
  assign new_n4156_ = new_n5211_ | new_n5406_;
  assign new_n4157_ = new_n5212_ & new_n5591_;
  assign new_n4158_ = new_n5201_ | new_n5593_;
  assign new_n4159_ = new_n4158_ & new_n4156_;
  assign new_n4160_ = new_n4157_ | new_n4155_;
  assign new_n4161_ = new_n5595_ | new_n5598_;
  assign new_n4162_ = new_n5228_ & new_n5590_;
  assign new_n4163_ = new_n5238_ | new_n5406_;
  assign new_n4164_ = new_n5239_ & new_n5591_;
  assign new_n4165_ = new_n5229_ | new_n5593_;
  assign new_n4166_ = new_n4165_ & new_n4163_;
  assign new_n4167_ = new_n4164_ | new_n4162_;
  assign new_n4168_ = new_n5602_ | new_n5598_;
  assign new_n4169_ = new_n5604_ | new_n5606_;
  assign new_n4170_ = new_n5609_ & new_n5611_;
  assign new_n4171_ = new_n5613_ & new_n5615_;
  assign new_n4172_ = new_n5617_ | new_n5606_;
  assign new_n4173_ = new_n5619_ & new_n5621_;
  assign new_n4174_ = new_n5623_ & new_n5625_;
  assign new_n4175_ = new_n5628_ & new_n5632_;
  assign new_n4176_ = new_n5628_ & new_n5634_;
  assign new_n4177_ = new_n5637_ | new_n5641_;
  assign new_n4178_ = new_n5644_ | new_n5648_;
  assign new_n4179_ = new_n5637_ | new_n5650_;
  assign new_n4180_ = new_n5644_ | new_n5652_;
  assign new_n4181_ = new_n5654_ & new_n5656_;
  assign new_n4182_ = new_n5658_ & new_n5660_;
  assign new_n4183_ = new_n5662_ & new_n5664_;
  assign new_n4184_ = new_n5666_ & new_n5668_;
  assign new_n4185_ = new_n5609_ | new_n5611_;
  assign new_n4186_ = new_n5613_ | new_n5615_;
  assign new_n4187_ = new_n5619_ | new_n5621_;
  assign new_n4188_ = new_n5623_ | new_n5625_;
  assign new_n4189_ = new_n5638_ & new_n5641_;
  assign new_n4190_ = new_n5645_ & new_n5648_;
  assign new_n4191_ = new_n5629_ | new_n5632_;
  assign new_n4192_ = new_n5638_ & new_n5650_;
  assign new_n4193_ = new_n5645_ & new_n5652_;
  assign new_n4194_ = new_n5629_ | new_n5634_;
  assign new_n4195_ = new_n5604_ & new_n5607_;
  assign new_n4196_ = new_n5617_ & new_n5607_;
  assign new_n4197_ = new_n5654_ | new_n5656_;
  assign new_n4198_ = new_n5658_ | new_n5660_;
  assign new_n4199_ = new_n5662_ | new_n5664_;
  assign new_n4200_ = new_n5666_ | new_n5668_;
  assign new_n4201_ = new_n5670_ & new_n2318_;
  assign new_n4202_ = new_n4201_ & new_n5673_;
  assign new_n4203_ = new_n5676_ & new_n2228_;
  assign new_n4204_ = new_n4203_ & new_n5673_;
  assign new_n4205_ = new_n5670_ & new_n2288_;
  assign new_n4206_ = new_n4205_ & new_n5679_;
  assign new_n4207_ = new_n5676_ & new_n2258_;
  assign new_n4208_ = new_n4207_ & new_n5679_;
  assign new_n4209_ = new_n4204_ | new_n4202_;
  assign new_n4210_ = new_n4209_ | new_n4206_;
  assign new_n4211_ = new_n4210_ | new_n4208_;
  assign new_n4212_ = new_n5671_ & new_n2322_;
  assign new_n4213_ = new_n4212_ & new_n5674_;
  assign new_n4214_ = new_n5677_ & new_n2232_;
  assign new_n4215_ = new_n4214_ & new_n5674_;
  assign new_n4216_ = new_n5671_ & new_n2292_;
  assign new_n4217_ = new_n4216_ & new_n5680_;
  assign new_n4218_ = new_n5677_ & new_n2262_;
  assign new_n4219_ = new_n4218_ & new_n5680_;
  assign new_n4220_ = new_n4215_ | new_n4213_;
  assign new_n4221_ = new_n4220_ | new_n4217_;
  assign new_n4222_ = new_n4221_ | new_n4219_;
  assign new_n4223_ = new_n5681_ | new_n5682_;
  assign new_n4224_ = new_n5681_ | new_n5683_;
  assign new_n4225_ = new_n5682_ | new_n5684_;
  assign new_n4226_ = new_n5684_ | new_n5683_;
  assign new_n4227_ = new_n4224_ & new_n4223_;
  assign new_n4228_ = new_n4227_ & new_n4225_;
  assign new_n4229_ = new_n4228_ & new_n4226_;
  assign new_n4230_ = new_n5114_ & new_n2334_;
  assign new_n4231_ = new_n4230_ & new_n5121_;
  assign new_n4232_ = new_n5128_ & new_n2244_;
  assign new_n4233_ = new_n4232_ & new_n5121_;
  assign new_n4234_ = new_n5114_ & new_n2304_;
  assign new_n4235_ = new_n4234_ & new_n5135_;
  assign new_n4236_ = new_n5128_ & new_n2274_;
  assign new_n4237_ = new_n4236_ & new_n5135_;
  assign new_n4238_ = new_n4233_ | new_n4231_;
  assign new_n4239_ = new_n4238_ | new_n4235_;
  assign new_n4240_ = new_n4239_ | new_n4237_;
  assign new_n4241_ = new_n4160_ & new_n5599_;
  assign new_n4242_ = new_n5595_ & new_n5685_;
  assign new_n4243_ = new_n4242_ | new_n4241_;
  assign new_n4244_ = new_n5686_ | new_n5689_;
  assign new_n4245_ = new_n3559_ | new_n5692_;
  assign new_n4246_ = new_n4245_ & new_n4244_;
  assign new_n4247_ = new_n4167_ & new_n5599_;
  assign new_n4248_ = new_n5602_ & new_n5685_;
  assign new_n4249_ = new_n4248_ | new_n4247_;
  assign new_n4250_ = new_n5693_ | new_n5689_;
  assign new_n4251_ = new_n3565_ | new_n5692_;
  assign new_n4252_ = new_n4251_ & new_n4250_;
  assign new_n4253_ = new_n5212_ | new_n5695_;
  assign new_n4254_ = new_n5201_ | new_n5698_;
  assign new_n4255_ = new_n4254_ & new_n4253_;
  assign new_n4256_ = new_n4255_ | new_n5702_;
  assign new_n4257_ = new_n5239_ | new_n5695_;
  assign new_n4258_ = new_n5229_ | new_n5698_;
  assign new_n4259_ = new_n4258_ & new_n4257_;
  assign new_n4260_ = new_n4259_ | new_n5702_;
  assign new_n4261_ = new_n5706_ & new_n2096_;
  assign new_n4262_ = new_n4261_ & new_n5714_;
  assign new_n4263_ = new_n5706_ & new_n2098_;
  assign new_n4264_ = new_n4263_ & new_n5714_;
  assign new_n4265_ = new_n5707_ & new_n2158_;
  assign new_n4266_ = new_n4265_ & new_n5724_;
  assign new_n4267_ = new_n5707_ & new_n2160_;
  assign new_n4268_ = new_n4267_ & new_n5724_;
  assign new_n4269_ = new_n5732_ & new_n2128_;
  assign new_n4270_ = new_n4269_ & new_n5725_;
  assign new_n4271_ = new_n5725_ & new_n5732_;
  assign new_n4272_ = new_n5495_ & new_n2238_;
  assign new_n4273_ = new_n4272_ & new_n5487_;
  assign new_n4274_ = new_n5495_ & new_n2268_;
  assign new_n4275_ = new_n4274_ & new_n5500_;
  assign new_n4276_ = new_n5478_ & new_n2298_;
  assign new_n4277_ = new_n4276_ & new_n5500_;
  assign new_n4278_ = new_n5733_ & new_n2190_;
  assign new_n4279_ = new_n4278_ & new_n5715_;
  assign new_n4280_ = new_n5733_ & new_n2192_;
  assign new_n4281_ = new_n4280_ & new_n5715_;
  assign new_n4282_ = new_n5735_ & new_n2194_;
  assign new_n4283_ = new_n4282_ & new_n5717_;
  assign new_n4284_ = new_n5709_ & new_n2100_;
  assign new_n4285_ = new_n4284_ & new_n5717_;
  assign new_n4286_ = new_n5735_ & new_n2130_;
  assign new_n4287_ = new_n4286_ & new_n5727_;
  assign new_n4288_ = new_n5709_ & new_n2162_;
  assign new_n4289_ = new_n4288_ & new_n5727_;
  assign new_n4290_ = new_n4285_ | new_n4283_;
  assign new_n4291_ = new_n4290_ | new_n4287_;
  assign new_n4292_ = new_n4291_ | new_n4289_;
  assign new_n4293_ = new_n5736_ & new_n2196_;
  assign new_n4294_ = new_n4293_ & new_n5718_;
  assign new_n4295_ = new_n5710_ & new_n2102_;
  assign new_n4296_ = new_n4295_ & new_n5718_;
  assign new_n4297_ = new_n5736_ & new_n2132_;
  assign new_n4298_ = new_n4297_ & new_n5728_;
  assign new_n4299_ = new_n5710_ & new_n2164_;
  assign new_n4300_ = new_n4299_ & new_n5728_;
  assign new_n4301_ = new_n4296_ | new_n4294_;
  assign new_n4302_ = new_n4301_ | new_n4298_;
  assign new_n4303_ = new_n4302_ | new_n4300_;
  assign new_n4304_ = new_n5478_ & new_n2328_;
  assign new_n4305_ = new_n4304_ & new_n5487_;
  assign G2531 = new_n5049_;
  assign G2532 = new_n5050_;
  assign G2533 = G2532;
  assign G2534 = new_n5740_;
  assign G2535 = G2534;
  assign G2536 = new_n5742_;
  assign G2537 = G2536;
  assign G2538 = new_n5741_;
  assign G2539 = new_n5060_;
  assign G2540 = new_n5057_;
  assign G2541 = new_n5058_;
  assign G2542 = new_n5059_;
  assign G2543 = new_n5056_;
  assign G2544 = new_n5053_;
  assign G2545 = new_n5054_;
  assign G2546 = new_n5055_;
  assign G2547 = new_n3246_;
  assign G2548 = new_n3248_;
  assign G2549 = new_n2342_;
  assign G2550 = new_n3249_;
  assign G2551 = new_n5051_;
  assign G2552 = new_n3251_;
  assign G2553 = new_n3252_;
  assign G2554 = new_n5743_;
  assign G2555 = G2554;
  assign G2556 = new_n5070_;
  assign G2557 = new_n2541_;
  assign G2558 = new_n2573_;
  assign G2559 = new_n2543_;
  assign G2560 = new_n2545_;
  assign G2561 = new_n5081_;
  assign G2562 = new_n2557_;
  assign G2563 = new_n3264_;
  assign G2564 = new_n3267_;
  assign G2565 = new_n3270_;
  assign G2566 = new_n5080_;
  assign G2567 = new_n5075_;
  assign G2568 = new_n2550_;
  assign G2569 = new_n2548_;
  assign G2570 = new_n2554_;
  assign G2571 = new_n2552_;
  assign G2572 = new_n2560_;
  assign G2573 = new_n5744_;
  assign G2574 = G2573;
  assign G2575 = new_n5745_;
  assign G2576 = G2575;
  assign G2577 = new_n3279_;
  assign G2578 = new_n5746_;
  assign G2579 = G2578;
  assign G2580 = new_n3291_;
  assign G2581 = ~new_n5098_;
  assign G2582 = new_n5096_;
  assign G2583 = new_n5097_;
  assign G2584 = new_n5747_;
  assign G2585 = G2584;
  assign G2586 = new_n3408_;
  assign G2587 = ~new_n5095_;
  assign G2588 = new_n5748_;
  assign G2589 = G2588;
  assign G2590 = ~new_n5094_;
  assign G2591 = new_n2706_;
  assign G2592 = new_n5099_;
  assign G2593 = new_n5749_;
  assign G2594 = G2593;
  assign n1416_li = new_n1576_;
  assign n1419_li = new_n1890_;
  assign n1422_li = new_n1892_;
  assign n1425_li = new_n1894_;
  assign n1428_li = new_n1578_;
  assign n1431_li = new_n1898_;
  assign n1434_li = new_n1900_;
  assign n1437_li = new_n1902_;
  assign n1440_li = new_n1580_;
  assign n1443_li = new_n1906_;
  assign n1446_li = new_n1908_;
  assign n1449_li = new_n1910_;
  assign n1452_li = new_n1582_;
  assign n1455_li = new_n1914_;
  assign n1458_li = new_n1916_;
  assign n1464_li = new_n1584_;
  assign n1467_li = new_n1920_;
  assign n1470_li = new_n1922_;
  assign n1476_li = new_n1586_;
  assign n1479_li = new_n1926_;
  assign n1482_li = new_n1928_;
  assign n1488_li = new_n1588_;
  assign n1491_li = new_n1932_;
  assign n1494_li = new_n1934_;
  assign n1497_li = new_n1936_;
  assign n1500_li = new_n1590_;
  assign n1512_li = new_n1592_;
  assign n1515_li = new_n1942_;
  assign n1518_li = new_n1944_;
  assign n1521_li = new_n1946_;
  assign n1524_li = new_n1594_;
  assign n1527_li = new_n1950_;
  assign n1530_li = new_n1952_;
  assign n1533_li = new_n1954_;
  assign n1536_li = new_n1596_;
  assign n1539_li = new_n1958_;
  assign n1542_li = new_n1960_;
  assign n1545_li = new_n1962_;
  assign n1548_li = new_n1598_;
  assign n1551_li = new_n1966_;
  assign n1554_li = new_n1968_;
  assign n1560_li = new_n1600_;
  assign n1563_li = new_n1972_;
  assign n1566_li = new_n1974_;
  assign n1572_li = new_n1602_;
  assign n1575_li = new_n1978_;
  assign n1578_li = new_n1980_;
  assign n1584_li = new_n1604_;
  assign n1587_li = new_n1984_;
  assign n1590_li = new_n1986_;
  assign n1596_li = new_n1606_;
  assign n1599_li = new_n1990_;
  assign n1602_li = new_n1992_;
  assign n1608_li = new_n1608_;
  assign n1611_li = new_n1996_;
  assign n1614_li = new_n1998_;
  assign n1620_li = new_n1610_;
  assign n1623_li = new_n2002_;
  assign n1626_li = new_n2004_;
  assign n1632_li = new_n1612_;
  assign n1635_li = new_n2008_;
  assign n1638_li = new_n2010_;
  assign n1644_li = new_n1614_;
  assign n1647_li = new_n2014_;
  assign n1650_li = new_n2016_;
  assign n1656_li = new_n1616_;
  assign n1659_li = new_n2020_;
  assign n1662_li = new_n2022_;
  assign n1668_li = new_n1618_;
  assign n1671_li = new_n2026_;
  assign n1674_li = new_n2028_;
  assign n1677_li = new_n2030_;
  assign n1680_li = new_n1620_;
  assign n1683_li = new_n2034_;
  assign n1686_li = new_n2036_;
  assign n1692_li = new_n1622_;
  assign n1695_li = new_n2040_;
  assign n1698_li = new_n2042_;
  assign n1704_li = new_n1624_;
  assign n1707_li = new_n2046_;
  assign n1710_li = new_n2048_;
  assign n1716_li = new_n1626_;
  assign n1719_li = new_n2052_;
  assign n1722_li = new_n2054_;
  assign n1728_li = new_n1628_;
  assign n1731_li = new_n2058_;
  assign n1734_li = new_n2060_;
  assign n1740_li = new_n1630_;
  assign n1743_li = new_n2064_;
  assign n1746_li = new_n2066_;
  assign n1749_li = new_n2068_;
  assign n1752_li = new_n1632_;
  assign n1755_li = new_n2072_;
  assign n1758_li = new_n2074_;
  assign n1761_li = new_n2076_;
  assign n1764_li = new_n1634_;
  assign n1776_li = new_n1636_;
  assign n1779_li = new_n2082_;
  assign n1788_li = new_n1638_;
  assign n1791_li = new_n2086_;
  assign n1794_li = new_n2088_;
  assign n1797_li = new_n2090_;
  assign n1800_li = new_n1640_;
  assign n1812_li = new_n1642_;
  assign n1824_li = new_n1644_;
  assign n1836_li = new_n1646_;
  assign n1848_li = new_n1648_;
  assign n1860_li = new_n1650_;
  assign n1872_li = new_n1652_;
  assign n1884_li = new_n1654_;
  assign n1896_li = new_n1656_;
  assign n1899_li = new_n2110_;
  assign n1908_li = new_n1658_;
  assign n1911_li = new_n2114_;
  assign n1920_li = new_n1660_;
  assign n1923_li = new_n2118_;
  assign n1926_li = new_n2120_;
  assign n1929_li = new_n2122_;
  assign n1932_li = new_n1662_;
  assign n1944_li = new_n1664_;
  assign n1956_li = new_n1666_;
  assign n1968_li = new_n1668_;
  assign n1980_li = new_n1670_;
  assign n1992_li = new_n1672_;
  assign n2004_li = new_n1674_;
  assign n2016_li = new_n1676_;
  assign n2019_li = new_n2140_;
  assign n2028_li = new_n1678_;
  assign n2031_li = new_n2144_;
  assign n2040_li = new_n1680_;
  assign n2043_li = new_n2148_;
  assign n2046_li = new_n2150_;
  assign n2049_li = new_n2152_;
  assign n2052_li = new_n1682_;
  assign n2064_li = new_n1684_;
  assign n2076_li = new_n1686_;
  assign n2088_li = new_n1688_;
  assign n2100_li = new_n1690_;
  assign n2112_li = new_n1692_;
  assign n2124_li = new_n1694_;
  assign n2136_li = new_n1696_;
  assign n2148_li = new_n1698_;
  assign n2151_li = new_n2172_;
  assign n2160_li = new_n1700_;
  assign n2163_li = new_n2176_;
  assign n2172_li = new_n1702_;
  assign n2175_li = new_n2180_;
  assign n2178_li = new_n2182_;
  assign n2181_li = new_n2184_;
  assign n2184_li = new_n1704_;
  assign n2196_li = new_n1706_;
  assign n2208_li = new_n1708_;
  assign n2220_li = new_n1710_;
  assign n2232_li = new_n1712_;
  assign n2244_li = new_n1714_;
  assign n2256_li = new_n1716_;
  assign n2268_li = new_n1718_;
  assign n2280_li = new_n1720_;
  assign n2283_li = new_n2204_;
  assign n2292_li = new_n1722_;
  assign n2295_li = new_n2208_;
  assign n2298_li = new_n2210_;
  assign n2301_li = new_n2212_;
  assign n2304_li = new_n1724_;
  assign n2316_li = new_n1726_;
  assign n2319_li = new_n2218_;
  assign n2322_li = new_n2220_;
  assign n2325_li = new_n2222_;
  assign n2328_li = new_n1728_;
  assign n2331_li = new_n2226_;
  assign n2340_li = new_n1730_;
  assign n2343_li = new_n2230_;
  assign n2376_li = new_n1736_;
  assign n2379_li = new_n2234_;
  assign n2388_li = new_n1738_;
  assign n2400_li = new_n1740_;
  assign n2412_li = new_n1742_;
  assign n2415_li = new_n2242_;
  assign n2424_li = new_n1744_;
  assign n2436_li = new_n1746_;
  assign n2439_li = new_n2248_;
  assign n2442_li = new_n2250_;
  assign n2445_li = new_n2252_;
  assign n2448_li = new_n1748_;
  assign n2451_li = new_n2256_;
  assign n2460_li = new_n1750_;
  assign n2463_li = new_n2260_;
  assign n2496_li = new_n1756_;
  assign n2499_li = new_n2264_;
  assign n2508_li = new_n1758_;
  assign n2520_li = new_n1760_;
  assign n2532_li = new_n1762_;
  assign n2535_li = new_n2272_;
  assign n2544_li = new_n1764_;
  assign n2556_li = new_n1766_;
  assign n2559_li = new_n2278_;
  assign n2562_li = new_n2280_;
  assign n2565_li = new_n2282_;
  assign n2568_li = new_n1768_;
  assign n2571_li = new_n2286_;
  assign n2580_li = new_n1770_;
  assign n2583_li = new_n2290_;
  assign n2616_li = new_n1776_;
  assign n2619_li = new_n2294_;
  assign n2628_li = new_n1778_;
  assign n2640_li = new_n1780_;
  assign n2652_li = new_n1782_;
  assign n2655_li = new_n2302_;
  assign n2664_li = new_n1784_;
  assign n2676_li = new_n1786_;
  assign n2679_li = new_n2308_;
  assign n2682_li = new_n2310_;
  assign n2685_li = new_n2312_;
  assign n2688_li = new_n1788_;
  assign n2691_li = new_n2316_;
  assign n2700_li = new_n1790_;
  assign n2703_li = new_n2320_;
  assign n2736_li = new_n1796_;
  assign n2739_li = new_n2324_;
  assign n2748_li = new_n1798_;
  assign n2760_li = new_n1800_;
  assign n2772_li = new_n1802_;
  assign n2775_li = new_n2332_;
  assign n2784_li = new_n1804_;
  assign n2787_li = new_n2336_;
  assign n2790_li = new_n2338_;
  assign n2793_li = new_n2340_;
  assign n2796_li = new_n1806_;
  assign n2799_li = new_n2344_;
  assign n2802_li = new_n2346_;
  assign n2805_li = new_n2348_;
  assign n2808_li = new_n1808_;
  assign n2820_li = new_n1810_;
  assign n2823_li = new_n2354_;
  assign n2826_li = new_n2356_;
  assign n2832_li = new_n1812_;
  assign n2835_li = new_n2360_;
  assign n2838_li = new_n2362_;
  assign n2841_li = new_n2364_;
  assign n2844_li = new_n1814_;
  assign n2856_li = new_n1816_;
  assign n2859_li = new_n2370_;
  assign n2862_li = new_n2372_;
  assign n2865_li = new_n2374_;
  assign n2868_li = new_n1818_;
  assign n2871_li = new_n2378_;
  assign n2874_li = new_n2380_;
  assign n2877_li = new_n2382_;
  assign n2880_li = new_n1820_;
  assign n2883_li = new_n2386_;
  assign n2886_li = new_n2388_;
  assign n2889_li = new_n2390_;
  assign n2892_li = new_n1822_;
  assign n2895_li = new_n2394_;
  assign n2898_li = new_n2396_;
  assign n2901_li = new_n2398_;
  assign n2904_li = new_n1824_;
  assign n2907_li = new_n2402_;
  assign n2916_li = new_n1826_;
  assign n2928_li = new_n1828_;
  assign n2940_li = new_n1830_;
  assign n2952_li = new_n1832_;
  assign n2955_li = new_n2412_;
  assign n2964_li = new_n1834_;
  assign n2976_li = new_n1836_;
  assign n2988_li = new_n1838_;
  assign n2991_li = new_n2420_;
  assign n3000_li = new_n1840_;
  assign n3003_li = new_n2424_;
  assign n3012_li = new_n1842_;
  assign n3015_li = new_n2428_;
  assign n3024_li = new_n1844_;
  assign n3027_li = new_n2432_;
  assign n3036_li = new_n1846_;
  assign n3039_li = new_n2436_;
  assign n3048_li = new_n1848_;
  assign n3051_li = new_n2440_;
  assign n3054_li = new_n2442_;
  assign n3057_li = new_n2444_;
  assign n3060_li = new_n1850_;
  assign n3072_li = new_n1852_;
  assign n3081_li = new_n5519_;
  assign n3084_li = new_n1854_;
  assign n3087_li = new_n2454_;
  assign n3093_li = new_n5515_;
  assign n3096_li = new_n1856_;
  assign n3105_li = new_n5526_;
  assign n3108_li = new_n1858_;
  assign n3117_li = new_n5525_;
  assign n3120_li = new_n1860_;
  assign n3123_li = new_n2468_;
  assign n3126_li = new_n2470_;
  assign n3129_li = new_n5751_;
  assign n3132_li = new_n1862_;
  assign n3135_li = new_n2476_;
  assign n3138_li = new_n2478_;
  assign n3141_li = new_n5753_;
  assign n3168_li = new_n1868_;
  assign n3171_li = new_n2484_;
  assign n3174_li = new_n2486_;
  assign n3177_li = new_n2488_;
  assign n3180_li = new_n1870_;
  assign n3183_li = new_n2492_;
  assign n3192_li = new_n1872_;
  assign n3195_li = new_n2496_;
  assign n3204_li = new_n1874_;
  assign n3207_li = new_n2500_;
  assign n3216_li = new_n1876_;
  assign n3219_li = new_n2504_;
  assign n3228_li = new_n1878_;
  assign n3231_li = new_n2508_;
  assign n3240_li = new_n1880_;
  assign n3243_li = new_n2512_;
  assign n3252_li = new_n1882_;
  assign n3255_li = new_n2516_;
  assign n3258_li = new_n2518_;
  assign n3264_li = new_n1884_;
  assign n3267_li = new_n2522_;
  assign n3270_li = new_n2524_;
  assign n3276_li = new_n1886_;
  assign n3279_li = new_n2528_;
  assign n3282_li = new_n2530_;
  assign n3288_li = new_n1888_;
  assign n3291_li = new_n2534_;
  assign n3294_li = new_n2536_;
  assign n4537_i2 = new_n5327_;
  assign n4538_i2 = new_n5583_;
  assign n4710_i2 = new_n5568_;
  assign n4711_i2 = new_n5567_;
  assign n4803_i2 = new_n2610_;
  assign n4804_i2 = new_n2612_;
  assign n4843_i2 = new_n2650_;
  assign n4844_i2 = new_n2652_;
  assign n4927_i2 = new_n5564_;
  assign n4928_i2 = new_n5103_;
  assign n4945_i2 = new_n2674_;
  assign n4946_i2 = new_n2676_;
  assign n5009_i2 = new_n2686_;
  assign n5178_i2 = new_n5565_;
  assign n5179_i2 = new_n2800_;
  assign n5477_i2 = new_n5332_;
  assign n5478_i2 = new_n5322_;
  assign n5479_i2 = new_n5330_;
  assign n5222_i2 = new_n2806_;
  assign n5223_i2 = new_n5755_;
  assign n5553_i2 = new_n5467_;
  assign n5554_i2 = new_n5459_;
  assign G491_i2 = new_n5576_;
  assign n2922_lo_buf_i2 = new_n5594_;
  assign n2946_lo_buf_i2 = new_n5219_;
  assign n2970_lo_buf_i2 = new_n5425_;
  assign n2982_lo_buf_i2 = new_n5431_;
  assign n3066_lo_buf_i2 = new_n5407_;
  assign n3078_lo_buf_i2 = new_n5215_;
  assign n3102_lo_buf_i2 = new_n5422_;
  assign n3114_lo_buf_i2 = new_n5428_;
  assign G1321_i2 = new_n5542_;
  assign G1033_i2 = new_n5440_;
  assign G1030_i2 = new_n5433_;
  assign G1072_i2 = new_n5452_;
  assign G1159_i2 = n5553_i2;
  assign G1152_i2 = n5554_i2;
  assign n2958_lo_buf_i2 = new_n5756_;
  assign n2994_lo_buf_i2 = new_n5384_;
  assign n3006_lo_buf_i2 = new_n5402_;
  assign n3030_lo_buf_i2 = new_n5757_;
  assign n3042_lo_buf_i2 = new_n5696_;
  assign n3090_lo_buf_i2 = new_n5758_;
  assign G370_i2 = n2922_lo_buf_i2;
  assign G447_i2 = n2946_lo_buf_i2;
  assign G455_i2 = n2970_lo_buf_i2;
  assign G459_i2 = n2982_lo_buf_i2;
  assign G497_i2 = n3066_lo_buf_i2;
  assign G503_i2 = n3078_lo_buf_i2;
  assign G511_i2 = n3102_lo_buf_i2;
  assign G515_i2 = n3114_lo_buf_i2;
  assign G1036_i2 = new_n5471_;
  assign G1062_i2 = new_n5447_;
  assign G1067_i2 = new_n5450_;
  assign G1014_i2 = new_n5690_;
  assign G1171_i2 = new_n5442_;
  assign G1166_i2 = new_n5435_;
  assign n3018_lo_buf_i2 = new_n5759_;
  assign G766_i2 = G491_i2;
  assign G451_i2 = n2958_lo_buf_i2;
  assign G463_i2 = n2994_lo_buf_i2;
  assign G467_i2 = n3006_lo_buf_i2;
  assign G475_i2 = n3030_lo_buf_i2;
  assign G479_i2 = n3042_lo_buf_i2;
  assign G507_i2 = n3090_lo_buf_i2;
  assign G1017_i2 = new_n5762_;
  assign G1008_i2 = new_n5601_;
  assign G1176_i2 = new_n5472_;
  assign G1144_i2 = G1014_i2;
  assign n2910_lo_buf_i2 = new_n5699_;
  assign G471_i2 = n3018_lo_buf_i2;
  assign G2138_i2 = new_n5686_;
  assign G2147_i2 = new_n5693_;
  assign G1148_i2 = G1017_i2;
  assign G1137_i2 = G1008_i2;
  assign G1329_i2 = new_n5691_;
  assign G374_i2 = new_n5480_;
  assign G386_i2 = new_n5489_;
  assign G663_i2 = G374_i2;
  assign G674_i2 = G386_i2;
  assign G578_i2 = n3129_li;
  assign G575_i2 = n3141_li;
  assign G2505_i2 = ~new_n5585_;
  assign G2508_i2 = ~new_n5584_;
  assign G987_i2 = new_n5764_;
  assign G984_i2 = new_n5765_;
  assign G1862_i2 = new_n5335_;
  assign G1859_i2 = new_n5337_;
  assign G1260_i2 = new_n5766_;
  assign G1865_i2 = new_n5767_;
  assign G2073_i2 = new_n5768_;
  assign G1402_i2 = new_n5769_;
  assign G2048_i2 = new_n5770_;
  assign G2276_i2 = new_n5771_;
  assign G366_i2 = n2910_lo_buf_i2;
  assign G2141_i2 = ~new_n5603_;
  assign G2008_i2 = ~new_n5610_;
  assign G2011_i2 = ~new_n5614_;
  assign G2150_i2 = ~new_n5616_;
  assign G2026_i2 = ~new_n5620_;
  assign G2029_i2 = ~new_n5624_;
  assign G2023_i2 = ~new_n5631_;
  assign G2041_i2 = ~new_n5633_;
  assign G2017_i2 = new_n5640_;
  assign G2020_i2 = new_n5647_;
  assign G2035_i2 = new_n5649_;
  assign G2038_i2 = new_n5651_;
  assign G2228_i2 = ~new_n5655_;
  assign G2231_i2 = ~new_n5659_;
  assign G2234_i2 = ~new_n5663_;
  assign G2237_i2 = ~new_n5667_;
  assign G1904_i2 = ~new_n5608_;
  assign G1907_i2 = ~new_n5612_;
  assign G1928_i2 = ~new_n5618_;
  assign G1931_i2 = ~new_n5622_;
  assign G1893_i2 = new_n5639_;
  assign G1896_i2 = new_n5646_;
  assign G1899_i2 = ~new_n5630_;
  assign G1937_i2 = G1893_i2;
  assign G1940_i2 = G1896_i2;
  assign G1943_i2 = G1899_i2;
  assign G1336_i2 = new_n5761_;
  assign G1996_i2 = ~new_n5653_;
  assign G1999_i2 = ~new_n5657_;
  assign G2002_i2 = ~new_n5661_;
  assign G2005_i2 = ~new_n5665_;
  assign G2014_i2 = new_n5773_;
  assign G2032_i2 = new_n5775_;
  assign G1076_i2 = new_n5777_;
  assign G1002_i2 = new_n5701_;
  assign G998_i2 = new_n5779_;
  assign G1890_i2 = ~new_n5782_;
  assign G1934_i2 = G1890_i2;
  assign G1044_i2 = new_n5589_;
  assign G1039_i2 = ~new_n5586_;
  assign n1770_lo_buf_i2 = new_n2080_;
  assign G342_i2 = new_n5738_;
  assign G354_i2 = new_n5720_;
  assign G1193_i2 = new_n5588_;
  assign n3234_lo_buf_i2 = new_n5785_;
  assign n3246_lo_buf_i2 = new_n5786_;
  assign G783_i2 = new_n2626_;
  assign G786_i2 = new_n2628_;
  assign G792_i2 = new_n2630_;
  assign G795_i2 = new_n2632_;
  assign G815_i2 = new_n2634_;
  assign G818_i2 = new_n2636_;
  assign G824_i2 = new_n2638_;
  assign G827_i2 = new_n2640_;
  assign G789_i2 = new_n2658_;
  assign G798_i2 = new_n2660_;
  assign G801_i2 = new_n2662_;
  assign G807_i2 = new_n2664_;
  assign G812_i2 = new_n2666_;
  assign G821_i2 = new_n2668_;
  assign G804_i2 = new_n2680_;
  assign G780_i2 = new_n2728_;
  assign G1231_i2 = n5223_i2;
  assign G1572_i2 = G1321_i2;
  assign G1377_i2 = new_n5460_;
  assign G1253_i2 = ~new_n4053_;
  assign G1359_i2 = new_n4055_;
  assign G1258_i2 = ~new_n4072_;
  assign G1367_i2 = new_n4074_;
  assign G1358_i2 = new_n4076_;
  assign G1366_i2 = new_n4078_;
  assign G2057_i2 = ~new_n4089_;
  assign G2117_i2 = new_n4091_;
  assign G2118_i2 = ~new_n4093_;
  assign G1254_i2 = ~new_n4095_;
  assign G1259_i2 = ~new_n4097_;
  assign G2058_i2 = ~new_n4099_;
  assign G405_i2 = new_n5481_;
  assign G417_i2 = new_n5490_;
  assign G1269_i2 = new_n4102_;
  assign G1275_i2 = new_n4105_;
  assign G1287_i2 = new_n4108_;
  assign G1266_i2 = new_n4111_;
  assign G1272_i2 = new_n4114_;
  assign G1278_i2 = new_n4117_;
  assign G1281_i2 = new_n4120_;
  assign G1284_i2 = new_n4123_;
  assign G1290_i2 = new_n4126_;
  assign G1293_i2 = new_n4129_;
  assign G1299_i2 = new_n4132_;
  assign G1305_i2 = new_n4135_;
  assign G1296_i2 = new_n4138_;
  assign G1302_i2 = new_n4141_;
  assign G1308_i2 = new_n4144_;
  assign G1311_i2 = new_n4147_;
  assign G811_i2 = new_n5750_;
  assign G810_i2 = new_n5752_;
  assign G1728_i2 = new_n4150_;
  assign G2512_i2 = ~new_n4151_;
  assign G1114_i2 = G987_i2;
  assign G1113_i2 = G984_i2;
  assign G1992_i2 = new_n5334_;
  assign G1991_i2 = new_n5336_;
  assign G1426_i2 = G1260_i2;
  assign G1966_i2 = G1865_i2;
  assign G2211_i2 = G2073_i2;
  assign G1509_i2 = G1402_i2;
  assign G2153_i2 = G2048_i2;
  assign G2329_i2 = G2276_i2;
  assign G1540_i2 = new_n5763_;
  assign G2167_i2 = G2014_i2;
  assign G2191_i2 = G2032_i2;
  assign G1234_i2 = G1076_i2;
  assign G1132_i2 = new_n5703_;
  assign G1129_i2 = G998_i2;
  assign G2088_i2 = ~new_n5783_;
  assign G2106_i2 = G2088_i2;
  assign G1314_i2 = ~new_n5789_;
  assign G636_i2 = G342_i2;
  assign G647_i2 = G354_i2;
  assign n3186_lo_buf_i2 = new_n2494_;
  assign n3198_lo_buf_i2 = new_n2498_;
  assign n3210_lo_buf_i2 = new_n2502_;
  assign n3222_lo_buf_i2 = new_n2506_;
  assign G1225_i2 = new_n5451_;
  assign G1342_i2 = new_n5466_;
  assign G1222_i2 = new_n5446_;
  assign G1228_i2 = new_n5449_;
  assign G1348_i2 = G1171_i2;
  assign G1345_i2 = G1166_i2;
  assign G1351_i2 = G1176_i2;
  assign G2242_i2 = new_n4161_;
  assign G2260_i2 = new_n4168_;
  assign G1374_i2 = new_n5600_;
  assign G1537_i2 = G1329_i2;
  assign G301_i2 = new_n5739_;
  assign G313_i2 = new_n5721_;
  assign G2365_i2 = ~new_n4169_;
  assign G2255_i2 = ~new_n4170_;
  assign G2253_i2 = ~new_n4171_;
  assign G2395_i2 = ~new_n4172_;
  assign G2272_i2 = ~new_n4173_;
  assign G2270_i2 = ~new_n4174_;
  assign G2245_i2 = ~new_n4175_;
  assign G2262_i2 = ~new_n4176_;
  assign G2249_i2 = new_n4177_;
  assign G2247_i2 = new_n4178_;
  assign G2266_i2 = new_n4179_;
  assign G2264_i2 = new_n4180_;
  assign G2403_i2 = ~new_n4181_;
  assign G2401_i2 = ~new_n4182_;
  assign G2410_i2 = ~new_n4183_;
  assign G2408_i2 = ~new_n4184_;
  assign G2306_i2 = ~new_n4185_;
  assign G2305_i2 = ~new_n4186_;
  assign G2314_i2 = ~new_n4187_;
  assign G2313_i2 = ~new_n4188_;
  assign G2303_i2 = new_n4189_;
  assign G2302_i2 = new_n4190_;
  assign G2301_i2 = ~new_n4191_;
  assign G2311_i2 = new_n4192_;
  assign G2310_i2 = new_n4193_;
  assign G2309_i2 = ~new_n4194_;
  assign G2404_i2 = ~new_n4195_;
  assign G2411_i2 = ~new_n4196_;
  assign G2420_i2 = ~new_n4197_;
  assign G2419_i2 = ~new_n4198_;
  assign G2433_i2 = ~new_n4199_;
  assign G2432_i2 = ~new_n4200_;
  assign G402_i2 = n3234_lo_buf_i2;
  assign G403_i2 = n3246_lo_buf_i2;
  assign G1053_i2 = new_n4211_;
  assign G1049_i2 = new_n4222_;
  assign G1058_i2 = new_n4229_;
  assign G1364_i2 = new_n5754_;
  assign G1079_i2 = new_n4240_;
  assign G1478_i2 = G1377_i2;
  assign G707_i2 = G405_i2;
  assign G718_i2 = G417_i2;
  assign G2417_i2 = new_n4243_;
  assign G2414_i2 = new_n4246_;
  assign G2431_i2 = new_n4249_;
  assign G2428_i2 = new_n4252_;
  assign G1653_i2 = G1540_i2;
  assign G2213_i2 = new_n4256_;
  assign G2221_i2 = new_n4260_;
  assign G2250_i2 = new_n5772_;
  assign G2267_i2 = new_n5774_;
  assign G1365_i2 = new_n5776_;
  assign G1368_i2 = G1132_i2;
  assign G1371_i2 = new_n5778_;
  assign G2218_i2 = ~new_n5784_;
  assign G2225_i2 = G2218_i2;
  assign n1503_lo_buf_i2 = new_n1940_;
  assign n1863_lo_buf_i2 = new_n2104_;
  assign n1887_lo_buf_i2 = new_n2108_;
  assign n1983_lo_buf_i2 = new_n2134_;
  assign n2007_lo_buf_i2 = new_n2138_;
  assign n2115_lo_buf_i2 = new_n2166_;
  assign n2139_lo_buf_i2 = new_n2170_;
  assign n2247_lo_buf_i2 = new_n2198_;
  assign n2271_lo_buf_i2 = new_n2202_;
  assign n2919_lo_buf_i2 = new_n2406_;
  assign n2943_lo_buf_i2 = new_n2410_;
  assign n2967_lo_buf_i2 = new_n2416_;
  assign n2979_lo_buf_i2 = new_n2418_;
  assign n3063_lo_buf_i2 = new_n2448_;
  assign n3075_lo_buf_i2 = new_n2450_;
  assign n3099_lo_buf_i2 = new_n2460_;
  assign n3111_lo_buf_i2 = new_n2464_;
  assign G878_i2 = new_n4262_;
  assign G875_i2 = new_n4264_;
  assign G661_i2 = new_n4266_;
  assign G660_i2 = new_n4268_;
  assign G879_i2 = new_n4270_;
  assign G876_i2 = new_n4271_;
  assign G1320_i2 = ~new_n5587_;
  assign G941_i2 = new_n4273_;
  assign G732_i2 = new_n4275_;
  assign G942_i2 = new_n4277_;
  assign G1493_i2 = G1314_i2;
  assign G1498_i2 = ~new_n5788_;
  assign G877_i2 = new_n4279_;
  assign G874_i2 = new_n4281_;
  assign n1806_lo_buf_i2 = new_n2094_;
  assign n1878_lo_buf_i2 = new_n2106_;
  assign n1938_lo_buf_i2 = new_n2126_;
  assign n1998_lo_buf_i2 = new_n2136_;
  assign n2058_lo_buf_i2 = new_n2156_;
  assign n2130_lo_buf_i2 = new_n2168_;
  assign n2190_lo_buf_i2 = new_n2188_;
  assign n2262_lo_buf_i2 = new_n2200_;
  assign n2310_lo_buf_i2 = new_n2216_;
  assign n2406_lo_buf_i2 = new_n2240_;
  assign n2430_lo_buf_i2 = new_n2246_;
  assign n2526_lo_buf_i2 = new_n2270_;
  assign n2550_lo_buf_i2 = new_n2276_;
  assign n2646_lo_buf_i2 = new_n2300_;
  assign n2670_lo_buf_i2 = new_n2306_;
  assign n2766_lo_buf_i2 = new_n2330_;
  assign G603_i2 = G301_i2;
  assign G614_i2 = G313_i2;
  assign G1026_i2 = new_n4292_;
  assign G1021_i2 = new_n4303_;
  assign G940_i2 = new_n4305_;
  assign G1636_i2 = ~new_n5790_;
  assign G1684_i2 = G1636_i2;
  assign n2352_lo_buf_i2 = new_n1732_;
  assign n2364_lo_buf_i2 = new_n1734_;
  assign n2472_lo_buf_i2 = new_n1752_;
  assign n2484_lo_buf_i2 = new_n1754_;
  assign n2592_lo_buf_i2 = new_n1772_;
  assign n2604_lo_buf_i2 = new_n1774_;
  assign n2712_lo_buf_i2 = new_n1792_;
  assign n2724_lo_buf_i2 = new_n1794_;
  assign n3150_lo_buf_i2 = new_n1864_;
  assign n3162_lo_buf_i2 = new_n1866_;
  assign new_n5047_ = new_n2377_;
  assign new_n5048_ = new_n2343_;
  assign new_n5049_ = new_n5048_;
  assign new_n5050_ = new_n5048_;
  assign new_n5051_ = new_n3250_;
  assign new_n5052_ = new_n5051_;
  assign new_n5053_ = new_n2285_;
  assign new_n5054_ = new_n2125_;
  assign new_n5055_ = new_n2255_;
  assign new_n5056_ = new_n2155_;
  assign new_n5057_ = new_n2315_;
  assign new_n5058_ = new_n2187_;
  assign new_n5059_ = new_n2225_;
  assign new_n5060_ = new_n2093_;
  assign new_n5061_ = new_n3258_;
  assign new_n5062_ = new_n3255_;
  assign new_n5063_ = new_n2384_;
  assign new_n5064_ = new_n5063_;
  assign new_n5065_ = new_n2385_;
  assign new_n5066_ = new_n5065_;
  assign new_n5067_ = new_n3265_;
  assign new_n5068_ = new_n3262_;
  assign new_n5069_ = new_n5068_;
  assign new_n5070_ = new_n5068_;
  assign new_n5071_ = new_n2392_;
  assign new_n5072_ = new_n5071_;
  assign new_n5073_ = new_n5072_;
  assign new_n5074_ = new_n5071_;
  assign new_n5075_ = new_n2564_;
  assign new_n5076_ = new_n2393_;
  assign new_n5077_ = new_n5076_;
  assign new_n5078_ = new_n5077_;
  assign new_n5079_ = new_n5076_;
  assign new_n5080_ = new_n2562_;
  assign new_n5081_ = new_n2547_;
  assign new_n5082_ = new_n3283_;
  assign new_n5083_ = new_n2571_;
  assign new_n5084_ = new_n3287_;
  assign new_n5085_ = new_n1949_;
  assign new_n5086_ = new_n2925_;
  assign new_n5087_ = new_n2856_;
  assign new_n5088_ = new_n2924_;
  assign new_n5089_ = new_n2857_;
  assign new_n5090_ = new_n2568_;
  assign new_n5091_ = new_n5090_;
  assign new_n5092_ = new_n2079_;
  assign new_n5093_ = new_n2926_;
  assign new_n5094_ = new_n3434_;
  assign new_n5095_ = new_n3412_;
  assign new_n5096_ = new_n3310_;
  assign new_n5097_ = new_n3325_;
  assign new_n5098_ = new_n3295_;
  assign new_n5099_ = new_n3437_;
  assign new_n5100_ = new_n2673_;
  assign new_n5101_ = new_n2672_;
  assign new_n5102_ = new_n5101_;
  assign new_n5103_ = new_n5101_;
  assign new_n5104_ = new_n2966_;
  assign new_n5105_ = new_n2968_;
  assign new_n5106_ = new_n2813_;
  assign new_n5107_ = new_n2815_;
  assign new_n5108_ = new_n3084_;
  assign new_n5109_ = new_n5108_;
  assign new_n5110_ = new_n5109_;
  assign new_n5111_ = new_n5109_;
  assign new_n5112_ = new_n5108_;
  assign new_n5113_ = new_n5112_;
  assign new_n5114_ = new_n5112_;
  assign new_n5115_ = new_n3086_;
  assign new_n5116_ = new_n5115_;
  assign new_n5117_ = new_n5116_;
  assign new_n5118_ = new_n5116_;
  assign new_n5119_ = new_n5115_;
  assign new_n5120_ = new_n5119_;
  assign new_n5121_ = new_n5119_;
  assign new_n5122_ = new_n2885_;
  assign new_n5123_ = new_n5122_;
  assign new_n5124_ = new_n5123_;
  assign new_n5125_ = new_n5123_;
  assign new_n5126_ = new_n5122_;
  assign new_n5127_ = new_n5126_;
  assign new_n5128_ = new_n5126_;
  assign new_n5129_ = new_n2887_;
  assign new_n5130_ = new_n5129_;
  assign new_n5131_ = new_n5130_;
  assign new_n5132_ = new_n5130_;
  assign new_n5133_ = new_n5129_;
  assign new_n5134_ = new_n5133_;
  assign new_n5135_ = new_n5133_;
  assign new_n5136_ = new_n3210_;
  assign new_n5137_ = new_n5136_;
  assign new_n5138_ = new_n5137_;
  assign new_n5139_ = new_n5138_;
  assign new_n5140_ = new_n5138_;
  assign new_n5141_ = new_n5137_;
  assign new_n5142_ = new_n5136_;
  assign new_n5143_ = new_n5142_;
  assign new_n5144_ = new_n5142_;
  assign new_n5145_ = new_n3211_;
  assign new_n5146_ = new_n5145_;
  assign new_n5147_ = new_n5146_;
  assign new_n5148_ = new_n5146_;
  assign new_n5149_ = new_n5145_;
  assign new_n5150_ = new_n3212_;
  assign new_n5151_ = new_n5150_;
  assign new_n5152_ = new_n5151_;
  assign new_n5153_ = new_n5152_;
  assign new_n5154_ = new_n5152_;
  assign new_n5155_ = new_n5151_;
  assign new_n5156_ = new_n5150_;
  assign new_n5157_ = new_n5156_;
  assign new_n5158_ = new_n5156_;
  assign new_n5159_ = new_n3213_;
  assign new_n5160_ = new_n5159_;
  assign new_n5161_ = new_n5160_;
  assign new_n5162_ = new_n5160_;
  assign new_n5163_ = new_n5159_;
  assign new_n5164_ = new_n3001_;
  assign new_n5165_ = new_n5164_;
  assign new_n5166_ = new_n5165_;
  assign new_n5167_ = new_n5166_;
  assign new_n5168_ = new_n5166_;
  assign new_n5169_ = new_n5165_;
  assign new_n5170_ = new_n5164_;
  assign new_n5171_ = new_n5170_;
  assign new_n5172_ = new_n5170_;
  assign new_n5173_ = new_n3000_;
  assign new_n5174_ = new_n5173_;
  assign new_n5175_ = new_n5174_;
  assign new_n5176_ = new_n5174_;
  assign new_n5177_ = new_n5173_;
  assign new_n5178_ = new_n3003_;
  assign new_n5179_ = new_n5178_;
  assign new_n5180_ = new_n5179_;
  assign new_n5181_ = new_n5180_;
  assign new_n5182_ = new_n5180_;
  assign new_n5183_ = new_n5179_;
  assign new_n5184_ = new_n5178_;
  assign new_n5185_ = new_n5184_;
  assign new_n5186_ = new_n5184_;
  assign new_n5187_ = new_n3002_;
  assign new_n5188_ = new_n5187_;
  assign new_n5189_ = new_n5188_;
  assign new_n5190_ = new_n5188_;
  assign new_n5191_ = new_n5187_;
  assign new_n5192_ = new_n3220_;
  assign new_n5193_ = new_n5192_;
  assign new_n5194_ = new_n5193_;
  assign new_n5195_ = new_n5194_;
  assign new_n5196_ = new_n5194_;
  assign new_n5197_ = new_n5193_;
  assign new_n5198_ = new_n5197_;
  assign new_n5199_ = new_n5192_;
  assign new_n5200_ = new_n5199_;
  assign new_n5201_ = new_n5199_;
  assign new_n5202_ = new_n3145_;
  assign new_n5203_ = new_n3221_;
  assign new_n5204_ = new_n5203_;
  assign new_n5205_ = new_n5204_;
  assign new_n5206_ = new_n5205_;
  assign new_n5207_ = new_n5205_;
  assign new_n5208_ = new_n5204_;
  assign new_n5209_ = new_n5208_;
  assign new_n5210_ = new_n5203_;
  assign new_n5211_ = new_n5210_;
  assign new_n5212_ = new_n5210_;
  assign new_n5213_ = new_n3144_;
  assign new_n5214_ = new_n5213_;
  assign new_n5215_ = new_n5213_;
  assign new_n5216_ = new_n3137_;
  assign new_n5217_ = new_n3136_;
  assign new_n5218_ = new_n5217_;
  assign new_n5219_ = new_n5217_;
  assign new_n5220_ = new_n3222_;
  assign new_n5221_ = new_n5220_;
  assign new_n5222_ = new_n5221_;
  assign new_n5223_ = new_n5222_;
  assign new_n5224_ = new_n5222_;
  assign new_n5225_ = new_n5221_;
  assign new_n5226_ = new_n5225_;
  assign new_n5227_ = new_n5220_;
  assign new_n5228_ = new_n5227_;
  assign new_n5229_ = new_n5227_;
  assign new_n5230_ = new_n3223_;
  assign new_n5231_ = new_n5230_;
  assign new_n5232_ = new_n5231_;
  assign new_n5233_ = new_n5232_;
  assign new_n5234_ = new_n5232_;
  assign new_n5235_ = new_n5231_;
  assign new_n5236_ = new_n5235_;
  assign new_n5237_ = new_n5230_;
  assign new_n5238_ = new_n5237_;
  assign new_n5239_ = new_n5237_;
  assign new_n5240_ = new_n3567_;
  assign new_n5241_ = new_n5240_;
  assign new_n5242_ = new_n5240_;
  assign new_n5243_ = new_n3570_;
  assign new_n5244_ = new_n5243_;
  assign new_n5245_ = new_n3574_;
  assign new_n5246_ = new_n3585_;
  assign new_n5247_ = new_n5246_;
  assign new_n5248_ = new_n5247_;
  assign new_n5249_ = new_n5246_;
  assign new_n5250_ = new_n3584_;
  assign new_n5251_ = new_n5250_;
  assign new_n5252_ = new_n5251_;
  assign new_n5253_ = new_n5250_;
  assign new_n5254_ = new_n3591_;
  assign new_n5255_ = new_n5254_;
  assign new_n5256_ = new_n5254_;
  assign new_n5257_ = new_n3590_;
  assign new_n5258_ = new_n5257_;
  assign new_n5259_ = new_n5257_;
  assign new_n5260_ = new_n3599_;
  assign new_n5261_ = new_n5260_;
  assign new_n5262_ = new_n3598_;
  assign new_n5263_ = new_n5262_;
  assign new_n5264_ = new_n2782_;
  assign new_n5265_ = new_n2783_;
  assign new_n5266_ = new_n3609_;
  assign new_n5267_ = new_n3608_;
  assign new_n5268_ = new_n2690_;
  assign new_n5269_ = new_n5268_;
  assign new_n5270_ = new_n2691_;
  assign new_n5271_ = new_n5270_;
  assign new_n5272_ = new_n3091_;
  assign new_n5273_ = new_n3090_;
  assign new_n5274_ = new_n3581_;
  assign new_n5275_ = new_n3665_;
  assign new_n5276_ = new_n5275_;
  assign new_n5277_ = new_n5275_;
  assign new_n5278_ = new_n3668_;
  assign new_n5279_ = new_n5278_;
  assign new_n5280_ = new_n3672_;
  assign new_n5281_ = new_n3683_;
  assign new_n5282_ = new_n5281_;
  assign new_n5283_ = new_n5282_;
  assign new_n5284_ = new_n5281_;
  assign new_n5285_ = new_n3682_;
  assign new_n5286_ = new_n5285_;
  assign new_n5287_ = new_n5286_;
  assign new_n5288_ = new_n5285_;
  assign new_n5289_ = new_n3689_;
  assign new_n5290_ = new_n5289_;
  assign new_n5291_ = new_n5289_;
  assign new_n5292_ = new_n3688_;
  assign new_n5293_ = new_n5292_;
  assign new_n5294_ = new_n5292_;
  assign new_n5295_ = new_n3697_;
  assign new_n5296_ = new_n5295_;
  assign new_n5297_ = new_n3696_;
  assign new_n5298_ = new_n5297_;
  assign new_n5299_ = new_n3707_;
  assign new_n5300_ = new_n3706_;
  assign new_n5301_ = new_n3095_;
  assign new_n5302_ = new_n3094_;
  assign new_n5303_ = new_n3679_;
  assign new_n5304_ = new_n2988_;
  assign new_n5305_ = new_n2981_;
  assign new_n5306_ = new_n2989_;
  assign new_n5307_ = new_n2980_;
  assign new_n5308_ = new_n2990_;
  assign new_n5309_ = new_n2987_;
  assign new_n5310_ = new_n2991_;
  assign new_n5311_ = new_n2986_;
  assign new_n5312_ = new_n2526_;
  assign new_n5313_ = new_n2521_;
  assign new_n5314_ = new_n2527_;
  assign new_n5315_ = new_n2520_;
  assign new_n5316_ = new_n2679_;
  assign new_n5317_ = new_n2586_;
  assign new_n5318_ = new_n2678_;
  assign new_n5319_ = new_n2587_;
  assign new_n5320_ = new_n3074_;
  assign new_n5321_ = new_n5320_;
  assign new_n5322_ = new_n5320_;
  assign new_n5323_ = new_n2577_;
  assign new_n5324_ = new_n3075_;
  assign new_n5325_ = new_n2576_;
  assign new_n5326_ = new_n5325_;
  assign new_n5327_ = new_n5325_;
  assign new_n5328_ = new_n3077_;
  assign new_n5329_ = new_n3073_;
  assign new_n5330_ = new_n3076_;
  assign new_n5331_ = new_n5330_;
  assign new_n5332_ = new_n3072_;
  assign new_n5333_ = new_n5332_;
  assign new_n5334_ = new_n3773_;
  assign new_n5335_ = new_n5334_;
  assign new_n5336_ = new_n3779_;
  assign new_n5337_ = new_n5336_;
  assign new_n5338_ = new_n2972_;
  assign new_n5339_ = new_n2971_;
  assign new_n5340_ = new_n2973_;
  assign new_n5341_ = new_n2970_;
  assign new_n5342_ = new_n2976_;
  assign new_n5343_ = new_n2975_;
  assign new_n5344_ = new_n2977_;
  assign new_n5345_ = new_n2974_;
  assign new_n5346_ = new_n3824_;
  assign new_n5347_ = new_n3817_;
  assign new_n5348_ = new_n3829_;
  assign new_n5349_ = new_n3818_;
  assign new_n5350_ = new_n3830_;
  assign new_n5351_ = new_n3823_;
  assign new_n5352_ = new_n3080_;
  assign new_n5353_ = new_n2982_;
  assign new_n5354_ = new_n3081_;
  assign new_n5355_ = new_n2983_;
  assign new_n5356_ = new_n2985_;
  assign new_n5357_ = new_n2978_;
  assign new_n5358_ = new_n2984_;
  assign new_n5359_ = new_n2979_;
  assign new_n5360_ = new_n3852_;
  assign new_n5361_ = new_n3847_;
  assign new_n5362_ = new_n3859_;
  assign new_n5363_ = new_n3846_;
  assign new_n5364_ = new_n3858_;
  assign new_n5365_ = new_n3853_;
  assign new_n5366_ = new_n3110_;
  assign new_n5367_ = new_n3109_;
  assign new_n5368_ = new_n3111_;
  assign new_n5369_ = new_n3108_;
  assign new_n5370_ = new_n2998_;
  assign new_n5371_ = new_n2996_;
  assign new_n5372_ = new_n2999_;
  assign new_n5373_ = new_n2997_;
  assign new_n5374_ = new_n3882_;
  assign new_n5375_ = new_n3875_;
  assign new_n5376_ = new_n3887_;
  assign new_n5377_ = new_n3876_;
  assign new_n5378_ = new_n3888_;
  assign new_n5379_ = new_n3881_;
  assign new_n5380_ = new_n2457_;
  assign new_n5381_ = new_n2415_;
  assign new_n5382_ = new_n2422_;
  assign new_n5383_ = new_n5382_;
  assign new_n5384_ = new_n5382_;
  assign new_n5385_ = new_n3117_;
  assign new_n5386_ = new_n5385_;
  assign new_n5387_ = new_n5386_;
  assign new_n5388_ = new_n5387_;
  assign new_n5389_ = new_n5387_;
  assign new_n5390_ = new_n5386_;
  assign new_n5391_ = new_n5390_;
  assign new_n5392_ = new_n5390_;
  assign new_n5393_ = new_n5385_;
  assign new_n5394_ = new_n5393_;
  assign new_n5395_ = new_n5394_;
  assign new_n5396_ = new_n5394_;
  assign new_n5397_ = new_n5393_;
  assign new_n5398_ = new_n5397_;
  assign new_n5399_ = new_n5397_;
  assign new_n5400_ = new_n2426_;
  assign new_n5401_ = new_n5400_;
  assign new_n5402_ = new_n5400_;
  assign new_n5403_ = new_n3142_;
  assign new_n5404_ = new_n5403_;
  assign new_n5405_ = new_n5404_;
  assign new_n5406_ = new_n5404_;
  assign new_n5407_ = new_n5403_;
  assign new_n5408_ = new_n3918_;
  assign new_n5409_ = new_n5408_;
  assign new_n5410_ = new_n5408_;
  assign new_n5411_ = new_n2435_;
  assign new_n5412_ = new_n3917_;
  assign new_n5413_ = new_n5412_;
  assign new_n5414_ = new_n5413_;
  assign new_n5415_ = new_n5413_;
  assign new_n5416_ = new_n5412_;
  assign new_n5417_ = new_n5416_;
  assign new_n5418_ = new_n5416_;
  assign new_n5419_ = new_n2439_;
  assign new_n5420_ = new_n3146_;
  assign new_n5421_ = new_n5420_;
  assign new_n5422_ = new_n5420_;
  assign new_n5423_ = new_n3138_;
  assign new_n5424_ = new_n5423_;
  assign new_n5425_ = new_n5423_;
  assign new_n5426_ = new_n3148_;
  assign new_n5427_ = new_n5426_;
  assign new_n5428_ = new_n5426_;
  assign new_n5429_ = new_n3140_;
  assign new_n5430_ = new_n5429_;
  assign new_n5431_ = new_n5429_;
  assign new_n5432_ = new_n3451_;
  assign new_n5433_ = new_n5432_;
  assign new_n5434_ = new_n5433_;
  assign new_n5435_ = new_n5432_;
  assign new_n5436_ = new_n3171_;
  assign new_n5437_ = new_n5436_;
  assign new_n5438_ = new_n5436_;
  assign new_n5439_ = new_n3448_;
  assign new_n5440_ = new_n5439_;
  assign new_n5441_ = new_n5440_;
  assign new_n5442_ = new_n5439_;
  assign new_n5443_ = new_n3173_;
  assign new_n5444_ = new_n5443_;
  assign new_n5445_ = new_n5443_;
  assign new_n5446_ = new_n3476_;
  assign new_n5447_ = new_n5446_;
  assign new_n5448_ = new_n2965_;
  assign new_n5449_ = new_n3487_;
  assign new_n5450_ = new_n5449_;
  assign new_n5451_ = new_n3454_;
  assign new_n5452_ = new_n5451_;
  assign new_n5453_ = new_n2964_;
  assign new_n5454_ = new_n3216_;
  assign new_n5455_ = new_n5454_;
  assign new_n5456_ = new_n5455_;
  assign new_n5457_ = new_n5455_;
  assign new_n5458_ = new_n5454_;
  assign new_n5459_ = new_n5458_;
  assign new_n5460_ = new_n5458_;
  assign new_n5461_ = new_n3170_;
  assign new_n5462_ = new_n3214_;
  assign new_n5463_ = new_n5462_;
  assign new_n5464_ = new_n5463_;
  assign new_n5465_ = new_n5463_;
  assign new_n5466_ = new_n5462_;
  assign new_n5467_ = new_n5466_;
  assign new_n5468_ = new_n3172_;
  assign new_n5469_ = new_n2431_;
  assign new_n5470_ = new_n3465_;
  assign new_n5471_ = new_n5470_;
  assign new_n5472_ = new_n5470_;
  assign new_n5473_ = new_n3240_;
  assign new_n5474_ = new_n5473_;
  assign new_n5475_ = new_n5474_;
  assign new_n5476_ = new_n5475_;
  assign new_n5477_ = new_n5475_;
  assign new_n5478_ = new_n5474_;
  assign new_n5479_ = new_n5473_;
  assign new_n5480_ = new_n5479_;
  assign new_n5481_ = new_n5479_;
  assign new_n5482_ = new_n3242_;
  assign new_n5483_ = new_n5482_;
  assign new_n5484_ = new_n5483_;
  assign new_n5485_ = new_n5484_;
  assign new_n5486_ = new_n5484_;
  assign new_n5487_ = new_n5483_;
  assign new_n5488_ = new_n5482_;
  assign new_n5489_ = new_n5488_;
  assign new_n5490_ = new_n5488_;
  assign new_n5491_ = new_n3241_;
  assign new_n5492_ = new_n5491_;
  assign new_n5493_ = new_n5492_;
  assign new_n5494_ = new_n5492_;
  assign new_n5495_ = new_n5491_;
  assign new_n5496_ = new_n3243_;
  assign new_n5497_ = new_n5496_;
  assign new_n5498_ = new_n5497_;
  assign new_n5499_ = new_n5497_;
  assign new_n5500_ = new_n5496_;
  assign new_n5501_ = new_n2615_;
  assign new_n5502_ = new_n2590_;
  assign new_n5503_ = new_n2614_;
  assign new_n5504_ = new_n2591_;
  assign new_n5505_ = new_n2588_;
  assign new_n5506_ = new_n2532_;
  assign new_n5507_ = new_n2589_;
  assign new_n5508_ = new_n2533_;
  assign new_n5509_ = new_n4047_;
  assign new_n5510_ = new_n4041_;
  assign new_n5511_ = new_n4051_;
  assign new_n5512_ = new_n5511_;
  assign new_n5513_ = new_n5511_;
  assign new_n5514_ = new_n4048_;
  assign new_n5515_ = new_n2624_;
  assign new_n5516_ = new_n5515_;
  assign new_n5517_ = new_n2597_;
  assign new_n5518_ = new_n2625_;
  assign new_n5519_ = new_n2596_;
  assign new_n5520_ = new_n5519_;
  assign new_n5521_ = new_n2594_;
  assign new_n5522_ = new_n2538_;
  assign new_n5523_ = new_n2595_;
  assign new_n5524_ = new_n2539_;
  assign new_n5525_ = new_n2600_;
  assign new_n5526_ = new_n2598_;
  assign new_n5527_ = new_n4066_;
  assign new_n5528_ = new_n4060_;
  assign new_n5529_ = new_n4070_;
  assign new_n5530_ = new_n5529_;
  assign new_n5531_ = new_n5529_;
  assign new_n5532_ = new_n4067_;
  assign new_n5533_ = new_n4042_;
  assign new_n5534_ = new_n4061_;
  assign new_n5535_ = new_n2958_;
  assign new_n5536_ = new_n2957_;
  assign new_n5537_ = new_n2959_;
  assign new_n5538_ = new_n2956_;
  assign new_n5539_ = new_n4083_;
  assign new_n5540_ = new_n3445_;
  assign new_n5541_ = new_n5540_;
  assign new_n5542_ = new_n5540_;
  assign new_n5543_ = new_n4087_;
  assign new_n5544_ = new_n5543_;
  assign new_n5545_ = new_n5543_;
  assign new_n5546_ = new_n4084_;
  assign new_n5547_ = new_n3444_;
  assign new_n5548_ = new_n1970_;
  assign new_n5549_ = new_n5548_;
  assign new_n5550_ = new_n5549_;
  assign new_n5551_ = new_n5550_;
  assign new_n5552_ = new_n5549_;
  assign new_n5553_ = new_n5548_;
  assign new_n5554_ = new_n5553_;
  assign new_n5555_ = new_n5553_;
  assign new_n5556_ = new_n1971_;
  assign new_n5557_ = new_n5556_;
  assign new_n5558_ = new_n5557_;
  assign new_n5559_ = new_n5558_;
  assign new_n5560_ = new_n5557_;
  assign new_n5561_ = new_n5556_;
  assign new_n5562_ = new_n5561_;
  assign new_n5563_ = new_n5561_;
  assign new_n5564_ = new_n2670_;
  assign new_n5565_ = new_n2798_;
  assign new_n5566_ = new_n5565_;
  assign new_n5567_ = new_n2582_;
  assign new_n5568_ = new_n2580_;
  assign new_n5569_ = new_n2038_;
  assign new_n5570_ = new_n5569_;
  assign new_n5571_ = new_n5570_;
  assign new_n5572_ = new_n5571_;
  assign new_n5573_ = new_n5570_;
  assign new_n5574_ = new_n5569_;
  assign new_n5575_ = new_n5574_;
  assign new_n5576_ = new_n5574_;
  assign new_n5577_ = new_n2039_;
  assign new_n5578_ = new_n5577_;
  assign new_n5579_ = new_n5578_;
  assign new_n5580_ = new_n5578_;
  assign new_n5581_ = new_n5577_;
  assign new_n5582_ = new_n5581_;
  assign new_n5583_ = new_n2578_;
  assign new_n5584_ = new_n3761_;
  assign new_n5585_ = new_n3663_;
  assign new_n5586_ = new_n4036_;
  assign new_n5587_ = new_n4152_;
  assign new_n5588_ = new_n4025_;
  assign new_n5589_ = new_n5588_;
  assign new_n5590_ = new_n3143_;
  assign new_n5591_ = new_n3135_;
  assign new_n5592_ = new_n3134_;
  assign new_n5593_ = new_n5592_;
  assign new_n5594_ = new_n5592_;
  assign new_n5595_ = new_n4159_;
  assign new_n5596_ = new_n3553_;
  assign new_n5597_ = new_n5596_;
  assign new_n5598_ = new_n5597_;
  assign new_n5599_ = new_n5597_;
  assign new_n5600_ = new_n5596_;
  assign new_n5601_ = new_n5600_;
  assign new_n5602_ = new_n4166_;
  assign new_n5603_ = new_n3902_;
  assign new_n5604_ = new_n5603_;
  assign new_n5605_ = new_n3530_;
  assign new_n5606_ = new_n5605_;
  assign new_n5607_ = new_n5605_;
  assign new_n5608_ = new_n3947_;
  assign new_n5609_ = new_n5608_;
  assign new_n5610_ = new_n3904_;
  assign new_n5611_ = new_n5610_;
  assign new_n5612_ = new_n3949_;
  assign new_n5613_ = new_n5612_;
  assign new_n5614_ = new_n3906_;
  assign new_n5615_ = new_n5614_;
  assign new_n5616_ = new_n3909_;
  assign new_n5617_ = new_n5616_;
  assign new_n5618_ = new_n3951_;
  assign new_n5619_ = new_n5618_;
  assign new_n5620_ = new_n3911_;
  assign new_n5621_ = new_n5620_;
  assign new_n5622_ = new_n3953_;
  assign new_n5623_ = new_n5622_;
  assign new_n5624_ = new_n3913_;
  assign new_n5625_ = new_n5624_;
  assign new_n5626_ = new_n3959_;
  assign new_n5627_ = new_n5626_;
  assign new_n5628_ = new_n5627_;
  assign new_n5629_ = new_n5627_;
  assign new_n5630_ = new_n5626_;
  assign new_n5631_ = new_n3919_;
  assign new_n5632_ = new_n5631_;
  assign new_n5633_ = new_n3921_;
  assign new_n5634_ = new_n5633_;
  assign new_n5635_ = new_n3955_;
  assign new_n5636_ = new_n5635_;
  assign new_n5637_ = new_n5636_;
  assign new_n5638_ = new_n5636_;
  assign new_n5639_ = new_n5635_;
  assign new_n5640_ = new_n3923_;
  assign new_n5641_ = new_n5640_;
  assign new_n5642_ = new_n3957_;
  assign new_n5643_ = new_n5642_;
  assign new_n5644_ = new_n5643_;
  assign new_n5645_ = new_n5643_;
  assign new_n5646_ = new_n5642_;
  assign new_n5647_ = new_n3925_;
  assign new_n5648_ = new_n5647_;
  assign new_n5649_ = new_n3927_;
  assign new_n5650_ = new_n5649_;
  assign new_n5651_ = new_n3929_;
  assign new_n5652_ = new_n5651_;
  assign new_n5653_ = new_n3963_;
  assign new_n5654_ = new_n5653_;
  assign new_n5655_ = new_n3933_;
  assign new_n5656_ = new_n5655_;
  assign new_n5657_ = new_n3967_;
  assign new_n5658_ = new_n5657_;
  assign new_n5659_ = new_n3937_;
  assign new_n5660_ = new_n5659_;
  assign new_n5661_ = new_n3971_;
  assign new_n5662_ = new_n5661_;
  assign new_n5663_ = new_n3941_;
  assign new_n5664_ = new_n5663_;
  assign new_n5665_ = new_n3975_;
  assign new_n5666_ = new_n5665_;
  assign new_n5667_ = new_n3945_;
  assign new_n5668_ = new_n5667_;
  assign new_n5669_ = new_n2696_;
  assign new_n5670_ = new_n5669_;
  assign new_n5671_ = new_n5669_;
  assign new_n5672_ = new_n2698_;
  assign new_n5673_ = new_n5672_;
  assign new_n5674_ = new_n5672_;
  assign new_n5675_ = new_n2693_;
  assign new_n5676_ = new_n5675_;
  assign new_n5677_ = new_n5675_;
  assign new_n5678_ = new_n2695_;
  assign new_n5679_ = new_n5678_;
  assign new_n5680_ = new_n5678_;
  assign new_n5681_ = new_n2699_;
  assign new_n5682_ = new_n2697_;
  assign new_n5683_ = new_n2692_;
  assign new_n5684_ = new_n2694_;
  assign new_n5685_ = new_n3552_;
  assign new_n5686_ = new_n3558_;
  assign new_n5687_ = new_n3509_;
  assign new_n5688_ = new_n5687_;
  assign new_n5689_ = new_n5688_;
  assign new_n5690_ = new_n5688_;
  assign new_n5691_ = new_n5687_;
  assign new_n5692_ = new_n3508_;
  assign new_n5693_ = new_n3564_;
  assign new_n5694_ = new_n2438_;
  assign new_n5695_ = new_n5694_;
  assign new_n5696_ = new_n5694_;
  assign new_n5697_ = new_n2404_;
  assign new_n5698_ = new_n5697_;
  assign new_n5699_ = new_n5697_;
  assign new_n5700_ = new_n4001_;
  assign new_n5701_ = new_n5700_;
  assign new_n5702_ = new_n5701_;
  assign new_n5703_ = new_n5700_;
  assign new_n5704_ = new_n2353_;
  assign new_n5705_ = new_n5704_;
  assign new_n5706_ = new_n5705_;
  assign new_n5707_ = new_n5705_;
  assign new_n5708_ = new_n5704_;
  assign new_n5709_ = new_n5708_;
  assign new_n5710_ = new_n5708_;
  assign new_n5711_ = new_n2368_;
  assign new_n5712_ = new_n5711_;
  assign new_n5713_ = new_n5712_;
  assign new_n5714_ = new_n5713_;
  assign new_n5715_ = new_n5713_;
  assign new_n5716_ = new_n5712_;
  assign new_n5717_ = new_n5716_;
  assign new_n5718_ = new_n5716_;
  assign new_n5719_ = new_n5711_;
  assign new_n5720_ = new_n5719_;
  assign new_n5721_ = new_n5719_;
  assign new_n5722_ = new_n2369_;
  assign new_n5723_ = new_n5722_;
  assign new_n5724_ = new_n5723_;
  assign new_n5725_ = new_n5723_;
  assign new_n5726_ = new_n5722_;
  assign new_n5727_ = new_n5726_;
  assign new_n5728_ = new_n5726_;
  assign new_n5729_ = new_n2352_;
  assign new_n5730_ = new_n5729_;
  assign new_n5731_ = new_n5730_;
  assign new_n5732_ = new_n5731_;
  assign new_n5733_ = new_n5731_;
  assign new_n5734_ = new_n5730_;
  assign new_n5735_ = new_n5734_;
  assign new_n5736_ = new_n5734_;
  assign new_n5737_ = new_n5729_;
  assign new_n5738_ = new_n5737_;
  assign new_n5739_ = new_n5737_;
  assign new_n5740_ = new_n2401_;
  assign new_n5741_ = new_n2447_;
  assign new_n5742_ = new_n5741_;
  assign new_n5743_ = new_n3259_;
  assign new_n5744_ = new_n3273_;
  assign new_n5745_ = new_n3276_;
  assign new_n5746_ = new_n3282_;
  assign new_n5747_ = new_n3396_;
  assign new_n5748_ = new_n3430_;
  assign new_n5749_ = new_n3443_;
  assign new_n5750_ = new_n2472_;
  assign new_n5751_ = new_n5750_;
  assign new_n5752_ = new_n2480_;
  assign new_n5753_ = new_n5752_;
  assign new_n5754_ = new_n2808_;
  assign new_n5755_ = new_n5754_;
  assign new_n5756_ = new_n2414_;
  assign new_n5757_ = new_n2434_;
  assign new_n5758_ = new_n2456_;
  assign new_n5759_ = new_n2430_;
  assign new_n5760_ = new_n3531_;
  assign new_n5761_ = new_n5760_;
  assign new_n5762_ = new_n5761_;
  assign new_n5763_ = new_n5760_;
  assign new_n5764_ = new_n3764_;
  assign new_n5765_ = new_n3767_;
  assign new_n5766_ = new_n3794_;
  assign new_n5767_ = new_n3809_;
  assign new_n5768_ = new_n3812_;
  assign new_n5769_ = new_n3841_;
  assign new_n5770_ = new_n3870_;
  assign new_n5771_ = new_n3899_;
  assign new_n5772_ = new_n3977_;
  assign new_n5773_ = new_n5772_;
  assign new_n5774_ = new_n3979_;
  assign new_n5775_ = new_n5774_;
  assign new_n5776_ = new_n3990_;
  assign new_n5777_ = new_n5776_;
  assign new_n5778_ = new_n4012_;
  assign new_n5779_ = new_n5778_;
  assign new_n5780_ = new_n4014_;
  assign new_n5781_ = new_n5780_;
  assign new_n5782_ = new_n5781_;
  assign new_n5783_ = new_n5781_;
  assign new_n5784_ = new_n5780_;
  assign new_n5785_ = new_n2510_;
  assign new_n5786_ = new_n2514_;
  assign new_n5787_ = new_n4154_;
  assign new_n5788_ = new_n5787_;
  assign new_n5789_ = new_n5788_;
  assign new_n5790_ = new_n5787_;
  always @ (posedge clock) begin
    n1416_lo <= n1416_li;
    n1419_lo <= n1419_li;
    n1422_lo <= n1422_li;
    n1425_lo <= n1425_li;
    n1428_lo <= n1428_li;
    n1431_lo <= n1431_li;
    n1434_lo <= n1434_li;
    n1437_lo <= n1437_li;
    n1440_lo <= n1440_li;
    n1443_lo <= n1443_li;
    n1446_lo <= n1446_li;
    n1449_lo <= n1449_li;
    n1452_lo <= n1452_li;
    n1455_lo <= n1455_li;
    n1458_lo <= n1458_li;
    n1464_lo <= n1464_li;
    n1467_lo <= n1467_li;
    n1470_lo <= n1470_li;
    n1476_lo <= n1476_li;
    n1479_lo <= n1479_li;
    n1482_lo <= n1482_li;
    n1488_lo <= n1488_li;
    n1491_lo <= n1491_li;
    n1494_lo <= n1494_li;
    n1497_lo <= n1497_li;
    n1500_lo <= n1500_li;
    n1512_lo <= n1512_li;
    n1515_lo <= n1515_li;
    n1518_lo <= n1518_li;
    n1521_lo <= n1521_li;
    n1524_lo <= n1524_li;
    n1527_lo <= n1527_li;
    n1530_lo <= n1530_li;
    n1533_lo <= n1533_li;
    n1536_lo <= n1536_li;
    n1539_lo <= n1539_li;
    n1542_lo <= n1542_li;
    n1545_lo <= n1545_li;
    n1548_lo <= n1548_li;
    n1551_lo <= n1551_li;
    n1554_lo <= n1554_li;
    n1560_lo <= n1560_li;
    n1563_lo <= n1563_li;
    n1566_lo <= n1566_li;
    n1572_lo <= n1572_li;
    n1575_lo <= n1575_li;
    n1578_lo <= n1578_li;
    n1584_lo <= n1584_li;
    n1587_lo <= n1587_li;
    n1590_lo <= n1590_li;
    n1596_lo <= n1596_li;
    n1599_lo <= n1599_li;
    n1602_lo <= n1602_li;
    n1608_lo <= n1608_li;
    n1611_lo <= n1611_li;
    n1614_lo <= n1614_li;
    n1620_lo <= n1620_li;
    n1623_lo <= n1623_li;
    n1626_lo <= n1626_li;
    n1632_lo <= n1632_li;
    n1635_lo <= n1635_li;
    n1638_lo <= n1638_li;
    n1644_lo <= n1644_li;
    n1647_lo <= n1647_li;
    n1650_lo <= n1650_li;
    n1656_lo <= n1656_li;
    n1659_lo <= n1659_li;
    n1662_lo <= n1662_li;
    n1668_lo <= n1668_li;
    n1671_lo <= n1671_li;
    n1674_lo <= n1674_li;
    n1677_lo <= n1677_li;
    n1680_lo <= n1680_li;
    n1683_lo <= n1683_li;
    n1686_lo <= n1686_li;
    n1692_lo <= n1692_li;
    n1695_lo <= n1695_li;
    n1698_lo <= n1698_li;
    n1704_lo <= n1704_li;
    n1707_lo <= n1707_li;
    n1710_lo <= n1710_li;
    n1716_lo <= n1716_li;
    n1719_lo <= n1719_li;
    n1722_lo <= n1722_li;
    n1728_lo <= n1728_li;
    n1731_lo <= n1731_li;
    n1734_lo <= n1734_li;
    n1740_lo <= n1740_li;
    n1743_lo <= n1743_li;
    n1746_lo <= n1746_li;
    n1749_lo <= n1749_li;
    n1752_lo <= n1752_li;
    n1755_lo <= n1755_li;
    n1758_lo <= n1758_li;
    n1761_lo <= n1761_li;
    n1764_lo <= n1764_li;
    n1776_lo <= n1776_li;
    n1779_lo <= n1779_li;
    n1788_lo <= n1788_li;
    n1791_lo <= n1791_li;
    n1794_lo <= n1794_li;
    n1797_lo <= n1797_li;
    n1800_lo <= n1800_li;
    n1812_lo <= n1812_li;
    n1824_lo <= n1824_li;
    n1836_lo <= n1836_li;
    n1848_lo <= n1848_li;
    n1860_lo <= n1860_li;
    n1872_lo <= n1872_li;
    n1884_lo <= n1884_li;
    n1896_lo <= n1896_li;
    n1899_lo <= n1899_li;
    n1908_lo <= n1908_li;
    n1911_lo <= n1911_li;
    n1920_lo <= n1920_li;
    n1923_lo <= n1923_li;
    n1926_lo <= n1926_li;
    n1929_lo <= n1929_li;
    n1932_lo <= n1932_li;
    n1944_lo <= n1944_li;
    n1956_lo <= n1956_li;
    n1968_lo <= n1968_li;
    n1980_lo <= n1980_li;
    n1992_lo <= n1992_li;
    n2004_lo <= n2004_li;
    n2016_lo <= n2016_li;
    n2019_lo <= n2019_li;
    n2028_lo <= n2028_li;
    n2031_lo <= n2031_li;
    n2040_lo <= n2040_li;
    n2043_lo <= n2043_li;
    n2046_lo <= n2046_li;
    n2049_lo <= n2049_li;
    n2052_lo <= n2052_li;
    n2064_lo <= n2064_li;
    n2076_lo <= n2076_li;
    n2088_lo <= n2088_li;
    n2100_lo <= n2100_li;
    n2112_lo <= n2112_li;
    n2124_lo <= n2124_li;
    n2136_lo <= n2136_li;
    n2148_lo <= n2148_li;
    n2151_lo <= n2151_li;
    n2160_lo <= n2160_li;
    n2163_lo <= n2163_li;
    n2172_lo <= n2172_li;
    n2175_lo <= n2175_li;
    n2178_lo <= n2178_li;
    n2181_lo <= n2181_li;
    n2184_lo <= n2184_li;
    n2196_lo <= n2196_li;
    n2208_lo <= n2208_li;
    n2220_lo <= n2220_li;
    n2232_lo <= n2232_li;
    n2244_lo <= n2244_li;
    n2256_lo <= n2256_li;
    n2268_lo <= n2268_li;
    n2280_lo <= n2280_li;
    n2283_lo <= n2283_li;
    n2292_lo <= n2292_li;
    n2295_lo <= n2295_li;
    n2298_lo <= n2298_li;
    n2301_lo <= n2301_li;
    n2304_lo <= n2304_li;
    n2316_lo <= n2316_li;
    n2319_lo <= n2319_li;
    n2322_lo <= n2322_li;
    n2325_lo <= n2325_li;
    n2328_lo <= n2328_li;
    n2331_lo <= n2331_li;
    n2340_lo <= n2340_li;
    n2343_lo <= n2343_li;
    n2376_lo <= n2376_li;
    n2379_lo <= n2379_li;
    n2388_lo <= n2388_li;
    n2400_lo <= n2400_li;
    n2412_lo <= n2412_li;
    n2415_lo <= n2415_li;
    n2424_lo <= n2424_li;
    n2436_lo <= n2436_li;
    n2439_lo <= n2439_li;
    n2442_lo <= n2442_li;
    n2445_lo <= n2445_li;
    n2448_lo <= n2448_li;
    n2451_lo <= n2451_li;
    n2460_lo <= n2460_li;
    n2463_lo <= n2463_li;
    n2496_lo <= n2496_li;
    n2499_lo <= n2499_li;
    n2508_lo <= n2508_li;
    n2520_lo <= n2520_li;
    n2532_lo <= n2532_li;
    n2535_lo <= n2535_li;
    n2544_lo <= n2544_li;
    n2556_lo <= n2556_li;
    n2559_lo <= n2559_li;
    n2562_lo <= n2562_li;
    n2565_lo <= n2565_li;
    n2568_lo <= n2568_li;
    n2571_lo <= n2571_li;
    n2580_lo <= n2580_li;
    n2583_lo <= n2583_li;
    n2616_lo <= n2616_li;
    n2619_lo <= n2619_li;
    n2628_lo <= n2628_li;
    n2640_lo <= n2640_li;
    n2652_lo <= n2652_li;
    n2655_lo <= n2655_li;
    n2664_lo <= n2664_li;
    n2676_lo <= n2676_li;
    n2679_lo <= n2679_li;
    n2682_lo <= n2682_li;
    n2685_lo <= n2685_li;
    n2688_lo <= n2688_li;
    n2691_lo <= n2691_li;
    n2700_lo <= n2700_li;
    n2703_lo <= n2703_li;
    n2736_lo <= n2736_li;
    n2739_lo <= n2739_li;
    n2748_lo <= n2748_li;
    n2760_lo <= n2760_li;
    n2772_lo <= n2772_li;
    n2775_lo <= n2775_li;
    n2784_lo <= n2784_li;
    n2787_lo <= n2787_li;
    n2790_lo <= n2790_li;
    n2793_lo <= n2793_li;
    n2796_lo <= n2796_li;
    n2799_lo <= n2799_li;
    n2802_lo <= n2802_li;
    n2805_lo <= n2805_li;
    n2808_lo <= n2808_li;
    n2820_lo <= n2820_li;
    n2823_lo <= n2823_li;
    n2826_lo <= n2826_li;
    n2832_lo <= n2832_li;
    n2835_lo <= n2835_li;
    n2838_lo <= n2838_li;
    n2841_lo <= n2841_li;
    n2844_lo <= n2844_li;
    n2856_lo <= n2856_li;
    n2859_lo <= n2859_li;
    n2862_lo <= n2862_li;
    n2865_lo <= n2865_li;
    n2868_lo <= n2868_li;
    n2871_lo <= n2871_li;
    n2874_lo <= n2874_li;
    n2877_lo <= n2877_li;
    n2880_lo <= n2880_li;
    n2883_lo <= n2883_li;
    n2886_lo <= n2886_li;
    n2889_lo <= n2889_li;
    n2892_lo <= n2892_li;
    n2895_lo <= n2895_li;
    n2898_lo <= n2898_li;
    n2901_lo <= n2901_li;
    n2904_lo <= n2904_li;
    n2907_lo <= n2907_li;
    n2916_lo <= n2916_li;
    n2928_lo <= n2928_li;
    n2940_lo <= n2940_li;
    n2952_lo <= n2952_li;
    n2955_lo <= n2955_li;
    n2964_lo <= n2964_li;
    n2976_lo <= n2976_li;
    n2988_lo <= n2988_li;
    n2991_lo <= n2991_li;
    n3000_lo <= n3000_li;
    n3003_lo <= n3003_li;
    n3012_lo <= n3012_li;
    n3015_lo <= n3015_li;
    n3024_lo <= n3024_li;
    n3027_lo <= n3027_li;
    n3036_lo <= n3036_li;
    n3039_lo <= n3039_li;
    n3048_lo <= n3048_li;
    n3051_lo <= n3051_li;
    n3054_lo <= n3054_li;
    n3057_lo <= n3057_li;
    n3060_lo <= n3060_li;
    n3072_lo <= n3072_li;
    n3081_lo <= n3081_li;
    n3084_lo <= n3084_li;
    n3087_lo <= n3087_li;
    n3093_lo <= n3093_li;
    n3096_lo <= n3096_li;
    n3105_lo <= n3105_li;
    n3108_lo <= n3108_li;
    n3117_lo <= n3117_li;
    n3120_lo <= n3120_li;
    n3123_lo <= n3123_li;
    n3126_lo <= n3126_li;
    n3129_lo <= n3129_li;
    n3132_lo <= n3132_li;
    n3135_lo <= n3135_li;
    n3138_lo <= n3138_li;
    n3141_lo <= n3141_li;
    n3168_lo <= n3168_li;
    n3171_lo <= n3171_li;
    n3174_lo <= n3174_li;
    n3177_lo <= n3177_li;
    n3180_lo <= n3180_li;
    n3183_lo <= n3183_li;
    n3192_lo <= n3192_li;
    n3195_lo <= n3195_li;
    n3204_lo <= n3204_li;
    n3207_lo <= n3207_li;
    n3216_lo <= n3216_li;
    n3219_lo <= n3219_li;
    n3228_lo <= n3228_li;
    n3231_lo <= n3231_li;
    n3240_lo <= n3240_li;
    n3243_lo <= n3243_li;
    n3252_lo <= n3252_li;
    n3255_lo <= n3255_li;
    n3258_lo <= n3258_li;
    n3264_lo <= n3264_li;
    n3267_lo <= n3267_li;
    n3270_lo <= n3270_li;
    n3276_lo <= n3276_li;
    n3279_lo <= n3279_li;
    n3282_lo <= n3282_li;
    n3288_lo <= n3288_li;
    n3291_lo <= n3291_li;
    n3294_lo <= n3294_li;
    n4537_o2 <= n4537_i2;
    n4538_o2 <= n4538_i2;
    n4710_o2 <= n4710_i2;
    n4711_o2 <= n4711_i2;
    n1211_inv <= n4803_i2;
    n1214_inv <= n4804_i2;
    n1217_inv <= n4843_i2;
    n1220_inv <= n4844_i2;
    n4927_o2 <= n4927_i2;
    n4928_o2 <= n4928_i2;
    n1229_inv <= n4945_i2;
    n1232_inv <= n4946_i2;
    n1235_inv <= n5009_i2;
    n5178_o2 <= n5178_i2;
    n5179_o2 <= n5179_i2;
    n5477_o2 <= n5477_i2;
    n5478_o2 <= n5478_i2;
    n5479_o2 <= n5479_i2;
    n5222_o2 <= n5222_i2;
    n5223_o2 <= n5223_i2;
    n5553_o2 <= n5553_i2;
    n5554_o2 <= n5554_i2;
    G491_o2 <= G491_i2;
    n2922_lo_buf_o2 <= n2922_lo_buf_i2;
    n2946_lo_buf_o2 <= n2946_lo_buf_i2;
    n2970_lo_buf_o2 <= n2970_lo_buf_i2;
    n2982_lo_buf_o2 <= n2982_lo_buf_i2;
    n3066_lo_buf_o2 <= n3066_lo_buf_i2;
    n3078_lo_buf_o2 <= n3078_lo_buf_i2;
    n3102_lo_buf_o2 <= n3102_lo_buf_i2;
    n3114_lo_buf_o2 <= n3114_lo_buf_i2;
    G1321_o2 <= G1321_i2;
    G1033_o2 <= G1033_i2;
    G1030_o2 <= G1030_i2;
    G1072_o2 <= G1072_i2;
    n1304_inv <= G1159_i2;
    n1307_inv <= G1152_i2;
    n2958_lo_buf_o2 <= n2958_lo_buf_i2;
    n2994_lo_buf_o2 <= n2994_lo_buf_i2;
    n3006_lo_buf_o2 <= n3006_lo_buf_i2;
    n3030_lo_buf_o2 <= n3030_lo_buf_i2;
    n3042_lo_buf_o2 <= n3042_lo_buf_i2;
    n3090_lo_buf_o2 <= n3090_lo_buf_i2;
    n1328_inv <= G370_i2;
    n1331_inv <= G447_i2;
    n1334_inv <= G455_i2;
    n1337_inv <= G459_i2;
    n1340_inv <= G497_i2;
    n1343_inv <= G503_i2;
    n1346_inv <= G511_i2;
    n1349_inv <= G515_i2;
    G1036_o2 <= G1036_i2;
    G1062_o2 <= G1062_i2;
    G1067_o2 <= G1067_i2;
    G1014_o2 <= G1014_i2;
    n1364_inv <= G1171_i2;
    n1367_inv <= G1166_i2;
    n3018_lo_buf_o2 <= n3018_lo_buf_i2;
    G766_o2 <= G766_i2;
    n1376_inv <= G451_i2;
    n1379_inv <= G463_i2;
    n1382_inv <= G467_i2;
    n1385_inv <= G475_i2;
    n1388_inv <= G479_i2;
    n1391_inv <= G507_i2;
    G1017_o2 <= G1017_i2;
    G1008_o2 <= G1008_i2;
    n1400_inv <= G1176_i2;
    n1403_inv <= G1144_i2;
    n2910_lo_buf_o2 <= n2910_lo_buf_i2;
    n1409_inv <= G471_i2;
    G2138_o2 <= G2138_i2;
    G2147_o2 <= G2147_i2;
    n1418_inv <= G1148_i2;
    G1137_o2 <= G1137_i2;
    G1329_o2 <= G1329_i2;
    G374_o2 <= G374_i2;
    G386_o2 <= G386_i2;
    G663_o2 <= G663_i2;
    G674_o2 <= G674_i2;
    G578_o2 <= G578_i2;
    G575_o2 <= G575_i2;
    G2505_o2 <= G2505_i2;
    n1448_inv <= G2508_i2;
    G987_o2 <= G987_i2;
    G984_o2 <= G984_i2;
    G1862_o2 <= G1862_i2;
    G1859_o2 <= G1859_i2;
    G1260_o2 <= G1260_i2;
    G1865_o2 <= G1865_i2;
    G2073_o2 <= G2073_i2;
    G1402_o2 <= G1402_i2;
    G2048_o2 <= G2048_i2;
    G2276_o2 <= G2276_i2;
    n1481_inv <= G366_i2;
    G2141_o2 <= G2141_i2;
    G2008_o2 <= G2008_i2;
    G2011_o2 <= G2011_i2;
    G2150_o2 <= G2150_i2;
    G2026_o2 <= G2026_i2;
    G2029_o2 <= G2029_i2;
    G2023_o2 <= G2023_i2;
    G2041_o2 <= G2041_i2;
    G2017_o2 <= G2017_i2;
    G2020_o2 <= G2020_i2;
    G2035_o2 <= G2035_i2;
    G2038_o2 <= G2038_i2;
    G2228_o2 <= G2228_i2;
    G2231_o2 <= G2231_i2;
    G2234_o2 <= G2234_i2;
    G2237_o2 <= G2237_i2;
    G1904_o2 <= G1904_i2;
    G1907_o2 <= G1907_i2;
    G1928_o2 <= G1928_i2;
    G1931_o2 <= G1931_i2;
    G1893_o2 <= G1893_i2;
    G1896_o2 <= G1896_i2;
    G1899_o2 <= G1899_i2;
    G1937_o2 <= G1937_i2;
    G1940_o2 <= G1940_i2;
    G1943_o2 <= G1943_i2;
    G1336_o2 <= G1336_i2;
    G1996_o2 <= G1996_i2;
    G1999_o2 <= G1999_i2;
    G2002_o2 <= G2002_i2;
    G2005_o2 <= G2005_i2;
    G2014_o2 <= G2014_i2;
    G2032_o2 <= G2032_i2;
    G1076_o2 <= G1076_i2;
    G1002_o2 <= G1002_i2;
    G998_o2 <= G998_i2;
    G1890_o2 <= G1890_i2;
    G1934_o2 <= G1934_i2;
    G1044_o2 <= G1044_i2;
    G1039_o2 <= G1039_i2;
    n1770_lo_buf_o2 <= n1770_lo_buf_i2;
    G342_o2 <= G342_i2;
    G354_o2 <= G354_i2;
    G1193_o2 <= G1193_i2;
    n3234_lo_buf_o2 <= n3234_lo_buf_i2;
    n3246_lo_buf_o2 <= n3246_lo_buf_i2;
    G783_o2 <= G783_i2;
    G786_o2 <= G786_i2;
    G792_o2 <= G792_i2;
    G795_o2 <= G795_i2;
    G815_o2 <= G815_i2;
    G818_o2 <= G818_i2;
    G824_o2 <= G824_i2;
    G827_o2 <= G827_i2;
    G789_o2 <= G789_i2;
    G798_o2 <= G798_i2;
    G801_o2 <= G801_i2;
    G807_o2 <= G807_i2;
    G812_o2 <= G812_i2;
    G821_o2 <= G821_i2;
    G804_o2 <= G804_i2;
    G780_o2 <= G780_i2;
    G1231_o2 <= G1231_i2;
    G1572_o2 <= G1572_i2;
    G1377_o2 <= G1377_i2;
    G1253_o2 <= G1253_i2;
    G1359_o2 <= G1359_i2;
    G1258_o2 <= G1258_i2;
    G1367_o2 <= G1367_i2;
    G1358_o2 <= G1358_i2;
    G1366_o2 <= G1366_i2;
    G2057_o2 <= G2057_i2;
    G2117_o2 <= G2117_i2;
    G2118_o2 <= G2118_i2;
    G1254_o2 <= G1254_i2;
    G1259_o2 <= G1259_i2;
    G2058_o2 <= G2058_i2;
    G405_o2 <= G405_i2;
    G417_o2 <= G417_i2;
    G1269_o2 <= G1269_i2;
    G1275_o2 <= G1275_i2;
    G1287_o2 <= G1287_i2;
    G1266_o2 <= G1266_i2;
    G1272_o2 <= G1272_i2;
    G1278_o2 <= G1278_i2;
    G1281_o2 <= G1281_i2;
    G1284_o2 <= G1284_i2;
    G1290_o2 <= G1290_i2;
    G1293_o2 <= G1293_i2;
    G1299_o2 <= G1299_i2;
    G1305_o2 <= G1305_i2;
    G1296_o2 <= G1296_i2;
    G1302_o2 <= G1302_i2;
    G1308_o2 <= G1308_i2;
    G1311_o2 <= G1311_i2;
    G811_o2 <= G811_i2;
    G810_o2 <= G810_i2;
    G1728_o2 <= G1728_i2;
    G2512_o2 <= G2512_i2;
    G1114_o2 <= G1114_i2;
    G1113_o2 <= G1113_i2;
    G1992_o2 <= G1992_i2;
    G1991_o2 <= G1991_i2;
    G1426_o2 <= G1426_i2;
    G1966_o2 <= G1966_i2;
    G2211_o2 <= G2211_i2;
    G1509_o2 <= G1509_i2;
    G2153_o2 <= G2153_i2;
    G2329_o2 <= G2329_i2;
    G1540_o2 <= G1540_i2;
    G2167_o2 <= G2167_i2;
    G2191_o2 <= G2191_i2;
    G1234_o2 <= G1234_i2;
    G1132_o2 <= G1132_i2;
    G1129_o2 <= G1129_i2;
    G2088_o2 <= G2088_i2;
    G2106_o2 <= G2106_i2;
    G1314_o2 <= G1314_i2;
    G636_o2 <= G636_i2;
    G647_o2 <= G647_i2;
    n3186_lo_buf_o2 <= n3186_lo_buf_i2;
    n3198_lo_buf_o2 <= n3198_lo_buf_i2;
    n3210_lo_buf_o2 <= n3210_lo_buf_i2;
    n3222_lo_buf_o2 <= n3222_lo_buf_i2;
    G1225_o2 <= G1225_i2;
    G1342_o2 <= G1342_i2;
    G1222_o2 <= G1222_i2;
    G1228_o2 <= G1228_i2;
    G1348_o2 <= G1348_i2;
    G1345_o2 <= G1345_i2;
    G1351_o2 <= G1351_i2;
    G2242_o2 <= G2242_i2;
    G2260_o2 <= G2260_i2;
    G1374_o2 <= G1374_i2;
    G1537_o2 <= G1537_i2;
    G301_o2 <= G301_i2;
    G313_o2 <= G313_i2;
    G2365_o2 <= G2365_i2;
    G2255_o2 <= G2255_i2;
    G2253_o2 <= G2253_i2;
    G2395_o2 <= G2395_i2;
    G2272_o2 <= G2272_i2;
    G2270_o2 <= G2270_i2;
    G2245_o2 <= G2245_i2;
    G2262_o2 <= G2262_i2;
    G2249_o2 <= G2249_i2;
    G2247_o2 <= G2247_i2;
    G2266_o2 <= G2266_i2;
    G2264_o2 <= G2264_i2;
    G2403_o2 <= G2403_i2;
    G2401_o2 <= G2401_i2;
    G2410_o2 <= G2410_i2;
    G2408_o2 <= G2408_i2;
    G2306_o2 <= G2306_i2;
    G2305_o2 <= G2305_i2;
    G2314_o2 <= G2314_i2;
    G2313_o2 <= G2313_i2;
    G2303_o2 <= G2303_i2;
    G2302_o2 <= G2302_i2;
    G2301_o2 <= G2301_i2;
    G2311_o2 <= G2311_i2;
    G2310_o2 <= G2310_i2;
    G2309_o2 <= G2309_i2;
    G2404_o2 <= G2404_i2;
    G2411_o2 <= G2411_i2;
    G2420_o2 <= G2420_i2;
    G2419_o2 <= G2419_i2;
    G2433_o2 <= G2433_i2;
    G2432_o2 <= G2432_i2;
    G402_o2 <= G402_i2;
    G403_o2 <= G403_i2;
    G1053_o2 <= G1053_i2;
    G1049_o2 <= G1049_i2;
    n2003_inv <= G1058_i2;
    G1364_o2 <= G1364_i2;
    G1079_o2 <= G1079_i2;
    G1478_o2 <= G1478_i2;
    G707_o2 <= G707_i2;
    G718_o2 <= G718_i2;
    G2417_o2 <= G2417_i2;
    G2414_o2 <= G2414_i2;
    G2431_o2 <= G2431_i2;
    G2428_o2 <= G2428_i2;
    G1653_o2 <= G1653_i2;
    G2213_o2 <= G2213_i2;
    G2221_o2 <= G2221_i2;
    G2250_o2 <= G2250_i2;
    G2267_o2 <= G2267_i2;
    G1365_o2 <= G1365_i2;
    G1368_o2 <= G1368_i2;
    G1371_o2 <= G1371_i2;
    G2218_o2 <= G2218_i2;
    G2225_o2 <= G2225_i2;
    n1503_lo_buf_o2 <= n1503_lo_buf_i2;
    n1863_lo_buf_o2 <= n1863_lo_buf_i2;
    n1887_lo_buf_o2 <= n1887_lo_buf_i2;
    n1983_lo_buf_o2 <= n1983_lo_buf_i2;
    n2007_lo_buf_o2 <= n2007_lo_buf_i2;
    n2115_lo_buf_o2 <= n2115_lo_buf_i2;
    n2139_lo_buf_o2 <= n2139_lo_buf_i2;
    n2247_lo_buf_o2 <= n2247_lo_buf_i2;
    n2271_lo_buf_o2 <= n2271_lo_buf_i2;
    n2919_lo_buf_o2 <= n2919_lo_buf_i2;
    n2943_lo_buf_o2 <= n2943_lo_buf_i2;
    n2967_lo_buf_o2 <= n2967_lo_buf_i2;
    n2979_lo_buf_o2 <= n2979_lo_buf_i2;
    n3063_lo_buf_o2 <= n3063_lo_buf_i2;
    n3075_lo_buf_o2 <= n3075_lo_buf_i2;
    n3099_lo_buf_o2 <= n3099_lo_buf_i2;
    n3111_lo_buf_o2 <= n3111_lo_buf_i2;
    G878_o2 <= G878_i2;
    G875_o2 <= G875_i2;
    G661_o2 <= G661_i2;
    G660_o2 <= G660_i2;
    G879_o2 <= G879_i2;
    G876_o2 <= G876_i2;
    G1320_o2 <= G1320_i2;
    G941_o2 <= G941_i2;
    G732_o2 <= G732_i2;
    G942_o2 <= G942_i2;
    G1493_o2 <= G1493_i2;
    G1498_o2 <= G1498_i2;
    G877_o2 <= G877_i2;
    G874_o2 <= G874_i2;
    n1806_lo_buf_o2 <= n1806_lo_buf_i2;
    n1878_lo_buf_o2 <= n1878_lo_buf_i2;
    n1938_lo_buf_o2 <= n1938_lo_buf_i2;
    n1998_lo_buf_o2 <= n1998_lo_buf_i2;
    n2058_lo_buf_o2 <= n2058_lo_buf_i2;
    n2130_lo_buf_o2 <= n2130_lo_buf_i2;
    n2190_lo_buf_o2 <= n2190_lo_buf_i2;
    n2262_lo_buf_o2 <= n2262_lo_buf_i2;
    n2310_lo_buf_o2 <= n2310_lo_buf_i2;
    n2406_lo_buf_o2 <= n2406_lo_buf_i2;
    n2430_lo_buf_o2 <= n2430_lo_buf_i2;
    n2526_lo_buf_o2 <= n2526_lo_buf_i2;
    n2550_lo_buf_o2 <= n2550_lo_buf_i2;
    n2646_lo_buf_o2 <= n2646_lo_buf_i2;
    n2670_lo_buf_o2 <= n2670_lo_buf_i2;
    n2766_lo_buf_o2 <= n2766_lo_buf_i2;
    G603_o2 <= G603_i2;
    G614_o2 <= G614_i2;
    G1026_o2 <= G1026_i2;
    G1021_o2 <= G1021_i2;
    G940_o2 <= G940_i2;
    G1636_o2 <= G1636_i2;
    G1684_o2 <= G1684_i2;
    n2352_lo_buf_o2 <= n2352_lo_buf_i2;
    n2364_lo_buf_o2 <= n2364_lo_buf_i2;
    n2472_lo_buf_o2 <= n2472_lo_buf_i2;
    n2484_lo_buf_o2 <= n2484_lo_buf_i2;
    n2592_lo_buf_o2 <= n2592_lo_buf_i2;
    n2604_lo_buf_o2 <= n2604_lo_buf_i2;
    n2712_lo_buf_o2 <= n2712_lo_buf_i2;
    n2724_lo_buf_o2 <= n2724_lo_buf_i2;
    n3150_lo_buf_o2 <= n3150_lo_buf_i2;
    n3162_lo_buf_o2 <= n3162_lo_buf_i2;
  end
  initial begin
    n1416_lo <= 1'b0;
    n1419_lo <= 1'b0;
    n1422_lo <= 1'b0;
    n1425_lo <= 1'b0;
    n1428_lo <= 1'b0;
    n1431_lo <= 1'b0;
    n1434_lo <= 1'b0;
    n1437_lo <= 1'b0;
    n1440_lo <= 1'b0;
    n1443_lo <= 1'b0;
    n1446_lo <= 1'b0;
    n1449_lo <= 1'b0;
    n1452_lo <= 1'b0;
    n1455_lo <= 1'b0;
    n1458_lo <= 1'b0;
    n1464_lo <= 1'b0;
    n1467_lo <= 1'b0;
    n1470_lo <= 1'b0;
    n1476_lo <= 1'b0;
    n1479_lo <= 1'b0;
    n1482_lo <= 1'b0;
    n1488_lo <= 1'b0;
    n1491_lo <= 1'b0;
    n1494_lo <= 1'b0;
    n1497_lo <= 1'b0;
    n1500_lo <= 1'b0;
    n1512_lo <= 1'b0;
    n1515_lo <= 1'b0;
    n1518_lo <= 1'b0;
    n1521_lo <= 1'b0;
    n1524_lo <= 1'b0;
    n1527_lo <= 1'b0;
    n1530_lo <= 1'b0;
    n1533_lo <= 1'b0;
    n1536_lo <= 1'b0;
    n1539_lo <= 1'b0;
    n1542_lo <= 1'b0;
    n1545_lo <= 1'b0;
    n1548_lo <= 1'b0;
    n1551_lo <= 1'b0;
    n1554_lo <= 1'b0;
    n1560_lo <= 1'b0;
    n1563_lo <= 1'b0;
    n1566_lo <= 1'b0;
    n1572_lo <= 1'b0;
    n1575_lo <= 1'b0;
    n1578_lo <= 1'b0;
    n1584_lo <= 1'b0;
    n1587_lo <= 1'b0;
    n1590_lo <= 1'b0;
    n1596_lo <= 1'b0;
    n1599_lo <= 1'b0;
    n1602_lo <= 1'b0;
    n1608_lo <= 1'b0;
    n1611_lo <= 1'b0;
    n1614_lo <= 1'b0;
    n1620_lo <= 1'b0;
    n1623_lo <= 1'b0;
    n1626_lo <= 1'b0;
    n1632_lo <= 1'b0;
    n1635_lo <= 1'b0;
    n1638_lo <= 1'b0;
    n1644_lo <= 1'b0;
    n1647_lo <= 1'b0;
    n1650_lo <= 1'b0;
    n1656_lo <= 1'b0;
    n1659_lo <= 1'b0;
    n1662_lo <= 1'b0;
    n1668_lo <= 1'b0;
    n1671_lo <= 1'b0;
    n1674_lo <= 1'b0;
    n1677_lo <= 1'b0;
    n1680_lo <= 1'b0;
    n1683_lo <= 1'b0;
    n1686_lo <= 1'b0;
    n1692_lo <= 1'b0;
    n1695_lo <= 1'b0;
    n1698_lo <= 1'b0;
    n1704_lo <= 1'b0;
    n1707_lo <= 1'b0;
    n1710_lo <= 1'b0;
    n1716_lo <= 1'b0;
    n1719_lo <= 1'b0;
    n1722_lo <= 1'b0;
    n1728_lo <= 1'b0;
    n1731_lo <= 1'b0;
    n1734_lo <= 1'b0;
    n1740_lo <= 1'b0;
    n1743_lo <= 1'b0;
    n1746_lo <= 1'b0;
    n1749_lo <= 1'b0;
    n1752_lo <= 1'b0;
    n1755_lo <= 1'b0;
    n1758_lo <= 1'b0;
    n1761_lo <= 1'b0;
    n1764_lo <= 1'b0;
    n1776_lo <= 1'b0;
    n1779_lo <= 1'b0;
    n1788_lo <= 1'b0;
    n1791_lo <= 1'b0;
    n1794_lo <= 1'b0;
    n1797_lo <= 1'b0;
    n1800_lo <= 1'b0;
    n1812_lo <= 1'b0;
    n1824_lo <= 1'b0;
    n1836_lo <= 1'b0;
    n1848_lo <= 1'b0;
    n1860_lo <= 1'b0;
    n1872_lo <= 1'b0;
    n1884_lo <= 1'b0;
    n1896_lo <= 1'b0;
    n1899_lo <= 1'b0;
    n1908_lo <= 1'b0;
    n1911_lo <= 1'b0;
    n1920_lo <= 1'b0;
    n1923_lo <= 1'b0;
    n1926_lo <= 1'b0;
    n1929_lo <= 1'b0;
    n1932_lo <= 1'b0;
    n1944_lo <= 1'b0;
    n1956_lo <= 1'b0;
    n1968_lo <= 1'b0;
    n1980_lo <= 1'b0;
    n1992_lo <= 1'b0;
    n2004_lo <= 1'b0;
    n2016_lo <= 1'b0;
    n2019_lo <= 1'b0;
    n2028_lo <= 1'b0;
    n2031_lo <= 1'b0;
    n2040_lo <= 1'b0;
    n2043_lo <= 1'b0;
    n2046_lo <= 1'b0;
    n2049_lo <= 1'b0;
    n2052_lo <= 1'b0;
    n2064_lo <= 1'b0;
    n2076_lo <= 1'b0;
    n2088_lo <= 1'b0;
    n2100_lo <= 1'b0;
    n2112_lo <= 1'b0;
    n2124_lo <= 1'b0;
    n2136_lo <= 1'b0;
    n2148_lo <= 1'b0;
    n2151_lo <= 1'b0;
    n2160_lo <= 1'b0;
    n2163_lo <= 1'b0;
    n2172_lo <= 1'b0;
    n2175_lo <= 1'b0;
    n2178_lo <= 1'b0;
    n2181_lo <= 1'b0;
    n2184_lo <= 1'b0;
    n2196_lo <= 1'b0;
    n2208_lo <= 1'b0;
    n2220_lo <= 1'b0;
    n2232_lo <= 1'b0;
    n2244_lo <= 1'b0;
    n2256_lo <= 1'b0;
    n2268_lo <= 1'b0;
    n2280_lo <= 1'b0;
    n2283_lo <= 1'b0;
    n2292_lo <= 1'b0;
    n2295_lo <= 1'b0;
    n2298_lo <= 1'b0;
    n2301_lo <= 1'b0;
    n2304_lo <= 1'b0;
    n2316_lo <= 1'b0;
    n2319_lo <= 1'b0;
    n2322_lo <= 1'b0;
    n2325_lo <= 1'b0;
    n2328_lo <= 1'b0;
    n2331_lo <= 1'b0;
    n2340_lo <= 1'b0;
    n2343_lo <= 1'b0;
    n2376_lo <= 1'b0;
    n2379_lo <= 1'b0;
    n2388_lo <= 1'b0;
    n2400_lo <= 1'b0;
    n2412_lo <= 1'b0;
    n2415_lo <= 1'b0;
    n2424_lo <= 1'b0;
    n2436_lo <= 1'b0;
    n2439_lo <= 1'b0;
    n2442_lo <= 1'b0;
    n2445_lo <= 1'b0;
    n2448_lo <= 1'b0;
    n2451_lo <= 1'b0;
    n2460_lo <= 1'b0;
    n2463_lo <= 1'b0;
    n2496_lo <= 1'b0;
    n2499_lo <= 1'b0;
    n2508_lo <= 1'b0;
    n2520_lo <= 1'b0;
    n2532_lo <= 1'b0;
    n2535_lo <= 1'b0;
    n2544_lo <= 1'b0;
    n2556_lo <= 1'b0;
    n2559_lo <= 1'b0;
    n2562_lo <= 1'b0;
    n2565_lo <= 1'b0;
    n2568_lo <= 1'b0;
    n2571_lo <= 1'b0;
    n2580_lo <= 1'b0;
    n2583_lo <= 1'b0;
    n2616_lo <= 1'b0;
    n2619_lo <= 1'b0;
    n2628_lo <= 1'b0;
    n2640_lo <= 1'b0;
    n2652_lo <= 1'b0;
    n2655_lo <= 1'b0;
    n2664_lo <= 1'b0;
    n2676_lo <= 1'b0;
    n2679_lo <= 1'b0;
    n2682_lo <= 1'b0;
    n2685_lo <= 1'b0;
    n2688_lo <= 1'b0;
    n2691_lo <= 1'b0;
    n2700_lo <= 1'b0;
    n2703_lo <= 1'b0;
    n2736_lo <= 1'b0;
    n2739_lo <= 1'b0;
    n2748_lo <= 1'b0;
    n2760_lo <= 1'b0;
    n2772_lo <= 1'b0;
    n2775_lo <= 1'b0;
    n2784_lo <= 1'b0;
    n2787_lo <= 1'b0;
    n2790_lo <= 1'b0;
    n2793_lo <= 1'b0;
    n2796_lo <= 1'b0;
    n2799_lo <= 1'b0;
    n2802_lo <= 1'b0;
    n2805_lo <= 1'b0;
    n2808_lo <= 1'b0;
    n2820_lo <= 1'b0;
    n2823_lo <= 1'b0;
    n2826_lo <= 1'b0;
    n2832_lo <= 1'b0;
    n2835_lo <= 1'b0;
    n2838_lo <= 1'b0;
    n2841_lo <= 1'b0;
    n2844_lo <= 1'b0;
    n2856_lo <= 1'b0;
    n2859_lo <= 1'b0;
    n2862_lo <= 1'b0;
    n2865_lo <= 1'b0;
    n2868_lo <= 1'b0;
    n2871_lo <= 1'b0;
    n2874_lo <= 1'b0;
    n2877_lo <= 1'b0;
    n2880_lo <= 1'b0;
    n2883_lo <= 1'b0;
    n2886_lo <= 1'b0;
    n2889_lo <= 1'b0;
    n2892_lo <= 1'b0;
    n2895_lo <= 1'b0;
    n2898_lo <= 1'b0;
    n2901_lo <= 1'b0;
    n2904_lo <= 1'b0;
    n2907_lo <= 1'b0;
    n2916_lo <= 1'b0;
    n2928_lo <= 1'b0;
    n2940_lo <= 1'b0;
    n2952_lo <= 1'b0;
    n2955_lo <= 1'b0;
    n2964_lo <= 1'b0;
    n2976_lo <= 1'b0;
    n2988_lo <= 1'b0;
    n2991_lo <= 1'b0;
    n3000_lo <= 1'b0;
    n3003_lo <= 1'b0;
    n3012_lo <= 1'b0;
    n3015_lo <= 1'b0;
    n3024_lo <= 1'b0;
    n3027_lo <= 1'b0;
    n3036_lo <= 1'b0;
    n3039_lo <= 1'b0;
    n3048_lo <= 1'b0;
    n3051_lo <= 1'b0;
    n3054_lo <= 1'b0;
    n3057_lo <= 1'b0;
    n3060_lo <= 1'b0;
    n3072_lo <= 1'b0;
    n3081_lo <= 1'b0;
    n3084_lo <= 1'b0;
    n3087_lo <= 1'b0;
    n3093_lo <= 1'b0;
    n3096_lo <= 1'b0;
    n3105_lo <= 1'b0;
    n3108_lo <= 1'b0;
    n3117_lo <= 1'b0;
    n3120_lo <= 1'b0;
    n3123_lo <= 1'b0;
    n3126_lo <= 1'b0;
    n3129_lo <= 1'b0;
    n3132_lo <= 1'b0;
    n3135_lo <= 1'b0;
    n3138_lo <= 1'b0;
    n3141_lo <= 1'b0;
    n3168_lo <= 1'b0;
    n3171_lo <= 1'b0;
    n3174_lo <= 1'b0;
    n3177_lo <= 1'b0;
    n3180_lo <= 1'b0;
    n3183_lo <= 1'b0;
    n3192_lo <= 1'b0;
    n3195_lo <= 1'b0;
    n3204_lo <= 1'b0;
    n3207_lo <= 1'b0;
    n3216_lo <= 1'b0;
    n3219_lo <= 1'b0;
    n3228_lo <= 1'b0;
    n3231_lo <= 1'b0;
    n3240_lo <= 1'b0;
    n3243_lo <= 1'b0;
    n3252_lo <= 1'b0;
    n3255_lo <= 1'b0;
    n3258_lo <= 1'b0;
    n3264_lo <= 1'b0;
    n3267_lo <= 1'b0;
    n3270_lo <= 1'b0;
    n3276_lo <= 1'b0;
    n3279_lo <= 1'b0;
    n3282_lo <= 1'b0;
    n3288_lo <= 1'b0;
    n3291_lo <= 1'b0;
    n3294_lo <= 1'b0;
    n4537_o2 <= 1'b0;
    n4538_o2 <= 1'b0;
    n4710_o2 <= 1'b0;
    n4711_o2 <= 1'b0;
    n1211_inv <= 1'b0;
    n1214_inv <= 1'b0;
    n1217_inv <= 1'b0;
    n1220_inv <= 1'b0;
    n4927_o2 <= 1'b0;
    n4928_o2 <= 1'b0;
    n1229_inv <= 1'b0;
    n1232_inv <= 1'b0;
    n1235_inv <= 1'b0;
    n5178_o2 <= 1'b0;
    n5179_o2 <= 1'b0;
    n5477_o2 <= 1'b0;
    n5478_o2 <= 1'b0;
    n5479_o2 <= 1'b0;
    n5222_o2 <= 1'b0;
    n5223_o2 <= 1'b0;
    n5553_o2 <= 1'b0;
    n5554_o2 <= 1'b0;
    G491_o2 <= 1'b0;
    n2922_lo_buf_o2 <= 1'b0;
    n2946_lo_buf_o2 <= 1'b0;
    n2970_lo_buf_o2 <= 1'b0;
    n2982_lo_buf_o2 <= 1'b0;
    n3066_lo_buf_o2 <= 1'b0;
    n3078_lo_buf_o2 <= 1'b0;
    n3102_lo_buf_o2 <= 1'b0;
    n3114_lo_buf_o2 <= 1'b0;
    G1321_o2 <= 1'b0;
    G1033_o2 <= 1'b0;
    G1030_o2 <= 1'b0;
    G1072_o2 <= 1'b0;
    n1304_inv <= 1'b0;
    n1307_inv <= 1'b0;
    n2958_lo_buf_o2 <= 1'b0;
    n2994_lo_buf_o2 <= 1'b0;
    n3006_lo_buf_o2 <= 1'b0;
    n3030_lo_buf_o2 <= 1'b0;
    n3042_lo_buf_o2 <= 1'b0;
    n3090_lo_buf_o2 <= 1'b0;
    n1328_inv <= 1'b0;
    n1331_inv <= 1'b0;
    n1334_inv <= 1'b0;
    n1337_inv <= 1'b0;
    n1340_inv <= 1'b0;
    n1343_inv <= 1'b0;
    n1346_inv <= 1'b0;
    n1349_inv <= 1'b0;
    G1036_o2 <= 1'b0;
    G1062_o2 <= 1'b0;
    G1067_o2 <= 1'b0;
    G1014_o2 <= 1'b0;
    n1364_inv <= 1'b0;
    n1367_inv <= 1'b0;
    n3018_lo_buf_o2 <= 1'b0;
    G766_o2 <= 1'b0;
    n1376_inv <= 1'b0;
    n1379_inv <= 1'b0;
    n1382_inv <= 1'b0;
    n1385_inv <= 1'b0;
    n1388_inv <= 1'b0;
    n1391_inv <= 1'b0;
    G1017_o2 <= 1'b0;
    G1008_o2 <= 1'b0;
    n1400_inv <= 1'b0;
    n1403_inv <= 1'b0;
    n2910_lo_buf_o2 <= 1'b0;
    n1409_inv <= 1'b0;
    G2138_o2 <= 1'b0;
    G2147_o2 <= 1'b0;
    n1418_inv <= 1'b0;
    G1137_o2 <= 1'b0;
    G1329_o2 <= 1'b0;
    G374_o2 <= 1'b0;
    G386_o2 <= 1'b0;
    G663_o2 <= 1'b0;
    G674_o2 <= 1'b0;
    G578_o2 <= 1'b0;
    G575_o2 <= 1'b0;
    G2505_o2 <= 1'b0;
    n1448_inv <= 1'b0;
    G987_o2 <= 1'b0;
    G984_o2 <= 1'b0;
    G1862_o2 <= 1'b0;
    G1859_o2 <= 1'b0;
    G1260_o2 <= 1'b0;
    G1865_o2 <= 1'b0;
    G2073_o2 <= 1'b0;
    G1402_o2 <= 1'b0;
    G2048_o2 <= 1'b0;
    G2276_o2 <= 1'b0;
    n1481_inv <= 1'b0;
    G2141_o2 <= 1'b0;
    G2008_o2 <= 1'b0;
    G2011_o2 <= 1'b0;
    G2150_o2 <= 1'b0;
    G2026_o2 <= 1'b0;
    G2029_o2 <= 1'b0;
    G2023_o2 <= 1'b0;
    G2041_o2 <= 1'b0;
    G2017_o2 <= 1'b0;
    G2020_o2 <= 1'b0;
    G2035_o2 <= 1'b0;
    G2038_o2 <= 1'b0;
    G2228_o2 <= 1'b0;
    G2231_o2 <= 1'b0;
    G2234_o2 <= 1'b0;
    G2237_o2 <= 1'b0;
    G1904_o2 <= 1'b0;
    G1907_o2 <= 1'b0;
    G1928_o2 <= 1'b0;
    G1931_o2 <= 1'b0;
    G1893_o2 <= 1'b0;
    G1896_o2 <= 1'b0;
    G1899_o2 <= 1'b0;
    G1937_o2 <= 1'b0;
    G1940_o2 <= 1'b0;
    G1943_o2 <= 1'b0;
    G1336_o2 <= 1'b0;
    G1996_o2 <= 1'b0;
    G1999_o2 <= 1'b0;
    G2002_o2 <= 1'b0;
    G2005_o2 <= 1'b0;
    G2014_o2 <= 1'b0;
    G2032_o2 <= 1'b0;
    G1076_o2 <= 1'b0;
    G1002_o2 <= 1'b0;
    G998_o2 <= 1'b0;
    G1890_o2 <= 1'b0;
    G1934_o2 <= 1'b0;
    G1044_o2 <= 1'b0;
    G1039_o2 <= 1'b0;
    n1770_lo_buf_o2 <= 1'b0;
    G342_o2 <= 1'b0;
    G354_o2 <= 1'b0;
    G1193_o2 <= 1'b0;
    n3234_lo_buf_o2 <= 1'b0;
    n3246_lo_buf_o2 <= 1'b0;
    G783_o2 <= 1'b0;
    G786_o2 <= 1'b0;
    G792_o2 <= 1'b0;
    G795_o2 <= 1'b0;
    G815_o2 <= 1'b0;
    G818_o2 <= 1'b0;
    G824_o2 <= 1'b0;
    G827_o2 <= 1'b0;
    G789_o2 <= 1'b0;
    G798_o2 <= 1'b0;
    G801_o2 <= 1'b0;
    G807_o2 <= 1'b0;
    G812_o2 <= 1'b0;
    G821_o2 <= 1'b0;
    G804_o2 <= 1'b0;
    G780_o2 <= 1'b0;
    G1231_o2 <= 1'b0;
    G1572_o2 <= 1'b0;
    G1377_o2 <= 1'b0;
    G1253_o2 <= 1'b0;
    G1359_o2 <= 1'b0;
    G1258_o2 <= 1'b0;
    G1367_o2 <= 1'b0;
    G1358_o2 <= 1'b0;
    G1366_o2 <= 1'b0;
    G2057_o2 <= 1'b0;
    G2117_o2 <= 1'b0;
    G2118_o2 <= 1'b0;
    G1254_o2 <= 1'b0;
    G1259_o2 <= 1'b0;
    G2058_o2 <= 1'b0;
    G405_o2 <= 1'b0;
    G417_o2 <= 1'b0;
    G1269_o2 <= 1'b0;
    G1275_o2 <= 1'b0;
    G1287_o2 <= 1'b0;
    G1266_o2 <= 1'b0;
    G1272_o2 <= 1'b0;
    G1278_o2 <= 1'b0;
    G1281_o2 <= 1'b0;
    G1284_o2 <= 1'b0;
    G1290_o2 <= 1'b0;
    G1293_o2 <= 1'b0;
    G1299_o2 <= 1'b0;
    G1305_o2 <= 1'b0;
    G1296_o2 <= 1'b0;
    G1302_o2 <= 1'b0;
    G1308_o2 <= 1'b0;
    G1311_o2 <= 1'b0;
    G811_o2 <= 1'b0;
    G810_o2 <= 1'b0;
    G1728_o2 <= 1'b0;
    G2512_o2 <= 1'b0;
    G1114_o2 <= 1'b0;
    G1113_o2 <= 1'b0;
    G1992_o2 <= 1'b0;
    G1991_o2 <= 1'b0;
    G1426_o2 <= 1'b0;
    G1966_o2 <= 1'b0;
    G2211_o2 <= 1'b0;
    G1509_o2 <= 1'b0;
    G2153_o2 <= 1'b0;
    G2329_o2 <= 1'b0;
    G1540_o2 <= 1'b0;
    G2167_o2 <= 1'b0;
    G2191_o2 <= 1'b0;
    G1234_o2 <= 1'b0;
    G1132_o2 <= 1'b0;
    G1129_o2 <= 1'b0;
    G2088_o2 <= 1'b0;
    G2106_o2 <= 1'b0;
    G1314_o2 <= 1'b0;
    G636_o2 <= 1'b0;
    G647_o2 <= 1'b0;
    n3186_lo_buf_o2 <= 1'b0;
    n3198_lo_buf_o2 <= 1'b0;
    n3210_lo_buf_o2 <= 1'b0;
    n3222_lo_buf_o2 <= 1'b0;
    G1225_o2 <= 1'b0;
    G1342_o2 <= 1'b0;
    G1222_o2 <= 1'b0;
    G1228_o2 <= 1'b0;
    G1348_o2 <= 1'b0;
    G1345_o2 <= 1'b0;
    G1351_o2 <= 1'b0;
    G2242_o2 <= 1'b0;
    G2260_o2 <= 1'b0;
    G1374_o2 <= 1'b0;
    G1537_o2 <= 1'b0;
    G301_o2 <= 1'b0;
    G313_o2 <= 1'b0;
    G2365_o2 <= 1'b0;
    G2255_o2 <= 1'b0;
    G2253_o2 <= 1'b0;
    G2395_o2 <= 1'b0;
    G2272_o2 <= 1'b0;
    G2270_o2 <= 1'b0;
    G2245_o2 <= 1'b0;
    G2262_o2 <= 1'b0;
    G2249_o2 <= 1'b0;
    G2247_o2 <= 1'b0;
    G2266_o2 <= 1'b0;
    G2264_o2 <= 1'b0;
    G2403_o2 <= 1'b0;
    G2401_o2 <= 1'b0;
    G2410_o2 <= 1'b0;
    G2408_o2 <= 1'b0;
    G2306_o2 <= 1'b0;
    G2305_o2 <= 1'b0;
    G2314_o2 <= 1'b0;
    G2313_o2 <= 1'b0;
    G2303_o2 <= 1'b0;
    G2302_o2 <= 1'b0;
    G2301_o2 <= 1'b0;
    G2311_o2 <= 1'b0;
    G2310_o2 <= 1'b0;
    G2309_o2 <= 1'b0;
    G2404_o2 <= 1'b0;
    G2411_o2 <= 1'b0;
    G2420_o2 <= 1'b0;
    G2419_o2 <= 1'b0;
    G2433_o2 <= 1'b0;
    G2432_o2 <= 1'b0;
    G402_o2 <= 1'b0;
    G403_o2 <= 1'b0;
    G1053_o2 <= 1'b0;
    G1049_o2 <= 1'b0;
    n2003_inv <= 1'b0;
    G1364_o2 <= 1'b0;
    G1079_o2 <= 1'b0;
    G1478_o2 <= 1'b0;
    G707_o2 <= 1'b0;
    G718_o2 <= 1'b0;
    G2417_o2 <= 1'b0;
    G2414_o2 <= 1'b0;
    G2431_o2 <= 1'b0;
    G2428_o2 <= 1'b0;
    G1653_o2 <= 1'b0;
    G2213_o2 <= 1'b0;
    G2221_o2 <= 1'b0;
    G2250_o2 <= 1'b0;
    G2267_o2 <= 1'b0;
    G1365_o2 <= 1'b0;
    G1368_o2 <= 1'b0;
    G1371_o2 <= 1'b0;
    G2218_o2 <= 1'b0;
    G2225_o2 <= 1'b0;
    n1503_lo_buf_o2 <= 1'b0;
    n1863_lo_buf_o2 <= 1'b0;
    n1887_lo_buf_o2 <= 1'b0;
    n1983_lo_buf_o2 <= 1'b0;
    n2007_lo_buf_o2 <= 1'b0;
    n2115_lo_buf_o2 <= 1'b0;
    n2139_lo_buf_o2 <= 1'b0;
    n2247_lo_buf_o2 <= 1'b0;
    n2271_lo_buf_o2 <= 1'b0;
    n2919_lo_buf_o2 <= 1'b0;
    n2943_lo_buf_o2 <= 1'b0;
    n2967_lo_buf_o2 <= 1'b0;
    n2979_lo_buf_o2 <= 1'b0;
    n3063_lo_buf_o2 <= 1'b0;
    n3075_lo_buf_o2 <= 1'b0;
    n3099_lo_buf_o2 <= 1'b0;
    n3111_lo_buf_o2 <= 1'b0;
    G878_o2 <= 1'b0;
    G875_o2 <= 1'b0;
    G661_o2 <= 1'b0;
    G660_o2 <= 1'b0;
    G879_o2 <= 1'b0;
    G876_o2 <= 1'b0;
    G1320_o2 <= 1'b0;
    G941_o2 <= 1'b0;
    G732_o2 <= 1'b0;
    G942_o2 <= 1'b0;
    G1493_o2 <= 1'b0;
    G1498_o2 <= 1'b0;
    G877_o2 <= 1'b0;
    G874_o2 <= 1'b0;
    n1806_lo_buf_o2 <= 1'b0;
    n1878_lo_buf_o2 <= 1'b0;
    n1938_lo_buf_o2 <= 1'b0;
    n1998_lo_buf_o2 <= 1'b0;
    n2058_lo_buf_o2 <= 1'b0;
    n2130_lo_buf_o2 <= 1'b0;
    n2190_lo_buf_o2 <= 1'b0;
    n2262_lo_buf_o2 <= 1'b0;
    n2310_lo_buf_o2 <= 1'b0;
    n2406_lo_buf_o2 <= 1'b0;
    n2430_lo_buf_o2 <= 1'b0;
    n2526_lo_buf_o2 <= 1'b0;
    n2550_lo_buf_o2 <= 1'b0;
    n2646_lo_buf_o2 <= 1'b0;
    n2670_lo_buf_o2 <= 1'b0;
    n2766_lo_buf_o2 <= 1'b0;
    G603_o2 <= 1'b0;
    G614_o2 <= 1'b0;
    G1026_o2 <= 1'b0;
    G1021_o2 <= 1'b0;
    G940_o2 <= 1'b0;
    G1636_o2 <= 1'b0;
    G1684_o2 <= 1'b0;
    n2352_lo_buf_o2 <= 1'b0;
    n2364_lo_buf_o2 <= 1'b0;
    n2472_lo_buf_o2 <= 1'b0;
    n2484_lo_buf_o2 <= 1'b0;
    n2592_lo_buf_o2 <= 1'b0;
    n2604_lo_buf_o2 <= 1'b0;
    n2712_lo_buf_o2 <= 1'b0;
    n2724_lo_buf_o2 <= 1'b0;
    n3150_lo_buf_o2 <= 1'b0;
    n3162_lo_buf_o2 <= 1'b0;
  end
endmodule


