// Benchmark "c1908" written by ABC on Sun Oct 29 19:31:51 2023

module c1908 (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33,
    G1884, G1885, G1886, G1887, G1888, G1889, G1890, G1891, G1892, G1893,
    G1894, G1895, G1896, G1897, G1898, G1899, G1900, G1901, G1902, G1903,
    G1904, G1905, G1906, G1907, G1908  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33;
  output G1884, G1885, G1886, G1887, G1888, G1889, G1890, G1891, G1892, G1893,
    G1894, G1895, G1896, G1897, G1898, G1899, G1900, G1901, G1902, G1903,
    G1904, G1905, G1906, G1907, G1908;
  reg n940_lo, n943_lo, n946_lo, n949_lo, n952_lo, n955_lo, n958_lo,
    n961_lo, n964_lo, n967_lo, n970_lo, n973_lo, n976_lo, n979_lo, n982_lo,
    n985_lo, n988_lo, n991_lo, n994_lo, n997_lo, n1000_lo, n1003_lo,
    n1006_lo, n1009_lo, n1012_lo, n1015_lo, n1018_lo, n1021_lo, n1024_lo,
    n1027_lo, n1030_lo, n1033_lo, n1036_lo, n1039_lo, n1042_lo, n1045_lo,
    n1048_lo, n1051_lo, n1054_lo, n1057_lo, n1060_lo, n1063_lo, n1066_lo,
    n1069_lo, n1072_lo, n1075_lo, n1078_lo, n1081_lo, n1084_lo, n1087_lo,
    n1090_lo, n1093_lo, n1096_lo, n1099_lo, n1102_lo, n1105_lo, n1108_lo,
    n1111_lo, n1114_lo, n1117_lo, n1120_lo, n1123_lo, n1126_lo, n1129_lo,
    n1132_lo, n1135_lo, n1138_lo, n1141_lo, n1144_lo, n1147_lo, n1150_lo,
    n1153_lo, n1156_lo, n1159_lo, n1162_lo, n1165_lo, n1168_lo, n1171_lo,
    n1174_lo, n1177_lo, n1180_lo, n1183_lo, n1186_lo, n1189_lo, n1192_lo,
    n1195_lo, n1198_lo, n1201_lo, n1204_lo, n1207_lo, n1210_lo, n1213_lo,
    n1216_lo, n1219_lo, n1222_lo, n1225_lo, n1228_lo, n1231_lo, n1234_lo,
    n1237_lo, n1240_lo, n1243_lo, n1246_lo, n1249_lo, n1252_lo, n1255_lo,
    n1258_lo, n1261_lo, n1264_lo, n1267_lo, n1270_lo, n1273_lo, n1276_lo,
    n1279_lo, n1282_lo, n1285_lo, n1288_lo, n1291_lo, n1294_lo, n1297_lo,
    n1300_lo, n1303_lo, n1306_lo, n1309_lo, n1312_lo, n1315_lo, n1318_lo,
    n1321_lo, n1324_lo, n1327_lo, n1330_lo, n1333_lo;
  wire new_G112_, new_G116_, new_G119_, new_G123_, new_G128_, new_G131_,
    new_G134_, new_G138_, new_G142_, new_G147_, new_G151_, new_G154_,
    new_G157_, new_G161_, new_G165_, new_G169_, new_G173_, new_G174_,
    new_G175_, new_G178_, new_G179_, new_G182_, new_G185_, new_G188_,
    new_G191_, new_G194_, new_G197_, new_G198_, new_G199_, new_G202_,
    new_G205_, new_G212_, new_G219_, new_G222_, new_G225_, new_G228_,
    new_G235_, new_G238_, new_G241_, new_G248_, new_G253_, new_G260_,
    new_G265_, new_G268_, new_G271_, new_G274_, new_G277_, new_G280_,
    new_G283_, new_G286_, new_G289_, new_G292_, new_G295_, new_G298_,
    new_G301_, new_G304_, new_G307_, new_G310_, new_G313_, new_G314_,
    new_G315_, new_G316_, new_G317_, new_G318_, new_G319_, new_G320_,
    new_G321_, new_G322_, new_G323_, new_G324_, new_G325_, new_G326_,
    new_G327_, new_G328_, new_G329_, new_G330_, new_G331_, new_G332_,
    new_G333_, new_G334_, new_G335_, new_G338_, new_G341_, new_G344_,
    new_G347_, new_G350_, new_G353_, new_G356_, new_G359_, new_G362_,
    new_G365_, new_G368_, new_G371_, new_G374_, new_G377_, new_G380_,
    new_G381_, new_G382_, new_G387_, new_G391_, new_G395_, new_G398_,
    new_G401_, new_G404_, new_G407_, new_G410_, new_G413_, new_G416_,
    new_G419_, new_G422_, new_G425_, new_G428_, new_G431_, new_G434_,
    new_G437_, new_G440_, new_G443_, new_G446_, new_G449_, new_G452_,
    new_G455_, new_G458_, new_G461_, new_G464_, new_G467_, new_G470_,
    new_G473_, new_G476_, new_G479_, new_G482_, new_G485_, new_G488_,
    new_G491_, new_G494_, new_G497_, new_G500_, new_G503_, new_G506_,
    new_G509_, new_G512_, new_G515_, new_G518_, new_G521_, new_G524_,
    new_G527_, new_G530_, new_G533_, new_G534_, new_G535_, new_G536_,
    new_G537_, new_G538_, new_G539_, new_G540_, new_G541_, new_G542_,
    new_G543_, new_G544_, new_G545_, new_G546_, new_G550_, new_G554_,
    new_G557_, new_G560_, new_G561_, new_G562_, new_G563_, new_G564_,
    new_G565_, new_G566_, new_G567_, new_G568_, new_G569_, new_G570_,
    new_G573_, new_G582_, new_G585_, new_G586_, new_G589_, new_G590_,
    new_G593_, new_G594_, new_G597_, new_G598_, new_G601_, new_G602_,
    new_G605_, new_G606_, new_G609_, new_G612_, new_G615_, new_G616_,
    new_G619_, new_G620_, new_G623_, new_G624_, new_G627_, new_G628_,
    new_G631_, new_G632_, new_G635_, new_G636_, new_G637_, new_G638_,
    new_G639_, new_G640_, new_G641_, new_G644_, new_G645_, new_G648_,
    new_G649_, new_G650_, new_G651_, new_G652_, new_G653_, new_G654_,
    new_G655_, new_G656_, new_G657_, new_G660_, new_G663_, new_G666_,
    new_G669_, new_G672_, new_G675_, new_G678_, new_G681_, new_G684_,
    new_G687_, new_G690_, new_G693_, new_G696_, new_G699_, new_G700_,
    new_G701_, new_G702_, new_G703_, new_G704_, new_G705_, new_G706_,
    new_G707_, new_G708_, new_G709_, new_G710_, new_G711_, new_G712_,
    new_G713_, new_G714_, new_G715_, new_G716_, new_G717_, new_G718_,
    new_G719_, new_G720_, new_G721_, new_G722_, new_G723_, new_G724_,
    new_G725_, new_G726_, new_G727_, new_G728_, new_G729_, new_G730_,
    new_G731_, new_G734_, new_G735_, new_G738_, new_G755_, new_G772_,
    new_G773_, new_G774_, new_G775_, new_G776_, new_G777_, new_G778_,
    new_G779_, new_G780_, new_G781_, new_G782_, new_G783_, new_G784_,
    new_G785_, new_G786_, new_G787_, new_G788_, new_G789_, new_G790_,
    new_G791_, new_G792_, new_G793_, new_G794_, new_G795_, new_G796_,
    new_G797_, new_G798_, new_G799_, new_G802_, new_G805_, new_G806_,
    new_G807_, new_G808_, new_G809_, new_G810_, new_G813_, new_G816_,
    new_G819_, new_G822_, new_G825_, new_G828_, new_G831_, new_G834_,
    new_G835_, new_G836_, new_G837_, new_G838_, new_G839_, new_G840_,
    new_G841_, new_G842_, new_G843_, new_G844_, new_G845_, new_G848_,
    new_G849_, new_G850_, new_G851_, new_G854_, new_G855_, new_G856_,
    new_G857_, new_G858_, new_G859_, new_G860_, new_G861_, new_G864_,
    new_G867_, new_G870_, new_G873_, new_G876_, new_G879_, new_G882_,
    new_G885_, new_G888_, new_G891_, new_G894_, new_G895_, new_G896_,
    new_G897_, new_G898_, new_G901_, new_G904_, new_G905_, new_G906_,
    new_G907_, new_G908_, new_G909_, new_G910_, new_G911_, new_G914_,
    new_G917_, new_G918_, new_G919_, new_G920_, new_G921_, new_G924_,
    new_G925_, new_G926_, new_G927_, new_G928_, new_G929_, new_G930_,
    new_G931_, new_G932_, new_G933_, new_G934_, new_G935_, new_G936_,
    new_G937_, new_G938_, new_G939_, new_G940_, new_G941_, new_G942_,
    new_G943_, new_G944_, new_G945_, new_G946_, new_G947_, new_G948_,
    new_G951_, new_G952_, new_G953_, new_G956_, new_G959_, new_G962_,
    new_G963_, new_G964_, new_G965_, new_G966_, new_G967_, new_G968_,
    new_G969_, new_G970_, new_G971_, new_G972_, new_G973_, new_G974_,
    new_G975_, new_G976_, new_G977_, new_G980_, new_G981_, new_G984_,
    new_G987_, new_G988_, new_G989_, new_G993_, new_G994_, new_G995_,
    new_G996_, new_G997_, new_G998_, new_G999_, new_G1000_, new_G1003_,
    new_G1006_, new_G1009_, new_G1012_, new_G1015_, new_G1019_, new_G1022_,
    new_G1023_, new_G1024_, new_G1025_, new_G1028_, new_G1031_, new_G1034_,
    new_G1035_, new_G1036_, new_G1037_, new_G1038_, new_G1041_, new_G1044_,
    new_G1047_, new_G1050_, new_G1053_, new_G1056_, new_G1059_, new_G1062_,
    new_G1065_, new_G1066_, new_G1067_, new_G1068_, new_G1069_, new_G1072_,
    new_G1075_, new_G1078_, new_G1081_, new_G1084_, new_G1087_, new_G1090_,
    new_G1091_, new_G1092_, new_G1093_, new_G1094_, new_G1095_, new_G1096_,
    new_G1097_, new_G1098_, new_G1099_, new_G1100_, new_G1103_, new_G1104_,
    new_G1107_, new_G1110_, new_G1111_, new_G1112_, new_G1113_, new_G1114_,
    new_G1115_, new_G1116_, new_G1117_, new_G1118_, new_G1121_, new_G1124_,
    new_G1125_, new_G1126_, new_G1129_, new_G1130_, new_G1131_, new_G1132_,
    new_G1135_, new_G1138_, new_G1139_, new_G1140_, new_G1143_, new_G1144_,
    new_G1145_, new_G1148_, new_G1151_, new_G1152_, new_G1153_, new_G1154_,
    new_G1155_, new_G1156_, new_G1157_, new_G1158_, new_G1159_, new_G1160_,
    new_G1163_, new_G1166_, new_G1167_, new_G1168_, new_G1169_, new_G1170_,
    new_G1171_, new_G1174_, new_G1175_, new_G1176_, new_G1177_, new_G1178_,
    new_G1181_, new_G1182_, new_G1185_, new_G1186_, new_G1187_, new_G1188_,
    new_G1189_, new_G1192_, new_G1195_, new_G1198_, new_G1199_, new_G1200_,
    new_G1201_, new_G1202_, new_G1203_, new_G1204_, new_G1205_, new_G1208_,
    new_G1209_, new_G1212_, new_G1215_, new_G1216_, new_G1217_, new_G1218_,
    new_G1219_, new_G1220_, new_G1221_, new_G1222_, new_G1225_, new_G1226_,
    new_G1227_, new_G1230_, new_G1233_, new_G1236_, new_G1239_, new_G1240_,
    new_G1243_, new_G1244_, new_G1245_, new_G1246_, new_G1247_, new_G1250_,
    new_G1251_, new_G1252_, new_G1253_, new_G1256_, new_G1259_, new_G1260_,
    new_G1261_, new_G1262_, new_G1263_, new_G1264_, new_G1265_, new_G1266_,
    new_G1267_, new_G1268_, new_G1269_, new_G1270_, new_G1273_, new_G1276_,
    new_G1279_, new_G1280_, new_G1281_, new_G1282_, new_G1283_, new_G1284_,
    new_G1287_, new_G1290_, new_G1293_, new_G1296_, new_G1299_, new_G1302_,
    new_G1305_, new_G1308_, new_G1309_, new_G1310_, new_G1311_, new_G1312_,
    new_G1313_, new_G1316_, new_G1317_, new_G1320_, new_G1321_, new_G1322_,
    new_G1323_, new_G1324_, new_G1325_, new_G1326_, new_G1327_, new_G1328_,
    new_G1329_, new_G1330_, new_G1331_, new_G1332_, new_G1333_, new_G1334_,
    new_G1335_, new_G1336_, new_G1337_, new_G1338_, new_G1339_, new_G1340_,
    new_G1341_, new_G1342_, new_G1343_, new_G1344_, new_G1347_, new_G1350_,
    new_G1353_, new_G1354_, new_G1355_, new_G1356_, new_G1357_, new_G1358_,
    new_G1359_, new_G1362_, new_G1363_, new_G1366_, new_G1369_, new_G1370_,
    new_G1371_, new_G1374_, new_G1375_, new_G1378_, new_G1381_, new_G1382_,
    new_G1383_, new_G1386_, new_G1389_, new_G1392_, new_G1395_, new_G1410_,
    new_G1420_, new_G1434_, new_G1439_, new_G1442_, new_G1445_, new_G1448_,
    new_G1451_, new_G1454_, new_G1457_, new_G1458_, new_G1459_, new_G1460_,
    new_G1461_, new_G1462_, new_G1463_, new_G1464_, new_G1465_, new_G1466_,
    new_G1467_, new_G1468_, new_G1469_, new_G1470_, new_G1471_, new_G1472_,
    new_G1473_, new_G1474_, new_G1475_, new_G1476_, new_G1479_, new_G1480_,
    new_G1483_, new_G1484_, new_G1487_, new_G1488_, new_G1489_, new_G1490_,
    new_G1493_, new_G1496_, new_G1499_, new_G1502_, new_G1505_, new_G1508_,
    new_G1511_, new_G1522_, new_G1538_, new_G1549_, new_G1563_, new_G1576_,
    new_G1584_, new_G1598_, new_G1607_, new_G1608_, new_G1609_, new_G1624_,
    new_G1625_, new_G1642_, new_G1645_, new_G1648_, new_G1651_, new_G1654_,
    new_G1657_, new_G1660_, new_G1663_, new_G1666_, new_G1669_, new_G1672_,
    new_G1675_, new_G1678_, new_G1681_, new_G1684_, new_G1687_, new_G1690_,
    new_G1693_, new_G1696_, new_G1699_, new_G1702_, new_G1705_, new_G1708_,
    new_G1711_, new_G1712_, new_G1713_, new_G1714_, new_G1715_, new_G1716_,
    new_G1717_, new_G1718_, new_G1719_, new_G1722_, new_G1725_, new_G1728_,
    new_G1731_, new_G1734_, new_G1737_, new_G1740_, new_G1743_, new_G1746_,
    new_G1747_, new_G1748_, new_G1749_, new_G1750_, new_G1751_, new_G1752_,
    new_G1753_, new_G1754_, new_G1755_, new_G1756_, new_G1757_, new_G1758_,
    new_G1759_, new_G1760_, new_G1761_, new_G1762_, new_G1763_, new_G1764_,
    new_G1765_, new_G1766_, new_G1767_, new_G1768_, new_G1769_, new_G1770_,
    new_G1771_, new_G1772_, new_G1773_, new_G1774_, new_G1775_, new_G1776_,
    new_G1777_, new_G1778_, new_G1779_, new_G1780_, new_G1781_, new_G1782_,
    new_G1783_, new_G1784_, new_G1785_, new_G1786_, new_G1787_, new_G1788_,
    new_G1791_, new_G1794_, new_G1795_, new_G1796_, new_G1797_, new_G1798_,
    new_G1799_, new_G1800_, new_G1801_, new_G1802_, new_G1803_, new_G1806_,
    new_G1809_, new_G1810_, new_G1817_, new_G1818_, new_G1819_, new_G1820_,
    new_G1821_, new_G1822_, new_G1825_, new_G1828_, new_G1831_, new_G1834_,
    new_G1837_, new_G1838_, new_G1839_, new_G1842_, new_G1845_, new_G1848_,
    new_G1849_, new_G1850_, new_G1851_, new_G1852_, new_G1853_, new_G1854_,
    new_G1855_, new_G1856_, new_G1857_, new_G1858_, new_G1859_, new_G1860_,
    new_G1861_, new_G1862_, new_G1863_, new_G1864_, new_G1865_, new_G1866_,
    new_G1867_, new_G1868_, new_G1869_, new_G1870_, new_G1871_, new_G1872_,
    new_G1873_, new_G1874_, new_G1875_, new_G1876_, new_G1877_, new_G1880_,
    new_G1881_, new_G1882_, new_G1883_, n940_li, n943_li, n946_li, n949_li,
    n952_li, n955_li, n958_li, n961_li, n964_li, n967_li, n970_li, n973_li,
    n976_li, n979_li, n982_li, n985_li, n988_li, n991_li, n994_li, n997_li,
    n1000_li, n1003_li, n1006_li, n1009_li, n1012_li, n1015_li, n1018_li,
    n1021_li, n1024_li, n1027_li, n1030_li, n1033_li, n1036_li, n1039_li,
    n1042_li, n1045_li, n1048_li, n1051_li, n1054_li, n1057_li, n1060_li,
    n1063_li, n1066_li, n1069_li, n1072_li, n1075_li, n1078_li, n1081_li,
    n1084_li, n1087_li, n1090_li, n1093_li, n1096_li, n1099_li, n1102_li,
    n1105_li, n1108_li, n1111_li, n1114_li, n1117_li, n1120_li, n1123_li,
    n1126_li, n1129_li, n1132_li, n1135_li, n1138_li, n1141_li, n1144_li,
    n1147_li, n1150_li, n1153_li, n1156_li, n1159_li, n1162_li, n1165_li,
    n1168_li, n1171_li, n1174_li, n1177_li, n1180_li, n1183_li, n1186_li,
    n1189_li, n1192_li, n1195_li, n1198_li, n1201_li, n1204_li, n1207_li,
    n1210_li, n1213_li, n1216_li, n1219_li, n1222_li, n1225_li, n1228_li,
    n1231_li, n1234_li, n1237_li, n1240_li, n1243_li, n1246_li, n1249_li,
    n1252_li, n1255_li, n1258_li, n1261_li, n1264_li, n1267_li, n1270_li,
    n1273_li, n1276_li, n1279_li, n1282_li, n1285_li, n1288_li, n1291_li,
    n1294_li, n1297_li, n1300_li, n1303_li, n1306_li, n1309_li, n1312_li,
    n1315_li, n1318_li, n1321_li, n1324_li, n1327_li, n1330_li, n1333_li;
  assign new_G112_ = ~n949_lo;
  assign new_G116_ = ~n961_lo;
  assign new_G119_ = ~n973_lo;
  assign new_G123_ = ~n985_lo;
  assign new_G128_ = ~n997_lo;
  assign new_G131_ = ~n1009_lo;
  assign new_G134_ = ~n1021_lo;
  assign new_G138_ = ~n1033_lo;
  assign new_G142_ = ~n1045_lo;
  assign new_G147_ = ~n1057_lo;
  assign new_G151_ = ~n1069_lo;
  assign new_G154_ = ~n1081_lo;
  assign new_G157_ = ~n1093_lo;
  assign new_G161_ = ~n1105_lo;
  assign new_G165_ = ~n1117_lo;
  assign new_G169_ = ~n1129_lo;
  assign new_G173_ = ~n1189_lo | ~n1285_lo;
  assign new_G174_ = ~n1201_lo | ~n1297_lo;
  assign new_G175_ = ~n1225_lo;
  assign new_G178_ = ~n1225_lo;
  assign new_G179_ = ~n1213_lo;
  assign new_G182_ = ~n1213_lo;
  assign new_G185_ = ~n1237_lo;
  assign new_G188_ = ~n1249_lo;
  assign new_G191_ = ~n1261_lo;
  assign new_G194_ = ~n1273_lo;
  assign new_G197_ = ~n1333_lo;
  assign new_G198_ = ~n1333_lo;
  assign new_G199_ = ~n1285_lo;
  assign new_G202_ = ~n1297_lo;
  assign new_G205_ = ~n1309_lo;
  assign new_G212_ = ~n1309_lo;
  assign new_G219_ = ~n1309_lo;
  assign new_G222_ = ~n1309_lo;
  assign new_G225_ = ~n1321_lo;
  assign new_G228_ = ~n1321_lo;
  assign new_G235_ = ~n1321_lo;
  assign new_G238_ = ~n1333_lo;
  assign new_G241_ = ~n1333_lo;
  assign new_G248_ = ~n1333_lo;
  assign new_G253_ = ~n1333_lo;
  assign new_G260_ = ~n1333_lo;
  assign new_G265_ = ~n949_lo;
  assign new_G268_ = ~n961_lo;
  assign new_G271_ = ~n973_lo;
  assign new_G274_ = ~n985_lo;
  assign new_G277_ = ~n997_lo;
  assign new_G280_ = ~n1009_lo;
  assign new_G283_ = ~n1021_lo;
  assign new_G286_ = ~n1033_lo;
  assign new_G289_ = ~n1045_lo;
  assign new_G292_ = ~n1057_lo;
  assign new_G295_ = ~n1069_lo;
  assign new_G298_ = ~n1081_lo;
  assign new_G301_ = ~n1093_lo;
  assign new_G304_ = ~n1105_lo;
  assign new_G307_ = ~n1117_lo;
  assign new_G310_ = ~n1129_lo;
  assign new_G313_ = ~new_G265_;
  assign new_G314_ = ~new_G268_;
  assign new_G315_ = ~new_G271_;
  assign new_G316_ = ~new_G274_;
  assign new_G317_ = ~new_G277_;
  assign new_G318_ = ~new_G280_;
  assign new_G319_ = ~new_G283_;
  assign new_G320_ = ~new_G286_;
  assign new_G321_ = ~new_G289_;
  assign new_G322_ = ~new_G292_;
  assign new_G323_ = ~new_G295_;
  assign new_G324_ = ~new_G298_;
  assign new_G325_ = ~new_G301_;
  assign new_G326_ = ~new_G304_;
  assign new_G327_ = ~new_G307_;
  assign new_G328_ = ~new_G310_;
  assign new_G329_ = ~new_G228_ | ~new_G253_;
  assign new_G330_ = ~new_G228_ | ~new_G253_;
  assign new_G331_ = ~new_G228_ | ~new_G253_;
  assign new_G332_ = ~new_G228_ | ~new_G253_;
  assign new_G333_ = ~new_G228_ | ~new_G253_;
  assign new_G334_ = ~new_G228_ | ~new_G253_;
  assign new_G335_ = ~new_G112_;
  assign new_G338_ = ~new_G116_;
  assign new_G341_ = ~new_G128_;
  assign new_G344_ = ~new_G131_;
  assign new_G347_ = ~new_G147_;
  assign new_G350_ = ~new_G165_;
  assign new_G353_ = n1189_lo & new_G241_;
  assign new_G356_ = ~new_G142_;
  assign new_G359_ = ~new_G151_;
  assign new_G362_ = ~new_G154_;
  assign new_G365_ = n1201_lo & new_G241_;
  assign new_G368_ = ~new_G161_;
  assign new_G371_ = n1141_lo & new_G175_ & new_G241_;
  assign new_G374_ = ~new_G169_;
  assign new_G377_ = ~new_G161_;
  assign new_G380_ = ~new_G248_ | ~new_G199_;
  assign new_G381_ = ~new_G248_ | ~new_G202_;
  assign new_G382_ = ~new_G182_ | ~n1225_lo;
  assign new_G387_ = ~new_G182_ | ~new_G222_;
  assign new_G391_ = ~new_G178_ | ~new_G222_;
  assign new_G395_ = ~new_G123_;
  assign new_G398_ = ~new_G138_;
  assign new_G401_ = ~new_G142_;
  assign new_G404_ = ~new_G161_;
  assign new_G407_ = ~new_G112_;
  assign new_G410_ = ~new_G112_;
  assign new_G413_ = ~new_G116_;
  assign new_G416_ = ~new_G151_;
  assign new_G419_ = ~new_G119_;
  assign new_G422_ = n1165_lo & new_G179_ & new_G241_;
  assign new_G425_ = ~new_G154_;
  assign new_G428_ = ~new_G123_;
  assign new_G431_ = ~new_G157_;
  assign new_G434_ = n1177_lo & new_G179_ & new_G241_;
  assign new_G437_ = ~new_G185_;
  assign new_G440_ = ~new_G185_;
  assign new_G443_ = ~new_G188_;
  assign new_G446_ = ~new_G188_;
  assign new_G449_ = ~new_G191_;
  assign new_G452_ = ~new_G191_;
  assign new_G455_ = ~new_G194_;
  assign new_G458_ = ~new_G194_;
  assign new_G461_ = new_G173_ & new_G238_;
  assign new_G464_ = new_G174_ & new_G238_;
  assign new_G467_ = ~new_G119_;
  assign new_G470_ = ~new_G119_;
  assign new_G473_ = ~new_G134_;
  assign new_G476_ = ~new_G134_;
  assign new_G479_ = ~new_G169_;
  assign new_G482_ = ~new_G169_;
  assign new_G485_ = ~new_G157_;
  assign new_G488_ = ~new_G157_;
  assign new_G491_ = ~new_G123_;
  assign new_G494_ = ~new_G123_;
  assign new_G497_ = ~new_G128_;
  assign new_G500_ = ~new_G138_;
  assign new_G503_ = n1153_lo & new_G175_ & new_G241_;
  assign new_G506_ = ~new_G165_;
  assign new_G509_ = ~new_G142_;
  assign new_G512_ = ~new_G142_;
  assign new_G515_ = ~new_G131_;
  assign new_G518_ = ~new_G138_;
  assign new_G521_ = ~new_G147_;
  assign new_G524_ = ~new_G165_;
  assign new_G527_ = ~new_G134_;
  assign new_G530_ = ~new_G147_;
  assign new_G533_ = ~new_G461_;
  assign new_G534_ = ~new_G464_;
  assign new_G535_ = ~new_G395_;
  assign new_G536_ = ~new_G398_;
  assign new_G537_ = ~new_G401_;
  assign new_G538_ = ~new_G404_;
  assign new_G539_ = ~new_G410_;
  assign new_G540_ = ~new_G422_;
  assign new_G541_ = ~new_G428_;
  assign new_G542_ = ~new_G431_;
  assign new_G543_ = ~new_G434_;
  assign new_G544_ = n1141_lo & new_G391_;
  assign new_G545_ = n1165_lo & new_G387_;
  assign new_G546_ = ~n1153_lo | ~new_G391_;
  assign new_G550_ = ~n1177_lo | ~new_G387_;
  assign new_G554_ = ~n1141_lo | ~new_G391_;
  assign new_G557_ = ~n1165_lo | ~new_G387_;
  assign new_G560_ = ~new_G440_;
  assign new_G561_ = ~new_G437_;
  assign new_G562_ = ~new_G446_;
  assign new_G563_ = ~new_G443_;
  assign new_G564_ = ~new_G452_;
  assign new_G565_ = ~new_G449_;
  assign new_G566_ = ~new_G458_;
  assign new_G567_ = ~new_G455_;
  assign new_G568_ = ~new_G199_ | ~new_G219_ | ~new_G248_ | ~new_G382_;
  assign new_G569_ = ~new_G202_ | ~new_G219_ | ~new_G248_ | ~new_G382_;
  assign new_G570_ = ~new_G225_ | ~new_G260_ | ~new_G382_;
  assign new_G573_ = new_G225_ & new_G260_ & new_G382_;
  assign new_G582_ = ~new_G335_;
  assign new_G585_ = ~new_G467_;
  assign new_G586_ = ~new_G335_;
  assign new_G589_ = ~new_G470_;
  assign new_G590_ = ~new_G341_;
  assign new_G593_ = ~new_G473_;
  assign new_G594_ = ~new_G341_;
  assign new_G597_ = ~new_G476_;
  assign new_G598_ = ~new_G347_;
  assign new_G601_ = ~new_G479_;
  assign new_G602_ = ~new_G347_;
  assign new_G605_ = ~new_G482_;
  assign new_G606_ = ~new_G353_;
  assign new_G609_ = ~new_G353_;
  assign new_G612_ = ~new_G359_;
  assign new_G615_ = ~new_G485_;
  assign new_G616_ = ~new_G359_;
  assign new_G619_ = ~new_G488_;
  assign new_G620_ = ~new_G365_;
  assign new_G623_ = ~new_G491_;
  assign new_G624_ = ~new_G365_;
  assign new_G627_ = ~new_G494_;
  assign new_G628_ = ~new_G371_;
  assign new_G631_ = ~new_G407_;
  assign new_G632_ = ~new_G371_;
  assign new_G635_ = ~new_G497_;
  assign new_G636_ = ~new_G500_;
  assign new_G637_ = ~new_G413_;
  assign new_G638_ = ~new_G503_;
  assign new_G639_ = ~new_G506_;
  assign new_G640_ = ~new_G416_;
  assign new_G641_ = ~new_G374_;
  assign new_G644_ = ~new_G509_;
  assign new_G645_ = ~new_G374_;
  assign new_G648_ = ~new_G512_;
  assign new_G649_ = ~new_G515_;
  assign new_G650_ = ~new_G518_;
  assign new_G651_ = ~new_G419_;
  assign new_G652_ = ~new_G521_;
  assign new_G653_ = ~new_G524_;
  assign new_G654_ = ~new_G425_;
  assign new_G655_ = ~new_G527_;
  assign new_G656_ = ~new_G530_;
  assign new_G657_ = ~new_G338_;
  assign new_G660_ = ~new_G338_;
  assign new_G663_ = ~new_G344_;
  assign new_G666_ = ~new_G344_;
  assign new_G669_ = ~new_G350_;
  assign new_G672_ = ~new_G350_;
  assign new_G675_ = ~new_G356_;
  assign new_G678_ = ~new_G356_;
  assign new_G681_ = ~new_G362_;
  assign new_G684_ = ~new_G362_;
  assign new_G687_ = ~new_G368_;
  assign new_G690_ = ~new_G368_;
  assign new_G693_ = ~new_G377_;
  assign new_G696_ = ~new_G377_;
  assign new_G699_ = ~new_G398_ | ~new_G535_;
  assign new_G700_ = ~new_G395_ | ~new_G536_;
  assign new_G701_ = ~new_G404_ | ~new_G537_;
  assign new_G702_ = ~new_G401_ | ~new_G538_;
  assign new_G703_ = ~new_G434_ | ~new_G542_;
  assign new_G704_ = ~new_G431_ | ~new_G543_;
  assign new_G705_ = ~new_G500_ | ~new_G635_;
  assign new_G706_ = ~new_G497_ | ~new_G636_;
  assign new_G707_ = ~new_G506_ | ~new_G638_;
  assign new_G708_ = ~new_G503_ | ~new_G639_;
  assign new_G709_ = ~new_G518_ | ~new_G649_;
  assign new_G710_ = ~new_G515_ | ~new_G650_;
  assign new_G711_ = ~new_G524_ | ~new_G652_;
  assign new_G712_ = ~new_G521_ | ~new_G653_;
  assign new_G713_ = ~new_G530_ | ~new_G655_;
  assign new_G714_ = ~new_G527_ | ~new_G656_;
  assign new_G715_ = ~new_G586_;
  assign new_G716_ = ~new_G582_;
  assign new_G717_ = ~new_G699_ | ~new_G700_;
  assign new_G718_ = ~new_G590_;
  assign new_G719_ = ~new_G594_;
  assign new_G720_ = ~new_G602_;
  assign new_G721_ = ~new_G598_;
  assign new_G722_ = ~new_G609_;
  assign new_G723_ = ~new_G616_;
  assign new_G724_ = ~new_G624_;
  assign new_G725_ = ~new_G701_ | ~new_G702_;
  assign new_G726_ = ~new_G632_;
  assign new_G727_ = ~new_G632_ | ~new_G539_;
  assign new_G728_ = ~new_G645_;
  assign new_G729_ = ~new_G703_ | ~new_G704_;
  assign new_G730_ = ~new_G546_;
  assign new_G731_ = ~new_G546_;
  assign new_G734_ = ~new_G550_;
  assign new_G735_ = ~new_G550_;
  assign new_G738_ = ~new_G568_ | ~new_G570_;
  assign new_G755_ = ~new_G569_ | ~new_G570_;
  assign new_G772_ = ~new_G657_;
  assign new_G773_ = ~new_G657_ | ~new_G585_;
  assign new_G774_ = ~new_G660_;
  assign new_G775_ = ~new_G660_ | ~new_G589_;
  assign new_G776_ = ~new_G663_;
  assign new_G777_ = ~new_G663_ | ~new_G593_;
  assign new_G778_ = ~new_G666_;
  assign new_G779_ = ~new_G666_ | ~new_G597_;
  assign new_G780_ = ~new_G669_;
  assign new_G781_ = ~new_G669_ | ~new_G601_;
  assign new_G782_ = ~new_G672_;
  assign new_G783_ = ~new_G672_ | ~new_G605_;
  assign new_G784_ = ~new_G675_;
  assign new_G785_ = ~new_G606_;
  assign new_G786_ = ~new_G678_;
  assign new_G787_ = ~new_G681_;
  assign new_G788_ = ~new_G681_ | ~new_G615_;
  assign new_G789_ = ~new_G612_;
  assign new_G790_ = ~new_G684_;
  assign new_G791_ = ~new_G684_ | ~new_G619_;
  assign new_G792_ = ~new_G687_;
  assign new_G793_ = ~new_G687_ | ~new_G623_;
  assign new_G794_ = ~new_G620_;
  assign new_G795_ = ~new_G690_;
  assign new_G796_ = ~new_G690_ | ~new_G627_;
  assign new_G797_ = ~new_G628_;
  assign new_G798_ = ~new_G628_ | ~new_G631_;
  assign new_G799_ = ~new_G705_ | ~new_G706_;
  assign new_G802_ = ~new_G707_ | ~new_G708_;
  assign new_G805_ = ~new_G693_;
  assign new_G806_ = ~new_G693_ | ~new_G644_;
  assign new_G807_ = ~new_G641_;
  assign new_G808_ = ~new_G696_;
  assign new_G809_ = ~new_G696_ | ~new_G648_;
  assign new_G810_ = ~new_G709_ | ~new_G710_;
  assign new_G813_ = ~new_G711_ | ~new_G712_;
  assign new_G816_ = ~new_G713_ | ~new_G714_;
  assign new_G819_ = ~new_G554_;
  assign new_G822_ = ~new_G554_;
  assign new_G825_ = ~new_G557_;
  assign new_G828_ = ~new_G557_;
  assign new_G831_ = ~new_G717_;
  assign new_G834_ = ~new_G410_ | ~new_G726_;
  assign new_G835_ = ~new_G467_ | ~new_G772_;
  assign new_G836_ = ~new_G470_ | ~new_G774_;
  assign new_G837_ = ~new_G473_ | ~new_G776_;
  assign new_G838_ = ~new_G476_ | ~new_G778_;
  assign new_G839_ = ~new_G479_ | ~new_G780_;
  assign new_G840_ = ~new_G482_ | ~new_G782_;
  assign new_G841_ = ~new_G485_ | ~new_G787_;
  assign new_G842_ = ~new_G488_ | ~new_G790_;
  assign new_G843_ = ~new_G491_ | ~new_G792_;
  assign new_G844_ = ~new_G494_ | ~new_G795_;
  assign new_G845_ = ~new_G725_;
  assign new_G848_ = ~new_G407_ | ~new_G797_;
  assign new_G849_ = ~new_G509_ | ~new_G805_;
  assign new_G850_ = ~new_G512_ | ~new_G808_;
  assign new_G851_ = ~new_G729_;
  assign new_G854_ = ~new_G834_ | ~new_G727_;
  assign new_G855_ = ~new_G816_ | ~new_G541_;
  assign new_G856_ = ~new_G816_;
  assign new_G857_ = ~new_G822_;
  assign new_G858_ = ~new_G819_;
  assign new_G859_ = ~new_G828_;
  assign new_G860_ = ~new_G825_;
  assign new_G861_ = ~new_G835_ | ~new_G773_;
  assign new_G864_ = ~new_G836_ | ~new_G775_;
  assign new_G867_ = ~new_G837_ | ~new_G777_;
  assign new_G870_ = ~new_G838_ | ~new_G779_;
  assign new_G873_ = ~new_G839_ | ~new_G781_;
  assign new_G876_ = ~new_G840_ | ~new_G783_;
  assign new_G879_ = ~new_G841_ | ~new_G788_;
  assign new_G882_ = ~new_G842_ | ~new_G791_;
  assign new_G885_ = ~new_G843_ | ~new_G793_;
  assign new_G888_ = ~new_G844_ | ~new_G796_;
  assign new_G891_ = ~new_G848_ | ~new_G798_;
  assign new_G894_ = ~new_G799_;
  assign new_G895_ = ~new_G799_ | ~new_G637_;
  assign new_G896_ = ~new_G802_;
  assign new_G897_ = ~new_G802_ | ~new_G640_;
  assign new_G898_ = ~new_G849_ | ~new_G806_;
  assign new_G901_ = ~new_G850_ | ~new_G809_;
  assign new_G904_ = ~new_G810_;
  assign new_G905_ = ~new_G810_ | ~new_G651_;
  assign new_G906_ = ~new_G813_;
  assign new_G907_ = ~new_G813_ | ~new_G654_;
  assign new_G908_ = ~new_G845_;
  assign new_G909_ = ~new_G428_ | ~new_G856_;
  assign new_G910_ = ~new_G851_;
  assign new_G911_ = ~new_G831_;
  assign new_G914_ = ~new_G831_;
  assign new_G917_ = ~new_G413_ | ~new_G894_;
  assign new_G918_ = ~new_G416_ | ~new_G896_;
  assign new_G919_ = ~new_G419_ | ~new_G904_;
  assign new_G920_ = ~new_G425_ | ~new_G906_;
  assign new_G921_ = ~new_G854_;
  assign new_G924_ = ~new_G864_ | ~new_G715_;
  assign new_G925_ = ~new_G864_;
  assign new_G926_ = ~new_G861_ | ~new_G716_;
  assign new_G927_ = ~new_G861_;
  assign new_G928_ = ~new_G867_ | ~new_G718_;
  assign new_G929_ = ~new_G867_;
  assign new_G930_ = ~new_G870_ | ~new_G719_;
  assign new_G931_ = ~new_G870_;
  assign new_G932_ = ~new_G876_ | ~new_G720_;
  assign new_G933_ = ~new_G876_;
  assign new_G934_ = ~new_G873_ | ~new_G721_;
  assign new_G935_ = ~new_G873_;
  assign new_G936_ = ~new_G882_ | ~new_G723_;
  assign new_G937_ = ~new_G882_;
  assign new_G938_ = ~new_G888_ | ~new_G724_;
  assign new_G939_ = ~new_G888_;
  assign new_G940_ = ~new_G891_;
  assign new_G941_ = ~new_G901_ | ~new_G728_;
  assign new_G942_ = ~new_G901_;
  assign new_G943_ = ~new_G855_ | ~new_G909_;
  assign new_G944_ = ~new_G879_;
  assign new_G945_ = ~new_G879_ | ~new_G789_;
  assign new_G946_ = ~new_G885_;
  assign new_G947_ = ~new_G885_ | ~new_G794_;
  assign new_G948_ = ~new_G895_ | ~new_G917_;
  assign new_G951_ = ~new_G898_;
  assign new_G952_ = ~new_G898_ | ~new_G807_;
  assign new_G953_ = ~new_G897_ | ~new_G918_;
  assign new_G956_ = ~new_G907_ | ~new_G920_;
  assign new_G959_ = ~new_G905_ | ~new_G919_;
  assign new_G962_ = ~new_G586_ | ~new_G925_;
  assign new_G963_ = ~new_G582_ | ~new_G927_;
  assign new_G964_ = ~new_G590_ | ~new_G929_;
  assign new_G965_ = ~new_G914_;
  assign new_G966_ = ~new_G911_;
  assign new_G967_ = ~new_G594_ | ~new_G931_;
  assign new_G968_ = ~new_G602_ | ~new_G933_;
  assign new_G969_ = ~new_G598_ | ~new_G935_;
  assign new_G970_ = ~new_G616_ | ~new_G937_;
  assign new_G971_ = ~new_G624_ | ~new_G939_;
  assign new_G972_ = ~new_G645_ | ~new_G942_;
  assign new_G973_ = ~new_G921_;
  assign new_G974_ = ~new_G612_ | ~new_G944_;
  assign new_G975_ = ~new_G620_ | ~new_G946_;
  assign new_G976_ = ~new_G641_ | ~new_G951_;
  assign new_G977_ = ~new_G943_;
  assign new_G980_ = ~new_G924_ | ~new_G962_;
  assign new_G981_ = ~new_G926_ | ~new_G963_;
  assign new_G984_ = ~new_G928_ | ~new_G964_;
  assign new_G987_ = ~new_G930_ | ~new_G967_;
  assign new_G988_ = ~new_G932_ | ~new_G968_;
  assign new_G989_ = ~new_G934_ | ~new_G969_;
  assign new_G993_ = ~new_G936_ | ~new_G970_;
  assign new_G994_ = ~new_G938_ | ~new_G971_;
  assign new_G995_ = ~new_G948_;
  assign new_G996_ = ~new_G941_ | ~new_G972_;
  assign new_G997_ = ~new_G953_;
  assign new_G998_ = ~new_G956_;
  assign new_G999_ = ~new_G959_;
  assign new_G1000_ = ~new_G947_ | ~new_G975_;
  assign new_G1003_ = ~new_G945_ | ~new_G974_;
  assign new_G1006_ = ~new_G952_ | ~new_G976_;
  assign new_G1009_ = ~new_G980_;
  assign new_G1012_ = ~new_G988_;
  assign new_G1015_ = ~new_G993_;
  assign new_G1019_ = ~new_G987_;
  assign new_G1022_ = ~new_G959_ | ~new_G998_;
  assign new_G1023_ = ~new_G956_ | ~new_G999_;
  assign new_G1024_ = ~new_G977_;
  assign new_G1025_ = ~new_G994_;
  assign new_G1028_ = ~new_G996_;
  assign new_G1031_ = ~new_G989_;
  assign new_G1034_ = ~new_G1000_;
  assign new_G1035_ = ~new_G1003_;
  assign new_G1036_ = ~new_G1006_ | ~new_G997_;
  assign new_G1037_ = ~new_G1006_;
  assign new_G1038_ = ~new_G1022_ | ~new_G1023_;
  assign new_G1041_ = ~new_G984_;
  assign new_G1044_ = ~new_G984_;
  assign new_G1047_ = ~new_G989_;
  assign new_G1050_ = ~new_G989_;
  assign new_G1053_ = ~new_G981_;
  assign new_G1056_ = ~new_G981_;
  assign new_G1059_ = ~new_G1015_;
  assign new_G1062_ = ~new_G1012_;
  assign new_G1065_ = ~new_G1025_;
  assign new_G1066_ = ~new_G953_ | ~new_G1037_;
  assign new_G1067_ = ~new_G1028_ | ~new_G1024_;
  assign new_G1068_ = ~new_G1028_;
  assign new_G1069_ = ~new_G1019_;
  assign new_G1072_ = ~new_G1019_;
  assign new_G1075_ = ~new_G1009_;
  assign new_G1078_ = ~new_G1009_;
  assign new_G1081_ = ~new_G1012_;
  assign new_G1084_ = ~new_G1015_;
  assign new_G1087_ = ~new_G1015_;
  assign new_G1090_ = ~new_G1038_ | ~new_G540_;
  assign new_G1091_ = ~new_G1038_;
  assign new_G1092_ = ~new_G1041_;
  assign new_G1093_ = ~new_G1044_;
  assign new_G1094_ = ~new_G1047_ | ~new_G784_;
  assign new_G1095_ = ~new_G1047_;
  assign new_G1096_ = ~new_G1050_ | ~new_G786_;
  assign new_G1097_ = ~new_G1050_;
  assign new_G1098_ = ~new_G1053_;
  assign new_G1099_ = ~new_G1056_;
  assign new_G1100_ = ~new_G1036_ | ~new_G1066_;
  assign new_G1103_ = ~new_G977_ | ~new_G1068_;
  assign new_G1104_ = ~new_G1031_;
  assign new_G1107_ = ~new_G1031_;
  assign new_G1110_ = ~new_G422_ | ~new_G1091_;
  assign new_G1111_ = ~new_G1072_;
  assign new_G1112_ = ~new_G1075_ | ~new_G1092_;
  assign new_G1113_ = ~new_G1075_;
  assign new_G1114_ = ~new_G1078_ | ~new_G1093_;
  assign new_G1115_ = ~new_G1078_;
  assign new_G1116_ = ~new_G675_ | ~new_G1095_;
  assign new_G1117_ = ~new_G678_ | ~new_G1097_;
  assign new_G1118_ = ~new_G1059_;
  assign new_G1121_ = ~new_G1059_;
  assign new_G1124_ = ~new_G1081_ | ~new_G1035_;
  assign new_G1125_ = ~new_G1081_;
  assign new_G1126_ = ~new_G1067_ | ~new_G1103_;
  assign new_G1129_ = ~new_G1084_;
  assign new_G1130_ = ~new_G1069_;
  assign new_G1131_ = ~new_G1087_;
  assign new_G1132_ = ~new_G1062_;
  assign new_G1135_ = ~new_G1062_;
  assign new_G1138_ = ~new_G1100_ | ~new_G995_;
  assign new_G1139_ = ~new_G1100_;
  assign new_G1140_ = ~new_G1090_ | ~new_G1110_;
  assign new_G1143_ = ~new_G1041_ | ~new_G1113_;
  assign new_G1144_ = ~new_G1044_ | ~new_G1115_;
  assign new_G1145_ = ~new_G1094_ | ~new_G1116_;
  assign new_G1148_ = ~new_G1096_ | ~new_G1117_;
  assign new_G1151_ = ~new_G1003_ | ~new_G1125_;
  assign new_G1152_ = ~new_G1104_;
  assign new_G1153_ = ~new_G1104_ | ~new_G1129_;
  assign new_G1154_ = ~new_G1107_;
  assign new_G1155_ = ~new_G1107_ | ~new_G1131_;
  assign new_G1156_ = ~new_G1121_;
  assign new_G1157_ = ~new_G948_ | ~new_G1139_;
  assign new_G1158_ = ~new_G1126_ | ~new_G910_;
  assign new_G1159_ = ~new_G1126_;
  assign new_G1160_ = ~new_G1112_ | ~new_G1143_;
  assign new_G1163_ = ~new_G1114_ | ~new_G1144_;
  assign new_G1166_ = ~new_G1132_;
  assign new_G1167_ = ~new_G1132_ | ~new_G1098_;
  assign new_G1168_ = ~new_G1118_;
  assign new_G1169_ = ~new_G1135_;
  assign new_G1170_ = ~new_G1135_ | ~new_G1099_;
  assign new_G1171_ = ~new_G1124_ | ~new_G1151_;
  assign new_G1174_ = ~new_G1084_ | ~new_G1152_;
  assign new_G1175_ = ~new_G1087_ | ~new_G1154_;
  assign new_G1176_ = ~new_G1148_ | ~new_G722_;
  assign new_G1177_ = ~new_G1148_;
  assign new_G1178_ = ~new_G1138_ | ~new_G1157_;
  assign new_G1181_ = ~new_G851_ | ~new_G1159_;
  assign new_G1182_ = ~new_G1140_ | ~new_G212_;
  assign new_G1185_ = ~new_G1145_;
  assign new_G1186_ = ~new_G1145_ | ~new_G785_;
  assign new_G1187_ = ~new_G1053_ | ~new_G1166_;
  assign new_G1188_ = ~new_G1056_ | ~new_G1169_;
  assign new_G1189_ = ~new_G1174_ | ~new_G1153_;
  assign new_G1192_ = ~new_G1175_ | ~new_G1155_;
  assign new_G1195_ = ~new_G1140_;
  assign new_G1198_ = ~new_G1163_ | ~new_G965_;
  assign new_G1199_ = ~new_G1163_;
  assign new_G1200_ = ~new_G1160_ | ~new_G966_;
  assign new_G1201_ = ~new_G1160_;
  assign new_G1202_ = ~new_G609_ | ~new_G1177_;
  assign new_G1203_ = ~new_G1171_ | ~new_G908_;
  assign new_G1204_ = ~new_G1171_;
  assign new_G1205_ = ~new_G1158_ | ~new_G1181_;
  assign new_G1208_ = ~new_G606_ | ~new_G1185_;
  assign new_G1209_ = ~new_G1187_ | ~new_G1167_;
  assign new_G1212_ = ~new_G1188_ | ~new_G1170_;
  assign new_G1215_ = ~new_G914_ | ~new_G1199_;
  assign new_G1216_ = ~new_G911_ | ~new_G1201_;
  assign new_G1217_ = ~new_G1176_ | ~new_G1202_;
  assign new_G1218_ = ~new_G845_ | ~new_G1204_;
  assign new_G1219_ = ~new_G1192_ | ~new_G1111_;
  assign new_G1220_ = ~new_G1192_;
  assign new_G1221_ = ~new_G1195_;
  assign new_G1222_ = ~new_G1178_ | ~new_G212_;
  assign new_G1225_ = ~new_G1189_;
  assign new_G1226_ = ~new_G1189_ | ~new_G1130_;
  assign new_G1227_ = ~new_G1178_;
  assign new_G1230_ = ~new_G1182_;
  assign new_G1233_ = ~new_G1182_;
  assign new_G1236_ = ~new_G1186_ | ~new_G1208_;
  assign new_G1239_ = ~new_G1198_ | ~new_G1215_;
  assign new_G1240_ = ~new_G1200_ | ~new_G1216_;
  assign new_G1243_ = ~new_G1212_ | ~new_G1156_;
  assign new_G1244_ = ~new_G1212_;
  assign new_G1245_ = ~new_G1203_ | ~new_G1218_;
  assign new_G1246_ = ~new_G1072_ | ~new_G1220_;
  assign new_G1247_ = ~new_G1205_ | ~new_G212_;
  assign new_G1250_ = ~new_G1209_;
  assign new_G1251_ = ~new_G1209_ | ~new_G1168_;
  assign new_G1252_ = ~new_G1069_ | ~new_G1225_;
  assign new_G1253_ = ~new_G1217_;
  assign new_G1256_ = ~new_G1205_;
  assign new_G1259_ = ~new_G1239_;
  assign new_G1260_ = ~new_G1121_ | ~new_G1244_;
  assign new_G1261_ = ~new_G1245_;
  assign new_G1262_ = ~new_G1219_ | ~new_G1246_;
  assign new_G1263_ = ~new_G1227_;
  assign new_G1264_ = ~new_G1233_ | ~new_G566_;
  assign new_G1265_ = ~new_G1233_;
  assign new_G1266_ = ~new_G1230_ | ~new_G567_;
  assign new_G1267_ = ~new_G1230_;
  assign new_G1268_ = ~new_G1236_;
  assign new_G1269_ = ~new_G1118_ | ~new_G1250_;
  assign new_G1270_ = ~new_G1222_;
  assign new_G1273_ = ~new_G1222_;
  assign new_G1276_ = ~new_G1226_ | ~new_G1252_;
  assign new_G1279_ = ~new_G1243_ | ~new_G1260_;
  assign new_G1280_ = ~new_G1253_;
  assign new_G1281_ = ~new_G1256_;
  assign new_G1282_ = ~new_G458_ | ~new_G1265_;
  assign new_G1283_ = ~new_G455_ | ~new_G1267_;
  assign new_G1284_ = ~new_G1240_;
  assign new_G1287_ = ~new_G1262_;
  assign new_G1290_ = ~new_G1247_;
  assign new_G1293_ = ~new_G1247_;
  assign new_G1296_ = ~new_G1240_;
  assign new_G1299_ = ~new_G1251_ | ~new_G1269_;
  assign new_G1302_ = new_G1259_ & new_G380_;
  assign new_G1305_ = new_G381_ & new_G1261_;
  assign new_G1308_ = ~new_G1273_ | ~new_G564_;
  assign new_G1309_ = ~new_G1273_;
  assign new_G1310_ = ~new_G1270_ | ~new_G565_;
  assign new_G1311_ = ~new_G1270_;
  assign new_G1312_ = ~new_G1264_ | ~new_G1282_;
  assign new_G1313_ = ~new_G1266_ | ~new_G1283_;
  assign new_G1316_ = ~new_G1276_;
  assign new_G1317_ = ~new_G1279_;
  assign new_G1320_ = ~new_G1284_;
  assign new_G1321_ = ~new_G1284_ | ~new_G1280_;
  assign new_G1322_ = ~new_G1287_;
  assign new_G1323_ = ~new_G1287_ | ~new_G973_;
  assign new_G1324_ = ~new_G1293_ | ~new_G859_;
  assign new_G1325_ = ~new_G1293_;
  assign new_G1326_ = ~new_G1290_ | ~new_G860_;
  assign new_G1327_ = ~new_G1290_;
  assign new_G1328_ = ~new_G452_ | ~new_G1309_;
  assign new_G1329_ = ~new_G449_ | ~new_G1311_;
  assign new_G1330_ = ~new_G1312_;
  assign new_G1331_ = ~new_G1296_;
  assign new_G1332_ = ~new_G1296_ | ~new_G1268_;
  assign new_G1333_ = ~new_G1299_;
  assign new_G1334_ = ~new_G1299_ | ~new_G1065_;
  assign new_G1335_ = ~new_G1302_;
  assign new_G1336_ = ~new_G1305_;
  assign new_G1337_ = ~new_G1253_ | ~new_G1320_;
  assign new_G1338_ = ~new_G1317_;
  assign new_G1339_ = ~new_G1317_ | ~new_G1034_;
  assign new_G1340_ = ~new_G921_ | ~new_G1322_;
  assign new_G1341_ = ~new_G828_ | ~new_G1325_;
  assign new_G1342_ = ~new_G825_ | ~new_G1327_;
  assign new_G1343_ = ~new_G1308_ | ~new_G1328_;
  assign new_G1344_ = ~new_G1310_ | ~new_G1329_;
  assign new_G1347_ = ~new_G1313_;
  assign new_G1350_ = ~new_G1313_;
  assign new_G1353_ = ~new_G1236_ | ~new_G1331_;
  assign new_G1354_ = ~new_G1025_ | ~new_G1333_;
  assign new_G1355_ = ~new_G1337_ | ~new_G1321_;
  assign new_G1356_ = ~new_G1000_ | ~new_G1338_;
  assign new_G1357_ = ~new_G1340_ | ~new_G1323_;
  assign new_G1358_ = ~new_G1324_ | ~new_G1341_;
  assign new_G1359_ = ~new_G1326_ | ~new_G1342_;
  assign new_G1362_ = ~new_G1343_;
  assign new_G1363_ = ~new_G1353_ | ~new_G1332_;
  assign new_G1366_ = ~new_G1354_ | ~new_G1334_;
  assign new_G1369_ = ~new_G1355_;
  assign new_G1370_ = ~new_G1356_ | ~new_G1339_;
  assign new_G1371_ = ~new_G1357_ | ~new_G212_;
  assign new_G1374_ = ~new_G1358_;
  assign new_G1375_ = ~new_G1344_;
  assign new_G1378_ = ~new_G1344_;
  assign new_G1381_ = ~new_G1363_;
  assign new_G1382_ = ~new_G1366_;
  assign new_G1383_ = ~new_G1369_ | ~new_G212_;
  assign new_G1386_ = ~new_G1370_ | ~new_G212_;
  assign new_G1389_ = ~new_G1359_;
  assign new_G1392_ = ~new_G1359_;
  assign new_G1395_ = new_G1347_ & new_G1375_;
  assign new_G1410_ = new_G1350_ & new_G1375_;
  assign new_G1420_ = new_G1347_ & new_G1378_;
  assign new_G1434_ = new_G1350_ & new_G1378_;
  assign new_G1439_ = ~new_G1371_;
  assign new_G1442_ = ~new_G1371_;
  assign new_G1445_ = ~new_G1383_;
  assign new_G1448_ = ~new_G1383_;
  assign new_G1451_ = ~new_G1386_;
  assign new_G1454_ = ~new_G1386_;
  assign new_G1457_ = ~new_G1442_ | ~new_G562_;
  assign new_G1458_ = ~new_G1442_;
  assign new_G1459_ = ~new_G1439_ | ~new_G563_;
  assign new_G1460_ = ~new_G1439_;
  assign new_G1461_ = ~new_G1448_ | ~new_G857_;
  assign new_G1462_ = ~new_G1448_;
  assign new_G1463_ = ~new_G1445_ | ~new_G858_;
  assign new_G1464_ = ~new_G1445_;
  assign new_G1465_ = ~new_G1454_ | ~new_G560_;
  assign new_G1466_ = ~new_G1454_;
  assign new_G1467_ = ~new_G1451_ | ~new_G561_;
  assign new_G1468_ = ~new_G1451_;
  assign new_G1469_ = ~new_G446_ | ~new_G1458_;
  assign new_G1470_ = ~new_G443_ | ~new_G1460_;
  assign new_G1471_ = ~new_G822_ | ~new_G1462_;
  assign new_G1472_ = ~new_G819_ | ~new_G1464_;
  assign new_G1473_ = ~new_G440_ | ~new_G1466_;
  assign new_G1474_ = ~new_G437_ | ~new_G1468_;
  assign new_G1475_ = ~new_G1457_ | ~new_G1469_;
  assign new_G1476_ = ~new_G1459_ | ~new_G1470_;
  assign new_G1479_ = ~new_G1461_ | ~new_G1471_;
  assign new_G1480_ = ~new_G1463_ | ~new_G1472_;
  assign new_G1483_ = ~new_G1465_ | ~new_G1473_;
  assign new_G1484_ = ~new_G1467_ | ~new_G1474_;
  assign new_G1487_ = ~new_G1475_;
  assign new_G1488_ = ~new_G1479_;
  assign new_G1489_ = ~new_G1483_;
  assign new_G1490_ = ~new_G1476_;
  assign new_G1493_ = ~new_G1476_;
  assign new_G1496_ = ~new_G1480_;
  assign new_G1499_ = new_G731_ & new_G1480_;
  assign new_G1502_ = ~new_G1484_;
  assign new_G1505_ = new_G735_ & new_G1484_;
  assign new_G1508_ = ~new_G550_ | ~new_G1488_ | ~new_G1489_ | ~new_G1374_ | ~new_G1330_ | ~new_G1362_ | ~new_G1487_ | ~new_G546_;
  assign new_G1511_ = ~new_G1499_;
  assign new_G1522_ = ~new_G1499_;
  assign new_G1538_ = ~new_G1505_;
  assign new_G1549_ = ~new_G1505_;
  assign new_G1563_ = new_G1389_ & new_G1490_;
  assign new_G1576_ = new_G1392_ & new_G1490_;
  assign new_G1584_ = new_G1389_ & new_G1493_;
  assign new_G1598_ = new_G1392_ & new_G1493_;
  assign new_G1607_ = new_G260_ & new_G1508_ & new_G235_ & new_G235_;
  assign new_G1608_ = new_G730_ & new_G1496_;
  assign new_G1609_ = new_G731_ & new_G1496_;
  assign new_G1624_ = new_G734_ & new_G1502_;
  assign new_G1625_ = new_G735_ & new_G1502_;
  assign new_G1642_ = ~new_G1511_ | ~new_G1538_ | ~new_G1584_ | ~new_G1395_ | ~new_G738_;
  assign new_G1645_ = ~new_G1511_ | ~new_G1538_ | ~new_G1563_ | ~new_G1420_ | ~new_G738_;
  assign new_G1648_ = ~new_G1511_ | ~new_G1538_ | ~new_G1563_ | ~new_G1410_ | ~new_G738_;
  assign new_G1651_ = ~new_G1511_ | ~new_G1538_ | ~new_G1576_ | ~new_G1395_ | ~new_G738_;
  assign new_G1654_ = ~new_G1522_ | ~new_G1538_ | ~new_G1598_ | ~new_G1410_ | ~new_G755_;
  assign new_G1657_ = ~new_G1522_ | ~new_G1549_ | ~new_G1584_ | ~new_G1434_ | ~new_G755_;
  assign new_G1660_ = ~new_G1522_ | ~new_G1549_ | ~new_G1598_ | ~new_G1420_ | ~new_G755_;
  assign new_G1663_ = new_G1511_ & new_G1538_ & new_G1584_ & new_G1395_ & new_G738_;
  assign new_G1666_ = new_G1511_ & new_G1538_ & new_G1563_ & new_G1420_ & new_G738_;
  assign new_G1669_ = new_G1511_ & new_G1538_ & new_G1563_ & new_G1410_ & new_G738_;
  assign new_G1672_ = new_G1511_ & new_G1538_ & new_G1576_ & new_G1395_ & new_G738_;
  assign new_G1675_ = new_G1522_ & new_G1538_ & new_G1598_ & new_G1410_ & new_G755_;
  assign new_G1678_ = new_G1522_ & new_G1549_ & new_G1584_ & new_G1434_ & new_G755_;
  assign new_G1681_ = new_G1522_ & new_G1549_ & new_G1598_ & new_G1420_ & new_G755_;
  assign new_G1684_ = ~new_G1511_ | ~new_G1625_ | ~new_G1584_ | ~new_G1420_ | ~new_G738_;
  assign new_G1687_ = ~new_G1522_ | ~new_G1625_ | ~new_G1584_ | ~new_G1410_ | ~new_G738_;
  assign new_G1690_ = ~new_G1522_ | ~new_G1625_ | ~new_G1598_ | ~new_G1395_ | ~new_G738_;
  assign new_G1693_ = ~new_G1522_ | ~new_G1625_ | ~new_G1563_ | ~new_G1434_ | ~new_G738_;
  assign new_G1696_ = ~new_G1522_ | ~new_G1625_ | ~new_G1576_ | ~new_G1420_ | ~new_G755_;
  assign new_G1699_ = ~new_G1609_ | ~new_G1549_ | ~new_G1584_ | ~new_G1420_ | ~new_G755_;
  assign new_G1702_ = ~new_G1609_ | ~new_G1549_ | ~new_G1584_ | ~new_G1410_ | ~new_G755_;
  assign new_G1705_ = ~new_G1609_ | ~new_G1549_ | ~new_G1598_ | ~new_G1395_ | ~new_G755_;
  assign new_G1708_ = ~new_G1609_ | ~new_G1549_ | ~new_G1576_ | ~new_G1420_ | ~new_G755_;
  assign new_G1711_ = ~new_G1522_ | ~new_G1625_ | ~new_G1563_ | ~new_G1395_ | ~new_G573_;
  assign new_G1712_ = ~new_G1609_ | ~new_G1549_ | ~new_G1563_ | ~new_G1395_ | ~new_G573_;
  assign new_G1713_ = ~new_G1609_ | ~new_G1625_ | ~new_G1584_ | ~new_G1395_ | ~new_G573_;
  assign new_G1714_ = ~new_G1609_ | ~new_G1625_ | ~new_G1563_ | ~new_G1420_ | ~new_G573_;
  assign new_G1715_ = ~new_G1609_ | ~new_G1625_ | ~new_G1563_ | ~new_G1410_ | ~new_G573_;
  assign new_G1716_ = ~new_G1609_ | ~new_G1625_ | ~new_G1576_ | ~new_G1395_ | ~new_G573_;
  assign new_G1717_ = ~new_G1609_ | ~new_G1624_ | ~new_G1563_ | ~new_G1395_ | ~new_G573_;
  assign new_G1718_ = ~new_G1608_ | ~new_G1625_ | ~new_G1563_ | ~new_G1395_ | ~new_G573_;
  assign new_G1719_ = new_G1511_ & new_G1625_ & new_G1584_ & new_G1420_ & new_G738_;
  assign new_G1722_ = new_G1522_ & new_G1625_ & new_G1584_ & new_G1410_ & new_G738_;
  assign new_G1725_ = new_G1522_ & new_G1625_ & new_G1598_ & new_G1395_ & new_G738_;
  assign new_G1728_ = new_G1522_ & new_G1625_ & new_G1563_ & new_G1434_ & new_G738_;
  assign new_G1731_ = new_G1522_ & new_G1625_ & new_G1576_ & new_G1420_ & new_G755_;
  assign new_G1734_ = new_G1609_ & new_G1549_ & new_G1584_ & new_G1420_ & new_G755_;
  assign new_G1737_ = new_G1609_ & new_G1549_ & new_G1584_ & new_G1410_ & new_G755_;
  assign new_G1740_ = new_G1609_ & new_G1549_ & new_G1598_ & new_G1395_ & new_G755_;
  assign new_G1743_ = new_G1609_ & new_G1549_ & new_G1576_ & new_G1420_ & new_G755_;
  assign new_G1746_ = ~new_G1663_ | ~new_G313_;
  assign new_G1747_ = ~new_G1663_;
  assign new_G1748_ = ~new_G1666_ | ~new_G314_;
  assign new_G1749_ = ~new_G1666_;
  assign new_G1750_ = ~new_G1669_ | ~new_G315_;
  assign new_G1751_ = ~new_G1669_;
  assign new_G1752_ = ~new_G1672_ | ~new_G316_;
  assign new_G1753_ = ~new_G1672_;
  assign new_G1754_ = ~new_G1675_ | ~new_G322_;
  assign new_G1755_ = ~new_G1675_;
  assign new_G1756_ = ~new_G1678_ | ~new_G327_;
  assign new_G1757_ = ~new_G1678_;
  assign new_G1758_ = ~new_G1681_ | ~new_G328_;
  assign new_G1759_ = ~new_G1681_;
  assign new_G1760_ = new_G1718_ & new_G1717_ & new_G1716_ & new_G1711_ & new_G1712_ & new_G1713_ & new_G1714_ & new_G1715_;
  assign new_G1761_ = ~new_G265_ | ~new_G1747_;
  assign new_G1762_ = ~new_G268_ | ~new_G1749_;
  assign new_G1763_ = ~new_G271_ | ~new_G1751_;
  assign new_G1764_ = ~new_G274_ | ~new_G1753_;
  assign new_G1765_ = ~new_G1719_ | ~new_G317_;
  assign new_G1766_ = ~new_G1719_;
  assign new_G1767_ = ~new_G1722_ | ~new_G318_;
  assign new_G1768_ = ~new_G1722_;
  assign new_G1769_ = ~new_G1725_ | ~new_G319_;
  assign new_G1770_ = ~new_G1725_;
  assign new_G1771_ = ~new_G1728_ | ~new_G320_;
  assign new_G1772_ = ~new_G1728_;
  assign new_G1773_ = ~new_G1731_ | ~new_G321_;
  assign new_G1774_ = ~new_G1731_;
  assign new_G1775_ = ~new_G292_ | ~new_G1755_;
  assign new_G1776_ = ~new_G1734_ | ~new_G323_;
  assign new_G1777_ = ~new_G1734_;
  assign new_G1778_ = ~new_G1737_ | ~new_G324_;
  assign new_G1779_ = ~new_G1737_;
  assign new_G1780_ = ~new_G1740_ | ~new_G325_;
  assign new_G1781_ = ~new_G1740_;
  assign new_G1782_ = ~new_G1743_ | ~new_G326_;
  assign new_G1783_ = ~new_G1743_;
  assign new_G1784_ = ~new_G307_ | ~new_G1757_;
  assign new_G1785_ = ~new_G310_ | ~new_G1759_;
  assign new_G1786_ = ~new_G1693_ | ~new_G1690_ | ~new_G1687_ | ~new_G1642_ | ~new_G1645_ | ~new_G1648_ | ~new_G1651_ | ~new_G1684_;
  assign new_G1787_ = ~new_G1660_ | ~new_G1657_ | ~new_G1708_ | ~new_G1696_ | ~new_G1654_ | ~new_G1699_ | ~new_G1702_ | ~new_G1705_;
  assign new_G1788_ = new_G1693_ & new_G1690_ & new_G1687_ & new_G1642_ & new_G1645_ & new_G1648_ & new_G1651_ & new_G1684_;
  assign new_G1791_ = new_G1660_ & new_G1657_ & new_G1708_ & new_G1696_ & new_G1654_ & new_G1699_ & new_G1702_ & new_G1705_;
  assign new_G1794_ = ~new_G277_ | ~new_G1766_;
  assign new_G1795_ = ~new_G280_ | ~new_G1768_;
  assign new_G1796_ = ~new_G283_ | ~new_G1770_;
  assign new_G1797_ = ~new_G286_ | ~new_G1772_;
  assign new_G1798_ = ~new_G289_ | ~new_G1774_;
  assign new_G1799_ = ~new_G295_ | ~new_G1777_;
  assign new_G1800_ = ~new_G298_ | ~new_G1779_;
  assign new_G1801_ = ~new_G301_ | ~new_G1781_;
  assign new_G1802_ = ~new_G304_ | ~new_G1783_;
  assign new_G1803_ = new_G1786_ & new_G197_;
  assign new_G1806_ = new_G1787_ & new_G198_;
  assign new_G1809_ = new_G1788_ & new_G1791_ & new_G1760_;
  assign new_G1810_ = ~new_G1788_ | ~new_G1791_;
  assign new_G1817_ = new_G260_ & new_G1508_ & n1321_lo & new_G1809_;
  assign new_G1818_ = ~new_G1803_ | ~new_G1335_;
  assign new_G1819_ = ~new_G1803_;
  assign new_G1820_ = ~new_G1806_ | ~new_G1336_;
  assign new_G1821_ = ~new_G1806_;
  assign new_G1822_ = new_G544_ & new_G205_ & new_G1810_;
  assign new_G1825_ = n1237_lo & new_G205_ & new_G1810_;
  assign new_G1828_ = n1261_lo & new_G205_ & new_G1810_;
  assign new_G1831_ = n1273_lo & new_G205_ & new_G1810_;
  assign new_G1834_ = new_G545_ & new_G205_ & new_G1810_;
  assign new_G1837_ = ~new_G1302_ | ~new_G1819_;
  assign new_G1838_ = ~new_G1305_ | ~new_G1821_;
  assign new_G1839_ = n1249_lo & new_G205_ & new_G1810_;
  assign new_G1842_ = ~new_G1818_ | ~new_G1837_;
  assign new_G1845_ = ~new_G1820_ | ~new_G1838_;
  assign new_G1848_ = ~new_G1822_ | ~new_G1381_;
  assign new_G1849_ = ~new_G1825_ | ~new_G1382_;
  assign new_G1850_ = ~new_G1828_ | ~new_G1263_;
  assign new_G1851_ = ~new_G1831_ | ~new_G1221_;
  assign new_G1852_ = ~new_G1834_ | ~new_G1281_;
  assign new_G1853_ = ~new_G1822_;
  assign new_G1854_ = ~new_G1825_;
  assign new_G1855_ = ~new_G1828_;
  assign new_G1856_ = ~new_G1831_;
  assign new_G1857_ = ~new_G1834_;
  assign new_G1858_ = ~new_G1839_;
  assign new_G1859_ = ~new_G1839_ | ~new_G1316_;
  assign new_G1860_ = ~new_G1363_ | ~new_G1853_;
  assign new_G1861_ = ~new_G1366_ | ~new_G1854_;
  assign new_G1862_ = ~new_G1227_ | ~new_G1855_;
  assign new_G1863_ = ~new_G1195_ | ~new_G1856_;
  assign new_G1864_ = ~new_G1256_ | ~new_G1857_;
  assign new_G1865_ = ~new_G1842_ | ~new_G533_;
  assign new_G1866_ = ~new_G1842_;
  assign new_G1867_ = ~new_G1845_ | ~new_G534_;
  assign new_G1868_ = ~new_G1845_;
  assign new_G1869_ = ~new_G1276_ | ~new_G1858_;
  assign new_G1870_ = ~new_G1860_ | ~new_G1848_;
  assign new_G1871_ = ~new_G1861_ | ~new_G1849_;
  assign new_G1872_ = ~new_G1862_ | ~new_G1850_;
  assign new_G1873_ = ~new_G1863_ | ~new_G1851_;
  assign new_G1874_ = ~new_G1864_ | ~new_G1852_;
  assign new_G1875_ = ~new_G461_ | ~new_G1866_;
  assign new_G1876_ = ~new_G464_ | ~new_G1868_;
  assign new_G1877_ = ~new_G1869_ | ~new_G1859_;
  assign new_G1880_ = ~new_G1877_ | ~new_G940_;
  assign new_G1881_ = ~new_G1877_;
  assign new_G1882_ = ~new_G891_ | ~new_G1881_;
  assign new_G1883_ = ~new_G1880_ | ~new_G1882_;
  assign G1884 = ~new_G1746_ | ~new_G1761_;
  assign G1885 = ~new_G1748_ | ~new_G1762_;
  assign G1886 = ~new_G1750_ | ~new_G1763_;
  assign G1887 = ~new_G1752_ | ~new_G1764_;
  assign G1888 = ~new_G1754_ | ~new_G1775_;
  assign G1889 = ~new_G1756_ | ~new_G1784_;
  assign G1890 = ~new_G1758_ | ~new_G1785_;
  assign G1891 = ~new_G1765_ | ~new_G1794_;
  assign G1892 = ~new_G1767_ | ~new_G1795_;
  assign G1893 = ~new_G1769_ | ~new_G1796_;
  assign G1894 = ~new_G1771_ | ~new_G1797_;
  assign G1895 = ~new_G1773_ | ~new_G1798_;
  assign G1896 = ~new_G1776_ | ~new_G1799_;
  assign G1897 = ~new_G1778_ | ~new_G1800_;
  assign G1898 = ~new_G1780_ | ~new_G1801_;
  assign G1899 = ~new_G1782_ | ~new_G1802_;
  assign G1900 = ~new_G1607_ & ~new_G1817_;
  assign G1901 = new_G1870_ & new_G329_;
  assign G1902 = new_G330_ & new_G1871_;
  assign G1903 = new_G332_ & new_G1872_;
  assign G1904 = new_G1873_ & new_G333_;
  assign G1905 = new_G334_ & new_G1874_;
  assign G1906 = ~new_G1865_ | ~new_G1875_;
  assign G1907 = ~new_G1867_ | ~new_G1876_;
  assign G1908 = new_G1883_ & new_G331_;
  assign n940_li = G1;
  assign n943_li = n940_lo;
  assign n946_li = n943_lo;
  assign n949_li = n946_lo;
  assign n952_li = G2;
  assign n955_li = n952_lo;
  assign n958_li = n955_lo;
  assign n961_li = n958_lo;
  assign n964_li = G3;
  assign n967_li = n964_lo;
  assign n970_li = n967_lo;
  assign n973_li = n970_lo;
  assign n976_li = G4;
  assign n979_li = n976_lo;
  assign n982_li = n979_lo;
  assign n985_li = n982_lo;
  assign n988_li = G5;
  assign n991_li = n988_lo;
  assign n994_li = n991_lo;
  assign n997_li = n994_lo;
  assign n1000_li = G6;
  assign n1003_li = n1000_lo;
  assign n1006_li = n1003_lo;
  assign n1009_li = n1006_lo;
  assign n1012_li = G7;
  assign n1015_li = n1012_lo;
  assign n1018_li = n1015_lo;
  assign n1021_li = n1018_lo;
  assign n1024_li = G8;
  assign n1027_li = n1024_lo;
  assign n1030_li = n1027_lo;
  assign n1033_li = n1030_lo;
  assign n1036_li = G9;
  assign n1039_li = n1036_lo;
  assign n1042_li = n1039_lo;
  assign n1045_li = n1042_lo;
  assign n1048_li = G10;
  assign n1051_li = n1048_lo;
  assign n1054_li = n1051_lo;
  assign n1057_li = n1054_lo;
  assign n1060_li = G11;
  assign n1063_li = n1060_lo;
  assign n1066_li = n1063_lo;
  assign n1069_li = n1066_lo;
  assign n1072_li = G12;
  assign n1075_li = n1072_lo;
  assign n1078_li = n1075_lo;
  assign n1081_li = n1078_lo;
  assign n1084_li = G13;
  assign n1087_li = n1084_lo;
  assign n1090_li = n1087_lo;
  assign n1093_li = n1090_lo;
  assign n1096_li = G14;
  assign n1099_li = n1096_lo;
  assign n1102_li = n1099_lo;
  assign n1105_li = n1102_lo;
  assign n1108_li = G15;
  assign n1111_li = n1108_lo;
  assign n1114_li = n1111_lo;
  assign n1117_li = n1114_lo;
  assign n1120_li = G16;
  assign n1123_li = n1120_lo;
  assign n1126_li = n1123_lo;
  assign n1129_li = n1126_lo;
  assign n1132_li = G17;
  assign n1135_li = n1132_lo;
  assign n1138_li = n1135_lo;
  assign n1141_li = n1138_lo;
  assign n1144_li = G18;
  assign n1147_li = n1144_lo;
  assign n1150_li = n1147_lo;
  assign n1153_li = n1150_lo;
  assign n1156_li = G19;
  assign n1159_li = n1156_lo;
  assign n1162_li = n1159_lo;
  assign n1165_li = n1162_lo;
  assign n1168_li = G20;
  assign n1171_li = n1168_lo;
  assign n1174_li = n1171_lo;
  assign n1177_li = n1174_lo;
  assign n1180_li = G21;
  assign n1183_li = n1180_lo;
  assign n1186_li = n1183_lo;
  assign n1189_li = n1186_lo;
  assign n1192_li = G22;
  assign n1195_li = n1192_lo;
  assign n1198_li = n1195_lo;
  assign n1201_li = n1198_lo;
  assign n1204_li = G23;
  assign n1207_li = n1204_lo;
  assign n1210_li = n1207_lo;
  assign n1213_li = n1210_lo;
  assign n1216_li = G24;
  assign n1219_li = n1216_lo;
  assign n1222_li = n1219_lo;
  assign n1225_li = n1222_lo;
  assign n1228_li = G25;
  assign n1231_li = n1228_lo;
  assign n1234_li = n1231_lo;
  assign n1237_li = n1234_lo;
  assign n1240_li = G26;
  assign n1243_li = n1240_lo;
  assign n1246_li = n1243_lo;
  assign n1249_li = n1246_lo;
  assign n1252_li = G27;
  assign n1255_li = n1252_lo;
  assign n1258_li = n1255_lo;
  assign n1261_li = n1258_lo;
  assign n1264_li = G28;
  assign n1267_li = n1264_lo;
  assign n1270_li = n1267_lo;
  assign n1273_li = n1270_lo;
  assign n1276_li = G29;
  assign n1279_li = n1276_lo;
  assign n1282_li = n1279_lo;
  assign n1285_li = n1282_lo;
  assign n1288_li = G30;
  assign n1291_li = n1288_lo;
  assign n1294_li = n1291_lo;
  assign n1297_li = n1294_lo;
  assign n1300_li = G31;
  assign n1303_li = n1300_lo;
  assign n1306_li = n1303_lo;
  assign n1309_li = n1306_lo;
  assign n1312_li = G32;
  assign n1315_li = n1312_lo;
  assign n1318_li = n1315_lo;
  assign n1321_li = n1318_lo;
  assign n1324_li = G33;
  assign n1327_li = n1324_lo;
  assign n1330_li = n1327_lo;
  assign n1333_li = n1330_lo;
  always @ (posedge clock) begin
    n940_lo <= n940_li;
    n943_lo <= n943_li;
    n946_lo <= n946_li;
    n949_lo <= n949_li;
    n952_lo <= n952_li;
    n955_lo <= n955_li;
    n958_lo <= n958_li;
    n961_lo <= n961_li;
    n964_lo <= n964_li;
    n967_lo <= n967_li;
    n970_lo <= n970_li;
    n973_lo <= n973_li;
    n976_lo <= n976_li;
    n979_lo <= n979_li;
    n982_lo <= n982_li;
    n985_lo <= n985_li;
    n988_lo <= n988_li;
    n991_lo <= n991_li;
    n994_lo <= n994_li;
    n997_lo <= n997_li;
    n1000_lo <= n1000_li;
    n1003_lo <= n1003_li;
    n1006_lo <= n1006_li;
    n1009_lo <= n1009_li;
    n1012_lo <= n1012_li;
    n1015_lo <= n1015_li;
    n1018_lo <= n1018_li;
    n1021_lo <= n1021_li;
    n1024_lo <= n1024_li;
    n1027_lo <= n1027_li;
    n1030_lo <= n1030_li;
    n1033_lo <= n1033_li;
    n1036_lo <= n1036_li;
    n1039_lo <= n1039_li;
    n1042_lo <= n1042_li;
    n1045_lo <= n1045_li;
    n1048_lo <= n1048_li;
    n1051_lo <= n1051_li;
    n1054_lo <= n1054_li;
    n1057_lo <= n1057_li;
    n1060_lo <= n1060_li;
    n1063_lo <= n1063_li;
    n1066_lo <= n1066_li;
    n1069_lo <= n1069_li;
    n1072_lo <= n1072_li;
    n1075_lo <= n1075_li;
    n1078_lo <= n1078_li;
    n1081_lo <= n1081_li;
    n1084_lo <= n1084_li;
    n1087_lo <= n1087_li;
    n1090_lo <= n1090_li;
    n1093_lo <= n1093_li;
    n1096_lo <= n1096_li;
    n1099_lo <= n1099_li;
    n1102_lo <= n1102_li;
    n1105_lo <= n1105_li;
    n1108_lo <= n1108_li;
    n1111_lo <= n1111_li;
    n1114_lo <= n1114_li;
    n1117_lo <= n1117_li;
    n1120_lo <= n1120_li;
    n1123_lo <= n1123_li;
    n1126_lo <= n1126_li;
    n1129_lo <= n1129_li;
    n1132_lo <= n1132_li;
    n1135_lo <= n1135_li;
    n1138_lo <= n1138_li;
    n1141_lo <= n1141_li;
    n1144_lo <= n1144_li;
    n1147_lo <= n1147_li;
    n1150_lo <= n1150_li;
    n1153_lo <= n1153_li;
    n1156_lo <= n1156_li;
    n1159_lo <= n1159_li;
    n1162_lo <= n1162_li;
    n1165_lo <= n1165_li;
    n1168_lo <= n1168_li;
    n1171_lo <= n1171_li;
    n1174_lo <= n1174_li;
    n1177_lo <= n1177_li;
    n1180_lo <= n1180_li;
    n1183_lo <= n1183_li;
    n1186_lo <= n1186_li;
    n1189_lo <= n1189_li;
    n1192_lo <= n1192_li;
    n1195_lo <= n1195_li;
    n1198_lo <= n1198_li;
    n1201_lo <= n1201_li;
    n1204_lo <= n1204_li;
    n1207_lo <= n1207_li;
    n1210_lo <= n1210_li;
    n1213_lo <= n1213_li;
    n1216_lo <= n1216_li;
    n1219_lo <= n1219_li;
    n1222_lo <= n1222_li;
    n1225_lo <= n1225_li;
    n1228_lo <= n1228_li;
    n1231_lo <= n1231_li;
    n1234_lo <= n1234_li;
    n1237_lo <= n1237_li;
    n1240_lo <= n1240_li;
    n1243_lo <= n1243_li;
    n1246_lo <= n1246_li;
    n1249_lo <= n1249_li;
    n1252_lo <= n1252_li;
    n1255_lo <= n1255_li;
    n1258_lo <= n1258_li;
    n1261_lo <= n1261_li;
    n1264_lo <= n1264_li;
    n1267_lo <= n1267_li;
    n1270_lo <= n1270_li;
    n1273_lo <= n1273_li;
    n1276_lo <= n1276_li;
    n1279_lo <= n1279_li;
    n1282_lo <= n1282_li;
    n1285_lo <= n1285_li;
    n1288_lo <= n1288_li;
    n1291_lo <= n1291_li;
    n1294_lo <= n1294_li;
    n1297_lo <= n1297_li;
    n1300_lo <= n1300_li;
    n1303_lo <= n1303_li;
    n1306_lo <= n1306_li;
    n1309_lo <= n1309_li;
    n1312_lo <= n1312_li;
    n1315_lo <= n1315_li;
    n1318_lo <= n1318_li;
    n1321_lo <= n1321_li;
    n1324_lo <= n1324_li;
    n1327_lo <= n1327_li;
    n1330_lo <= n1330_li;
    n1333_lo <= n1333_li;
  end
  initial begin
    n940_lo <= 1'b0;
    n943_lo <= 1'b0;
    n946_lo <= 1'b0;
    n949_lo <= 1'b0;
    n952_lo <= 1'b0;
    n955_lo <= 1'b0;
    n958_lo <= 1'b0;
    n961_lo <= 1'b0;
    n964_lo <= 1'b0;
    n967_lo <= 1'b0;
    n970_lo <= 1'b0;
    n973_lo <= 1'b0;
    n976_lo <= 1'b0;
    n979_lo <= 1'b0;
    n982_lo <= 1'b0;
    n985_lo <= 1'b0;
    n988_lo <= 1'b0;
    n991_lo <= 1'b0;
    n994_lo <= 1'b0;
    n997_lo <= 1'b0;
    n1000_lo <= 1'b0;
    n1003_lo <= 1'b0;
    n1006_lo <= 1'b0;
    n1009_lo <= 1'b0;
    n1012_lo <= 1'b0;
    n1015_lo <= 1'b0;
    n1018_lo <= 1'b0;
    n1021_lo <= 1'b0;
    n1024_lo <= 1'b0;
    n1027_lo <= 1'b0;
    n1030_lo <= 1'b0;
    n1033_lo <= 1'b0;
    n1036_lo <= 1'b0;
    n1039_lo <= 1'b0;
    n1042_lo <= 1'b0;
    n1045_lo <= 1'b0;
    n1048_lo <= 1'b0;
    n1051_lo <= 1'b0;
    n1054_lo <= 1'b0;
    n1057_lo <= 1'b0;
    n1060_lo <= 1'b0;
    n1063_lo <= 1'b0;
    n1066_lo <= 1'b0;
    n1069_lo <= 1'b0;
    n1072_lo <= 1'b0;
    n1075_lo <= 1'b0;
    n1078_lo <= 1'b0;
    n1081_lo <= 1'b0;
    n1084_lo <= 1'b0;
    n1087_lo <= 1'b0;
    n1090_lo <= 1'b0;
    n1093_lo <= 1'b0;
    n1096_lo <= 1'b0;
    n1099_lo <= 1'b0;
    n1102_lo <= 1'b0;
    n1105_lo <= 1'b0;
    n1108_lo <= 1'b0;
    n1111_lo <= 1'b0;
    n1114_lo <= 1'b0;
    n1117_lo <= 1'b0;
    n1120_lo <= 1'b0;
    n1123_lo <= 1'b0;
    n1126_lo <= 1'b0;
    n1129_lo <= 1'b0;
    n1132_lo <= 1'b0;
    n1135_lo <= 1'b0;
    n1138_lo <= 1'b0;
    n1141_lo <= 1'b0;
    n1144_lo <= 1'b0;
    n1147_lo <= 1'b0;
    n1150_lo <= 1'b0;
    n1153_lo <= 1'b0;
    n1156_lo <= 1'b0;
    n1159_lo <= 1'b0;
    n1162_lo <= 1'b0;
    n1165_lo <= 1'b0;
    n1168_lo <= 1'b0;
    n1171_lo <= 1'b0;
    n1174_lo <= 1'b0;
    n1177_lo <= 1'b0;
    n1180_lo <= 1'b0;
    n1183_lo <= 1'b0;
    n1186_lo <= 1'b0;
    n1189_lo <= 1'b0;
    n1192_lo <= 1'b0;
    n1195_lo <= 1'b0;
    n1198_lo <= 1'b0;
    n1201_lo <= 1'b0;
    n1204_lo <= 1'b0;
    n1207_lo <= 1'b0;
    n1210_lo <= 1'b0;
    n1213_lo <= 1'b0;
    n1216_lo <= 1'b0;
    n1219_lo <= 1'b0;
    n1222_lo <= 1'b0;
    n1225_lo <= 1'b0;
    n1228_lo <= 1'b0;
    n1231_lo <= 1'b0;
    n1234_lo <= 1'b0;
    n1237_lo <= 1'b0;
    n1240_lo <= 1'b0;
    n1243_lo <= 1'b0;
    n1246_lo <= 1'b0;
    n1249_lo <= 1'b0;
    n1252_lo <= 1'b0;
    n1255_lo <= 1'b0;
    n1258_lo <= 1'b0;
    n1261_lo <= 1'b0;
    n1264_lo <= 1'b0;
    n1267_lo <= 1'b0;
    n1270_lo <= 1'b0;
    n1273_lo <= 1'b0;
    n1276_lo <= 1'b0;
    n1279_lo <= 1'b0;
    n1282_lo <= 1'b0;
    n1285_lo <= 1'b0;
    n1288_lo <= 1'b0;
    n1291_lo <= 1'b0;
    n1294_lo <= 1'b0;
    n1297_lo <= 1'b0;
    n1300_lo <= 1'b0;
    n1303_lo <= 1'b0;
    n1306_lo <= 1'b0;
    n1309_lo <= 1'b0;
    n1312_lo <= 1'b0;
    n1315_lo <= 1'b0;
    n1318_lo <= 1'b0;
    n1321_lo <= 1'b0;
    n1324_lo <= 1'b0;
    n1327_lo <= 1'b0;
    n1330_lo <= 1'b0;
    n1333_lo <= 1'b0;
  end
endmodule


