
module mymod
(
  A_0_,
  A_1_,
  A_2_,
  A_3_,
  A_4_,
  A_5_,
  A_6_,
  A_7_,
  B_0_,
  B_1_,
  B_2_,
  B_3_,
  B_4_,
  B_5_,
  B_6_,
  B_7_,
  SUM_0_,
  SUM_1_,
  SUM_2_,
  SUM_3_,
  SUM_4_,
  SUM_5_,
  SUM_6_,
  SUM_7_
);

  input A_0_;input A_1_;input A_2_;input A_3_;input A_4_;input A_5_;input A_6_;input A_7_;input B_0_;input B_1_;input B_2_;input B_3_;input B_4_;input B_5_;input B_6_;input B_7_;
  output SUM_0_;output SUM_1_;output SUM_2_;output SUM_3_;output SUM_4_;output SUM_5_;output SUM_6_;output SUM_7_;
  wire A_0__p;
  wire A_0__n;
  wire A_1__p;
  wire A_1__n;
  wire A_2__p;
  wire A_2__n;
  wire A_3__p;
  wire A_3__n;
  wire A_4__p;
  wire A_4__n;
  wire A_5__p;
  wire A_5__n;
  wire A_6__p;
  wire A_6__n;
  wire A_7__p;
  wire A_7__n;
  wire B_0__p;
  wire B_0__n;
  wire B_1__p;
  wire B_1__n;
  wire B_2__p;
  wire B_2__n;
  wire B_3__p;
  wire B_3__n;
  wire B_4__p;
  wire B_4__n;
  wire B_5__p;
  wire B_5__n;
  wire B_6__p;
  wire B_6__n;
  wire B_7__p;
  wire B_7__n;
  wire g17_p;
  wire g17_n;
  wire g18_p;
  wire g18_n;
  wire g19_p;
  wire g19_n;
  wire g20_p;
  wire g20_n;
  wire g21_p;
  wire g21_n;
  wire g22_p;
  wire g22_n;
  wire g23_p;
  wire g23_n;
  wire g24_p;
  wire g24_n;
  wire g25_p;
  wire g25_n;
  wire g26_p;
  wire g26_n;
  wire g27_p;
  wire g27_n;
  wire g28_p;
  wire g28_n;
  wire g29_p;
  wire g29_n;
  wire g30_p;
  wire g30_n;
  wire g31_p;
  wire g31_n;
  wire g32_p;
  wire g32_n;
  wire g33_p;
  wire g33_n;
  wire g34_p;
  wire g34_n;
  wire g35_p;
  wire g35_n;
  wire g36_p;
  wire g36_n;
  wire g37_p;
  wire g37_n;
  wire g38_p;
  wire g38_n;
  wire g39_p;
  wire g39_n;
  wire g40_p;
  wire g40_n;
  wire g41_p;
  wire g41_n;
  wire g42_p;
  wire g42_n;
  wire g43_p;
  wire g43_n;
  wire g44_p;
  wire g44_n;
  wire g45_p;
  wire g45_n;
  wire g46_p;
  wire g46_n;
  wire g47_p;
  wire g47_n;
  wire g48_p;
  wire g48_n;
  wire g49_p;
  wire g49_n;
  wire g50_p;
  wire g50_n;
  wire g51_p;
  wire g51_n;
  wire g52_p;
  wire g52_n;
  wire g53_p;
  wire g53_n;
  wire g54_p;
  wire g54_n;
  wire g55_p;
  wire g55_n;
  wire g56_p;
  wire g56_n;
  wire g57_p;
  wire g57_n;
  wire g58_p;
  wire g58_n;
  wire g59_p;
  wire g59_n;
  wire g60_p;
  wire g60_n;
  wire g61_p;
  wire g61_n;
  wire g62_p;
  wire g62_n;
  wire g63_p;
  wire g63_n;
  wire g64_p;
  wire g64_n;
  wire g65_p;
  wire g65_n;
  wire g66_p;
  wire g66_n;
  wire g67_p;
  wire g67_n;
  wire g68_p;
  wire g68_n;
  wire g69_p;
  wire g69_n;
  wire g70_p;
  wire g70_n;
  wire g71_p;
  wire g71_n;
  wire g72_p;
  wire g72_n;
  wire g73_p;
  wire g73_n;
  wire g74_p;
  wire g74_n;
  wire g75_p;
  wire g75_n;
  wire g76_p;
  wire g76_n;
  wire g77_p;
  wire g77_n;
  wire g78_p;
  wire g78_n;
  wire g79_p;
  wire g79_n;
  wire g80_p;
  wire g80_n;
  wire g81_p;
  wire g81_n;
  wire g82_p;
  wire g82_n;
  wire g83_p;
  wire g83_n;
  wire g84_p;
  wire g84_n;
  wire A_6__p_spl_;
  wire B_6__p_spl_;
  wire A_6__n_spl_;
  wire B_6__n_spl_;
  wire A_5__p_spl_;
  wire B_5__p_spl_;
  wire A_5__n_spl_;
  wire B_5__n_spl_;
  wire A_4__p_spl_;
  wire B_4__p_spl_;
  wire A_4__n_spl_;
  wire B_4__n_spl_;
  wire g19_n_spl_;
  wire g19_p_spl_;
  wire A_3__p_spl_;
  wire B_3__p_spl_;
  wire A_3__n_spl_;
  wire B_3__n_spl_;
  wire A_2__p_spl_;
  wire B_2__p_spl_;
  wire A_2__n_spl_;
  wire B_2__n_spl_;
  wire A_1__p_spl_;
  wire B_1__p_spl_;
  wire A_1__n_spl_;
  wire B_1__n_spl_;
  wire A_0__p_spl_;
  wire B_0__p_spl_;
  wire g27_n_spl_;
  wire g28_p_spl_;
  wire g27_p_spl_;
  wire g28_n_spl_;
  wire g28_n_spl_0;
  wire g26_n_spl_;
  wire g26_p_spl_;
  wire g25_n_spl_;
  wire g30_n_spl_;
  wire g25_p_spl_;
  wire g30_p_spl_;
  wire g24_n_spl_;
  wire g24_p_spl_;
  wire g23_n_spl_;
  wire g32_n_spl_;
  wire g23_p_spl_;
  wire g32_p_spl_;
  wire g22_n_spl_;
  wire g22_p_spl_;
  wire g21_p_spl_;
  wire g34_n_spl_;
  wire g35_n_spl_;
  wire g18_n_spl_;
  wire g18_p_spl_;
  wire g36_n_spl_;
  wire g38_p_spl_;
  wire g39_n_spl_;
  wire g17_p_spl_;
  wire g40_n_spl_;
  wire g42_p_spl_;
  wire A_7__n_spl_;
  wire B_7__n_spl_;
  wire g44_n_spl_;
  wire g44_n_spl_0;
  wire g45_p_spl_;
  wire g47_n_spl_;
  wire g48_n_spl_;
  wire g48_n_spl_0;
  wire g48_n_spl_00;
  wire g48_n_spl_01;
  wire g48_n_spl_1;
  wire g48_n_spl_10;
  wire g46_p_spl_;
  wire g46_p_spl_0;
  wire g46_p_spl_00;
  wire g46_p_spl_01;
  wire g46_p_spl_1;
  wire g46_p_spl_10;

  buf

  (
    A_0__p,
    A_0_
  );


  not

  (
    A_0__n,
    A_0_
  );


  buf

  (
    A_1__p,
    A_1_
  );


  not

  (
    A_1__n,
    A_1_
  );


  buf

  (
    A_2__p,
    A_2_
  );


  not

  (
    A_2__n,
    A_2_
  );


  buf

  (
    A_3__p,
    A_3_
  );


  not

  (
    A_3__n,
    A_3_
  );


  buf

  (
    A_4__p,
    A_4_
  );


  not

  (
    A_4__n,
    A_4_
  );


  buf

  (
    A_5__p,
    A_5_
  );


  not

  (
    A_5__n,
    A_5_
  );


  buf

  (
    A_6__p,
    A_6_
  );


  not

  (
    A_6__n,
    A_6_
  );


  buf

  (
    A_7__p,
    A_7_
  );


  not

  (
    A_7__n,
    A_7_
  );


  buf

  (
    B_0__p,
    B_0_
  );


  not

  (
    B_0__n,
    B_0_
  );


  buf

  (
    B_1__p,
    B_1_
  );


  not

  (
    B_1__n,
    B_1_
  );


  buf

  (
    B_2__p,
    B_2_
  );


  not

  (
    B_2__n,
    B_2_
  );


  buf

  (
    B_3__p,
    B_3_
  );


  not

  (
    B_3__n,
    B_3_
  );


  buf

  (
    B_4__p,
    B_4_
  );


  not

  (
    B_4__n,
    B_4_
  );


  buf

  (
    B_5__p,
    B_5_
  );


  not

  (
    B_5__n,
    B_5_
  );


  buf

  (
    B_6__p,
    B_6_
  );


  not

  (
    B_6__n,
    B_6_
  );


  buf

  (
    B_7__p,
    B_7_
  );


  not

  (
    B_7__n,
    B_7_
  );


  and

  (
    g17_p,
    A_6__p_spl_,
    B_6__p_spl_
  );


  or

  (
    g17_n,
    A_6__n_spl_,
    B_6__n_spl_
  );


  and

  (
    g18_p,
    A_5__p_spl_,
    B_5__p_spl_
  );


  or

  (
    g18_n,
    A_5__n_spl_,
    B_5__n_spl_
  );


  and

  (
    g19_p,
    A_4__p_spl_,
    B_4__p_spl_
  );


  or

  (
    g19_n,
    A_4__n_spl_,
    B_4__n_spl_
  );


  and

  (
    g20_p,
    A_4__n_spl_,
    B_4__n_spl_
  );


  or

  (
    g20_n,
    A_4__p_spl_,
    B_4__p_spl_
  );


  and

  (
    g21_p,
    g19_n_spl_,
    g20_n
  );


  or

  (
    g21_n,
    g19_p_spl_,
    g20_p
  );


  and

  (
    g22_p,
    A_3__p_spl_,
    B_3__p_spl_
  );


  or

  (
    g22_n,
    A_3__n_spl_,
    B_3__n_spl_
  );


  and

  (
    g23_p,
    A_3__n_spl_,
    B_3__n_spl_
  );


  or

  (
    g23_n,
    A_3__p_spl_,
    B_3__p_spl_
  );


  and

  (
    g24_p,
    A_2__p_spl_,
    B_2__p_spl_
  );


  or

  (
    g24_n,
    A_2__n_spl_,
    B_2__n_spl_
  );


  and

  (
    g25_p,
    A_2__n_spl_,
    B_2__n_spl_
  );


  or

  (
    g25_n,
    A_2__p_spl_,
    B_2__p_spl_
  );


  and

  (
    g26_p,
    A_1__p_spl_,
    B_1__p_spl_
  );


  or

  (
    g26_n,
    A_1__n_spl_,
    B_1__n_spl_
  );


  and

  (
    g27_p,
    A_1__n_spl_,
    B_1__n_spl_
  );


  or

  (
    g27_n,
    A_1__p_spl_,
    B_1__p_spl_
  );


  and

  (
    g28_p,
    A_0__p_spl_,
    B_0__p_spl_
  );


  or

  (
    g28_n,
    A_0__n,
    B_0__n
  );


  and

  (
    g29_p,
    g27_n_spl_,
    g28_p_spl_
  );


  or

  (
    g29_n,
    g27_p_spl_,
    g28_n_spl_0
  );


  and

  (
    g30_p,
    g26_n_spl_,
    g29_n
  );


  or

  (
    g30_n,
    g26_p_spl_,
    g29_p
  );


  and

  (
    g31_p,
    g25_n_spl_,
    g30_n_spl_
  );


  or

  (
    g31_n,
    g25_p_spl_,
    g30_p_spl_
  );


  and

  (
    g32_p,
    g24_n_spl_,
    g31_n
  );


  or

  (
    g32_n,
    g24_p_spl_,
    g31_p
  );


  and

  (
    g33_p,
    g23_n_spl_,
    g32_n_spl_
  );


  or

  (
    g33_n,
    g23_p_spl_,
    g32_p_spl_
  );


  and

  (
    g34_p,
    g22_n_spl_,
    g33_n
  );


  or

  (
    g34_n,
    g22_p_spl_,
    g33_p
  );


  and

  (
    g35_p,
    g21_p_spl_,
    g34_n_spl_
  );


  or

  (
    g35_n,
    g21_n,
    g34_p
  );


  and

  (
    g36_p,
    g19_n_spl_,
    g35_n_spl_
  );


  or

  (
    g36_n,
    g19_p_spl_,
    g35_p
  );


  and

  (
    g37_p,
    A_5__n_spl_,
    B_5__n_spl_
  );


  or

  (
    g37_n,
    A_5__p_spl_,
    B_5__p_spl_
  );


  and

  (
    g38_p,
    g18_n_spl_,
    g37_n
  );


  or

  (
    g38_n,
    g18_p_spl_,
    g37_p
  );


  and

  (
    g39_p,
    g36_n_spl_,
    g38_p_spl_
  );


  or

  (
    g39_n,
    g36_p,
    g38_n
  );


  and

  (
    g40_p,
    g18_n_spl_,
    g39_n_spl_
  );


  or

  (
    g40_n,
    g18_p_spl_,
    g39_p
  );


  and

  (
    g41_p,
    A_6__n_spl_,
    B_6__n_spl_
  );


  or

  (
    g41_n,
    A_6__p_spl_,
    B_6__p_spl_
  );


  and

  (
    g42_p,
    g17_n,
    g41_n
  );


  or

  (
    g42_n,
    g17_p_spl_,
    g41_p
  );


  and

  (
    g43_p,
    g40_n_spl_,
    g42_p_spl_
  );


  or

  (
    g43_n,
    g40_p,
    g42_n
  );


  or

  (
    g44_n,
    g17_p_spl_,
    g43_p
  );


  and

  (
    g45_p,
    A_7__n_spl_,
    B_7__n_spl_
  );


  and

  (
    g46_p,
    g44_n_spl_0,
    g45_p_spl_
  );


  or

  (
    g47_n,
    A_7__n_spl_,
    B_7__n_spl_
  );


  or

  (
    g48_n,
    g44_n_spl_0,
    g47_n_spl_
  );


  or

  (
    g49_n,
    A_0__p_spl_,
    B_0__p_spl_
  );


  and

  (
    g50_p,
    g28_n_spl_0,
    g49_n
  );


  and

  (
    g51_p,
    g48_n_spl_00,
    g50_p
  );


  or

  (
    g52_n,
    g46_p_spl_00,
    g51_p
  );


  and

  (
    g53_p,
    g26_n_spl_,
    g27_n_spl_
  );


  or

  (
    g53_n,
    g26_p_spl_,
    g27_p_spl_
  );


  or

  (
    g54_n,
    g28_n_spl_,
    g53_n
  );


  or

  (
    g55_n,
    g28_p_spl_,
    g53_p
  );


  and

  (
    g56_p,
    g54_n,
    g55_n
  );


  and

  (
    g57_p,
    g48_n_spl_00,
    g56_p
  );


  or

  (
    g58_n,
    g46_p_spl_00,
    g57_p
  );


  and

  (
    g59_p,
    g24_n_spl_,
    g25_n_spl_
  );


  or

  (
    g59_n,
    g24_p_spl_,
    g25_p_spl_
  );


  and

  (
    g60_p,
    g30_p_spl_,
    g59_p
  );


  and

  (
    g61_p,
    g30_n_spl_,
    g59_n
  );


  or

  (
    g62_n,
    g60_p,
    g61_p
  );


  and

  (
    g63_p,
    g48_n_spl_01,
    g62_n
  );


  or

  (
    g64_n,
    g46_p_spl_01,
    g63_p
  );


  and

  (
    g65_p,
    g22_n_spl_,
    g23_n_spl_
  );


  or

  (
    g65_n,
    g22_p_spl_,
    g23_p_spl_
  );


  or

  (
    g66_n,
    g32_p_spl_,
    g65_n
  );


  or

  (
    g67_n,
    g32_n_spl_,
    g65_p
  );


  and

  (
    g68_p,
    g66_n,
    g67_n
  );


  and

  (
    g69_p,
    g48_n_spl_01,
    g68_p
  );


  or

  (
    g70_n,
    g46_p_spl_01,
    g69_p
  );


  or

  (
    g71_n,
    g21_p_spl_,
    g34_n_spl_
  );


  and

  (
    g72_p,
    g35_n_spl_,
    g71_n
  );


  and

  (
    g73_p,
    g48_n_spl_10,
    g72_p
  );


  or

  (
    g74_n,
    g46_p_spl_10,
    g73_p
  );


  or

  (
    g75_n,
    g36_n_spl_,
    g38_p_spl_
  );


  and

  (
    g76_p,
    g39_n_spl_,
    g75_n
  );


  and

  (
    g77_p,
    g48_n_spl_10,
    g76_p
  );


  or

  (
    g78_n,
    g46_p_spl_10,
    g77_p
  );


  or

  (
    g79_n,
    g40_n_spl_,
    g42_p_spl_
  );


  and

  (
    g80_p,
    g43_n,
    g79_n
  );


  and

  (
    g81_p,
    g48_n_spl_1,
    g80_p
  );


  or

  (
    g82_n,
    g46_p_spl_1,
    g81_p
  );


  or

  (
    g83_n,
    g44_n_spl_,
    g45_p_spl_
  );


  and

  (
    g84_p,
    g47_n_spl_,
    g83_n
  );


  buf

  (
    SUM_0_,
    g52_n
  );


  buf

  (
    SUM_1_,
    g58_n
  );


  buf

  (
    SUM_2_,
    g64_n
  );


  buf

  (
    SUM_3_,
    g70_n
  );


  buf

  (
    SUM_4_,
    g74_n
  );


  buf

  (
    SUM_5_,
    g78_n
  );


  buf

  (
    SUM_6_,
    g82_n
  );


  not

  (
    SUM_7_,
    g84_p
  );


  buf

  (
    A_6__p_spl_,
    A_6__p
  );


  buf

  (
    B_6__p_spl_,
    B_6__p
  );


  buf

  (
    A_6__n_spl_,
    A_6__n
  );


  buf

  (
    B_6__n_spl_,
    B_6__n
  );


  buf

  (
    A_5__p_spl_,
    A_5__p
  );


  buf

  (
    B_5__p_spl_,
    B_5__p
  );


  buf

  (
    A_5__n_spl_,
    A_5__n
  );


  buf

  (
    B_5__n_spl_,
    B_5__n
  );


  buf

  (
    A_4__p_spl_,
    A_4__p
  );


  buf

  (
    B_4__p_spl_,
    B_4__p
  );


  buf

  (
    A_4__n_spl_,
    A_4__n
  );


  buf

  (
    B_4__n_spl_,
    B_4__n
  );


  buf

  (
    g19_n_spl_,
    g19_n
  );


  buf

  (
    g19_p_spl_,
    g19_p
  );


  buf

  (
    A_3__p_spl_,
    A_3__p
  );


  buf

  (
    B_3__p_spl_,
    B_3__p
  );


  buf

  (
    A_3__n_spl_,
    A_3__n
  );


  buf

  (
    B_3__n_spl_,
    B_3__n
  );


  buf

  (
    A_2__p_spl_,
    A_2__p
  );


  buf

  (
    B_2__p_spl_,
    B_2__p
  );


  buf

  (
    A_2__n_spl_,
    A_2__n
  );


  buf

  (
    B_2__n_spl_,
    B_2__n
  );


  buf

  (
    A_1__p_spl_,
    A_1__p
  );


  buf

  (
    B_1__p_spl_,
    B_1__p
  );


  buf

  (
    A_1__n_spl_,
    A_1__n
  );


  buf

  (
    B_1__n_spl_,
    B_1__n
  );


  buf

  (
    A_0__p_spl_,
    A_0__p
  );


  buf

  (
    B_0__p_spl_,
    B_0__p
  );


  buf

  (
    g27_n_spl_,
    g27_n
  );


  buf

  (
    g28_p_spl_,
    g28_p
  );


  buf

  (
    g27_p_spl_,
    g27_p
  );


  buf

  (
    g28_n_spl_,
    g28_n
  );


  buf

  (
    g28_n_spl_0,
    g28_n_spl_
  );


  buf

  (
    g26_n_spl_,
    g26_n
  );


  buf

  (
    g26_p_spl_,
    g26_p
  );


  buf

  (
    g25_n_spl_,
    g25_n
  );


  buf

  (
    g30_n_spl_,
    g30_n
  );


  buf

  (
    g25_p_spl_,
    g25_p
  );


  buf

  (
    g30_p_spl_,
    g30_p
  );


  buf

  (
    g24_n_spl_,
    g24_n
  );


  buf

  (
    g24_p_spl_,
    g24_p
  );


  buf

  (
    g23_n_spl_,
    g23_n
  );


  buf

  (
    g32_n_spl_,
    g32_n
  );


  buf

  (
    g23_p_spl_,
    g23_p
  );


  buf

  (
    g32_p_spl_,
    g32_p
  );


  buf

  (
    g22_n_spl_,
    g22_n
  );


  buf

  (
    g22_p_spl_,
    g22_p
  );


  buf

  (
    g21_p_spl_,
    g21_p
  );


  buf

  (
    g34_n_spl_,
    g34_n
  );


  buf

  (
    g35_n_spl_,
    g35_n
  );


  buf

  (
    g18_n_spl_,
    g18_n
  );


  buf

  (
    g18_p_spl_,
    g18_p
  );


  buf

  (
    g36_n_spl_,
    g36_n
  );


  buf

  (
    g38_p_spl_,
    g38_p
  );


  buf

  (
    g39_n_spl_,
    g39_n
  );


  buf

  (
    g17_p_spl_,
    g17_p
  );


  buf

  (
    g40_n_spl_,
    g40_n
  );


  buf

  (
    g42_p_spl_,
    g42_p
  );


  buf

  (
    A_7__n_spl_,
    A_7__n
  );


  buf

  (
    B_7__n_spl_,
    B_7__n
  );


  buf

  (
    g44_n_spl_,
    g44_n
  );


  buf

  (
    g44_n_spl_0,
    g44_n_spl_
  );


  buf

  (
    g45_p_spl_,
    g45_p
  );


  buf

  (
    g47_n_spl_,
    g47_n
  );


  buf

  (
    g48_n_spl_,
    g48_n
  );


  buf

  (
    g48_n_spl_0,
    g48_n_spl_
  );


  buf

  (
    g48_n_spl_00,
    g48_n_spl_0
  );


  buf

  (
    g48_n_spl_01,
    g48_n_spl_0
  );


  buf

  (
    g48_n_spl_1,
    g48_n_spl_
  );


  buf

  (
    g48_n_spl_10,
    g48_n_spl_1
  );


  buf

  (
    g46_p_spl_,
    g46_p
  );


  buf

  (
    g46_p_spl_0,
    g46_p_spl_
  );


  buf

  (
    g46_p_spl_00,
    g46_p_spl_0
  );


  buf

  (
    g46_p_spl_01,
    g46_p_spl_0
  );


  buf

  (
    g46_p_spl_1,
    g46_p_spl_
  );


  buf

  (
    g46_p_spl_10,
    g46_p_spl_1
  );


endmodule
