// Benchmark "mymod" written by ABC on Sun Oct 29 19:31:50 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58,
    G59, G60,
    G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, G865, G866,
    G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, G877, G878,
    G879, G880  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G58, G59, G60;
  output G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, G865,
    G866, G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, G877,
    G878, G879, G880;
  reg n480_lo, n492_lo, n495_lo, n498_lo, n501_lo, n504_lo, n516_lo,
    n528_lo, n531_lo, n540_lo, n543_lo, n546_lo, n549_lo, n552_lo, n564_lo,
    n579_lo, n600_lo, n603_lo, n606_lo, n609_lo, n612_lo, n615_lo, n618_lo,
    n621_lo, n627_lo, n630_lo, n633_lo, n639_lo, n642_lo, n645_lo, n648_lo,
    n660_lo, n663_lo, n672_lo, n675_lo, n678_lo, n681_lo, n684_lo, n687_lo,
    n690_lo, n693_lo, n696_lo, n699_lo, n702_lo, n705_lo, n708_lo, n711_lo,
    n714_lo, n717_lo, n720_lo, n723_lo, n726_lo, n729_lo, n732_lo, n735_lo,
    n738_lo, n741_lo, n744_lo, n747_lo, n750_lo, n756_lo, n759_lo, n762_lo,
    n768_lo, n771_lo, n774_lo, n780_lo, n783_lo, n786_lo, n792_lo, n795_lo,
    n804_lo, n807_lo, n816_lo, n819_lo, n828_lo, n831_lo, n843_lo, n846_lo,
    n849_lo, n852_lo, n855_lo, n858_lo, n861_lo, n864_lo, n867_lo, n870_lo,
    n879_lo, n891_lo, n903_lo, n915_lo, n918_lo, n927_lo, n951_lo, n954_lo,
    n957_lo, n960_lo, n963_lo, n966_lo, n972_lo, n975_lo, n978_lo, n984_lo,
    n987_lo, n990_lo, n996_lo, n999_lo, n1002_lo, n1008_lo, n1011_lo,
    n1014_lo, n1020_lo, n1023_lo, n1026_lo, n1032_lo, n1035_lo, n1038_lo,
    n1044_lo, n1047_lo, n1050_lo, n1053_lo, n1056_lo, n1059_lo, n1062_lo,
    n1065_lo, n1068_lo, n1071_lo, n1074_lo, n1077_lo, n1080_lo, n1083_lo,
    n1086_lo, n1089_lo, n1092_lo, n1095_lo, n1098_lo, n1101_lo, n1104_lo,
    n1107_lo, n1110_lo, n1113_lo, n1116_lo, n1119_lo, n1122_lo, n1125_lo,
    n1128_lo, n1131_lo, n1134_lo, n1137_lo, n1140_lo, n1143_lo, n1146_lo,
    n1149_lo, n1152_lo, n1155_lo, n1158_lo, n1167_lo, n1170_lo, n1173_lo,
    n1176_lo, n1179_lo, n1529_o2, n1616_o2, n1655_o2, n1656_o2, n1657_o2,
    n1730_o2, n1731_o2, n1732_o2, n1729_o2, n1805_o2, n1808_o2, n1807_o2,
    n1809_o2, n1663_o2, n1664_o2, n1704_o2, n1705_o2, n1706_o2, n1707_o2,
    n1708_o2, n1709_o2, G280_o2, G655_o2, G663_o2, G672_o2, G538_o2,
    n1780_o2, n1781_o2, n1797_o2, n1798_o2, n1799_o2, n1800_o2, G578_o2,
    n1828_o2, n801_lo_buf_o2, G693_o2, G702_o2, G712_o2, G685_o2, G658_o2,
    G667_o2, G677_o2, G650_o2, G798_o2, n1017_lo_buf_o2, n1029_lo_buf_o2,
    n1041_lo_buf_o2, G558_o2, G562_o2, G566_o2, n1835_o2, n1836_o2,
    n1837_o2, n765_lo_buf_o2, n777_lo_buf_o2, n789_lo_buf_o2, G617_o2,
    G626_o2, G636_o2, n489_lo_buf_o2, n513_lo_buf_o2, n561_lo_buf_o2,
    n597_lo_buf_o2, n657_lo_buf_o2, G276_o2, n1005_lo_buf_o2,
    n1161_lo_buf_o2, G620_o2, G629_o2, G639_o2, G554_o2, G690_o2, G698_o2,
    G707_o2, G319_o2, G389_o2, n753_lo_buf_o2, G647_o2, G769_o2, G785_o2,
    G808_o2, G445_o2, G448_o2, G477_o2, G480_o2, G436_o2, G786_o2, G787_o2,
    G826_o2, G827_o2, G825_o2, G610_o2, n537_lo_buf_o2, n669_lo_buf_o2,
    n969_lo_buf_o2, n981_lo_buf_o2, n993_lo_buf_o2, G309_o2, G461_o2,
    G487_o2, G460_o2, G468_o2, G287_o2, G613_o2, n585_lo_buf_o2,
    n813_lo_buf_o2, n825_lo_buf_o2, n837_lo_buf_o2, n897_lo_buf_o2,
    n909_lo_buf_o2, n933_lo_buf_o2, G451_o2, G682_o2, G756_o2, G542_o2,
    G546_o2, G550_o2, G310_o2, n798_lo_buf_o2, n882_lo_buf_o2, G427_o2,
    G497_o2, G499_o2, G501_o2, G498_o2, G500_o2, G502_o2, G369_o2,
    n939_lo_buf_o2, n486_lo_buf_o2, n510_lo_buf_o2, n558_lo_buf_o2,
    n594_lo_buf_o2, n654_lo_buf_o2, n477_lo_buf_o2, n525_lo_buf_o2,
    n573_lo_buf_o2;
  wire new_n683_, new_n685_, new_n687_, new_n689_, new_n691_, new_n693_,
    new_n695_, new_n697_, new_n699_, new_n701_, new_n703_, new_n705_,
    new_n707_, new_n709_, new_n711_, new_n713_, new_n715_, new_n717_,
    new_n719_, new_n721_, new_n723_, new_n725_, new_n727_, new_n729_,
    new_n731_, new_n733_, new_n735_, new_n737_, new_n739_, new_n741_,
    new_n743_, new_n745_, new_n747_, new_n749_, new_n751_, new_n753_,
    new_n755_, new_n757_, new_n759_, new_n761_, new_n763_, new_n765_,
    new_n767_, new_n769_, new_n771_, new_n773_, new_n775_, new_n777_,
    new_n779_, new_n781_, new_n783_, new_n785_, new_n787_, new_n789_,
    new_n791_, new_n793_, new_n795_, new_n797_, new_n799_, new_n801_,
    new_n803_, new_n804_, new_n806_, new_n807_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n825_,
    new_n827_, new_n830_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n847_, new_n850_, new_n851_, new_n853_, new_n856_,
    new_n857_, new_n859_, new_n861_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n875_, new_n878_, new_n879_, new_n881_, new_n883_, new_n886_,
    new_n887_, new_n889_, new_n891_, new_n893_, new_n895_, new_n897_,
    new_n899_, new_n901_, new_n903_, new_n905_, new_n907_, new_n909_,
    new_n911_, new_n913_, new_n915_, new_n917_, new_n919_, new_n921_,
    new_n924_, new_n925_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n942_, new_n943_, new_n946_, new_n947_, new_n950_, new_n951_,
    new_n954_, new_n955_, new_n957_, new_n959_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n969_, new_n971_, new_n972_,
    new_n973_, new_n975_, new_n976_, new_n977_, new_n979_, new_n981_,
    new_n983_, new_n986_, new_n987_, new_n989_, new_n991_, new_n993_,
    new_n994_, new_n996_, new_n997_, new_n999_, new_n1002_, new_n1003_,
    new_n1005_, new_n1008_, new_n1009_, new_n1011_, new_n1014_, new_n1015_,
    new_n1017_, new_n1018_, new_n1020_, new_n1021_, new_n1023_, new_n1024_,
    new_n1026_, new_n1027_, new_n1029_, new_n1030_, new_n1032_, new_n1033_,
    new_n1035_, new_n1036_, new_n1038_, new_n1039_, new_n1041_, new_n1043_,
    new_n1045_, new_n1046_, new_n1047_, new_n1049_, new_n1051_, new_n1054_,
    new_n1055_, new_n1057_, new_n1059_, new_n1062_, new_n1063_, new_n1065_,
    new_n1067_, new_n1070_, new_n1071_, new_n1073_, new_n1075_, new_n1078_,
    new_n1079_, new_n1081_, new_n1083_, new_n1086_, new_n1087_, new_n1089_,
    new_n1091_, new_n1094_, new_n1095_, new_n1097_, new_n1099_, new_n1102_,
    new_n1103_, new_n1105_, new_n1107_, new_n1110_, new_n1111_, new_n1113_,
    new_n1114_, new_n1115_, new_n1117_, new_n1119_, new_n1122_, new_n1123_,
    new_n1126_, new_n1128_, new_n1130_, new_n1132_, new_n1134_, new_n1136_,
    new_n1138_, new_n1140_, new_n1142_, new_n1144_, new_n1146_, new_n1148_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1155_, new_n1156_,
    new_n1157_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1165_, new_n1168_, new_n1170_, new_n1172_, new_n1174_, new_n1176_,
    new_n1177_, new_n1179_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1190_, new_n1191_, new_n1193_,
    new_n1194_, new_n1196_, new_n1198_, new_n1200_, new_n1202_, new_n1204_,
    new_n1206_, new_n1208_, new_n1210_, new_n1212_, new_n1213_, new_n1214_,
    new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1221_,
    new_n1223_, new_n1225_, new_n1227_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1245_,
    new_n1246_, new_n1247_, new_n1249_, new_n1251_, new_n1253_, new_n1255_,
    new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1267_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1276_, new_n1277_,
    new_n1278_, new_n1280_, new_n1282_, new_n1284_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1296_, new_n1298_, new_n1300_, new_n1302_, new_n1304_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1311_, new_n1313_,
    new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_,
    new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1337_, new_n1339_, new_n1342_, new_n1344_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1361_, new_n1362_, new_n1364_, new_n1366_,
    new_n1368_, new_n1370_, new_n1372_, new_n1374_, new_n1376_, new_n1378_,
    new_n1379_, new_n1381_, new_n1382_, new_n1383_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n2141_, new_n2142_,
    new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_,
    new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_,
    new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_,
    new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_,
    new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_,
    new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_,
    new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_,
    new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_,
    new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_,
    new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_,
    new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_,
    new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_,
    new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_,
    new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_,
    new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_,
    new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_,
    new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_,
    new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_,
    new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_,
    new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_,
    new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_,
    new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_,
    new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_,
    new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_,
    new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, n480_li, n492_li, n495_li, n498_li, n501_li,
    n504_li, n516_li, n528_li, n531_li, n540_li, n543_li, n546_li, n549_li,
    n552_li, n564_li, n579_li, n600_li, n603_li, n606_li, n609_li, n612_li,
    n615_li, n618_li, n621_li, n627_li, n630_li, n633_li, n639_li, n642_li,
    n645_li, n648_li, n660_li, n663_li, n672_li, n675_li, n678_li, n681_li,
    n684_li, n687_li, n690_li, n693_li, n696_li, n699_li, n702_li, n705_li,
    n708_li, n711_li, n714_li, n717_li, n720_li, n723_li, n726_li, n729_li,
    n732_li, n735_li, n738_li, n741_li, n744_li, n747_li, n750_li, n756_li,
    n759_li, n762_li, n768_li, n771_li, n774_li, n780_li, n783_li, n786_li,
    n792_li, n795_li, n804_li, n807_li, n816_li, n819_li, n828_li, n831_li,
    n843_li, n846_li, n849_li, n852_li, n855_li, n858_li, n861_li, n864_li,
    n867_li, n870_li, n879_li, n891_li, n903_li, n915_li, n918_li, n927_li,
    n951_li, n954_li, n957_li, n960_li, n963_li, n966_li, n972_li, n975_li,
    n978_li, n984_li, n987_li, n990_li, n996_li, n999_li, n1002_li,
    n1008_li, n1011_li, n1014_li, n1020_li, n1023_li, n1026_li, n1032_li,
    n1035_li, n1038_li, n1044_li, n1047_li, n1050_li, n1053_li, n1056_li,
    n1059_li, n1062_li, n1065_li, n1068_li, n1071_li, n1074_li, n1077_li,
    n1080_li, n1083_li, n1086_li, n1089_li, n1092_li, n1095_li, n1098_li,
    n1101_li, n1104_li, n1107_li, n1110_li, n1113_li, n1116_li, n1119_li,
    n1122_li, n1125_li, n1128_li, n1131_li, n1134_li, n1137_li, n1140_li,
    n1143_li, n1146_li, n1149_li, n1152_li, n1155_li, n1158_li, n1167_li,
    n1170_li, n1173_li, n1176_li, n1179_li, n1529_i2, n1616_i2, n1655_i2,
    n1656_i2, n1657_i2, n1730_i2, n1731_i2, n1732_i2, n1729_i2, n1805_i2,
    n1808_i2, n1807_i2, n1809_i2, n1663_i2, n1664_i2, n1704_i2, n1705_i2,
    n1706_i2, n1707_i2, n1708_i2, n1709_i2, G280_i2, G655_i2, G663_i2,
    G672_i2, G538_i2, n1780_i2, n1781_i2, n1797_i2, n1798_i2, n1799_i2,
    n1800_i2, G578_i2, n1828_i2, n801_lo_buf_i2, G693_i2, G702_i2, G712_i2,
    G685_i2, G658_i2, G667_i2, G677_i2, G650_i2, G798_i2, n1017_lo_buf_i2,
    n1029_lo_buf_i2, n1041_lo_buf_i2, G558_i2, G562_i2, G566_i2, n1835_i2,
    n1836_i2, n1837_i2, n765_lo_buf_i2, n777_lo_buf_i2, n789_lo_buf_i2,
    G617_i2, G626_i2, G636_i2, n489_lo_buf_i2, n513_lo_buf_i2,
    n561_lo_buf_i2, n597_lo_buf_i2, n657_lo_buf_i2, G276_i2,
    n1005_lo_buf_i2, n1161_lo_buf_i2, G620_i2, G629_i2, G639_i2, G554_i2,
    G690_i2, G698_i2, G707_i2, G319_i2, G389_i2, n753_lo_buf_i2, G647_i2,
    G769_i2, G785_i2, G808_i2, G445_i2, G448_i2, G477_i2, G480_i2, G436_i2,
    G786_i2, G787_i2, G826_i2, G827_i2, G825_i2, G610_i2, n537_lo_buf_i2,
    n669_lo_buf_i2, n969_lo_buf_i2, n981_lo_buf_i2, n993_lo_buf_i2,
    G309_i2, G461_i2, G487_i2, G460_i2, G468_i2, G287_i2, G613_i2,
    n585_lo_buf_i2, n813_lo_buf_i2, n825_lo_buf_i2, n837_lo_buf_i2,
    n897_lo_buf_i2, n909_lo_buf_i2, n933_lo_buf_i2, G451_i2, G682_i2,
    G756_i2, G542_i2, G546_i2, G550_i2, G310_i2, n798_lo_buf_i2,
    n882_lo_buf_i2, G427_i2, G497_i2, G499_i2, G501_i2, G498_i2, G500_i2,
    G502_i2, G369_i2, n939_lo_buf_i2, n486_lo_buf_i2, n510_lo_buf_i2,
    n558_lo_buf_i2, n594_lo_buf_i2, n654_lo_buf_i2, n477_lo_buf_i2,
    n525_lo_buf_i2, n573_lo_buf_i2;
  assign new_n683_ = G1;
  assign new_n685_ = G2;
  assign new_n687_ = G3;
  assign new_n689_ = G4;
  assign new_n691_ = G5;
  assign new_n693_ = G6;
  assign new_n695_ = G7;
  assign new_n697_ = G8;
  assign new_n699_ = G9;
  assign new_n701_ = G10;
  assign new_n703_ = G11;
  assign new_n705_ = G12;
  assign new_n707_ = G13;
  assign new_n709_ = G14;
  assign new_n711_ = G15;
  assign new_n713_ = G16;
  assign new_n715_ = G17;
  assign new_n717_ = G18;
  assign new_n719_ = G19;
  assign new_n721_ = G20;
  assign new_n723_ = G21;
  assign new_n725_ = G22;
  assign new_n727_ = G23;
  assign new_n729_ = G24;
  assign new_n731_ = G25;
  assign new_n733_ = G26;
  assign new_n735_ = G27;
  assign new_n737_ = G28;
  assign new_n739_ = G29;
  assign new_n741_ = G30;
  assign new_n743_ = G31;
  assign new_n745_ = G32;
  assign new_n747_ = G33;
  assign new_n749_ = G34;
  assign new_n751_ = G35;
  assign new_n753_ = G36;
  assign new_n755_ = G37;
  assign new_n757_ = G38;
  assign new_n759_ = G39;
  assign new_n761_ = G40;
  assign new_n763_ = G41;
  assign new_n765_ = G42;
  assign new_n767_ = G43;
  assign new_n769_ = G44;
  assign new_n771_ = G45;
  assign new_n773_ = G46;
  assign new_n775_ = G47;
  assign new_n777_ = G48;
  assign new_n779_ = G49;
  assign new_n781_ = G50;
  assign new_n783_ = G51;
  assign new_n785_ = G52;
  assign new_n787_ = G53;
  assign new_n789_ = G54;
  assign new_n791_ = G55;
  assign new_n793_ = G56;
  assign new_n795_ = G57;
  assign new_n797_ = G58;
  assign new_n799_ = G59;
  assign new_n801_ = G60;
  assign new_n803_ = n480_lo;
  assign new_n804_ = ~n480_lo;
  assign new_n806_ = ~n492_lo;
  assign new_n807_ = n495_lo;
  assign new_n809_ = n498_lo;
  assign new_n811_ = n501_lo;
  assign new_n812_ = ~n501_lo;
  assign new_n813_ = n504_lo;
  assign new_n814_ = ~n504_lo;
  assign new_n815_ = n516_lo;
  assign new_n816_ = ~n516_lo;
  assign new_n817_ = n528_lo;
  assign new_n818_ = ~n528_lo;
  assign new_n819_ = n531_lo;
  assign new_n820_ = ~n531_lo;
  assign new_n822_ = ~n540_lo;
  assign new_n823_ = n543_lo;
  assign new_n825_ = n546_lo;
  assign new_n827_ = n549_lo;
  assign new_n830_ = ~n552_lo;
  assign new_n832_ = ~n564_lo;
  assign new_n833_ = n579_lo;
  assign new_n834_ = ~n579_lo;
  assign new_n835_ = n600_lo;
  assign new_n836_ = ~n600_lo;
  assign new_n837_ = n603_lo;
  assign new_n839_ = n606_lo;
  assign new_n841_ = n609_lo;
  assign new_n842_ = ~n609_lo;
  assign new_n844_ = ~n612_lo;
  assign new_n845_ = n615_lo;
  assign new_n847_ = n618_lo;
  assign new_n850_ = ~n621_lo;
  assign new_n851_ = n627_lo;
  assign new_n853_ = n630_lo;
  assign new_n856_ = ~n633_lo;
  assign new_n857_ = n639_lo;
  assign new_n859_ = n642_lo;
  assign new_n861_ = n645_lo;
  assign new_n864_ = ~n648_lo;
  assign new_n865_ = n660_lo;
  assign new_n866_ = ~n660_lo;
  assign new_n867_ = n663_lo;
  assign new_n868_ = ~n663_lo;
  assign new_n869_ = n672_lo;
  assign new_n870_ = ~n672_lo;
  assign new_n871_ = n675_lo;
  assign new_n873_ = n678_lo;
  assign new_n875_ = n681_lo;
  assign new_n878_ = ~n684_lo;
  assign new_n879_ = n687_lo;
  assign new_n881_ = n690_lo;
  assign new_n883_ = n693_lo;
  assign new_n886_ = ~n696_lo;
  assign new_n887_ = n699_lo;
  assign new_n889_ = n702_lo;
  assign new_n891_ = n705_lo;
  assign new_n893_ = n708_lo;
  assign new_n895_ = n711_lo;
  assign new_n897_ = n714_lo;
  assign new_n899_ = n717_lo;
  assign new_n901_ = n720_lo;
  assign new_n903_ = n723_lo;
  assign new_n905_ = n726_lo;
  assign new_n907_ = n729_lo;
  assign new_n909_ = n732_lo;
  assign new_n911_ = n735_lo;
  assign new_n913_ = n738_lo;
  assign new_n915_ = n741_lo;
  assign new_n917_ = n744_lo;
  assign new_n919_ = n747_lo;
  assign new_n921_ = n750_lo;
  assign new_n924_ = ~n756_lo;
  assign new_n925_ = n759_lo;
  assign new_n927_ = n762_lo;
  assign new_n928_ = ~n762_lo;
  assign new_n930_ = ~n768_lo;
  assign new_n931_ = n771_lo;
  assign new_n933_ = n774_lo;
  assign new_n934_ = ~n774_lo;
  assign new_n936_ = ~n780_lo;
  assign new_n937_ = n783_lo;
  assign new_n939_ = n786_lo;
  assign new_n940_ = ~n786_lo;
  assign new_n942_ = ~n792_lo;
  assign new_n943_ = n795_lo;
  assign new_n946_ = ~n804_lo;
  assign new_n947_ = n807_lo;
  assign new_n950_ = ~n816_lo;
  assign new_n951_ = n819_lo;
  assign new_n954_ = ~n828_lo;
  assign new_n955_ = n831_lo;
  assign new_n957_ = n843_lo;
  assign new_n959_ = n846_lo;
  assign new_n961_ = n849_lo;
  assign new_n963_ = n852_lo;
  assign new_n964_ = ~n852_lo;
  assign new_n965_ = n855_lo;
  assign new_n967_ = n858_lo;
  assign new_n969_ = n861_lo;
  assign new_n971_ = n864_lo;
  assign new_n972_ = ~n864_lo;
  assign new_n973_ = n867_lo;
  assign new_n975_ = n870_lo;
  assign new_n976_ = ~n870_lo;
  assign new_n977_ = n879_lo;
  assign new_n979_ = n891_lo;
  assign new_n981_ = n903_lo;
  assign new_n983_ = n915_lo;
  assign new_n986_ = ~n918_lo;
  assign new_n987_ = n927_lo;
  assign new_n989_ = n951_lo;
  assign new_n991_ = n954_lo;
  assign new_n993_ = n957_lo;
  assign new_n994_ = ~n957_lo;
  assign new_n996_ = ~n960_lo;
  assign new_n997_ = n963_lo;
  assign new_n999_ = n966_lo;
  assign new_n1002_ = ~n972_lo;
  assign new_n1003_ = n975_lo;
  assign new_n1005_ = n978_lo;
  assign new_n1008_ = ~n984_lo;
  assign new_n1009_ = n987_lo;
  assign new_n1011_ = n990_lo;
  assign new_n1014_ = ~n996_lo;
  assign new_n1015_ = n999_lo;
  assign new_n1017_ = n1002_lo;
  assign new_n1018_ = ~n1002_lo;
  assign new_n1020_ = ~n1008_lo;
  assign new_n1021_ = n1011_lo;
  assign new_n1023_ = n1014_lo;
  assign new_n1024_ = ~n1014_lo;
  assign new_n1026_ = ~n1020_lo;
  assign new_n1027_ = n1023_lo;
  assign new_n1029_ = n1026_lo;
  assign new_n1030_ = ~n1026_lo;
  assign new_n1032_ = ~n1032_lo;
  assign new_n1033_ = n1035_lo;
  assign new_n1035_ = n1038_lo;
  assign new_n1036_ = ~n1038_lo;
  assign new_n1038_ = ~n1044_lo;
  assign new_n1039_ = n1047_lo;
  assign new_n1041_ = n1050_lo;
  assign new_n1043_ = n1053_lo;
  assign new_n1045_ = n1056_lo;
  assign new_n1046_ = ~n1056_lo;
  assign new_n1047_ = n1059_lo;
  assign new_n1049_ = n1062_lo;
  assign new_n1051_ = n1065_lo;
  assign new_n1054_ = ~n1068_lo;
  assign new_n1055_ = n1071_lo;
  assign new_n1057_ = n1074_lo;
  assign new_n1059_ = n1077_lo;
  assign new_n1062_ = ~n1080_lo;
  assign new_n1063_ = n1083_lo;
  assign new_n1065_ = n1086_lo;
  assign new_n1067_ = n1089_lo;
  assign new_n1070_ = ~n1092_lo;
  assign new_n1071_ = n1095_lo;
  assign new_n1073_ = n1098_lo;
  assign new_n1075_ = n1101_lo;
  assign new_n1078_ = ~n1104_lo;
  assign new_n1079_ = n1107_lo;
  assign new_n1081_ = n1110_lo;
  assign new_n1083_ = n1113_lo;
  assign new_n1086_ = ~n1116_lo;
  assign new_n1087_ = n1119_lo;
  assign new_n1089_ = n1122_lo;
  assign new_n1091_ = n1125_lo;
  assign new_n1094_ = ~n1128_lo;
  assign new_n1095_ = n1131_lo;
  assign new_n1097_ = n1134_lo;
  assign new_n1099_ = n1137_lo;
  assign new_n1102_ = ~n1140_lo;
  assign new_n1103_ = n1143_lo;
  assign new_n1105_ = n1146_lo;
  assign new_n1107_ = n1149_lo;
  assign new_n1110_ = ~n1152_lo;
  assign new_n1111_ = n1155_lo;
  assign new_n1113_ = n1158_lo;
  assign new_n1114_ = ~n1158_lo;
  assign new_n1115_ = n1167_lo;
  assign new_n1117_ = n1170_lo;
  assign new_n1119_ = n1173_lo;
  assign new_n1122_ = ~n1176_lo;
  assign new_n1123_ = n1179_lo;
  assign new_n1126_ = ~n1529_o2;
  assign new_n1128_ = ~n1616_o2;
  assign new_n1130_ = ~n1655_o2;
  assign new_n1132_ = ~n1656_o2;
  assign new_n1134_ = ~n1657_o2;
  assign new_n1136_ = ~n1730_o2;
  assign new_n1138_ = ~n1731_o2;
  assign new_n1140_ = ~n1732_o2;
  assign new_n1142_ = ~n1729_o2;
  assign new_n1144_ = ~n1805_o2;
  assign new_n1146_ = ~n1808_o2;
  assign new_n1148_ = ~n1807_o2;
  assign new_n1150_ = ~n1809_o2;
  assign new_n1151_ = n1663_o2;
  assign new_n1152_ = ~n1663_o2;
  assign new_n1153_ = n1664_o2;
  assign new_n1155_ = n1704_o2;
  assign new_n1156_ = ~n1704_o2;
  assign new_n1157_ = n1705_o2;
  assign new_n1159_ = n1706_o2;
  assign new_n1160_ = ~n1706_o2;
  assign new_n1161_ = n1707_o2;
  assign new_n1162_ = ~n1707_o2;
  assign new_n1163_ = n1708_o2;
  assign new_n1165_ = n1709_o2;
  assign new_n1168_ = ~G280_o2;
  assign new_n1170_ = ~G655_o2;
  assign new_n1172_ = ~G663_o2;
  assign new_n1174_ = ~G672_o2;
  assign new_n1176_ = ~G538_o2;
  assign new_n1177_ = n1780_o2;
  assign new_n1179_ = n1781_o2;
  assign new_n1182_ = ~n1797_o2;
  assign new_n1183_ = n1798_o2;
  assign new_n1184_ = ~n1798_o2;
  assign new_n1185_ = n1799_o2;
  assign new_n1186_ = ~n1799_o2;
  assign new_n1187_ = n1800_o2;
  assign new_n1188_ = ~n1800_o2;
  assign new_n1190_ = ~G578_o2;
  assign new_n1191_ = n1828_o2;
  assign new_n1193_ = n801_lo_buf_o2;
  assign new_n1194_ = ~n801_lo_buf_o2;
  assign new_n1196_ = ~G693_o2;
  assign new_n1198_ = ~G702_o2;
  assign new_n1200_ = ~G712_o2;
  assign new_n1202_ = ~G685_o2;
  assign new_n1204_ = ~G658_o2;
  assign new_n1206_ = ~G667_o2;
  assign new_n1208_ = ~G677_o2;
  assign new_n1210_ = ~G650_o2;
  assign new_n1212_ = ~G798_o2;
  assign new_n1213_ = n1017_lo_buf_o2;
  assign new_n1214_ = ~n1017_lo_buf_o2;
  assign new_n1215_ = n1029_lo_buf_o2;
  assign new_n1216_ = ~n1029_lo_buf_o2;
  assign new_n1217_ = n1041_lo_buf_o2;
  assign new_n1218_ = ~n1041_lo_buf_o2;
  assign new_n1219_ = G558_o2;
  assign new_n1221_ = G562_o2;
  assign new_n1223_ = G566_o2;
  assign new_n1225_ = n1835_o2;
  assign new_n1227_ = n1836_o2;
  assign new_n1230_ = ~n1837_o2;
  assign new_n1231_ = n765_lo_buf_o2;
  assign new_n1232_ = ~n765_lo_buf_o2;
  assign new_n1233_ = n777_lo_buf_o2;
  assign new_n1234_ = ~n777_lo_buf_o2;
  assign new_n1235_ = n789_lo_buf_o2;
  assign new_n1236_ = ~n789_lo_buf_o2;
  assign new_n1237_ = G617_o2;
  assign new_n1238_ = ~G617_o2;
  assign new_n1239_ = G626_o2;
  assign new_n1240_ = ~G626_o2;
  assign new_n1241_ = G636_o2;
  assign new_n1242_ = ~G636_o2;
  assign new_n1243_ = n489_lo_buf_o2;
  assign new_n1245_ = n513_lo_buf_o2;
  assign new_n1246_ = ~n513_lo_buf_o2;
  assign new_n1247_ = n561_lo_buf_o2;
  assign new_n1249_ = n597_lo_buf_o2;
  assign new_n1251_ = n657_lo_buf_o2;
  assign new_n1253_ = G276_o2;
  assign new_n1255_ = n1005_lo_buf_o2;
  assign new_n1256_ = ~n1005_lo_buf_o2;
  assign new_n1257_ = n1161_lo_buf_o2;
  assign new_n1258_ = ~n1161_lo_buf_o2;
  assign new_n1259_ = G620_o2;
  assign new_n1260_ = ~G620_o2;
  assign new_n1261_ = G629_o2;
  assign new_n1262_ = ~G629_o2;
  assign new_n1263_ = G639_o2;
  assign new_n1264_ = ~G639_o2;
  assign new_n1265_ = G554_o2;
  assign new_n1267_ = G690_o2;
  assign new_n1269_ = G698_o2;
  assign new_n1270_ = ~G698_o2;
  assign new_n1271_ = G707_o2;
  assign new_n1272_ = ~G707_o2;
  assign new_n1273_ = G319_o2;
  assign new_n1276_ = ~G389_o2;
  assign new_n1277_ = n753_lo_buf_o2;
  assign new_n1278_ = ~n753_lo_buf_o2;
  assign new_n1280_ = ~G647_o2;
  assign new_n1282_ = ~G769_o2;
  assign new_n1284_ = ~G785_o2;
  assign new_n1286_ = ~G808_o2;
  assign new_n1287_ = G445_o2;
  assign new_n1288_ = ~G445_o2;
  assign new_n1289_ = G448_o2;
  assign new_n1290_ = ~G448_o2;
  assign new_n1291_ = G477_o2;
  assign new_n1292_ = ~G477_o2;
  assign new_n1293_ = G480_o2;
  assign new_n1294_ = ~G480_o2;
  assign new_n1296_ = ~G436_o2;
  assign new_n1298_ = ~G786_o2;
  assign new_n1300_ = ~G787_o2;
  assign new_n1302_ = ~G826_o2;
  assign new_n1304_ = ~G827_o2;
  assign new_n1306_ = ~G825_o2;
  assign new_n1307_ = G610_o2;
  assign new_n1308_ = ~G610_o2;
  assign new_n1309_ = n537_lo_buf_o2;
  assign new_n1311_ = n669_lo_buf_o2;
  assign new_n1313_ = n969_lo_buf_o2;
  assign new_n1314_ = ~n969_lo_buf_o2;
  assign new_n1315_ = n981_lo_buf_o2;
  assign new_n1316_ = ~n981_lo_buf_o2;
  assign new_n1317_ = n993_lo_buf_o2;
  assign new_n1318_ = ~n993_lo_buf_o2;
  assign new_n1319_ = G309_o2;
  assign new_n1320_ = ~G309_o2;
  assign new_n1321_ = G461_o2;
  assign new_n1322_ = ~G461_o2;
  assign new_n1323_ = G487_o2;
  assign new_n1324_ = ~G487_o2;
  assign new_n1325_ = G460_o2;
  assign new_n1326_ = ~G460_o2;
  assign new_n1327_ = G468_o2;
  assign new_n1330_ = ~G287_o2;
  assign new_n1331_ = G613_o2;
  assign new_n1332_ = ~G613_o2;
  assign new_n1333_ = n585_lo_buf_o2;
  assign new_n1334_ = ~n585_lo_buf_o2;
  assign new_n1335_ = n813_lo_buf_o2;
  assign new_n1337_ = n825_lo_buf_o2;
  assign new_n1339_ = n837_lo_buf_o2;
  assign new_n1342_ = ~n897_lo_buf_o2;
  assign new_n1344_ = ~n909_lo_buf_o2;
  assign new_n1346_ = ~n933_lo_buf_o2;
  assign new_n1347_ = G451_o2;
  assign new_n1348_ = ~G451_o2;
  assign new_n1349_ = G682_o2;
  assign new_n1350_ = ~G682_o2;
  assign new_n1351_ = G756_o2;
  assign new_n1352_ = ~G756_o2;
  assign new_n1353_ = G542_o2;
  assign new_n1354_ = ~G542_o2;
  assign new_n1355_ = G546_o2;
  assign new_n1356_ = ~G546_o2;
  assign new_n1357_ = G550_o2;
  assign new_n1358_ = ~G550_o2;
  assign new_n1359_ = G310_o2;
  assign new_n1361_ = n798_lo_buf_o2;
  assign new_n1362_ = ~n798_lo_buf_o2;
  assign new_n1364_ = ~n882_lo_buf_o2;
  assign new_n1366_ = ~G427_o2;
  assign new_n1368_ = ~G497_o2;
  assign new_n1370_ = ~G499_o2;
  assign new_n1372_ = ~G501_o2;
  assign new_n1374_ = ~G498_o2;
  assign new_n1376_ = ~G500_o2;
  assign new_n1378_ = ~G502_o2;
  assign new_n1379_ = G369_o2;
  assign new_n1381_ = n939_lo_buf_o2;
  assign new_n1382_ = ~n939_lo_buf_o2;
  assign new_n1383_ = n486_lo_buf_o2;
  assign new_n1385_ = n510_lo_buf_o2;
  assign new_n1386_ = ~n510_lo_buf_o2;
  assign new_n1387_ = n558_lo_buf_o2;
  assign new_n1388_ = ~n558_lo_buf_o2;
  assign new_n1389_ = n594_lo_buf_o2;
  assign new_n1390_ = ~n594_lo_buf_o2;
  assign new_n1391_ = n654_lo_buf_o2;
  assign new_n1392_ = ~n654_lo_buf_o2;
  assign new_n1393_ = n477_lo_buf_o2;
  assign new_n1394_ = ~n477_lo_buf_o2;
  assign new_n1395_ = n525_lo_buf_o2;
  assign new_n1396_ = ~n525_lo_buf_o2;
  assign new_n1397_ = n573_lo_buf_o2;
  assign new_n1398_ = ~n573_lo_buf_o2;
  assign new_n1399_ = new_n866_ | new_n2142_;
  assign new_n1400_ = new_n1399_ | new_n2144_;
  assign new_n1401_ = new_n2145_ | new_n2142_;
  assign new_n1402_ = new_n2146_ | new_n2147_;
  assign new_n1403_ = new_n2146_ | new_n2144_;
  assign new_n1404_ = new_n886_ | new_n878_;
  assign new_n1405_ = new_n806_ | new_n2148_;
  assign new_n1406_ = new_n1405_ | new_n2149_;
  assign new_n1407_ = new_n1406_ | new_n2150_;
  assign new_n1408_ = new_n817_ & new_n803_;
  assign new_n1409_ = new_n818_ | new_n2148_;
  assign new_n1410_ = new_n1408_ & new_n813_;
  assign new_n1411_ = new_n1409_ | new_n2149_;
  assign new_n1412_ = new_n1410_ & new_n815_;
  assign new_n1413_ = new_n1411_ | new_n2150_;
  assign new_n1414_ = new_n1412_ & new_n2152_;
  assign new_n1415_ = new_n865_ & new_n835_;
  assign new_n1416_ = new_n1415_ & new_n869_;
  assign new_n1417_ = new_n2153_ | new_n2145_;
  assign new_n1418_ = new_n2154_ | new_n2147_;
  assign new_n1419_ = new_n2154_ | new_n2143_;
  assign new_n1420_ = new_n901_ | new_n893_;
  assign new_n1421_ = new_n2155_ & new_n917_;
  assign new_n1422_ = new_n1413_ | new_n2152_;
  assign new_n1423_ = new_n2156_ | new_n2141_;
  assign new_n1424_ = new_n1423_ | new_n2157_;
  assign new_n1425_ = new_n2156_ | new_n2153_;
  assign new_n1426_ = new_n1425_ | new_n864_;
  assign new_n1427_ = new_n1426_ | new_n2157_;
  assign new_n1428_ = new_n2155_ & new_n909_;
  assign new_n1429_ = new_n2158_ & new_n2160_;
  assign new_n1430_ = new_n2162_ | new_n2164_;
  assign new_n1431_ = new_n2162_ & new_n2164_;
  assign new_n1432_ = new_n2158_ | new_n2160_;
  assign new_n1433_ = new_n1432_ & new_n1430_;
  assign new_n1434_ = new_n1431_ | new_n1429_;
  assign new_n1435_ = new_n2166_ & new_n2167_;
  assign new_n1436_ = new_n2168_ | new_n2169_;
  assign new_n1437_ = new_n2168_ & new_n2169_;
  assign new_n1438_ = new_n2166_ | new_n2167_;
  assign new_n1439_ = new_n1438_ & new_n1436_;
  assign new_n1440_ = new_n1437_ | new_n1435_;
  assign new_n1441_ = new_n1440_ & new_n1434_;
  assign new_n1442_ = new_n1439_ & new_n1433_;
  assign new_n1443_ = new_n1442_ | new_n1441_;
  assign new_n1444_ = new_n2170_ & new_n2161_;
  assign new_n1445_ = new_n2171_ | new_n2165_;
  assign new_n1446_ = new_n2171_ & new_n2165_;
  assign new_n1447_ = new_n2170_ | new_n2161_;
  assign new_n1448_ = new_n1447_ & new_n1445_;
  assign new_n1449_ = new_n1446_ | new_n1444_;
  assign new_n1450_ = new_n2172_ & new_n2173_;
  assign new_n1451_ = new_n2174_ | new_n2175_;
  assign new_n1452_ = new_n2174_ & new_n2175_;
  assign new_n1453_ = new_n2172_ | new_n2173_;
  assign new_n1454_ = new_n1453_ & new_n1451_;
  assign new_n1455_ = new_n1452_ | new_n1450_;
  assign new_n1456_ = new_n1455_ & new_n1449_;
  assign new_n1457_ = new_n1454_ & new_n1448_;
  assign new_n1458_ = new_n1457_ | new_n1456_;
  assign new_n1459_ = new_n2178_ | new_n954_;
  assign new_n1460_ = new_n1282_ | new_n2185_;
  assign new_n1461_ = new_n1460_ & new_n1459_;
  assign new_n1462_ = new_n1200_ | new_n2192_;
  assign new_n1463_ = new_n1140_ | new_n2199_;
  assign new_n1464_ = new_n1463_ & new_n1462_;
  assign new_n1465_ = new_n1122_ | new_n2205_;
  assign new_n1466_ = new_n1134_ | new_n2208_;
  assign new_n1467_ = new_n1466_ & new_n1465_;
  assign new_n1468_ = new_n2215_ | new_n1038_;
  assign new_n1469_ = new_n1464_ & new_n1461_;
  assign new_n1470_ = new_n1469_ & new_n1467_;
  assign new_n1471_ = new_n1470_ & new_n1468_;
  assign new_n1472_ = new_n2178_ | new_n942_;
  assign new_n1473_ = new_n1284_ | new_n2185_;
  assign new_n1474_ = new_n1473_ & new_n1472_;
  assign new_n1475_ = new_n1202_ | new_n2192_;
  assign new_n1476_ = new_n1144_ | new_n2199_;
  assign new_n1477_ = new_n1476_ & new_n1475_;
  assign new_n1478_ = new_n1142_ | new_n2208_;
  assign new_n1479_ = new_n2215_ | new_n1020_;
  assign new_n1480_ = new_n1479_ & new_n1478_;
  assign new_n1481_ = new_n1477_ & new_n1474_;
  assign new_n1482_ = new_n1481_ & new_n1480_;
  assign new_n1483_ = new_n2179_ | new_n946_;
  assign new_n1484_ = new_n1298_ | new_n2186_;
  assign new_n1485_ = new_n1484_ & new_n1483_;
  assign new_n1486_ = new_n1196_ | new_n2193_;
  assign new_n1487_ = new_n1136_ | new_n2200_;
  assign new_n1488_ = new_n1487_ & new_n1486_;
  assign new_n1489_ = new_n1102_ | new_n2205_;
  assign new_n1490_ = new_n1130_ | new_n2209_;
  assign new_n1491_ = new_n1490_ & new_n1489_;
  assign new_n1492_ = new_n2216_ | new_n1026_;
  assign new_n1493_ = new_n1488_ & new_n1485_;
  assign new_n1494_ = new_n1493_ & new_n1491_;
  assign new_n1495_ = new_n1494_ & new_n1492_;
  assign new_n1496_ = new_n2179_ | new_n950_;
  assign new_n1497_ = new_n1300_ | new_n2186_;
  assign new_n1498_ = new_n1497_ & new_n1496_;
  assign new_n1499_ = new_n1198_ | new_n2193_;
  assign new_n1500_ = new_n1138_ | new_n2200_;
  assign new_n1501_ = new_n1500_ & new_n1499_;
  assign new_n1502_ = new_n1110_ | new_n2204_;
  assign new_n1503_ = new_n1132_ | new_n2209_;
  assign new_n1504_ = new_n1503_ & new_n1502_;
  assign new_n1505_ = new_n2216_ | new_n1032_;
  assign new_n1506_ = new_n1501_ & new_n1498_;
  assign new_n1507_ = new_n1506_ & new_n1504_;
  assign new_n1508_ = new_n1507_ & new_n1505_;
  assign new_n1509_ = new_n1212_ | new_n1190_;
  assign new_n1510_ = new_n1509_ & new_n2220_;
  assign new_n1511_ = new_n2181_ | new_n936_;
  assign new_n1512_ = new_n1286_ | new_n2188_;
  assign new_n1513_ = new_n1512_ & new_n1511_;
  assign new_n1514_ = new_n1208_ | new_n2195_;
  assign new_n1515_ = new_n1174_ | new_n2202_;
  assign new_n1516_ = new_n1515_ & new_n1514_;
  assign new_n1517_ = new_n1150_ | new_n2211_;
  assign new_n1518_ = new_n2218_ | new_n1014_;
  assign new_n1519_ = new_n1518_ & new_n1517_;
  assign new_n1520_ = new_n1516_ & new_n1513_;
  assign new_n1521_ = new_n1520_ & new_n1519_;
  assign new_n1522_ = new_n1128_ | new_n2181_;
  assign new_n1523_ = new_n1306_ | new_n2188_;
  assign new_n1524_ = new_n1523_ & new_n1522_;
  assign new_n1525_ = new_n1210_ | new_n2195_;
  assign new_n1526_ = new_n2220_ | new_n2202_;
  assign new_n1527_ = new_n1526_ & new_n1525_;
  assign new_n1528_ = new_n1176_ | new_n2211_;
  assign new_n1529_ = new_n2218_ | new_n996_;
  assign new_n1530_ = new_n1529_ & new_n1528_;
  assign new_n1531_ = new_n1527_ & new_n1524_;
  assign new_n1532_ = new_n1531_ & new_n1530_;
  assign new_n1533_ = new_n2182_ | new_n924_;
  assign new_n1534_ = new_n1302_ | new_n2189_;
  assign new_n1535_ = new_n1534_ & new_n1533_;
  assign new_n1536_ = new_n1204_ | new_n2196_;
  assign new_n1537_ = new_n1170_ | new_n2203_;
  assign new_n1538_ = new_n1537_ & new_n1536_;
  assign new_n1539_ = new_n1148_ | new_n2212_;
  assign new_n1540_ = new_n2219_ | new_n1002_;
  assign new_n1541_ = new_n1540_ & new_n1539_;
  assign new_n1542_ = new_n1538_ & new_n1535_;
  assign new_n1543_ = new_n1542_ & new_n1541_;
  assign new_n1544_ = new_n2182_ | new_n930_;
  assign new_n1545_ = new_n1304_ | new_n2189_;
  assign new_n1546_ = new_n1545_ & new_n1544_;
  assign new_n1547_ = new_n1206_ | new_n2196_;
  assign new_n1548_ = new_n1172_ | new_n2203_;
  assign new_n1549_ = new_n1548_ & new_n1547_;
  assign new_n1550_ = new_n1146_ | new_n2212_;
  assign new_n1551_ = new_n2219_ | new_n1008_;
  assign new_n1552_ = new_n1551_ & new_n1550_;
  assign new_n1553_ = new_n1549_ & new_n1546_;
  assign new_n1554_ = new_n1553_ & new_n1552_;
  assign new_n1555_ = new_n1156_ | new_n1152_;
  assign new_n1556_ = new_n1555_ | new_n812_;
  assign new_n1557_ = new_n1556_ | new_n1182_;
  assign new_n1558_ = new_n2222_ & new_n2225_;
  assign new_n1559_ = new_n2227_ | new_n2229_;
  assign new_n1560_ = new_n2232_ & new_n2235_;
  assign new_n1561_ = new_n2237_ | new_n2239_;
  assign new_n1562_ = new_n2242_ & new_n2245_;
  assign new_n1563_ = new_n2247_ | new_n2249_;
  assign new_n1564_ = new_n1324_ & new_n1320_;
  assign new_n1565_ = new_n1323_ | new_n1319_;
  assign new_n1566_ = new_n1326_ & new_n1322_;
  assign new_n1567_ = new_n1325_ | new_n1321_;
  assign new_n1568_ = new_n1566_ & new_n1564_;
  assign new_n1569_ = new_n1567_ | new_n1565_;
  assign new_n1570_ = new_n2251_ & new_n2253_;
  assign new_n1571_ = new_n2256_ | new_n2259_;
  assign new_n1572_ = new_n1259_ & new_n1238_;
  assign new_n1573_ = new_n1260_ | new_n1237_;
  assign new_n1574_ = new_n2262_ & new_n1240_;
  assign new_n1575_ = new_n2264_ | new_n1239_;
  assign new_n1576_ = new_n2266_ & new_n1242_;
  assign new_n1577_ = new_n2268_ | new_n1241_;
  assign new_n1578_ = new_n2269_ & new_n1308_;
  assign new_n1579_ = new_n2270_ | new_n1307_;
  assign new_n1580_ = new_n2227_ & new_n2229_;
  assign new_n1581_ = new_n2222_ | new_n2225_;
  assign new_n1582_ = new_n2272_ & new_n2273_;
  assign new_n1583_ = new_n2275_ | new_n2277_;
  assign new_n1584_ = new_n2237_ & new_n2239_;
  assign new_n1585_ = new_n2232_ | new_n2235_;
  assign new_n1586_ = new_n2279_ & new_n2282_;
  assign new_n1587_ = new_n2284_ | new_n2287_;
  assign new_n1588_ = new_n2247_ & new_n2249_;
  assign new_n1589_ = new_n2242_ | new_n2245_;
  assign new_n1590_ = new_n2290_ & new_n2293_;
  assign new_n1591_ = new_n2296_ | new_n2300_;
  assign new_n1592_ = new_n2256_ & new_n2259_;
  assign new_n1593_ = new_n2251_ | new_n2253_;
  assign new_n1594_ = new_n1593_ & new_n2302_;
  assign new_n1595_ = new_n2303_ | new_n1570_;
  assign new_n1596_ = new_n2272_ & new_n2287_;
  assign new_n1597_ = new_n2275_ | new_n2282_;
  assign new_n1598_ = new_n2279_ & new_n2271_;
  assign new_n1599_ = new_n2284_ | new_n2274_;
  assign new_n1600_ = new_n2304_ & new_n2300_;
  assign new_n1601_ = new_n2305_ | new_n2293_;
  assign new_n1602_ = new_n2306_ & new_n2269_;
  assign new_n1603_ = new_n2307_ | new_n2270_;
  assign new_n1604_ = new_n1603_ & new_n1350_;
  assign new_n1605_ = new_n1602_ | new_n2308_;
  assign new_n1606_ = new_n2304_ & new_n2290_;
  assign new_n1607_ = new_n2305_ | new_n2296_;
  assign new_n1608_ = new_n1606_ & new_n2310_;
  assign new_n1609_ = new_n1607_ | new_n2313_;
  assign new_n1610_ = new_n1597_ & new_n2273_;
  assign new_n1611_ = new_n1596_ | new_n2277_;
  assign new_n1612_ = new_n1610_ & new_n1601_;
  assign new_n1613_ = new_n1611_ | new_n1600_;
  assign new_n1614_ = new_n1612_ & new_n1609_;
  assign new_n1615_ = new_n1613_ | new_n1608_;
  assign new_n1616_ = new_n2315_ | new_n1366_;
  assign new_n1617_ = new_n1374_ & new_n1368_;
  assign new_n1618_ = new_n1617_ & new_n2317_;
  assign new_n1619_ = new_n1376_ & new_n1370_;
  assign new_n1620_ = new_n1619_ & new_n2317_;
  assign new_n1621_ = new_n1378_ & new_n1372_;
  assign new_n1622_ = new_n1621_ & new_n2318_;
  assign new_n1623_ = new_n2320_ | new_n2321_;
  assign new_n1624_ = new_n2323_ | new_n2324_;
  assign new_n1625_ = new_n2326_ | new_n2327_;
  assign new_n1626_ = new_n2328_ & new_n2330_;
  assign new_n1627_ = new_n1396_ | new_n2331_;
  assign new_n1628_ = new_n1626_ & new_n2333_;
  assign new_n1629_ = new_n1627_ | new_n1398_;
  assign new_n1630_ = new_n2320_ & new_n2321_;
  assign new_n1631_ = new_n2323_ & new_n2324_;
  assign new_n1632_ = new_n2326_ & new_n2327_;
  assign new_n1633_ = new_n2334_ | new_n1327_;
  assign new_n1634_ = new_n1362_ | new_n2336_;
  assign new_n1635_ = new_n1634_ & new_n1633_;
  assign new_n1636_ = new_n1635_ & new_n2318_;
  assign new_n1637_ = new_n2338_ | new_n1382_;
  assign new_n1638_ = new_n2339_ | new_n2341_;
  assign new_n1639_ = new_n1577_ | new_n2343_;
  assign new_n1640_ = new_n1639_ & new_n1638_;
  assign new_n1641_ = new_n2344_ | new_n2306_;
  assign new_n1642_ = new_n1579_ | new_n2307_;
  assign new_n1643_ = new_n1642_ & new_n1641_;
  assign new_n1644_ = new_n2310_ | new_n2345_;
  assign new_n1645_ = new_n2313_ | new_n1591_;
  assign new_n1646_ = new_n1645_ & new_n1644_;
  assign new_n1647_ = new_n2347_ & new_n2349_;
  assign new_n1648_ = new_n2350_ | new_n2351_;
  assign new_n1649_ = new_n2350_ & new_n2351_;
  assign new_n1650_ = new_n2347_ | new_n2349_;
  assign new_n1651_ = new_n1650_ & new_n1648_;
  assign new_n1652_ = new_n1649_ | new_n1647_;
  assign new_n1653_ = new_n2353_ & new_n2355_;
  assign new_n1654_ = new_n2356_ | new_n2357_;
  assign new_n1655_ = new_n2356_ & new_n2357_;
  assign new_n1656_ = new_n2353_ | new_n2355_;
  assign new_n1657_ = new_n1656_ & new_n1654_;
  assign new_n1658_ = new_n1655_ | new_n1653_;
  assign new_n1659_ = new_n1657_ | new_n1651_;
  assign new_n1660_ = new_n1658_ | new_n1652_;
  assign new_n1661_ = new_n1660_ & new_n1659_;
  assign new_n1662_ = new_n2359_ & new_n2361_;
  assign new_n1663_ = new_n2362_ | new_n2363_;
  assign new_n1664_ = new_n2362_ & new_n2363_;
  assign new_n1665_ = new_n2359_ | new_n2361_;
  assign new_n1666_ = new_n1665_ & new_n1663_;
  assign new_n1667_ = new_n1664_ | new_n1662_;
  assign new_n1668_ = new_n2364_ & new_n2366_;
  assign new_n1669_ = new_n2367_ | new_n2368_;
  assign new_n1670_ = new_n2367_ & new_n2368_;
  assign new_n1671_ = new_n2364_ | new_n2366_;
  assign new_n1672_ = new_n1671_ & new_n1669_;
  assign new_n1673_ = new_n1670_ | new_n1668_;
  assign new_n1674_ = new_n1672_ | new_n1666_;
  assign new_n1675_ = new_n1673_ | new_n1667_;
  assign new_n1676_ = new_n1675_ & new_n1674_;
  assign new_n1677_ = new_n2224_ & new_n2258_;
  assign new_n1678_ = new_n2230_ | new_n2254_;
  assign new_n1679_ = new_n2230_ & new_n2254_;
  assign new_n1680_ = new_n2226_ | new_n2260_;
  assign new_n1681_ = new_n1680_ & new_n1678_;
  assign new_n1682_ = new_n1679_ | new_n1677_;
  assign new_n1683_ = new_n2244_ & new_n2234_;
  assign new_n1684_ = new_n2250_ | new_n2240_;
  assign new_n1685_ = new_n2250_ & new_n2240_;
  assign new_n1686_ = new_n2246_ | new_n2236_;
  assign new_n1687_ = new_n1686_ & new_n1684_;
  assign new_n1688_ = new_n1685_ | new_n1683_;
  assign new_n1689_ = new_n1687_ | new_n1681_;
  assign new_n1690_ = new_n1688_ | new_n1682_;
  assign new_n1691_ = new_n1690_ & new_n1689_;
  assign new_n1692_ = new_n2370_ & new_n2372_;
  assign new_n1693_ = new_n2373_ | new_n2374_;
  assign new_n1694_ = new_n2373_ & new_n2374_;
  assign new_n1695_ = new_n2370_ | new_n2372_;
  assign new_n1696_ = new_n1695_ & new_n1693_;
  assign new_n1697_ = new_n1694_ | new_n1692_;
  assign new_n1698_ = new_n2376_ & new_n2378_;
  assign new_n1699_ = new_n2379_ | new_n2380_;
  assign new_n1700_ = new_n2379_ & new_n2380_;
  assign new_n1701_ = new_n2376_ | new_n2378_;
  assign new_n1702_ = new_n1701_ & new_n1699_;
  assign new_n1703_ = new_n1700_ | new_n1698_;
  assign new_n1704_ = new_n1702_ | new_n1696_;
  assign new_n1705_ = new_n1703_ | new_n1697_;
  assign new_n1706_ = new_n1705_ & new_n1704_;
  assign new_n1707_ = new_n1162_ | new_n1160_;
  assign new_n1708_ = new_n1707_ | new_n842_;
  assign new_n1709_ = new_n1708_ | new_n850_;
  assign new_n1710_ = new_n1709_ | new_n2381_;
  assign new_n1711_ = new_n1710_ | new_n856_;
  assign new_n1712_ = new_n2383_ & new_n2262_;
  assign new_n1713_ = new_n2384_ | new_n2264_;
  assign new_n1714_ = new_n2266_ & new_n2261_;
  assign new_n1715_ = new_n2268_ | new_n2263_;
  assign new_n1716_ = new_n1714_ & new_n2341_;
  assign new_n1717_ = new_n1715_ | new_n2343_;
  assign new_n1718_ = new_n1713_ & new_n1270_;
  assign new_n1719_ = new_n1712_ | new_n2385_;
  assign new_n1720_ = new_n1718_ & new_n1717_;
  assign new_n1721_ = new_n1719_ | new_n1716_;
  assign new_n1722_ = new_n1721_ | new_n2386_;
  assign new_n1723_ = new_n1720_ | new_n1573_;
  assign new_n1724_ = new_n1723_ & new_n1722_;
  assign new_n1725_ = new_n2265_ & new_n2340_;
  assign new_n1726_ = new_n2267_ | new_n2342_;
  assign new_n1727_ = new_n1726_ & new_n2384_;
  assign new_n1728_ = new_n1725_ | new_n2383_;
  assign new_n1729_ = new_n1728_ | new_n2387_;
  assign new_n1730_ = new_n1727_ | new_n1575_;
  assign new_n1731_ = new_n1730_ & new_n1729_;
  assign new_n1732_ = new_n2280_ & new_n2299_;
  assign new_n1733_ = new_n2285_ | new_n2294_;
  assign new_n1734_ = new_n2291_ & new_n2280_;
  assign new_n1735_ = new_n2297_ | new_n2285_;
  assign new_n1736_ = new_n1734_ & new_n2311_;
  assign new_n1737_ = new_n1735_ | new_n2314_;
  assign new_n1738_ = new_n1733_ & new_n2281_;
  assign new_n1739_ = new_n1732_ | new_n2288_;
  assign new_n1740_ = new_n1738_ & new_n1737_;
  assign new_n1741_ = new_n1739_ | new_n1736_;
  assign new_n1742_ = new_n1741_ | new_n2388_;
  assign new_n1743_ = new_n1740_ | new_n1583_;
  assign new_n1744_ = new_n1743_ & new_n1742_;
  assign new_n1745_ = new_n2311_ & new_n2291_;
  assign new_n1746_ = new_n2314_ | new_n2297_;
  assign new_n1747_ = new_n1746_ & new_n2294_;
  assign new_n1748_ = new_n1745_ | new_n2301_;
  assign new_n1749_ = new_n1748_ | new_n2389_;
  assign new_n1750_ = new_n1747_ | new_n1587_;
  assign new_n1751_ = new_n1750_ & new_n1749_;
  assign new_n1752_ = new_n2390_ | new_n2391_;
  assign new_n1753_ = new_n1614_ | new_n1595_;
  assign new_n1754_ = new_n1753_ & new_n1752_;
  assign new_n1755_ = new_n2393_ | new_n2394_;
  assign new_n1756_ = new_n2395_ & new_n975_;
  assign new_n1757_ = new_n2396_ | new_n2397_;
  assign new_n1758_ = new_n1757_ | new_n1330_;
  assign new_n1759_ = new_n1758_ | new_n1359_;
  assign new_n1760_ = new_n1347_ & new_n2398_;
  assign new_n1761_ = new_n2396_ | new_n1273_;
  assign new_n1762_ = new_n1761_ | new_n1334_;
  assign new_n1763_ = new_n2400_ | new_n2334_;
  assign new_n1764_ = new_n2402_ & new_n2404_;
  assign new_n1765_ = new_n1764_ & new_n2407_;
  assign new_n1766_ = new_n1765_ | new_n2331_;
  assign new_n1767_ = new_n2409_ | new_n820_;
  assign new_n1768_ = new_n1767_ | new_n868_;
  assign new_n1769_ = new_n2393_ & new_n2394_;
  assign new_n1770_ = new_n2410_ | new_n2407_;
  assign new_n1771_ = new_n2411_ | new_n1386_;
  assign new_n1772_ = new_n1771_ & new_n1770_;
  assign new_n1773_ = new_n1772_ & new_n2412_;
  assign new_n1774_ = new_n1773_ & new_n1381_;
  assign new_n1775_ = new_n1774_ & new_n2404_;
  assign new_n1776_ = new_n2330_ & new_n2413_;
  assign new_n1777_ = new_n1776_ & new_n2333_;
  assign new_n1778_ = new_n1777_ & new_n2408_;
  assign new_n1779_ = new_n2409_ | new_n2338_;
  assign new_n1780_ = new_n1779_ | new_n2411_;
  assign new_n1781_ = new_n1780_ & new_n1778_;
  assign new_n1782_ = new_n1781_ | new_n1775_;
  assign new_n1783_ = new_n2415_ | new_n2417_;
  assign new_n1784_ = new_n2418_ | new_n2415_;
  assign new_n1785_ = new_n2419_ | new_n2421_;
  assign new_n1786_ = new_n2419_ | new_n2422_;
  assign new_n1787_ = new_n1786_ | new_n1114_;
  assign new_n1788_ = new_n1783_ & new_n2424_;
  assign new_n1789_ = new_n1788_ & new_n1785_;
  assign new_n1790_ = new_n1789_ & new_n1787_;
  assign new_n1791_ = new_n1230_ | new_n2426_;
  assign new_n1792_ = new_n2336_ | new_n928_;
  assign new_n1793_ = new_n1792_ & new_n1791_;
  assign new_n1794_ = new_n2400_ | new_n1342_;
  assign new_n1795_ = new_n1794_ & new_n2428_;
  assign new_n1796_ = new_n1795_ & new_n1793_;
  assign new_n1797_ = new_n2397_ | new_n2426_;
  assign new_n1798_ = new_n2337_ | new_n934_;
  assign new_n1799_ = new_n1798_ & new_n1797_;
  assign new_n1800_ = new_n2401_ | new_n1344_;
  assign new_n1801_ = new_n1800_ & new_n2428_;
  assign new_n1802_ = new_n1801_ & new_n1799_;
  assign new_n1803_ = new_n986_ | new_n2425_;
  assign new_n1804_ = new_n2337_ | new_n940_;
  assign new_n1805_ = new_n1804_ & new_n1803_;
  assign new_n1806_ = new_n2401_ | new_n1346_;
  assign new_n1807_ = new_n1806_ & new_n2429_;
  assign new_n1808_ = new_n1807_ & new_n1805_;
  assign new_n1809_ = new_n2430_ | new_n1629_;
  assign new_n1810_ = new_n1809_ | new_n834_;
  assign new_n1811_ = new_n2432_ & new_n2434_;
  assign new_n1812_ = new_n2432_ & new_n2435_;
  assign new_n1813_ = new_n2433_ & new_n2436_;
  assign new_n1814_ = new_n2438_ & new_n2440_;
  assign new_n1815_ = new_n2438_ & new_n2441_;
  assign new_n1816_ = new_n2439_ & new_n2442_;
  assign G855 = new_n1400_;
  assign G856 = new_n1402_;
  assign G857 = new_n2151_;
  assign G858 = new_n1404_;
  assign G859 = new_n1407_;
  assign G860 = new_n1414_;
  assign G861 = new_n1416_;
  assign G862 = ~new_n1418_;
  assign G863 = ~new_n1419_;
  assign G864 = ~new_n1421_;
  assign G865 = ~new_n1422_;
  assign G866 = new_n1126_;
  assign G867 = new_n1424_;
  assign G868 = new_n1427_;
  assign G869 = ~new_n1428_;
  assign G870 = new_n1443_;
  assign G871 = new_n1458_;
  assign G872 = new_n1471_;
  assign G873 = new_n1482_;
  assign G874 = new_n1495_;
  assign G875 = new_n1508_;
  assign G876 = new_n1510_;
  assign G877 = new_n1521_;
  assign G878 = new_n1532_;
  assign G879 = new_n1543_;
  assign G880 = new_n1554_;
  assign n480_li = new_n1151_;
  assign n492_li = new_n1155_;
  assign n495_li = new_n687_;
  assign n498_li = new_n807_;
  assign n501_li = new_n809_;
  assign n504_li = new_n811_;
  assign n516_li = new_n1157_;
  assign n528_li = new_n1153_;
  assign n531_li = new_n693_;
  assign n540_li = new_n1177_;
  assign n543_li = new_n695_;
  assign n546_li = new_n823_;
  assign n549_li = new_n825_;
  assign n552_li = new_n827_;
  assign n564_li = new_n1159_;
  assign n579_li = new_n701_;
  assign n600_li = new_n1161_;
  assign n603_li = new_n705_;
  assign n606_li = new_n837_;
  assign n609_li = new_n839_;
  assign n612_li = new_n841_;
  assign n615_li = new_n707_;
  assign n618_li = new_n845_;
  assign n621_li = new_n847_;
  assign n627_li = new_n709_;
  assign n630_li = new_n851_;
  assign n633_li = new_n853_;
  assign n639_li = new_n711_;
  assign n642_li = new_n857_;
  assign n645_li = new_n859_;
  assign n648_li = new_n861_;
  assign n660_li = new_n1163_;
  assign n663_li = new_n715_;
  assign n672_li = new_n1179_;
  assign n675_li = new_n717_;
  assign n678_li = new_n871_;
  assign n681_li = new_n873_;
  assign n684_li = new_n875_;
  assign n687_li = new_n719_;
  assign n690_li = new_n879_;
  assign n693_li = new_n881_;
  assign n696_li = new_n883_;
  assign n699_li = new_n721_;
  assign n702_li = new_n887_;
  assign n705_li = new_n889_;
  assign n708_li = new_n891_;
  assign n711_li = new_n723_;
  assign n714_li = new_n895_;
  assign n717_li = new_n897_;
  assign n720_li = new_n899_;
  assign n723_li = new_n725_;
  assign n726_li = new_n903_;
  assign n729_li = new_n905_;
  assign n732_li = new_n907_;
  assign n735_li = new_n727_;
  assign n738_li = new_n911_;
  assign n741_li = new_n913_;
  assign n744_li = new_n915_;
  assign n747_li = new_n729_;
  assign n750_li = new_n919_;
  assign n756_li = new_n2346_;
  assign n759_li = new_n731_;
  assign n762_li = new_n925_;
  assign n768_li = new_n2348_;
  assign n771_li = new_n733_;
  assign n774_li = new_n931_;
  assign n780_li = new_n2354_;
  assign n783_li = new_n735_;
  assign n786_li = new_n937_;
  assign n792_li = new_n2352_;
  assign n795_li = new_n737_;
  assign n804_li = new_n2358_;
  assign n807_li = new_n739_;
  assign n816_li = new_n2360_;
  assign n819_li = new_n741_;
  assign n828_li = new_n2365_;
  assign n831_li = new_n743_;
  assign n843_li = new_n745_;
  assign n846_li = new_n957_;
  assign n849_li = new_n959_;
  assign n852_li = new_n961_;
  assign n855_li = new_n747_;
  assign n858_li = new_n965_;
  assign n861_li = new_n967_;
  assign n864_li = new_n969_;
  assign n867_li = new_n749_;
  assign n870_li = new_n973_;
  assign n879_li = new_n751_;
  assign n891_li = new_n753_;
  assign n903_li = new_n755_;
  assign n915_li = new_n757_;
  assign n918_li = new_n983_;
  assign n927_li = new_n759_;
  assign n951_li = new_n763_;
  assign n954_li = new_n989_;
  assign n957_li = new_n991_;
  assign n960_li = new_n2260_;
  assign n963_li = new_n765_;
  assign n966_li = new_n997_;
  assign n972_li = new_n2226_;
  assign n975_li = new_n767_;
  assign n978_li = new_n1003_;
  assign n984_li = new_n2236_;
  assign n987_li = new_n769_;
  assign n990_li = new_n1009_;
  assign n996_li = new_n2246_;
  assign n999_li = new_n771_;
  assign n1002_li = new_n1015_;
  assign n1008_li = new_n2369_;
  assign n1011_li = new_n773_;
  assign n1014_li = new_n1021_;
  assign n1020_li = new_n2371_;
  assign n1023_li = new_n775_;
  assign n1026_li = new_n1027_;
  assign n1032_li = new_n2377_;
  assign n1035_li = new_n777_;
  assign n1038_li = new_n1033_;
  assign n1044_li = new_n2375_;
  assign n1047_li = new_n779_;
  assign n1050_li = new_n1039_;
  assign n1053_li = new_n1041_;
  assign n1056_li = new_n1043_;
  assign n1059_li = new_n781_;
  assign n1062_li = new_n1047_;
  assign n1065_li = new_n1049_;
  assign n1068_li = new_n1051_;
  assign n1071_li = new_n783_;
  assign n1074_li = new_n1055_;
  assign n1077_li = new_n1057_;
  assign n1080_li = new_n1059_;
  assign n1083_li = new_n785_;
  assign n1086_li = new_n1063_;
  assign n1089_li = new_n1065_;
  assign n1092_li = new_n1067_;
  assign n1095_li = new_n787_;
  assign n1098_li = new_n1071_;
  assign n1101_li = new_n1073_;
  assign n1104_li = new_n1075_;
  assign n1107_li = new_n789_;
  assign n1110_li = new_n1079_;
  assign n1113_li = new_n1081_;
  assign n1116_li = new_n1083_;
  assign n1119_li = new_n791_;
  assign n1122_li = new_n1087_;
  assign n1125_li = new_n1089_;
  assign n1128_li = new_n1091_;
  assign n1131_li = new_n793_;
  assign n1134_li = new_n1095_;
  assign n1137_li = new_n1097_;
  assign n1140_li = new_n1099_;
  assign n1143_li = new_n795_;
  assign n1146_li = new_n1103_;
  assign n1149_li = new_n1105_;
  assign n1152_li = new_n1107_;
  assign n1155_li = new_n797_;
  assign n1158_li = new_n1111_;
  assign n1167_li = new_n799_;
  assign n1170_li = new_n1115_;
  assign n1173_li = new_n1117_;
  assign n1176_li = new_n1119_;
  assign n1179_li = new_n801_;
  assign n1529_i2 = new_n1165_;
  assign n1616_i2 = new_n1191_;
  assign n1655_i2 = new_n1219_;
  assign n1656_i2 = new_n1221_;
  assign n1657_i2 = new_n1223_;
  assign n1730_i2 = new_n1267_;
  assign n1731_i2 = new_n2385_;
  assign n1732_i2 = new_n2382_;
  assign n1729_i2 = new_n1265_;
  assign n1805_i2 = new_n2308_;
  assign n1808_i2 = new_n2231_;
  assign n1807_i2 = new_n2221_;
  assign n1809_i2 = new_n2241_;
  assign n1663_i2 = new_n1225_;
  assign n1664_i2 = new_n1227_;
  assign n1704_i2 = new_n2395_;
  assign n1705_i2 = new_n1245_;
  assign n1706_i2 = new_n1247_;
  assign n1707_i2 = new_n1249_;
  assign n1708_i2 = new_n1251_;
  assign n1709_i2 = new_n1253_;
  assign G280_i2 = ~new_n2381_;
  assign G655_i2 = new_n2276_;
  assign G663_i2 = new_n2288_;
  assign G672_i2 = new_n2301_;
  assign G538_i2 = new_n2255_;
  assign n1780_i2 = new_n1309_;
  assign n1781_i2 = new_n1311_;
  assign n1797_i2 = new_n1333_;
  assign n1798_i2 = new_n1335_;
  assign n1799_i2 = new_n1337_;
  assign n1800_i2 = new_n1339_;
  assign G578_i2 = new_n2302_;
  assign n1828_i2 = new_n2315_;
  assign n801_lo_buf_i2 = new_n1361_;
  assign G693_i2 = new_n2386_;
  assign G702_i2 = new_n2387_;
  assign G712_i2 = new_n2339_;
  assign G685_i2 = new_n2344_;
  assign G658_i2 = new_n2388_;
  assign G667_i2 = new_n2389_;
  assign G677_i2 = new_n2345_;
  assign G650_i2 = new_n2391_;
  assign G798_i2 = new_n2390_;
  assign n1017_lo_buf_i2 = new_n1023_;
  assign n1029_lo_buf_i2 = new_n1029_;
  assign n1041_lo_buf_i2 = new_n1035_;
  assign G558_i2 = ~new_n2319_;
  assign G562_i2 = ~new_n2322_;
  assign G566_i2 = ~new_n2325_;
  assign n1835_i2 = new_n2329_;
  assign n1836_i2 = new_n2328_;
  assign n1837_i2 = new_n2332_;
  assign n765_lo_buf_i2 = new_n927_;
  assign n777_lo_buf_i2 = new_n933_;
  assign n789_lo_buf_i2 = new_n939_;
  assign G617_i2 = ~new_n2424_;
  assign G626_i2 = ~new_n2417_;
  assign G636_i2 = ~new_n2421_;
  assign n489_lo_buf_i2 = new_n2413_;
  assign n513_lo_buf_i2 = new_n2408_;
  assign n561_lo_buf_i2 = new_n2410_;
  assign n597_lo_buf_i2 = new_n2412_;
  assign n657_lo_buf_i2 = new_n1391_;
  assign G276_i2 = new_n2405_;
  assign n1005_lo_buf_i2 = new_n1017_;
  assign n1161_lo_buf_i2 = new_n1113_;
  assign G620_i2 = ~new_n2414_;
  assign G629_i2 = ~new_n2418_;
  assign G639_i2 = ~new_n2422_;
  assign G554_i2 = ~new_n2392_;
  assign G690_i2 = ~new_n2423_;
  assign G698_i2 = ~new_n2416_;
  assign G707_i2 = ~new_n2420_;
  assign G319_i2 = ~new_n2402_;
  assign G389_i2 = G276_i2;
  assign n753_lo_buf_i2 = new_n2398_;
  assign G647_i2 = new_n2303_;
  assign G769_i2 = new_n1640_;
  assign G785_i2 = new_n1643_;
  assign G808_i2 = new_n1646_;
  assign G445_i2 = new_n1661_;
  assign G448_i2 = new_n1676_;
  assign G477_i2 = new_n1691_;
  assign G480_i2 = new_n1706_;
  assign G436_i2 = ~new_n1711_;
  assign G786_i2 = new_n1724_;
  assign G787_i2 = new_n1731_;
  assign G826_i2 = new_n1744_;
  assign G827_i2 = new_n1751_;
  assign G825_i2 = new_n1754_;
  assign G610_i2 = ~new_n2443_;
  assign n537_lo_buf_i2 = new_n819_;
  assign n669_lo_buf_i2 = new_n867_;
  assign n969_lo_buf_i2 = new_n999_;
  assign n981_lo_buf_i2 = new_n1005_;
  assign n993_lo_buf_i2 = new_n1011_;
  assign G309_i2 = new_n1756_;
  assign G461_i2 = ~new_n2429_;
  assign G487_i2 = new_n1760_;
  assign G460_i2 = ~new_n1763_;
  assign G468_i2 = ~new_n2433_;
  assign G287_i2 = ~new_n2430_;
  assign G613_i2 = ~new_n1769_;
  assign n585_lo_buf_i2 = new_n833_;
  assign n813_lo_buf_i2 = new_n2440_;
  assign n825_lo_buf_i2 = new_n2441_;
  assign n837_lo_buf_i2 = new_n2442_;
  assign n897_lo_buf_i2 = new_n2434_;
  assign n909_lo_buf_i2 = new_n2435_;
  assign n933_lo_buf_i2 = new_n2436_;
  assign G451_i2 = new_n2439_;
  assign G682_i2 = G610_i2;
  assign G756_i2 = ~new_n1790_;
  assign G542_i2 = ~new_n1796_;
  assign G546_i2 = ~new_n1802_;
  assign G550_i2 = ~new_n1808_;
  assign G310_i2 = new_n2444_;
  assign n798_lo_buf_i2 = new_n943_;
  assign n882_lo_buf_i2 = new_n977_;
  assign G427_i2 = ~new_n1810_;
  assign G497_i2 = new_n1811_;
  assign G499_i2 = new_n1812_;
  assign G501_i2 = new_n1813_;
  assign G498_i2 = new_n1814_;
  assign G500_i2 = new_n1815_;
  assign G502_i2 = new_n1816_;
  assign G369_i2 = G310_i2;
  assign n939_lo_buf_i2 = new_n761_;
  assign n486_lo_buf_i2 = new_n685_;
  assign n510_lo_buf_i2 = new_n689_;
  assign n558_lo_buf_i2 = new_n697_;
  assign n594_lo_buf_i2 = new_n703_;
  assign n654_lo_buf_i2 = new_n713_;
  assign n477_lo_buf_i2 = new_n683_;
  assign n525_lo_buf_i2 = new_n691_;
  assign n573_lo_buf_i2 = new_n699_;
  assign new_n2141_ = new_n822_;
  assign new_n2142_ = new_n2141_;
  assign new_n2143_ = new_n832_;
  assign new_n2144_ = new_n2143_;
  assign new_n2145_ = new_n830_;
  assign new_n2146_ = new_n1401_;
  assign new_n2147_ = new_n870_;
  assign new_n2148_ = new_n804_;
  assign new_n2149_ = new_n814_;
  assign new_n2150_ = new_n816_;
  assign new_n2151_ = new_n1403_;
  assign new_n2152_ = new_n2151_;
  assign new_n2153_ = new_n836_;
  assign new_n2154_ = new_n1417_;
  assign new_n2155_ = new_n1420_;
  assign new_n2156_ = new_n844_;
  assign new_n2157_ = new_n1168_;
  assign new_n2158_ = new_n1287_;
  assign new_n2159_ = new_n963_;
  assign new_n2160_ = new_n2159_;
  assign new_n2161_ = new_n2159_;
  assign new_n2162_ = new_n1288_;
  assign new_n2163_ = new_n964_;
  assign new_n2164_ = new_n2163_;
  assign new_n2165_ = new_n2163_;
  assign new_n2166_ = new_n1289_;
  assign new_n2167_ = new_n971_;
  assign new_n2168_ = new_n1290_;
  assign new_n2169_ = new_n972_;
  assign new_n2170_ = new_n1291_;
  assign new_n2171_ = new_n1292_;
  assign new_n2172_ = new_n1293_;
  assign new_n2173_ = new_n1045_;
  assign new_n2174_ = new_n1294_;
  assign new_n2175_ = new_n1046_;
  assign new_n2176_ = new_n1054_;
  assign new_n2177_ = new_n2176_;
  assign new_n2178_ = new_n2177_;
  assign new_n2179_ = new_n2177_;
  assign new_n2180_ = new_n2176_;
  assign new_n2181_ = new_n2180_;
  assign new_n2182_ = new_n2180_;
  assign new_n2183_ = new_n1062_;
  assign new_n2184_ = new_n2183_;
  assign new_n2185_ = new_n2184_;
  assign new_n2186_ = new_n2184_;
  assign new_n2187_ = new_n2183_;
  assign new_n2188_ = new_n2187_;
  assign new_n2189_ = new_n2187_;
  assign new_n2190_ = new_n1070_;
  assign new_n2191_ = new_n2190_;
  assign new_n2192_ = new_n2191_;
  assign new_n2193_ = new_n2191_;
  assign new_n2194_ = new_n2190_;
  assign new_n2195_ = new_n2194_;
  assign new_n2196_ = new_n2194_;
  assign new_n2197_ = new_n1078_;
  assign new_n2198_ = new_n2197_;
  assign new_n2199_ = new_n2198_;
  assign new_n2200_ = new_n2198_;
  assign new_n2201_ = new_n2197_;
  assign new_n2202_ = new_n2201_;
  assign new_n2203_ = new_n2201_;
  assign new_n2204_ = new_n1094_;
  assign new_n2205_ = new_n2204_;
  assign new_n2206_ = new_n1086_;
  assign new_n2207_ = new_n2206_;
  assign new_n2208_ = new_n2207_;
  assign new_n2209_ = new_n2207_;
  assign new_n2210_ = new_n2206_;
  assign new_n2211_ = new_n2210_;
  assign new_n2212_ = new_n2210_;
  assign new_n2213_ = new_n1296_;
  assign new_n2214_ = new_n2213_;
  assign new_n2215_ = new_n2214_;
  assign new_n2216_ = new_n2214_;
  assign new_n2217_ = new_n2213_;
  assign new_n2218_ = new_n2217_;
  assign new_n2219_ = new_n2217_;
  assign new_n2220_ = new_n1280_;
  assign new_n2221_ = new_n1353_;
  assign new_n2222_ = new_n2221_;
  assign new_n2223_ = new_n1313_;
  assign new_n2224_ = new_n2223_;
  assign new_n2225_ = new_n2224_;
  assign new_n2226_ = new_n2223_;
  assign new_n2227_ = new_n1354_;
  assign new_n2228_ = new_n1314_;
  assign new_n2229_ = new_n2228_;
  assign new_n2230_ = new_n2228_;
  assign new_n2231_ = new_n1355_;
  assign new_n2232_ = new_n2231_;
  assign new_n2233_ = new_n1315_;
  assign new_n2234_ = new_n2233_;
  assign new_n2235_ = new_n2234_;
  assign new_n2236_ = new_n2233_;
  assign new_n2237_ = new_n1356_;
  assign new_n2238_ = new_n1316_;
  assign new_n2239_ = new_n2238_;
  assign new_n2240_ = new_n2238_;
  assign new_n2241_ = new_n1357_;
  assign new_n2242_ = new_n2241_;
  assign new_n2243_ = new_n1317_;
  assign new_n2244_ = new_n2243_;
  assign new_n2245_ = new_n2244_;
  assign new_n2246_ = new_n2243_;
  assign new_n2247_ = new_n1358_;
  assign new_n2248_ = new_n1318_;
  assign new_n2249_ = new_n2248_;
  assign new_n2250_ = new_n2248_;
  assign new_n2251_ = new_n1568_;
  assign new_n2252_ = new_n994_;
  assign new_n2253_ = new_n2252_;
  assign new_n2254_ = new_n2252_;
  assign new_n2255_ = new_n1569_;
  assign new_n2256_ = new_n2255_;
  assign new_n2257_ = new_n993_;
  assign new_n2258_ = new_n2257_;
  assign new_n2259_ = new_n2258_;
  assign new_n2260_ = new_n2257_;
  assign new_n2261_ = new_n1261_;
  assign new_n2262_ = new_n2261_;
  assign new_n2263_ = new_n1262_;
  assign new_n2264_ = new_n2263_;
  assign new_n2265_ = new_n1263_;
  assign new_n2266_ = new_n2265_;
  assign new_n2267_ = new_n1264_;
  assign new_n2268_ = new_n2267_;
  assign new_n2269_ = new_n1331_;
  assign new_n2270_ = new_n1332_;
  assign new_n2271_ = new_n1581_;
  assign new_n2272_ = new_n2271_;
  assign new_n2273_ = new_n1559_;
  assign new_n2274_ = new_n1580_;
  assign new_n2275_ = new_n2274_;
  assign new_n2276_ = new_n1558_;
  assign new_n2277_ = new_n2276_;
  assign new_n2278_ = new_n1585_;
  assign new_n2279_ = new_n2278_;
  assign new_n2280_ = new_n2278_;
  assign new_n2281_ = new_n1561_;
  assign new_n2282_ = new_n2281_;
  assign new_n2283_ = new_n1584_;
  assign new_n2284_ = new_n2283_;
  assign new_n2285_ = new_n2283_;
  assign new_n2286_ = new_n1560_;
  assign new_n2287_ = new_n2286_;
  assign new_n2288_ = new_n2286_;
  assign new_n2289_ = new_n1589_;
  assign new_n2290_ = new_n2289_;
  assign new_n2291_ = new_n2289_;
  assign new_n2292_ = new_n1563_;
  assign new_n2293_ = new_n2292_;
  assign new_n2294_ = new_n2292_;
  assign new_n2295_ = new_n1588_;
  assign new_n2296_ = new_n2295_;
  assign new_n2297_ = new_n2295_;
  assign new_n2298_ = new_n1562_;
  assign new_n2299_ = new_n2298_;
  assign new_n2300_ = new_n2299_;
  assign new_n2301_ = new_n2298_;
  assign new_n2302_ = new_n1571_;
  assign new_n2303_ = new_n1592_;
  assign new_n2304_ = new_n1598_;
  assign new_n2305_ = new_n1599_;
  assign new_n2306_ = new_n1351_;
  assign new_n2307_ = new_n1352_;
  assign new_n2308_ = new_n1349_;
  assign new_n2309_ = new_n1605_;
  assign new_n2310_ = new_n2309_;
  assign new_n2311_ = new_n2309_;
  assign new_n2312_ = new_n1604_;
  assign new_n2313_ = new_n2312_;
  assign new_n2314_ = new_n2312_;
  assign new_n2315_ = new_n1379_;
  assign new_n2316_ = new_n1616_;
  assign new_n2317_ = new_n2316_;
  assign new_n2318_ = new_n2316_;
  assign new_n2319_ = new_n1618_;
  assign new_n2320_ = new_n2319_;
  assign new_n2321_ = new_n1024_;
  assign new_n2322_ = new_n1620_;
  assign new_n2323_ = new_n2322_;
  assign new_n2324_ = new_n1030_;
  assign new_n2325_ = new_n1622_;
  assign new_n2326_ = new_n2325_;
  assign new_n2327_ = new_n1036_;
  assign new_n2328_ = new_n1395_;
  assign new_n2329_ = new_n1393_;
  assign new_n2330_ = new_n2329_;
  assign new_n2331_ = new_n1394_;
  assign new_n2332_ = new_n1397_;
  assign new_n2333_ = new_n2332_;
  assign new_n2334_ = new_n1364_;
  assign new_n2335_ = new_n1348_;
  assign new_n2336_ = new_n2335_;
  assign new_n2337_ = new_n2335_;
  assign new_n2338_ = new_n1390_;
  assign new_n2339_ = new_n1576_;
  assign new_n2340_ = new_n1257_;
  assign new_n2341_ = new_n2340_;
  assign new_n2342_ = new_n1258_;
  assign new_n2343_ = new_n2342_;
  assign new_n2344_ = new_n1578_;
  assign new_n2345_ = new_n1590_;
  assign new_n2346_ = new_n1277_;
  assign new_n2347_ = new_n2346_;
  assign new_n2348_ = new_n1231_;
  assign new_n2349_ = new_n2348_;
  assign new_n2350_ = new_n1278_;
  assign new_n2351_ = new_n1232_;
  assign new_n2352_ = new_n1235_;
  assign new_n2353_ = new_n2352_;
  assign new_n2354_ = new_n1233_;
  assign new_n2355_ = new_n2354_;
  assign new_n2356_ = new_n1236_;
  assign new_n2357_ = new_n1234_;
  assign new_n2358_ = new_n1193_;
  assign new_n2359_ = new_n2358_;
  assign new_n2360_ = new_n1183_;
  assign new_n2361_ = new_n2360_;
  assign new_n2362_ = new_n1194_;
  assign new_n2363_ = new_n1184_;
  assign new_n2364_ = new_n1187_;
  assign new_n2365_ = new_n1185_;
  assign new_n2366_ = new_n2365_;
  assign new_n2367_ = new_n1188_;
  assign new_n2368_ = new_n1186_;
  assign new_n2369_ = new_n1255_;
  assign new_n2370_ = new_n2369_;
  assign new_n2371_ = new_n1213_;
  assign new_n2372_ = new_n2371_;
  assign new_n2373_ = new_n1256_;
  assign new_n2374_ = new_n1214_;
  assign new_n2375_ = new_n1217_;
  assign new_n2376_ = new_n2375_;
  assign new_n2377_ = new_n1215_;
  assign new_n2378_ = new_n2377_;
  assign new_n2379_ = new_n1218_;
  assign new_n2380_ = new_n1216_;
  assign new_n2381_ = new_n1557_;
  assign new_n2382_ = new_n1271_;
  assign new_n2383_ = new_n2382_;
  assign new_n2384_ = new_n1272_;
  assign new_n2385_ = new_n1269_;
  assign new_n2386_ = new_n1572_;
  assign new_n2387_ = new_n1574_;
  assign new_n2388_ = new_n1582_;
  assign new_n2389_ = new_n1586_;
  assign new_n2390_ = new_n1615_;
  assign new_n2391_ = new_n1594_;
  assign new_n2392_ = new_n1636_;
  assign new_n2393_ = new_n2392_;
  assign new_n2394_ = new_n1018_;
  assign new_n2395_ = new_n1243_;
  assign new_n2396_ = new_n1276_;
  assign new_n2397_ = new_n1246_;
  assign new_n2398_ = new_n921_;
  assign new_n2399_ = new_n1762_;
  assign new_n2400_ = new_n2399_;
  assign new_n2401_ = new_n2399_;
  assign new_n2402_ = new_n1637_;
  assign new_n2403_ = new_n1628_;
  assign new_n2404_ = new_n2403_;
  assign new_n2405_ = new_n2403_;
  assign new_n2406_ = new_n1385_;
  assign new_n2407_ = new_n2406_;
  assign new_n2408_ = new_n2406_;
  assign new_n2409_ = new_n1392_;
  assign new_n2410_ = new_n1387_;
  assign new_n2411_ = new_n1388_;
  assign new_n2412_ = new_n1389_;
  assign new_n2413_ = new_n1383_;
  assign new_n2414_ = new_n1630_;
  assign new_n2415_ = new_n2414_;
  assign new_n2416_ = new_n1624_;
  assign new_n2417_ = new_n2416_;
  assign new_n2418_ = new_n1631_;
  assign new_n2419_ = new_n1784_;
  assign new_n2420_ = new_n1625_;
  assign new_n2421_ = new_n2420_;
  assign new_n2422_ = new_n1632_;
  assign new_n2423_ = new_n1623_;
  assign new_n2424_ = new_n2423_;
  assign new_n2425_ = new_n976_;
  assign new_n2426_ = new_n2425_;
  assign new_n2427_ = new_n1759_;
  assign new_n2428_ = new_n2427_;
  assign new_n2429_ = new_n2427_;
  assign new_n2430_ = new_n1768_;
  assign new_n2431_ = new_n1766_;
  assign new_n2432_ = new_n2431_;
  assign new_n2433_ = new_n2431_;
  assign new_n2434_ = new_n979_;
  assign new_n2435_ = new_n981_;
  assign new_n2436_ = new_n987_;
  assign new_n2437_ = new_n1782_;
  assign new_n2438_ = new_n2437_;
  assign new_n2439_ = new_n2437_;
  assign new_n2440_ = new_n947_;
  assign new_n2441_ = new_n951_;
  assign new_n2442_ = new_n955_;
  assign new_n2443_ = new_n1755_;
  assign new_n2444_ = new_n1123_;
  always @ (posedge clock) begin
    n480_lo <= n480_li;
    n492_lo <= n492_li;
    n495_lo <= n495_li;
    n498_lo <= n498_li;
    n501_lo <= n501_li;
    n504_lo <= n504_li;
    n516_lo <= n516_li;
    n528_lo <= n528_li;
    n531_lo <= n531_li;
    n540_lo <= n540_li;
    n543_lo <= n543_li;
    n546_lo <= n546_li;
    n549_lo <= n549_li;
    n552_lo <= n552_li;
    n564_lo <= n564_li;
    n579_lo <= n579_li;
    n600_lo <= n600_li;
    n603_lo <= n603_li;
    n606_lo <= n606_li;
    n609_lo <= n609_li;
    n612_lo <= n612_li;
    n615_lo <= n615_li;
    n618_lo <= n618_li;
    n621_lo <= n621_li;
    n627_lo <= n627_li;
    n630_lo <= n630_li;
    n633_lo <= n633_li;
    n639_lo <= n639_li;
    n642_lo <= n642_li;
    n645_lo <= n645_li;
    n648_lo <= n648_li;
    n660_lo <= n660_li;
    n663_lo <= n663_li;
    n672_lo <= n672_li;
    n675_lo <= n675_li;
    n678_lo <= n678_li;
    n681_lo <= n681_li;
    n684_lo <= n684_li;
    n687_lo <= n687_li;
    n690_lo <= n690_li;
    n693_lo <= n693_li;
    n696_lo <= n696_li;
    n699_lo <= n699_li;
    n702_lo <= n702_li;
    n705_lo <= n705_li;
    n708_lo <= n708_li;
    n711_lo <= n711_li;
    n714_lo <= n714_li;
    n717_lo <= n717_li;
    n720_lo <= n720_li;
    n723_lo <= n723_li;
    n726_lo <= n726_li;
    n729_lo <= n729_li;
    n732_lo <= n732_li;
    n735_lo <= n735_li;
    n738_lo <= n738_li;
    n741_lo <= n741_li;
    n744_lo <= n744_li;
    n747_lo <= n747_li;
    n750_lo <= n750_li;
    n756_lo <= n756_li;
    n759_lo <= n759_li;
    n762_lo <= n762_li;
    n768_lo <= n768_li;
    n771_lo <= n771_li;
    n774_lo <= n774_li;
    n780_lo <= n780_li;
    n783_lo <= n783_li;
    n786_lo <= n786_li;
    n792_lo <= n792_li;
    n795_lo <= n795_li;
    n804_lo <= n804_li;
    n807_lo <= n807_li;
    n816_lo <= n816_li;
    n819_lo <= n819_li;
    n828_lo <= n828_li;
    n831_lo <= n831_li;
    n843_lo <= n843_li;
    n846_lo <= n846_li;
    n849_lo <= n849_li;
    n852_lo <= n852_li;
    n855_lo <= n855_li;
    n858_lo <= n858_li;
    n861_lo <= n861_li;
    n864_lo <= n864_li;
    n867_lo <= n867_li;
    n870_lo <= n870_li;
    n879_lo <= n879_li;
    n891_lo <= n891_li;
    n903_lo <= n903_li;
    n915_lo <= n915_li;
    n918_lo <= n918_li;
    n927_lo <= n927_li;
    n951_lo <= n951_li;
    n954_lo <= n954_li;
    n957_lo <= n957_li;
    n960_lo <= n960_li;
    n963_lo <= n963_li;
    n966_lo <= n966_li;
    n972_lo <= n972_li;
    n975_lo <= n975_li;
    n978_lo <= n978_li;
    n984_lo <= n984_li;
    n987_lo <= n987_li;
    n990_lo <= n990_li;
    n996_lo <= n996_li;
    n999_lo <= n999_li;
    n1002_lo <= n1002_li;
    n1008_lo <= n1008_li;
    n1011_lo <= n1011_li;
    n1014_lo <= n1014_li;
    n1020_lo <= n1020_li;
    n1023_lo <= n1023_li;
    n1026_lo <= n1026_li;
    n1032_lo <= n1032_li;
    n1035_lo <= n1035_li;
    n1038_lo <= n1038_li;
    n1044_lo <= n1044_li;
    n1047_lo <= n1047_li;
    n1050_lo <= n1050_li;
    n1053_lo <= n1053_li;
    n1056_lo <= n1056_li;
    n1059_lo <= n1059_li;
    n1062_lo <= n1062_li;
    n1065_lo <= n1065_li;
    n1068_lo <= n1068_li;
    n1071_lo <= n1071_li;
    n1074_lo <= n1074_li;
    n1077_lo <= n1077_li;
    n1080_lo <= n1080_li;
    n1083_lo <= n1083_li;
    n1086_lo <= n1086_li;
    n1089_lo <= n1089_li;
    n1092_lo <= n1092_li;
    n1095_lo <= n1095_li;
    n1098_lo <= n1098_li;
    n1101_lo <= n1101_li;
    n1104_lo <= n1104_li;
    n1107_lo <= n1107_li;
    n1110_lo <= n1110_li;
    n1113_lo <= n1113_li;
    n1116_lo <= n1116_li;
    n1119_lo <= n1119_li;
    n1122_lo <= n1122_li;
    n1125_lo <= n1125_li;
    n1128_lo <= n1128_li;
    n1131_lo <= n1131_li;
    n1134_lo <= n1134_li;
    n1137_lo <= n1137_li;
    n1140_lo <= n1140_li;
    n1143_lo <= n1143_li;
    n1146_lo <= n1146_li;
    n1149_lo <= n1149_li;
    n1152_lo <= n1152_li;
    n1155_lo <= n1155_li;
    n1158_lo <= n1158_li;
    n1167_lo <= n1167_li;
    n1170_lo <= n1170_li;
    n1173_lo <= n1173_li;
    n1176_lo <= n1176_li;
    n1179_lo <= n1179_li;
    n1529_o2 <= n1529_i2;
    n1616_o2 <= n1616_i2;
    n1655_o2 <= n1655_i2;
    n1656_o2 <= n1656_i2;
    n1657_o2 <= n1657_i2;
    n1730_o2 <= n1730_i2;
    n1731_o2 <= n1731_i2;
    n1732_o2 <= n1732_i2;
    n1729_o2 <= n1729_i2;
    n1805_o2 <= n1805_i2;
    n1808_o2 <= n1808_i2;
    n1807_o2 <= n1807_i2;
    n1809_o2 <= n1809_i2;
    n1663_o2 <= n1663_i2;
    n1664_o2 <= n1664_i2;
    n1704_o2 <= n1704_i2;
    n1705_o2 <= n1705_i2;
    n1706_o2 <= n1706_i2;
    n1707_o2 <= n1707_i2;
    n1708_o2 <= n1708_i2;
    n1709_o2 <= n1709_i2;
    G280_o2 <= G280_i2;
    G655_o2 <= G655_i2;
    G663_o2 <= G663_i2;
    G672_o2 <= G672_i2;
    G538_o2 <= G538_i2;
    n1780_o2 <= n1780_i2;
    n1781_o2 <= n1781_i2;
    n1797_o2 <= n1797_i2;
    n1798_o2 <= n1798_i2;
    n1799_o2 <= n1799_i2;
    n1800_o2 <= n1800_i2;
    G578_o2 <= G578_i2;
    n1828_o2 <= n1828_i2;
    n801_lo_buf_o2 <= n801_lo_buf_i2;
    G693_o2 <= G693_i2;
    G702_o2 <= G702_i2;
    G712_o2 <= G712_i2;
    G685_o2 <= G685_i2;
    G658_o2 <= G658_i2;
    G667_o2 <= G667_i2;
    G677_o2 <= G677_i2;
    G650_o2 <= G650_i2;
    G798_o2 <= G798_i2;
    n1017_lo_buf_o2 <= n1017_lo_buf_i2;
    n1029_lo_buf_o2 <= n1029_lo_buf_i2;
    n1041_lo_buf_o2 <= n1041_lo_buf_i2;
    G558_o2 <= G558_i2;
    G562_o2 <= G562_i2;
    G566_o2 <= G566_i2;
    n1835_o2 <= n1835_i2;
    n1836_o2 <= n1836_i2;
    n1837_o2 <= n1837_i2;
    n765_lo_buf_o2 <= n765_lo_buf_i2;
    n777_lo_buf_o2 <= n777_lo_buf_i2;
    n789_lo_buf_o2 <= n789_lo_buf_i2;
    G617_o2 <= G617_i2;
    G626_o2 <= G626_i2;
    G636_o2 <= G636_i2;
    n489_lo_buf_o2 <= n489_lo_buf_i2;
    n513_lo_buf_o2 <= n513_lo_buf_i2;
    n561_lo_buf_o2 <= n561_lo_buf_i2;
    n597_lo_buf_o2 <= n597_lo_buf_i2;
    n657_lo_buf_o2 <= n657_lo_buf_i2;
    G276_o2 <= G276_i2;
    n1005_lo_buf_o2 <= n1005_lo_buf_i2;
    n1161_lo_buf_o2 <= n1161_lo_buf_i2;
    G620_o2 <= G620_i2;
    G629_o2 <= G629_i2;
    G639_o2 <= G639_i2;
    G554_o2 <= G554_i2;
    G690_o2 <= G690_i2;
    G698_o2 <= G698_i2;
    G707_o2 <= G707_i2;
    G319_o2 <= G319_i2;
    G389_o2 <= G389_i2;
    n753_lo_buf_o2 <= n753_lo_buf_i2;
    G647_o2 <= G647_i2;
    G769_o2 <= G769_i2;
    G785_o2 <= G785_i2;
    G808_o2 <= G808_i2;
    G445_o2 <= G445_i2;
    G448_o2 <= G448_i2;
    G477_o2 <= G477_i2;
    G480_o2 <= G480_i2;
    G436_o2 <= G436_i2;
    G786_o2 <= G786_i2;
    G787_o2 <= G787_i2;
    G826_o2 <= G826_i2;
    G827_o2 <= G827_i2;
    G825_o2 <= G825_i2;
    G610_o2 <= G610_i2;
    n537_lo_buf_o2 <= n537_lo_buf_i2;
    n669_lo_buf_o2 <= n669_lo_buf_i2;
    n969_lo_buf_o2 <= n969_lo_buf_i2;
    n981_lo_buf_o2 <= n981_lo_buf_i2;
    n993_lo_buf_o2 <= n993_lo_buf_i2;
    G309_o2 <= G309_i2;
    G461_o2 <= G461_i2;
    G487_o2 <= G487_i2;
    G460_o2 <= G460_i2;
    G468_o2 <= G468_i2;
    G287_o2 <= G287_i2;
    G613_o2 <= G613_i2;
    n585_lo_buf_o2 <= n585_lo_buf_i2;
    n813_lo_buf_o2 <= n813_lo_buf_i2;
    n825_lo_buf_o2 <= n825_lo_buf_i2;
    n837_lo_buf_o2 <= n837_lo_buf_i2;
    n897_lo_buf_o2 <= n897_lo_buf_i2;
    n909_lo_buf_o2 <= n909_lo_buf_i2;
    n933_lo_buf_o2 <= n933_lo_buf_i2;
    G451_o2 <= G451_i2;
    G682_o2 <= G682_i2;
    G756_o2 <= G756_i2;
    G542_o2 <= G542_i2;
    G546_o2 <= G546_i2;
    G550_o2 <= G550_i2;
    G310_o2 <= G310_i2;
    n798_lo_buf_o2 <= n798_lo_buf_i2;
    n882_lo_buf_o2 <= n882_lo_buf_i2;
    G427_o2 <= G427_i2;
    G497_o2 <= G497_i2;
    G499_o2 <= G499_i2;
    G501_o2 <= G501_i2;
    G498_o2 <= G498_i2;
    G500_o2 <= G500_i2;
    G502_o2 <= G502_i2;
    G369_o2 <= G369_i2;
    n939_lo_buf_o2 <= n939_lo_buf_i2;
    n486_lo_buf_o2 <= n486_lo_buf_i2;
    n510_lo_buf_o2 <= n510_lo_buf_i2;
    n558_lo_buf_o2 <= n558_lo_buf_i2;
    n594_lo_buf_o2 <= n594_lo_buf_i2;
    n654_lo_buf_o2 <= n654_lo_buf_i2;
    n477_lo_buf_o2 <= n477_lo_buf_i2;
    n525_lo_buf_o2 <= n525_lo_buf_i2;
    n573_lo_buf_o2 <= n573_lo_buf_i2;
  end
  initial begin
    n480_lo <= 1'b0;
    n492_lo <= 1'b0;
    n495_lo <= 1'b0;
    n498_lo <= 1'b0;
    n501_lo <= 1'b0;
    n504_lo <= 1'b0;
    n516_lo <= 1'b0;
    n528_lo <= 1'b0;
    n531_lo <= 1'b0;
    n540_lo <= 1'b0;
    n543_lo <= 1'b0;
    n546_lo <= 1'b0;
    n549_lo <= 1'b0;
    n552_lo <= 1'b0;
    n564_lo <= 1'b0;
    n579_lo <= 1'b0;
    n600_lo <= 1'b0;
    n603_lo <= 1'b0;
    n606_lo <= 1'b0;
    n609_lo <= 1'b0;
    n612_lo <= 1'b0;
    n615_lo <= 1'b0;
    n618_lo <= 1'b0;
    n621_lo <= 1'b0;
    n627_lo <= 1'b0;
    n630_lo <= 1'b0;
    n633_lo <= 1'b0;
    n639_lo <= 1'b0;
    n642_lo <= 1'b0;
    n645_lo <= 1'b0;
    n648_lo <= 1'b0;
    n660_lo <= 1'b0;
    n663_lo <= 1'b0;
    n672_lo <= 1'b0;
    n675_lo <= 1'b0;
    n678_lo <= 1'b0;
    n681_lo <= 1'b0;
    n684_lo <= 1'b0;
    n687_lo <= 1'b0;
    n690_lo <= 1'b0;
    n693_lo <= 1'b0;
    n696_lo <= 1'b0;
    n699_lo <= 1'b0;
    n702_lo <= 1'b0;
    n705_lo <= 1'b0;
    n708_lo <= 1'b0;
    n711_lo <= 1'b0;
    n714_lo <= 1'b0;
    n717_lo <= 1'b0;
    n720_lo <= 1'b0;
    n723_lo <= 1'b0;
    n726_lo <= 1'b0;
    n729_lo <= 1'b0;
    n732_lo <= 1'b0;
    n735_lo <= 1'b0;
    n738_lo <= 1'b0;
    n741_lo <= 1'b0;
    n744_lo <= 1'b0;
    n747_lo <= 1'b0;
    n750_lo <= 1'b0;
    n756_lo <= 1'b0;
    n759_lo <= 1'b0;
    n762_lo <= 1'b0;
    n768_lo <= 1'b0;
    n771_lo <= 1'b0;
    n774_lo <= 1'b0;
    n780_lo <= 1'b0;
    n783_lo <= 1'b0;
    n786_lo <= 1'b0;
    n792_lo <= 1'b0;
    n795_lo <= 1'b0;
    n804_lo <= 1'b0;
    n807_lo <= 1'b0;
    n816_lo <= 1'b0;
    n819_lo <= 1'b0;
    n828_lo <= 1'b0;
    n831_lo <= 1'b0;
    n843_lo <= 1'b0;
    n846_lo <= 1'b0;
    n849_lo <= 1'b0;
    n852_lo <= 1'b0;
    n855_lo <= 1'b0;
    n858_lo <= 1'b0;
    n861_lo <= 1'b0;
    n864_lo <= 1'b0;
    n867_lo <= 1'b0;
    n870_lo <= 1'b0;
    n879_lo <= 1'b0;
    n891_lo <= 1'b0;
    n903_lo <= 1'b0;
    n915_lo <= 1'b0;
    n918_lo <= 1'b0;
    n927_lo <= 1'b0;
    n951_lo <= 1'b0;
    n954_lo <= 1'b0;
    n957_lo <= 1'b0;
    n960_lo <= 1'b0;
    n963_lo <= 1'b0;
    n966_lo <= 1'b0;
    n972_lo <= 1'b0;
    n975_lo <= 1'b0;
    n978_lo <= 1'b0;
    n984_lo <= 1'b0;
    n987_lo <= 1'b0;
    n990_lo <= 1'b0;
    n996_lo <= 1'b0;
    n999_lo <= 1'b0;
    n1002_lo <= 1'b0;
    n1008_lo <= 1'b0;
    n1011_lo <= 1'b0;
    n1014_lo <= 1'b0;
    n1020_lo <= 1'b0;
    n1023_lo <= 1'b0;
    n1026_lo <= 1'b0;
    n1032_lo <= 1'b0;
    n1035_lo <= 1'b0;
    n1038_lo <= 1'b0;
    n1044_lo <= 1'b0;
    n1047_lo <= 1'b0;
    n1050_lo <= 1'b0;
    n1053_lo <= 1'b0;
    n1056_lo <= 1'b0;
    n1059_lo <= 1'b0;
    n1062_lo <= 1'b0;
    n1065_lo <= 1'b0;
    n1068_lo <= 1'b0;
    n1071_lo <= 1'b0;
    n1074_lo <= 1'b0;
    n1077_lo <= 1'b0;
    n1080_lo <= 1'b0;
    n1083_lo <= 1'b0;
    n1086_lo <= 1'b0;
    n1089_lo <= 1'b0;
    n1092_lo <= 1'b0;
    n1095_lo <= 1'b0;
    n1098_lo <= 1'b0;
    n1101_lo <= 1'b0;
    n1104_lo <= 1'b0;
    n1107_lo <= 1'b0;
    n1110_lo <= 1'b0;
    n1113_lo <= 1'b0;
    n1116_lo <= 1'b0;
    n1119_lo <= 1'b0;
    n1122_lo <= 1'b0;
    n1125_lo <= 1'b0;
    n1128_lo <= 1'b0;
    n1131_lo <= 1'b0;
    n1134_lo <= 1'b0;
    n1137_lo <= 1'b0;
    n1140_lo <= 1'b0;
    n1143_lo <= 1'b0;
    n1146_lo <= 1'b0;
    n1149_lo <= 1'b0;
    n1152_lo <= 1'b0;
    n1155_lo <= 1'b0;
    n1158_lo <= 1'b0;
    n1167_lo <= 1'b0;
    n1170_lo <= 1'b0;
    n1173_lo <= 1'b0;
    n1176_lo <= 1'b0;
    n1179_lo <= 1'b0;
    n1529_o2 <= 1'b0;
    n1616_o2 <= 1'b0;
    n1655_o2 <= 1'b0;
    n1656_o2 <= 1'b0;
    n1657_o2 <= 1'b0;
    n1730_o2 <= 1'b0;
    n1731_o2 <= 1'b0;
    n1732_o2 <= 1'b0;
    n1729_o2 <= 1'b0;
    n1805_o2 <= 1'b0;
    n1808_o2 <= 1'b0;
    n1807_o2 <= 1'b0;
    n1809_o2 <= 1'b0;
    n1663_o2 <= 1'b0;
    n1664_o2 <= 1'b0;
    n1704_o2 <= 1'b0;
    n1705_o2 <= 1'b0;
    n1706_o2 <= 1'b0;
    n1707_o2 <= 1'b0;
    n1708_o2 <= 1'b0;
    n1709_o2 <= 1'b0;
    G280_o2 <= 1'b0;
    G655_o2 <= 1'b0;
    G663_o2 <= 1'b0;
    G672_o2 <= 1'b0;
    G538_o2 <= 1'b0;
    n1780_o2 <= 1'b0;
    n1781_o2 <= 1'b0;
    n1797_o2 <= 1'b0;
    n1798_o2 <= 1'b0;
    n1799_o2 <= 1'b0;
    n1800_o2 <= 1'b0;
    G578_o2 <= 1'b0;
    n1828_o2 <= 1'b0;
    n801_lo_buf_o2 <= 1'b0;
    G693_o2 <= 1'b0;
    G702_o2 <= 1'b0;
    G712_o2 <= 1'b0;
    G685_o2 <= 1'b0;
    G658_o2 <= 1'b0;
    G667_o2 <= 1'b0;
    G677_o2 <= 1'b0;
    G650_o2 <= 1'b0;
    G798_o2 <= 1'b0;
    n1017_lo_buf_o2 <= 1'b0;
    n1029_lo_buf_o2 <= 1'b0;
    n1041_lo_buf_o2 <= 1'b0;
    G558_o2 <= 1'b0;
    G562_o2 <= 1'b0;
    G566_o2 <= 1'b0;
    n1835_o2 <= 1'b0;
    n1836_o2 <= 1'b0;
    n1837_o2 <= 1'b0;
    n765_lo_buf_o2 <= 1'b0;
    n777_lo_buf_o2 <= 1'b0;
    n789_lo_buf_o2 <= 1'b0;
    G617_o2 <= 1'b0;
    G626_o2 <= 1'b0;
    G636_o2 <= 1'b0;
    n489_lo_buf_o2 <= 1'b0;
    n513_lo_buf_o2 <= 1'b0;
    n561_lo_buf_o2 <= 1'b0;
    n597_lo_buf_o2 <= 1'b0;
    n657_lo_buf_o2 <= 1'b0;
    G276_o2 <= 1'b0;
    n1005_lo_buf_o2 <= 1'b0;
    n1161_lo_buf_o2 <= 1'b0;
    G620_o2 <= 1'b0;
    G629_o2 <= 1'b0;
    G639_o2 <= 1'b0;
    G554_o2 <= 1'b0;
    G690_o2 <= 1'b0;
    G698_o2 <= 1'b0;
    G707_o2 <= 1'b0;
    G319_o2 <= 1'b0;
    G389_o2 <= 1'b0;
    n753_lo_buf_o2 <= 1'b0;
    G647_o2 <= 1'b0;
    G769_o2 <= 1'b0;
    G785_o2 <= 1'b0;
    G808_o2 <= 1'b0;
    G445_o2 <= 1'b0;
    G448_o2 <= 1'b0;
    G477_o2 <= 1'b0;
    G480_o2 <= 1'b0;
    G436_o2 <= 1'b0;
    G786_o2 <= 1'b0;
    G787_o2 <= 1'b0;
    G826_o2 <= 1'b0;
    G827_o2 <= 1'b0;
    G825_o2 <= 1'b0;
    G610_o2 <= 1'b0;
    n537_lo_buf_o2 <= 1'b0;
    n669_lo_buf_o2 <= 1'b0;
    n969_lo_buf_o2 <= 1'b0;
    n981_lo_buf_o2 <= 1'b0;
    n993_lo_buf_o2 <= 1'b0;
    G309_o2 <= 1'b0;
    G461_o2 <= 1'b0;
    G487_o2 <= 1'b0;
    G460_o2 <= 1'b0;
    G468_o2 <= 1'b0;
    G287_o2 <= 1'b0;
    G613_o2 <= 1'b0;
    n585_lo_buf_o2 <= 1'b0;
    n813_lo_buf_o2 <= 1'b0;
    n825_lo_buf_o2 <= 1'b0;
    n837_lo_buf_o2 <= 1'b0;
    n897_lo_buf_o2 <= 1'b0;
    n909_lo_buf_o2 <= 1'b0;
    n933_lo_buf_o2 <= 1'b0;
    G451_o2 <= 1'b0;
    G682_o2 <= 1'b0;
    G756_o2 <= 1'b0;
    G542_o2 <= 1'b0;
    G546_o2 <= 1'b0;
    G550_o2 <= 1'b0;
    G310_o2 <= 1'b0;
    n798_lo_buf_o2 <= 1'b0;
    n882_lo_buf_o2 <= 1'b0;
    G427_o2 <= 1'b0;
    G497_o2 <= 1'b0;
    G499_o2 <= 1'b0;
    G501_o2 <= 1'b0;
    G498_o2 <= 1'b0;
    G500_o2 <= 1'b0;
    G502_o2 <= 1'b0;
    G369_o2 <= 1'b0;
    n939_lo_buf_o2 <= 1'b0;
    n486_lo_buf_o2 <= 1'b0;
    n510_lo_buf_o2 <= 1'b0;
    n558_lo_buf_o2 <= 1'b0;
    n594_lo_buf_o2 <= 1'b0;
    n654_lo_buf_o2 <= 1'b0;
    n477_lo_buf_o2 <= 1'b0;
    n525_lo_buf_o2 <= 1'b0;
    n573_lo_buf_o2 <= 1'b0;
  end
endmodule


