// Benchmark "mymod" written by ABC on Wed Nov  1 23:37:48 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33,
    G1884, G1885, G1886, G1887, G1888, G1889, G1890, G1891, G1892, G1893,
    G1894, G1895, G1896, G1897, G1898, G1899, G1900, G1901, G1902, G1903,
    G1904, G1905, G1906, G1907, G1908  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33;
  output G1884, G1885, G1886, G1887, G1888, G1889, G1890, G1891, G1892, G1893,
    G1894, G1895, G1896, G1897, G1898, G1899, G1900, G1901, G1902, G1903,
    G1904, G1905, G1906, G1907, G1908;
  reg n940_lo, n949_lo, n961_lo, n973_lo, n976_lo, n985_lo, n988_lo,
    n997_lo, n1009_lo, n1021_lo, n1033_lo, n1045_lo, n1057_lo, n1060_lo,
    n1069_lo, n1081_lo, n1093_lo, n1105_lo, n1117_lo, n1120_lo, n1129_lo,
    n1132_lo, n1156_lo, n1168_lo, n1180_lo, n1189_lo, n1192_lo, n1195_lo,
    n1201_lo, n1204_lo, n1228_lo, n1231_lo, n1234_lo, n1237_lo, n1240_lo,
    n1243_lo, n1249_lo, n1252_lo, n1255_lo, n1261_lo, n1264_lo, n1267_lo,
    n1273_lo, n1276_lo, n1279_lo, n1282_lo, n1285_lo, n1288_lo, n1291_lo,
    n1294_lo, n1297_lo, n1300_lo, n1303_lo, n1309_lo, n1312_lo, n1315_lo,
    n1318_lo, n1321_lo, n1333_lo, n1225_o2, n1229_o2, n1228_o2, n1259_o2,
    n1272_o2, n1269_o2, n1307_o2, n1201_o2, n1202_o2, n1203_o2, n1204_o2,
    n622_o2, n1205_o2, n1206_o2, n497_o2, n1212_o2, n1213_o2, n1214_o2,
    n1215_o2, n1216_o2, n1217_o2, n1218_o2, n1219_o2, n1242_o2, n1243_o2,
    n1273_o2, n1274_o2, n1275_o2, n1276_o2, n1277_o2, n1286_o2, n1299_o2,
    n601_o2, n625_o2, n463_o2, lo082_buf_o2, n455_o2, n642_o2, n459_o2,
    n501_o2, n599_o2, n485_o2, lo086_buf_o2, lo122_buf_o2, n502_o2,
    n627_o2, lo038_buf_o2, lo046_buf_o2, lo050_buf_o2, lo058_buf_o2,
    lo070_buf_o2, lo094_buf_o2, n462_o2, lo006_buf_o2, lo010_buf_o2,
    lo022_buf_o2, lo026_buf_o2, lo030_buf_o2, lo034_buf_o2, lo054_buf_o2,
    lo130_buf_o2, n547_o2, n424_inv, n617_o2, lo042_buf_o2, lo062_buf_o2,
    lo110_buf_o2, n733_o2, n734_o2, n570_o2, n461_o2, n644_o2, n628_o2,
    n528_o2, n460_inv, lo002_buf_o2, lo014_buf_o2, lo018_buf_o2,
    lo078_buf_o2, lo090_buf_o2, n513_o2, lo102_buf_o2, lo106_buf_o2,
    n600_o2, n529_o2, n593_o2, lo066_buf_o2, n549_o2, n550_o2, n571_o2,
    n572_o2, n495_o2, n496_o2, n620_o2, n482_o2, lo081_buf_o2, n576_o2,
    n520_o2, n521_o2, n562_o2, n508_o2, n509_o2, lo074_buf_o2, n539_o2,
    n536_o2, n516_o2, n491_o2, n557_o2, n586_o2, n483_o2, n484_o2,
    lo004_buf_o2, lo008_buf_o2, lo020_buf_o2, lo024_buf_o2, lo028_buf_o2,
    lo032_buf_o2, lo052_buf_o2, lo128_buf_o2, lo037_buf_o2, lo045_buf_o2,
    lo049_buf_o2, lo057_buf_o2, lo069_buf_o2, lo093_buf_o2;
  wire new_new_n427__, new_new_n429__, new_new_n431__, new_new_n433__,
    new_new_n435__, new_new_n437__, new_new_n439__, new_new_n441__,
    new_new_n443__, new_new_n445__, new_new_n447__, new_new_n449__,
    new_new_n451__, new_new_n453__, new_new_n455__, new_new_n457__,
    new_new_n459__, new_new_n461__, new_new_n463__, new_new_n465__,
    new_new_n467__, new_new_n469__, new_new_n471__, new_new_n473__,
    new_new_n475__, new_new_n477__, new_new_n479__, new_new_n481__,
    new_new_n483__, new_new_n485__, new_new_n487__, new_new_n489__,
    new_new_n491__, new_new_n493__, new_new_n494__, new_new_n495__,
    new_new_n496__, new_new_n497__, new_new_n498__, new_new_n499__,
    new_new_n500__, new_new_n501__, new_new_n502__, new_new_n503__,
    new_new_n504__, new_new_n505__, new_new_n506__, new_new_n507__,
    new_new_n508__, new_new_n509__, new_new_n510__, new_new_n511__,
    new_new_n512__, new_new_n513__, new_new_n514__, new_new_n515__,
    new_new_n516__, new_new_n517__, new_new_n518__, new_new_n519__,
    new_new_n520__, new_new_n521__, new_new_n522__, new_new_n523__,
    new_new_n524__, new_new_n525__, new_new_n526__, new_new_n527__,
    new_new_n528__, new_new_n529__, new_new_n530__, new_new_n531__,
    new_new_n532__, new_new_n533__, new_new_n534__, new_new_n535__,
    new_new_n537__, new_new_n539__, new_new_n541__, new_new_n543__,
    new_new_n544__, new_new_n545__, new_new_n547__, new_new_n548__,
    new_new_n549__, new_new_n550__, new_new_n551__, new_new_n552__,
    new_new_n553__, new_new_n555__, new_new_n557__, new_new_n558__,
    new_new_n559__, new_new_n560__, new_new_n561__, new_new_n563__,
    new_new_n566__, new_new_n567__, new_new_n569__, new_new_n571__,
    new_new_n573__, new_new_n575__, new_new_n576__, new_new_n577__,
    new_new_n579__, new_new_n581__, new_new_n583__, new_new_n585__,
    new_new_n586__, new_new_n587__, new_new_n589__, new_new_n591__,
    new_new_n593__, new_new_n594__, new_new_n595__, new_new_n597__,
    new_new_n598__, new_new_n599__, new_new_n600__, new_new_n601__,
    new_new_n603__, new_new_n605__, new_new_n607__, new_new_n609__,
    new_new_n610__, new_new_n612__, new_new_n613__, new_new_n614__,
    new_new_n615__, new_new_n617__, new_new_n620__, new_new_n622__,
    new_new_n623__, new_new_n624__, new_new_n625__, new_new_n627__,
    new_new_n629__, new_new_n631__, new_new_n633__, new_new_n634__,
    new_new_n636__, new_new_n637__, new_new_n639__, new_new_n640__,
    new_new_n641__, new_new_n643__, new_new_n645__, new_new_n647__,
    new_new_n649__, new_new_n651__, new_new_n653__, new_new_n655__,
    new_new_n657__, new_new_n659__, new_new_n661__, new_new_n663__,
    new_new_n665__, new_new_n668__, new_new_n670__, new_new_n671__,
    new_new_n672__, new_new_n673__, new_new_n674__, new_new_n675__,
    new_new_n676__, new_new_n677__, new_new_n678__, new_new_n679__,
    new_new_n680__, new_new_n681__, new_new_n683__, new_new_n684__,
    new_new_n685__, new_new_n686__, new_new_n687__, new_new_n689__,
    new_new_n690__, new_new_n691__, new_new_n692__, new_new_n693__,
    new_new_n694__, new_new_n695__, new_new_n697__, new_new_n698__,
    new_new_n699__, new_new_n700__, new_new_n701__, new_new_n702__,
    new_new_n703__, new_new_n705__, new_new_n707__, new_new_n708__,
    new_new_n709__, new_new_n711__, new_new_n713__, new_new_n716__,
    new_new_n717__, new_new_n718__, new_new_n719__, new_new_n721__,
    new_new_n723__, new_new_n725__, new_new_n726__, new_new_n727__,
    new_new_n728__, new_new_n729__, new_new_n730__, new_new_n731__,
    new_new_n732__, new_new_n733__, new_new_n735__, new_new_n737__,
    new_new_n739__, new_new_n741__, new_new_n743__, new_new_n745__,
    new_new_n746__, new_new_n747__, new_new_n748__, new_new_n749__,
    new_new_n751__, new_new_n752__, new_new_n753__, new_new_n754__,
    new_new_n755__, new_new_n756__, new_new_n757__, new_new_n759__,
    new_new_n761__, new_new_n762__, new_new_n763__, new_new_n764__,
    new_new_n765__, new_new_n767__, new_new_n769__, new_new_n770__,
    new_new_n771__, new_new_n773__, new_new_n774__, new_new_n775__,
    new_new_n776__, new_new_n777__, new_new_n778__, new_new_n779__,
    new_new_n780__, new_new_n781__, new_new_n782__, new_new_n783__,
    new_new_n786__, new_new_n788__, new_new_n789__, new_new_n792__,
    new_new_n793__, new_new_n794__, new_new_n795__, new_new_n796__,
    new_new_n797__, new_new_n798__, new_new_n799__, new_new_n800__,
    new_new_n801__, new_new_n802__, new_new_n803__, new_new_n804__,
    new_new_n805__, new_new_n806__, new_new_n807__, new_new_n808__,
    new_new_n809__, new_new_n810__, new_new_n811__, new_new_n812__,
    new_new_n813__, new_new_n814__, new_new_n815__, new_new_n816__,
    new_new_n817__, new_new_n818__, new_new_n819__, new_new_n820__,
    new_new_n821__, new_new_n822__, new_new_n823__, new_new_n824__,
    new_new_n825__, new_new_n826__, new_new_n827__, new_new_n828__,
    new_new_n829__, new_new_n830__, new_new_n831__, new_new_n832__,
    new_new_n833__, new_new_n834__, new_new_n835__, new_new_n836__,
    new_new_n837__, new_new_n838__, new_new_n839__, new_new_n840__,
    new_new_n841__, new_new_n842__, new_new_n843__, new_new_n844__,
    new_new_n845__, new_new_n846__, new_new_n847__, new_new_n848__,
    new_new_n849__, new_new_n850__, new_new_n851__, new_new_n852__,
    new_new_n853__, new_new_n854__, new_new_n855__, new_new_n856__,
    new_new_n857__, new_new_n858__, new_new_n859__, new_new_n860__,
    new_new_n861__, new_new_n862__, new_new_n863__, new_new_n864__,
    new_new_n865__, new_new_n866__, new_new_n867__, new_new_n868__,
    new_new_n869__, new_new_n870__, new_new_n871__, new_new_n872__,
    new_new_n873__, new_new_n874__, new_new_n875__, new_new_n876__,
    new_new_n877__, new_new_n878__, new_new_n879__, new_new_n880__,
    new_new_n881__, new_new_n882__, new_new_n883__, new_new_n884__,
    new_new_n885__, new_new_n886__, new_new_n887__, new_new_n888__,
    new_new_n889__, new_new_n890__, new_new_n891__, new_new_n892__,
    new_new_n893__, new_new_n894__, new_new_n895__, new_new_n896__,
    new_new_n897__, new_new_n898__, new_new_n899__, new_new_n900__,
    new_new_n901__, new_new_n902__, new_new_n903__, new_new_n904__,
    new_new_n905__, new_new_n906__, new_new_n907__, new_new_n908__,
    new_new_n909__, new_new_n910__, new_new_n911__, new_new_n912__,
    new_new_n913__, new_new_n914__, new_new_n915__, new_new_n916__,
    new_new_n917__, new_new_n918__, new_new_n919__, new_new_n920__,
    new_new_n921__, new_new_n922__, new_new_n923__, new_new_n924__,
    new_new_n925__, new_new_n926__, new_new_n927__, new_new_n928__,
    new_new_n929__, new_new_n930__, new_new_n931__, new_new_n932__,
    new_new_n933__, new_new_n934__, new_new_n935__, new_new_n936__,
    new_new_n937__, new_new_n938__, new_new_n939__, new_new_n940__,
    new_new_n941__, new_new_n942__, new_new_n943__, new_new_n944__,
    new_new_n945__, new_new_n946__, new_new_n947__, new_new_n948__,
    new_new_n949__, new_new_n950__, new_new_n951__, new_new_n952__,
    new_new_n953__, new_new_n954__, new_new_n955__, new_new_n956__,
    new_new_n957__, new_new_n958__, new_new_n959__, new_new_n960__,
    new_new_n961__, new_new_n962__, new_new_n963__, new_new_n964__,
    new_new_n965__, new_new_n966__, new_new_n967__, new_new_n968__,
    new_new_n969__, new_new_n970__, new_new_n971__, new_new_n972__,
    new_new_n973__, new_new_n974__, new_new_n975__, new_new_n976__,
    new_new_n977__, new_new_n978__, new_new_n979__, new_new_n980__,
    new_new_n981__, new_new_n982__, new_new_n983__, new_new_n984__,
    new_new_n985__, new_new_n986__, new_new_n987__, new_new_n988__,
    new_new_n989__, new_new_n990__, new_new_n991__, new_new_n992__,
    new_new_n993__, new_new_n994__, new_new_n995__, new_new_n996__,
    new_new_n997__, new_new_n998__, new_new_n999__, new_new_n1000__,
    new_new_n1001__, new_new_n1002__, new_new_n1003__, new_new_n1004__,
    new_new_n1005__, new_new_n1006__, new_new_n1007__, new_new_n1008__,
    new_new_n1009__, new_new_n1010__, new_new_n1011__, new_new_n1012__,
    new_new_n1013__, new_new_n1014__, new_new_n1015__, new_new_n1016__,
    new_new_n1017__, new_new_n1018__, new_new_n1019__, new_new_n1020__,
    new_new_n1021__, new_new_n1022__, new_new_n1023__, new_new_n1024__,
    new_new_n1025__, new_new_n1026__, new_new_n1027__, new_new_n1028__,
    new_new_n1029__, new_new_n1030__, new_new_n1031__, new_new_n1032__,
    new_new_n1033__, new_new_n1034__, new_new_n1035__, new_new_n1036__,
    new_new_n1037__, new_new_n1038__, new_new_n1039__, new_new_n1040__,
    new_new_n1041__, new_new_n1042__, new_new_n1043__, new_new_n1044__,
    new_new_n1045__, new_new_n1046__, new_new_n1047__, new_new_n1048__,
    new_new_n1049__, new_new_n1050__, new_new_n1051__, new_new_n1052__,
    new_new_n1053__, new_new_n1054__, new_new_n1055__, new_new_n1056__,
    new_new_n1057__, new_new_n1058__, new_new_n1059__, new_new_n1060__,
    new_new_n1061__, new_new_n1062__, new_new_n1063__, new_new_n1064__,
    new_new_n1065__, new_new_n1066__, new_new_n1067__, new_new_n1068__,
    new_new_n1069__, new_new_n1070__, new_new_n1071__, new_new_n1072__,
    new_new_n1073__, new_new_n1074__, new_new_n1075__, new_new_n1076__,
    new_new_n1077__, new_new_n1078__, new_new_n1079__, new_new_n1080__,
    new_new_n1081__, new_new_n1082__, new_new_n1083__, new_new_n1084__,
    new_new_n1085__, new_new_n1086__, new_new_n1087__, new_new_n1088__,
    new_new_n1089__, new_new_n1090__, new_new_n1091__, new_new_n1092__,
    new_new_n1093__, new_new_n1094__, new_new_n1095__, new_new_n1096__,
    new_new_n1097__, new_new_n1098__, new_new_n1099__, new_new_n1100__,
    new_new_n1101__, new_new_n1102__, new_new_n1103__, new_new_n1104__,
    new_new_n1105__, new_new_n1106__, new_new_n1107__, new_new_n1108__,
    new_new_n1109__, new_new_n1110__, new_new_n1111__, new_new_n1112__,
    new_new_n1113__, new_new_n1114__, new_new_n1115__, new_new_n1116__,
    new_new_n1117__, new_new_n1118__, new_new_n1119__, new_new_n1120__,
    new_new_n1121__, new_new_n1122__, new_new_n1123__, new_new_n1124__,
    new_new_n1125__, new_new_n1126__, new_new_n1127__, new_new_n1128__,
    new_new_n1129__, new_new_n1130__, new_new_n1131__, new_new_n1132__,
    new_new_n1133__, new_new_n1134__, new_new_n1135__, new_new_n1136__,
    new_new_n1137__, new_new_n1138__, new_new_n1139__, new_new_n1140__,
    new_new_n1141__, new_new_n1142__, new_new_n1143__, new_new_n1144__,
    new_new_n1145__, new_new_n1146__, new_new_n1147__, new_new_n1148__,
    new_new_n1149__, new_new_n1150__, new_new_n1151__, new_new_n1152__,
    new_new_n1153__, new_new_n1154__, new_new_n1155__, new_new_n1156__,
    new_new_n1157__, new_new_n1158__, new_new_n1159__, new_new_n1160__,
    new_new_n1161__, new_new_n1162__, new_new_n1163__, new_new_n1164__,
    new_new_n1165__, new_new_n1166__, new_new_n1167__, new_new_n1168__,
    new_new_n1169__, new_new_n1170__, new_new_n1171__, new_new_n1172__,
    new_new_n1173__, new_new_n1174__, new_new_n1175__, new_new_n1176__,
    new_new_n1177__, new_new_n1178__, new_new_n1179__, new_new_n1180__,
    new_new_n1181__, new_new_n1182__, new_new_n1183__, new_new_n1184__,
    new_new_n1185__, new_new_n1186__, new_new_n1187__, new_new_n1188__,
    new_new_n1189__, new_new_n1190__, new_new_n1191__, new_new_n1192__,
    new_new_n1193__, new_new_n1194__, new_new_n1195__, new_new_n1196__,
    new_new_n1197__, new_new_n1198__, new_new_n1199__, new_new_n1200__,
    new_new_n1201__, new_new_n1202__, new_new_n1203__, new_new_n1204__,
    new_new_n1205__, new_new_n1206__, new_new_n1207__, new_new_n1208__,
    new_new_n1209__, new_new_n1210__, new_new_n1211__, new_new_n1212__,
    new_new_n1213__, new_new_n1214__, new_new_n1215__, new_new_n1216__,
    new_new_n1217__, new_new_n1218__, new_new_n1219__, new_new_n1220__,
    new_new_n1221__, new_new_n1222__, new_new_n1223__, new_new_n1224__,
    new_new_n1225__, new_new_n1226__, new_new_n1227__, new_new_n1228__,
    new_new_n1229__, new_new_n1230__, new_new_n1231__, new_new_n1232__,
    new_new_n1233__, new_new_n1234__, new_new_n1235__, new_new_n1236__,
    new_new_n1237__, new_new_n1238__, new_new_n1239__, new_new_n1240__,
    new_new_n1241__, new_new_n1242__, new_new_n1243__, new_new_n1244__,
    new_new_n1245__, new_new_n1246__, new_new_n1247__, new_new_n1248__,
    new_new_n1249__, new_new_n1250__, new_new_n1251__, new_new_n1252__,
    new_new_n1253__, new_new_n1254__, new_new_n1464__, new_new_n1465__,
    new_new_n1466__, new_new_n1467__, new_new_n1468__, new_new_n1469__,
    new_new_n1470__, new_new_n1471__, new_new_n1472__, new_new_n1473__,
    new_new_n1474__, new_new_n1475__, new_new_n1476__, new_new_n1477__,
    new_new_n1478__, new_new_n1479__, new_new_n1480__, new_new_n1481__,
    new_new_n1482__, new_new_n1483__, new_new_n1484__, new_new_n1485__,
    new_new_n1486__, new_new_n1487__, new_new_n1488__, new_new_n1489__,
    new_new_n1490__, new_new_n1491__, new_new_n1492__, new_new_n1493__,
    new_new_n1494__, new_new_n1495__, new_new_n1496__, new_new_n1497__,
    new_new_n1498__, new_new_n1499__, new_new_n1500__, new_new_n1501__,
    new_new_n1502__, new_new_n1503__, new_new_n1504__, new_new_n1505__,
    new_new_n1506__, new_new_n1507__, new_new_n1508__, new_new_n1509__,
    new_new_n1510__, new_new_n1511__, new_new_n1512__, new_new_n1513__,
    new_new_n1514__, new_new_n1515__, new_new_n1516__, new_new_n1517__,
    new_new_n1518__, new_new_n1519__, new_new_n1520__, new_new_n1521__,
    new_new_n1522__, new_new_n1523__, new_new_n1524__, new_new_n1525__,
    new_new_n1526__, new_new_n1527__, new_new_n1528__, new_new_n1529__,
    new_new_n1530__, new_new_n1531__, new_new_n1532__, new_new_n1533__,
    new_new_n1534__, new_new_n1535__, new_new_n1536__, new_new_n1537__,
    new_new_n1538__, new_new_n1539__, new_new_n1540__, new_new_n1541__,
    new_new_n1542__, new_new_n1543__, new_new_n1544__, new_new_n1545__,
    new_new_n1546__, new_new_n1547__, new_new_n1548__, new_new_n1549__,
    new_new_n1550__, new_new_n1551__, new_new_n1552__, new_new_n1553__,
    new_new_n1554__, new_new_n1555__, new_new_n1556__, new_new_n1557__,
    new_new_n1558__, new_new_n1559__, new_new_n1560__, new_new_n1561__,
    new_new_n1562__, new_new_n1563__, new_new_n1564__, new_new_n1565__,
    new_new_n1566__, new_new_n1567__, new_new_n1568__, new_new_n1569__,
    new_new_n1570__, new_new_n1571__, new_new_n1572__, new_new_n1573__,
    new_new_n1574__, new_new_n1575__, new_new_n1576__, new_new_n1577__,
    new_new_n1578__, new_new_n1579__, new_new_n1580__, new_new_n1581__,
    new_new_n1582__, new_new_n1583__, new_new_n1584__, new_new_n1585__,
    new_new_n1586__, new_new_n1587__, new_new_n1588__, new_new_n1589__,
    new_new_n1590__, new_new_n1591__, new_new_n1592__, new_new_n1593__,
    new_new_n1594__, new_new_n1595__, new_new_n1596__, new_new_n1597__,
    new_new_n1598__, new_new_n1599__, new_new_n1600__, new_new_n1601__,
    new_new_n1602__, new_new_n1603__, new_new_n1604__, new_new_n1605__,
    new_new_n1606__, new_new_n1607__, new_new_n1608__, new_new_n1609__,
    new_new_n1610__, new_new_n1611__, new_new_n1612__, new_new_n1613__,
    new_new_n1614__, new_new_n1615__, new_new_n1616__, new_new_n1617__,
    new_new_n1618__, new_new_n1619__, new_new_n1620__, new_new_n1621__,
    new_new_n1622__, new_new_n1623__, new_new_n1624__, new_new_n1625__,
    new_new_n1626__, new_new_n1627__, new_new_n1628__, new_new_n1629__,
    new_new_n1630__, new_new_n1631__, new_new_n1632__, new_new_n1633__,
    new_new_n1634__, new_new_n1635__, new_new_n1636__, new_new_n1637__,
    new_new_n1638__, new_new_n1639__, new_new_n1640__, new_new_n1641__,
    new_new_n1642__, new_new_n1643__, new_new_n1644__, new_new_n1645__,
    new_new_n1646__, new_new_n1647__, new_new_n1648__, new_new_n1649__,
    new_new_n1650__, new_new_n1651__, new_new_n1652__, new_new_n1653__,
    new_new_n1654__, new_new_n1655__, new_new_n1656__, new_new_n1657__,
    new_new_n1658__, new_new_n1659__, new_new_n1660__, new_new_n1661__,
    new_new_n1662__, new_new_n1663__, new_new_n1664__, new_new_n1665__,
    new_new_n1666__, new_new_n1667__, new_new_n1668__, new_new_n1669__,
    new_new_n1670__, new_new_n1671__, new_new_n1672__, new_new_n1673__,
    new_new_n1674__, new_new_n1675__, new_new_n1676__, new_new_n1677__,
    new_new_n1678__, new_new_n1679__, new_new_n1680__, new_new_n1681__,
    new_new_n1682__, new_new_n1683__, new_new_n1684__, new_new_n1685__,
    new_new_n1686__, new_new_n1687__, new_new_n1688__, new_new_n1689__,
    new_new_n1690__, new_new_n1691__, new_new_n1692__, new_new_n1693__,
    new_new_n1694__, new_new_n1695__, new_new_n1696__, new_new_n1697__,
    new_new_n1698__, new_new_n1699__, new_new_n1700__, new_new_n1701__,
    new_new_n1702__, new_new_n1703__, new_new_n1704__, new_new_n1705__,
    new_new_n1706__, new_new_n1707__, new_new_n1708__, new_new_n1709__,
    new_new_n1710__, new_new_n1711__, new_new_n1712__, new_new_n1713__,
    new_new_n1714__, new_new_n1715__, new_new_n1716__, new_new_n1717__,
    new_new_n1718__, new_new_n1719__, new_new_n1720__, new_new_n1721__,
    new_new_n1722__, new_new_n1723__, new_new_n1724__, new_new_n1725__,
    new_new_n1726__, new_new_n1727__, new_new_n1728__, new_new_n1729__,
    new_new_n1730__, new_new_n1731__, new_new_n1732__, new_new_n1733__,
    new_new_n1734__, new_new_n1735__, new_new_n1736__, new_new_n1737__,
    new_new_n1738__, new_new_n1739__, new_new_n1740__, new_new_n1741__,
    new_new_n1742__, new_new_n1743__, new_new_n1744__, new_new_n1745__,
    new_new_n1746__, n2688, n2691, n2694, n2697, n2700, n2703, n2706,
    n2709, n2712, n2715, n2718, n2721, n2724, n2727, n2730, n2733, n2736,
    n2739, n2742, n2745, n2748, n2751, n2754, n2757, n2760, n2763, n2766,
    n2769, n2772, n2775, n2778, n2781, n2784, n2787, n2790, n2793, n2796,
    n2799, n2802, n2805, n2808, n2811, n2814, n2817, n2820, n2823, n2826,
    n2829, n2832, n2835, n2838, n2841, n2844, n2847, n2850, n2853, n2856,
    n2859, n2862, n2865, n2868, n2871, n2874, n2877, n2880, n2883, n2886,
    n2889, n2892, n2895, n2898, n2901, n2904, n2907, n2910, n2913, n2916,
    n2919, n2922, n2925, n2928, n2931, n2934, n2937, n2940, n2943, n2946,
    n2949, n2952, n2955, n2958, n2961, n2964, n2967, n2970, n2973, n2976,
    n2979, n2982, n2985, n2988, n2991, n2994, n2997, n3000, n3003, n3006,
    n3009, n3012, n3015, n3018, n3021, n3024, n3027, n3030, n3033, n3036,
    n3039, n3042, n3045, n3048, n3051, n3054, n3057, n3060, n3063, n3066,
    n3069, n3072, n3075, n3078, n3081, n3084, n3087, n3090, n3093, n3096,
    n3099, n3102, n3105, n3108, n3111, n3114, n3117, n3120, n3123, n3126,
    n3129, n3132, n3135, n3138, n3141, n3144, n3147, n3150, n3153, n3156,
    n3159, n3162, n3165, n3168, n3171, n3174, n3177, n3180, n3183, n3186,
    n3189, n3192, n3195, n3198, n3201, n3204, n3207, n3210, n3213, n3216,
    n3219, n3222, n3225, n3228, n3231, n3234, n3237;
  buf1  g0000(.din(G1), .dout(new_new_n427__));
  buf1  g0001(.din(G2), .dout(new_new_n429__));
  buf1  g0002(.din(G3), .dout(new_new_n431__));
  buf1  g0003(.din(G4), .dout(new_new_n433__));
  buf1  g0004(.din(G5), .dout(new_new_n435__));
  buf1  g0005(.din(G6), .dout(new_new_n437__));
  buf1  g0006(.din(G7), .dout(new_new_n439__));
  buf1  g0007(.din(G8), .dout(new_new_n441__));
  buf1  g0008(.din(G9), .dout(new_new_n443__));
  buf1  g0009(.din(G10), .dout(new_new_n445__));
  buf1  g0010(.din(G11), .dout(new_new_n447__));
  buf1  g0011(.din(G12), .dout(new_new_n449__));
  buf1  g0012(.din(G13), .dout(new_new_n451__));
  buf1  g0013(.din(G14), .dout(new_new_n453__));
  buf1  g0014(.din(G15), .dout(new_new_n455__));
  buf1  g0015(.din(G16), .dout(new_new_n457__));
  buf1  g0016(.din(G17), .dout(new_new_n459__));
  buf1  g0017(.din(G18), .dout(new_new_n461__));
  buf1  g0018(.din(G19), .dout(new_new_n463__));
  buf1  g0019(.din(G20), .dout(new_new_n465__));
  buf1  g0020(.din(G21), .dout(new_new_n467__));
  buf1  g0021(.din(G22), .dout(new_new_n469__));
  buf1  g0022(.din(G23), .dout(new_new_n471__));
  buf1  g0023(.din(G24), .dout(new_new_n473__));
  buf1  g0024(.din(G25), .dout(new_new_n475__));
  buf1  g0025(.din(G26), .dout(new_new_n477__));
  buf1  g0026(.din(G27), .dout(new_new_n479__));
  buf1  g0027(.din(G28), .dout(new_new_n481__));
  buf1  g0028(.din(G29), .dout(new_new_n483__));
  buf1  g0029(.din(G30), .dout(new_new_n485__));
  buf1  g0030(.din(G31), .dout(new_new_n487__));
  buf1  g0031(.din(G32), .dout(new_new_n489__));
  buf1  g0032(.din(G33), .dout(new_new_n491__));
  buf1  g0033(.din(n940_lo), .dout(new_new_n493__));
  not1  g0034(.din(n940_lo), .dout(new_new_n494__));
  buf1  g0035(.din(n949_lo), .dout(new_new_n495__));
  not1  g0036(.din(n949_lo), .dout(new_new_n496__));
  buf1  g0037(.din(n961_lo), .dout(new_new_n497__));
  not1  g0038(.din(n961_lo), .dout(new_new_n498__));
  buf1  g0039(.din(n973_lo), .dout(new_new_n499__));
  not1  g0040(.din(n973_lo), .dout(new_new_n500__));
  buf1  g0041(.din(n976_lo), .dout(new_new_n501__));
  not1  g0042(.din(n976_lo), .dout(new_new_n502__));
  buf1  g0043(.din(n985_lo), .dout(new_new_n503__));
  not1  g0044(.din(n985_lo), .dout(new_new_n504__));
  buf1  g0045(.din(n988_lo), .dout(new_new_n505__));
  not1  g0046(.din(n988_lo), .dout(new_new_n506__));
  buf1  g0047(.din(n997_lo), .dout(new_new_n507__));
  not1  g0048(.din(n997_lo), .dout(new_new_n508__));
  buf1  g0049(.din(n1009_lo), .dout(new_new_n509__));
  not1  g0050(.din(n1009_lo), .dout(new_new_n510__));
  buf1  g0051(.din(n1021_lo), .dout(new_new_n511__));
  not1  g0052(.din(n1021_lo), .dout(new_new_n512__));
  buf1  g0053(.din(n1033_lo), .dout(new_new_n513__));
  not1  g0054(.din(n1033_lo), .dout(new_new_n514__));
  buf1  g0055(.din(n1045_lo), .dout(new_new_n515__));
  not1  g0056(.din(n1045_lo), .dout(new_new_n516__));
  buf1  g0057(.din(n1057_lo), .dout(new_new_n517__));
  not1  g0058(.din(n1057_lo), .dout(new_new_n518__));
  buf1  g0059(.din(n1060_lo), .dout(new_new_n519__));
  not1  g0060(.din(n1060_lo), .dout(new_new_n520__));
  buf1  g0061(.din(n1069_lo), .dout(new_new_n521__));
  not1  g0062(.din(n1069_lo), .dout(new_new_n522__));
  buf1  g0063(.din(n1081_lo), .dout(new_new_n523__));
  not1  g0064(.din(n1081_lo), .dout(new_new_n524__));
  buf1  g0065(.din(n1093_lo), .dout(new_new_n525__));
  not1  g0066(.din(n1093_lo), .dout(new_new_n526__));
  buf1  g0067(.din(n1105_lo), .dout(new_new_n527__));
  not1  g0068(.din(n1105_lo), .dout(new_new_n528__));
  buf1  g0069(.din(n1117_lo), .dout(new_new_n529__));
  not1  g0070(.din(n1117_lo), .dout(new_new_n530__));
  buf1  g0071(.din(n1120_lo), .dout(new_new_n531__));
  not1  g0072(.din(n1120_lo), .dout(new_new_n532__));
  buf1  g0073(.din(n1129_lo), .dout(new_new_n533__));
  not1  g0074(.din(n1129_lo), .dout(new_new_n534__));
  buf1  g0075(.din(n1132_lo), .dout(new_new_n535__));
  buf1  g0076(.din(n1156_lo), .dout(new_new_n537__));
  buf1  g0077(.din(n1168_lo), .dout(new_new_n539__));
  buf1  g0078(.din(n1180_lo), .dout(new_new_n541__));
  buf1  g0079(.din(n1189_lo), .dout(new_new_n543__));
  not1  g0080(.din(n1189_lo), .dout(new_new_n544__));
  buf1  g0081(.din(n1192_lo), .dout(new_new_n545__));
  buf1  g0082(.din(n1195_lo), .dout(new_new_n547__));
  not1  g0083(.din(n1195_lo), .dout(new_new_n548__));
  buf1  g0084(.din(n1201_lo), .dout(new_new_n549__));
  not1  g0085(.din(n1201_lo), .dout(new_new_n550__));
  buf1  g0086(.din(n1204_lo), .dout(new_new_n551__));
  not1  g0087(.din(n1204_lo), .dout(new_new_n552__));
  buf1  g0088(.din(n1228_lo), .dout(new_new_n553__));
  buf1  g0089(.din(n1231_lo), .dout(new_new_n555__));
  buf1  g0090(.din(n1234_lo), .dout(new_new_n557__));
  not1  g0091(.din(n1234_lo), .dout(new_new_n558__));
  buf1  g0092(.din(n1237_lo), .dout(new_new_n559__));
  not1  g0093(.din(n1237_lo), .dout(new_new_n560__));
  buf1  g0094(.din(n1240_lo), .dout(new_new_n561__));
  buf1  g0095(.din(n1243_lo), .dout(new_new_n563__));
  not1  g0096(.din(n1249_lo), .dout(new_new_n566__));
  buf1  g0097(.din(n1252_lo), .dout(new_new_n567__));
  buf1  g0098(.din(n1255_lo), .dout(new_new_n569__));
  buf1  g0099(.din(n1261_lo), .dout(new_new_n571__));
  buf1  g0100(.din(n1264_lo), .dout(new_new_n573__));
  buf1  g0101(.din(n1267_lo), .dout(new_new_n575__));
  not1  g0102(.din(n1267_lo), .dout(new_new_n576__));
  buf1  g0103(.din(n1273_lo), .dout(new_new_n577__));
  buf1  g0104(.din(n1276_lo), .dout(new_new_n579__));
  buf1  g0105(.din(n1279_lo), .dout(new_new_n581__));
  buf1  g0106(.din(n1282_lo), .dout(new_new_n583__));
  buf1  g0107(.din(n1285_lo), .dout(new_new_n585__));
  not1  g0108(.din(n1285_lo), .dout(new_new_n586__));
  buf1  g0109(.din(n1288_lo), .dout(new_new_n587__));
  buf1  g0110(.din(n1291_lo), .dout(new_new_n589__));
  buf1  g0111(.din(n1294_lo), .dout(new_new_n591__));
  buf1  g0112(.din(n1297_lo), .dout(new_new_n593__));
  not1  g0113(.din(n1297_lo), .dout(new_new_n594__));
  buf1  g0114(.din(n1300_lo), .dout(new_new_n595__));
  buf1  g0115(.din(n1303_lo), .dout(new_new_n597__));
  not1  g0116(.din(n1303_lo), .dout(new_new_n598__));
  buf1  g0117(.din(n1309_lo), .dout(new_new_n599__));
  not1  g0118(.din(n1309_lo), .dout(new_new_n600__));
  buf1  g0119(.din(n1312_lo), .dout(new_new_n601__));
  buf1  g0120(.din(n1315_lo), .dout(new_new_n603__));
  buf1  g0121(.din(n1318_lo), .dout(new_new_n605__));
  buf1  g0122(.din(n1321_lo), .dout(new_new_n607__));
  buf1  g0123(.din(n1333_lo), .dout(new_new_n609__));
  not1  g0124(.din(n1333_lo), .dout(new_new_n610__));
  not1  g0125(.din(n1225_o2), .dout(new_new_n612__));
  buf1  g0126(.din(n1229_o2), .dout(new_new_n613__));
  not1  g0127(.din(n1229_o2), .dout(new_new_n614__));
  buf1  g0128(.din(n1228_o2), .dout(new_new_n615__));
  buf1  g0129(.din(n1259_o2), .dout(new_new_n617__));
  not1  g0130(.din(n1272_o2), .dout(new_new_n620__));
  not1  g0131(.din(n1269_o2), .dout(new_new_n622__));
  buf1  g0132(.din(n1307_o2), .dout(new_new_n623__));
  not1  g0133(.din(n1307_o2), .dout(new_new_n624__));
  buf1  g0134(.din(n1201_o2), .dout(new_new_n625__));
  buf1  g0135(.din(n1202_o2), .dout(new_new_n627__));
  buf1  g0136(.din(n1203_o2), .dout(new_new_n629__));
  buf1  g0137(.din(n1204_o2), .dout(new_new_n631__));
  buf1  g0138(.din(n622_o2), .dout(new_new_n633__));
  not1  g0139(.din(n622_o2), .dout(new_new_n634__));
  not1  g0140(.din(n1205_o2), .dout(new_new_n636__));
  buf1  g0141(.din(n1206_o2), .dout(new_new_n637__));
  buf1  g0142(.din(n497_o2), .dout(new_new_n639__));
  not1  g0143(.din(n497_o2), .dout(new_new_n640__));
  buf1  g0144(.din(n1212_o2), .dout(new_new_n641__));
  buf1  g0145(.din(n1213_o2), .dout(new_new_n643__));
  buf1  g0146(.din(n1214_o2), .dout(new_new_n645__));
  buf1  g0147(.din(n1215_o2), .dout(new_new_n647__));
  buf1  g0148(.din(n1216_o2), .dout(new_new_n649__));
  buf1  g0149(.din(n1217_o2), .dout(new_new_n651__));
  buf1  g0150(.din(n1218_o2), .dout(new_new_n653__));
  buf1  g0151(.din(n1219_o2), .dout(new_new_n655__));
  buf1  g0152(.din(n1242_o2), .dout(new_new_n657__));
  buf1  g0153(.din(n1243_o2), .dout(new_new_n659__));
  buf1  g0154(.din(n1273_o2), .dout(new_new_n661__));
  buf1  g0155(.din(n1274_o2), .dout(new_new_n663__));
  buf1  g0156(.din(n1275_o2), .dout(new_new_n665__));
  not1  g0157(.din(n1276_o2), .dout(new_new_n668__));
  not1  g0158(.din(n1277_o2), .dout(new_new_n670__));
  buf1  g0159(.din(n1286_o2), .dout(new_new_n671__));
  not1  g0160(.din(n1286_o2), .dout(new_new_n672__));
  buf1  g0161(.din(n1299_o2), .dout(new_new_n673__));
  not1  g0162(.din(n1299_o2), .dout(new_new_n674__));
  buf1  g0163(.din(n601_o2), .dout(new_new_n675__));
  not1  g0164(.din(n601_o2), .dout(new_new_n676__));
  buf1  g0165(.din(n625_o2), .dout(new_new_n677__));
  not1  g0166(.din(n625_o2), .dout(new_new_n678__));
  buf1  g0167(.din(n463_o2), .dout(new_new_n679__));
  not1  g0168(.din(n463_o2), .dout(new_new_n680__));
  buf1  g0169(.din(lo082_buf_o2), .dout(new_new_n681__));
  buf1  g0170(.din(n455_o2), .dout(new_new_n683__));
  not1  g0171(.din(n455_o2), .dout(new_new_n684__));
  buf1  g0172(.din(n642_o2), .dout(new_new_n685__));
  not1  g0173(.din(n642_o2), .dout(new_new_n686__));
  buf1  g0174(.din(n459_o2), .dout(new_new_n687__));
  buf1  g0175(.din(n501_o2), .dout(new_new_n689__));
  not1  g0176(.din(n501_o2), .dout(new_new_n690__));
  buf1  g0177(.din(n599_o2), .dout(new_new_n691__));
  not1  g0178(.din(n599_o2), .dout(new_new_n692__));
  buf1  g0179(.din(n485_o2), .dout(new_new_n693__));
  not1  g0180(.din(n485_o2), .dout(new_new_n694__));
  buf1  g0181(.din(lo086_buf_o2), .dout(new_new_n695__));
  buf1  g0182(.din(lo122_buf_o2), .dout(new_new_n697__));
  not1  g0183(.din(lo122_buf_o2), .dout(new_new_n698__));
  buf1  g0184(.din(n502_o2), .dout(new_new_n699__));
  not1  g0185(.din(n502_o2), .dout(new_new_n700__));
  buf1  g0186(.din(n627_o2), .dout(new_new_n701__));
  not1  g0187(.din(n627_o2), .dout(new_new_n702__));
  buf1  g0188(.din(lo038_buf_o2), .dout(new_new_n703__));
  buf1  g0189(.din(lo046_buf_o2), .dout(new_new_n705__));
  buf1  g0190(.din(lo050_buf_o2), .dout(new_new_n707__));
  not1  g0191(.din(lo050_buf_o2), .dout(new_new_n708__));
  buf1  g0192(.din(lo058_buf_o2), .dout(new_new_n709__));
  buf1  g0193(.din(lo070_buf_o2), .dout(new_new_n711__));
  buf1  g0194(.din(lo094_buf_o2), .dout(new_new_n713__));
  not1  g0195(.din(n462_o2), .dout(new_new_n716__));
  buf1  g0196(.din(lo006_buf_o2), .dout(new_new_n717__));
  not1  g0197(.din(lo006_buf_o2), .dout(new_new_n718__));
  buf1  g0198(.din(lo010_buf_o2), .dout(new_new_n719__));
  buf1  g0199(.din(lo022_buf_o2), .dout(new_new_n721__));
  buf1  g0200(.din(lo026_buf_o2), .dout(new_new_n723__));
  buf1  g0201(.din(lo030_buf_o2), .dout(new_new_n725__));
  not1  g0202(.din(lo030_buf_o2), .dout(new_new_n726__));
  buf1  g0203(.din(lo034_buf_o2), .dout(new_new_n727__));
  not1  g0204(.din(lo034_buf_o2), .dout(new_new_n728__));
  buf1  g0205(.din(lo054_buf_o2), .dout(new_new_n729__));
  not1  g0206(.din(lo054_buf_o2), .dout(new_new_n730__));
  buf1  g0207(.din(lo130_buf_o2), .dout(new_new_n731__));
  not1  g0208(.din(lo130_buf_o2), .dout(new_new_n732__));
  buf1  g0209(.din(n547_o2), .dout(new_new_n733__));
  buf1  g0210(.din(n424_inv), .dout(new_new_n735__));
  buf1  g0211(.din(n617_o2), .dout(new_new_n737__));
  buf1  g0212(.din(lo042_buf_o2), .dout(new_new_n739__));
  buf1  g0213(.din(lo062_buf_o2), .dout(new_new_n741__));
  buf1  g0214(.din(lo110_buf_o2), .dout(new_new_n743__));
  buf1  g0215(.din(n733_o2), .dout(new_new_n745__));
  not1  g0216(.din(n733_o2), .dout(new_new_n746__));
  buf1  g0217(.din(n734_o2), .dout(new_new_n747__));
  not1  g0218(.din(n734_o2), .dout(new_new_n748__));
  buf1  g0219(.din(n570_o2), .dout(new_new_n749__));
  buf1  g0220(.din(n461_o2), .dout(new_new_n751__));
  not1  g0221(.din(n461_o2), .dout(new_new_n752__));
  buf1  g0222(.din(n644_o2), .dout(new_new_n753__));
  not1  g0223(.din(n644_o2), .dout(new_new_n754__));
  buf1  g0224(.din(n628_o2), .dout(new_new_n755__));
  not1  g0225(.din(n628_o2), .dout(new_new_n756__));
  buf1  g0226(.din(n528_o2), .dout(new_new_n757__));
  buf1  g0227(.din(n460_inv), .dout(new_new_n759__));
  buf1  g0228(.din(lo002_buf_o2), .dout(new_new_n761__));
  not1  g0229(.din(lo002_buf_o2), .dout(new_new_n762__));
  buf1  g0230(.din(lo014_buf_o2), .dout(new_new_n763__));
  not1  g0231(.din(lo014_buf_o2), .dout(new_new_n764__));
  buf1  g0232(.din(lo018_buf_o2), .dout(new_new_n765__));
  buf1  g0233(.din(lo078_buf_o2), .dout(new_new_n767__));
  buf1  g0234(.din(lo090_buf_o2), .dout(new_new_n769__));
  not1  g0235(.din(lo090_buf_o2), .dout(new_new_n770__));
  buf1  g0236(.din(n513_o2), .dout(new_new_n771__));
  buf1  g0237(.din(lo102_buf_o2), .dout(new_new_n773__));
  not1  g0238(.din(lo102_buf_o2), .dout(new_new_n774__));
  buf1  g0239(.din(lo106_buf_o2), .dout(new_new_n775__));
  not1  g0240(.din(lo106_buf_o2), .dout(new_new_n776__));
  buf1  g0241(.din(n600_o2), .dout(new_new_n777__));
  not1  g0242(.din(n600_o2), .dout(new_new_n778__));
  buf1  g0243(.din(n529_o2), .dout(new_new_n779__));
  not1  g0244(.din(n529_o2), .dout(new_new_n780__));
  buf1  g0245(.din(n593_o2), .dout(new_new_n781__));
  not1  g0246(.din(n593_o2), .dout(new_new_n782__));
  buf1  g0247(.din(lo066_buf_o2), .dout(new_new_n783__));
  not1  g0248(.din(n549_o2), .dout(new_new_n786__));
  not1  g0249(.din(n550_o2), .dout(new_new_n788__));
  buf1  g0250(.din(n571_o2), .dout(new_new_n789__));
  not1  g0251(.din(n572_o2), .dout(new_new_n792__));
  buf1  g0252(.din(n495_o2), .dout(new_new_n793__));
  not1  g0253(.din(n495_o2), .dout(new_new_n794__));
  buf1  g0254(.din(n496_o2), .dout(new_new_n795__));
  not1  g0255(.din(n496_o2), .dout(new_new_n796__));
  buf1  g0256(.din(n620_o2), .dout(new_new_n797__));
  not1  g0257(.din(n620_o2), .dout(new_new_n798__));
  buf1  g0258(.din(n482_o2), .dout(new_new_n799__));
  not1  g0259(.din(n482_o2), .dout(new_new_n800__));
  buf1  g0260(.din(lo081_buf_o2), .dout(new_new_n801__));
  not1  g0261(.din(lo081_buf_o2), .dout(new_new_n802__));
  buf1  g0262(.din(n576_o2), .dout(new_new_n803__));
  not1  g0263(.din(n576_o2), .dout(new_new_n804__));
  buf1  g0264(.din(n520_o2), .dout(new_new_n805__));
  not1  g0265(.din(n520_o2), .dout(new_new_n806__));
  buf1  g0266(.din(n521_o2), .dout(new_new_n807__));
  not1  g0267(.din(n521_o2), .dout(new_new_n808__));
  buf1  g0268(.din(n562_o2), .dout(new_new_n809__));
  not1  g0269(.din(n562_o2), .dout(new_new_n810__));
  buf1  g0270(.din(n508_o2), .dout(new_new_n811__));
  not1  g0271(.din(n508_o2), .dout(new_new_n812__));
  buf1  g0272(.din(n509_o2), .dout(new_new_n813__));
  not1  g0273(.din(n509_o2), .dout(new_new_n814__));
  buf1  g0274(.din(lo074_buf_o2), .dout(new_new_n815__));
  not1  g0275(.din(lo074_buf_o2), .dout(new_new_n816__));
  buf1  g0276(.din(n539_o2), .dout(new_new_n817__));
  not1  g0277(.din(n539_o2), .dout(new_new_n818__));
  buf1  g0278(.din(n536_o2), .dout(new_new_n819__));
  not1  g0279(.din(n536_o2), .dout(new_new_n820__));
  buf1  g0280(.din(n516_o2), .dout(new_new_n821__));
  not1  g0281(.din(n516_o2), .dout(new_new_n822__));
  buf1  g0282(.din(n491_o2), .dout(new_new_n823__));
  not1  g0283(.din(n491_o2), .dout(new_new_n824__));
  buf1  g0284(.din(n557_o2), .dout(new_new_n825__));
  not1  g0285(.din(n557_o2), .dout(new_new_n826__));
  buf1  g0286(.din(n586_o2), .dout(new_new_n827__));
  not1  g0287(.din(n586_o2), .dout(new_new_n828__));
  buf1  g0288(.din(n483_o2), .dout(new_new_n829__));
  not1  g0289(.din(n483_o2), .dout(new_new_n830__));
  buf1  g0290(.din(n484_o2), .dout(new_new_n831__));
  not1  g0291(.din(n484_o2), .dout(new_new_n832__));
  buf1  g0292(.din(lo004_buf_o2), .dout(new_new_n833__));
  not1  g0293(.din(lo004_buf_o2), .dout(new_new_n834__));
  buf1  g0294(.din(lo008_buf_o2), .dout(new_new_n835__));
  not1  g0295(.din(lo008_buf_o2), .dout(new_new_n836__));
  buf1  g0296(.din(lo020_buf_o2), .dout(new_new_n837__));
  not1  g0297(.din(lo020_buf_o2), .dout(new_new_n838__));
  buf1  g0298(.din(lo024_buf_o2), .dout(new_new_n839__));
  not1  g0299(.din(lo024_buf_o2), .dout(new_new_n840__));
  buf1  g0300(.din(lo028_buf_o2), .dout(new_new_n841__));
  not1  g0301(.din(lo028_buf_o2), .dout(new_new_n842__));
  buf1  g0302(.din(lo032_buf_o2), .dout(new_new_n843__));
  not1  g0303(.din(lo032_buf_o2), .dout(new_new_n844__));
  buf1  g0304(.din(lo052_buf_o2), .dout(new_new_n845__));
  not1  g0305(.din(lo052_buf_o2), .dout(new_new_n846__));
  buf1  g0306(.din(lo128_buf_o2), .dout(new_new_n847__));
  not1  g0307(.din(lo128_buf_o2), .dout(new_new_n848__));
  buf1  g0308(.din(lo037_buf_o2), .dout(new_new_n849__));
  not1  g0309(.din(lo037_buf_o2), .dout(new_new_n850__));
  buf1  g0310(.din(lo045_buf_o2), .dout(new_new_n851__));
  not1  g0311(.din(lo045_buf_o2), .dout(new_new_n852__));
  buf1  g0312(.din(lo049_buf_o2), .dout(new_new_n853__));
  not1  g0313(.din(lo049_buf_o2), .dout(new_new_n854__));
  buf1  g0314(.din(lo057_buf_o2), .dout(new_new_n855__));
  not1  g0315(.din(lo057_buf_o2), .dout(new_new_n856__));
  buf1  g0316(.din(lo069_buf_o2), .dout(new_new_n857__));
  not1  g0317(.din(lo069_buf_o2), .dout(new_new_n858__));
  buf1  g0318(.din(lo093_buf_o2), .dout(new_new_n859__));
  not1  g0319(.din(lo093_buf_o2), .dout(new_new_n860__));
  and1  g0320(.dina(new_new_n1464__), .dinb(new_new_n1465__), .dout(new_new_n861__));
  or1   g0321(.dina(new_new_n1466__), .dinb(new_new_n1467__), .dout(new_new_n862__));
  and1  g0322(.dina(new_new_n496__), .dinb(new_new_n1470__), .dout(new_new_n863__));
  and1  g0323(.dina(new_new_n495__), .dinb(new_new_n1476__), .dout(new_new_n864__));
  or1   g0324(.dina(new_new_n863__), .dinb(new_new_n864__), .dout(new_new_n865__));
  and1  g0325(.dina(new_new_n498__), .dinb(new_new_n1470__), .dout(new_new_n866__));
  and1  g0326(.dina(new_new_n497__), .dinb(new_new_n1476__), .dout(new_new_n867__));
  or1   g0327(.dina(new_new_n866__), .dinb(new_new_n867__), .dout(new_new_n868__));
  and1  g0328(.dina(new_new_n500__), .dinb(new_new_n1471__), .dout(new_new_n869__));
  and1  g0329(.dina(new_new_n499__), .dinb(new_new_n1477__), .dout(new_new_n870__));
  or1   g0330(.dina(new_new_n869__), .dinb(new_new_n870__), .dout(new_new_n871__));
  and1  g0331(.dina(new_new_n504__), .dinb(new_new_n1471__), .dout(new_new_n872__));
  and1  g0332(.dina(new_new_n503__), .dinb(new_new_n1477__), .dout(new_new_n873__));
  or1   g0333(.dina(new_new_n872__), .dinb(new_new_n873__), .dout(new_new_n874__));
  and1  g0334(.dina(new_new_n1481__), .dinb(new_new_n1465__), .dout(new_new_n875__));
  or1   g0335(.dina(new_new_n1483__), .dinb(new_new_n1467__), .dout(new_new_n876__));
  and1  g0336(.dina(new_new_n518__), .dinb(new_new_n1486__), .dout(new_new_n877__));
  and1  g0337(.dina(new_new_n517__), .dinb(new_new_n1491__), .dout(new_new_n878__));
  or1   g0338(.dina(new_new_n877__), .dinb(new_new_n878__), .dout(new_new_n879__));
  and1  g0339(.dina(new_new_n530__), .dinb(new_new_n1486__), .dout(new_new_n880__));
  and1  g0340(.dina(new_new_n529__), .dinb(new_new_n1491__), .dout(new_new_n881__));
  or1   g0341(.dina(new_new_n880__), .dinb(new_new_n881__), .dout(new_new_n882__));
  and1  g0342(.dina(new_new_n534__), .dinb(new_new_n1487__), .dout(new_new_n883__));
  and1  g0343(.dina(new_new_n533__), .dinb(new_new_n1492__), .dout(new_new_n884__));
  or1   g0344(.dina(new_new_n883__), .dinb(new_new_n884__), .dout(new_new_n885__));
  and1  g0345(.dina(new_new_n679__), .dinb(new_new_n1494__), .dout(new_new_n886__));
  or1   g0346(.dina(new_new_n1495__), .dinb(new_new_n689__), .dout(new_new_n887__));
  and1  g0347(.dina(new_new_n701__), .dinb(new_new_n886__), .dout(new_new_n888__));
  or1   g0348(.dina(new_new_n702__), .dinb(new_new_n887__), .dout(new_new_n889__));
  and1  g0349(.dina(new_new_n1464__), .dinb(new_new_n1496__), .dout(new_new_n890__));
  or1   g0350(.dina(new_new_n1466__), .dinb(new_new_n1497__), .dout(new_new_n891__));
  and1  g0351(.dina(new_new_n508__), .dinb(new_new_n1499__), .dout(new_new_n892__));
  and1  g0352(.dina(new_new_n507__), .dinb(new_new_n1502__), .dout(new_new_n893__));
  or1   g0353(.dina(new_new_n892__), .dinb(new_new_n893__), .dout(new_new_n894__));
  and1  g0354(.dina(new_new_n510__), .dinb(new_new_n1499__), .dout(new_new_n895__));
  and1  g0355(.dina(new_new_n509__), .dinb(new_new_n1502__), .dout(new_new_n896__));
  or1   g0356(.dina(new_new_n895__), .dinb(new_new_n896__), .dout(new_new_n897__));
  and1  g0357(.dina(new_new_n512__), .dinb(new_new_n1500__), .dout(new_new_n898__));
  and1  g0358(.dina(new_new_n511__), .dinb(new_new_n1503__), .dout(new_new_n899__));
  or1   g0359(.dina(new_new_n898__), .dinb(new_new_n899__), .dout(new_new_n900__));
  and1  g0360(.dina(new_new_n514__), .dinb(new_new_n1500__), .dout(new_new_n901__));
  and1  g0361(.dina(new_new_n513__), .dinb(new_new_n1503__), .dout(new_new_n902__));
  or1   g0362(.dina(new_new_n901__), .dinb(new_new_n902__), .dout(new_new_n903__));
  and1  g0363(.dina(new_new_n1481__), .dinb(new_new_n1496__), .dout(new_new_n904__));
  or1   g0364(.dina(new_new_n1483__), .dinb(new_new_n1497__), .dout(new_new_n905__));
  and1  g0365(.dina(new_new_n515__), .dinb(new_new_n904__), .dout(new_new_n906__));
  and1  g0366(.dina(new_new_n516__), .dinb(new_new_n905__), .dout(new_new_n907__));
  or1   g0367(.dina(new_new_n906__), .dinb(new_new_n907__), .dout(new_new_n908__));
  and1  g0368(.dina(new_new_n675__), .dinb(new_new_n1480__), .dout(new_new_n909__));
  or1   g0369(.dina(new_new_n1504__), .dinb(new_new_n1482__), .dout(new_new_n910__));
  and1  g0370(.dina(new_new_n1505__), .dinb(new_new_n909__), .dout(new_new_n911__));
  or1   g0371(.dina(new_new_n678__), .dinb(new_new_n910__), .dout(new_new_n912__));
  and1  g0372(.dina(new_new_n700__), .dinb(new_new_n911__), .dout(new_new_n913__));
  or1   g0373(.dina(new_new_n699__), .dinb(new_new_n912__), .dout(new_new_n914__));
  and1  g0374(.dina(new_new_n1506__), .dinb(new_new_n913__), .dout(new_new_n915__));
  or1   g0375(.dina(new_new_n692__), .dinb(new_new_n914__), .dout(new_new_n916__));
  and1  g0376(.dina(new_new_n522__), .dinb(new_new_n1508__), .dout(new_new_n917__));
  and1  g0377(.dina(new_new_n521__), .dinb(new_new_n1511__), .dout(new_new_n918__));
  or1   g0378(.dina(new_new_n917__), .dinb(new_new_n918__), .dout(new_new_n919__));
  and1  g0379(.dina(new_new_n524__), .dinb(new_new_n1508__), .dout(new_new_n920__));
  and1  g0380(.dina(new_new_n523__), .dinb(new_new_n1511__), .dout(new_new_n921__));
  or1   g0381(.dina(new_new_n920__), .dinb(new_new_n921__), .dout(new_new_n922__));
  and1  g0382(.dina(new_new_n526__), .dinb(new_new_n1509__), .dout(new_new_n923__));
  and1  g0383(.dina(new_new_n525__), .dinb(new_new_n1512__), .dout(new_new_n924__));
  or1   g0384(.dina(new_new_n923__), .dinb(new_new_n924__), .dout(new_new_n925__));
  and1  g0385(.dina(new_new_n528__), .dinb(new_new_n1509__), .dout(new_new_n926__));
  and1  g0386(.dina(new_new_n527__), .dinb(new_new_n1512__), .dout(new_new_n927__));
  or1   g0387(.dina(new_new_n926__), .dinb(new_new_n927__), .dout(new_new_n928__));
  and1  g0388(.dina(new_new_n1473__), .dinb(new_new_n1487__), .dout(new_new_n929__));
  or1   g0389(.dina(new_new_n1479__), .dinb(new_new_n1492__), .dout(new_new_n930__));
  and1  g0390(.dina(new_new_n607__), .dinb(new_new_n1515__), .dout(new_new_n931__));
  and1  g0391(.dina(new_new_n1504__), .dinb(new_new_n1495__), .dout(new_new_n932__));
  and1  g0392(.dina(new_new_n1494__), .dinb(new_new_n932__), .dout(new_new_n933__));
  and1  g0393(.dina(new_new_n1505__), .dinb(new_new_n933__), .dout(new_new_n934__));
  and1  g0394(.dina(new_new_n1506__), .dinb(new_new_n934__), .dout(new_new_n935__));
  or1   g0395(.dina(new_new_n1519__), .dinb(new_new_n935__), .dout(new_new_n936__));
  or1   g0396(.dina(new_new_n931__), .dinb(new_new_n936__), .dout(new_new_n937__));
  and1  g0397(.dina(new_new_n1522__), .dinb(new_new_n633__), .dout(new_new_n938__));
  or1   g0398(.dina(new_new_n1525__), .dinb(new_new_n634__), .dout(new_new_n939__));
  and1  g0399(.dina(new_new_n1515__), .dinb(new_new_n938__), .dout(new_new_n940__));
  or1   g0400(.dina(new_new_n1527__), .dinb(new_new_n939__), .dout(new_new_n941__));
  and1  g0401(.dina(new_new_n624__), .dinb(new_new_n941__), .dout(new_new_n942__));
  and1  g0402(.dina(new_new_n623__), .dinb(new_new_n940__), .dout(new_new_n943__));
  or1   g0403(.dina(new_new_n942__), .dinb(new_new_n943__), .dout(new_new_n944__));
  and1  g0404(.dina(new_new_n1530__), .dinb(new_new_n944__), .dout(new_new_n945__));
  and1  g0405(.dina(new_new_n559__), .dinb(new_new_n1522__), .dout(new_new_n946__));
  or1   g0406(.dina(new_new_n560__), .dinb(new_new_n1525__), .dout(new_new_n947__));
  and1  g0407(.dina(new_new_n1516__), .dinb(new_new_n946__), .dout(new_new_n948__));
  or1   g0408(.dina(new_new_n1527__), .dinb(new_new_n947__), .dout(new_new_n949__));
  and1  g0409(.dina(new_new_n639__), .dinb(new_new_n949__), .dout(new_new_n950__));
  and1  g0410(.dina(new_new_n640__), .dinb(new_new_n948__), .dout(new_new_n951__));
  or1   g0411(.dina(new_new_n950__), .dinb(new_new_n951__), .dout(new_new_n952__));
  and1  g0412(.dina(new_new_n1530__), .dinb(new_new_n952__), .dout(new_new_n953__));
  and1  g0413(.dina(new_new_n571__), .dinb(new_new_n1521__), .dout(new_new_n954__));
  and1  g0414(.dina(new_new_n1516__), .dinb(new_new_n954__), .dout(new_new_n955__));
  or1   g0415(.dina(new_new_n622__), .dinb(new_new_n955__), .dout(new_new_n956__));
  and1  g0416(.dina(new_new_n1531__), .dinb(new_new_n956__), .dout(new_new_n957__));
  and1  g0417(.dina(new_new_n577__), .dinb(new_new_n1523__), .dout(new_new_n958__));
  and1  g0418(.dina(new_new_n1517__), .dinb(new_new_n958__), .dout(new_new_n959__));
  or1   g0419(.dina(new_new_n612__), .dinb(new_new_n959__), .dout(new_new_n960__));
  and1  g0420(.dina(new_new_n1531__), .dinb(new_new_n960__), .dout(new_new_n961__));
  and1  g0421(.dina(new_new_n1523__), .dinb(new_new_n617__), .dout(new_new_n962__));
  and1  g0422(.dina(new_new_n1517__), .dinb(new_new_n962__), .dout(new_new_n963__));
  or1   g0423(.dina(new_new_n615__), .dinb(new_new_n963__), .dout(new_new_n964__));
  and1  g0424(.dina(new_new_n1532__), .dinb(new_new_n964__), .dout(new_new_n965__));
  and1  g0425(.dina(new_new_n543__), .dinb(new_new_n585__), .dout(new_new_n966__));
  or1   g0426(.dina(new_new_n544__), .dinb(new_new_n586__), .dout(new_new_n967__));
  and1  g0427(.dina(new_new_n1533__), .dinb(new_new_n967__), .dout(new_new_n968__));
  or1   g0428(.dina(new_new_n1519__), .dinb(new_new_n966__), .dout(new_new_n969__));
  and1  g0429(.dina(new_new_n613__), .dinb(new_new_n683__), .dout(new_new_n970__));
  or1   g0430(.dina(new_new_n614__), .dinb(new_new_n684__), .dout(new_new_n971__));
  and1  g0431(.dina(new_new_n1479__), .dinb(new_new_n1534__), .dout(new_new_n972__));
  or1   g0432(.dina(new_new_n1473__), .dinb(new_new_n1535__), .dout(new_new_n973__));
  and1  g0433(.dina(new_new_n1472__), .dinb(new_new_n1535__), .dout(new_new_n974__));
  or1   g0434(.dina(new_new_n1478__), .dinb(new_new_n1534__), .dout(new_new_n975__));
  and1  g0435(.dina(new_new_n973__), .dinb(new_new_n975__), .dout(new_new_n976__));
  or1   g0436(.dina(new_new_n972__), .dinb(new_new_n974__), .dout(new_new_n977__));
  and1  g0437(.dina(new_new_n969__), .dinb(new_new_n977__), .dout(new_new_n978__));
  and1  g0438(.dina(new_new_n968__), .dinb(new_new_n976__), .dout(new_new_n979__));
  or1   g0439(.dina(new_new_n978__), .dinb(new_new_n979__), .dout(new_new_n980__));
  and1  g0440(.dina(new_new_n549__), .dinb(new_new_n593__), .dout(new_new_n981__));
  or1   g0441(.dina(new_new_n550__), .dinb(new_new_n594__), .dout(new_new_n982__));
  and1  g0442(.dina(new_new_n1533__), .dinb(new_new_n982__), .dout(new_new_n983__));
  or1   g0443(.dina(new_new_n1518__), .dinb(new_new_n981__), .dout(new_new_n984__));
  and1  g0444(.dina(new_new_n746__), .dinb(new_new_n748__), .dout(new_new_n985__));
  or1   g0445(.dina(new_new_n745__), .dinb(new_new_n747__), .dout(new_new_n986__));
  and1  g0446(.dina(new_new_n685__), .dinb(new_new_n986__), .dout(new_new_n987__));
  or1   g0447(.dina(new_new_n686__), .dinb(new_new_n985__), .dout(new_new_n988__));
  and1  g0448(.dina(new_new_n1493__), .dinb(new_new_n1536__), .dout(new_new_n989__));
  or1   g0449(.dina(new_new_n1488__), .dinb(new_new_n1537__), .dout(new_new_n990__));
  and1  g0450(.dina(new_new_n1488__), .dinb(new_new_n1537__), .dout(new_new_n991__));
  or1   g0451(.dina(new_new_n1493__), .dinb(new_new_n1536__), .dout(new_new_n992__));
  and1  g0452(.dina(new_new_n990__), .dinb(new_new_n992__), .dout(new_new_n993__));
  or1   g0453(.dina(new_new_n989__), .dinb(new_new_n991__), .dout(new_new_n994__));
  and1  g0454(.dina(new_new_n984__), .dinb(new_new_n994__), .dout(new_new_n995__));
  and1  g0455(.dina(new_new_n983__), .dinb(new_new_n993__), .dout(new_new_n996__));
  or1   g0456(.dina(new_new_n995__), .dinb(new_new_n996__), .dout(new_new_n997__));
  or1   g0457(.dina(new_new_n566__), .dinb(new_new_n1524__), .dout(new_new_n998__));
  or1   g0458(.dina(new_new_n1526__), .dinb(new_new_n998__), .dout(new_new_n999__));
  and1  g0459(.dina(new_new_n620__), .dinb(new_new_n999__), .dout(new_new_n1000__));
  and1  g0460(.dina(new_new_n1532__), .dinb(new_new_n1000__), .dout(new_new_n1001__));
  and1  g0461(.dina(new_new_n673__), .dinb(new_new_n777__), .dout(new_new_n1002__));
  or1   g0462(.dina(new_new_n674__), .dinb(new_new_n1538__), .dout(new_new_n1003__));
  and1  g0463(.dina(new_new_n794__), .dinb(new_new_n796__), .dout(new_new_n1004__));
  or1   g0464(.dina(new_new_n793__), .dinb(new_new_n795__), .dout(new_new_n1005__));
  or1   g0465(.dina(new_new_n636__), .dinb(new_new_n1538__), .dout(new_new_n1006__));
  and1  g0466(.dina(new_new_n1539__), .dinb(new_new_n798__), .dout(new_new_n1007__));
  or1   g0467(.dina(new_new_n1541__), .dinb(new_new_n1543__), .dout(new_new_n1008__));
  or1   g0468(.dina(new_new_n1544__), .dinb(new_new_n1008__), .dout(new_new_n1009__));
  or1   g0469(.dina(new_new_n1003__), .dinb(new_new_n1007__), .dout(new_new_n1010__));
  and1  g0470(.dina(new_new_n1009__), .dinb(new_new_n1010__), .dout(new_new_n1011__));
  or1   g0471(.dina(new_new_n668__), .dinb(new_new_n716__), .dout(new_new_n1012__));
  or1   g0472(.dina(new_new_n1545__), .dinb(new_new_n1547__), .dout(new_new_n1013__));
  or1   g0473(.dina(new_new_n1549__), .dinb(new_new_n1547__), .dout(new_new_n1014__));
  or1   g0474(.dina(new_new_n1550__), .dinb(new_new_n1548__), .dout(new_new_n1015__));
  and1  g0475(.dina(new_new_n1539__), .dinb(new_new_n1551__), .dout(new_new_n1016__));
  or1   g0476(.dina(new_new_n1541__), .dinb(new_new_n1004__), .dout(new_new_n1017__));
  or1   g0477(.dina(new_new_n1552__), .dinb(new_new_n1017__), .dout(new_new_n1018__));
  or1   g0478(.dina(new_new_n558__), .dinb(new_new_n1016__), .dout(new_new_n1019__));
  and1  g0479(.dina(new_new_n1018__), .dinb(new_new_n1019__), .dout(new_new_n1020__));
  or1   g0480(.dina(new_new_n1553__), .dinb(new_new_n780__), .dout(new_new_n1021__));
  and1  g0481(.dina(new_new_n786__), .dinb(new_new_n788__), .dout(new_new_n1022__));
  and1  g0482(.dina(new_new_n789__), .dinb(new_new_n792__), .dout(new_new_n1023__));
  and1  g0483(.dina(new_new_n1022__), .dinb(new_new_n1023__), .dout(new_new_n1024__));
  and1  g0484(.dina(new_new_n1021__), .dinb(new_new_n1024__), .dout(new_new_n1025__));
  or1   g0485(.dina(new_new_n774__), .dinb(new_new_n782__), .dout(new_new_n1026__));
  or1   g0486(.dina(new_new_n1554__), .dinb(new_new_n781__), .dout(new_new_n1027__));
  or1   g0487(.dina(new_new_n776__), .dinb(new_new_n779__), .dout(new_new_n1028__));
  and1  g0488(.dina(new_new_n1027__), .dinb(new_new_n1028__), .dout(new_new_n1029__));
  and1  g0489(.dina(new_new_n1026__), .dinb(new_new_n1029__), .dout(new_new_n1030__));
  and1  g0490(.dina(new_new_n1025__), .dinb(new_new_n1030__), .dout(new_new_n1031__));
  and1  g0491(.dina(new_new_n830__), .dinb(new_new_n832__), .dout(new_new_n1032__));
  or1   g0492(.dina(new_new_n829__), .dinb(new_new_n831__), .dout(new_new_n1033__));
  or1   g0493(.dina(new_new_n1555__), .dinb(new_new_n1556__), .dout(new_new_n1034__));
  or1   g0494(.dina(new_new_n1557__), .dinb(new_new_n1558__), .dout(new_new_n1035__));
  and1  g0495(.dina(new_new_n1559__), .dinb(new_new_n1035__), .dout(new_new_n1036__));
  or1   g0496(.dina(new_new_n1561__), .dinb(new_new_n1564__), .dout(new_new_n1037__));
  and1  g0497(.dina(new_new_n1565__), .dinb(new_new_n1566__), .dout(new_new_n1038__));
  or1   g0498(.dina(new_new_n1567__), .dinb(new_new_n1568__), .dout(new_new_n1039__));
  and1  g0499(.dina(new_new_n1567__), .dinb(new_new_n1568__), .dout(new_new_n1040__));
  or1   g0500(.dina(new_new_n1565__), .dinb(new_new_n1566__), .dout(new_new_n1041__));
  and1  g0501(.dina(new_new_n1039__), .dinb(new_new_n1041__), .dout(new_new_n1042__));
  or1   g0502(.dina(new_new_n1038__), .dinb(new_new_n1040__), .dout(new_new_n1043__));
  and1  g0503(.dina(new_new_n770__), .dinb(new_new_n1569__), .dout(new_new_n1044__));
  or1   g0504(.dina(new_new_n1564__), .dinb(new_new_n816__), .dout(new_new_n1045__));
  and1  g0505(.dina(new_new_n1571__), .dinb(new_new_n1044__), .dout(new_new_n1046__));
  or1   g0506(.dina(new_new_n1575__), .dinb(new_new_n1045__), .dout(new_new_n1047__));
  and1  g0507(.dina(new_new_n1043__), .dinb(new_new_n1047__), .dout(new_new_n1048__));
  and1  g0508(.dina(new_new_n1042__), .dinb(new_new_n1046__), .dout(new_new_n1049__));
  or1   g0509(.dina(new_new_n1048__), .dinb(new_new_n1049__), .dout(new_new_n1050__));
  and1  g0510(.dina(new_new_n1578__), .dinb(new_new_n1580__), .dout(new_new_n1051__));
  or1   g0511(.dina(new_new_n1582__), .dinb(new_new_n1584__), .dout(new_new_n1052__));
  and1  g0512(.dina(new_new_n1582__), .dinb(new_new_n1584__), .dout(new_new_n1053__));
  or1   g0513(.dina(new_new_n1578__), .dinb(new_new_n1580__), .dout(new_new_n1054__));
  and1  g0514(.dina(new_new_n1052__), .dinb(new_new_n1054__), .dout(new_new_n1055__));
  or1   g0515(.dina(new_new_n1051__), .dinb(new_new_n1053__), .dout(new_new_n1056__));
  and1  g0516(.dina(new_new_n1585__), .dinb(new_new_n1586__), .dout(new_new_n1057__));
  or1   g0517(.dina(new_new_n1588__), .dinb(new_new_n1589__), .dout(new_new_n1058__));
  and1  g0518(.dina(new_new_n1588__), .dinb(new_new_n1589__), .dout(new_new_n1059__));
  or1   g0519(.dina(new_new_n1585__), .dinb(new_new_n1586__), .dout(new_new_n1060__));
  and1  g0520(.dina(new_new_n1058__), .dinb(new_new_n1060__), .dout(new_new_n1061__));
  or1   g0521(.dina(new_new_n1057__), .dinb(new_new_n1059__), .dout(new_new_n1062__));
  or1   g0522(.dina(new_new_n1055__), .dinb(new_new_n1061__), .dout(new_new_n1063__));
  or1   g0523(.dina(new_new_n1056__), .dinb(new_new_n1062__), .dout(new_new_n1064__));
  and1  g0524(.dina(new_new_n1063__), .dinb(new_new_n1064__), .dout(new_new_n1065__));
  and1  g0525(.dina(new_new_n1591__), .dinb(new_new_n1593__), .dout(new_new_n1066__));
  or1   g0526(.dina(new_new_n1596__), .dinb(new_new_n1598__), .dout(new_new_n1067__));
  and1  g0527(.dina(new_new_n1596__), .dinb(new_new_n1598__), .dout(new_new_n1068__));
  or1   g0528(.dina(new_new_n1591__), .dinb(new_new_n1593__), .dout(new_new_n1069__));
  and1  g0529(.dina(new_new_n1067__), .dinb(new_new_n1069__), .dout(new_new_n1070__));
  or1   g0530(.dina(new_new_n1066__), .dinb(new_new_n1068__), .dout(new_new_n1071__));
  and1  g0531(.dina(new_new_n1600__), .dinb(new_new_n1603__), .dout(new_new_n1072__));
  or1   g0532(.dina(new_new_n1606__), .dinb(new_new_n1608__), .dout(new_new_n1073__));
  and1  g0533(.dina(new_new_n1606__), .dinb(new_new_n1608__), .dout(new_new_n1074__));
  or1   g0534(.dina(new_new_n1600__), .dinb(new_new_n1603__), .dout(new_new_n1075__));
  and1  g0535(.dina(new_new_n1073__), .dinb(new_new_n1075__), .dout(new_new_n1076__));
  or1   g0536(.dina(new_new_n1072__), .dinb(new_new_n1074__), .dout(new_new_n1077__));
  and1  g0537(.dina(new_new_n1610__), .dinb(new_new_n1611__), .dout(new_new_n1078__));
  or1   g0538(.dina(new_new_n1612__), .dinb(new_new_n1613__), .dout(new_new_n1079__));
  and1  g0539(.dina(new_new_n1612__), .dinb(new_new_n1613__), .dout(new_new_n1080__));
  or1   g0540(.dina(new_new_n1610__), .dinb(new_new_n1611__), .dout(new_new_n1081__));
  and1  g0541(.dina(new_new_n1079__), .dinb(new_new_n1081__), .dout(new_new_n1082__));
  or1   g0542(.dina(new_new_n1078__), .dinb(new_new_n1080__), .dout(new_new_n1083__));
  and1  g0543(.dina(new_new_n672__), .dinb(new_new_n693__), .dout(new_new_n1084__));
  and1  g0544(.dina(new_new_n671__), .dinb(new_new_n694__), .dout(new_new_n1085__));
  and1  g0545(.dina(new_new_n1569__), .dinb(new_new_n1614__), .dout(new_new_n1086__));
  and1  g0546(.dina(new_new_n637__), .dinb(new_new_n670__), .dout(new_new_n1087__));
  or1   g0547(.dina(new_new_n1542__), .dinb(new_new_n1615__), .dout(new_new_n1088__));
  or1   g0548(.dina(new_new_n1616__), .dinb(new_new_n1617__), .dout(new_new_n1089__));
  or1   g0549(.dina(new_new_n1618__), .dinb(new_new_n1615__), .dout(new_new_n1090__));
  and1  g0550(.dina(new_new_n1089__), .dinb(new_new_n1619__), .dout(new_new_n1091__));
  or1   g0551(.dina(new_new_n1620__), .dinb(new_new_n1617__), .dout(new_new_n1092__));
  and1  g0552(.dina(new_new_n1619__), .dinb(new_new_n1092__), .dout(new_new_n1093__));
  and1  g0553(.dina(new_new_n1621__), .dinb(new_new_n1622__), .dout(new_new_n1094__));
  and1  g0554(.dina(new_new_n812__), .dinb(new_new_n814__), .dout(new_new_n1095__));
  or1   g0555(.dina(new_new_n811__), .dinb(new_new_n813__), .dout(new_new_n1096__));
  and1  g0556(.dina(new_new_n1583__), .dinb(new_new_n1623__), .dout(new_new_n1097__));
  or1   g0557(.dina(new_new_n1579__), .dinb(new_new_n1624__), .dout(new_new_n1098__));
  and1  g0558(.dina(new_new_n1579__), .dinb(new_new_n1624__), .dout(new_new_n1099__));
  or1   g0559(.dina(new_new_n1583__), .dinb(new_new_n1623__), .dout(new_new_n1100__));
  and1  g0560(.dina(new_new_n1098__), .dinb(new_new_n1100__), .dout(new_new_n1101__));
  or1   g0561(.dina(new_new_n1097__), .dinb(new_new_n1099__), .dout(new_new_n1102__));
  and1  g0562(.dina(new_new_n806__), .dinb(new_new_n808__), .dout(new_new_n1103__));
  or1   g0563(.dina(new_new_n805__), .dinb(new_new_n807__), .dout(new_new_n1104__));
  and1  g0564(.dina(new_new_n1625__), .dinb(new_new_n1626__), .dout(new_new_n1105__));
  or1   g0565(.dina(new_new_n1628__), .dinb(new_new_n1629__), .dout(new_new_n1106__));
  and1  g0566(.dina(new_new_n1628__), .dinb(new_new_n1629__), .dout(new_new_n1107__));
  or1   g0567(.dina(new_new_n1625__), .dinb(new_new_n1626__), .dout(new_new_n1108__));
  and1  g0568(.dina(new_new_n1106__), .dinb(new_new_n1108__), .dout(new_new_n1109__));
  or1   g0569(.dina(new_new_n1105__), .dinb(new_new_n1107__), .dout(new_new_n1110__));
  and1  g0570(.dina(new_new_n1102__), .dinb(new_new_n1109__), .dout(new_new_n1111__));
  and1  g0571(.dina(new_new_n1101__), .dinb(new_new_n1110__), .dout(new_new_n1112__));
  or1   g0572(.dina(new_new_n1111__), .dinb(new_new_n1112__), .dout(new_new_n1113__));
  and1  g0573(.dina(new_new_n1571__), .dinb(new_new_n803__), .dout(new_new_n1114__));
  or1   g0574(.dina(new_new_n1575__), .dinb(new_new_n804__), .dout(new_new_n1115__));
  and1  g0575(.dina(new_new_n1631__), .dinb(new_new_n1632__), .dout(new_new_n1116__));
  or1   g0576(.dina(new_new_n1633__), .dinb(new_new_n1634__), .dout(new_new_n1117__));
  and1  g0577(.dina(new_new_n1633__), .dinb(new_new_n1634__), .dout(new_new_n1118__));
  or1   g0578(.dina(new_new_n1631__), .dinb(new_new_n1632__), .dout(new_new_n1119__));
  and1  g0579(.dina(new_new_n1117__), .dinb(new_new_n1119__), .dout(new_new_n1120__));
  or1   g0580(.dina(new_new_n1116__), .dinb(new_new_n1118__), .dout(new_new_n1121__));
  and1  g0581(.dina(new_new_n1594__), .dinb(new_new_n1636__), .dout(new_new_n1122__));
  or1   g0582(.dina(new_new_n1599__), .dinb(new_new_n1638__), .dout(new_new_n1123__));
  and1  g0583(.dina(new_new_n1599__), .dinb(new_new_n1638__), .dout(new_new_n1124__));
  or1   g0584(.dina(new_new_n1594__), .dinb(new_new_n1636__), .dout(new_new_n1125__));
  and1  g0585(.dina(new_new_n1123__), .dinb(new_new_n1125__), .dout(new_new_n1126__));
  or1   g0586(.dina(new_new_n1122__), .dinb(new_new_n1124__), .dout(new_new_n1127__));
  and1  g0587(.dina(new_new_n1120__), .dinb(new_new_n1127__), .dout(new_new_n1128__));
  and1  g0588(.dina(new_new_n1121__), .dinb(new_new_n1126__), .dout(new_new_n1129__));
  or1   g0589(.dina(new_new_n1128__), .dinb(new_new_n1129__), .dout(new_new_n1130__));
  and1  g0590(.dina(new_new_n1640__), .dinb(new_new_n1641__), .dout(new_new_n1131__));
  or1   g0591(.dina(new_new_n1643__), .dinb(new_new_n1645__), .dout(new_new_n1132__));
  and1  g0592(.dina(new_new_n1643__), .dinb(new_new_n1645__), .dout(new_new_n1133__));
  or1   g0593(.dina(new_new_n1640__), .dinb(new_new_n1641__), .dout(new_new_n1134__));
  and1  g0594(.dina(new_new_n1132__), .dinb(new_new_n1134__), .dout(new_new_n1135__));
  or1   g0595(.dina(new_new_n1131__), .dinb(new_new_n1133__), .dout(new_new_n1136__));
  or1   g0596(.dina(new_new_n1561__), .dinb(new_new_n1646__), .dout(new_new_n1137__));
  and1  g0597(.dina(new_new_n1648__), .dinb(new_new_n1649__), .dout(new_new_n1138__));
  and1  g0598(.dina(new_new_n1648__), .dinb(new_new_n1650__), .dout(new_new_n1139__));
  and1  g0599(.dina(new_new_n1647__), .dinb(new_new_n1651__), .dout(new_new_n1140__));
  and1  g0600(.dina(new_new_n1652__), .dinb(new_new_n1653__), .dout(new_new_n1141__));
  or1   g0601(.dina(new_new_n1652__), .dinb(new_new_n1653__), .dout(new_new_n1142__));
  or1   g0602(.dina(new_new_n1562__), .dinb(new_new_n1654__), .dout(new_new_n1143__));
  or1   g0603(.dina(new_new_n1656__), .dinb(new_new_n1657__), .dout(new_new_n1144__));
  and1  g0604(.dina(new_new_n1656__), .dinb(new_new_n1657__), .dout(new_new_n1145__));
  and1  g0605(.dina(new_new_n1658__), .dinb(new_new_n1572__), .dout(new_new_n1146__));
  or1   g0606(.dina(new_new_n548__), .dinb(new_new_n1574__), .dout(new_new_n1147__));
  and1  g0607(.dina(new_new_n1659__), .dinb(new_new_n1609__), .dout(new_new_n1148__));
  or1   g0608(.dina(new_new_n1661__), .dinb(new_new_n1602__), .dout(new_new_n1149__));
  and1  g0609(.dina(new_new_n1661__), .dinb(new_new_n1604__), .dout(new_new_n1150__));
  or1   g0610(.dina(new_new_n1659__), .dinb(new_new_n1609__), .dout(new_new_n1151__));
  and1  g0611(.dina(new_new_n1149__), .dinb(new_new_n1151__), .dout(new_new_n1152__));
  or1   g0612(.dina(new_new_n1148__), .dinb(new_new_n1150__), .dout(new_new_n1153__));
  and1  g0613(.dina(new_new_n1146__), .dinb(new_new_n1153__), .dout(new_new_n1154__));
  and1  g0614(.dina(new_new_n1147__), .dinb(new_new_n1152__), .dout(new_new_n1155__));
  or1   g0615(.dina(new_new_n1154__), .dinb(new_new_n1155__), .dout(new_new_n1156__));
  or1   g0616(.dina(new_new_n1595__), .dinb(new_new_n1639__), .dout(new_new_n1157__));
  or1   g0617(.dina(new_new_n1590__), .dinb(new_new_n1635__), .dout(new_new_n1158__));
  and1  g0618(.dina(new_new_n1157__), .dinb(new_new_n1158__), .dout(new_new_n1159__));
  and1  g0619(.dina(new_new_n1662__), .dinb(new_new_n1663__), .dout(new_new_n1160__));
  or1   g0620(.dina(new_new_n1662__), .dinb(new_new_n1663__), .dout(new_new_n1161__));
  and1  g0621(.dina(new_new_n1572__), .dinb(new_new_n1664__), .dout(new_new_n1162__));
  or1   g0622(.dina(new_new_n1576__), .dinb(new_new_n802__), .dout(new_new_n1163__));
  and1  g0623(.dina(new_new_n1666__), .dinb(new_new_n1667__), .dout(new_new_n1164__));
  or1   g0624(.dina(new_new_n1668__), .dinb(new_new_n1669__), .dout(new_new_n1165__));
  and1  g0625(.dina(new_new_n1668__), .dinb(new_new_n1669__), .dout(new_new_n1166__));
  or1   g0626(.dina(new_new_n1666__), .dinb(new_new_n1667__), .dout(new_new_n1167__));
  and1  g0627(.dina(new_new_n1165__), .dinb(new_new_n1167__), .dout(new_new_n1168__));
  or1   g0628(.dina(new_new_n1164__), .dinb(new_new_n1166__), .dout(new_new_n1169__));
  and1  g0629(.dina(new_new_n1670__), .dinb(new_new_n1671__), .dout(new_new_n1170__));
  or1   g0630(.dina(new_new_n1672__), .dinb(new_new_n1673__), .dout(new_new_n1171__));
  and1  g0631(.dina(new_new_n1672__), .dinb(new_new_n1673__), .dout(new_new_n1172__));
  or1   g0632(.dina(new_new_n1670__), .dinb(new_new_n1671__), .dout(new_new_n1173__));
  and1  g0633(.dina(new_new_n1171__), .dinb(new_new_n1173__), .dout(new_new_n1174__));
  or1   g0634(.dina(new_new_n1170__), .dinb(new_new_n1172__), .dout(new_new_n1175__));
  and1  g0635(.dina(new_new_n1083__), .dinb(new_new_n1174__), .dout(new_new_n1176__));
  and1  g0636(.dina(new_new_n1674__), .dinb(new_new_n1175__), .dout(new_new_n1177__));
  or1   g0637(.dina(new_new_n1176__), .dinb(new_new_n1177__), .dout(new_new_n1178__));
  and1  g0638(.dina(new_new_n1677__), .dinb(new_new_n1680__), .dout(new_new_n1179__));
  or1   g0639(.dina(new_new_n1682__), .dinb(new_new_n1685__), .dout(new_new_n1180__));
  and1  g0640(.dina(new_new_n1682__), .dinb(new_new_n1685__), .dout(new_new_n1181__));
  or1   g0641(.dina(new_new_n1677__), .dinb(new_new_n1680__), .dout(new_new_n1182__));
  and1  g0642(.dina(new_new_n1180__), .dinb(new_new_n1182__), .dout(new_new_n1183__));
  or1   g0643(.dina(new_new_n1179__), .dinb(new_new_n1181__), .dout(new_new_n1184__));
  and1  g0644(.dina(new_new_n1688__), .dinb(new_new_n1689__), .dout(new_new_n1185__));
  and1  g0645(.dina(new_new_n1690__), .dinb(new_new_n1691__), .dout(new_new_n1186__));
  or1   g0646(.dina(new_new_n1185__), .dinb(new_new_n1186__), .dout(new_new_n1187__));
  and1  g0647(.dina(new_new_n1692__), .dinb(new_new_n1693__), .dout(new_new_n1188__));
  and1  g0648(.dina(new_new_n1695__), .dinb(new_new_n1697__), .dout(new_new_n1189__));
  and1  g0649(.dina(new_new_n1698__), .dinb(new_new_n1700__), .dout(new_new_n1190__));
  and1  g0650(.dina(new_new_n1702__), .dinb(new_new_n552__), .dout(new_new_n1191__));
  and1  g0651(.dina(new_new_n1703__), .dinb(new_new_n1191__), .dout(new_new_n1192__));
  and1  g0652(.dina(new_new_n1704__), .dinb(new_new_n1693__), .dout(new_new_n1193__));
  or1   g0653(.dina(new_new_n858__), .dinb(new_new_n1705__), .dout(new_new_n1194__));
  and1  g0654(.dina(new_new_n1703__), .dinb(new_new_n1193__), .dout(new_new_n1195__));
  or1   g0655(.dina(new_new_n1706__), .dinb(new_new_n1194__), .dout(new_new_n1196__));
  and1  g0656(.dina(new_new_n1686__), .dinb(new_new_n1196__), .dout(new_new_n1197__));
  and1  g0657(.dina(new_new_n1679__), .dinb(new_new_n1195__), .dout(new_new_n1198__));
  or1   g0658(.dina(new_new_n1197__), .dinb(new_new_n1198__), .dout(new_new_n1199__));
  and1  g0659(.dina(new_new_n1708__), .dinb(new_new_n1709__), .dout(new_new_n1200__));
  or1   g0660(.dina(new_new_n1708__), .dinb(new_new_n1709__), .dout(new_new_n1201__));
  and1  g0661(.dina(new_new_n1711__), .dinb(new_new_n1689__), .dout(new_new_n1202__));
  and1  g0662(.dina(new_new_n1713__), .dinb(new_new_n1691__), .dout(new_new_n1203__));
  or1   g0663(.dina(new_new_n1202__), .dinb(new_new_n1203__), .dout(new_new_n1204__));
  and1  g0664(.dina(new_new_n1717__), .dinb(new_new_n1697__), .dout(new_new_n1205__));
  or1   g0665(.dina(new_new_n1720__), .dinb(new_new_n1700__), .dout(new_new_n1206__));
  and1  g0666(.dina(new_new_n1720__), .dinb(new_new_n1701__), .dout(new_new_n1207__));
  or1   g0667(.dina(new_new_n1717__), .dinb(new_new_n1696__), .dout(new_new_n1208__));
  and1  g0668(.dina(new_new_n1206__), .dinb(new_new_n1208__), .dout(new_new_n1209__));
  or1   g0669(.dina(new_new_n1205__), .dinb(new_new_n1207__), .dout(new_new_n1210__));
  and1  g0670(.dina(new_new_n1723__), .dinb(new_new_n1210__), .dout(new_new_n1211__));
  and1  g0671(.dina(new_new_n1725__), .dinb(new_new_n1209__), .dout(new_new_n1212__));
  or1   g0672(.dina(new_new_n1211__), .dinb(new_new_n1212__), .dout(new_new_n1213__));
  and1  g0673(.dina(new_new_n1688__), .dinb(new_new_n1136__), .dout(new_new_n1214__));
  and1  g0674(.dina(new_new_n1690__), .dinb(new_new_n1727__), .dout(new_new_n1215__));
  or1   g0675(.dina(new_new_n1214__), .dinb(new_new_n1215__), .dout(new_new_n1216__));
  and1  g0676(.dina(new_new_n1728__), .dinb(new_new_n1723__), .dout(new_new_n1217__));
  or1   g0677(.dina(new_new_n1730__), .dinb(new_new_n1725__), .dout(new_new_n1218__));
  and1  g0678(.dina(new_new_n1730__), .dinb(new_new_n1726__), .dout(new_new_n1219__));
  or1   g0679(.dina(new_new_n1728__), .dinb(new_new_n1722__), .dout(new_new_n1220__));
  and1  g0680(.dina(new_new_n1218__), .dinb(new_new_n1220__), .dout(new_new_n1221__));
  or1   g0681(.dina(new_new_n1217__), .dinb(new_new_n1219__), .dout(new_new_n1222__));
  and1  g0682(.dina(new_new_n1731__), .dinb(new_new_n1222__), .dout(new_new_n1223__));
  and1  g0683(.dina(new_new_n494__), .dinb(new_new_n1221__), .dout(new_new_n1224__));
  or1   g0684(.dina(new_new_n1223__), .dinb(new_new_n1224__), .dout(new_new_n1225__));
  and1  g0685(.dina(new_new_n1734__), .dinb(new_new_n1683__), .dout(new_new_n1226__));
  or1   g0686(.dina(new_new_n1737__), .dinb(new_new_n1676__), .dout(new_new_n1227__));
  and1  g0687(.dina(new_new_n1737__), .dinb(new_new_n1678__), .dout(new_new_n1228__));
  or1   g0688(.dina(new_new_n1734__), .dinb(new_new_n1683__), .dout(new_new_n1229__));
  and1  g0689(.dina(new_new_n1227__), .dinb(new_new_n1229__), .dout(new_new_n1230__));
  or1   g0690(.dina(new_new_n1226__), .dinb(new_new_n1228__), .dout(new_new_n1231__));
  and1  g0691(.dina(new_new_n502__), .dinb(new_new_n1231__), .dout(new_new_n1232__));
  and1  g0692(.dina(new_new_n1739__), .dinb(new_new_n1230__), .dout(new_new_n1233__));
  or1   g0693(.dina(new_new_n1232__), .dinb(new_new_n1233__), .dout(new_new_n1234__));
  and1  g0694(.dina(new_new_n1721__), .dinb(new_new_n1738__), .dout(new_new_n1235__));
  or1   g0695(.dina(new_new_n1716__), .dinb(new_new_n1733__), .dout(new_new_n1236__));
  and1  g0696(.dina(new_new_n1718__), .dinb(new_new_n1735__), .dout(new_new_n1237__));
  or1   g0697(.dina(new_new_n1721__), .dinb(new_new_n1738__), .dout(new_new_n1238__));
  and1  g0698(.dina(new_new_n1236__), .dinb(new_new_n1238__), .dout(new_new_n1239__));
  or1   g0699(.dina(new_new_n1235__), .dinb(new_new_n1237__), .dout(new_new_n1240__));
  and1  g0700(.dina(new_new_n1695__), .dinb(new_new_n1240__), .dout(new_new_n1241__));
  and1  g0701(.dina(new_new_n1698__), .dinb(new_new_n1239__), .dout(new_new_n1242__));
  or1   g0702(.dina(new_new_n1241__), .dinb(new_new_n1242__), .dout(new_new_n1243__));
  and1  g0703(.dina(new_new_n1711__), .dinb(new_new_n1740__), .dout(new_new_n1244__));
  or1   g0704(.dina(new_new_n1713__), .dinb(new_new_n1742__), .dout(new_new_n1245__));
  and1  g0705(.dina(new_new_n1714__), .dinb(new_new_n1742__), .dout(new_new_n1246__));
  or1   g0706(.dina(new_new_n1710__), .dinb(new_new_n1740__), .dout(new_new_n1247__));
  and1  g0707(.dina(new_new_n1245__), .dinb(new_new_n1247__), .dout(new_new_n1248__));
  or1   g0708(.dina(new_new_n1244__), .dinb(new_new_n1246__), .dout(new_new_n1249__));
  and1  g0709(.dina(new_new_n1743__), .dinb(new_new_n1249__), .dout(new_new_n1250__));
  and1  g0710(.dina(new_new_n1707__), .dinb(new_new_n1248__), .dout(new_new_n1251__));
  or1   g0711(.dina(new_new_n1250__), .dinb(new_new_n1251__), .dout(new_new_n1252__));
  and1  g0712(.dina(new_new_n1745__), .dinb(new_new_n1746__), .dout(new_new_n1253__));
  or1   g0713(.dina(new_new_n1745__), .dinb(new_new_n1746__), .dout(new_new_n1254__));
  buf1  g0714(.din(new_new_n865__), .dout(G1884));
  buf1  g0715(.din(new_new_n868__), .dout(G1885));
  buf1  g0716(.din(new_new_n871__), .dout(G1886));
  buf1  g0717(.din(new_new_n874__), .dout(G1887));
  buf1  g0718(.din(new_new_n879__), .dout(G1888));
  buf1  g0719(.din(new_new_n882__), .dout(G1889));
  buf1  g0720(.din(new_new_n885__), .dout(G1890));
  buf1  g0721(.din(new_new_n894__), .dout(G1891));
  buf1  g0722(.din(new_new_n897__), .dout(G1892));
  buf1  g0723(.din(new_new_n900__), .dout(G1893));
  buf1  g0724(.din(new_new_n903__), .dout(G1894));
  buf1  g0725(.din(new_new_n908__), .dout(G1895));
  buf1  g0726(.din(new_new_n919__), .dout(G1896));
  buf1  g0727(.din(new_new_n922__), .dout(G1897));
  buf1  g0728(.din(new_new_n925__), .dout(G1898));
  buf1  g0729(.din(new_new_n928__), .dout(G1899));
  buf1  g0730(.din(new_new_n937__), .dout(G1900));
  buf1  g0731(.din(new_new_n945__), .dout(G1901));
  buf1  g0732(.din(new_new_n953__), .dout(G1902));
  buf1  g0733(.din(new_new_n957__), .dout(G1903));
  buf1  g0734(.din(new_new_n961__), .dout(G1904));
  buf1  g0735(.din(new_new_n965__), .dout(G1905));
  buf1  g0736(.din(new_new_n980__), .dout(G1906));
  buf1  g0737(.din(new_new_n997__), .dout(G1907));
  buf1  g0738(.din(new_new_n1001__), .dout(G1908));
  buf1  g0739(.din(new_new_n427__), .dout(n2688));
  buf1  g0740(.din(new_new_n661__), .dout(n2691));
  buf1  g0741(.din(new_new_n641__), .dout(n2694));
  buf1  g0742(.din(new_new_n643__), .dout(n2697));
  buf1  g0743(.din(new_new_n433__), .dout(n2700));
  buf1  g0744(.din(new_new_n663__), .dout(n2703));
  buf1  g0745(.din(new_new_n435__), .dout(n2706));
  buf1  g0746(.din(new_new_n665__), .dout(n2709));
  buf1  g0747(.din(new_new_n645__), .dout(n2712));
  buf1  g0748(.din(new_new_n647__), .dout(n2715));
  buf1  g0749(.din(new_new_n649__), .dout(n2718));
  buf1  g0750(.din(new_new_n651__), .dout(n2721));
  buf1  g0751(.din(new_new_n625__), .dout(n2724));
  buf1  g0752(.din(new_new_n447__), .dout(n2727));
  buf1  g0753(.din(new_new_n657__), .dout(n2730));
  buf1  g0754(.din(new_new_n627__), .dout(n2733));
  buf1  g0755(.din(new_new_n629__), .dout(n2736));
  buf1  g0756(.din(new_new_n653__), .dout(n2739));
  buf1  g0757(.din(new_new_n631__), .dout(n2742));
  buf1  g0758(.din(new_new_n457__), .dout(n2745));
  buf1  g0759(.din(new_new_n659__), .dout(n2748));
  buf1  g0760(.din(new_new_n459__), .dout(n2751));
  buf1  g0761(.din(new_new_n463__), .dout(n2754));
  buf1  g0762(.din(new_new_n465__), .dout(n2757));
  buf1  g0763(.din(new_new_n467__), .dout(n2760));
  buf1  g0764(.din(new_new_n681__), .dout(n2763));
  buf1  g0765(.din(new_new_n469__), .dout(n2766));
  buf1  g0766(.din(new_new_n545__), .dout(n2769));
  buf1  g0767(.din(new_new_n695__), .dout(n2772));
  buf1  g0768(.din(new_new_n471__), .dout(n2775));
  buf1  g0769(.din(new_new_n475__), .dout(n2778));
  buf1  g0770(.din(new_new_n553__), .dout(n2781));
  buf1  g0771(.din(new_new_n555__), .dout(n2784));
  buf1  g0772(.din(new_new_n1552__), .dout(n2787));
  buf1  g0773(.din(new_new_n477__), .dout(n2790));
  buf1  g0774(.din(new_new_n561__), .dout(n2793));
  buf1  g0775(.din(new_new_n1554__), .dout(n2796));
  buf1  g0776(.din(new_new_n479__), .dout(n2799));
  buf1  g0777(.din(new_new_n567__), .dout(n2802));
  buf1  g0778(.din(new_new_n1553__), .dout(n2805));
  buf1  g0779(.din(new_new_n481__), .dout(n2808));
  buf1  g0780(.din(new_new_n573__), .dout(n2811));
  buf1  g0781(.din(new_new_n743__), .dout(n2814));
  buf1  g0782(.din(new_new_n483__), .dout(n2817));
  buf1  g0783(.din(new_new_n579__), .dout(n2820));
  buf1  g0784(.din(new_new_n581__), .dout(n2823));
  buf1  g0785(.din(new_new_n1545__), .dout(n2826));
  buf1  g0786(.din(new_new_n485__), .dout(n2829));
  buf1  g0787(.din(new_new_n587__), .dout(n2832));
  buf1  g0788(.din(new_new_n589__), .dout(n2835));
  buf1  g0789(.din(new_new_n1549__), .dout(n2838));
  buf1  g0790(.din(new_new_n487__), .dout(n2841));
  buf1  g0791(.din(new_new_n595__), .dout(n2844));
  buf1  g0792(.din(new_new_n1542__), .dout(n2847));
  buf1  g0793(.din(new_new_n489__), .dout(n2850));
  buf1  g0794(.din(new_new_n601__), .dout(n2853));
  buf1  g0795(.din(new_new_n603__), .dout(n2856));
  buf1  g0796(.din(new_new_n1550__), .dout(n2859));
  buf1  g0797(.din(new_new_n1548__), .dout(n2862));
  buf1  g0798(.din(new_new_n733__), .dout(n2865));
  buf1  g0799(.din(new_new_n737__), .dout(n2868));
  buf1  g0800(.din(new_new_n735__), .dout(n2871));
  buf1  g0801(.din(new_new_n749__), .dout(n2874));
  buf1  g0802(.din(new_new_n759__), .dout(n2877));
  buf1  g0803(.din(new_new_n757__), .dout(n2880));
  buf1  g0804(.din(new_new_n1543__), .dout(n2883));
  buf1  g0805(.din(new_new_n703__), .dout(n2886));
  buf1  g0806(.din(new_new_n705__), .dout(n2889));
  buf1  g0807(.din(new_new_n1587__), .dout(n2892));
  buf1  g0808(.din(new_new_n709__), .dout(n2895));
  buf1  g0809(.din(new_new_n1544__), .dout(n2898));
  buf1  g0810(.din(new_new_n711__), .dout(n2901));
  buf1  g0811(.din(new_new_n1646__), .dout(n2904));
  buf1  g0812(.din(new_new_n1551__), .dout(n2907));
  buf1  g0813(.din(new_new_n1627__), .dout(n2910));
  buf1  g0814(.din(new_new_n719__), .dout(n2913));
  buf1  g0815(.din(new_new_n721__), .dout(n2916));
  buf1  g0816(.din(new_new_n723__), .dout(n2919));
  buf1  g0817(.din(new_new_n1605__), .dout(n2922));
  buf1  g0818(.din(new_new_n1665__), .dout(n2925));
  buf1  g0819(.din(new_new_n1660__), .dout(n2928));
  buf1  g0820(.din(new_new_n1576__), .dout(n2931));
  buf1  g0821(.din(new_new_n739__), .dout(n2934));
  buf1  g0822(.din(new_new_n741__), .dout(n2937));
  buf1  g0823(.din(new_new_n1630__), .dout(n2940));
  buf1  g0824(.din(new_new_n1604__), .dout(n2943));
  buf1  g0825(.din(new_new_n765__), .dout(n2946));
  buf1  g0826(.din(new_new_n767__), .dout(n2949));
  buf1  g0827(.din(new_new_n1563__), .dout(n2952));
  buf1  g0828(.din(new_new_n771__), .dout(n2955));
  buf1  g0829(.din(new_new_n783__), .dout(n2958));
  not1  g0830(.din(new_new_n1557__), .dout(n2961));
  buf1  g0831(.din(new_new_n1558__), .dout(n2964));
  not1  g0832(.din(new_new_n1555__), .dout(n2967));
  buf1  g0833(.din(new_new_n1664__), .dout(n2970));
  buf1  g0834(.din(new_new_n1616__), .dout(n2973));
  buf1  g0835(.din(new_new_n1620__), .dout(n2976));
  buf1  g0836(.din(new_new_n1618__), .dout(n2979));
  not1  g0837(.din(new_new_n1556__), .dout(n2982));
  buf1  g0838(.din(new_new_n1559__), .dout(n2985));
  buf1  g0839(.din(new_new_n1639__), .dout(n2988));
  buf1  g0840(.din(new_new_n1658__), .dout(n2991));
  buf1  g0841(.din(new_new_n1562__), .dout(n2994));
  not1  g0842(.din(new_new_n1621__), .dout(n2997));
  buf1  g0843(.din(new_new_n1622__), .dout(n3000));
  buf1  g0844(.din(new_new_n1678__), .dout(n3003));
  buf1  g0845(.din(new_new_n1714__), .dout(n3006));
  buf1  g0846(.din(new_new_n1741__), .dout(n3009));
  buf1  g0847(.din(new_new_n1686__), .dout(n3012));
  buf1  g0848(.din(new_new_n1704__), .dout(n3015));
  buf1  g0849(.din(new_new_n1705__), .dout(n3018));
  buf1  g0850(.din(new_new_n1614__), .dout(n3021));
  buf1  g0851(.din(new_new_n1729__), .dout(n3024));
  buf1  g0852(.din(new_new_n1726__), .dout(n3027));
  buf1  g0853(.din(new_new_n1718__), .dout(n3030));
  buf1  g0854(.din(new_new_n1735__), .dout(n3033));
  buf1  g0855(.din(new_new_n1701__), .dout(n3036));
  buf1  g0856(.din(new_new_n1642__), .dout(n3039));
  buf1  g0857(.din(new_new_n1644__), .dout(n3042));
  buf1  g0858(.din(new_new_n1706__), .dout(n3045));
  buf1  g0859(.din(new_new_n1651__), .dout(n3048));
  buf1  g0860(.din(new_new_n1654__), .dout(n3051));
  buf1  g0861(.din(new_new_n1674__), .dout(n3054));
  buf1  g0862(.din(new_new_n1743__), .dout(n3057));
  buf1  g0863(.din(new_new_n1687__), .dout(n3060));
  buf1  g0864(.din(new_new_n575__), .dout(n3063));
  buf1  g0865(.din(new_new_n1084__), .dout(n3066));
  buf1  g0866(.din(new_new_n1085__), .dout(n3069));
  buf1  g0867(.din(new_new_n1655__), .dout(n3072));
  buf1  g0868(.din(new_new_n1091__), .dout(n3075));
  buf1  g0869(.din(new_new_n1093__), .dout(n3078));
  buf1  g0870(.din(new_new_n1094__), .dout(n3081));
  buf1  g0871(.din(new_new_n1649__), .dout(n3084));
  not1  g0872(.din(new_new_n1650__), .dout(n3087));
  buf1  g0873(.din(new_new_n1731__), .dout(n3090));
  buf1  g0874(.din(new_new_n1739__), .dout(n3093));
  buf1  g0875(.din(new_new_n1694__), .dout(n3096));
  buf1  g0876(.din(new_new_n1702__), .dout(n3099));
  buf1  g0877(.din(new_new_n551__), .dout(n3102));
  buf1  g0878(.din(new_new_n1727__), .dout(n3105));
  buf1  g0879(.din(new_new_n563__), .dout(n3108));
  buf1  g0880(.din(new_new_n569__), .dout(n3111));
  buf1  g0881(.din(new_new_n1137__), .dout(n3114));
  buf1  g0882(.din(new_new_n1138__), .dout(n3117));
  not1  g0883(.din(new_new_n1139__), .dout(n3120));
  buf1  g0884(.din(new_new_n1692__), .dout(n3123));
  buf1  g0885(.din(new_new_n1141__), .dout(n3126));
  not1  g0886(.din(new_new_n1142__), .dout(n3129));
  buf1  g0887(.din(new_new_n1144__), .dout(n3132));
  buf1  g0888(.din(new_new_n1145__), .dout(n3135));
  buf1  g0889(.din(new_new_n1160__), .dout(n3138));
  not1  g0890(.din(new_new_n1161__), .dout(n3141));
  buf1  g0891(.din(new_new_n1178__), .dout(n3144));
  not1  g0892(.din(new_new_n1744__), .dout(n3147));
  buf1  g0893(.din(new_new_n541__), .dout(n3150));
  buf1  g0894(.din(new_new_n1188__), .dout(n3153));
  buf1  g0895(.din(new_new_n1189__), .dout(n3156));
  buf1  g0896(.din(new_new_n1190__), .dout(n3159));
  buf1  g0897(.din(new_new_n1192__), .dout(n3162));
  buf1  g0898(.din(new_new_n1200__), .dout(n3165));
  not1  g0899(.din(new_new_n1201__), .dout(n3168));
  buf1  g0900(.din(new_new_n537__), .dout(n3171));
  buf1  g0901(.din(new_new_n1204__), .dout(n3174));
  buf1  g0902(.din(new_new_n1213__), .dout(n3177));
  buf1  g0903(.din(new_new_n1216__), .dout(n3180));
  buf1  g0904(.din(new_new_n1225__), .dout(n3183));
  buf1  g0905(.din(new_new_n1234__), .dout(n3186));
  buf1  g0906(.din(new_new_n1243__), .dout(n3189));
  buf1  g0907(.din(new_new_n1253__), .dout(n3192));
  not1  g0908(.din(new_new_n1254__), .dout(n3195));
  buf1  g0909(.din(new_new_n429__), .dout(n3198));
  buf1  g0910(.din(new_new_n431__), .dout(n3201));
  buf1  g0911(.din(new_new_n437__), .dout(n3204));
  buf1  g0912(.din(new_new_n439__), .dout(n3207));
  buf1  g0913(.din(new_new_n441__), .dout(n3210));
  buf1  g0914(.din(new_new_n443__), .dout(n3213));
  buf1  g0915(.din(new_new_n453__), .dout(n3216));
  buf1  g0916(.din(new_new_n491__), .dout(n3219));
  buf1  g0917(.din(new_new_n445__), .dout(n3222));
  buf1  g0918(.din(new_new_n449__), .dout(n3225));
  buf1  g0919(.din(new_new_n451__), .dout(n3228));
  buf1  g0920(.din(new_new_n455__), .dout(n3231));
  buf1  g0921(.din(new_new_n461__), .dout(n3234));
  buf1  g0922(.din(new_new_n473__), .dout(n3237));
  buf1  g0923(.din(new_new_n752__), .dout(new_new_n1464__));
  buf1  g0924(.din(new_new_n755__), .dout(new_new_n1465__));
  buf1  g0925(.din(new_new_n751__), .dout(new_new_n1466__));
  buf1  g0926(.din(new_new_n756__), .dout(new_new_n1467__));
  buf1  g0927(.din(new_new_n862__), .dout(new_new_n1468__));
  buf1  g0928(.din(new_new_n1468__), .dout(new_new_n1469__));
  buf1  g0929(.din(new_new_n1469__), .dout(new_new_n1470__));
  buf1  g0930(.din(new_new_n1469__), .dout(new_new_n1471__));
  buf1  g0931(.din(new_new_n1468__), .dout(new_new_n1472__));
  buf1  g0932(.din(new_new_n1472__), .dout(new_new_n1473__));
  buf1  g0933(.din(new_new_n861__), .dout(new_new_n1474__));
  buf1  g0934(.din(new_new_n1474__), .dout(new_new_n1475__));
  buf1  g0935(.din(new_new_n1475__), .dout(new_new_n1476__));
  buf1  g0936(.din(new_new_n1475__), .dout(new_new_n1477__));
  buf1  g0937(.din(new_new_n1474__), .dout(new_new_n1478__));
  buf1  g0938(.din(new_new_n1478__), .dout(new_new_n1479__));
  buf1  g0939(.din(new_new_n754__), .dout(new_new_n1480__));
  buf1  g0940(.din(new_new_n1480__), .dout(new_new_n1481__));
  buf1  g0941(.din(new_new_n753__), .dout(new_new_n1482__));
  buf1  g0942(.din(new_new_n1482__), .dout(new_new_n1483__));
  buf1  g0943(.din(new_new_n876__), .dout(new_new_n1484__));
  buf1  g0944(.din(new_new_n1484__), .dout(new_new_n1485__));
  buf1  g0945(.din(new_new_n1485__), .dout(new_new_n1486__));
  buf1  g0946(.din(new_new_n1485__), .dout(new_new_n1487__));
  buf1  g0947(.din(new_new_n1484__), .dout(new_new_n1488__));
  buf1  g0948(.din(new_new_n875__), .dout(new_new_n1489__));
  buf1  g0949(.din(new_new_n1489__), .dout(new_new_n1490__));
  buf1  g0950(.din(new_new_n1490__), .dout(new_new_n1491__));
  buf1  g0951(.din(new_new_n1490__), .dout(new_new_n1492__));
  buf1  g0952(.din(new_new_n1489__), .dout(new_new_n1493__));
  buf1  g0953(.din(new_new_n690__), .dout(new_new_n1494__));
  buf1  g0954(.din(new_new_n680__), .dout(new_new_n1495__));
  buf1  g0955(.din(new_new_n888__), .dout(new_new_n1496__));
  buf1  g0956(.din(new_new_n889__), .dout(new_new_n1497__));
  buf1  g0957(.din(new_new_n891__), .dout(new_new_n1498__));
  buf1  g0958(.din(new_new_n1498__), .dout(new_new_n1499__));
  buf1  g0959(.din(new_new_n1498__), .dout(new_new_n1500__));
  buf1  g0960(.din(new_new_n890__), .dout(new_new_n1501__));
  buf1  g0961(.din(new_new_n1501__), .dout(new_new_n1502__));
  buf1  g0962(.din(new_new_n1501__), .dout(new_new_n1503__));
  buf1  g0963(.din(new_new_n676__), .dout(new_new_n1504__));
  buf1  g0964(.din(new_new_n677__), .dout(new_new_n1505__));
  buf1  g0965(.din(new_new_n691__), .dout(new_new_n1506__));
  buf1  g0966(.din(new_new_n916__), .dout(new_new_n1507__));
  buf1  g0967(.din(new_new_n1507__), .dout(new_new_n1508__));
  buf1  g0968(.din(new_new_n1507__), .dout(new_new_n1509__));
  buf1  g0969(.din(new_new_n915__), .dout(new_new_n1510__));
  buf1  g0970(.din(new_new_n1510__), .dout(new_new_n1511__));
  buf1  g0971(.din(new_new_n1510__), .dout(new_new_n1512__));
  buf1  g0972(.din(new_new_n930__), .dout(new_new_n1513__));
  buf1  g0973(.din(new_new_n1513__), .dout(new_new_n1514__));
  buf1  g0974(.din(new_new_n1514__), .dout(new_new_n1515__));
  buf1  g0975(.din(new_new_n1514__), .dout(new_new_n1516__));
  buf1  g0976(.din(new_new_n1513__), .dout(new_new_n1517__));
  buf1  g0977(.din(new_new_n609__), .dout(new_new_n1518__));
  buf1  g0978(.din(new_new_n1518__), .dout(new_new_n1519__));
  buf1  g0979(.din(new_new_n600__), .dout(new_new_n1520__));
  buf1  g0980(.din(new_new_n1520__), .dout(new_new_n1521__));
  buf1  g0981(.din(new_new_n1521__), .dout(new_new_n1522__));
  buf1  g0982(.din(new_new_n1520__), .dout(new_new_n1523__));
  buf1  g0983(.din(new_new_n599__), .dout(new_new_n1524__));
  buf1  g0984(.din(new_new_n1524__), .dout(new_new_n1525__));
  buf1  g0985(.din(new_new_n929__), .dout(new_new_n1526__));
  buf1  g0986(.din(new_new_n1526__), .dout(new_new_n1527__));
  buf1  g0987(.din(new_new_n687__), .dout(new_new_n1528__));
  buf1  g0988(.din(new_new_n1528__), .dout(new_new_n1529__));
  buf1  g0989(.din(new_new_n1529__), .dout(new_new_n1530__));
  buf1  g0990(.din(new_new_n1529__), .dout(new_new_n1531__));
  buf1  g0991(.din(new_new_n1528__), .dout(new_new_n1532__));
  buf1  g0992(.din(new_new_n610__), .dout(new_new_n1533__));
  buf1  g0993(.din(new_new_n971__), .dout(new_new_n1534__));
  buf1  g0994(.din(new_new_n970__), .dout(new_new_n1535__));
  buf1  g0995(.din(new_new_n988__), .dout(new_new_n1536__));
  buf1  g0996(.din(new_new_n987__), .dout(new_new_n1537__));
  buf1  g0997(.din(new_new_n778__), .dout(new_new_n1538__));
  buf1  g0998(.din(new_new_n698__), .dout(new_new_n1539__));
  buf1  g0999(.din(new_new_n697__), .dout(new_new_n1540__));
  buf1  g1000(.din(new_new_n1540__), .dout(new_new_n1541__));
  buf1  g1001(.din(new_new_n1540__), .dout(new_new_n1542__));
  buf1  g1002(.din(new_new_n797__), .dout(new_new_n1543__));
  buf1  g1003(.din(new_new_n1002__), .dout(new_new_n1544__));
  buf1  g1004(.din(new_new_n583__), .dout(new_new_n1545__));
  buf1  g1005(.din(new_new_n655__), .dout(new_new_n1546__));
  buf1  g1006(.din(new_new_n1546__), .dout(new_new_n1547__));
  buf1  g1007(.din(new_new_n1546__), .dout(new_new_n1548__));
  buf1  g1008(.din(new_new_n591__), .dout(new_new_n1549__));
  buf1  g1009(.din(new_new_n605__), .dout(new_new_n1550__));
  buf1  g1010(.din(new_new_n1005__), .dout(new_new_n1551__));
  buf1  g1011(.din(new_new_n557__), .dout(new_new_n1552__));
  buf1  g1012(.din(new_new_n775__), .dout(new_new_n1553__));
  buf1  g1013(.din(new_new_n773__), .dout(new_new_n1554__));
  buf1  g1014(.din(new_new_n1012__), .dout(new_new_n1555__));
  buf1  g1015(.din(new_new_n1020__), .dout(new_new_n1556__));
  buf1  g1016(.din(new_new_n1006__), .dout(new_new_n1557__));
  buf1  g1017(.din(new_new_n1011__), .dout(new_new_n1558__));
  buf1  g1018(.din(new_new_n1031__), .dout(new_new_n1559__));
  buf1  g1019(.din(new_new_n597__), .dout(new_new_n1560__));
  buf1  g1020(.din(new_new_n1560__), .dout(new_new_n1561__));
  buf1  g1021(.din(new_new_n1560__), .dout(new_new_n1562__));
  buf1  g1022(.din(new_new_n769__), .dout(new_new_n1563__));
  buf1  g1023(.din(new_new_n1563__), .dout(new_new_n1564__));
  buf1  g1024(.din(new_new_n818__), .dout(new_new_n1565__));
  buf1  g1025(.din(new_new_n819__), .dout(new_new_n1566__));
  buf1  g1026(.din(new_new_n817__), .dout(new_new_n1567__));
  buf1  g1027(.din(new_new_n820__), .dout(new_new_n1568__));
  buf1  g1028(.din(new_new_n815__), .dout(new_new_n1569__));
  buf1  g1029(.din(new_new_n732__), .dout(new_new_n1570__));
  buf1  g1030(.din(new_new_n1570__), .dout(new_new_n1571__));
  buf1  g1031(.din(new_new_n1570__), .dout(new_new_n1572__));
  buf1  g1032(.din(new_new_n731__), .dout(new_new_n1573__));
  buf1  g1033(.din(new_new_n1573__), .dout(new_new_n1574__));
  buf1  g1034(.din(new_new_n1574__), .dout(new_new_n1575__));
  buf1  g1035(.din(new_new_n1573__), .dout(new_new_n1576__));
  buf1  g1036(.din(new_new_n822__), .dout(new_new_n1577__));
  buf1  g1037(.din(new_new_n1577__), .dout(new_new_n1578__));
  buf1  g1038(.din(new_new_n1577__), .dout(new_new_n1579__));
  buf1  g1039(.din(new_new_n825__), .dout(new_new_n1580__));
  buf1  g1040(.din(new_new_n821__), .dout(new_new_n1581__));
  buf1  g1041(.din(new_new_n1581__), .dout(new_new_n1582__));
  buf1  g1042(.din(new_new_n1581__), .dout(new_new_n1583__));
  buf1  g1043(.din(new_new_n826__), .dout(new_new_n1584__));
  buf1  g1044(.din(new_new_n708__), .dout(new_new_n1585__));
  buf1  g1045(.din(new_new_n809__), .dout(new_new_n1586__));
  buf1  g1046(.din(new_new_n707__), .dout(new_new_n1587__));
  buf1  g1047(.din(new_new_n1587__), .dout(new_new_n1588__));
  buf1  g1048(.din(new_new_n810__), .dout(new_new_n1589__));
  buf1  g1049(.din(new_new_n823__), .dout(new_new_n1590__));
  buf1  g1050(.din(new_new_n1590__), .dout(new_new_n1591__));
  buf1  g1051(.din(new_new_n827__), .dout(new_new_n1592__));
  buf1  g1052(.din(new_new_n1592__), .dout(new_new_n1593__));
  buf1  g1053(.din(new_new_n1592__), .dout(new_new_n1594__));
  buf1  g1054(.din(new_new_n824__), .dout(new_new_n1595__));
  buf1  g1055(.din(new_new_n1595__), .dout(new_new_n1596__));
  buf1  g1056(.din(new_new_n828__), .dout(new_new_n1597__));
  buf1  g1057(.din(new_new_n1597__), .dout(new_new_n1598__));
  buf1  g1058(.din(new_new_n1597__), .dout(new_new_n1599__));
  buf1  g1059(.din(new_new_n726__), .dout(new_new_n1600__));
  buf1  g1060(.din(new_new_n763__), .dout(new_new_n1601__));
  buf1  g1061(.din(new_new_n1601__), .dout(new_new_n1602__));
  buf1  g1062(.din(new_new_n1602__), .dout(new_new_n1603__));
  buf1  g1063(.din(new_new_n1601__), .dout(new_new_n1604__));
  buf1  g1064(.din(new_new_n725__), .dout(new_new_n1605__));
  buf1  g1065(.din(new_new_n1605__), .dout(new_new_n1606__));
  buf1  g1066(.din(new_new_n764__), .dout(new_new_n1607__));
  buf1  g1067(.din(new_new_n1607__), .dout(new_new_n1608__));
  buf1  g1068(.din(new_new_n1607__), .dout(new_new_n1609__));
  buf1  g1069(.din(new_new_n1071__), .dout(new_new_n1610__));
  buf1  g1070(.din(new_new_n1076__), .dout(new_new_n1611__));
  buf1  g1071(.din(new_new_n1070__), .dout(new_new_n1612__));
  buf1  g1072(.din(new_new_n1077__), .dout(new_new_n1613__));
  buf1  g1073(.din(new_new_n1037__), .dout(new_new_n1614__));
  buf1  g1074(.din(new_new_n1087__), .dout(new_new_n1615__));
  buf1  g1075(.din(new_new_n1013__), .dout(new_new_n1616__));
  buf1  g1076(.din(new_new_n1088__), .dout(new_new_n1617__));
  buf1  g1077(.din(new_new_n1015__), .dout(new_new_n1618__));
  buf1  g1078(.din(new_new_n1090__), .dout(new_new_n1619__));
  buf1  g1079(.din(new_new_n1014__), .dout(new_new_n1620__));
  buf1  g1080(.din(new_new_n1034__), .dout(new_new_n1621__));
  buf1  g1081(.din(new_new_n1036__), .dout(new_new_n1622__));
  buf1  g1082(.din(new_new_n1095__), .dout(new_new_n1623__));
  buf1  g1083(.din(new_new_n1096__), .dout(new_new_n1624__));
  buf1  g1084(.din(new_new_n718__), .dout(new_new_n1625__));
  buf1  g1085(.din(new_new_n1104__), .dout(new_new_n1626__));
  buf1  g1086(.din(new_new_n717__), .dout(new_new_n1627__));
  buf1  g1087(.din(new_new_n1627__), .dout(new_new_n1628__));
  buf1  g1088(.din(new_new_n1103__), .dout(new_new_n1629__));
  buf1  g1089(.din(new_new_n761__), .dout(new_new_n1630__));
  buf1  g1090(.din(new_new_n1630__), .dout(new_new_n1631__));
  buf1  g1091(.din(new_new_n1114__), .dout(new_new_n1632__));
  buf1  g1092(.din(new_new_n762__), .dout(new_new_n1633__));
  buf1  g1093(.din(new_new_n1115__), .dout(new_new_n1634__));
  buf1  g1094(.din(new_new_n1032__), .dout(new_new_n1635__));
  buf1  g1095(.din(new_new_n1635__), .dout(new_new_n1636__));
  buf1  g1096(.din(new_new_n1033__), .dout(new_new_n1637__));
  buf1  g1097(.din(new_new_n1637__), .dout(new_new_n1638__));
  buf1  g1098(.din(new_new_n1637__), .dout(new_new_n1639__));
  buf1  g1099(.din(new_new_n844__), .dout(new_new_n1640__));
  buf1  g1100(.din(new_new_n846__), .dout(new_new_n1641__));
  buf1  g1101(.din(new_new_n843__), .dout(new_new_n1642__));
  buf1  g1102(.din(new_new_n1642__), .dout(new_new_n1643__));
  buf1  g1103(.din(new_new_n845__), .dout(new_new_n1644__));
  buf1  g1104(.din(new_new_n1644__), .dout(new_new_n1645__));
  buf1  g1105(.din(new_new_n713__), .dout(new_new_n1646__));
  buf1  g1106(.din(new_new_n598__), .dout(new_new_n1647__));
  buf1  g1107(.din(new_new_n1647__), .dout(new_new_n1648__));
  buf1  g1108(.din(new_new_n1113__), .dout(new_new_n1649__));
  buf1  g1109(.din(new_new_n1130__), .dout(new_new_n1650__));
  buf1  g1110(.din(new_new_n1050__), .dout(new_new_n1651__));
  buf1  g1111(.din(new_new_n576__), .dout(new_new_n1652__));
  buf1  g1112(.din(new_new_n1140__), .dout(new_new_n1653__));
  buf1  g1113(.din(new_new_n1065__), .dout(new_new_n1654__));
  buf1  g1114(.din(new_new_n1086__), .dout(new_new_n1655__));
  buf1  g1115(.din(new_new_n1655__), .dout(new_new_n1656__));
  buf1  g1116(.din(new_new_n1143__), .dout(new_new_n1657__));
  buf1  g1117(.din(new_new_n547__), .dout(new_new_n1658__));
  buf1  g1118(.din(new_new_n730__), .dout(new_new_n1659__));
  buf1  g1119(.din(new_new_n729__), .dout(new_new_n1660__));
  buf1  g1120(.din(new_new_n1660__), .dout(new_new_n1661__));
  buf1  g1121(.din(new_new_n1156__), .dout(new_new_n1662__));
  buf1  g1122(.din(new_new_n1159__), .dout(new_new_n1663__));
  buf1  g1123(.din(new_new_n801__), .dout(new_new_n1664__));
  buf1  g1124(.din(new_new_n727__), .dout(new_new_n1665__));
  buf1  g1125(.din(new_new_n1665__), .dout(new_new_n1666__));
  buf1  g1126(.din(new_new_n800__), .dout(new_new_n1667__));
  buf1  g1127(.din(new_new_n728__), .dout(new_new_n1668__));
  buf1  g1128(.din(new_new_n799__), .dout(new_new_n1669__));
  buf1  g1129(.din(new_new_n1162__), .dout(new_new_n1670__));
  buf1  g1130(.din(new_new_n1169__), .dout(new_new_n1671__));
  buf1  g1131(.din(new_new_n1163__), .dout(new_new_n1672__));
  buf1  g1132(.din(new_new_n1168__), .dout(new_new_n1673__));
  buf1  g1133(.din(new_new_n1082__), .dout(new_new_n1674__));
  buf1  g1134(.din(new_new_n849__), .dout(new_new_n1675__));
  buf1  g1135(.din(new_new_n1675__), .dout(new_new_n1676__));
  buf1  g1136(.din(new_new_n1676__), .dout(new_new_n1677__));
  buf1  g1137(.din(new_new_n1675__), .dout(new_new_n1678__));
  buf1  g1138(.din(new_new_n856__), .dout(new_new_n1679__));
  buf1  g1139(.din(new_new_n1679__), .dout(new_new_n1680__));
  buf1  g1140(.din(new_new_n850__), .dout(new_new_n1681__));
  buf1  g1141(.din(new_new_n1681__), .dout(new_new_n1682__));
  buf1  g1142(.din(new_new_n1681__), .dout(new_new_n1683__));
  buf1  g1143(.din(new_new_n855__), .dout(new_new_n1684__));
  buf1  g1144(.din(new_new_n1684__), .dout(new_new_n1685__));
  buf1  g1145(.din(new_new_n1684__), .dout(new_new_n1686__));
  buf1  g1146(.din(new_new_n531__), .dout(new_new_n1687__));
  buf1  g1147(.din(new_new_n1687__), .dout(new_new_n1688__));
  buf1  g1148(.din(new_new_n1184__), .dout(new_new_n1689__));
  buf1  g1149(.din(new_new_n532__), .dout(new_new_n1690__));
  buf1  g1150(.din(new_new_n1183__), .dout(new_new_n1691__));
  buf1  g1151(.din(new_new_n535__), .dout(new_new_n1692__));
  buf1  g1152(.din(new_new_n860__), .dout(new_new_n1693__));
  buf1  g1153(.din(new_new_n505__), .dout(new_new_n1694__));
  buf1  g1154(.din(new_new_n1694__), .dout(new_new_n1695__));
  buf1  g1155(.din(new_new_n842__), .dout(new_new_n1696__));
  buf1  g1156(.din(new_new_n1696__), .dout(new_new_n1697__));
  buf1  g1157(.din(new_new_n506__), .dout(new_new_n1698__));
  buf1  g1158(.din(new_new_n841__), .dout(new_new_n1699__));
  buf1  g1159(.din(new_new_n1699__), .dout(new_new_n1700__));
  buf1  g1160(.din(new_new_n1699__), .dout(new_new_n1701__));
  buf1  g1161(.din(new_new_n539__), .dout(new_new_n1702__));
  buf1  g1162(.din(new_new_n848__), .dout(new_new_n1703__));
  buf1  g1163(.din(new_new_n857__), .dout(new_new_n1704__));
  buf1  g1164(.din(new_new_n859__), .dout(new_new_n1705__));
  buf1  g1165(.din(new_new_n847__), .dout(new_new_n1706__));
  buf1  g1166(.din(new_new_n520__), .dout(new_new_n1707__));
  buf1  g1167(.din(new_new_n1707__), .dout(new_new_n1708__));
  buf1  g1168(.din(new_new_n1199__), .dout(new_new_n1709__));
  buf1  g1169(.din(new_new_n852__), .dout(new_new_n1710__));
  buf1  g1170(.din(new_new_n1710__), .dout(new_new_n1711__));
  buf1  g1171(.din(new_new_n851__), .dout(new_new_n1712__));
  buf1  g1172(.din(new_new_n1712__), .dout(new_new_n1713__));
  buf1  g1173(.din(new_new_n1712__), .dout(new_new_n1714__));
  buf1  g1174(.din(new_new_n837__), .dout(new_new_n1715__));
  buf1  g1175(.din(new_new_n1715__), .dout(new_new_n1716__));
  buf1  g1176(.din(new_new_n1716__), .dout(new_new_n1717__));
  buf1  g1177(.din(new_new_n1715__), .dout(new_new_n1718__));
  buf1  g1178(.din(new_new_n838__), .dout(new_new_n1719__));
  buf1  g1179(.din(new_new_n1719__), .dout(new_new_n1720__));
  buf1  g1180(.din(new_new_n1719__), .dout(new_new_n1721__));
  buf1  g1181(.din(new_new_n836__), .dout(new_new_n1722__));
  buf1  g1182(.din(new_new_n1722__), .dout(new_new_n1723__));
  buf1  g1183(.din(new_new_n835__), .dout(new_new_n1724__));
  buf1  g1184(.din(new_new_n1724__), .dout(new_new_n1725__));
  buf1  g1185(.din(new_new_n1724__), .dout(new_new_n1726__));
  buf1  g1186(.din(new_new_n1135__), .dout(new_new_n1727__));
  buf1  g1187(.din(new_new_n834__), .dout(new_new_n1728__));
  buf1  g1188(.din(new_new_n833__), .dout(new_new_n1729__));
  buf1  g1189(.din(new_new_n1729__), .dout(new_new_n1730__));
  buf1  g1190(.din(new_new_n493__), .dout(new_new_n1731__));
  buf1  g1191(.din(new_new_n839__), .dout(new_new_n1732__));
  buf1  g1192(.din(new_new_n1732__), .dout(new_new_n1733__));
  buf1  g1193(.din(new_new_n1733__), .dout(new_new_n1734__));
  buf1  g1194(.din(new_new_n1732__), .dout(new_new_n1735__));
  buf1  g1195(.din(new_new_n840__), .dout(new_new_n1736__));
  buf1  g1196(.din(new_new_n1736__), .dout(new_new_n1737__));
  buf1  g1197(.din(new_new_n1736__), .dout(new_new_n1738__));
  buf1  g1198(.din(new_new_n501__), .dout(new_new_n1739__));
  buf1  g1199(.din(new_new_n854__), .dout(new_new_n1740__));
  buf1  g1200(.din(new_new_n853__), .dout(new_new_n1741__));
  buf1  g1201(.din(new_new_n1741__), .dout(new_new_n1742__));
  buf1  g1202(.din(new_new_n519__), .dout(new_new_n1743__));
  buf1  g1203(.din(new_new_n1187__), .dout(new_new_n1744__));
  buf1  g1204(.din(new_new_n1744__), .dout(new_new_n1745__));
  buf1  g1205(.din(new_new_n1252__), .dout(new_new_n1746__));
  always @ (posedge clock) begin
    n940_lo <= n2688;
    n949_lo <= n2691;
    n961_lo <= n2694;
    n973_lo <= n2697;
    n976_lo <= n2700;
    n985_lo <= n2703;
    n988_lo <= n2706;
    n997_lo <= n2709;
    n1009_lo <= n2712;
    n1021_lo <= n2715;
    n1033_lo <= n2718;
    n1045_lo <= n2721;
    n1057_lo <= n2724;
    n1060_lo <= n2727;
    n1069_lo <= n2730;
    n1081_lo <= n2733;
    n1093_lo <= n2736;
    n1105_lo <= n2739;
    n1117_lo <= n2742;
    n1120_lo <= n2745;
    n1129_lo <= n2748;
    n1132_lo <= n2751;
    n1156_lo <= n2754;
    n1168_lo <= n2757;
    n1180_lo <= n2760;
    n1189_lo <= n2763;
    n1192_lo <= n2766;
    n1195_lo <= n2769;
    n1201_lo <= n2772;
    n1204_lo <= n2775;
    n1228_lo <= n2778;
    n1231_lo <= n2781;
    n1234_lo <= n2784;
    n1237_lo <= n2787;
    n1240_lo <= n2790;
    n1243_lo <= n2793;
    n1249_lo <= n2796;
    n1252_lo <= n2799;
    n1255_lo <= n2802;
    n1261_lo <= n2805;
    n1264_lo <= n2808;
    n1267_lo <= n2811;
    n1273_lo <= n2814;
    n1276_lo <= n2817;
    n1279_lo <= n2820;
    n1282_lo <= n2823;
    n1285_lo <= n2826;
    n1288_lo <= n2829;
    n1291_lo <= n2832;
    n1294_lo <= n2835;
    n1297_lo <= n2838;
    n1300_lo <= n2841;
    n1303_lo <= n2844;
    n1309_lo <= n2847;
    n1312_lo <= n2850;
    n1315_lo <= n2853;
    n1318_lo <= n2856;
    n1321_lo <= n2859;
    n1333_lo <= n2862;
    n1225_o2 <= n2865;
    n1229_o2 <= n2868;
    n1228_o2 <= n2871;
    n1259_o2 <= n2874;
    n1272_o2 <= n2877;
    n1269_o2 <= n2880;
    n1307_o2 <= n2883;
    n1201_o2 <= n2886;
    n1202_o2 <= n2889;
    n1203_o2 <= n2892;
    n1204_o2 <= n2895;
    n622_o2 <= n2898;
    n1205_o2 <= n2901;
    n1206_o2 <= n2904;
    n497_o2 <= n2907;
    n1212_o2 <= n2910;
    n1213_o2 <= n2913;
    n1214_o2 <= n2916;
    n1215_o2 <= n2919;
    n1216_o2 <= n2922;
    n1217_o2 <= n2925;
    n1218_o2 <= n2928;
    n1219_o2 <= n2931;
    n1242_o2 <= n2934;
    n1243_o2 <= n2937;
    n1273_o2 <= n2940;
    n1274_o2 <= n2943;
    n1275_o2 <= n2946;
    n1276_o2 <= n2949;
    n1277_o2 <= n2952;
    n1286_o2 <= n2955;
    n1299_o2 <= n2958;
    n601_o2 <= n2961;
    n625_o2 <= n2964;
    n463_o2 <= n2967;
    lo082_buf_o2 <= n2970;
    n455_o2 <= n2973;
    n642_o2 <= n2976;
    n459_o2 <= n2979;
    n501_o2 <= n2982;
    n599_o2 <= n2985;
    n485_o2 <= n2988;
    lo086_buf_o2 <= n2991;
    lo122_buf_o2 <= n2994;
    n502_o2 <= n2997;
    n627_o2 <= n3000;
    lo038_buf_o2 <= n3003;
    lo046_buf_o2 <= n3006;
    lo050_buf_o2 <= n3009;
    lo058_buf_o2 <= n3012;
    lo070_buf_o2 <= n3015;
    lo094_buf_o2 <= n3018;
    n462_o2 <= n3021;
    lo006_buf_o2 <= n3024;
    lo010_buf_o2 <= n3027;
    lo022_buf_o2 <= n3030;
    lo026_buf_o2 <= n3033;
    lo030_buf_o2 <= n3036;
    lo034_buf_o2 <= n3039;
    lo054_buf_o2 <= n3042;
    lo130_buf_o2 <= n3045;
    n547_o2 <= n3048;
    n424_inv <= n3051;
    n617_o2 <= n3054;
    lo042_buf_o2 <= n3057;
    lo062_buf_o2 <= n3060;
    lo110_buf_o2 <= n3063;
    n733_o2 <= n3066;
    n734_o2 <= n3069;
    n570_o2 <= n3072;
    n461_o2 <= n3075;
    n644_o2 <= n3078;
    n628_o2 <= n3081;
    n528_o2 <= n3084;
    n460_inv <= n3087;
    lo002_buf_o2 <= n3090;
    lo014_buf_o2 <= n3093;
    lo018_buf_o2 <= n3096;
    lo078_buf_o2 <= n3099;
    lo090_buf_o2 <= n3102;
    n513_o2 <= n3105;
    lo102_buf_o2 <= n3108;
    lo106_buf_o2 <= n3111;
    n600_o2 <= n3114;
    n529_o2 <= n3117;
    n593_o2 <= n3120;
    lo066_buf_o2 <= n3123;
    n549_o2 <= n3126;
    n550_o2 <= n3129;
    n571_o2 <= n3132;
    n572_o2 <= n3135;
    n495_o2 <= n3138;
    n496_o2 <= n3141;
    n620_o2 <= n3144;
    n482_o2 <= n3147;
    lo081_buf_o2 <= n3150;
    n576_o2 <= n3153;
    n520_o2 <= n3156;
    n521_o2 <= n3159;
    n562_o2 <= n3162;
    n508_o2 <= n3165;
    n509_o2 <= n3168;
    lo074_buf_o2 <= n3171;
    n539_o2 <= n3174;
    n536_o2 <= n3177;
    n516_o2 <= n3180;
    n491_o2 <= n3183;
    n557_o2 <= n3186;
    n586_o2 <= n3189;
    n483_o2 <= n3192;
    n484_o2 <= n3195;
    lo004_buf_o2 <= n3198;
    lo008_buf_o2 <= n3201;
    lo020_buf_o2 <= n3204;
    lo024_buf_o2 <= n3207;
    lo028_buf_o2 <= n3210;
    lo032_buf_o2 <= n3213;
    lo052_buf_o2 <= n3216;
    lo128_buf_o2 <= n3219;
    lo037_buf_o2 <= n3222;
    lo045_buf_o2 <= n3225;
    lo049_buf_o2 <= n3228;
    lo057_buf_o2 <= n3231;
    lo069_buf_o2 <= n3234;
    lo093_buf_o2 <= n3237;
  end
  initial begin
    n940_lo <= 1'b0;
    n949_lo <= 1'b0;
    n961_lo <= 1'b0;
    n973_lo <= 1'b0;
    n976_lo <= 1'b0;
    n985_lo <= 1'b0;
    n988_lo <= 1'b0;
    n997_lo <= 1'b0;
    n1009_lo <= 1'b0;
    n1021_lo <= 1'b0;
    n1033_lo <= 1'b0;
    n1045_lo <= 1'b0;
    n1057_lo <= 1'b0;
    n1060_lo <= 1'b0;
    n1069_lo <= 1'b0;
    n1081_lo <= 1'b0;
    n1093_lo <= 1'b0;
    n1105_lo <= 1'b0;
    n1117_lo <= 1'b0;
    n1120_lo <= 1'b0;
    n1129_lo <= 1'b0;
    n1132_lo <= 1'b0;
    n1156_lo <= 1'b0;
    n1168_lo <= 1'b0;
    n1180_lo <= 1'b0;
    n1189_lo <= 1'b0;
    n1192_lo <= 1'b0;
    n1195_lo <= 1'b0;
    n1201_lo <= 1'b0;
    n1204_lo <= 1'b0;
    n1228_lo <= 1'b0;
    n1231_lo <= 1'b0;
    n1234_lo <= 1'b0;
    n1237_lo <= 1'b0;
    n1240_lo <= 1'b0;
    n1243_lo <= 1'b0;
    n1249_lo <= 1'b0;
    n1252_lo <= 1'b0;
    n1255_lo <= 1'b0;
    n1261_lo <= 1'b0;
    n1264_lo <= 1'b0;
    n1267_lo <= 1'b0;
    n1273_lo <= 1'b0;
    n1276_lo <= 1'b0;
    n1279_lo <= 1'b0;
    n1282_lo <= 1'b0;
    n1285_lo <= 1'b0;
    n1288_lo <= 1'b0;
    n1291_lo <= 1'b0;
    n1294_lo <= 1'b0;
    n1297_lo <= 1'b0;
    n1300_lo <= 1'b0;
    n1303_lo <= 1'b0;
    n1309_lo <= 1'b0;
    n1312_lo <= 1'b0;
    n1315_lo <= 1'b0;
    n1318_lo <= 1'b0;
    n1321_lo <= 1'b0;
    n1333_lo <= 1'b0;
    n1225_o2 <= 1'b0;
    n1229_o2 <= 1'b0;
    n1228_o2 <= 1'b0;
    n1259_o2 <= 1'b0;
    n1272_o2 <= 1'b0;
    n1269_o2 <= 1'b0;
    n1307_o2 <= 1'b0;
    n1201_o2 <= 1'b0;
    n1202_o2 <= 1'b0;
    n1203_o2 <= 1'b0;
    n1204_o2 <= 1'b0;
    n622_o2 <= 1'b0;
    n1205_o2 <= 1'b0;
    n1206_o2 <= 1'b0;
    n497_o2 <= 1'b0;
    n1212_o2 <= 1'b0;
    n1213_o2 <= 1'b0;
    n1214_o2 <= 1'b0;
    n1215_o2 <= 1'b0;
    n1216_o2 <= 1'b0;
    n1217_o2 <= 1'b0;
    n1218_o2 <= 1'b0;
    n1219_o2 <= 1'b0;
    n1242_o2 <= 1'b0;
    n1243_o2 <= 1'b0;
    n1273_o2 <= 1'b0;
    n1274_o2 <= 1'b0;
    n1275_o2 <= 1'b0;
    n1276_o2 <= 1'b0;
    n1277_o2 <= 1'b0;
    n1286_o2 <= 1'b0;
    n1299_o2 <= 1'b0;
    n601_o2 <= 1'b0;
    n625_o2 <= 1'b0;
    n463_o2 <= 1'b0;
    lo082_buf_o2 <= 1'b0;
    n455_o2 <= 1'b0;
    n642_o2 <= 1'b0;
    n459_o2 <= 1'b0;
    n501_o2 <= 1'b0;
    n599_o2 <= 1'b0;
    n485_o2 <= 1'b0;
    lo086_buf_o2 <= 1'b0;
    lo122_buf_o2 <= 1'b0;
    n502_o2 <= 1'b0;
    n627_o2 <= 1'b0;
    lo038_buf_o2 <= 1'b0;
    lo046_buf_o2 <= 1'b0;
    lo050_buf_o2 <= 1'b0;
    lo058_buf_o2 <= 1'b0;
    lo070_buf_o2 <= 1'b0;
    lo094_buf_o2 <= 1'b0;
    n462_o2 <= 1'b0;
    lo006_buf_o2 <= 1'b0;
    lo010_buf_o2 <= 1'b0;
    lo022_buf_o2 <= 1'b0;
    lo026_buf_o2 <= 1'b0;
    lo030_buf_o2 <= 1'b0;
    lo034_buf_o2 <= 1'b0;
    lo054_buf_o2 <= 1'b0;
    lo130_buf_o2 <= 1'b0;
    n547_o2 <= 1'b0;
    n424_inv <= 1'b0;
    n617_o2 <= 1'b0;
    lo042_buf_o2 <= 1'b0;
    lo062_buf_o2 <= 1'b0;
    lo110_buf_o2 <= 1'b0;
    n733_o2 <= 1'b0;
    n734_o2 <= 1'b0;
    n570_o2 <= 1'b0;
    n461_o2 <= 1'b0;
    n644_o2 <= 1'b0;
    n628_o2 <= 1'b0;
    n528_o2 <= 1'b0;
    n460_inv <= 1'b0;
    lo002_buf_o2 <= 1'b0;
    lo014_buf_o2 <= 1'b0;
    lo018_buf_o2 <= 1'b0;
    lo078_buf_o2 <= 1'b0;
    lo090_buf_o2 <= 1'b0;
    n513_o2 <= 1'b0;
    lo102_buf_o2 <= 1'b0;
    lo106_buf_o2 <= 1'b0;
    n600_o2 <= 1'b0;
    n529_o2 <= 1'b0;
    n593_o2 <= 1'b0;
    lo066_buf_o2 <= 1'b0;
    n549_o2 <= 1'b0;
    n550_o2 <= 1'b0;
    n571_o2 <= 1'b0;
    n572_o2 <= 1'b0;
    n495_o2 <= 1'b0;
    n496_o2 <= 1'b0;
    n620_o2 <= 1'b0;
    n482_o2 <= 1'b0;
    lo081_buf_o2 <= 1'b0;
    n576_o2 <= 1'b0;
    n520_o2 <= 1'b0;
    n521_o2 <= 1'b0;
    n562_o2 <= 1'b0;
    n508_o2 <= 1'b0;
    n509_o2 <= 1'b0;
    lo074_buf_o2 <= 1'b0;
    n539_o2 <= 1'b0;
    n536_o2 <= 1'b0;
    n516_o2 <= 1'b0;
    n491_o2 <= 1'b0;
    n557_o2 <= 1'b0;
    n586_o2 <= 1'b0;
    n483_o2 <= 1'b0;
    n484_o2 <= 1'b0;
    lo004_buf_o2 <= 1'b0;
    lo008_buf_o2 <= 1'b0;
    lo020_buf_o2 <= 1'b0;
    lo024_buf_o2 <= 1'b0;
    lo028_buf_o2 <= 1'b0;
    lo032_buf_o2 <= 1'b0;
    lo052_buf_o2 <= 1'b0;
    lo128_buf_o2 <= 1'b0;
    lo037_buf_o2 <= 1'b0;
    lo045_buf_o2 <= 1'b0;
    lo049_buf_o2 <= 1'b0;
    lo057_buf_o2 <= 1'b0;
    lo069_buf_o2 <= 1'b0;
    lo093_buf_o2 <= 1'b0;
  end
endmodule


