module c2670(G1,G10,G100,G101,G102,G103,G104,G105,G106,G107,G108,G109,G11,
  G110,G111,G112,G113,G114,G115,G116,G117,G118,G119,G12,G120,G121,G122,G123,
  G124,G125,G126,G127,G128,G129,G13,G130,G131,G132,G133,G134,G135,G136,G137,
  G138,G139,G14,G140,G141,G142,G143,G144,G145,G146,G147,G148,G149,G15,G150,
  G151,G152,G153,G154,G155,G156,G157,G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,
  G25,G2531,G2532,G2533,G2534,G2535,G2536,G2537,G2538,G2539,G2540,G2541,G2542,
  G2543,G2544,G2545,G2546,G2547,G2548,G2549,G2550,G2551,G2552,G2553,G2554,
  G2555,G2556,G2557,G2558,G2559,G2560,G2561,G2562,G2563,G2564,G2565,G2566,
  G2567,G2568,G2569,G2570,G2571,G2572,G2573,G2574,G2575,G2576,G2577,G2578,
  G2579,G2580,G2581,G2582,G2583,G2584,G2585,G2586,G2587,G2588,G2589,G2590,
  G2591,G2592,G2593,G2594,G26,G27,G28,G29,G3,G30,G31,G32,G33,G34,G35,G36,G37,
  G38,G39,G4,G40,G41,G42,G43,G44,G45,G46,G47,G48,G49,G5,G50,G51,G52,G53,G54,
  G55,G56,G57,G58,G59,G6,G60,G61,G62,G63,G64,G65,G66,G67,G68,G69,G7,G70,G71,
  G72,G73,G74,G75,G76,G77,G78,G79,G8,G80,G81,G82,G83,G84,G85,G86,G87,G88,G89,
  G9,G90,G91,G92,G93,G94,G95,G96,G97,G98,G99);
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
  G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,
  G40,G41,G42,G43,G44,G45,G46,G47,G48,G49,G50,G51,G52,G53,G54,G55,G56,G57,G58,
  G59,G60,G61,G62,G63,G64,G65,G66,G67,G68,G69,G70,G71,G72,G73,G74,G75,G76,G77,
  G78,G79,G80,G81,G82,G83,G84,G85,G86,G87,G88,G89,G90,G91,G92,G93,G94,G95,G96,
  G97,G98,G99,G100,G101,G102,G103,G104,G105,G106,G107,G108,G109,G110,G111,G112,
  G113,G114,G115,G116,G117,G118,G119,G120,G121,G122,G123,G124,G125,G126,G127,
  G128,G129,G130,G131,G132,G133,G134,G135,G136,G137,G138,G139,G140,G141,G142,
  G143,G144,G145,G146,G147,G148,G149,G150,G151,G152,G153,G154,G155,G156,G157;
output G2531,G2532,G2533,G2534,G2535,G2536,G2537,G2538,G2539,G2540,G2541,G2542,
  G2543,G2544,G2545,G2546,G2547,G2548,G2549,G2550,G2551,G2552,G2553,G2554,
  G2555,G2556,G2557,G2558,G2559,G2560,G2561,G2562,G2563,G2564,G2565,G2566,
  G2567,G2568,G2569,G2570,G2571,G2572,G2573,G2574,G2575,G2576,G2577,G2578,
  G2579,G2580,G2581,G2582,G2583,G2584,G2585,G2586,G2587,G2588,G2589,G2590,
  G2591,G2592,G2593,G2594;

  wire G282,G283,G284,G285,G286,G287,G288,G291,G292,G295,G298,G301,G313,G325,
    G329,G335,G336,G339,G342,G354,G366,G370,G374,G386,G398,G399,G400,G401,G402,
    G403,G404,G405,G417,G429,G435,G442,G443,G447,G451,G455,G459,G463,G467,G471,
    G475,G479,G485,G491,G497,G503,G507,G511,G515,G519,G522,G525,G526,G527,G530,
    G533,G536,G539,G542,G545,G548,G551,G554,G557,G560,G563,G566,G569,G572,G575,
    G578,G581,G584,G585,G586,G587,G588,G589,G590,G591,G592,G593,G594,G595,G598,
    G603,G614,G625,G626,G627,G628,G629,G630,G631,G636,G647,G658,G659,G660,G661,
    G662,G663,G674,G685,G686,G687,G688,G689,G690,G694,G698,G701,G702,G703,G704,
    G705,G706,G707,G718,G729,G730,G731,G732,G733,G734,G739,G745,G746,G747,G748,
    G749,G750,G751,G756,G761,G766,G771,G772,G773,G774,G775,G776,G777,G780,G783,
    G786,G789,G792,G795,G798,G801,G804,G807,G810,G811,G812,G815,G818,G821,G824,
    G827,G830,G831,G832,G833,G834,G835,G836,G837,G838,G839,G840,G841,G842,G843,
    G844,G845,G846,G847,G848,G849,G850,G851,G852,G853,G854,G855,G856,G857,G858,
    G859,G860,G861,G862,G863,G864,G865,G866,G867,G868,G869,G870,G871,G872,G873,
    G874,G875,G876,G877,G878,G879,G880,G881,G882,G883,G884,G885,G886,G887,G888,
    G889,G890,G891,G892,G893,G894,G895,G896,G897,G898,G901,G904,G908,G912,G915,
    G918,G921,G922,G923,G924,G925,G926,G927,G928,G929,G930,G931,G932,G933,G934,
    G935,G936,G937,G938,G939,G940,G941,G942,G943,G944,G945,G946,G947,G948,G949,
    G950,G951,G952,G953,G954,G955,G959,G963,G966,G967,G968,G969,G970,G971,G972,
    G973,G974,G975,G976,G977,G978,G979,G980,G983,G984,G987,G990,G993,G998,
    G1002,G1008,G1014,G1017,G1021,G1026,G1030,G1033,G1036,G1039,G1044,G1049,
    G1053,G1058,G1062,G1067,G1072,G1076,G1079,G1082,G1085,G1088,G1089,G1090,
    G1093,G1096,G1097,G1098,G1101,G1104,G1107,G1110,G1111,G1112,G1113,G1114,
    G1115,G1116,G1117,G1118,G1119,G1120,G1123,G1126,G1127,G1128,G1129,G1132,
    G1137,G1144,G1148,G1152,G1159,G1166,G1171,G1176,G1181,G1184,G1187,G1190,
    G1193,G1196,G1197,G1198,G1199,G1200,G1201,G1202,G1203,G1204,G1205,G1206,
    G1207,G1208,G1209,G1210,G1211,G1212,G1213,G1214,G1215,G1216,G1219,G1220,
    G1221,G1222,G1225,G1228,G1231,G1234,G1237,G1240,G1243,G1246,G1249,G1250,
    G1251,G1252,G1253,G1254,G1255,G1256,G1257,G1258,G1259,G1260,G1263,G1266,
    G1269,G1272,G1275,G1278,G1281,G1284,G1287,G1290,G1293,G1296,G1299,G1302,
    G1305,G1308,G1311,G1314,G1320,G1321,G1326,G1327,G1328,G1329,G1336,G1342,
    G1345,G1348,G1351,G1354,G1355,G1356,G1357,G1358,G1359,G1360,G1361,G1362,
    G1363,G1364,G1365,G1366,G1367,G1368,G1371,G1374,G1377,G1380,G1383,G1384,
    G1387,G1390,G1393,G1396,G1399,G1402,G1405,G1406,G1407,G1408,G1409,G1412,
    G1415,G1418,G1421,G1424,G1425,G1426,G1427,G1428,G1429,G1430,G1431,G1432,
    G1433,G1434,G1435,G1436,G1437,G1438,G1439,G1440,G1441,G1442,G1443,G1444,
    G1445,G1446,G1447,G1448,G1449,G1450,G1451,G1452,G1453,G1454,G1455,G1456,
    G1457,G1458,G1459,G1460,G1461,G1462,G1463,G1464,G1465,G1466,G1467,G1468,
    G1469,G1470,G1471,G1472,G1475,G1476,G1477,G1478,G1479,G1483,G1484,G1485,
    G1486,G1487,G1488,G1493,G1497,G1498,G1502,G1507,G1508,G1509,G1510,G1511,
    G1512,G1513,G1514,G1515,G1516,G1517,G1518,G1519,G1520,G1524,G1528,G1531,
    G1532,G1533,G1534,G1535,G1536,G1537,G1540,G1543,G1546,G1549,G1552,G1555,
    G1556,G1557,G1560,G1563,G1566,G1569,G1572,G1575,G1578,G1581,G1584,G1587,
    G1590,G1593,G1596,G1599,G1600,G1601,G1602,G1603,G1606,G1607,G1610,G1613,
    G1616,G1619,G1620,G1621,G1622,G1623,G1624,G1625,G1626,G1627,G1628,G1629,
    G1630,G1631,G1632,G1633,G1634,G1635,G1636,G1640,G1641,G1642,G1643,G1644,
    G1645,G1646,G1650,G1651,G1652,G1653,G1654,G1657,G1661,G1662,G1663,G1664,
    G1665,G1666,G1667,G1668,G1669,G1670,G1675,G1676,G1681,G1682,G1683,G1684,
    G1688,G1689,G1690,G1691,G1692,G1693,G1694,G1695,G1696,G1697,G1698,G1699,
    G1700,G1701,G1702,G1703,G1704,G1705,G1706,G1709,G1712,G1715,G1718,G1719,
    G1720,G1721,G1722,G1723,G1724,G1725,G1726,G1727,G1728,G1731,G1732,G1733,
    G1734,G1735,G1736,G1737,G1738,G1739,G1744,G1749,G1750,G1751,G1752,G1753,
    G1754,G1755,G1756,G1761,G1766,G1767,G1768,G1769,G1770,G1771,G1772,G1773,
    G1774,G1775,G1776,G1777,G1778,G1779,G1780,G1781,G1782,G1785,G1789,G1792,
    G1795,G1798,G1799,G1800,G1801,G1802,G1805,G1811,G1814,G1815,G1816,G1822,
    G1823,G1824,G1825,G1826,G1829,G1835,G1840,G1846,G1851,G1854,G1857,G1858,
    G1859,G1862,G1865,G1868,G1869,G1870,G1871,G1872,G1873,G1874,G1875,G1876,
    G1877,G1878,G1879,G1880,G1881,G1882,G1883,G1884,G1887,G1888,G1889,G1890,
    G1893,G1896,G1899,G1902,G1903,G1904,G1907,G1910,G1913,G1916,G1919,G1922,
    G1925,G1926,G1927,G1928,G1931,G1934,G1937,G1940,G1943,G1946,G1947,G1948,
    G1953,G1954,G1955,G1956,G1961,G1962,G1963,G1964,G1965,G1966,G1967,G1970,
    G1971,G1972,G1973,G1974,G1975,G1976,G1977,G1978,G1981,G1982,G1983,G1984,
    G1985,G1986,G1987,G1988,G1989,G1990,G1991,G1992,G1993,G1996,G1999,G2002,
    G2005,G2008,G2011,G2014,G2017,G2020,G2023,G2026,G2029,G2032,G2035,G2038,
    G2041,G2044,G2045,G2046,G2047,G2048,G2051,G2052,G2053,G2054,G2055,G2056,
    G2057,G2058,G2059,G2060,G2061,G2062,G2063,G2064,G2065,G2066,G2067,G2068,
    G2069,G2070,G2071,G2072,G2073,G2076,G2079,G2082,G2085,G2088,G2091,G2094,
    G2097,G2100,G2103,G2106,G2109,G2112,G2115,G2116,G2117,G2118,G2119,G2120,
    G2121,G2122,G2123,G2124,G2125,G2126,G2127,G2128,G2129,G2130,G2131,G2132,
    G2133,G2134,G2135,G2138,G2141,G2144,G2147,G2150,G2153,G2154,G2155,G2156,
    G2157,G2158,G2161,G2164,G2167,G2170,G2173,G2176,G2179,G2182,G2185,G2188,
    G2191,G2194,G2197,G2200,G2203,G2206,G2207,G2208,G2209,G2210,G2211,G2212,
    G2213,G2214,G2215,G2216,G2217,G2218,G2219,G2220,G2221,G2222,G2223,G2224,
    G2225,G2226,G2227,G2228,G2231,G2234,G2237,G2240,G2241,G2242,G2243,G2244,
    G2245,G2246,G2247,G2248,G2249,G2250,G2251,G2252,G2253,G2254,G2255,G2256,
    G2257,G2258,G2259,G2260,G2261,G2262,G2263,G2264,G2265,G2266,G2267,G2268,
    G2269,G2270,G2271,G2272,G2273,G2274,G2275,G2276,G2279,G2282,G2285,G2288,
    G2291,G2294,G2297,G2300,G2301,G2302,G2303,G2304,G2305,G2306,G2307,G2308,
    G2309,G2310,G2311,G2312,G2313,G2314,G2315,G2316,G2317,G2320,G2323,G2326,
    G2329,G2330,G2331,G2332,G2333,G2334,G2335,G2336,G2337,G2340,G2345,G2349,
    G2352,G2353,G2359,G2364,G2365,G2366,G2367,G2368,G2369,G2370,G2375,G2379,
    G2382,G2383,G2389,G2394,G2395,G2396,G2397,G2398,G2399,G2400,G2401,G2402,
    G2403,G2404,G2405,G2406,G2407,G2408,G2409,G2410,G2411,G2412,G2413,G2414,
    G2417,G2418,G2419,G2420,G2421,G2422,G2423,G2424,G2425,G2426,G2427,G2428,
    G2431,G2432,G2433,G2434,G2435,G2436,G2437,G2438,G2439,G2440,G2441,G2442,
    G2443,G2447,G2450,G2451,G2454,G2458,G2461,G2462,G2465,G2466,G2467,G2470,
    G2473,G2474,G2475,G2476,G2477,G2478,G2479,G2480,G2481,G2482,G2483,G2484,
    G2485,G2486,G2487,G2488,G2489,G2490,G2491,G2492,G2495,G2496,G2499,G2500,
    G2501,G2502,G2503,G2504,G2505,G2508,G2512,G2515,G2516,G2517,G2520,G2523,
    G2524,G2527,G2528;

  and (G282,G1,G3);
  not (G283,G118);
  not (G284,G127);
  and (G285,G142,G141,G140,G139);
  not (G286,G282);
  and (G287,G2,G11,G121);
  not (G288,G121);
  and (G291,G29,G29);
  not (G292,G115);
  not (G295,G8);
  not (G298,G8);
  not (G301,G117);
  not (G313,G120);
  not (G325,G122);
  not (G329,G123);
  and (G335,G9,G123);
  and (G336,G106,G64,G76,G32);
  and (G339,G96,G43,G86,G53);
  not (G342,G117);
  not (G354,G120);
  not (G366,G125);
  not (G370,G126);
  not (G374,G145);
  not (G386,G146);
  not (G398,G148);
  not (G399,G149);
  not (G400,G150);
  not (G401,G151);
  not (G402,G152);
  not (G403,G153);
  not (G404,G156);
  not (G405,G145);
  not (G417,G146);
  not (G429,G12);
  not (G435,G12);
  not (G442,G157);
  and (G443,G7,G121);
  not (G447,G128);
  not (G451,G129);
  not (G455,G130);
  not (G459,G131);
  not (G463,G132);
  not (G467,G133);
  not (G471,G134);
  not (G475,G135);
  not (G479,G136);
  not (G485,G23);
  not (G491,G23);
  not (G497,G138);
  not (G503,G139);
  not (G507,G140);
  not (G511,G141);
  not (G515,G142);
  not (G519,G143);
  not (G522,G144);
  not (G525,G154);
  not (G526,G155);
  not (G527,G126);
  not (G530,G125);
  not (G533,G128);
  not (G536,G130);
  not (G539,G129);
  not (G542,G132);
  not (G545,G131);
  not (G548,G134);
  not (G551,G133);
  not (G554,G136);
  not (G557,G135);
  not (G560,G138);
  not (G563,G140);
  not (G566,G139);
  not (G569,G142);
  not (G572,G141);
  not (G575,G144);
  not (G578,G143);
  not (G581,G291);
  nand (G584,G149,G398);
  nand (G585,G148,G399);
  nand (G586,G151,G400);
  nand (G587,G150,G401);
  nand (G588,G153,G402);
  nand (G589,G152,G403);
  nand (G590,G155,G525);
  nand (G591,G154,G526);
  and (G592,G147,G443);
  not (G593,G336);
  not (G594,G339);
  and (G595,G339,G336);
  not (G598,G295);
  not (G603,G301);
  not (G614,G313);
  and (G625,G62,G301,G313);
  and (G626,G52,G301,G313);
  and (G627,G61,G301,G313);
  and (G628,G60,G301,G313);
  and (G629,G59,G301,G313);
  and (G630,G9,G329);
  not (G631,G295);
  not (G636,G342);
  not (G647,G354);
  and (G658,G58,G342,G354);
  and (G659,G57,G342,G354);
  and (G660,G56,G342,G354);
  and (G661,G55,G342,G354);
  and (G662,G54,G342,G354);
  not (G663,G374);
  not (G674,G386);
  and (G685,G90,G374,G386);
  and (G686,G89,G374,G386);
  and (G687,G88,G374,G386);
  and (G688,G87,G374,G386);
  and (G689,G374,G386);
  nand (G690,G584,G585);
  nand (G694,G586,G587);
  nand (G698,G588,G589);
  not (G701,G533);
  nand (G702,G533,G404);
  not (G703,G536);
  not (G704,G539);
  not (G705,G542);
  not (G706,G545);
  not (G707,G405);
  not (G718,G417);
  and (G729,G94,G405,G417);
  and (G730,G85,G405,G417);
  and (G731,G93,G405,G417);
  and (G732,G92,G405,G417);
  and (G733,G91,G405,G417);
  not (G734,G429);
  not (G739,G435);
  not (G745,G560);
  nand (G746,G560,G442);
  not (G747,G563);
  not (G748,G566);
  not (G749,G569);
  not (G750,G572);
  not (G751,G298);
  not (G756,G298);
  not (G761,G485);
  not (G766,G491);
  not (G771,G527);
  not (G772,G530);
  not (G773,G548);
  not (G774,G551);
  not (G775,G554);
  not (G776,G557);
  nand (G777,G590,G591);
  not (G780,G366);
  not (G783,G370);
  not (G786,G447);
  not (G789,G451);
  not (G792,G455);
  not (G795,G459);
  not (G798,G463);
  not (G801,G467);
  not (G804,G471);
  not (G807,G475);
  not (G810,G575);
  not (G811,G578);
  not (G812,G479);
  not (G815,G497);
  not (G818,G503);
  not (G821,G507);
  not (G824,G511);
  not (G827,G515);
  and (G830,G147,G593);
  and (G831,G119,G594);
  or (G832,G630,G335);
  nand (G833,G156,G701);
  nand (G834,G539,G703);
  nand (G835,G536,G704);
  nand (G836,G545,G705);
  nand (G837,G542,G706);
  nand (G838,G157,G745);
  nand (G839,G566,G747);
  nand (G840,G563,G748);
  nand (G841,G572,G749);
  nand (G842,G569,G750);
  nand (G843,G530,G771);
  nand (G844,G527,G772);
  nand (G845,G551,G773);
  nand (G846,G548,G774);
  nand (G847,G557,G775);
  nand (G848,G554,G776);
  nand (G849,G578,G810);
  nand (G850,G575,G811);
  not (G851,G830);
  not (G852,G831);
  and (G853,G73,G603,G614);
  and (G854,G41,G301,G614);
  and (G855,G51,G603,G313);
  and (G856,G63,G603,G614);
  and (G857,G31,G301,G614);
  and (G858,G42,G603,G313);
  and (G859,G72,G603,G614);
  and (G860,G40,G301,G614);
  and (G861,G50,G603,G313);
  and (G862,G71,G603,G614);
  and (G863,G39,G301,G614);
  and (G864,G49,G603,G313);
  and (G865,G70,G603,G614);
  and (G866,G38,G301,G614);
  and (G867,G48,G603,G313);
  and (G868,G69,G636,G647);
  and (G869,G37,G342,G647);
  and (G870,G47,G636,G354);
  and (G871,G68,G636,G647);
  and (G872,G36,G342,G647);
  and (G873,G46,G636,G354);
  and (G874,G67,G636,G647);
  and (G875,G35,G342,G647);
  and (G876,G636,G354);
  and (G877,G66,G636,G647);
  and (G878,G34,G342,G647);
  and (G879,G45,G636,G354);
  and (G880,G65,G636,G647);
  and (G881,G33,G342,G647);
  and (G882,G44,G636,G354);
  and (G883,G110,G663,G674);
  and (G884,G80,G374,G674);
  and (G885,G100,G663,G386);
  and (G886,G109,G663,G674);
  and (G887,G79,G374,G674);
  and (G888,G99,G663,G386);
  and (G889,G108,G663,G674);
  and (G890,G78,G374,G674);
  and (G891,G98,G663,G386);
  and (G892,G107,G663,G674);
  and (G893,G77,G374,G674);
  and (G894,G97,G663,G386);
  and (G895,G663,G674);
  and (G896,G374,G674);
  and (G897,G663,G386);
  not (G898,G690);
  not (G901,G694);
  nand (G904,G833,G702);
  nand (G908,G834,G835);
  nand (G912,G836,G837);
  not (G915,G698);
  not (G918,G698);
  not (G921,G780);
  not (G922,G783);
  not (G923,G786);
  not (G924,G789);
  not (G925,G792);
  not (G926,G795);
  not (G927,G798);
  not (G928,G801);
  not (G929,G804);
  not (G930,G807);
  and (G931,G114,G707,G718);
  and (G932,G84,G405,G718);
  and (G933,G104,G707,G417);
  and (G934,G105,G707,G718);
  and (G935,G75,G405,G718);
  and (G936,G95,G707,G417);
  and (G937,G113,G707,G718);
  and (G938,G83,G405,G718);
  and (G939,G103,G707,G417);
  and (G940,G112,G707,G718);
  and (G941,G82,G405,G718);
  and (G942,G102,G707,G417);
  and (G943,G111,G707,G718);
  and (G944,G81,G405,G718);
  and (G945,G101,G707,G417);
  and (G946,G13,G734);
  and (G947,G4,G734);
  and (G948,G14,G734);
  and (G949,G5,G734);
  and (G950,G15,G739);
  and (G951,G16,G739);
  and (G952,G17,G739);
  and (G953,G6,G739);
  and (G954,G18,G739);
  nand (G955,G838,G746);
  nand (G959,G839,G840);
  nand (G963,G841,G842);
  and (G966,G19,G761);
  and (G967,G24,G761);
  and (G968,G20,G761);
  and (G969,G25,G761);
  and (G970,G21,G766);
  and (G971,G26,G766);
  and (G972,G27,G766);
  and (G973,G22,G766);
  not (G974,G812);
  not (G975,G815);
  not (G976,G818);
  not (G977,G821);
  not (G978,G824);
  not (G979,G827);
  nand (G980,G843,G844);
  not (G983,G777);
  nand (G984,G847,G848);
  nand (G987,G845,G846);
  nand (G990,G849,G850);
  and (G993,G851,G852);
  or (G998,G853,G854,G855,G625);
  or (G1002,G856,G857,G858,G626);
  or (G1008,G859,G860,G861,G627);
  or (G1014,G862,G863,G864,G628);
  or (G1017,G865,G866,G867,G629);
  or (G1021,G868,G869,G870,G658);
  or (G1026,G871,G872,G873,G659);
  or (G1030,G874,G875,G876,G660);
  or (G1033,G877,G878,G879,G661);
  or (G1036,G880,G881,G882,G662);
  or (G1039,G883,G884,G885,G685);
  or (G1044,G886,G887,G888,G686);
  or (G1049,G889,G890,G891,G687);
  or (G1053,G892,G893,G894,G688);
  or (G1058,G895,G896,G897,G689);
  or (G1062,G934,G935,G936,G730);
  or (G1067,G937,G938,G939,G731);
  or (G1072,G940,G941,G942,G732);
  or (G1076,G943,G944,G945,G733);
  or (G1079,G931,G932,G933,G729);
  not (G1082,G904);
  not (G1085,G908);
  not (G1088,G915);
  not (G1089,G918);
  not (G1090,G912);
  not (G1093,G912);
  and (G1096,G694,G690,G915);
  and (G1097,G901,G898,G918);
  not (G1098,G955);
  not (G1101,G959);
  not (G1104,G963);
  not (G1107,G963);
  not (G1110,G990);
  not (G1111,G980);
  nand (G1112,G980,G983);
  not (G1113,G984);
  not (G1114,G987);
  and (G1115,G998,G122);
  and (G1116,G1008,G122);
  and (G1117,G1002,G122);
  and (G1118,G288,G116,G28,G993);
  and (G1119,G288,G116,G993,G286);
  not (G1120,G998);
  not (G1123,G1008);
  and (G1126,G1002,G329);
  and (G1127,G1008,G329);
  and (G1128,G1021,G123);
  not (G1129,G998);
  not (G1132,G1002);
  not (G1137,G1008);
  not (G1144,G1014);
  not (G1148,G1017);
  not (G1152,G1021);
  not (G1159,G1026);
  not (G1166,G1030);
  not (G1171,G1033);
  not (G1176,G1036);
  nand (G1181,G519,G1053);
  nand (G1184,G522,G1058);
  not (G1187,G1072);
  and (G1190,G1039,G284);
  not (G1193,G1044);
  and (G1196,G898,G694,G1088);
  and (G1197,G690,G901,G1089);
  and (G1198,G1002,G429);
  and (G1199,G1008,G429);
  and (G1200,G1014,G429);
  and (G1201,G1017,G429);
  and (G1202,G1021,G435);
  and (G1203,G1026,G435);
  and (G1204,G1030,G435);
  and (G1205,G1033,G435);
  and (G1206,G1036,G435);
  not (G1207,G1079);
  and (G1208,G1062,G485);
  and (G1209,G1067,G485);
  and (G1210,G1072,G485);
  and (G1211,G1076,G485);
  and (G1212,G1039,G491);
  and (G1213,G1044,G491);
  and (G1214,G1049,G491);
  and (G1215,G1053,G491);
  not (G1216,G1002);
  nand (G1219,G777,G1111);
  nand (G1220,G987,G1113);
  nand (G1221,G984,G1114);
  not (G1222,G1062);
  not (G1225,G1072);
  not (G1228,G1067);
  not (G1231,G1039);
  not (G1234,G1076);
  not (G1237,G1049);
  not (G1240,G1044);
  not (G1243,G1058);
  not (G1246,G1053);
  not (G1249,G1090);
  not (G1250,G1093);
  nor (G1251,G1196,G1096);
  nor (G1252,G1197,G1097);
  and (G1253,G908,G904,G1090);
  and (G1254,G1085,G1082,G1093);
  or (G1255,G973,G1215);
  not (G1256,G1104);
  not (G1257,G1107);
  and (G1258,G959,G955,G1104);
  and (G1259,G1101,G1098,G1107);
  nand (G1260,G1219,G1112);
  nand (G1263,G1220,G1221);
  or (G1266,G946,G1198);
  or (G1269,G947,G1199);
  or (G1272,G948,G1200);
  or (G1275,G949,G1201);
  or (G1278,G950,G1202);
  or (G1281,G951,G1203);
  or (G1284,G952,G1204);
  or (G1287,G953,G1205);
  or (G1290,G954,G1206);
  or (G1293,G966,G1208);
  or (G1296,G967,G1209);
  or (G1299,G968,G1210);
  or (G1302,G969,G1211);
  or (G1305,G970,G1212);
  or (G1308,G971,G1213);
  or (G1311,G972,G1214);
  and (G1314,G1193,G1190,G30);
  not (G1320,G1190);
  nand (G1321,G283,G1123);
  and (G1326,G1120,G329);
  and (G1327,G1148,G123);
  and (G1328,G1144,G329);
  not (G1329,G1144);
  not (G1336,G1148);
  not (G1342,G1159);
  not (G1345,G1166);
  not (G1348,G1171);
  not (G1351,G1176);
  and (G1354,G519,G1181);
  and (G1355,G1181,G1053);
  and (G1356,G522,G1184);
  and (G1357,G1184,G1058);
  and (G1358,G1082,G908,G1249);
  and (G1359,G904,G1085,G1250);
  not (G1360,G1222);
  nand (G1361,G1222,G1207);
  not (G1362,G1225);
  not (G1363,G1228);
  not (G1364,G1231);
  not (G1365,G1234);
  and (G1366,G1098,G959,G1256);
  and (G1367,G955,G1101,G1257);
  not (G1368,G1132);
  not (G1371,G1129);
  not (G1374,G1137);
  not (G1377,G1152);
  not (G1380,G1123);
  not (G1383,G1216);
  not (G1384,G1132);
  not (G1387,G1129);
  not (G1390,G1137);
  not (G1393,G1120);
  not (G1396,G1137);
  not (G1399,G1137);
  nand (G1402,G1252,G1251);
  not (G1405,G1237);
  not (G1406,G1240);
  not (G1407,G1243);
  not (G1408,G1246);
  and (G1409,G30,G1193,G1320);
  or (G1412,G1127,G1327);
  or (G1415,G1328,G1128);
  or (G1418,G1354,G1355);
  or (G1421,G1356,G1357);
  nor (G1424,G1358,G1253);
  nor (G1425,G1359,G1254);
  not (G1426,G1260);
  not (G1427,G1263);
  nand (G1428,G1266,G921);
  not (G1429,G1266);
  nand (G1430,G1269,G922);
  not (G1431,G1269);
  nand (G1432,G1272,G923);
  not (G1433,G1272);
  nand (G1434,G1275,G924);
  not (G1435,G1275);
  nand (G1436,G1278,G925);
  not (G1437,G1278);
  nand (G1438,G1281,G926);
  not (G1439,G1281);
  nand (G1440,G1284,G927);
  not (G1441,G1284);
  nand (G1442,G1287,G928);
  not (G1443,G1287);
  nand (G1444,G1290,G929);
  not (G1445,G1290);
  nand (G1446,G1293,G930);
  not (G1447,G1293);
  nand (G1448,G1079,G1360);
  nand (G1449,G1228,G1362);
  nand (G1450,G1225,G1363);
  nand (G1451,G1234,G1364);
  nand (G1452,G1231,G1365);
  nor (G1453,G1366,G1258);
  nor (G1454,G1367,G1259);
  nand (G1455,G1296,G974);
  not (G1456,G1296);
  nand (G1457,G1299,G975);
  not (G1458,G1299);
  nand (G1459,G1302,G976);
  not (G1460,G1302);
  nand (G1461,G1305,G977);
  not (G1462,G1305);
  nand (G1463,G1308,G978);
  not (G1464,G1308);
  nand (G1465,G1311,G979);
  not (G1466,G1311);
  nand (G1467,G1240,G1405);
  nand (G1468,G1237,G1406);
  nand (G1469,G1246,G1407);
  nand (G1470,G1243,G1408);
  and (G1471,G1321,G325);
  not (G1472,G1314);
  not (G1475,G1368);
  not (G1476,G1371);
  not (G1477,G1374);
  not (G1478,G1377);
  not (G1479,G1321);
  not (G1483,G1384);
  not (G1484,G1387);
  not (G1485,G1390);
  not (G1486,G1393);
  not (G1487,G1396);
  not (G1488,G1314);
  not (G1493,G1314);
  and (G1497,G1321,G123);
  not (G1498,G1314);
  not (G1502,G1314);
  nand (G1507,G1402,G1426);
  not (G1508,G1399);
  not (G1509,G1402);
  nand (G1510,G780,G1429);
  nand (G1511,G783,G1431);
  nand (G1512,G786,G1433);
  nand (G1513,G789,G1435);
  nand (G1514,G792,G1437);
  nand (G1515,G795,G1439);
  nand (G1516,G798,G1441);
  nand (G1517,G801,G1443);
  nand (G1518,G804,G1445);
  nand (G1519,G807,G1447);
  nand (G1520,G1448,G1361);
  nand (G1524,G1449,G1450);
  nand (G1528,G1451,G1452);
  nand (G1531,G812,G1456);
  nand (G1532,G815,G1458);
  nand (G1533,G818,G1460);
  nand (G1534,G821,G1462);
  nand (G1535,G824,G1464);
  nand (G1536,G827,G1466);
  not (G1537,G1329);
  not (G1540,G1336);
  not (G1543,G1345);
  not (G1546,G1342);
  not (G1549,G1351);
  not (G1552,G1348);
  not (G1555,G1380);
  nand (G1556,G1380,G1383);
  not (G1557,G1329);
  not (G1560,G1345);
  not (G1563,G1342);
  not (G1566,G1351);
  not (G1569,G1348);
  not (G1572,G1321);
  not (G1575,G1329);
  not (G1578,G1336);
  not (G1581,G1329);
  not (G1584,G1336);
  nand (G1587,G1425,G1424);
  nand (G1590,G1469,G1470);
  nand (G1593,G1467,G1468);
  nand (G1596,G1454,G1453);
  nand (G1599,G1371,G1475);
  nand (G1600,G1368,G1476);
  nand (G1601,G1387,G1483);
  nand (G1602,G1384,G1484);
  or (G1603,G1126,G1497);
  nand (G1606,G1260,G1509);
  not (G1607,G1418);
  not (G1610,G1421);
  not (G1613,G1409);
  not (G1616,G1409);
  nand (G1619,G1428,G1510);
  nand (G1620,G1430,G1511);
  nand (G1621,G1432,G1512);
  nand (G1622,G1434,G1513);
  nand (G1623,G1436,G1514);
  nand (G1624,G1438,G1515);
  nand (G1625,G1440,G1516);
  nand (G1626,G1442,G1517);
  nand (G1627,G1444,G1518);
  nand (G1628,G1446,G1519);
  nand (G1629,G1455,G1531);
  nand (G1630,G1457,G1532);
  nand (G1631,G1459,G1533);
  nand (G1632,G1461,G1534);
  nand (G1633,G1463,G1535);
  nand (G1634,G1465,G1536);
  nand (G1635,G1216,G1555);
  not (G1636,G1472);
  and (G1640,G1176,G1488);
  and (G1641,G1062,G1488);
  and (G1642,G1067,G1488);
  and (G1643,G1187,G1488);
  and (G1644,G1152,G1493);
  and (G1645,G1159,G1493);
  nand (G1646,G1599,G1600);
  not (G1650,G1537);
  nand (G1651,G1537,G1477);
  nand (G1652,G1540,G1478);
  not (G1653,G1540);
  not (G1654,G1479);
  nand (G1657,G1601,G1602);
  not (G1661,G1557);
  nand (G1662,G1557,G1485);
  not (G1663,G1575);
  and (G1664,G1152,G1498);
  and (G1665,G1159,G1498);
  and (G1666,G1176,G1502);
  and (G1667,G1062,G1502);
  and (G1668,G1067,G1502);
  and (G1669,G1187,G1502);
  not (G1670,G1493);
  not (G1675,G1578);
  not (G1676,G1498);
  nand (G1681,G1606,G1507);
  not (G1682,G1581);
  not (G1683,G1584);
  not (G1684,G1472);
  not (G1688,G1587);
  nand (G1689,G1587,G1427);
  not (G1690,G1628);
  not (G1691,G1627);
  not (G1692,G1626);
  not (G1693,G1625);
  not (G1694,G1624);
  not (G1695,G1623);
  not (G1696,G1622);
  not (G1697,G1621);
  not (G1698,G1620);
  not (G1699,G1619);
  not (G1700,G1634);
  not (G1701,G1633);
  not (G1702,G1632);
  not (G1703,G1631);
  not (G1704,G1630);
  not (G1705,G1629);
  not (G1706,G1520);
  not (G1709,G1524);
  not (G1712,G1528);
  not (G1715,G1528);
  not (G1718,G1596);
  nand (G1719,G1596,G1110);
  not (G1720,G1543);
  not (G1721,G1546);
  not (G1722,G1549);
  not (G1723,G1552);
  not (G1724,G1560);
  not (G1725,G1563);
  not (G1726,G1566);
  not (G1727,G1569);
  nand (G1728,G1635,G1556);
  not (G1731,G1572);
  not (G1732,G1590);
  not (G1733,G1593);
  and (G1734,G1421,G1610);
  and (G1735,G1418,G1607);
  nand (G1736,G1374,G1650);
  nand (G1737,G1377,G1653);
  nand (G1738,G1390,G1661);
  not (G1739,G1613);
  not (G1744,G1613);
  not (G1749,G1681);
  nand (G1750,G1263,G1688);
  and (G1751,G1690,G1691,G1692,G1693,G1694);
  and (G1752,G1695,G1696,G1697,G1698,G1699);
  and (G1753,G1255,G1700);
  and (G1754,G1701,G1702,G1703,G1704,G1705);
  nand (G1755,G990,G1718);
  not (G1756,G1616);
  not (G1761,G1616);
  nand (G1766,G1546,G1720);
  nand (G1767,G1543,G1721);
  nand (G1768,G1552,G1722);
  nand (G1769,G1549,G1723);
  nand (G1770,G1563,G1724);
  nand (G1771,G1560,G1725);
  nand (G1772,G1569,G1726);
  nand (G1773,G1566,G1727);
  nand (G1774,G1593,G1732);
  nand (G1775,G1590,G1733);
  or (G1776,G1734,G1610);
  or (G1777,G1735,G1607);
  and (G1778,G1152,G1670);
  and (G1779,G1159,G1670);
  and (G1780,G1166,G1670);
  and (G1781,G1171,G1670);
  not (G1782,G1646);
  nand (G1785,G1736,G1651);
  nand (G1789,G1652,G1737);
  not (G1792,G1657);
  nand (G1795,G1738,G1662);
  and (G1798,G1152,G1676);
  and (G1799,G1159,G1676);
  and (G1800,G1166,G1676);
  and (G1801,G1171,G1676);
  and (G1802,G1749,G10);
  not (G1805,G1636);
  nand (G1811,G1750,G1689);
  and (G1814,G1751,G1752);
  and (G1815,G1753,G1754);
  not (G1816,G1684);
  not (G1822,G1712);
  not (G1823,G1715);
  and (G1824,G1524,G1520,G1712);
  and (G1825,G1709,G1706,G1715);
  nand (G1826,G1755,G1719);
  not (G1829,G1636);
  not (G1835,G1636);
  not (G1840,G1684);
  not (G1846,G1684);
  nand (G1851,G1768,G1769);
  nand (G1854,G1766,G1767);
  not (G1857,G1728);
  nand (G1858,G1728,G1731);
  nand (G1859,G1772,G1773);
  nand (G1862,G1770,G1771);
  nand (G1865,G1774,G1775);
  and (G1868,G1640,G1739);
  and (G1869,G1641,G1739);
  and (G1870,G1642,G1739);
  and (G1871,G1643,G1739);
  or (G1872,G1778,G1644);
  or (G1873,G1779,G1645);
  and (G1874,G1780,G598);
  and (G1875,G1781,G598);
  or (G1876,G1798,G1664);
  or (G1877,G1799,G1665);
  and (G1878,G1800,G631);
  and (G1879,G1801,G631);
  and (G1880,G1666,G1744);
  and (G1881,G1667,G1744);
  and (G1882,G1668,G1744);
  and (G1883,G1669,G1744);
  and (G1884,G1814,G1815,G832);
  and (G1887,G1706,G1524,G1822);
  and (G1888,G1520,G1709,G1823);
  nand (G1889,G1572,G1857);
  not (G1890,G1868);
  not (G1893,G1869);
  not (G1896,G1870);
  not (G1899,G1871);
  and (G1902,G1872,G598);
  and (G1903,G1873,G598);
  not (G1904,G1874);
  not (G1907,G1875);
  not (G1910,G1785);
  not (G1913,G1789);
  not (G1916,G1789);
  not (G1919,G1795);
  not (G1922,G1795);
  and (G1925,G366,G1805);
  and (G1926,G1876,G631);
  and (G1927,G1877,G631);
  not (G1928,G1878);
  not (G1931,G1879);
  not (G1934,G1880);
  not (G1937,G1881);
  not (G1940,G1882);
  not (G1943,G1883);
  not (G1946,G1802);
  and (G1947,G366,G1816);
  not (G1948,G1805);
  and (G1953,G370,G1805);
  and (G1954,G447,G1805);
  and (G1955,G451,G1805);
  not (G1956,G1816);
  and (G1961,G370,G1816);
  and (G1962,G447,G1816);
  and (G1963,G451,G1816);
  nor (G1964,G1887,G1824);
  nor (G1965,G1888,G1825);
  not (G1966,G1865);
  not (G1967,G1829);
  and (G1970,G455,G1829);
  and (G1971,G459,G1829);
  and (G1972,G463,G1829);
  and (G1973,G467,G1829);
  and (G1974,G471,G1835);
  and (G1975,G475,G1835);
  and (G1976,G479,G1835);
  and (G1977,G497,G1835);
  not (G1978,G1840);
  and (G1981,G455,G1840);
  and (G1982,G459,G1840);
  and (G1983,G463,G1840);
  and (G1984,G467,G1840);
  and (G1985,G471,G1846);
  and (G1986,G475,G1846);
  and (G1987,G479,G1846);
  and (G1988,G497,G1846);
  not (G1989,G1851);
  not (G1990,G1854);
  not (G1991,G1859);
  not (G1992,G1862);
  nand (G1993,G1858,G1889);
  not (G1996,G1902);
  not (G1999,G1903);
  not (G2002,G1926);
  not (G2005,G1927);
  and (G2008,G1972,G751);
  and (G2011,G1973,G751);
  and (G2014,G1974,G1756);
  and (G2017,G1975,G1756);
  and (G2020,G1976,G1756);
  and (G2023,G1977,G1756);
  and (G2026,G1983,G756);
  and (G2029,G1984,G756);
  and (G2032,G1985,G1761);
  and (G2035,G1986,G1761);
  and (G2038,G1987,G1761);
  and (G2041,G1988,G1761);
  nand (G2044,G1854,G1989);
  nand (G2045,G1851,G1990);
  nand (G2046,G1862,G1991);
  nand (G2047,G1859,G1992);
  nand (G2048,G1965,G1964);
  not (G2051,G1913);
  not (G2052,G1916);
  not (G2053,G1919);
  not (G2054,G1922);
  and (G2055,G1785,G1646,G1913);
  and (G2056,G1910,G1782,G1916);
  and (G2057,G1657,G1479,G1919);
  and (G2058,G1792,G1654,G1922);
  nand (G2059,G1993,G1486);
  not (G2060,G1993);
  and (G2061,G479,G1948);
  and (G2062,G479,G1956);
  and (G2063,G497,G1948);
  and (G2064,G503,G1948);
  and (G2065,G507,G1948);
  and (G2066,G497,G1956);
  and (G2067,G503,G1956);
  and (G2068,G507,G1956);
  and (G2069,G511,G1967);
  and (G2070,G515,G1967);
  and (G2071,G511,G1978);
  and (G2072,G515,G1978);
  nand (G2073,G2044,G2045);
  nand (G2076,G2046,G2047);
  not (G2079,G1899);
  not (G2082,G1896);
  not (G2085,G1893);
  not (G2088,G1890);
  not (G2091,G1907);
  not (G2094,G1904);
  not (G2097,G1943);
  not (G2100,G1940);
  not (G2103,G1937);
  not (G2106,G1934);
  not (G2109,G1931);
  not (G2112,G1928);
  and (G2115,G1782,G1785,G2051);
  and (G2116,G1646,G1910,G2052);
  and (G2117,G1654,G1657,G2053);
  and (G2118,G1479,G1792,G2054);
  nand (G2119,G1393,G2060);
  or (G2120,G2061,G1925);
  nand (G2121,G2048,G1966);
  and (G2122,G2023,G1899);
  and (G2123,G2020,G1896);
  and (G2124,G2017,G1893);
  and (G2125,G1890,G2014);
  and (G2126,G2011,G1907);
  and (G2127,G2008,G1904);
  or (G2128,G2062,G1947);
  and (G2129,G2041,G1943);
  and (G2130,G2038,G1940);
  and (G2131,G2035,G1937);
  and (G2132,G1934,G2032);
  and (G2133,G2029,G1931);
  and (G2134,G2026,G1928);
  or (G2135,G2063,G1953);
  or (G2138,G2064,G1954);
  or (G2141,G2065,G1955);
  or (G2144,G2066,G1961);
  or (G2147,G2067,G1962);
  or (G2150,G2068,G1963);
  not (G2153,G2048);
  or (G2154,G2069,G1970);
  or (G2155,G2070,G1971);
  or (G2156,G2071,G1981);
  or (G2157,G2072,G1982);
  not (G2158,G2023);
  not (G2161,G2020);
  not (G2164,G2017);
  not (G2167,G2014);
  not (G2170,G2011);
  not (G2173,G2008);
  not (G2176,G1999);
  not (G2179,G1996);
  not (G2182,G2041);
  not (G2185,G2038);
  not (G2188,G2035);
  not (G2191,G2032);
  not (G2194,G2029);
  not (G2197,G2026);
  not (G2200,G2005);
  not (G2203,G2002);
  nand (G2206,G2059,G2119);
  nor (G2207,G2115,G2055);
  nor (G2208,G2116,G2056);
  nor (G2209,G2117,G2057);
  nor (G2210,G2118,G2058);
  not (G2211,G2073);
  not (G2212,G2076);
  and (G2213,G2120,G1132);
  nand (G2214,G1865,G2153);
  not (G2215,G2079);
  not (G2216,G2082);
  not (G2217,G2085);
  not (G2218,G2088);
  not (G2219,G2091);
  not (G2220,G2094);
  and (G2221,G2128,G1132);
  not (G2222,G2097);
  not (G2223,G2100);
  not (G2224,G2103);
  not (G2225,G2106);
  not (G2226,G2109);
  not (G2227,G2112);
  and (G2228,G2154,G751);
  and (G2231,G2155,G751);
  and (G2234,G2156,G756);
  and (G2237,G2157,G756);
  and (G2240,G2206,G325);
  and (G2241,G2138,G1329);
  and (G2242,G2135,G1137);
  nand (G2243,G2214,G2121);
  not (G2244,G2158);
  nand (G2245,G2158,G2215);
  not (G2246,G2161);
  nand (G2247,G2161,G2216);
  not (G2248,G2164);
  nand (G2249,G2164,G2217);
  not (G2250,G2167);
  nand (G2251,G2167,G2218);
  not (G2252,G2170);
  nand (G2253,G2170,G2219);
  not (G2254,G2173);
  nand (G2255,G2173,G2220);
  not (G2256,G2176);
  not (G2257,G2179);
  and (G2258,G2141,G1336);
  and (G2259,G2147,G1329);
  and (G2260,G2144,G1137);
  not (G2261,G2182);
  nand (G2262,G2182,G2222);
  not (G2263,G2185);
  nand (G2264,G2185,G2223);
  not (G2265,G2188);
  nand (G2266,G2188,G2224);
  not (G2267,G2191);
  nand (G2268,G2191,G2225);
  not (G2269,G2194);
  nand (G2270,G2194,G2226);
  not (G2271,G2197);
  nand (G2272,G2197,G2227);
  not (G2273,G2200);
  not (G2274,G2203);
  and (G2275,G2150,G1336);
  nand (G2276,G2208,G2207);
  nand (G2279,G2210,G2209);
  not (G2282,G2138);
  not (G2285,G2135);
  not (G2288,G2141);
  not (G2291,G2147);
  not (G2294,G2144);
  not (G2297,G2150);
  not (G2300,G2243);
  nand (G2301,G2079,G2244);
  nand (G2302,G2082,G2246);
  nand (G2303,G2085,G2248);
  nand (G2304,G2088,G2250);
  nand (G2305,G2091,G2252);
  nand (G2306,G2094,G2254);
  and (G2307,G2231,G1999);
  and (G2308,G2228,G1996);
  nand (G2309,G2097,G2261);
  nand (G2310,G2100,G2263);
  nand (G2311,G2103,G2265);
  nand (G2312,G2106,G2267);
  nand (G2313,G2109,G2269);
  nand (G2314,G2112,G2271);
  and (G2315,G2237,G2005);
  and (G2316,G2234,G2002);
  not (G2317,G2231);
  not (G2320,G2228);
  not (G2323,G2237);
  not (G2326,G2234);
  not (G2329,G2276);
  nand (G2330,G2276,G2211);
  not (G2331,G2279);
  nand (G2332,G2279,G2212);
  not (G2333,G2282);
  nand (G2334,G2282,G1663);
  nand (G2335,G2285,G1487);
  not (G2336,G2285);
  and (G2337,G2300,G581);
  nand (G2340,G2301,G2245);
  nand (G2345,G2302,G2247);
  nand (G2349,G2303,G2249);
  nand (G2352,G2304,G2251);
  nand (G2353,G2305,G2253);
  nand (G2359,G2306,G2255);
  not (G2364,G2288);
  nand (G2365,G2288,G1675);
  not (G2366,G2291);
  nand (G2367,G2291,G1682);
  nand (G2368,G2294,G1508);
  not (G2369,G2294);
  nand (G2370,G2309,G2262);
  nand (G2375,G2310,G2264);
  nand (G2379,G2311,G2266);
  nand (G2382,G2312,G2268);
  nand (G2383,G2313,G2270);
  nand (G2389,G2314,G2272);
  not (G2394,G2297);
  nand (G2395,G2297,G1683);
  nand (G2396,G2073,G2329);
  nand (G2397,G2076,G2331);
  nand (G2398,G1575,G2333);
  nand (G2399,G1396,G2336);
  not (G2400,G2317);
  nand (G2401,G2317,G2256);
  not (G2402,G2320);
  nand (G2403,G2320,G2257);
  nand (G2404,G1578,G2364);
  nand (G2405,G1581,G2366);
  nand (G2406,G1399,G2369);
  not (G2407,G2323);
  nand (G2408,G2323,G2273);
  not (G2409,G2326);
  nand (G2410,G2326,G2274);
  nand (G2411,G1584,G2394);
  nand (G2412,G2396,G2330);
  nand (G2413,G2397,G2332);
  nand (G2414,G2398,G2334);
  nand (G2417,G2399,G2335);
  not (G2418,G2337);
  nand (G2419,G2176,G2400);
  nand (G2420,G2179,G2402);
  nand (G2421,G2404,G2365);
  and (G2422,G2345,G2352,G2349,G2340);
  and (G2423,G2340,G2123);
  and (G2424,G2345,G2340,G2124);
  and (G2425,G2349,G2340,G2125,G2345);
  and (G2426,G2353,G2127);
  and (G2427,G2359,G2353,G2307);
  nand (G2428,G2405,G2367);
  nand (G2431,G2406,G2368);
  nand (G2432,G2200,G2407);
  nand (G2433,G2203,G2409);
  nand (G2434,G2411,G2395);
  and (G2435,G2375,G2382,G2379,G2370);
  and (G2436,G2370,G2130);
  and (G2437,G2375,G2370,G2131);
  and (G2438,G2379,G2370,G2132,G2375);
  and (G2439,G2383,G2134);
  and (G2440,G2389,G2383,G2315);
  not (G2441,G2412);
  and (G2442,G2413,G123);
  nand (G2443,G2419,G2401);
  nand (G2447,G2420,G2403);
  not (G2450,G2422);
  or (G2451,G2122,G2423,G2424,G2425);
  nand (G2454,G2432,G2408);
  nand (G2458,G2433,G2410);
  not (G2461,G2435);
  or (G2462,G2129,G2436,G2437,G2438);
  and (G2465,G2414,G2242);
  and (G2466,G2417,G2414,G2213);
  or (G2467,G1326,G2442);
  and (G2470,G2441,G581);
  and (G2473,G2428,G2260);
  and (G2474,G2431,G2428,G2221);
  or (G2475,G2241,G2465,G2466);
  not (G2476,G2451);
  and (G2477,G2359,G2421,G2443,G2353,G2447);
  and (G2478,G2443,G2353,G2308,G2359);
  and (G2479,G2447,G2443,G2353,G2258,G2359);
  or (G2480,G2259,G2473,G2474);
  not (G2481,G2462);
  and (G2482,G2389,G2434,G2454,G2383,G2458);
  and (G2483,G2454,G2383,G2316,G2389);
  and (G2484,G2458,G2454,G2383,G2275,G2389);
  or (G2485,G2126,G2426,G2427,G2478,G2479);
  and (G2486,G2477,G2475);
  nand (G2487,G2476,G2450);
  not (G2488,G2470);
  or (G2489,G2133,G2439,G2440,G2483,G2484);
  and (G2490,G2482,G2480);
  nand (G2491,G2481,G2461);
  or (G2492,G2485,G2486);
  and (G2495,G2418,G2488,G1826);
  or (G2496,G2489,G2490);
  not (G2499,G2492);
  and (G2500,G2487,G2492);
  not (G2501,G2496);
  and (G2502,G2491,G2496);
  and (G2503,G2451,G2499);
  and (G2504,G2462,G2501);
  or (G2505,G2503,G2500);
  or (G2508,G2504,G2502);
  nand (G2512,G2508,G2505);
  and (G2515,G2508,G2512);
  and (G2516,G2512,G2505);
  or (G2517,G2515,G2516);
  not (G2520,G2517);
  and (G2523,G2517,G2520);
  or (G2524,G2523,G2520);
  and (G2527,G1811,G1946,G2524);
  and (G2528,G2495,G2527,G993);
  not (G2531,G115);
  not (G2532,G115);
  not (G2533,G115);
  not (G2534,G124);
  not (G2535,G124);
  not (G2536,G137);
  not (G2537,G137);
  not (G2538,G137);
  not (G2539,G32);
  not (G2540,G106);
  not (G2541,G64);
  not (G2542,G76);
  not (G2543,G53);
  not (G2544,G96);
  not (G2545,G43);
  not (G2546,G86);
  not (G2547,G285);
  not (G2548,G287);
  not (G2549,G292);
  and (G2550,G74,G292);
  not (G2551,G443);
  nand (G2552,G119,G443);
  not (G2553,G592);
  not (G2554,G595);
  not (G2555,G595);
  not (G2556,G993);
  not (G2557,G1044);
  not (G2558,G1049);
  not (G2559,G1039);
  not (G2560,G1026);
  not (G2561,G1021);
  not (G2562,G1017);
  or (G2563,G325,G1117);
  not (G2564,G1118);
  not (G2565,G1119);
  not (G2566,G1144);
  not (G2567,G1148);
  not (G2568,G1152);
  not (G2569,G1159);
  not (G2570,G1166);
  not (G2571,G1171);
  not (G2572,G1176);
  not (G2573,G1412);
  not (G2574,G1412);
  not (G2575,G1415);
  not (G2576,G1415);
  or (G2577,G1471,G1116);
  not (G2578,G1603);
  not (G2579,G1603);
  nand (G2580,G1776,G1777);
  not (G2581,G1802);
  not (G2582,G1826);
  not (G2583,G1811);
  not (G2584,G1884);
  not (G2585,G1884);
  or (G2586,G2240,G1115);
  not (G2587,G2337);
  not (G2588,G2467);
  not (G2589,G2467);
  not (G2590,G2470);
  not (G2591,G2508);
  not (G2592,G2524);
  not (G2593,G2528);
  not (G2594,G2528);

endmodule
