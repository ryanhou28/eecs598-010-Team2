

module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G426,
  G427,
  G428,
  G429,
  G430,
  G431,
  G432
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;
  output G426;output G427;output G428;output G429;output G430;output G431;output G432;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire g37_p;
  wire g37_n;
  wire g38_p;
  wire g38_n;
  wire g39_p;
  wire g39_n;
  wire g40_p;
  wire g40_n;
  wire g41_p;
  wire g41_n;
  wire g42_p;
  wire g42_n;
  wire g43_p;
  wire g43_n;
  wire g44_p;
  wire g44_n;
  wire g45_p;
  wire g45_n;
  wire g46_p;
  wire g46_n;
  wire g47_p;
  wire g47_n;
  wire g48_p;
  wire g48_n;
  wire g49_p;
  wire g49_n;
  wire g50_p;
  wire g50_n;
  wire g51_p;
  wire g51_n;
  wire g52_p;
  wire g52_n;
  wire g53_p;
  wire g53_n;
  wire g54_p;
  wire g54_n;
  wire g55_p;
  wire g55_n;
  wire g56_p;
  wire g56_n;
  wire g57_p;
  wire g57_n;
  wire g58_p;
  wire g58_n;
  wire g59_p;
  wire g59_n;
  wire g60_p;
  wire g60_n;
  wire g61_p;
  wire g61_n;
  wire g62_p;
  wire g62_n;
  wire g63_p;
  wire g63_n;
  wire g64_p;
  wire g64_n;
  wire g65_p;
  wire g65_n;
  wire g66_p;
  wire g66_n;
  wire g67_p;
  wire g67_n;
  wire g68_p;
  wire g68_n;
  wire g69_p;
  wire g69_n;
  wire g70_p;
  wire g70_n;
  wire g71_p;
  wire g71_n;
  wire g72_p;
  wire g72_n;
  wire g73_p;
  wire g73_n;
  wire g74_p;
  wire g74_n;
  wire g75_p;
  wire g75_n;
  wire g76_p;
  wire g76_n;
  wire g77_p;
  wire g77_n;
  wire g78_p;
  wire g78_n;
  wire g79_p;
  wire g79_n;
  wire g80_p;
  wire g80_n;
  wire g81_p;
  wire g81_n;
  wire g82_p;
  wire g82_n;
  wire g83_p;
  wire g83_n;
  wire g84_p;
  wire g84_n;
  wire g85_p;
  wire g85_n;
  wire g86_p;
  wire g86_n;
  wire g87_p;
  wire g87_n;
  wire g88_p;
  wire g88_n;
  wire g89_p;
  wire g89_n;
  wire g90_p;
  wire g90_n;
  wire g91_p;
  wire g91_n;
  wire g92_p;
  wire g92_n;
  wire g93_p;
  wire g93_n;
  wire g94_p;
  wire g94_n;
  wire g95_p;
  wire g95_n;
  wire g96_p;
  wire g96_n;
  wire g97_p;
  wire g97_n;
  wire g98_p;
  wire g98_n;
  wire g99_p;
  wire g99_n;
  wire g100_p;
  wire g100_n;
  wire g101_p;
  wire g101_n;
  wire g102_p;
  wire g102_n;
  wire g103_p;
  wire g103_n;
  wire g104_p;
  wire g104_n;
  wire g105_p;
  wire g105_n;
  wire g106_p;
  wire g106_n;
  wire g107_p;
  wire g107_n;
  wire g108_p;
  wire g108_n;
  wire g109_p;
  wire g109_n;
  wire g110_p;
  wire g110_n;
  wire g111_p;
  wire g111_n;
  wire g112_p;
  wire g112_n;
  wire g113_p;
  wire g113_n;
  wire g114_p;
  wire g114_n;
  wire g115_p;
  wire g115_n;
  wire g116_p;
  wire g116_n;
  wire g117_p;
  wire g117_n;
  wire g118_p;
  wire g118_n;
  wire g119_p;
  wire g119_n;
  wire g120_p;
  wire g120_n;
  wire g121_p;
  wire g121_n;
  wire g122_p;
  wire g122_n;
  wire g123_p;
  wire g123_n;
  wire g124_p;
  wire g124_n;
  wire g125_p;
  wire g125_n;
  wire g126_p;
  wire g126_n;
  wire g127_p;
  wire g127_n;
  wire g128_p;
  wire g128_n;
  wire g129_p;
  wire g129_n;
  wire g130_p;
  wire g130_n;
  wire g131_p;
  wire g131_n;
  wire g132_p;
  wire g132_n;
  wire g133_p;
  wire g133_n;
  wire g134_p;
  wire g134_n;
  wire g135_p;
  wire g135_n;
  wire g136_p;
  wire g136_n;
  wire g137_p;
  wire g137_n;
  wire g138_p;
  wire g138_n;
  wire g139_p;
  wire g139_n;
  wire g140_p;
  wire g140_n;
  wire g141_p;
  wire g141_n;
  wire g142_p;
  wire g142_n;
  wire g143_p;
  wire g143_n;
  wire g144_p;
  wire g144_n;
  wire g145_p;
  wire g145_n;
  wire g146_p;
  wire g146_n;
  wire g147_p;
  wire g147_n;
  wire g148_p;
  wire g148_n;
  wire g149_p;
  wire g149_n;
  wire g150_p;
  wire g150_n;
  wire g151_p;
  wire g151_n;
  wire g152_p;
  wire g152_n;
  wire g153_p;
  wire g153_n;
  wire g154_p;
  wire g154_n;
  wire g155_p;
  wire g155_n;
  wire g156_p;
  wire g156_n;
  wire g157_p;
  wire g157_n;
  wire g158_p;
  wire g158_n;
  wire g159_p;
  wire g159_n;

wire G1_spl_, G2_spl_, G3_spl_, G4_spl_, G5_spl_, G6_spl_, G7_spl_, G8_spl_, G9_spl_, G10_spl_, G11_spl_, G12_spl_, G13_spl_, G14_spl_, G15_spl_, G16_spl_, G17_spl_, G18_spl_, G19_spl_, G20_spl_, G21_spl_, G22_spl_, G23_spl_, G24_spl_, G25_spl_, G26_spl_, G27_spl_, G28_spl_, G29_spl_, G30_spl_, G31_spl_, G32_spl_, G33_spl_, G34_spl_, G35_spl_, G36_spl_, G10_p_spl_, G8_n_spl_, G10_n_spl_, G8_p_spl_, G6_p_spl_, G4_n_spl_, G6_n_spl_, G4_p_spl_, G26_p_spl_, G24_n_spl_, G26_n_spl_, G24_p_spl_, G18_p_spl_, G16_n_spl_, G18_n_spl_, G16_p_spl_, G14_p_spl_, G12_n_spl_, G14_n_spl_, G12_p_spl_, G30_p_spl_, G28_n_spl_, G30_n_spl_, G28_p_spl_, G2_p_spl_, G1_n_spl_, G2_n_spl_, G1_p_spl_, G22_p_spl_, G20_n_spl_, G22_n_spl_, G20_p_spl_, G34_p_spl_, G32_n_spl_, G34_n_spl_, G32_p_spl_, g53_n_spl_, g53_n_spl_0, g53_n_spl_00, g53_n_spl_000, g53_n_spl_001, g53_n_spl_01, g53_n_spl_1, g53_n_spl_10, g53_n_spl_11, g53_p_spl_, g53_p_spl_0, g53_p_spl_00, g53_p_spl_000, g53_p_spl_01, g53_p_spl_1, g53_p_spl_10, g53_p_spl_11, g55_p_spl_, G27_n_spl_, g55_n_spl_, G27_p_spl_, g58_p_spl_, G31_n_spl_, g58_n_spl_, G31_p_spl_, g61_p_spl_, G19_n_spl_, g61_n_spl_, G19_p_spl_, g66_p_spl_, G11_n_spl_, g66_n_spl_, G11_p_spl_, g69_p_spl_, G35_n_spl_, g69_n_spl_, G35_p_spl_, g73_p_spl_, G23_n_spl_, g73_n_spl_, G23_p_spl_, g76_p_spl_, G7_n_spl_, g76_n_spl_, G7_p_spl_, g80_p_spl_, G3_n_spl_, g80_n_spl_, G3_p_spl_, g83_p_spl_, G15_n_spl_, g83_n_spl_, G15_p_spl_, g88_n_spl_, g88_n_spl_0, g88_n_spl_00, g88_n_spl_000, g88_n_spl_001, g88_n_spl_01, g88_n_spl_1, g88_n_spl_10, g88_n_spl_11, g88_p_spl_, g88_p_spl_0, g88_p_spl_00, g88_p_spl_000, g88_p_spl_01, g88_p_spl_1, g88_p_spl_10, g88_p_spl_11, g90_p_spl_, G29_n_spl_, g90_n_spl_, G29_p_spl_, g93_n_spl_, G33_p_spl_, g96_p_spl_, G21_n_spl_, g96_n_spl_, G21_p_spl_, g101_p_spl_, G13_n_spl_, g101_n_spl_, G13_p_spl_, g104_n_spl_, G36_p_spl_, g108_n_spl_, G25_p_spl_, g111_n_spl_, G9_p_spl_, g115_p_spl_, G5_n_spl_, g118_p_spl_, G17_n_spl_, g118_n_spl_, G17_p_spl_, g123_p_spl_, g123_p_spl_0, g123_p_spl_00, g123_p_spl_1, g123_n_spl_, g123_n_spl_0, g123_n_spl_00, g123_n_spl_000, g123_n_spl_01, g123_n_spl_1, g123_n_spl_10, g123_n_spl_11, g127_n_spl_, g134_n_spl_, g130_p_spl_, g140_n_spl_, g145_n_spl_, g143_n_spl_, g136_p_spl_, g129_p_spl_, g135_n_spl_, g151_n_spl_;

buf (G1_p, G1_spl_);
not (G1_n, G1_spl_);
buf (G2_p, G2_spl_);
not (G2_n, G2_spl_);
buf (G3_p, G3_spl_);
not (G3_n, G3_spl_);
buf (G4_p, G4_spl_);
not (G4_n, G4_spl_);
buf (G5_p, G5_spl_);
not (G5_n, G5_spl_);
buf (G6_p, G6_spl_);
not (G6_n, G6_spl_);
buf (G7_p, G7_spl_);
not (G7_n, G7_spl_);
buf (G8_p, G8_spl_);
not (G8_n, G8_spl_);
buf (G9_p, G9_spl_);
not (G9_n, G9_spl_);
buf (G10_p, G10_spl_);
not (G10_n, G10_spl_);
buf (G11_p, G11_spl_);
not (G11_n, G11_spl_);
buf (G12_p, G12_spl_);
not (G12_n, G12_spl_);
buf (G13_p, G13_spl_);
not (G13_n, G13_spl_);
buf (G14_p, G14_spl_);
not (G14_n, G14_spl_);
buf (G15_p, G15_spl_);
not (G15_n, G15_spl_);
buf (G16_p, G16_spl_);
not (G16_n, G16_spl_);
buf (G17_p, G17_spl_);
not (G17_n, G17_spl_);
buf (G18_p, G18_spl_);
not (G18_n, G18_spl_);
buf (G19_p, G19_spl_);
not (G19_n, G19_spl_);
buf (G20_p, G20_spl_);
not (G20_n, G20_spl_);
buf (G21_p, G21_spl_);
not (G21_n, G21_spl_);
buf (G22_p, G22_spl_);
not (G22_n, G22_spl_);
buf (G23_p, G23_spl_);
not (G23_n, G23_spl_);
buf (G24_p, G24_spl_);
not (G24_n, G24_spl_);
buf (G25_p, G25_spl_);
not (G25_n, G25_spl_);
buf (G26_p, G26_spl_);
not (G26_n, G26_spl_);
buf (G27_p, G27_spl_);
not (G27_n, G27_spl_);
buf (G28_p, G28_spl_);
not (G28_n, G28_spl_);
buf (G29_p, G29_spl_);
not (G29_n, G29_spl_);
buf (G30_p, G30_spl_);
not (G30_n, G30_spl_);
buf (G31_p, G31_spl_);
not (G31_n, G31_spl_);
buf (G32_p, G32_spl_);
not (G32_n, G32_spl_);
buf (G33_p, G33_spl_);
not (G33_n, G33_spl_);
buf (G34_p, G34_spl_);
not (G34_n, G34_spl_);
buf (G35_p, G35_spl_);
not (G35_n, G35_spl_);
buf (G36_p, G36_spl_);
not (G36_n, G36_spl_);
and (g37_p, G10_p_spl_, G8_n_spl_);
or (g37_n, G10_n_spl_, G8_p_spl_);
and (g38_p, G6_p_spl_, G4_n_spl_);
or (g38_n, G6_n_spl_, G4_p_spl_);
and (g39_p, G26_p_spl_, G24_n_spl_);
or (g39_n, G26_n_spl_, G24_p_spl_);
and (g40_p, g39_n, g38_n);
or (g40_n, g39_p, g38_p);
and (g41_p, g40_p, g37_n);
or (g41_n, g40_n, g37_p);
and (g42_p, G18_p_spl_, G16_n_spl_);
or (g42_n, G18_n_spl_, G16_p_spl_);
and (g43_p, G14_p_spl_, G12_n_spl_);
or (g43_n, G14_n_spl_, G12_p_spl_);
and (g44_p, g43_n, g42_n);
or (g44_n, g43_p, g42_p);
and (g45_p, G30_p_spl_, G28_n_spl_);
or (g45_n, G30_n_spl_, G28_p_spl_);
and (g46_p, G2_p_spl_, G1_n_spl_);
or (g46_n, G2_n_spl_, G1_p_spl_);
and (g47_p, g46_n, g45_n);
or (g47_n, g46_p, g45_p);
and (g48_p, G22_p_spl_, G20_n_spl_);
or (g48_n, G22_n_spl_, G20_p_spl_);
and (g49_p, G34_p_spl_, G32_n_spl_);
or (g49_n, G34_n_spl_, G32_p_spl_);
and (g50_p, g49_n, g48_n);
or (g50_n, g49_p, g48_p);
and (g51_p, g50_p, g47_p);
or (g51_n, g50_n, g47_n);
and (g52_p, g51_p, g44_p);
or (g52_n, g51_n, g44_n);
and (g53_p, g52_p, g41_p);
or (g53_n, g52_n, g41_n);
and (g54_p, g53_n_spl_000, G24_p_spl_);
or (g54_n, g53_p_spl_000, G24_n_spl_);
and (g55_p, g54_n, G26_p_spl_);
or (g55_n, g54_p, G26_n_spl_);
and (g56_p, g55_p_spl_, G27_n_spl_);
or (g56_n, g55_n_spl_, G27_p_spl_);
and (g57_p, g53_n_spl_000, G28_p_spl_);
or (g57_n, g53_p_spl_000, G28_n_spl_);
and (g58_p, g57_n, G30_p_spl_);
or (g58_n, g57_p, G30_n_spl_);
and (g59_p, g58_p_spl_, G31_n_spl_);
or (g59_n, g58_n_spl_, G31_p_spl_);
and (g60_p, g53_n_spl_001, G16_p_spl_);
or (g60_n, g53_p_spl_00, G16_n_spl_);
and (g61_p, g60_n, G18_p_spl_);
or (g61_n, g60_p, G18_n_spl_);
and (g62_p, g61_p_spl_, G19_n_spl_);
or (g62_n, g61_n_spl_, G19_p_spl_);
and (g63_p, g62_n, g59_n);
or (g63_n, g62_p, g59_p);
and (g64_p, g63_p, g56_n);
or (g64_n, g63_n, g56_p);
and (g65_p, g53_n_spl_001, G8_p_spl_);
or (g65_n, g53_p_spl_01, G8_n_spl_);
and (g66_p, g65_n, G10_p_spl_);
or (g66_n, g65_p, G10_n_spl_);
and (g67_p, g66_p_spl_, G11_n_spl_);
or (g67_n, g66_n_spl_, G11_p_spl_);
and (g68_p, g53_n_spl_01, G32_p_spl_);
or (g68_n, g53_p_spl_01, G32_n_spl_);
and (g69_p, g68_n, G34_p_spl_);
or (g69_n, g68_p, G34_n_spl_);
and (g70_p, g69_p_spl_, G35_n_spl_);
or (g70_n, g69_n_spl_, G35_p_spl_);
and (g71_p, g70_n, g67_n);
or (g71_n, g70_p, g67_p);
and (g72_p, g53_n_spl_01, G20_p_spl_);
or (g72_n, g53_p_spl_10, G20_n_spl_);
and (g73_p, g72_n, G22_p_spl_);
or (g73_n, g72_p, G22_n_spl_);
and (g74_p, g73_p_spl_, G23_n_spl_);
or (g74_n, g73_n_spl_, G23_p_spl_);
and (g75_p, g53_n_spl_10, G4_p_spl_);
or (g75_n, g53_p_spl_10, G4_n_spl_);
and (g76_p, g75_n, G6_p_spl_);
or (g76_n, g75_p, G6_n_spl_);
and (g77_p, g76_p_spl_, G7_n_spl_);
or (g77_n, g76_n_spl_, G7_p_spl_);
and (g78_p, g77_n, g74_n);
or (g78_n, g77_p, g74_p);
and (g79_p, g53_n_spl_10, G1_p_spl_);
or (g79_n, g53_p_spl_11, G1_n_spl_);
and (g80_p, g79_n, G2_p_spl_);
or (g80_n, g79_p, G2_n_spl_);
and (g81_p, g80_p_spl_, G3_n_spl_);
or (g81_n, g80_n_spl_, G3_p_spl_);
and (g82_p, g53_n_spl_11, G12_p_spl_);
or (g82_n, g53_p_spl_11, G12_n_spl_);
and (g83_p, g82_n, G14_p_spl_);
or (g83_n, g82_p, G14_n_spl_);
and (g84_p, g83_p_spl_, G15_n_spl_);
or (g84_n, g83_n_spl_, G15_p_spl_);
and (g85_p, g84_n, g81_n);
or (g85_n, g84_p, g81_p);
and (g86_p, g85_p, g78_p);
or (g86_n, g85_n, g78_n);
and (g87_p, g86_p, g71_p);
or (g87_n, g86_n, g71_n);
and (g88_p, g87_p, g64_p);
or (g88_n, g87_n, g64_n);
and (g89_p, g88_n_spl_000, G27_p_spl_);
or (g89_n, g88_p_spl_000, G27_n_spl_);
and (g90_p, g89_n, g55_p_spl_);
or (g90_n, g89_p, g55_n_spl_);
and (g91_p, g90_p_spl_, G29_n_spl_);
or (g91_n, g90_n_spl_, G29_p_spl_);
and (g92_p, g88_n_spl_000, G31_p_spl_);
or (g92_n, g88_p_spl_000, G31_n_spl_);
and (g93_p, g92_n, g58_p_spl_);
or (g93_n, g92_p, g58_n_spl_);
and (g94_p, g93_p, G33_n);
or (g94_n, g93_n_spl_, G33_p_spl_);
and (g95_p, g88_n_spl_001, G19_p_spl_);
or (g95_n, g88_p_spl_00, G19_n_spl_);
and (g96_p, g95_n, g61_p_spl_);
or (g96_n, g95_p, g61_n_spl_);
and (g97_p, g96_p_spl_, G21_n_spl_);
or (g97_n, g96_n_spl_, G21_p_spl_);
and (g98_p, g97_n, g94_n);
or (g98_n, g97_p, g94_p);
and (g99_p, g98_p, g91_n);
or (g99_n, g98_n, g91_p);
and (g100_p, g88_n_spl_001, G11_p_spl_);
or (g100_n, g88_p_spl_01, G11_n_spl_);
and (g101_p, g100_n, g66_p_spl_);
or (g101_n, g100_p, g66_n_spl_);
and (g102_p, g101_p_spl_, G13_n_spl_);
or (g102_n, g101_n_spl_, G13_p_spl_);
and (g103_p, g88_n_spl_01, G35_p_spl_);
or (g103_n, g88_p_spl_01, G35_n_spl_);
and (g104_p, g103_n, g69_p_spl_);
or (g104_n, g103_p, g69_n_spl_);
and (g105_p, g104_p, G36_n);
or (g105_n, g104_n_spl_, G36_p_spl_);
and (g106_p, g105_n, g102_n);
or (g106_n, g105_p, g102_p);
and (g107_p, g88_n_spl_01, G23_p_spl_);
or (g107_n, g88_p_spl_10, G23_n_spl_);
and (g108_p, g107_n, g73_p_spl_);
or (g108_n, g107_p, g73_n_spl_);
and (g109_p, g108_p, G25_n);
or (g109_n, g108_n_spl_, G25_p_spl_);
and (g110_p, g88_n_spl_10, G7_p_spl_);
or (g110_n, g88_p_spl_10, G7_n_spl_);
and (g111_p, g110_n, g76_p_spl_);
or (g111_n, g110_p, g76_n_spl_);
and (g112_p, g111_p, G9_n);
or (g112_n, g111_n_spl_, G9_p_spl_);
and (g113_p, g112_n, g109_n);
or (g113_n, g112_p, g109_p);
and (g114_p, g88_n_spl_10, G3_p_spl_);
or (g114_n, g88_p_spl_11, G3_n_spl_);
and (g115_p, g114_n, g80_p_spl_);
or (g115_n, g114_p, g80_n_spl_);
and (g116_p, g115_p_spl_, G5_n_spl_);
or (g116_n, g115_n, G5_p);
and (g117_p, g88_n_spl_11, G15_p_spl_);
or (g117_n, g88_p_spl_11, G15_n_spl_);
and (g118_p, g117_n, g83_p_spl_);
or (g118_n, g117_p, g83_n_spl_);
and (g119_p, g118_p_spl_, G17_n_spl_);
or (g119_n, g118_n_spl_, G17_p_spl_);
and (g120_p, g119_n, g116_n);
or (g120_n, g119_p, g116_p);
and (g121_p, g120_p, g113_p);
or (g121_n, g120_n, g113_n);
and (g122_p, g121_p, g106_p);
or (g122_n, g121_n, g106_n);
and (g123_p, g122_p, g99_p);
or (g123_n, g122_n, g99_n);
or (g124_n, g123_p_spl_00, G5_n_spl_);
and (g125_p, g124_n, g115_p_spl_);
and (g126_p, g123_n_spl_000, G9_p_spl_);
or (g127_n, g126_p, g111_n_spl_);
and (g128_p, g123_n_spl_000, G13_p_spl_);
or (g128_n, g123_p_spl_00, G13_n_spl_);
and (g129_p, g128_n, g101_p_spl_);
or (g129_n, g128_p, g101_n_spl_);
and (g130_p, g129_n, g127_n_spl_);
and (g131_p, g123_n_spl_00, G21_p_spl_);
or (g131_n, g123_p_spl_0, G21_n_spl_);
and (g132_p, g131_n, g96_p_spl_);
or (g132_n, g131_p, g96_n_spl_);
and (g133_p, g123_n_spl_01, G17_p_spl_);
or (g133_n, g123_p_spl_1, G17_n_spl_);
and (g134_p, g133_n, g118_p_spl_);
or (g134_n, g133_p, g118_n_spl_);
and (g135_p, g134_n_spl_, g132_n);
or (g135_n, g134_p, g132_p);
and (g136_p, g135_p, g130_p_spl_);
and (g137_p, g123_n_spl_01, G36_p_spl_);
or (g138_n, g137_p, g104_n_spl_);
and (g139_p, g123_n_spl_10, G33_p_spl_);
or (g140_n, g139_p, g93_n_spl_);
and (g141_p, g140_n_spl_, g138_n);
and (g142_p, g123_n_spl_10, G29_p_spl_);
or (g142_n, g123_p_spl_1, G29_n_spl_);
and (g143_p, g142_n, g90_p_spl_);
or (g143_n, g142_p, g90_n_spl_);
and (g144_p, g123_n_spl_11, G25_p_spl_);
or (g145_n, g144_p, g108_n_spl_);
and (g146_p, g145_n_spl_, g143_n_spl_);
and (g147_p, g146_p, g141_p);
and (g148_p, g147_p, g136_p_spl_);
or (g149_n, g148_p, g125_p);
or (g150_n, g145_n_spl_, g129_p_spl_);
or (g151_n, g150_n, g135_n_spl_);
or (g152_n, g143_n_spl_, g135_n_spl_);
and (g153_p, g152_n, g130_p_spl_);
and (g154_p, g153_p, g151_n_spl_);
or (g155_n, g143_p, g140_n_spl_);
and (g156_p, g155_n, g134_n_spl_);
or (g157_n, g156_p, g129_p_spl_);
and (g158_p, g151_n_spl_, g127_n_spl_);
and (g159_p, g158_p, g157_n);
buf (G426, g53_n_spl_11);
buf (G427, g88_n_spl_11);
buf (G428, g123_n_spl_11);
not (G429, g149_n);
not (G430, g136_p_spl_);
not (G431, g154_p);
not (G432, g159_p);
/*splt*/ buf (G1_spl_, G1);
/*splt*/ buf (G2_spl_, G2);
/*splt*/ buf (G3_spl_, G3);
/*splt*/ buf (G4_spl_, G4);
/*splt*/ buf (G5_spl_, G5);
/*splt*/ buf (G6_spl_, G6);
/*splt*/ buf (G7_spl_, G7);
/*splt*/ buf (G8_spl_, G8);
/*splt*/ buf (G9_spl_, G9);
/*splt*/ buf (G10_spl_, G10);
/*splt*/ buf (G11_spl_, G11);
/*splt*/ buf (G12_spl_, G12);
/*splt*/ buf (G13_spl_, G13);
/*splt*/ buf (G14_spl_, G14);
/*splt*/ buf (G15_spl_, G15);
/*splt*/ buf (G16_spl_, G16);
/*splt*/ buf (G17_spl_, G17);
/*splt*/ buf (G18_spl_, G18);
/*splt*/ buf (G19_spl_, G19);
/*splt*/ buf (G20_spl_, G20);
/*splt*/ buf (G21_spl_, G21);
/*splt*/ buf (G22_spl_, G22);
/*splt*/ buf (G23_spl_, G23);
/*splt*/ buf (G24_spl_, G24);
/*splt*/ buf (G25_spl_, G25);
/*splt*/ buf (G26_spl_, G26);
/*splt*/ buf (G27_spl_, G27);
/*splt*/ buf (G28_spl_, G28);
/*splt*/ buf (G29_spl_, G29);
/*splt*/ buf (G30_spl_, G30);
/*splt*/ buf (G31_spl_, G31);
/*splt*/ buf (G32_spl_, G32);
/*splt*/ buf (G33_spl_, G33);
/*splt*/ buf (G34_spl_, G34);
/*splt*/ buf (G35_spl_, G35);
/*splt*/ buf (G36_spl_, G36);
/*splt*/ buf (G10_p_spl_, G10_p);
/*splt*/ buf (G8_n_spl_, G8_n);
/*splt*/ buf (G10_n_spl_, G10_n);
/*splt*/ buf (G8_p_spl_, G8_p);
/*splt*/ buf (G6_p_spl_, G6_p);
/*splt*/ buf (G4_n_spl_, G4_n);
/*splt*/ buf (G6_n_spl_, G6_n);
/*splt*/ buf (G4_p_spl_, G4_p);
/*splt*/ buf (G26_p_spl_, G26_p);
/*splt*/ buf (G24_n_spl_, G24_n);
/*splt*/ buf (G26_n_spl_, G26_n);
/*splt*/ buf (G24_p_spl_, G24_p);
/*splt*/ buf (G18_p_spl_, G18_p);
/*splt*/ buf (G16_n_spl_, G16_n);
/*splt*/ buf (G18_n_spl_, G18_n);
/*splt*/ buf (G16_p_spl_, G16_p);
/*splt*/ buf (G14_p_spl_, G14_p);
/*splt*/ buf (G12_n_spl_, G12_n);
/*splt*/ buf (G14_n_spl_, G14_n);
/*splt*/ buf (G12_p_spl_, G12_p);
/*splt*/ buf (G30_p_spl_, G30_p);
/*splt*/ buf (G28_n_spl_, G28_n);
/*splt*/ buf (G30_n_spl_, G30_n);
/*splt*/ buf (G28_p_spl_, G28_p);
/*splt*/ buf (G2_p_spl_, G2_p);
/*splt*/ buf (G1_n_spl_, G1_n);
/*splt*/ buf (G2_n_spl_, G2_n);
/*splt*/ buf (G1_p_spl_, G1_p);
/*splt*/ buf (G22_p_spl_, G22_p);
/*splt*/ buf (G20_n_spl_, G20_n);
/*splt*/ buf (G22_n_spl_, G22_n);
/*splt*/ buf (G20_p_spl_, G20_p);
/*splt*/ buf (G34_p_spl_, G34_p);
/*splt*/ buf (G32_n_spl_, G32_n);
/*splt*/ buf (G34_n_spl_, G34_n);
/*splt*/ buf (G32_p_spl_, G32_p);
/*splt*/ buf (g53_n_spl_, g53_n);
/*splt*/ buf (g53_n_spl_0, g53_n_spl_);
/*splt*/ buf (g53_n_spl_00, g53_n_spl_0);
/*splt*/ buf (g53_n_spl_000, g53_n_spl_00);
/*splt*/ buf (g53_n_spl_001, g53_n_spl_00);
/*splt*/ buf (g53_n_spl_01, g53_n_spl_0);
/*splt*/ buf (g53_n_spl_1, g53_n_spl_);
/*splt*/ buf (g53_n_spl_10, g53_n_spl_1);
/*splt*/ buf (g53_n_spl_11, g53_n_spl_1);
/*splt*/ buf (g53_p_spl_, g53_p);
/*splt*/ buf (g53_p_spl_0, g53_p_spl_);
/*splt*/ buf (g53_p_spl_00, g53_p_spl_0);
/*splt*/ buf (g53_p_spl_000, g53_p_spl_00);
/*splt*/ buf (g53_p_spl_01, g53_p_spl_0);
/*splt*/ buf (g53_p_spl_1, g53_p_spl_);
/*splt*/ buf (g53_p_spl_10, g53_p_spl_1);
/*splt*/ buf (g53_p_spl_11, g53_p_spl_1);
/*splt*/ buf (g55_p_spl_, g55_p);
/*splt*/ buf (G27_n_spl_, G27_n);
/*splt*/ buf (g55_n_spl_, g55_n);
/*splt*/ buf (G27_p_spl_, G27_p);
/*splt*/ buf (g58_p_spl_, g58_p);
/*splt*/ buf (G31_n_spl_, G31_n);
/*splt*/ buf (g58_n_spl_, g58_n);
/*splt*/ buf (G31_p_spl_, G31_p);
/*splt*/ buf (g61_p_spl_, g61_p);
/*splt*/ buf (G19_n_spl_, G19_n);
/*splt*/ buf (g61_n_spl_, g61_n);
/*splt*/ buf (G19_p_spl_, G19_p);
/*splt*/ buf (g66_p_spl_, g66_p);
/*splt*/ buf (G11_n_spl_, G11_n);
/*splt*/ buf (g66_n_spl_, g66_n);
/*splt*/ buf (G11_p_spl_, G11_p);
/*splt*/ buf (g69_p_spl_, g69_p);
/*splt*/ buf (G35_n_spl_, G35_n);
/*splt*/ buf (g69_n_spl_, g69_n);
/*splt*/ buf (G35_p_spl_, G35_p);
/*splt*/ buf (g73_p_spl_, g73_p);
/*splt*/ buf (G23_n_spl_, G23_n);
/*splt*/ buf (g73_n_spl_, g73_n);
/*splt*/ buf (G23_p_spl_, G23_p);
/*splt*/ buf (g76_p_spl_, g76_p);
/*splt*/ buf (G7_n_spl_, G7_n);
/*splt*/ buf (g76_n_spl_, g76_n);
/*splt*/ buf (G7_p_spl_, G7_p);
/*splt*/ buf (g80_p_spl_, g80_p);
/*splt*/ buf (G3_n_spl_, G3_n);
/*splt*/ buf (g80_n_spl_, g80_n);
/*splt*/ buf (G3_p_spl_, G3_p);
/*splt*/ buf (g83_p_spl_, g83_p);
/*splt*/ buf (G15_n_spl_, G15_n);
/*splt*/ buf (g83_n_spl_, g83_n);
/*splt*/ buf (G15_p_spl_, G15_p);
/*splt*/ buf (g88_n_spl_, g88_n);
/*splt*/ buf (g88_n_spl_0, g88_n_spl_);
/*splt*/ buf (g88_n_spl_00, g88_n_spl_0);
/*splt*/ buf (g88_n_spl_000, g88_n_spl_00);
/*splt*/ buf (g88_n_spl_001, g88_n_spl_00);
/*splt*/ buf (g88_n_spl_01, g88_n_spl_0);
/*splt*/ buf (g88_n_spl_1, g88_n_spl_);
/*splt*/ buf (g88_n_spl_10, g88_n_spl_1);
/*splt*/ buf (g88_n_spl_11, g88_n_spl_1);
/*splt*/ buf (g88_p_spl_, g88_p);
/*splt*/ buf (g88_p_spl_0, g88_p_spl_);
/*splt*/ buf (g88_p_spl_00, g88_p_spl_0);
/*splt*/ buf (g88_p_spl_000, g88_p_spl_00);
/*splt*/ buf (g88_p_spl_01, g88_p_spl_0);
/*splt*/ buf (g88_p_spl_1, g88_p_spl_);
/*splt*/ buf (g88_p_spl_10, g88_p_spl_1);
/*splt*/ buf (g88_p_spl_11, g88_p_spl_1);
/*splt*/ buf (g90_p_spl_, g90_p);
/*splt*/ buf (G29_n_spl_, G29_n);
/*splt*/ buf (g90_n_spl_, g90_n);
/*splt*/ buf (G29_p_spl_, G29_p);
/*splt*/ buf (g93_n_spl_, g93_n);
/*splt*/ buf (G33_p_spl_, G33_p);
/*splt*/ buf (g96_p_spl_, g96_p);
/*splt*/ buf (G21_n_spl_, G21_n);
/*splt*/ buf (g96_n_spl_, g96_n);
/*splt*/ buf (G21_p_spl_, G21_p);
/*splt*/ buf (g101_p_spl_, g101_p);
/*splt*/ buf (G13_n_spl_, G13_n);
/*splt*/ buf (g101_n_spl_, g101_n);
/*splt*/ buf (G13_p_spl_, G13_p);
/*splt*/ buf (g104_n_spl_, g104_n);
/*splt*/ buf (G36_p_spl_, G36_p);
/*splt*/ buf (g108_n_spl_, g108_n);
/*splt*/ buf (G25_p_spl_, G25_p);
/*splt*/ buf (g111_n_spl_, g111_n);
/*splt*/ buf (G9_p_spl_, G9_p);
/*splt*/ buf (g115_p_spl_, g115_p);
/*splt*/ buf (G5_n_spl_, G5_n);
/*splt*/ buf (g118_p_spl_, g118_p);
/*splt*/ buf (G17_n_spl_, G17_n);
/*splt*/ buf (g118_n_spl_, g118_n);
/*splt*/ buf (G17_p_spl_, G17_p);
/*splt*/ buf (g123_p_spl_, g123_p);
/*splt*/ buf (g123_p_spl_0, g123_p_spl_);
/*splt*/ buf (g123_p_spl_00, g123_p_spl_0);
/*splt*/ buf (g123_p_spl_1, g123_p_spl_);
/*splt*/ buf (g123_n_spl_, g123_n);
/*splt*/ buf (g123_n_spl_0, g123_n_spl_);
/*splt*/ buf (g123_n_spl_00, g123_n_spl_0);
/*splt*/ buf (g123_n_spl_000, g123_n_spl_00);
/*splt*/ buf (g123_n_spl_01, g123_n_spl_0);
/*splt*/ buf (g123_n_spl_1, g123_n_spl_);
/*splt*/ buf (g123_n_spl_10, g123_n_spl_1);
/*splt*/ buf (g123_n_spl_11, g123_n_spl_1);
/*splt*/ buf (g127_n_spl_, g127_n);
/*splt*/ buf (g134_n_spl_, g134_n);
/*splt*/ buf (g130_p_spl_, g130_p);
/*splt*/ buf (g140_n_spl_, g140_n);
/*splt*/ buf (g145_n_spl_, g145_n);
/*splt*/ buf (g143_n_spl_, g143_n);
/*splt*/ buf (g136_p_spl_, g136_p);
/*splt*/ buf (g129_p_spl_, g129_p);
/*splt*/ buf (g135_n_spl_, g135_n);
/*splt*/ buf (g151_n_spl_, g151_n);

endmodule
