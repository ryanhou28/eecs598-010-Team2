// Benchmark "mymod" written by ABC on Sun Oct 29 23:44:44 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58,
    G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70, G71, G72,
    G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86,
    G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G109, G110, G111, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G124,
    G125, G126, G127, G128, G129, G130, G131, G132, G133, G134, G135, G136,
    G137, G138, G139, G140, G141, G142, G143, G144, G145, G146, G147, G148,
    G149, G150, G151, G152, G153, G154, G155, G156, G157,
    G2531, G2532, G2533, G2534, G2535, G2536, G2537, G2538, G2539, G2540,
    G2541, G2542, G2543, G2544, G2545, G2546, G2547, G2548, G2549, G2550,
    G2551, G2552, G2553, G2554, G2555, G2556, G2557, G2558, G2559, G2560,
    G2561, G2562, G2563, G2564, G2565, G2566, G2567, G2568, G2569, G2570,
    G2571, G2572, G2573, G2574, G2575, G2576, G2577, G2578, G2579, G2580,
    G2581, G2582, G2583, G2584, G2585, G2586, G2587, G2588, G2589, G2590,
    G2591, G2592, G2593, G2594  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G70,
    G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G97, G98,
    G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G110,
    G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G133, G134,
    G135, G136, G137, G138, G139, G140, G141, G142, G143, G144, G145, G146,
    G147, G148, G149, G150, G151, G152, G153, G154, G155, G156, G157;
  output G2531, G2532, G2533, G2534, G2535, G2536, G2537, G2538, G2539, G2540,
    G2541, G2542, G2543, G2544, G2545, G2546, G2547, G2548, G2549, G2550,
    G2551, G2552, G2553, G2554, G2555, G2556, G2557, G2558, G2559, G2560,
    G2561, G2562, G2563, G2564, G2565, G2566, G2567, G2568, G2569, G2570,
    G2571, G2572, G2573, G2574, G2575, G2576, G2577, G2578, G2579, G2580,
    G2581, G2582, G2583, G2584, G2585, G2586, G2587, G2588, G2589, G2590,
    G2591, G2592, G2593, G2594;
  reg n1416_lo, n1419_lo, n1422_lo, n1425_lo, n1428_lo, n1431_lo, n1434_lo,
    n1437_lo, n1440_lo, n1443_lo, n1446_lo, n1449_lo, n1452_lo, n1455_lo,
    n1458_lo, n1464_lo, n1467_lo, n1470_lo, n1476_lo, n1479_lo, n1482_lo,
    n1488_lo, n1491_lo, n1494_lo, n1497_lo, n1500_lo, n1503_lo, n1512_lo,
    n1515_lo, n1518_lo, n1521_lo, n1524_lo, n1527_lo, n1530_lo, n1533_lo,
    n1536_lo, n1539_lo, n1542_lo, n1545_lo, n1548_lo, n1551_lo, n1554_lo,
    n1560_lo, n1563_lo, n1566_lo, n1572_lo, n1575_lo, n1578_lo, n1584_lo,
    n1587_lo, n1590_lo, n1596_lo, n1599_lo, n1602_lo, n1608_lo, n1611_lo,
    n1614_lo, n1620_lo, n1623_lo, n1626_lo, n1632_lo, n1635_lo, n1638_lo,
    n1644_lo, n1647_lo, n1650_lo, n1656_lo, n1659_lo, n1662_lo, n1668_lo,
    n1671_lo, n1674_lo, n1680_lo, n1683_lo, n1686_lo, n1692_lo, n1695_lo,
    n1698_lo, n1704_lo, n1707_lo, n1710_lo, n1716_lo, n1719_lo, n1722_lo,
    n1728_lo, n1731_lo, n1734_lo, n1740_lo, n1743_lo, n1746_lo, n1749_lo,
    n1752_lo, n1755_lo, n1758_lo, n1761_lo, n1764_lo, n1776_lo, n1788_lo,
    n1791_lo, n1794_lo, n1797_lo, n1800_lo, n1803_lo, n1812_lo, n1815_lo,
    n1824_lo, n1827_lo, n1836_lo, n1839_lo, n1848_lo, n1851_lo, n1860_lo,
    n1872_lo, n1875_lo, n1884_lo, n1896_lo, n1899_lo, n1908_lo, n1920_lo,
    n1923_lo, n1926_lo, n1929_lo, n1932_lo, n1935_lo, n1944_lo, n1947_lo,
    n1956_lo, n1959_lo, n1962_lo, n1968_lo, n1971_lo, n1980_lo, n1983_lo,
    n1992_lo, n1995_lo, n2004_lo, n2016_lo, n2019_lo, n2028_lo, n2040_lo,
    n2043_lo, n2046_lo, n2049_lo, n2052_lo, n2055_lo, n2064_lo, n2067_lo,
    n2076_lo, n2079_lo, n2088_lo, n2091_lo, n2100_lo, n2103_lo, n2112_lo,
    n2115_lo, n2124_lo, n2127_lo, n2136_lo, n2148_lo, n2151_lo, n2160_lo,
    n2172_lo, n2175_lo, n2178_lo, n2181_lo, n2184_lo, n2187_lo, n2196_lo,
    n2199_lo, n2208_lo, n2211_lo, n2220_lo, n2223_lo, n2232_lo, n2235_lo,
    n2244_lo, n2247_lo, n2256_lo, n2259_lo, n2268_lo, n2280_lo, n2283_lo,
    n2292_lo, n2295_lo, n2298_lo, n2301_lo, n2304_lo, n2307_lo, n2316_lo,
    n2319_lo, n2322_lo, n2325_lo, n2328_lo, n2331_lo, n2340_lo, n2343_lo,
    n2376_lo, n2379_lo, n2388_lo, n2391_lo, n2400_lo, n2403_lo, n2412_lo,
    n2415_lo, n2424_lo, n2427_lo, n2436_lo, n2439_lo, n2442_lo, n2445_lo,
    n2448_lo, n2451_lo, n2460_lo, n2463_lo, n2496_lo, n2499_lo, n2508_lo,
    n2511_lo, n2520_lo, n2523_lo, n2532_lo, n2535_lo, n2544_lo, n2547_lo,
    n2556_lo, n2559_lo, n2562_lo, n2565_lo, n2568_lo, n2571_lo, n2580_lo,
    n2583_lo, n2616_lo, n2619_lo, n2628_lo, n2631_lo, n2640_lo, n2643_lo,
    n2652_lo, n2655_lo, n2664_lo, n2667_lo, n2676_lo, n2679_lo, n2682_lo,
    n2685_lo, n2688_lo, n2691_lo, n2700_lo, n2703_lo, n2736_lo, n2739_lo,
    n2748_lo, n2751_lo, n2760_lo, n2763_lo, n2772_lo, n2775_lo, n2784_lo,
    n2787_lo, n2790_lo, n2793_lo, n2796_lo, n2799_lo, n2802_lo, n2805_lo,
    n2808_lo, n2820_lo, n2823_lo, n2826_lo, n2829_lo, n2832_lo, n2835_lo,
    n2838_lo, n2841_lo, n2844_lo, n2856_lo, n2859_lo, n2862_lo, n2865_lo,
    n2868_lo, n2871_lo, n2874_lo, n2877_lo, n2880_lo, n2883_lo, n2886_lo,
    n2889_lo, n2892_lo, n2895_lo, n2898_lo, n2901_lo, n2904_lo, n2907_lo,
    n2916_lo, n2919_lo, n2925_lo, n2928_lo, n2940_lo, n2943_lo, n2952_lo,
    n2955_lo, n2961_lo, n2964_lo, n2967_lo, n2970_lo, n2976_lo, n2979_lo,
    n2982_lo, n2988_lo, n2991_lo, n2994_lo, n2997_lo, n3000_lo, n3003_lo,
    n3006_lo, n3012_lo, n3015_lo, n3018_lo, n3021_lo, n3024_lo, n3027_lo,
    n3030_lo, n3033_lo, n3036_lo, n3039_lo, n3045_lo, n3048_lo, n3051_lo,
    n3054_lo, n3057_lo, n3060_lo, n3063_lo, n3069_lo, n3072_lo, n3075_lo,
    n3081_lo, n3084_lo, n3087_lo, n3093_lo, n3096_lo, n3099_lo, n3102_lo,
    n3105_lo, n3108_lo, n3111_lo, n3114_lo, n3117_lo, n3120_lo, n3123_lo,
    n3126_lo, n3129_lo, n3132_lo, n3135_lo, n3138_lo, n3141_lo, n3156_lo,
    n3168_lo, n3171_lo, n3174_lo, n3177_lo, n3180_lo, n3183_lo, n3192_lo,
    n3195_lo, n3204_lo, n3207_lo, n3210_lo, n3216_lo, n3219_lo, n3222_lo,
    n3228_lo, n3231_lo, n3240_lo, n3243_lo, n3252_lo, n3255_lo, n3258_lo,
    n3264_lo, n3267_lo, n3270_lo, n3276_lo, n3279_lo, n3282_lo, n3288_lo,
    n3291_lo, n3294_lo, n3603_o2, n3604_o2, n1391_inv, n3798_o2, n3846_o2,
    n4019_o2, n4017_o2, n2177_o2, n2150_o2, n2154_o2, n2184_o2, n2515_o2,
    n3837_o2, n2167_o2, n2118_o2, n2186_o2, n2174_o2, n3964_o2, n4005_o2,
    n4006_o2, n1445_inv, n2176_o2, n2227_o2, n2236_o2, n2245_o2, n2518_o2,
    n4023_o2, n1466_inv, n4038_o2, n4039_o2, n1475_inv, n2119_o2, n2275_o2,
    n2595_o2, n2594_o2, lo498_buf_o2, lo502_buf_o2, lo550_buf_o2, n2596_o2,
    n2593_o2, n2668_o2, lo542_buf_o2, n2667_o2, n2404_o2, n2410_o2,
    n2419_o2, n2392_o2, n2369_o2, n2397_o2, n2601_o2, n2658_o2, n2574_o2,
    n2205_o2, lo510_buf_o2, lo514_buf_o2, lo554_buf_o2, lo558_buf_o2,
    lo578_buf_o2, n2254_o2, n2421_o2, n2422_o2, n2130_o2, n2127_o2,
    n2131_o2, n2128_o2, n2264_o2, n2467_o2, n2471_o2, n2488_o2, n2478_o2,
    n2486_o2, n2485_o2, n2498_o2, n2495_o2, n2496_o2, n2458_o2, n2643_o2,
    n2462_o2, n2468_o2, n2639_o2, n2499_o2, n2472_o2, n2474_o2, n2489_o2,
    n2321_o2, n2322_o2, n2640_o2, n2642_o2, n2187_o2, n2373_o2, n2603_o2,
    n2388_o2, n2437_o2, n2356_o2, n2452_o2, n2347_o2, n2329_o2, n2669_o2,
    n2332_o2, n2664_o2, n2665_o2, n2653_o2, n2654_o2, n2636_o2, n2660_o2,
    n2318_o2, n2319_o2, n2586_o2, n2587_o2, n2288_o2, n2344_o2, n2530_o2,
    n2303_o2, n2566_o2, n2567_o2, n2554_o2, n2194_o2, lo582_buf_o2,
    lo030_buf_o2, lo174_buf_o2, lo178_buf_o2, lo186_buf_o2, lo266_buf_o2,
    lo306_buf_o2, lo346_buf_o2, lo386_buf_o2, lo426_buf_o2, lo590_buf_o2,
    lo594_buf_o2, lo606_buf_o2, lo610_buf_o2, n2238_o2, n2229_o2, n2242_o2,
    n2233_o2, n2168_o2, n2237_o2, n2228_o2, n2172_o2, n2223_o2, n2222_o2,
    n2170_o2, n2181_o2, n2510_o2, n2621_o2, lo466_buf_o2, lo478_buf_o2,
    n2149_o2, n2429_o2, n2444_o2, n2153_o2, n2433_o2, n2448_o2, n2367_o2,
    n2386_o2, n2539_o2, n2183_o2, n2220_o2, n2514_o2, n2196_o2, n2616_o2,
    n2612_o2, n2627_o2, n2140_o2, n1877_inv, lo149_buf_o2, lo197_buf_o2,
    lo118_buf_o2, lo158_buf_o2, lo166_buf_o2, lo242_buf_o2, lo286_buf_o2,
    lo506_buf_o2, n2198_o2, n2202_o2, n2197_o2, n1913_inv, n2146_o2,
    n1919_inv, lo312_buf_o2, lo316_buf_o2, lo352_buf_o2, lo356_buf_o2,
    lo392_buf_o2, lo396_buf_o2, lo432_buf_o2, lo436_buf_o2, lo576_buf_o2;
  wire new_n1372_, new_n1374_, new_n1376_, new_n1378_, new_n1380_,
    new_n1382_, new_n1384_, new_n1386_, new_n1388_, new_n1390_, new_n1392_,
    new_n1394_, new_n1396_, new_n1398_, new_n1400_, new_n1402_, new_n1404_,
    new_n1406_, new_n1408_, new_n1410_, new_n1412_, new_n1414_, new_n1416_,
    new_n1418_, new_n1420_, new_n1422_, new_n1424_, new_n1426_, new_n1428_,
    new_n1430_, new_n1432_, new_n1434_, new_n1436_, new_n1438_, new_n1440_,
    new_n1442_, new_n1444_, new_n1446_, new_n1448_, new_n1450_, new_n1452_,
    new_n1454_, new_n1456_, new_n1458_, new_n1460_, new_n1462_, new_n1464_,
    new_n1466_, new_n1468_, new_n1470_, new_n1472_, new_n1474_, new_n1476_,
    new_n1478_, new_n1480_, new_n1482_, new_n1484_, new_n1486_, new_n1488_,
    new_n1490_, new_n1492_, new_n1494_, new_n1496_, new_n1498_, new_n1500_,
    new_n1502_, new_n1504_, new_n1506_, new_n1508_, new_n1510_, new_n1512_,
    new_n1514_, new_n1516_, new_n1518_, new_n1520_, new_n1522_, new_n1524_,
    new_n1526_, new_n1528_, new_n1530_, new_n1532_, new_n1534_, new_n1536_,
    new_n1538_, new_n1540_, new_n1542_, new_n1544_, new_n1546_, new_n1548_,
    new_n1550_, new_n1552_, new_n1554_, new_n1556_, new_n1558_, new_n1560_,
    new_n1562_, new_n1564_, new_n1566_, new_n1568_, new_n1570_, new_n1572_,
    new_n1574_, new_n1576_, new_n1578_, new_n1580_, new_n1582_, new_n1584_,
    new_n1586_, new_n1588_, new_n1590_, new_n1592_, new_n1594_, new_n1596_,
    new_n1598_, new_n1600_, new_n1602_, new_n1604_, new_n1606_, new_n1608_,
    new_n1610_, new_n1612_, new_n1614_, new_n1616_, new_n1618_, new_n1620_,
    new_n1622_, new_n1624_, new_n1626_, new_n1628_, new_n1630_, new_n1632_,
    new_n1634_, new_n1636_, new_n1638_, new_n1640_, new_n1642_, new_n1644_,
    new_n1646_, new_n1648_, new_n1650_, new_n1652_, new_n1654_, new_n1656_,
    new_n1658_, new_n1660_, new_n1662_, new_n1664_, new_n1666_, new_n1668_,
    new_n1670_, new_n1672_, new_n1674_, new_n1676_, new_n1678_, new_n1680_,
    new_n1682_, new_n1684_, new_n1686_, new_n1688_, new_n1690_, new_n1692_,
    new_n1694_, new_n1696_, new_n1698_, new_n1701_, new_n1702_, new_n1704_,
    new_n1706_, new_n1708_, new_n1710_, new_n1712_, new_n1714_, new_n1716_,
    new_n1718_, new_n1720_, new_n1722_, new_n1724_, new_n1726_, new_n1728_,
    new_n1730_, new_n1732_, new_n1735_, new_n1736_, new_n1738_, new_n1740_,
    new_n1742_, new_n1744_, new_n1747_, new_n1748_, new_n1750_, new_n1752_,
    new_n1754_, new_n1756_, new_n1758_, new_n1760_, new_n1763_, new_n1764_,
    new_n1766_, new_n1768_, new_n1769_, new_n1770_, new_n1772_, new_n1774_,
    new_n1776_, new_n1778_, new_n1780_, new_n1782_, new_n1784_, new_n1786_,
    new_n1788_, new_n1790_, new_n1792_, new_n1794_, new_n1796_, new_n1798_,
    new_n1800_, new_n1802_, new_n1804_, new_n1806_, new_n1808_, new_n1810_,
    new_n1812_, new_n1814_, new_n1816_, new_n1818_, new_n1820_, new_n1822_,
    new_n1824_, new_n1826_, new_n1828_, new_n1830_, new_n1832_, new_n1834_,
    new_n1835_, new_n1836_, new_n1838_, new_n1840_, new_n1842_, new_n1844_,
    new_n1846_, new_n1848_, new_n1850_, new_n1852_, new_n1854_, new_n1856_,
    new_n1858_, new_n1860_, new_n1862_, new_n1864_, new_n1867_, new_n1868_,
    new_n1870_, new_n1872_, new_n1875_, new_n1876_, new_n1878_, new_n1880_,
    new_n1882_, new_n1884_, new_n1887_, new_n1888_, new_n1890_, new_n1892_,
    new_n1894_, new_n1896_, new_n1899_, new_n1900_, new_n1903_, new_n1904_,
    new_n1907_, new_n1908_, new_n1910_, new_n1912_, new_n1914_, new_n1916_,
    new_n1918_, new_n1920_, new_n1922_, new_n1924_, new_n1926_, new_n1929_,
    new_n1930_, new_n1932_, new_n1934_, new_n1936_, new_n1938_, new_n1940_,
    new_n1942_, new_n1943_, new_n1944_, new_n1946_, new_n1948_, new_n1951_,
    new_n1952_, new_n1954_, new_n1956_, new_n1958_, new_n1960_, new_n1962_,
    new_n1964_, new_n1966_, new_n1968_, new_n1971_, new_n1972_, new_n1974_,
    new_n1976_, new_n1978_, new_n1980_, new_n1982_, new_n1984_, new_n1986_,
    new_n1988_, new_n1990_, new_n1992_, new_n1995_, new_n1996_, new_n1998_,
    new_n2000_, new_n2002_, new_n2004_, new_n2006_, new_n2008_, new_n2010_,
    new_n2012_, new_n2015_, new_n2016_, new_n2018_, new_n2020_, new_n2022_,
    new_n2024_, new_n2026_, new_n2028_, new_n2031_, new_n2032_, new_n2035_,
    new_n2036_, new_n2039_, new_n2040_, new_n2042_, new_n2044_, new_n2046_,
    new_n2048_, new_n2050_, new_n2052_, new_n2054_, new_n2056_, new_n2058_,
    new_n2060_, new_n2062_, new_n2064_, new_n2066_, new_n2069_, new_n2070_,
    new_n2072_, new_n2074_, new_n2076_, new_n2078_, new_n2080_, new_n2082_,
    new_n2084_, new_n2086_, new_n2088_, new_n2090_, new_n2092_, new_n2094_,
    new_n2096_, new_n2098_, new_n2100_, new_n2102_, new_n2105_, new_n2106_,
    new_n2108_, new_n2110_, new_n2112_, new_n2114_, new_n2116_, new_n2118_,
    new_n2120_, new_n2122_, new_n2124_, new_n2126_, new_n2128_, new_n2130_,
    new_n2132_, new_n2134_, new_n2136_, new_n2138_, new_n2141_, new_n2142_,
    new_n2144_, new_n2146_, new_n2148_, new_n2150_, new_n2152_, new_n2154_,
    new_n2156_, new_n2158_, new_n2160_, new_n2162_, new_n2164_, new_n2166_,
    new_n2168_, new_n2170_, new_n2172_, new_n2174_, new_n2177_, new_n2178_,
    new_n2180_, new_n2182_, new_n2184_, new_n2186_, new_n2188_, new_n2190_,
    new_n2192_, new_n2194_, new_n2196_, new_n2198_, new_n2200_, new_n2202_,
    new_n2204_, new_n2206_, new_n2208_, new_n2209_, new_n2210_, new_n2212_,
    new_n2214_, new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2222_,
    new_n2224_, new_n2226_, new_n2227_, new_n2228_, new_n2230_, new_n2232_,
    new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2240_,
    new_n2242_, new_n2244_, new_n2245_, new_n2246_, new_n2248_, new_n2250_,
    new_n2252_, new_n2253_, new_n2254_, new_n2256_, new_n2258_, new_n2260_,
    new_n2261_, new_n2262_, new_n2264_, new_n2266_, new_n2269_, new_n2270_,
    new_n2272_, new_n2274_, new_n2276_, new_n2279_, new_n2280_, new_n2282_,
    new_n2284_, new_n2286_, new_n2288_, new_n2290_, new_n2291_, new_n2292_,
    new_n2294_, new_n2296_, new_n2297_, new_n2298_, new_n2300_, new_n2302_,
    new_n2303_, new_n2304_, new_n2306_, new_n2308_, new_n2309_, new_n2310_,
    new_n2312_, new_n2314_, new_n2316_, new_n2317_, new_n2318_, new_n2320_,
    new_n2322_, new_n2323_, new_n2325_, new_n2326_, new_n2328_, new_n2330_,
    new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2336_, new_n2338_,
    new_n2339_, new_n2340_, new_n2342_, new_n2344_, new_n2347_, new_n2348_,
    new_n2350_, new_n2352_, new_n2353_, new_n2354_, new_n2356_, new_n2358_,
    new_n2360_, new_n2362_, new_n2365_, new_n2366_, new_n2368_, new_n2370_,
    new_n2371_, new_n2372_, new_n2374_, new_n2376_, new_n2378_, new_n2379_,
    new_n2380_, new_n2381_, new_n2382_, new_n2384_, new_n2386_, new_n2387_,
    new_n2388_, new_n2389_, new_n2390_, new_n2392_, new_n2394_, new_n2395_,
    new_n2396_, new_n2398_, new_n2399_, new_n2400_, new_n2402_, new_n2404_,
    new_n2406_, new_n2407_, new_n2408_, new_n2410_, new_n2412_, new_n2414_,
    new_n2416_, new_n2418_, new_n2420_, new_n2421_, new_n2422_, new_n2424_,
    new_n2426_, new_n2427_, new_n2428_, new_n2430_, new_n2432_, new_n2434_,
    new_n2436_, new_n2438_, new_n2440_, new_n2441_, new_n2442_, new_n2444_,
    new_n2446_, new_n2447_, new_n2448_, new_n2450_, new_n2452_, new_n2453_,
    new_n2454_, new_n2456_, new_n2458_, new_n2459_, new_n2461_, new_n2463_,
    new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_,
    new_n2472_, new_n2473_, new_n2474_, new_n2477_, new_n2479_, new_n2480_,
    new_n2482_, new_n2484_, new_n2485_, new_n2487_, new_n2489_, new_n2490_,
    new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_,
    new_n2499_, new_n2501_, new_n2502_, new_n2504_, new_n2506_, new_n2508_,
    new_n2510_, new_n2511_, new_n2512_, new_n2514_, new_n2516_, new_n2517_,
    new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2523_, new_n2524_,
    new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_,
    new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2546_, new_n2548_, new_n2551_, new_n2552_, new_n2555_, new_n2557_,
    new_n2559_, new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_,
    new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_,
    new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_,
    new_n2579_, new_n2581_, new_n2583_, new_n2585_, new_n2587_, new_n2589_,
    new_n2590_, new_n2591_, new_n2592_, new_n2594_, new_n2596_, new_n2598_,
    new_n2600_, new_n2602_, new_n2604_, new_n2606_, new_n2608_, new_n2610_,
    new_n2612_, new_n2613_, new_n2614_, new_n2616_, new_n2618_, new_n2619_,
    new_n2620_, new_n2622_, new_n2624_, new_n2626_, new_n2628_, new_n2629_,
    new_n2630_, new_n2631_, new_n2632_, new_n2634_, new_n2636_, new_n2637_,
    new_n2638_, new_n2639_, new_n2640_, new_n2642_, new_n2643_, new_n2644_,
    new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_,
    new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_,
    new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2662_, new_n2663_,
    new_n2664_, new_n2666_, new_n2668_, new_n2670_, new_n2671_, new_n2672_,
    new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_,
    new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_,
    new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_,
    new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_,
    new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_,
    new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_,
    new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_,
    new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_,
    new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_,
    new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_,
    new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_,
    new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_,
    new_n2745_, new_n2746_, new_n2747_, new_n2749_, new_n2750_, new_n2751_,
    new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_,
    new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_,
    new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_,
    new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_,
    new_n2776_, new_n2777_, new_n2778_, new_n2781_, new_n2783_, new_n2785_,
    new_n2786_, new_n2788_, new_n2791_, new_n2792_, new_n2794_, new_n2795_,
    new_n2796_, new_n2798_, new_n2800_, new_n2802_, new_n2804_, new_n2805_,
    new_n2806_, new_n2808_, new_n2810_, new_n2812_, new_n2813_, new_n2814_,
    new_n2815_, new_n2816_, new_n2817_, new_n2819_, new_n2820_, new_n2823_,
    new_n2824_, new_n2827_, new_n2828_, new_n2831_, new_n2832_, new_n2834_,
    new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_,
    new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_,
    new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_,
    new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_,
    new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_,
    new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_,
    new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_,
    new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_,
    new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_,
    new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_,
    new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_,
    new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_,
    new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_,
    new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_,
    new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_,
    new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_,
    new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_,
    new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_,
    new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_,
    new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_,
    new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_,
    new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_,
    new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_,
    new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_,
    new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_,
    new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_,
    new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_,
    new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_,
    new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_,
    new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_,
    new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_, new_n3020_,
    new_n3021_, new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_,
    new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_,
    new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_,
    new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_,
    new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_,
    new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_,
    new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_,
    new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_,
    new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_,
    new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_,
    new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_,
    new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_,
    new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_,
    new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_,
    new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_,
    new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_,
    new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_,
    new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_,
    new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_,
    new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_,
    new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_,
    new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_,
    new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_,
    new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_,
    new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_,
    new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_,
    new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_,
    new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_,
    new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_,
    new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_,
    new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_,
    new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_,
    new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_,
    new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_,
    new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_,
    new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_,
    new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_,
    new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_,
    new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_,
    new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_,
    new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_,
    new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_,
    new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_,
    new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_,
    new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_,
    new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_,
    new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_,
    new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_,
    new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_,
    new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_,
    new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_,
    new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_,
    new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_,
    new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_,
    new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_,
    new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_,
    new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_,
    new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_,
    new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_,
    new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_,
    new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_,
    new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_,
    new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_,
    new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_,
    new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_,
    new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_,
    new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_,
    new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_,
    new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_,
    new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_,
    new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_,
    new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_,
    new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_,
    new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_,
    new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_,
    new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_,
    new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_,
    new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_,
    new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_,
    new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_,
    new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_,
    new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_,
    new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_,
    new_n3519_, new_n3520_, new_n3521_, new_n4161_, new_n4162_, new_n4163_,
    new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_,
    new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_,
    new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_,
    new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_,
    new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_,
    new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_,
    new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_,
    new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_,
    new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_,
    new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_,
    new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_,
    new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_,
    new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_,
    new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_,
    new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_,
    new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_,
    new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_,
    new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_,
    new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_,
    new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_,
    new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_,
    new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_,
    new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_,
    new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_,
    new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_,
    new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_,
    new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_,
    new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_,
    new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_,
    new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_,
    new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_,
    new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_,
    new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_,
    new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_,
    new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_,
    new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_,
    new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_,
    new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_,
    new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_,
    new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_,
    new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_,
    new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_,
    new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_,
    new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_,
    new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_,
    new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_,
    new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_,
    new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_,
    new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_,
    new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_,
    new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_,
    new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_,
    new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_,
    new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_,
    new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_,
    new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_,
    new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_,
    new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_,
    new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_,
    new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_,
    new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_,
    new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_,
    new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_,
    new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_,
    new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_,
    new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_,
    new_n4614_, new_n4615_, n4649_li000_li000, n4652_li001_li001,
    n4655_li002_li002, n4658_li003_li003, n4661_li004_li004,
    n4664_li005_li005, n4667_li006_li006, n4670_li007_li007,
    n4673_li008_li008, n4676_li009_li009, n4679_li010_li010,
    n4682_li011_li011, n4685_li012_li012, n4688_li013_li013,
    n4691_li014_li014, n4697_li016_li016, n4700_li017_li017,
    n4703_li018_li018, n4709_li020_li020, n4712_li021_li021,
    n4715_li022_li022, n4721_li024_li024, n4724_li025_li025,
    n4727_li026_li026, n4730_li027_li027, n4733_li028_li028,
    n4736_li029_li029, n4745_li032_li032, n4748_li033_li033,
    n4751_li034_li034, n4754_li035_li035, n4757_li036_li036,
    n4760_li037_li037, n4763_li038_li038, n4766_li039_li039,
    n4769_li040_li040, n4772_li041_li041, n4775_li042_li042,
    n4778_li043_li043, n4781_li044_li044, n4784_li045_li045,
    n4787_li046_li046, n4793_li048_li048, n4796_li049_li049,
    n4799_li050_li050, n4805_li052_li052, n4808_li053_li053,
    n4811_li054_li054, n4817_li056_li056, n4820_li057_li057,
    n4823_li058_li058, n4829_li060_li060, n4832_li061_li061,
    n4835_li062_li062, n4841_li064_li064, n4844_li065_li065,
    n4847_li066_li066, n4853_li068_li068, n4856_li069_li069,
    n4859_li070_li070, n4865_li072_li072, n4868_li073_li073,
    n4871_li074_li074, n4877_li076_li076, n4880_li077_li077,
    n4883_li078_li078, n4889_li080_li080, n4892_li081_li081,
    n4895_li082_li082, n4901_li084_li084, n4904_li085_li085,
    n4907_li086_li086, n4913_li088_li088, n4916_li089_li089,
    n4919_li090_li090, n4925_li092_li092, n4928_li093_li093,
    n4931_li094_li094, n4937_li096_li096, n4940_li097_li097,
    n4943_li098_li098, n4949_li100_li100, n4952_li101_li101,
    n4955_li102_li102, n4961_li104_li104, n4964_li105_li105,
    n4967_li106_li106, n4973_li108_li108, n4976_li109_li109,
    n4979_li110_li110, n4982_li111_li111, n4985_li112_li112,
    n4988_li113_li113, n4991_li114_li114, n4994_li115_li115,
    n4997_li116_li116, n5009_li120_li120, n5021_li124_li124,
    n5024_li125_li125, n5027_li126_li126, n5030_li127_li127,
    n5033_li128_li128, n5036_li129_li129, n5045_li132_li132,
    n5048_li133_li133, n5057_li136_li136, n5060_li137_li137,
    n5069_li140_li140, n5072_li141_li141, n5081_li144_li144,
    n5084_li145_li145, n5093_li148_li148, n5105_li152_li152,
    n5108_li153_li153, n5117_li156_li156, n5129_li160_li160,
    n5132_li161_li161, n5141_li164_li164, n5153_li168_li168,
    n5156_li169_li169, n5159_li170_li170, n5162_li171_li171,
    n5165_li172_li172, n5168_li173_li173, n5177_li176_li176,
    n5180_li177_li177, n5189_li180_li180, n5192_li181_li181,
    n5195_li182_li182, n5201_li184_li184, n5204_li185_li185,
    n5213_li188_li188, n5216_li189_li189, n5225_li192_li192,
    n5228_li193_li193, n5237_li196_li196, n5249_li200_li200,
    n5252_li201_li201, n5261_li204_li204, n5273_li208_li208,
    n5276_li209_li209, n5279_li210_li210, n5282_li211_li211,
    n5285_li212_li212, n5288_li213_li213, n5297_li216_li216,
    n5300_li217_li217, n5309_li220_li220, n5312_li221_li221,
    n5321_li224_li224, n5324_li225_li225, n5333_li228_li228,
    n5336_li229_li229, n5345_li232_li232, n5348_li233_li233,
    n5357_li236_li236, n5360_li237_li237, n5369_li240_li240,
    n5381_li244_li244, n5384_li245_li245, n5393_li248_li248,
    n5405_li252_li252, n5408_li253_li253, n5411_li254_li254,
    n5414_li255_li255, n5417_li256_li256, n5420_li257_li257,
    n5429_li260_li260, n5432_li261_li261, n5441_li264_li264,
    n5444_li265_li265, n5453_li268_li268, n5456_li269_li269,
    n5465_li272_li272, n5468_li273_li273, n5477_li276_li276,
    n5480_li277_li277, n5489_li280_li280, n5492_li281_li281,
    n5501_li284_li284, n5513_li288_li288, n5516_li289_li289,
    n5525_li292_li292, n5528_li293_li293, n5531_li294_li294,
    n5534_li295_li295, n5537_li296_li296, n5540_li297_li297,
    n5549_li300_li300, n5552_li301_li301, n5555_li302_li302,
    n5558_li303_li303, n5561_li304_li304, n5564_li305_li305,
    n5573_li308_li308, n5576_li309_li309, n5609_li320_li320,
    n5612_li321_li321, n5621_li324_li324, n5624_li325_li325,
    n5633_li328_li328, n5636_li329_li329, n5645_li332_li332,
    n5648_li333_li333, n5657_li336_li336, n5660_li337_li337,
    n5669_li340_li340, n5672_li341_li341, n5675_li342_li342,
    n5678_li343_li343, n5681_li344_li344, n5684_li345_li345,
    n5693_li348_li348, n5696_li349_li349, n5729_li360_li360,
    n5732_li361_li361, n5741_li364_li364, n5744_li365_li365,
    n5753_li368_li368, n5756_li369_li369, n5765_li372_li372,
    n5768_li373_li373, n5777_li376_li376, n5780_li377_li377,
    n5789_li380_li380, n5792_li381_li381, n5795_li382_li382,
    n5798_li383_li383, n5801_li384_li384, n5804_li385_li385,
    n5813_li388_li388, n5816_li389_li389, n5849_li400_li400,
    n5852_li401_li401, n5861_li404_li404, n5864_li405_li405,
    n5873_li408_li408, n5876_li409_li409, n5885_li412_li412,
    n5888_li413_li413, n5897_li416_li416, n5900_li417_li417,
    n5909_li420_li420, n5912_li421_li421, n5915_li422_li422,
    n5918_li423_li423, n5921_li424_li424, n5924_li425_li425,
    n5933_li428_li428, n5936_li429_li429, n5969_li440_li440,
    n5972_li441_li441, n5981_li444_li444, n5984_li445_li445,
    n5993_li448_li448, n5996_li449_li449, n6005_li452_li452,
    n6008_li453_li453, n6017_li456_li456, n6020_li457_li457,
    n6023_li458_li458, n6026_li459_li459, n6029_li460_li460,
    n6032_li461_li461, n6035_li462_li462, n6038_li463_li463,
    n6041_li464_li464, n6053_li468_li468, n6056_li469_li469,
    n6059_li470_li470, n6062_li471_li471, n6065_li472_li472,
    n6068_li473_li473, n6071_li474_li474, n6074_li475_li475,
    n6077_li476_li476, n6089_li480_li480, n6092_li481_li481,
    n6095_li482_li482, n6098_li483_li483, n6101_li484_li484,
    n6104_li485_li485, n6107_li486_li486, n6110_li487_li487,
    n6113_li488_li488, n6116_li489_li489, n6119_li490_li490,
    n6122_li491_li491, n6125_li492_li492, n6128_li493_li493,
    n6131_li494_li494, n6134_li495_li495, n6137_li496_li496,
    n6140_li497_li497, n6149_li500_li500, n6152_li501_li501,
    n6158_li503_li503, n6161_li504_li504, n6173_li508_li508,
    n6176_li509_li509, n6185_li512_li512, n6188_li513_li513,
    n6194_li515_li515, n6197_li516_li516, n6200_li517_li517,
    n6203_li518_li518, n6209_li520_li520, n6212_li521_li521,
    n6215_li522_li522, n6221_li524_li524, n6224_li525_li525,
    n6227_li526_li526, n6230_li527_li527, n6233_li528_li528,
    n6236_li529_li529, n6239_li530_li530, n6245_li532_li532,
    n6248_li533_li533, n6251_li534_li534, n6254_li535_li535,
    n6257_li536_li536, n6260_li537_li537, n6263_li538_li538,
    n6266_li539_li539, n6269_li540_li540, n6272_li541_li541,
    n6278_li543_li543, n6281_li544_li544, n6284_li545_li545,
    n6287_li546_li546, n6290_li547_li547, n6293_li548_li548,
    n6296_li549_li549, n6302_li551_li551, n6305_li552_li552,
    n6308_li553_li553, n6314_li555_li555, n6317_li556_li556,
    n6320_li557_li557, n6326_li559_li559, n6329_li560_li560,
    n6332_li561_li561, n6335_li562_li562, n6338_li563_li563,
    n6341_li564_li564, n6344_li565_li565, n6347_li566_li566,
    n6350_li567_li567, n6353_li568_li568, n6356_li569_li569,
    n6359_li570_li570, n6362_li571_li571, n6365_li572_li572,
    n6368_li573_li573, n6371_li574_li574, n6374_li575_li575,
    n6389_li580_li580, n6401_li584_li584, n6404_li585_li585,
    n6407_li586_li586, n6410_li587_li587, n6413_li588_li588,
    n6416_li589_li589, n6425_li592_li592, n6428_li593_li593,
    n6437_li596_li596, n6440_li597_li597, n6443_li598_li598,
    n6449_li600_li600, n6452_li601_li601, n6455_li602_li602,
    n6461_li604_li604, n6464_li605_li605, n6473_li608_li608,
    n6476_li609_li609, n6485_li612_li612, n6488_li613_li613,
    n6491_li614_li614, n6497_li616_li616, n6500_li617_li617,
    n6503_li618_li618, n6509_li620_li620, n6512_li621_li621,
    n6515_li622_li622, n6521_li624_li624, n6524_li625_li625,
    n6527_li626_li626, n3603_i2, n3604_i2, n3618_i2, n3798_i2, n3846_i2,
    n4019_i2, n4017_i2, n2177_i2, n2150_i2, n2154_i2, n2184_i2, n2515_i2,
    n3837_i2, n2167_i2, n2118_i2, n2186_i2, n2174_i2, n3964_i2, n4005_i2,
    n4006_i2, n2195_i2, n2176_i2, n2227_i2, n2236_i2, n2245_i2, n2518_i2,
    n4023_i2, n4024_i2, n4038_i2, n4039_i2, n4040_i2, n2119_i2, n2275_i2,
    n2595_i2, n2594_i2, lo498_buf_i2, lo502_buf_i2, lo550_buf_i2, n2596_i2,
    n2593_i2, n2668_i2, lo542_buf_i2, n2667_i2, n2404_i2, n2410_i2,
    n2419_i2, n2392_i2, n2369_i2, n2397_i2, n2601_i2, n2658_i2, n2574_i2,
    n2205_i2, lo510_buf_i2, lo514_buf_i2, lo554_buf_i2, lo558_buf_i2,
    lo578_buf_i2, n2254_i2, n2421_i2, n2422_i2, n2130_i2, n2127_i2,
    n2131_i2, n2128_i2, n2264_i2, n2467_i2, n2471_i2, n2488_i2, n2478_i2,
    n2486_i2, n2485_i2, n2498_i2, n2495_i2, n2496_i2, n2458_i2, n2643_i2,
    n2462_i2, n2468_i2, n2639_i2, n2499_i2, n2472_i2, n2474_i2, n2489_i2,
    n2321_i2, n2322_i2, n2640_i2, n2642_i2, n2187_i2, n2373_i2, n2603_i2,
    n2388_i2, n2437_i2, n2356_i2, n2452_i2, n2347_i2, n2329_i2, n2669_i2,
    n2332_i2, n2664_i2, n2665_i2, n2653_i2, n2654_i2, n2636_i2, n2660_i2,
    n2318_i2, n2319_i2, n2586_i2, n2587_i2, n2288_i2, n2344_i2, n2530_i2,
    n2303_i2, n2566_i2, n2567_i2, n2554_i2, n2194_i2, lo582_buf_i2,
    lo030_buf_i2, lo174_buf_i2, lo178_buf_i2, lo186_buf_i2, lo266_buf_i2,
    lo306_buf_i2, lo346_buf_i2, lo386_buf_i2, lo426_buf_i2, lo590_buf_i2,
    lo594_buf_i2, lo606_buf_i2, lo610_buf_i2, n2238_i2, n2229_i2, n2242_i2,
    n2233_i2, n2168_i2, n2237_i2, n2228_i2, n2172_i2, n2223_i2, n2222_i2,
    n2170_i2, n2181_i2, n2510_i2, n2621_i2, lo466_buf_i2, lo478_buf_i2,
    n2149_i2, n2429_i2, n2444_i2, n2153_i2, n2433_i2, n2448_i2, n2367_i2,
    n2386_i2, n2539_i2, n2183_i2, n2220_i2, n2514_i2, n2196_i2, n2616_i2,
    n2612_i2, n2627_i2, n2140_i2, n2144_i2, lo149_buf_i2, lo197_buf_i2,
    lo118_buf_i2, lo158_buf_i2, lo166_buf_i2, lo242_buf_i2, lo286_buf_i2,
    lo506_buf_i2, n2198_i2, n2202_i2, n2197_i2, n2166_i2, n2146_i2,
    n2165_i2, lo312_buf_i2, lo316_buf_i2, lo352_buf_i2, lo356_buf_i2,
    lo392_buf_i2, lo396_buf_i2, lo432_buf_i2, lo436_buf_i2, lo576_buf_i2;
  assign new_n1372_ = G1;
  assign new_n1374_ = G2;
  assign new_n1376_ = G3;
  assign new_n1378_ = G4;
  assign new_n1380_ = G5;
  assign new_n1382_ = G6;
  assign new_n1384_ = G7;
  assign new_n1386_ = G8;
  assign new_n1388_ = G9;
  assign new_n1390_ = G10;
  assign new_n1392_ = G11;
  assign new_n1394_ = G12;
  assign new_n1396_ = G13;
  assign new_n1398_ = G14;
  assign new_n1400_ = G15;
  assign new_n1402_ = G16;
  assign new_n1404_ = G17;
  assign new_n1406_ = G18;
  assign new_n1408_ = G19;
  assign new_n1410_ = G20;
  assign new_n1412_ = G21;
  assign new_n1414_ = G22;
  assign new_n1416_ = G23;
  assign new_n1418_ = G24;
  assign new_n1420_ = G25;
  assign new_n1422_ = G26;
  assign new_n1424_ = G27;
  assign new_n1426_ = G28;
  assign new_n1428_ = G29;
  assign new_n1430_ = G30;
  assign new_n1432_ = G31;
  assign new_n1434_ = G32;
  assign new_n1436_ = G33;
  assign new_n1438_ = G34;
  assign new_n1440_ = G35;
  assign new_n1442_ = G36;
  assign new_n1444_ = G37;
  assign new_n1446_ = G38;
  assign new_n1448_ = G39;
  assign new_n1450_ = G40;
  assign new_n1452_ = G41;
  assign new_n1454_ = G42;
  assign new_n1456_ = G43;
  assign new_n1458_ = G44;
  assign new_n1460_ = G45;
  assign new_n1462_ = G46;
  assign new_n1464_ = G47;
  assign new_n1466_ = G48;
  assign new_n1468_ = G49;
  assign new_n1470_ = G50;
  assign new_n1472_ = G51;
  assign new_n1474_ = G52;
  assign new_n1476_ = G53;
  assign new_n1478_ = G54;
  assign new_n1480_ = G55;
  assign new_n1482_ = G56;
  assign new_n1484_ = G57;
  assign new_n1486_ = G58;
  assign new_n1488_ = G59;
  assign new_n1490_ = G60;
  assign new_n1492_ = G61;
  assign new_n1494_ = G62;
  assign new_n1496_ = G63;
  assign new_n1498_ = G64;
  assign new_n1500_ = G65;
  assign new_n1502_ = G66;
  assign new_n1504_ = G67;
  assign new_n1506_ = G68;
  assign new_n1508_ = G69;
  assign new_n1510_ = G70;
  assign new_n1512_ = G71;
  assign new_n1514_ = G72;
  assign new_n1516_ = G73;
  assign new_n1518_ = G74;
  assign new_n1520_ = G75;
  assign new_n1522_ = G76;
  assign new_n1524_ = G77;
  assign new_n1526_ = G78;
  assign new_n1528_ = G79;
  assign new_n1530_ = G80;
  assign new_n1532_ = G81;
  assign new_n1534_ = G82;
  assign new_n1536_ = G83;
  assign new_n1538_ = G84;
  assign new_n1540_ = G85;
  assign new_n1542_ = G86;
  assign new_n1544_ = G87;
  assign new_n1546_ = G88;
  assign new_n1548_ = G89;
  assign new_n1550_ = G90;
  assign new_n1552_ = G91;
  assign new_n1554_ = G92;
  assign new_n1556_ = G93;
  assign new_n1558_ = G94;
  assign new_n1560_ = G95;
  assign new_n1562_ = G96;
  assign new_n1564_ = G97;
  assign new_n1566_ = G98;
  assign new_n1568_ = G99;
  assign new_n1570_ = G100;
  assign new_n1572_ = G101;
  assign new_n1574_ = G102;
  assign new_n1576_ = G103;
  assign new_n1578_ = G104;
  assign new_n1580_ = G105;
  assign new_n1582_ = G106;
  assign new_n1584_ = G107;
  assign new_n1586_ = G108;
  assign new_n1588_ = G109;
  assign new_n1590_ = G110;
  assign new_n1592_ = G111;
  assign new_n1594_ = G112;
  assign new_n1596_ = G113;
  assign new_n1598_ = G114;
  assign new_n1600_ = G115;
  assign new_n1602_ = G116;
  assign new_n1604_ = G117;
  assign new_n1606_ = G118;
  assign new_n1608_ = G119;
  assign new_n1610_ = G120;
  assign new_n1612_ = G121;
  assign new_n1614_ = G122;
  assign new_n1616_ = G123;
  assign new_n1618_ = G124;
  assign new_n1620_ = G125;
  assign new_n1622_ = G126;
  assign new_n1624_ = G127;
  assign new_n1626_ = G128;
  assign new_n1628_ = G129;
  assign new_n1630_ = G130;
  assign new_n1632_ = G131;
  assign new_n1634_ = G132;
  assign new_n1636_ = G133;
  assign new_n1638_ = G134;
  assign new_n1640_ = G135;
  assign new_n1642_ = G136;
  assign new_n1644_ = G137;
  assign new_n1646_ = G138;
  assign new_n1648_ = G139;
  assign new_n1650_ = G140;
  assign new_n1652_ = G141;
  assign new_n1654_ = G142;
  assign new_n1656_ = G143;
  assign new_n1658_ = G144;
  assign new_n1660_ = G145;
  assign new_n1662_ = G146;
  assign new_n1664_ = G147;
  assign new_n1666_ = G148;
  assign new_n1668_ = G149;
  assign new_n1670_ = G150;
  assign new_n1672_ = G151;
  assign new_n1674_ = G152;
  assign new_n1676_ = G153;
  assign new_n1678_ = G154;
  assign new_n1680_ = G155;
  assign new_n1682_ = G156;
  assign new_n1684_ = G157;
  assign new_n1686_ = n1416_lo;
  assign new_n1688_ = n1419_lo;
  assign new_n1690_ = n1422_lo;
  assign new_n1692_ = n1425_lo;
  assign new_n1694_ = n1428_lo;
  assign new_n1696_ = n1431_lo;
  assign new_n1698_ = n1434_lo;
  assign new_n1701_ = ~n1437_lo;
  assign new_n1702_ = n1440_lo;
  assign new_n1704_ = n1443_lo;
  assign new_n1706_ = n1446_lo;
  assign new_n1708_ = n1449_lo;
  assign new_n1710_ = n1452_lo;
  assign new_n1712_ = n1455_lo;
  assign new_n1714_ = n1458_lo;
  assign new_n1716_ = n1464_lo;
  assign new_n1718_ = n1467_lo;
  assign new_n1720_ = n1470_lo;
  assign new_n1722_ = n1476_lo;
  assign new_n1724_ = n1479_lo;
  assign new_n1726_ = n1482_lo;
  assign new_n1728_ = n1488_lo;
  assign new_n1730_ = n1491_lo;
  assign new_n1732_ = n1494_lo;
  assign new_n1735_ = ~n1497_lo;
  assign new_n1736_ = n1500_lo;
  assign new_n1738_ = n1503_lo;
  assign new_n1740_ = n1512_lo;
  assign new_n1742_ = n1515_lo;
  assign new_n1744_ = n1518_lo;
  assign new_n1747_ = ~n1521_lo;
  assign new_n1748_ = n1524_lo;
  assign new_n1750_ = n1527_lo;
  assign new_n1752_ = n1530_lo;
  assign new_n1754_ = n1533_lo;
  assign new_n1756_ = n1536_lo;
  assign new_n1758_ = n1539_lo;
  assign new_n1760_ = n1542_lo;
  assign new_n1763_ = ~n1545_lo;
  assign new_n1764_ = n1548_lo;
  assign new_n1766_ = n1551_lo;
  assign new_n1768_ = n1554_lo;
  assign new_n1769_ = ~n1554_lo;
  assign new_n1770_ = n1560_lo;
  assign new_n1772_ = n1563_lo;
  assign new_n1774_ = n1566_lo;
  assign new_n1776_ = n1572_lo;
  assign new_n1778_ = n1575_lo;
  assign new_n1780_ = n1578_lo;
  assign new_n1782_ = n1584_lo;
  assign new_n1784_ = n1587_lo;
  assign new_n1786_ = n1590_lo;
  assign new_n1788_ = n1596_lo;
  assign new_n1790_ = n1599_lo;
  assign new_n1792_ = n1602_lo;
  assign new_n1794_ = n1608_lo;
  assign new_n1796_ = n1611_lo;
  assign new_n1798_ = n1614_lo;
  assign new_n1800_ = n1620_lo;
  assign new_n1802_ = n1623_lo;
  assign new_n1804_ = n1626_lo;
  assign new_n1806_ = n1632_lo;
  assign new_n1808_ = n1635_lo;
  assign new_n1810_ = n1638_lo;
  assign new_n1812_ = n1644_lo;
  assign new_n1814_ = n1647_lo;
  assign new_n1816_ = n1650_lo;
  assign new_n1818_ = n1656_lo;
  assign new_n1820_ = n1659_lo;
  assign new_n1822_ = n1662_lo;
  assign new_n1824_ = n1668_lo;
  assign new_n1826_ = n1671_lo;
  assign new_n1828_ = n1674_lo;
  assign new_n1830_ = n1680_lo;
  assign new_n1832_ = n1683_lo;
  assign new_n1834_ = n1686_lo;
  assign new_n1835_ = ~n1686_lo;
  assign new_n1836_ = n1692_lo;
  assign new_n1838_ = n1695_lo;
  assign new_n1840_ = n1698_lo;
  assign new_n1842_ = n1704_lo;
  assign new_n1844_ = n1707_lo;
  assign new_n1846_ = n1710_lo;
  assign new_n1848_ = n1716_lo;
  assign new_n1850_ = n1719_lo;
  assign new_n1852_ = n1722_lo;
  assign new_n1854_ = n1728_lo;
  assign new_n1856_ = n1731_lo;
  assign new_n1858_ = n1734_lo;
  assign new_n1860_ = n1740_lo;
  assign new_n1862_ = n1743_lo;
  assign new_n1864_ = n1746_lo;
  assign new_n1867_ = ~n1749_lo;
  assign new_n1868_ = n1752_lo;
  assign new_n1870_ = n1755_lo;
  assign new_n1872_ = n1758_lo;
  assign new_n1875_ = ~n1761_lo;
  assign new_n1876_ = n1764_lo;
  assign new_n1878_ = n1776_lo;
  assign new_n1880_ = n1788_lo;
  assign new_n1882_ = n1791_lo;
  assign new_n1884_ = n1794_lo;
  assign new_n1887_ = ~n1797_lo;
  assign new_n1888_ = n1800_lo;
  assign new_n1890_ = n1803_lo;
  assign new_n1892_ = n1812_lo;
  assign new_n1894_ = n1815_lo;
  assign new_n1896_ = n1824_lo;
  assign new_n1899_ = ~n1827_lo;
  assign new_n1900_ = n1836_lo;
  assign new_n1903_ = ~n1839_lo;
  assign new_n1904_ = n1848_lo;
  assign new_n1907_ = ~n1851_lo;
  assign new_n1908_ = n1860_lo;
  assign new_n1910_ = n1872_lo;
  assign new_n1912_ = n1875_lo;
  assign new_n1914_ = n1884_lo;
  assign new_n1916_ = n1896_lo;
  assign new_n1918_ = n1899_lo;
  assign new_n1920_ = n1908_lo;
  assign new_n1922_ = n1920_lo;
  assign new_n1924_ = n1923_lo;
  assign new_n1926_ = n1926_lo;
  assign new_n1929_ = ~n1929_lo;
  assign new_n1930_ = n1932_lo;
  assign new_n1932_ = n1935_lo;
  assign new_n1934_ = n1944_lo;
  assign new_n1936_ = n1947_lo;
  assign new_n1938_ = n1956_lo;
  assign new_n1940_ = n1959_lo;
  assign new_n1942_ = n1962_lo;
  assign new_n1943_ = ~n1962_lo;
  assign new_n1944_ = n1968_lo;
  assign new_n1946_ = n1971_lo;
  assign new_n1948_ = n1980_lo;
  assign new_n1951_ = ~n1983_lo;
  assign new_n1952_ = n1992_lo;
  assign new_n1954_ = n1995_lo;
  assign new_n1956_ = n2004_lo;
  assign new_n1958_ = n2016_lo;
  assign new_n1960_ = n2019_lo;
  assign new_n1962_ = n2028_lo;
  assign new_n1964_ = n2040_lo;
  assign new_n1966_ = n2043_lo;
  assign new_n1968_ = n2046_lo;
  assign new_n1971_ = ~n2049_lo;
  assign new_n1972_ = n2052_lo;
  assign new_n1974_ = n2055_lo;
  assign new_n1976_ = n2064_lo;
  assign new_n1978_ = n2067_lo;
  assign new_n1980_ = n2076_lo;
  assign new_n1982_ = n2079_lo;
  assign new_n1984_ = n2088_lo;
  assign new_n1986_ = n2091_lo;
  assign new_n1988_ = n2100_lo;
  assign new_n1990_ = n2103_lo;
  assign new_n1992_ = n2112_lo;
  assign new_n1995_ = ~n2115_lo;
  assign new_n1996_ = n2124_lo;
  assign new_n1998_ = n2127_lo;
  assign new_n2000_ = n2136_lo;
  assign new_n2002_ = n2148_lo;
  assign new_n2004_ = n2151_lo;
  assign new_n2006_ = n2160_lo;
  assign new_n2008_ = n2172_lo;
  assign new_n2010_ = n2175_lo;
  assign new_n2012_ = n2178_lo;
  assign new_n2015_ = ~n2181_lo;
  assign new_n2016_ = n2184_lo;
  assign new_n2018_ = n2187_lo;
  assign new_n2020_ = n2196_lo;
  assign new_n2022_ = n2199_lo;
  assign new_n2024_ = n2208_lo;
  assign new_n2026_ = n2211_lo;
  assign new_n2028_ = n2220_lo;
  assign new_n2031_ = ~n2223_lo;
  assign new_n2032_ = n2232_lo;
  assign new_n2035_ = ~n2235_lo;
  assign new_n2036_ = n2244_lo;
  assign new_n2039_ = ~n2247_lo;
  assign new_n2040_ = n2256_lo;
  assign new_n2042_ = n2259_lo;
  assign new_n2044_ = n2268_lo;
  assign new_n2046_ = n2280_lo;
  assign new_n2048_ = n2283_lo;
  assign new_n2050_ = n2292_lo;
  assign new_n2052_ = n2295_lo;
  assign new_n2054_ = n2298_lo;
  assign new_n2056_ = n2301_lo;
  assign new_n2058_ = n2304_lo;
  assign new_n2060_ = n2307_lo;
  assign new_n2062_ = n2316_lo;
  assign new_n2064_ = n2319_lo;
  assign new_n2066_ = n2322_lo;
  assign new_n2069_ = ~n2325_lo;
  assign new_n2070_ = n2328_lo;
  assign new_n2072_ = n2331_lo;
  assign new_n2074_ = n2340_lo;
  assign new_n2076_ = n2343_lo;
  assign new_n2078_ = n2376_lo;
  assign new_n2080_ = n2379_lo;
  assign new_n2082_ = n2388_lo;
  assign new_n2084_ = n2391_lo;
  assign new_n2086_ = n2400_lo;
  assign new_n2088_ = n2403_lo;
  assign new_n2090_ = n2412_lo;
  assign new_n2092_ = n2415_lo;
  assign new_n2094_ = n2424_lo;
  assign new_n2096_ = n2427_lo;
  assign new_n2098_ = n2436_lo;
  assign new_n2100_ = n2439_lo;
  assign new_n2102_ = n2442_lo;
  assign new_n2105_ = ~n2445_lo;
  assign new_n2106_ = n2448_lo;
  assign new_n2108_ = n2451_lo;
  assign new_n2110_ = n2460_lo;
  assign new_n2112_ = n2463_lo;
  assign new_n2114_ = n2496_lo;
  assign new_n2116_ = n2499_lo;
  assign new_n2118_ = n2508_lo;
  assign new_n2120_ = n2511_lo;
  assign new_n2122_ = n2520_lo;
  assign new_n2124_ = n2523_lo;
  assign new_n2126_ = n2532_lo;
  assign new_n2128_ = n2535_lo;
  assign new_n2130_ = n2544_lo;
  assign new_n2132_ = n2547_lo;
  assign new_n2134_ = n2556_lo;
  assign new_n2136_ = n2559_lo;
  assign new_n2138_ = n2562_lo;
  assign new_n2141_ = ~n2565_lo;
  assign new_n2142_ = n2568_lo;
  assign new_n2144_ = n2571_lo;
  assign new_n2146_ = n2580_lo;
  assign new_n2148_ = n2583_lo;
  assign new_n2150_ = n2616_lo;
  assign new_n2152_ = n2619_lo;
  assign new_n2154_ = n2628_lo;
  assign new_n2156_ = n2631_lo;
  assign new_n2158_ = n2640_lo;
  assign new_n2160_ = n2643_lo;
  assign new_n2162_ = n2652_lo;
  assign new_n2164_ = n2655_lo;
  assign new_n2166_ = n2664_lo;
  assign new_n2168_ = n2667_lo;
  assign new_n2170_ = n2676_lo;
  assign new_n2172_ = n2679_lo;
  assign new_n2174_ = n2682_lo;
  assign new_n2177_ = ~n2685_lo;
  assign new_n2178_ = n2688_lo;
  assign new_n2180_ = n2691_lo;
  assign new_n2182_ = n2700_lo;
  assign new_n2184_ = n2703_lo;
  assign new_n2186_ = n2736_lo;
  assign new_n2188_ = n2739_lo;
  assign new_n2190_ = n2748_lo;
  assign new_n2192_ = n2751_lo;
  assign new_n2194_ = n2760_lo;
  assign new_n2196_ = n2763_lo;
  assign new_n2198_ = n2772_lo;
  assign new_n2200_ = n2775_lo;
  assign new_n2202_ = n2784_lo;
  assign new_n2204_ = n2787_lo;
  assign new_n2206_ = n2790_lo;
  assign new_n2208_ = n2793_lo;
  assign new_n2209_ = ~n2793_lo;
  assign new_n2210_ = n2796_lo;
  assign new_n2212_ = n2799_lo;
  assign new_n2214_ = n2802_lo;
  assign new_n2217_ = ~n2805_lo;
  assign new_n2218_ = n2808_lo;
  assign new_n2219_ = ~n2808_lo;
  assign new_n2220_ = n2820_lo;
  assign new_n2222_ = n2823_lo;
  assign new_n2224_ = n2826_lo;
  assign new_n2226_ = n2829_lo;
  assign new_n2227_ = ~n2829_lo;
  assign new_n2228_ = n2832_lo;
  assign new_n2230_ = n2835_lo;
  assign new_n2232_ = n2838_lo;
  assign new_n2234_ = n2841_lo;
  assign new_n2235_ = ~n2841_lo;
  assign new_n2236_ = n2844_lo;
  assign new_n2237_ = ~n2844_lo;
  assign new_n2238_ = n2856_lo;
  assign new_n2240_ = n2859_lo;
  assign new_n2242_ = n2862_lo;
  assign new_n2244_ = n2865_lo;
  assign new_n2245_ = ~n2865_lo;
  assign new_n2246_ = n2868_lo;
  assign new_n2248_ = n2871_lo;
  assign new_n2250_ = n2874_lo;
  assign new_n2252_ = n2877_lo;
  assign new_n2253_ = ~n2877_lo;
  assign new_n2254_ = n2880_lo;
  assign new_n2256_ = n2883_lo;
  assign new_n2258_ = n2886_lo;
  assign new_n2260_ = n2889_lo;
  assign new_n2261_ = ~n2889_lo;
  assign new_n2262_ = n2892_lo;
  assign new_n2264_ = n2895_lo;
  assign new_n2266_ = n2898_lo;
  assign new_n2269_ = ~n2901_lo;
  assign new_n2270_ = n2904_lo;
  assign new_n2272_ = n2907_lo;
  assign new_n2274_ = n2916_lo;
  assign new_n2276_ = n2919_lo;
  assign new_n2279_ = ~n2925_lo;
  assign new_n2280_ = n2928_lo;
  assign new_n2282_ = n2940_lo;
  assign new_n2284_ = n2943_lo;
  assign new_n2286_ = n2952_lo;
  assign new_n2288_ = n2955_lo;
  assign new_n2290_ = n2961_lo;
  assign new_n2291_ = ~n2961_lo;
  assign new_n2292_ = n2964_lo;
  assign new_n2294_ = n2967_lo;
  assign new_n2296_ = n2970_lo;
  assign new_n2297_ = ~n2970_lo;
  assign new_n2298_ = n2976_lo;
  assign new_n2300_ = n2979_lo;
  assign new_n2302_ = n2982_lo;
  assign new_n2303_ = ~n2982_lo;
  assign new_n2304_ = n2988_lo;
  assign new_n2306_ = n2991_lo;
  assign new_n2308_ = n2994_lo;
  assign new_n2309_ = ~n2994_lo;
  assign new_n2310_ = n2997_lo;
  assign new_n2312_ = n3000_lo;
  assign new_n2314_ = n3003_lo;
  assign new_n2316_ = n3006_lo;
  assign new_n2317_ = ~n3006_lo;
  assign new_n2318_ = n3012_lo;
  assign new_n2320_ = n3015_lo;
  assign new_n2322_ = n3018_lo;
  assign new_n2323_ = ~n3018_lo;
  assign new_n2325_ = ~n3021_lo;
  assign new_n2326_ = n3024_lo;
  assign new_n2328_ = n3027_lo;
  assign new_n2330_ = n3030_lo;
  assign new_n2331_ = ~n3030_lo;
  assign new_n2332_ = n3033_lo;
  assign new_n2333_ = ~n3033_lo;
  assign new_n2334_ = n3036_lo;
  assign new_n2336_ = n3039_lo;
  assign new_n2338_ = n3045_lo;
  assign new_n2339_ = ~n3045_lo;
  assign new_n2340_ = n3048_lo;
  assign new_n2342_ = n3051_lo;
  assign new_n2344_ = n3054_lo;
  assign new_n2347_ = ~n3057_lo;
  assign new_n2348_ = n3060_lo;
  assign new_n2350_ = n3063_lo;
  assign new_n2352_ = n3069_lo;
  assign new_n2353_ = ~n3069_lo;
  assign new_n2354_ = n3072_lo;
  assign new_n2356_ = n3075_lo;
  assign new_n2358_ = n3081_lo;
  assign new_n2360_ = n3084_lo;
  assign new_n2362_ = n3087_lo;
  assign new_n2365_ = ~n3093_lo;
  assign new_n2366_ = n3096_lo;
  assign new_n2368_ = n3099_lo;
  assign new_n2370_ = n3102_lo;
  assign new_n2371_ = ~n3102_lo;
  assign new_n2372_ = n3105_lo;
  assign new_n2374_ = n3108_lo;
  assign new_n2376_ = n3111_lo;
  assign new_n2378_ = n3114_lo;
  assign new_n2379_ = ~n3114_lo;
  assign new_n2380_ = n3117_lo;
  assign new_n2381_ = ~n3117_lo;
  assign new_n2382_ = n3120_lo;
  assign new_n2384_ = n3123_lo;
  assign new_n2386_ = n3126_lo;
  assign new_n2387_ = ~n3126_lo;
  assign new_n2388_ = n3129_lo;
  assign new_n2389_ = ~n3129_lo;
  assign new_n2390_ = n3132_lo;
  assign new_n2392_ = n3135_lo;
  assign new_n2394_ = n3138_lo;
  assign new_n2395_ = ~n3138_lo;
  assign new_n2396_ = n3141_lo;
  assign new_n2398_ = n3156_lo;
  assign new_n2399_ = ~n3156_lo;
  assign new_n2400_ = n3168_lo;
  assign new_n2402_ = n3171_lo;
  assign new_n2404_ = n3174_lo;
  assign new_n2406_ = n3177_lo;
  assign new_n2407_ = ~n3177_lo;
  assign new_n2408_ = n3180_lo;
  assign new_n2410_ = n3183_lo;
  assign new_n2412_ = n3192_lo;
  assign new_n2414_ = n3195_lo;
  assign new_n2416_ = n3204_lo;
  assign new_n2418_ = n3207_lo;
  assign new_n2420_ = n3210_lo;
  assign new_n2421_ = ~n3210_lo;
  assign new_n2422_ = n3216_lo;
  assign new_n2424_ = n3219_lo;
  assign new_n2426_ = n3222_lo;
  assign new_n2427_ = ~n3222_lo;
  assign new_n2428_ = n3228_lo;
  assign new_n2430_ = n3231_lo;
  assign new_n2432_ = n3240_lo;
  assign new_n2434_ = n3243_lo;
  assign new_n2436_ = n3252_lo;
  assign new_n2438_ = n3255_lo;
  assign new_n2440_ = n3258_lo;
  assign new_n2441_ = ~n3258_lo;
  assign new_n2442_ = n3264_lo;
  assign new_n2444_ = n3267_lo;
  assign new_n2446_ = n3270_lo;
  assign new_n2447_ = ~n3270_lo;
  assign new_n2448_ = n3276_lo;
  assign new_n2450_ = n3279_lo;
  assign new_n2452_ = n3282_lo;
  assign new_n2453_ = ~n3282_lo;
  assign new_n2454_ = n3288_lo;
  assign new_n2456_ = n3291_lo;
  assign new_n2458_ = n3294_lo;
  assign new_n2459_ = ~n3294_lo;
  assign new_n2461_ = ~n3603_o2;
  assign new_n2463_ = ~n3604_o2;
  assign new_n2465_ = ~n1391_inv;
  assign new_n2466_ = n3798_o2;
  assign new_n2467_ = ~n3798_o2;
  assign new_n2468_ = n3846_o2;
  assign new_n2469_ = ~n3846_o2;
  assign new_n2470_ = n4019_o2;
  assign new_n2472_ = n4017_o2;
  assign new_n2473_ = ~n4017_o2;
  assign new_n2474_ = n2177_o2;
  assign new_n2477_ = ~n2150_o2;
  assign new_n2479_ = ~n2154_o2;
  assign new_n2480_ = n2184_o2;
  assign new_n2482_ = n2515_o2;
  assign new_n2484_ = n3837_o2;
  assign new_n2485_ = ~n3837_o2;
  assign new_n2487_ = ~n2167_o2;
  assign new_n2489_ = ~n2118_o2;
  assign new_n2490_ = n2186_o2;
  assign new_n2493_ = ~n2174_o2;
  assign new_n2494_ = n3964_o2;
  assign new_n2495_ = ~n3964_o2;
  assign new_n2496_ = n4005_o2;
  assign new_n2497_ = ~n4005_o2;
  assign new_n2498_ = n4006_o2;
  assign new_n2499_ = ~n4006_o2;
  assign new_n2501_ = ~n1445_inv;
  assign new_n2502_ = n2176_o2;
  assign new_n2504_ = n2227_o2;
  assign new_n2506_ = n2236_o2;
  assign new_n2508_ = n2245_o2;
  assign new_n2510_ = n2518_o2;
  assign new_n2511_ = ~n2518_o2;
  assign new_n2512_ = n4023_o2;
  assign new_n2514_ = n1466_inv;
  assign new_n2516_ = n4038_o2;
  assign new_n2517_ = ~n4038_o2;
  assign new_n2518_ = n4039_o2;
  assign new_n2519_ = ~n4039_o2;
  assign new_n2520_ = n1475_inv;
  assign new_n2521_ = ~n1475_inv;
  assign new_n2523_ = ~n2119_o2;
  assign new_n2524_ = n2275_o2;
  assign new_n2525_ = ~n2275_o2;
  assign new_n2526_ = n2595_o2;
  assign new_n2527_ = ~n2595_o2;
  assign new_n2528_ = n2594_o2;
  assign new_n2529_ = ~n2594_o2;
  assign new_n2530_ = lo498_buf_o2;
  assign new_n2531_ = ~lo498_buf_o2;
  assign new_n2532_ = lo502_buf_o2;
  assign new_n2533_ = ~lo502_buf_o2;
  assign new_n2534_ = lo550_buf_o2;
  assign new_n2535_ = ~lo550_buf_o2;
  assign new_n2536_ = n2596_o2;
  assign new_n2537_ = ~n2596_o2;
  assign new_n2538_ = n2593_o2;
  assign new_n2541_ = ~n2668_o2;
  assign new_n2542_ = lo542_buf_o2;
  assign new_n2543_ = ~lo542_buf_o2;
  assign new_n2544_ = n2667_o2;
  assign new_n2546_ = n2404_o2;
  assign new_n2548_ = n2410_o2;
  assign new_n2551_ = ~n2419_o2;
  assign new_n2552_ = n2392_o2;
  assign new_n2555_ = ~n2369_o2;
  assign new_n2557_ = ~n2397_o2;
  assign new_n2559_ = ~n2601_o2;
  assign new_n2561_ = ~n2658_o2;
  assign new_n2562_ = n2574_o2;
  assign new_n2563_ = ~n2574_o2;
  assign new_n2564_ = n2205_o2;
  assign new_n2565_ = ~n2205_o2;
  assign new_n2566_ = lo510_buf_o2;
  assign new_n2567_ = ~lo510_buf_o2;
  assign new_n2568_ = lo514_buf_o2;
  assign new_n2569_ = ~lo514_buf_o2;
  assign new_n2570_ = lo554_buf_o2;
  assign new_n2571_ = ~lo554_buf_o2;
  assign new_n2572_ = lo558_buf_o2;
  assign new_n2573_ = ~lo558_buf_o2;
  assign new_n2574_ = lo578_buf_o2;
  assign new_n2575_ = ~lo578_buf_o2;
  assign new_n2576_ = n2254_o2;
  assign new_n2577_ = ~n2254_o2;
  assign new_n2579_ = ~n2421_o2;
  assign new_n2581_ = ~n2422_o2;
  assign new_n2583_ = ~n2130_o2;
  assign new_n2585_ = ~n2127_o2;
  assign new_n2587_ = ~n2131_o2;
  assign new_n2589_ = ~n2128_o2;
  assign new_n2590_ = n2264_o2;
  assign new_n2591_ = ~n2264_o2;
  assign new_n2592_ = n2467_o2;
  assign new_n2594_ = n2471_o2;
  assign new_n2596_ = n2488_o2;
  assign new_n2598_ = n2478_o2;
  assign new_n2600_ = n2486_o2;
  assign new_n2602_ = n2485_o2;
  assign new_n2604_ = n2498_o2;
  assign new_n2606_ = n2495_o2;
  assign new_n2608_ = n2496_o2;
  assign new_n2610_ = n2458_o2;
  assign new_n2612_ = n2643_o2;
  assign new_n2613_ = ~n2643_o2;
  assign new_n2614_ = n2462_o2;
  assign new_n2616_ = n2468_o2;
  assign new_n2618_ = n2639_o2;
  assign new_n2619_ = ~n2639_o2;
  assign new_n2620_ = n2499_o2;
  assign new_n2622_ = n2472_o2;
  assign new_n2624_ = n2474_o2;
  assign new_n2626_ = n2489_o2;
  assign new_n2628_ = n2321_o2;
  assign new_n2629_ = ~n2321_o2;
  assign new_n2630_ = n2322_o2;
  assign new_n2631_ = ~n2322_o2;
  assign new_n2632_ = n2640_o2;
  assign new_n2634_ = n2642_o2;
  assign new_n2636_ = n2187_o2;
  assign new_n2637_ = ~n2187_o2;
  assign new_n2638_ = n2373_o2;
  assign new_n2639_ = ~n2373_o2;
  assign new_n2640_ = n2603_o2;
  assign new_n2642_ = n2388_o2;
  assign new_n2643_ = ~n2388_o2;
  assign new_n2644_ = n2437_o2;
  assign new_n2645_ = ~n2437_o2;
  assign new_n2646_ = n2356_o2;
  assign new_n2647_ = ~n2356_o2;
  assign new_n2648_ = n2452_o2;
  assign new_n2649_ = ~n2452_o2;
  assign new_n2650_ = n2347_o2;
  assign new_n2651_ = ~n2347_o2;
  assign new_n2652_ = n2329_o2;
  assign new_n2653_ = ~n2329_o2;
  assign new_n2654_ = n2669_o2;
  assign new_n2655_ = ~n2669_o2;
  assign new_n2656_ = n2332_o2;
  assign new_n2657_ = ~n2332_o2;
  assign new_n2658_ = n2664_o2;
  assign new_n2659_ = ~n2664_o2;
  assign new_n2660_ = n2665_o2;
  assign new_n2662_ = n2653_o2;
  assign new_n2663_ = ~n2653_o2;
  assign new_n2664_ = n2654_o2;
  assign new_n2666_ = n2636_o2;
  assign new_n2668_ = n2660_o2;
  assign new_n2670_ = n2318_o2;
  assign new_n2671_ = ~n2318_o2;
  assign new_n2672_ = n2319_o2;
  assign new_n2673_ = ~n2319_o2;
  assign new_n2674_ = n2586_o2;
  assign new_n2675_ = ~n2586_o2;
  assign new_n2676_ = n2587_o2;
  assign new_n2677_ = ~n2587_o2;
  assign new_n2678_ = n2288_o2;
  assign new_n2679_ = ~n2288_o2;
  assign new_n2680_ = n2344_o2;
  assign new_n2681_ = ~n2344_o2;
  assign new_n2682_ = n2530_o2;
  assign new_n2683_ = ~n2530_o2;
  assign new_n2684_ = n2303_o2;
  assign new_n2685_ = ~n2303_o2;
  assign new_n2686_ = n2566_o2;
  assign new_n2687_ = ~n2566_o2;
  assign new_n2688_ = n2567_o2;
  assign new_n2689_ = ~n2567_o2;
  assign new_n2690_ = n2554_o2;
  assign new_n2691_ = ~n2554_o2;
  assign new_n2692_ = n2194_o2;
  assign new_n2693_ = ~n2194_o2;
  assign new_n2694_ = lo582_buf_o2;
  assign new_n2695_ = ~lo582_buf_o2;
  assign new_n2696_ = lo030_buf_o2;
  assign new_n2697_ = ~lo030_buf_o2;
  assign new_n2698_ = lo174_buf_o2;
  assign new_n2699_ = ~lo174_buf_o2;
  assign new_n2700_ = lo178_buf_o2;
  assign new_n2701_ = ~lo178_buf_o2;
  assign new_n2702_ = lo186_buf_o2;
  assign new_n2703_ = ~lo186_buf_o2;
  assign new_n2704_ = lo266_buf_o2;
  assign new_n2705_ = ~lo266_buf_o2;
  assign new_n2706_ = lo306_buf_o2;
  assign new_n2707_ = ~lo306_buf_o2;
  assign new_n2708_ = lo346_buf_o2;
  assign new_n2709_ = ~lo346_buf_o2;
  assign new_n2710_ = lo386_buf_o2;
  assign new_n2711_ = ~lo386_buf_o2;
  assign new_n2712_ = lo426_buf_o2;
  assign new_n2713_ = ~lo426_buf_o2;
  assign new_n2714_ = lo590_buf_o2;
  assign new_n2715_ = ~lo590_buf_o2;
  assign new_n2716_ = lo594_buf_o2;
  assign new_n2717_ = ~lo594_buf_o2;
  assign new_n2718_ = lo606_buf_o2;
  assign new_n2719_ = ~lo606_buf_o2;
  assign new_n2720_ = lo610_buf_o2;
  assign new_n2721_ = ~lo610_buf_o2;
  assign new_n2722_ = n2238_o2;
  assign new_n2723_ = ~n2238_o2;
  assign new_n2724_ = n2229_o2;
  assign new_n2725_ = ~n2229_o2;
  assign new_n2726_ = n2242_o2;
  assign new_n2727_ = ~n2242_o2;
  assign new_n2728_ = n2233_o2;
  assign new_n2729_ = ~n2233_o2;
  assign new_n2730_ = n2168_o2;
  assign new_n2731_ = ~n2168_o2;
  assign new_n2732_ = n2237_o2;
  assign new_n2733_ = ~n2237_o2;
  assign new_n2734_ = n2228_o2;
  assign new_n2735_ = ~n2228_o2;
  assign new_n2736_ = n2172_o2;
  assign new_n2737_ = ~n2172_o2;
  assign new_n2738_ = n2223_o2;
  assign new_n2739_ = ~n2223_o2;
  assign new_n2740_ = n2222_o2;
  assign new_n2741_ = ~n2222_o2;
  assign new_n2742_ = n2170_o2;
  assign new_n2743_ = ~n2170_o2;
  assign new_n2744_ = n2181_o2;
  assign new_n2745_ = ~n2181_o2;
  assign new_n2746_ = n2510_o2;
  assign new_n2747_ = ~n2510_o2;
  assign new_n2749_ = ~n2621_o2;
  assign new_n2750_ = lo466_buf_o2;
  assign new_n2751_ = ~lo466_buf_o2;
  assign new_n2752_ = lo478_buf_o2;
  assign new_n2753_ = ~lo478_buf_o2;
  assign new_n2754_ = n2149_o2;
  assign new_n2755_ = ~n2149_o2;
  assign new_n2756_ = n2429_o2;
  assign new_n2757_ = ~n2429_o2;
  assign new_n2758_ = n2444_o2;
  assign new_n2759_ = ~n2444_o2;
  assign new_n2760_ = n2153_o2;
  assign new_n2761_ = ~n2153_o2;
  assign new_n2762_ = n2433_o2;
  assign new_n2763_ = ~n2433_o2;
  assign new_n2764_ = n2448_o2;
  assign new_n2765_ = ~n2448_o2;
  assign new_n2766_ = n2367_o2;
  assign new_n2767_ = ~n2367_o2;
  assign new_n2768_ = n2386_o2;
  assign new_n2769_ = ~n2386_o2;
  assign new_n2770_ = n2539_o2;
  assign new_n2771_ = ~n2539_o2;
  assign new_n2772_ = n2183_o2;
  assign new_n2773_ = ~n2183_o2;
  assign new_n2774_ = n2220_o2;
  assign new_n2775_ = ~n2220_o2;
  assign new_n2776_ = n2514_o2;
  assign new_n2777_ = ~n2514_o2;
  assign new_n2778_ = n2196_o2;
  assign new_n2781_ = ~n2616_o2;
  assign new_n2783_ = ~n2612_o2;
  assign new_n2785_ = ~n2627_o2;
  assign new_n2786_ = n2140_o2;
  assign new_n2788_ = n1877_inv;
  assign new_n2791_ = ~lo149_buf_o2;
  assign new_n2792_ = lo197_buf_o2;
  assign new_n2794_ = lo118_buf_o2;
  assign new_n2795_ = ~lo118_buf_o2;
  assign new_n2796_ = lo158_buf_o2;
  assign new_n2798_ = lo166_buf_o2;
  assign new_n2800_ = lo242_buf_o2;
  assign new_n2802_ = lo286_buf_o2;
  assign new_n2804_ = lo506_buf_o2;
  assign new_n2805_ = ~lo506_buf_o2;
  assign new_n2806_ = n2198_o2;
  assign new_n2808_ = n2202_o2;
  assign new_n2810_ = n2197_o2;
  assign new_n2812_ = n1913_inv;
  assign new_n2813_ = ~n1913_inv;
  assign new_n2814_ = n2146_o2;
  assign new_n2815_ = ~n2146_o2;
  assign new_n2816_ = n1919_inv;
  assign new_n2817_ = ~n1919_inv;
  assign new_n2819_ = ~lo312_buf_o2;
  assign new_n2820_ = lo316_buf_o2;
  assign new_n2823_ = ~lo352_buf_o2;
  assign new_n2824_ = lo356_buf_o2;
  assign new_n2827_ = ~lo392_buf_o2;
  assign new_n2828_ = lo396_buf_o2;
  assign new_n2831_ = ~lo432_buf_o2;
  assign new_n2832_ = lo436_buf_o2;
  assign new_n2834_ = lo576_buf_o2;
  assign new_n2835_ = ~lo576_buf_o2;
  assign new_n2836_ = new_n2523_ | new_n2489_;
  assign new_n2837_ = new_n1763_ | new_n1701_;
  assign new_n2838_ = new_n2837_ | new_n4161_;
  assign new_n2839_ = new_n4163_ & new_n2056_;
  assign new_n2840_ = new_n4161_ | new_n1735_;
  assign new_n2841_ = new_n4166_ | new_n2235_;
  assign new_n2842_ = new_n4166_ | new_n2407_;
  assign new_n2843_ = new_n2589_ | new_n2585_;
  assign new_n2844_ = new_n2587_ | new_n2583_;
  assign new_n2845_ = new_n4167_ | new_n4168_;
  assign new_n2846_ = new_n4167_ & new_n2406_;
  assign new_n2847_ = new_n4168_ & new_n2234_;
  assign new_n2848_ = new_n2847_ | new_n2846_;
  assign new_n2849_ = new_n2463_ & new_n2461_;
  assign new_n2850_ = new_n2479_ & new_n2477_;
  assign new_n2851_ = new_n2493_ & new_n2487_;
  assign new_n2852_ = new_n2480_ | new_n2474_;
  assign new_n2853_ = new_n2466_ | new_n4170_;
  assign new_n2854_ = new_n2244_ | new_n2217_;
  assign new_n2855_ = new_n2854_ | new_n4172_;
  assign new_n2856_ = new_n4173_ | new_n1867_;
  assign new_n2857_ = new_n1708_ & new_n1692_;
  assign new_n2858_ = new_n2857_ | new_n4173_;
  assign new_n2859_ = new_n4174_ | new_n4176_;
  assign new_n2860_ = new_n4178_ | new_n4180_;
  assign new_n2861_ = new_n2860_ & new_n2859_;
  assign new_n2862_ = new_n2473_ & new_n4180_;
  assign new_n2863_ = new_n4182_ & new_n4176_;
  assign new_n2864_ = new_n2863_ | new_n2862_;
  assign new_n2865_ = new_n4170_ & new_n4183_;
  assign new_n2866_ = new_n2865_ | new_n4184_;
  assign new_n2867_ = new_n2467_ | new_n4177_;
  assign new_n2868_ = new_n4186_ | new_n4181_;
  assign new_n2869_ = new_n2868_ & new_n2867_;
  assign new_n2870_ = new_n2525_ | new_n2388_;
  assign new_n2871_ = new_n2524_ | new_n2389_;
  assign new_n2872_ = new_n2871_ & new_n2870_;
  assign new_n2873_ = new_n2872_ | new_n2396_;
  assign new_n2874_ = new_n2685_ | new_n2679_;
  assign new_n2875_ = new_n2684_ | new_n2678_;
  assign new_n2876_ = new_n2875_ & new_n1754_;
  assign new_n2877_ = new_n2876_ & new_n2874_;
  assign new_n2878_ = new_n2673_ & new_n2671_;
  assign new_n2879_ = new_n2672_ | new_n2670_;
  assign new_n2880_ = new_n2631_ & new_n2629_;
  assign new_n2881_ = new_n2630_ | new_n2628_;
  assign new_n2882_ = new_n2880_ | new_n2879_;
  assign new_n2883_ = new_n2881_ | new_n2878_;
  assign new_n2884_ = new_n2883_ & new_n2882_;
  assign new_n2885_ = new_n4187_ & new_n4188_;
  assign new_n2886_ = new_n4189_ | new_n4190_;
  assign new_n2887_ = new_n4189_ & new_n4190_;
  assign new_n2888_ = new_n4187_ | new_n4188_;
  assign new_n2889_ = new_n2888_ & new_n2886_;
  assign new_n2890_ = new_n2887_ | new_n2885_;
  assign new_n2891_ = new_n4191_ & new_n4192_;
  assign new_n2892_ = new_n4193_ | new_n4194_;
  assign new_n2893_ = new_n4193_ & new_n4194_;
  assign new_n2894_ = new_n4191_ | new_n4192_;
  assign new_n2895_ = new_n2894_ & new_n2892_;
  assign new_n2896_ = new_n2893_ | new_n2891_;
  assign new_n2897_ = new_n2896_ | new_n2889_;
  assign new_n2898_ = new_n2895_ | new_n2890_;
  assign new_n2899_ = new_n2898_ & new_n2897_;
  assign new_n2900_ = new_n2646_ & new_n2381_;
  assign new_n2901_ = new_n2555_ & new_n2358_;
  assign new_n2902_ = new_n2638_ & new_n2291_;
  assign new_n2903_ = new_n2902_ | new_n2901_;
  assign new_n2904_ = new_n2903_ | new_n2900_;
  assign new_n2905_ = new_n2643_ & new_n2332_;
  assign new_n2906_ = new_n2552_ & new_n2365_;
  assign new_n2907_ = new_n2906_ | new_n2905_;
  assign new_n2908_ = new_n2557_ & new_n2372_;
  assign new_n2909_ = new_n2642_ & new_n2333_;
  assign new_n2910_ = new_n2909_ | new_n2908_;
  assign new_n2911_ = new_n2910_ | new_n2907_;
  assign new_n2912_ = new_n2546_ & new_n2279_;
  assign new_n2913_ = new_n2639_ & new_n2290_;
  assign new_n2914_ = new_n2913_ | new_n2912_;
  assign new_n2915_ = new_n2548_ & new_n2325_;
  assign new_n2916_ = new_n2647_ & new_n2380_;
  assign new_n2917_ = new_n2916_ | new_n2915_;
  assign new_n2918_ = new_n2917_ | new_n2914_;
  assign new_n2919_ = new_n2918_ | new_n2911_;
  assign new_n2920_ = new_n2919_ | new_n2904_;
  assign new_n2921_ = new_n2551_ & new_n2310_;
  assign new_n2922_ = new_n2581_ & new_n2579_;
  assign new_n2923_ = new_n2922_ | new_n1747_;
  assign new_n2924_ = new_n2923_ | new_n2921_;
  assign new_n2925_ = new_n2644_ & new_n2353_;
  assign new_n2926_ = new_n2645_ & new_n2352_;
  assign new_n2927_ = new_n2926_ | new_n2925_;
  assign new_n2928_ = new_n2649_ & new_n2338_;
  assign new_n2929_ = new_n2648_ & new_n2339_;
  assign new_n2930_ = new_n2929_ | new_n2928_;
  assign new_n2931_ = new_n2930_ | new_n2927_;
  assign new_n2932_ = new_n2931_ | new_n2924_;
  assign new_n2933_ = new_n2614_ | new_n2610_;
  assign new_n2934_ = new_n2616_ | new_n2592_;
  assign new_n2935_ = new_n2934_ | new_n2933_;
  assign new_n2936_ = new_n2622_ | new_n2594_;
  assign new_n2937_ = new_n2624_ | new_n2598_;
  assign new_n2938_ = new_n2937_ | new_n2936_;
  assign new_n2939_ = new_n2938_ | new_n2935_;
  assign new_n2940_ = new_n2602_ | new_n2600_;
  assign new_n2941_ = new_n2626_ | new_n2596_;
  assign new_n2942_ = new_n2941_ | new_n2940_;
  assign new_n2943_ = new_n2608_ | new_n2606_;
  assign new_n2944_ = new_n2620_ | new_n2604_;
  assign new_n2945_ = new_n2944_ | new_n2943_;
  assign new_n2946_ = new_n2945_ | new_n2942_;
  assign new_n2947_ = new_n2946_ | new_n2939_;
  assign new_n2948_ = new_n2947_ | new_n2932_;
  assign new_n2949_ = new_n2948_ | new_n2920_;
  assign new_n2950_ = new_n4174_ & new_n4183_;
  assign new_n2951_ = new_n4184_ | new_n2227_;
  assign new_n2952_ = new_n2950_ & new_n2511_;
  assign new_n2953_ = new_n2951_ & new_n2510_;
  assign new_n2954_ = new_n2953_ | new_n2952_;
  assign new_n2955_ = new_n2954_ & new_n4169_;
  assign new_n2956_ = new_n4195_ & new_n2252_;
  assign new_n2957_ = new_n2956_ | new_n2955_;
  assign new_n2958_ = new_n2690_ | new_n2682_;
  assign new_n2959_ = new_n2691_ | new_n2683_;
  assign new_n2960_ = new_n2959_ & new_n4196_;
  assign new_n2961_ = new_n2960_ & new_n2958_;
  assign new_n2962_ = new_n4195_ | new_n4177_;
  assign new_n2963_ = new_n2689_ & new_n2687_;
  assign new_n2964_ = new_n2688_ | new_n2686_;
  assign new_n2965_ = new_n4197_ & new_n4198_;
  assign new_n2966_ = new_n4186_ | new_n4199_;
  assign new_n2967_ = new_n4185_ & new_n4199_;
  assign new_n2968_ = new_n4197_ | new_n4198_;
  assign new_n2969_ = new_n2968_ & new_n2966_;
  assign new_n2970_ = new_n2967_ | new_n2965_;
  assign new_n2971_ = new_n2969_ | new_n4200_;
  assign new_n2972_ = new_n2970_ | new_n4201_;
  assign new_n2973_ = new_n2972_ & new_n2971_;
  assign new_n2974_ = new_n2973_ | new_n4181_;
  assign new_n2975_ = new_n2974_ & new_n2962_;
  assign new_n2976_ = new_n2677_ & new_n2674_;
  assign new_n2977_ = new_n2676_ | new_n2675_;
  assign new_n2978_ = new_n2977_ | new_n4200_;
  assign new_n2979_ = new_n2976_ | new_n4201_;
  assign new_n2980_ = new_n2979_ & new_n4196_;
  assign new_n2981_ = new_n2980_ & new_n2978_;
  assign new_n2982_ = new_n2559_ | new_n2538_;
  assign new_n2983_ = new_n2666_ | new_n2640_;
  assign new_n2984_ = new_n2983_ & new_n2982_;
  assign new_n2985_ = new_n2632_ | new_n2618_;
  assign new_n2986_ = new_n2634_ | new_n2612_;
  assign new_n2987_ = new_n2986_ | new_n4202_;
  assign new_n2988_ = new_n2987_ | new_n2984_;
  assign new_n2989_ = new_n4202_ | new_n2613_;
  assign new_n2990_ = new_n2989_ & new_n2619_;
  assign new_n2991_ = new_n2990_ & new_n2988_;
  assign new_n2992_ = new_n2664_ | new_n2662_;
  assign new_n2993_ = new_n4203_ | new_n4204_;
  assign new_n2994_ = new_n2660_ | new_n2658_;
  assign new_n2995_ = new_n2544_ & new_n2541_;
  assign new_n2996_ = new_n2995_ | new_n2654_;
  assign new_n2997_ = new_n2996_ | new_n4205_;
  assign new_n2998_ = new_n2997_ | new_n4206_;
  assign new_n2999_ = new_n2998_ | new_n2991_;
  assign new_n3000_ = new_n4204_ | new_n2655_;
  assign new_n3001_ = new_n3000_ | new_n4205_;
  assign new_n3002_ = new_n3001_ & new_n2561_;
  assign new_n3003_ = new_n3002_ | new_n4203_;
  assign new_n3004_ = new_n4206_ | new_n2659_;
  assign new_n3005_ = new_n3004_ & new_n2663_;
  assign new_n3006_ = new_n3005_ & new_n3003_;
  assign new_n3007_ = new_n3006_ & new_n2999_;
  assign new_n3008_ = new_n4207_ | new_n4208_;
  assign new_n3009_ = new_n3008_ | new_n4209_;
  assign new_n3010_ = new_n4210_ | new_n4172_;
  assign new_n3011_ = new_n3010_ | new_n4211_;
  assign new_n3012_ = new_n3011_ | new_n3009_;
  assign new_n3013_ = new_n2702_ & new_n4213_;
  assign new_n3014_ = new_n2703_ | new_n4216_;
  assign new_n3015_ = new_n2754_ & new_n4220_;
  assign new_n3016_ = new_n2755_ | new_n4227_;
  assign new_n3017_ = new_n2760_ & new_n4227_;
  assign new_n3018_ = new_n2761_ | new_n4220_;
  assign new_n3019_ = new_n2773_ & new_n2744_;
  assign new_n3020_ = new_n2772_ | new_n2745_;
  assign new_n3021_ = new_n2777_ & new_n2747_;
  assign new_n3022_ = new_n2776_ | new_n2746_;
  assign new_n3023_ = new_n4213_ & new_n1942_;
  assign new_n3024_ = new_n4216_ | new_n1943_;
  assign new_n3025_ = new_n4233_ & new_n4235_;
  assign new_n3026_ = new_n4237_ | new_n4239_;
  assign new_n3027_ = new_n3020_ & new_n3014_;
  assign new_n3028_ = new_n4240_ | new_n4241_;
  assign new_n3029_ = new_n2731_ & new_n4244_;
  assign new_n3030_ = new_n2730_ | new_n4249_;
  assign new_n3031_ = new_n2743_ & new_n2737_;
  assign new_n3032_ = new_n2742_ | new_n2736_;
  assign new_n3033_ = new_n3031_ & new_n3030_;
  assign new_n3034_ = new_n3032_ | new_n3029_;
  assign new_n3035_ = new_n2693_ & new_n2637_;
  assign new_n3036_ = new_n2692_ | new_n2636_;
  assign new_n3037_ = new_n3034_ & new_n3024_;
  assign new_n3038_ = new_n4252_ | new_n4253_;
  assign new_n3039_ = new_n2740_ & new_n2739_;
  assign new_n3040_ = new_n2741_ | new_n2738_;
  assign new_n3041_ = new_n3040_ & new_n4254_;
  assign new_n3042_ = new_n3039_ | new_n4255_;
  assign new_n3043_ = new_n2705_ & new_n4249_;
  assign new_n3044_ = new_n2704_ | new_n4244_;
  assign new_n3045_ = new_n3043_ & new_n4255_;
  assign new_n3046_ = new_n3044_ | new_n4254_;
  assign new_n3047_ = new_n3046_ & new_n3042_;
  assign new_n3048_ = new_n3045_ | new_n3041_;
  assign new_n3049_ = new_n2735_ & new_n2725_;
  assign new_n3050_ = new_n2734_ | new_n2724_;
  assign new_n3051_ = new_n3050_ & new_n4250_;
  assign new_n3052_ = new_n3049_ | new_n4245_;
  assign new_n3053_ = new_n2700_ & new_n4214_;
  assign new_n3054_ = new_n2701_ | new_n4217_;
  assign new_n3055_ = new_n2728_ & new_n4245_;
  assign new_n3056_ = new_n2729_ | new_n4250_;
  assign new_n3057_ = new_n3056_ & new_n3054_;
  assign new_n3058_ = new_n3055_ | new_n3053_;
  assign new_n3059_ = new_n3057_ & new_n3052_;
  assign new_n3060_ = new_n3058_ | new_n3051_;
  assign new_n3061_ = new_n2733_ & new_n2723_;
  assign new_n3062_ = new_n2732_ | new_n2722_;
  assign new_n3063_ = new_n3062_ & new_n4251_;
  assign new_n3064_ = new_n3061_ | new_n4246_;
  assign new_n3065_ = new_n2698_ & new_n4214_;
  assign new_n3066_ = new_n2699_ | new_n4217_;
  assign new_n3067_ = new_n2726_ & new_n4246_;
  assign new_n3068_ = new_n2727_ | new_n4251_;
  assign new_n3069_ = new_n3068_ & new_n3066_;
  assign new_n3070_ = new_n3067_ | new_n3065_;
  assign new_n3071_ = new_n3069_ & new_n3064_;
  assign new_n3072_ = new_n3070_ | new_n3063_;
  assign new_n3073_ = new_n4257_ & new_n4258_;
  assign new_n3074_ = new_n4259_ | new_n4261_;
  assign new_n3075_ = new_n4259_ & new_n4261_;
  assign new_n3076_ = new_n4257_ | new_n4258_;
  assign new_n3077_ = new_n3076_ & new_n3074_;
  assign new_n3078_ = new_n3075_ | new_n3073_;
  assign new_n3079_ = new_n4263_ | new_n4265_;
  assign new_n3080_ = new_n2706_ & new_n4267_;
  assign new_n3081_ = new_n2707_ | new_n4270_;
  assign new_n3082_ = new_n2712_ & new_n4270_;
  assign new_n3083_ = new_n2713_ | new_n4267_;
  assign new_n3084_ = new_n3083_ & new_n3081_;
  assign new_n3085_ = new_n3082_ | new_n3080_;
  assign new_n3086_ = new_n3085_ & new_n4221_;
  assign new_n3087_ = new_n3084_ | new_n4228_;
  assign new_n3088_ = new_n2708_ & new_n4268_;
  assign new_n3089_ = new_n2709_ | new_n4271_;
  assign new_n3090_ = new_n2710_ & new_n4271_;
  assign new_n3091_ = new_n2711_ | new_n4268_;
  assign new_n3092_ = new_n3091_ & new_n3089_;
  assign new_n3093_ = new_n3090_ | new_n3088_;
  assign new_n3094_ = new_n3093_ & new_n4228_;
  assign new_n3095_ = new_n3092_ | new_n4221_;
  assign new_n3096_ = new_n3095_ & new_n3087_;
  assign new_n3097_ = new_n3094_ | new_n3086_;
  assign new_n3098_ = new_n2815_ & new_n2794_;
  assign new_n3099_ = new_n4272_ | new_n2795_;
  assign new_n3100_ = new_n4273_ & new_n2805_;
  assign new_n3101_ = new_n2817_ | new_n2804_;
  assign new_n3102_ = new_n4274_ & new_n4275_;
  assign new_n3103_ = new_n3101_ | new_n3099_;
  assign new_n3104_ = new_n4277_ | new_n4279_;
  assign new_n3105_ = new_n2529_ & new_n2526_;
  assign new_n3106_ = new_n2528_ | new_n2527_;
  assign new_n3107_ = new_n4282_ | new_n4285_;
  assign new_n3108_ = new_n4288_ & new_n4290_;
  assign new_n3109_ = new_n4294_ & new_n1714_;
  assign new_n3110_ = new_n4301_ & new_n4306_;
  assign new_n3111_ = new_n3110_ | new_n3109_;
  assign new_n3112_ = new_n1804_ & new_n4294_;
  assign new_n3113_ = new_n4312_ & new_n4306_;
  assign new_n3114_ = new_n3113_ | new_n3112_;
  assign new_n3115_ = new_n1798_ & new_n4293_;
  assign new_n3116_ = new_n4314_ & new_n4305_;
  assign new_n3117_ = new_n3116_ | new_n3115_;
  assign new_n3118_ = new_n4317_ & new_n1822_;
  assign new_n3119_ = new_n4323_ & new_n4327_;
  assign new_n3120_ = new_n3119_ | new_n3118_;
  assign new_n3121_ = new_n1846_ & new_n4317_;
  assign new_n3122_ = new_n4333_ & new_n4327_;
  assign new_n3123_ = new_n3122_ | new_n3121_;
  assign new_n3124_ = new_n1852_ & new_n4318_;
  assign new_n3125_ = new_n4335_ & new_n4328_;
  assign new_n3126_ = new_n3125_ | new_n3124_;
  assign new_n3127_ = new_n4336_ & new_n2537_;
  assign new_n3128_ = new_n4338_ & new_n4342_;
  assign new_n3129_ = new_n4336_ & new_n2536_;
  assign new_n3130_ = new_n4345_ & new_n4263_;
  assign new_n3131_ = new_n3130_ | new_n3128_;
  assign new_n3132_ = new_n2758_ & new_n4223_;
  assign new_n3133_ = new_n2759_ | new_n4230_;
  assign new_n3134_ = new_n2764_ & new_n4230_;
  assign new_n3135_ = new_n2765_ | new_n4223_;
  assign new_n3136_ = new_n3135_ & new_n3133_;
  assign new_n3137_ = new_n3134_ | new_n3132_;
  assign new_n3138_ = new_n4348_ & new_n4288_;
  assign new_n3139_ = new_n4351_ | new_n4282_;
  assign new_n3140_ = new_n4287_ & new_n4352_;
  assign new_n3141_ = new_n4281_ | new_n4354_;
  assign new_n3142_ = new_n3141_ | new_n3138_;
  assign new_n3143_ = new_n4357_ & new_n4301_;
  assign new_n3144_ = new_n4360_ | new_n4361_;
  assign new_n3145_ = new_n4360_ & new_n4361_;
  assign new_n3146_ = new_n4357_ | new_n4300_;
  assign new_n3147_ = new_n3146_ & new_n3144_;
  assign new_n3148_ = new_n3145_ | new_n3143_;
  assign new_n3149_ = new_n3147_ & new_n4362_;
  assign new_n3150_ = new_n3148_ & new_n3077_;
  assign new_n3151_ = new_n3150_ | new_n3149_;
  assign new_n3152_ = new_n2810_ | new_n2806_;
  assign new_n3153_ = new_n3152_ & new_n4366_;
  assign new_n3154_ = new_n4375_ & new_n2798_;
  assign new_n3155_ = new_n2808_ & new_n4379_;
  assign new_n3156_ = new_n3155_ | new_n3154_;
  assign new_n3157_ = new_n3156_ | new_n3153_;
  assign new_n3158_ = new_n2802_ & new_n4384_;
  assign new_n3159_ = new_n2796_ & new_n4393_;
  assign new_n3160_ = new_n3159_ | new_n3158_;
  assign new_n3161_ = new_n3160_ & new_n4366_;
  assign new_n3162_ = new_n4375_ & new_n2792_;
  assign new_n3163_ = new_n2800_ & new_n4393_;
  assign new_n3164_ = new_n3163_ & new_n4379_;
  assign new_n3165_ = new_n3164_ | new_n3162_;
  assign new_n3166_ = new_n3165_ | new_n3161_;
  assign new_n3167_ = new_n4318_ & new_n1828_;
  assign new_n3168_ = new_n4405_ & new_n4328_;
  assign new_n3169_ = new_n4406_ & new_n4407_;
  assign new_n3170_ = new_n4408_ & new_n4409_;
  assign new_n3171_ = new_n4410_ & new_n4411_;
  assign new_n3172_ = new_n4412_ & new_n4413_;
  assign new_n3173_ = new_n4302_ | new_n4414_;
  assign new_n3174_ = new_n1774_ & new_n4295_;
  assign new_n3175_ = new_n4262_ & new_n4307_;
  assign new_n3176_ = new_n3175_ | new_n3174_;
  assign new_n3177_ = new_n4415_ | new_n4417_;
  assign new_n3178_ = new_n4415_ & new_n4417_;
  assign new_n3179_ = new_n4419_ | new_n4421_;
  assign new_n3180_ = new_n1780_ & new_n4295_;
  assign new_n3181_ = new_n4358_ & new_n4307_;
  assign new_n3182_ = new_n3181_ | new_n3180_;
  assign new_n3183_ = new_n4422_ | new_n4424_;
  assign new_n3184_ = new_n4422_ & new_n4424_;
  assign new_n3185_ = new_n1786_ & new_n4297_;
  assign new_n3186_ = new_n4427_ & new_n4309_;
  assign new_n3187_ = new_n3186_ | new_n3185_;
  assign new_n3188_ = new_n4429_ & new_n4431_;
  assign new_n3189_ = new_n4429_ | new_n4431_;
  assign new_n3190_ = new_n1792_ & new_n4297_;
  assign new_n3191_ = new_n4277_ & new_n4309_;
  assign new_n3192_ = new_n3191_ | new_n3190_;
  assign new_n3193_ = new_n4433_ & new_n4342_;
  assign new_n3194_ = new_n4433_ | new_n4341_;
  assign new_n3195_ = new_n4434_ & new_n4436_;
  assign new_n3196_ = new_n4338_ & new_n4436_;
  assign new_n3197_ = new_n4298_ & new_n1726_;
  assign new_n3198_ = new_n4439_ & new_n4310_;
  assign new_n3199_ = new_n3198_ | new_n3197_;
  assign new_n3200_ = new_n4440_ & new_n4442_;
  assign new_n3201_ = new_n4440_ | new_n4442_;
  assign new_n3202_ = new_n4339_ & new_n4443_;
  assign new_n3203_ = new_n4444_ | new_n4445_;
  assign new_n3204_ = new_n4446_ & new_n4239_;
  assign new_n3205_ = new_n4447_ | new_n4237_;
  assign new_n3206_ = new_n4448_ & new_n4265_;
  assign new_n3207_ = new_n2395_ & new_n4449_;
  assign new_n3208_ = new_n4450_ & new_n2387_;
  assign new_n3209_ = new_n4345_ & new_n4451_;
  assign new_n3210_ = new_n4346_ & new_n4452_;
  assign new_n3211_ = new_n2813_ | new_n1951_;
  assign new_n3212_ = new_n4298_ & new_n1720_;
  assign new_n3213_ = new_n4454_ & new_n4310_;
  assign new_n3214_ = new_n3213_ | new_n3212_;
  assign new_n3215_ = new_n4456_ | new_n4457_;
  assign new_n3216_ = new_n4320_ & new_n1810_;
  assign new_n3217_ = new_n4459_ & new_n4330_;
  assign new_n3218_ = new_n3217_ | new_n3216_;
  assign new_n3219_ = new_n4320_ & new_n1816_;
  assign new_n3220_ = new_n2756_ & new_n4224_;
  assign new_n3221_ = new_n2757_ | new_n4231_;
  assign new_n3222_ = new_n2762_ & new_n4231_;
  assign new_n3223_ = new_n2763_ | new_n4224_;
  assign new_n3224_ = new_n3223_ & new_n3221_;
  assign new_n3225_ = new_n3222_ | new_n3220_;
  assign new_n3226_ = new_n4461_ & new_n4330_;
  assign new_n3227_ = new_n3226_ | new_n3219_;
  assign new_n3228_ = new_n1858_ & new_n4321_;
  assign new_n3229_ = new_n3018_ & new_n3016_;
  assign new_n3230_ = new_n4463_ | new_n4464_;
  assign new_n3231_ = new_n4466_ & new_n4331_;
  assign new_n3232_ = new_n3231_ | new_n3228_;
  assign new_n3233_ = new_n1840_ & new_n4321_;
  assign new_n3234_ = new_n4348_ & new_n4331_;
  assign new_n3235_ = new_n3234_ | new_n3233_;
  assign new_n3236_ = new_n4467_ & new_n4432_;
  assign new_n3237_ = new_n2569_ & new_n2296_;
  assign new_n3238_ = new_n3237_ | new_n3236_;
  assign new_n3239_ = new_n4445_ & new_n2316_;
  assign new_n3240_ = new_n4285_ & new_n4443_;
  assign new_n3241_ = new_n3240_ | new_n3239_;
  assign new_n3242_ = new_n4468_ | new_n4469_;
  assign new_n3243_ = new_n4352_ & new_n4470_;
  assign new_n3244_ = new_n4354_ & new_n4471_;
  assign new_n3245_ = new_n3244_ | new_n3243_;
  assign new_n3246_ = new_n4283_ | new_n4473_;
  assign new_n3247_ = new_n4289_ & new_n4471_;
  assign new_n3248_ = new_n4474_ & new_n4475_;
  assign new_n3249_ = new_n4474_ | new_n4475_;
  assign new_n3250_ = new_n4461_ | new_n4283_;
  assign new_n3251_ = new_n4289_ & new_n4477_;
  assign new_n3252_ = new_n4478_ & new_n4479_;
  assign new_n3253_ = new_n4478_ | new_n4479_;
  assign new_n3254_ = new_n4427_ | new_n4279_;
  assign new_n3255_ = new_n4339_ & new_n4432_;
  assign new_n3256_ = new_n4346_ & new_n4264_;
  assign new_n3257_ = new_n3256_ | new_n3255_;
  assign new_n3258_ = new_n4480_ & new_n4481_;
  assign new_n3259_ = new_n4480_ | new_n4481_;
  assign new_n3260_ = new_n4482_ & new_n4454_;
  assign new_n3261_ = new_n4483_ & new_n4358_;
  assign new_n3262_ = new_n2785_ & new_n2749_;
  assign new_n3263_ = new_n3262_ | new_n3261_;
  assign new_n3264_ = new_n4482_ | new_n4455_;
  assign new_n3265_ = new_n4483_ | new_n4359_;
  assign new_n3266_ = new_n3265_ & new_n3264_;
  assign new_n3267_ = new_n3266_ & new_n3263_;
  assign new_n3268_ = new_n3267_ | new_n3260_;
  assign new_n3269_ = new_n3268_ & new_n3259_;
  assign new_n3270_ = new_n3269_ | new_n3258_;
  assign new_n3271_ = new_n3140_ | new_n3139_;
  assign new_n3272_ = new_n3271_ & new_n4484_;
  assign new_n3273_ = new_n4485_ | new_n4486_;
  assign new_n3274_ = new_n3273_ & new_n4487_;
  assign new_n3275_ = new_n4236_ & new_n4238_;
  assign new_n3276_ = new_n4233_ | new_n4235_;
  assign new_n3277_ = new_n3276_ & new_n3026_;
  assign new_n3278_ = new_n3275_ | new_n4488_;
  assign new_n3279_ = new_n4477_ & new_n4489_;
  assign new_n3280_ = new_n4491_ | new_n4492_;
  assign new_n3281_ = new_n4491_ & new_n4492_;
  assign new_n3282_ = new_n4476_ | new_n4489_;
  assign new_n3283_ = new_n3282_ & new_n3280_;
  assign new_n3284_ = new_n3281_ | new_n3279_;
  assign new_n3285_ = new_n3284_ | new_n3277_;
  assign new_n3286_ = new_n3283_ | new_n3278_;
  assign new_n3287_ = new_n3286_ & new_n3285_;
  assign new_n3288_ = new_n4493_ | new_n4494_;
  assign new_n3289_ = new_n4493_ & new_n4494_;
  assign new_n3290_ = new_n4495_ & new_n4428_;
  assign new_n3291_ = new_n3035_ & new_n3027_;
  assign new_n3292_ = new_n3291_ | new_n3290_;
  assign new_n3293_ = new_n4496_ & new_n4498_;
  assign new_n3294_ = new_n4496_ | new_n4498_;
  assign new_n3295_ = new_n4499_ & new_n4500_;
  assign new_n3296_ = new_n4501_ | new_n4502_;
  assign new_n3297_ = new_n4501_ & new_n4502_;
  assign new_n3298_ = new_n4499_ | new_n4500_;
  assign new_n3299_ = new_n3298_ & new_n3296_;
  assign new_n3300_ = new_n3297_ | new_n3295_;
  assign new_n3301_ = new_n4421_ & new_n4503_;
  assign new_n3302_ = new_n4505_ | new_n4418_;
  assign new_n3303_ = new_n4505_ & new_n4418_;
  assign new_n3304_ = new_n4420_ | new_n4503_;
  assign new_n3305_ = new_n3304_ & new_n3302_;
  assign new_n3306_ = new_n3303_ | new_n3301_;
  assign new_n3307_ = new_n3305_ & new_n3300_;
  assign new_n3308_ = new_n3306_ & new_n3299_;
  assign new_n3309_ = new_n3308_ | new_n3307_;
  assign new_n3310_ = new_n4437_ & new_n4506_;
  assign new_n3311_ = new_n4508_ | new_n4343_;
  assign new_n3312_ = new_n4508_ & new_n4343_;
  assign new_n3313_ = new_n4437_ | new_n4506_;
  assign new_n3314_ = new_n3313_ & new_n3311_;
  assign new_n3315_ = new_n3312_ | new_n3310_;
  assign new_n3316_ = new_n4425_ & new_n4509_;
  assign new_n3317_ = new_n4510_ | new_n4511_;
  assign new_n3318_ = new_n4510_ & new_n4511_;
  assign new_n3319_ = new_n4425_ | new_n4509_;
  assign new_n3320_ = new_n3319_ & new_n3317_;
  assign new_n3321_ = new_n3318_ | new_n3316_;
  assign new_n3322_ = new_n3320_ & new_n3314_;
  assign new_n3323_ = new_n3321_ & new_n3315_;
  assign new_n3324_ = new_n3323_ | new_n3322_;
  assign new_n3325_ = new_n4466_ & new_n4512_;
  assign new_n3326_ = new_n4513_ | new_n4335_;
  assign new_n3327_ = new_n4513_ & new_n4334_;
  assign new_n3328_ = new_n4465_ | new_n4512_;
  assign new_n3329_ = new_n3328_ & new_n3326_;
  assign new_n3330_ = new_n3327_ | new_n3325_;
  assign new_n3331_ = new_n3329_ | new_n3096_;
  assign new_n3332_ = new_n3330_ | new_n4405_;
  assign new_n3333_ = new_n3332_ & new_n3331_;
  assign new_n3334_ = new_n4514_ & new_n4515_;
  assign new_n3335_ = new_n4516_ | new_n4517_;
  assign new_n3336_ = new_n4516_ & new_n4517_;
  assign new_n3337_ = new_n4514_ | new_n4515_;
  assign new_n3338_ = new_n3337_ & new_n3335_;
  assign new_n3339_ = new_n3336_ | new_n3334_;
  assign new_n3340_ = new_n4518_ & new_n4519_;
  assign new_n3341_ = new_n4520_ | new_n4521_;
  assign new_n3342_ = new_n4520_ & new_n4521_;
  assign new_n3343_ = new_n4518_ | new_n4519_;
  assign new_n3344_ = new_n3343_ & new_n3341_;
  assign new_n3345_ = new_n3342_ | new_n3340_;
  assign new_n3346_ = new_n4522_ & new_n4523_;
  assign new_n3347_ = new_n4524_ | new_n4525_;
  assign new_n3348_ = new_n4524_ & new_n4525_;
  assign new_n3349_ = new_n4522_ | new_n4523_;
  assign new_n3350_ = new_n3349_ & new_n3347_;
  assign new_n3351_ = new_n3348_ | new_n3346_;
  assign new_n3352_ = new_n4526_ & new_n4527_;
  assign new_n3353_ = new_n4528_ | new_n4529_;
  assign new_n3354_ = new_n4528_ & new_n4529_;
  assign new_n3355_ = new_n4526_ | new_n4527_;
  assign new_n3356_ = new_n3355_ & new_n3353_;
  assign new_n3357_ = new_n3354_ | new_n3352_;
  assign new_n3358_ = new_n3357_ | new_n3350_;
  assign new_n3359_ = new_n3356_ | new_n3351_;
  assign new_n3360_ = new_n3359_ & new_n3358_;
  assign new_n3361_ = new_n4314_ & new_n3037_;
  assign new_n3362_ = new_n4452_ & new_n4278_;
  assign new_n3363_ = new_n3362_ | new_n3361_;
  assign new_n3364_ = new_n4290_ | new_n4439_;
  assign new_n3365_ = new_n4312_ | new_n4451_;
  assign new_n3366_ = new_n3365_ & new_n3364_;
  assign new_n3367_ = new_n4530_ & new_n4531_;
  assign new_n3368_ = new_n4530_ | new_n4531_;
  assign new_n3369_ = new_n4532_ & new_n4459_;
  assign new_n3370_ = new_n4533_ | new_n4473_;
  assign new_n3371_ = new_n4533_ & new_n4472_;
  assign new_n3372_ = new_n4532_ | new_n4458_;
  assign new_n3373_ = new_n3372_ & new_n3370_;
  assign new_n3374_ = new_n3371_ | new_n3369_;
  assign new_n3375_ = new_n4333_ & new_n4534_;
  assign new_n3376_ = new_n4535_ | new_n4323_;
  assign new_n3377_ = new_n4535_ & new_n4324_;
  assign new_n3378_ = new_n4332_ | new_n4534_;
  assign new_n3379_ = new_n3378_ & new_n3376_;
  assign new_n3380_ = new_n3377_ | new_n3375_;
  assign new_n3381_ = new_n4536_ & new_n4537_;
  assign new_n3382_ = new_n4538_ | new_n4539_;
  assign new_n3383_ = new_n4538_ & new_n4539_;
  assign new_n3384_ = new_n4536_ | new_n4537_;
  assign new_n3385_ = new_n3384_ & new_n3382_;
  assign new_n3386_ = new_n3383_ | new_n3381_;
  assign new_n3387_ = new_n4540_ & new_n4349_;
  assign new_n3388_ = new_n4462_ | new_n4351_;
  assign new_n3389_ = new_n4462_ & new_n4350_;
  assign new_n3390_ = new_n4540_ | new_n4349_;
  assign new_n3391_ = new_n3390_ & new_n3388_;
  assign new_n3392_ = new_n3389_ | new_n3387_;
  assign new_n3393_ = new_n3391_ & new_n3386_;
  assign new_n3394_ = new_n3392_ & new_n3385_;
  assign new_n3395_ = new_n3394_ | new_n3393_;
  assign new_n3396_ = new_n4384_ | new_n1995_;
  assign new_n3397_ = new_n3396_ & new_n4378_;
  assign new_n3398_ = new_n2791_ & new_n4394_;
  assign new_n3399_ = new_n3398_ & new_n4367_;
  assign new_n3400_ = new_n4385_ & new_n2039_;
  assign new_n3401_ = new_n3400_ | new_n3399_;
  assign new_n3402_ = new_n3401_ | new_n3397_;
  assign new_n3403_ = new_n4394_ & new_n1890_;
  assign new_n3404_ = new_n4396_ & new_n1894_;
  assign new_n3405_ = new_n4396_ & new_n1974_;
  assign new_n3406_ = new_n4397_ & new_n1978_;
  assign new_n3407_ = new_n4397_ & new_n1986_;
  assign new_n3408_ = new_n4385_ & new_n2018_;
  assign new_n3409_ = new_n4386_ & new_n2022_;
  assign new_n3410_ = new_n4386_ & new_n2031_;
  assign new_n3411_ = new_n4367_ & new_n1899_;
  assign new_n3412_ = new_n4369_ | new_n1982_;
  assign new_n3413_ = new_n4400_ & new_n1903_;
  assign new_n3414_ = new_n3413_ & new_n4369_;
  assign new_n3415_ = new_n4400_ & new_n1990_;
  assign new_n3416_ = new_n3415_ | new_n4368_;
  assign new_n3417_ = new_n4388_ & new_n2048_;
  assign new_n3418_ = new_n4401_ & new_n1918_;
  assign new_n3419_ = new_n3418_ | new_n3417_;
  assign new_n3420_ = new_n3419_ & new_n4371_;
  assign new_n3421_ = new_n4542_ | new_n4544_;
  assign new_n3422_ = new_n4547_ | new_n4549_;
  assign new_n3423_ = new_n3422_ & new_n3421_;
  assign new_n3424_ = new_n4550_ & new_n4552_;
  assign new_n3425_ = new_n4556_ & new_n2076_;
  assign new_n3426_ = new_n4567_ & new_n2184_;
  assign new_n3427_ = new_n3426_ | new_n3425_;
  assign new_n3428_ = new_n4556_ & new_n2084_;
  assign new_n3429_ = new_n4567_ & new_n2192_;
  assign new_n3430_ = new_n3429_ | new_n3428_;
  assign new_n3431_ = new_n4557_ & new_n2088_;
  assign new_n3432_ = new_n4568_ & new_n2196_;
  assign new_n3433_ = new_n3432_ | new_n3431_;
  assign new_n3434_ = new_n4557_ & new_n2112_;
  assign new_n3435_ = new_n4568_ & new_n2148_;
  assign new_n3436_ = new_n3435_ | new_n3434_;
  assign new_n3437_ = new_n4559_ & new_n2120_;
  assign new_n3438_ = new_n4570_ & new_n2156_;
  assign new_n3439_ = new_n3438_ | new_n3437_;
  assign new_n3440_ = new_n4559_ & new_n2124_;
  assign new_n3441_ = new_n4570_ & new_n2160_;
  assign new_n3442_ = new_n3441_ | new_n3440_;
  assign new_n3443_ = new_n4560_ & new_n2080_;
  assign new_n3444_ = new_n4571_ & new_n2188_;
  assign new_n3445_ = new_n3444_ | new_n3443_;
  assign new_n3446_ = new_n3445_ & new_n4577_;
  assign new_n3447_ = new_n4560_ & new_n2116_;
  assign new_n3448_ = new_n4571_ & new_n2152_;
  assign new_n3449_ = new_n3448_ | new_n3447_;
  assign new_n3450_ = new_n3449_ & new_n4580_;
  assign new_n3451_ = new_n3450_ | new_n3446_;
  assign new_n3452_ = new_n4562_ & new_n2060_;
  assign new_n3453_ = new_n4574_ & new_n2168_;
  assign new_n3454_ = new_n3453_ | new_n3452_;
  assign new_n3455_ = new_n3454_ & new_n4577_;
  assign new_n3456_ = new_n4562_ & new_n2096_;
  assign new_n3457_ = new_n4574_ & new_n2132_;
  assign new_n3458_ = new_n3457_ | new_n3456_;
  assign new_n3459_ = new_n3458_ & new_n4580_;
  assign new_n3460_ = new_n3459_ | new_n3455_;
  assign new_n3461_ = new_n4563_ & new_n2092_;
  assign new_n3462_ = new_n4573_ & new_n2200_;
  assign new_n3463_ = new_n3462_ | new_n3461_;
  assign new_n3464_ = new_n3463_ & new_n4578_;
  assign new_n3465_ = new_n4563_ & new_n2128_;
  assign new_n3466_ = new_n4575_ & new_n2164_;
  assign new_n3467_ = new_n3466_ | new_n3465_;
  assign new_n3468_ = new_n3467_ & new_n4579_;
  assign new_n3469_ = new_n3468_ | new_n3464_;
  assign new_n3470_ = new_n4401_ & new_n1907_;
  assign new_n3471_ = new_n3470_ & new_n4371_;
  assign new_n3472_ = new_n4388_ & new_n2035_;
  assign new_n3473_ = new_n3472_ | new_n3471_;
  assign new_n3474_ = new_n4389_ & new_n2042_;
  assign new_n3475_ = new_n4403_ & new_n1912_;
  assign new_n3476_ = new_n3475_ | new_n3474_;
  assign new_n3477_ = new_n3476_ & new_n4372_;
  assign new_n3478_ = new_n4374_ & new_n1954_;
  assign new_n3479_ = new_n4403_ & new_n1998_;
  assign new_n3480_ = new_n3479_ & new_n4380_;
  assign new_n3481_ = new_n3480_ | new_n3478_;
  assign new_n3482_ = new_n3481_ | new_n3477_;
  assign new_n3483_ = new_n4376_ & new_n1960_;
  assign new_n3484_ = new_n4402_ & new_n2004_;
  assign new_n3485_ = new_n3484_ & new_n4380_;
  assign new_n3486_ = new_n3485_ | new_n3483_;
  assign new_n3487_ = new_n4581_ & new_n4582_;
  assign new_n3488_ = new_n4542_ | new_n4583_;
  assign new_n3489_ = new_n4547_ | new_n4584_;
  assign new_n3490_ = new_n3489_ & new_n3488_;
  assign new_n3491_ = new_n4543_ | new_n4585_;
  assign new_n3492_ = new_n4546_ | new_n4586_;
  assign new_n3493_ = new_n3492_ & new_n3491_;
  assign new_n3494_ = new_n4550_ | new_n4552_;
  assign new_n3495_ = new_n4548_ & new_n4587_;
  assign new_n3496_ = new_n4543_ & new_n4588_;
  assign new_n3497_ = new_n3496_ | new_n4589_;
  assign new_n3498_ = new_n3497_ | new_n3495_;
  assign new_n3499_ = new_n3498_ & new_n3494_;
  assign new_n3500_ = new_n4592_ | new_n2819_;
  assign new_n3501_ = new_n4595_ | new_n2831_;
  assign new_n3502_ = new_n3501_ & new_n3500_;
  assign new_n3503_ = new_n3502_ | new_n4597_;
  assign new_n3504_ = new_n4592_ | new_n2823_;
  assign new_n3505_ = new_n4595_ | new_n2827_;
  assign new_n3506_ = new_n3505_ & new_n3504_;
  assign new_n3507_ = new_n3506_ | new_n4599_;
  assign new_n3508_ = new_n4600_ & new_n1878_;
  assign new_n3509_ = new_n4600_ & new_n1962_;
  assign new_n3510_ = new_n4602_ & new_n2006_;
  assign new_n3511_ = new_n2237_ & new_n4602_;
  assign new_n3512_ = new_n4603_ & new_n4604_;
  assign new_n3513_ = new_n4596_ & new_n2820_;
  assign new_n3514_ = new_n4591_ & new_n2832_;
  assign new_n3515_ = new_n3514_ | new_n3513_;
  assign new_n3516_ = new_n3515_ & new_n4599_;
  assign new_n3517_ = new_n4596_ & new_n2824_;
  assign new_n3518_ = new_n4593_ & new_n2828_;
  assign new_n3519_ = new_n3518_ | new_n3517_;
  assign new_n3520_ = new_n3519_ & new_n4597_;
  assign new_n3521_ = new_n3520_ | new_n3516_;
  assign G2531 = new_n4163_;
  assign G2532 = new_n4164_;
  assign G2533 = G2532;
  assign G2534 = new_n4605_;
  assign G2535 = G2534;
  assign G2536 = new_n4607_;
  assign G2537 = G2536;
  assign G2538 = new_n4606_;
  assign G2539 = new_n1887_;
  assign G2540 = new_n2177_;
  assign G2541 = new_n2015_;
  assign G2542 = new_n2069_;
  assign G2543 = new_n1971_;
  assign G2544 = new_n2141_;
  assign G2545 = new_n1929_;
  assign G2546 = new_n2105_;
  assign G2547 = new_n2836_;
  assign G2548 = new_n2838_;
  assign G2549 = new_n2208_;
  assign G2550 = new_n2839_;
  assign G2551 = new_n4165_;
  assign G2552 = new_n2841_;
  assign G2553 = new_n2842_;
  assign G2554 = new_n4608_;
  assign G2555 = G2554;
  assign G2556 = new_n4171_;
  assign G2557 = new_n2849_;
  assign G2558 = new_n2850_;
  assign G2559 = new_n2465_;
  assign G2560 = new_n2851_;
  assign G2561 = ~new_n4182_;
  assign G2562 = new_n2501_;
  assign G2563 = new_n2853_;
  assign G2564 = new_n2856_;
  assign G2565 = new_n2858_;
  assign G2566 = new_n2472_;
  assign G2567 = new_n4178_;
  assign G2568 = new_n2490_;
  assign G2569 = new_n2502_;
  assign G2570 = new_n2504_;
  assign G2571 = new_n2506_;
  assign G2572 = new_n2508_;
  assign G2573 = new_n4609_;
  assign G2574 = G2573;
  assign G2575 = ~new_n4610_;
  assign G2576 = G2575;
  assign G2577 = new_n2866_;
  assign G2578 = new_n4611_;
  assign G2579 = G2578;
  assign G2580 = new_n2873_;
  assign G2581 = ~new_n4208_;
  assign G2582 = new_n4207_;
  assign G2583 = new_n4209_;
  assign G2584 = new_n4612_;
  assign G2585 = G2584;
  assign G2586 = new_n2957_;
  assign G2587 = ~new_n4210_;
  assign G2588 = new_n4613_;
  assign G2589 = G2588;
  assign G2590 = ~new_n4211_;
  assign G2591 = new_n3007_;
  assign G2592 = new_n4615_;
  assign G2593 = new_n4614_;
  assign G2594 = G2593;
  assign n4649_li000_li000 = new_n1372_;
  assign n4652_li001_li001 = new_n1686_;
  assign n4655_li002_li002 = new_n1688_;
  assign n4658_li003_li003 = new_n1690_;
  assign n4661_li004_li004 = new_n1374_;
  assign n4664_li005_li005 = new_n1694_;
  assign n4667_li006_li006 = new_n1696_;
  assign n4670_li007_li007 = new_n1698_;
  assign n4673_li008_li008 = new_n1376_;
  assign n4676_li009_li009 = new_n1702_;
  assign n4679_li010_li010 = new_n1704_;
  assign n4682_li011_li011 = new_n1706_;
  assign n4685_li012_li012 = new_n1378_;
  assign n4688_li013_li013 = new_n1710_;
  assign n4691_li014_li014 = new_n1712_;
  assign n4697_li016_li016 = new_n1380_;
  assign n4700_li017_li017 = new_n1716_;
  assign n4703_li018_li018 = new_n1718_;
  assign n4709_li020_li020 = new_n1382_;
  assign n4712_li021_li021 = new_n1722_;
  assign n4715_li022_li022 = new_n1724_;
  assign n4721_li024_li024 = new_n1384_;
  assign n4724_li025_li025 = new_n1728_;
  assign n4727_li026_li026 = new_n1730_;
  assign n4730_li027_li027 = new_n1732_;
  assign n4733_li028_li028 = new_n1386_;
  assign n4736_li029_li029 = new_n1736_;
  assign n4745_li032_li032 = new_n1388_;
  assign n4748_li033_li033 = new_n1740_;
  assign n4751_li034_li034 = new_n1742_;
  assign n4754_li035_li035 = new_n1744_;
  assign n4757_li036_li036 = new_n1390_;
  assign n4760_li037_li037 = new_n1748_;
  assign n4763_li038_li038 = new_n1750_;
  assign n4766_li039_li039 = new_n1752_;
  assign n4769_li040_li040 = new_n1392_;
  assign n4772_li041_li041 = new_n1756_;
  assign n4775_li042_li042 = new_n1758_;
  assign n4778_li043_li043 = new_n1760_;
  assign n4781_li044_li044 = new_n1394_;
  assign n4784_li045_li045 = new_n1764_;
  assign n4787_li046_li046 = new_n1766_;
  assign n4793_li048_li048 = new_n1396_;
  assign n4796_li049_li049 = new_n1770_;
  assign n4799_li050_li050 = new_n1772_;
  assign n4805_li052_li052 = new_n1398_;
  assign n4808_li053_li053 = new_n1776_;
  assign n4811_li054_li054 = new_n1778_;
  assign n4817_li056_li056 = new_n1400_;
  assign n4820_li057_li057 = new_n1782_;
  assign n4823_li058_li058 = new_n1784_;
  assign n4829_li060_li060 = new_n1402_;
  assign n4832_li061_li061 = new_n1788_;
  assign n4835_li062_li062 = new_n1790_;
  assign n4841_li064_li064 = new_n1404_;
  assign n4844_li065_li065 = new_n1794_;
  assign n4847_li066_li066 = new_n1796_;
  assign n4853_li068_li068 = new_n1406_;
  assign n4856_li069_li069 = new_n1800_;
  assign n4859_li070_li070 = new_n1802_;
  assign n4865_li072_li072 = new_n1408_;
  assign n4868_li073_li073 = new_n1806_;
  assign n4871_li074_li074 = new_n1808_;
  assign n4877_li076_li076 = new_n1410_;
  assign n4880_li077_li077 = new_n1812_;
  assign n4883_li078_li078 = new_n1814_;
  assign n4889_li080_li080 = new_n1412_;
  assign n4892_li081_li081 = new_n1818_;
  assign n4895_li082_li082 = new_n1820_;
  assign n4901_li084_li084 = new_n1414_;
  assign n4904_li085_li085 = new_n1824_;
  assign n4907_li086_li086 = new_n1826_;
  assign n4913_li088_li088 = new_n1416_;
  assign n4916_li089_li089 = new_n1830_;
  assign n4919_li090_li090 = new_n1832_;
  assign n4925_li092_li092 = new_n1418_;
  assign n4928_li093_li093 = new_n1836_;
  assign n4931_li094_li094 = new_n1838_;
  assign n4937_li096_li096 = new_n1420_;
  assign n4940_li097_li097 = new_n1842_;
  assign n4943_li098_li098 = new_n1844_;
  assign n4949_li100_li100 = new_n1422_;
  assign n4952_li101_li101 = new_n1848_;
  assign n4955_li102_li102 = new_n1850_;
  assign n4961_li104_li104 = new_n1424_;
  assign n4964_li105_li105 = new_n1854_;
  assign n4967_li106_li106 = new_n1856_;
  assign n4973_li108_li108 = new_n1426_;
  assign n4976_li109_li109 = new_n1860_;
  assign n4979_li110_li110 = new_n1862_;
  assign n4982_li111_li111 = new_n1864_;
  assign n4985_li112_li112 = new_n1428_;
  assign n4988_li113_li113 = new_n1868_;
  assign n4991_li114_li114 = new_n1870_;
  assign n4994_li115_li115 = new_n1872_;
  assign n4997_li116_li116 = new_n1430_;
  assign n5009_li120_li120 = new_n1432_;
  assign n5021_li124_li124 = new_n1434_;
  assign n5024_li125_li125 = new_n1880_;
  assign n5027_li126_li126 = new_n1882_;
  assign n5030_li127_li127 = new_n4407_;
  assign n5033_li128_li128 = new_n1436_;
  assign n5036_li129_li129 = new_n1888_;
  assign n5045_li132_li132 = new_n1438_;
  assign n5048_li133_li133 = new_n1892_;
  assign n5057_li136_li136 = new_n1440_;
  assign n5060_li137_li137 = new_n1896_;
  assign n5069_li140_li140 = new_n1442_;
  assign n5072_li141_li141 = new_n1900_;
  assign n5081_li144_li144 = new_n1444_;
  assign n5084_li145_li145 = new_n1904_;
  assign n5093_li148_li148 = new_n1446_;
  assign n5105_li152_li152 = new_n1448_;
  assign n5108_li153_li153 = new_n1910_;
  assign n5117_li156_li156 = new_n1450_;
  assign n5129_li160_li160 = new_n1452_;
  assign n5132_li161_li161 = new_n1916_;
  assign n5141_li164_li164 = new_n1454_;
  assign n5153_li168_li168 = new_n1456_;
  assign n5156_li169_li169 = new_n1922_;
  assign n5159_li170_li170 = new_n1924_;
  assign n5162_li171_li171 = new_n4409_;
  assign n5165_li172_li172 = new_n1458_;
  assign n5168_li173_li173 = new_n1930_;
  assign n5177_li176_li176 = new_n1460_;
  assign n5180_li177_li177 = new_n1934_;
  assign n5189_li180_li180 = new_n1462_;
  assign n5192_li181_li181 = new_n1938_;
  assign n5195_li182_li182 = new_n1940_;
  assign n5201_li184_li184 = new_n1464_;
  assign n5204_li185_li185 = new_n1944_;
  assign n5213_li188_li188 = new_n1466_;
  assign n5216_li189_li189 = new_n1948_;
  assign n5225_li192_li192 = new_n1468_;
  assign n5228_li193_li193 = new_n1952_;
  assign n5237_li196_li196 = new_n1470_;
  assign n5249_li200_li200 = new_n1472_;
  assign n5252_li201_li201 = new_n1958_;
  assign n5261_li204_li204 = new_n1474_;
  assign n5273_li208_li208 = new_n1476_;
  assign n5276_li209_li209 = new_n1964_;
  assign n5279_li210_li210 = new_n1966_;
  assign n5282_li211_li211 = new_n4408_;
  assign n5285_li212_li212 = new_n1478_;
  assign n5288_li213_li213 = new_n1972_;
  assign n5297_li216_li216 = new_n1480_;
  assign n5300_li217_li217 = new_n1976_;
  assign n5309_li220_li220 = new_n1482_;
  assign n5312_li221_li221 = new_n1980_;
  assign n5321_li224_li224 = new_n1484_;
  assign n5324_li225_li225 = new_n1984_;
  assign n5333_li228_li228 = new_n1486_;
  assign n5336_li229_li229 = new_n1988_;
  assign n5345_li232_li232 = new_n1488_;
  assign n5348_li233_li233 = new_n1992_;
  assign n5357_li236_li236 = new_n1490_;
  assign n5360_li237_li237 = new_n1996_;
  assign n5369_li240_li240 = new_n1492_;
  assign n5381_li244_li244 = new_n1494_;
  assign n5384_li245_li245 = new_n2002_;
  assign n5393_li248_li248 = new_n1496_;
  assign n5405_li252_li252 = new_n1498_;
  assign n5408_li253_li253 = new_n2008_;
  assign n5411_li254_li254 = new_n2010_;
  assign n5414_li255_li255 = new_n4406_;
  assign n5417_li256_li256 = new_n1500_;
  assign n5420_li257_li257 = new_n2016_;
  assign n5429_li260_li260 = new_n1502_;
  assign n5432_li261_li261 = new_n2020_;
  assign n5441_li264_li264 = new_n1504_;
  assign n5444_li265_li265 = new_n2024_;
  assign n5453_li268_li268 = new_n1506_;
  assign n5456_li269_li269 = new_n2028_;
  assign n5465_li272_li272 = new_n1508_;
  assign n5468_li273_li273 = new_n2032_;
  assign n5477_li276_li276 = new_n1510_;
  assign n5480_li277_li277 = new_n2036_;
  assign n5489_li280_li280 = new_n1512_;
  assign n5492_li281_li281 = new_n2040_;
  assign n5501_li284_li284 = new_n1514_;
  assign n5513_li288_li288 = new_n1516_;
  assign n5516_li289_li289 = new_n2046_;
  assign n5525_li292_li292 = new_n1518_;
  assign n5528_li293_li293 = new_n2050_;
  assign n5531_li294_li294 = new_n2052_;
  assign n5534_li295_li295 = new_n2054_;
  assign n5537_li296_li296 = new_n1520_;
  assign n5540_li297_li297 = new_n2058_;
  assign n5549_li300_li300 = new_n1522_;
  assign n5552_li301_li301 = new_n2062_;
  assign n5555_li302_li302 = new_n2064_;
  assign n5558_li303_li303 = new_n4411_;
  assign n5561_li304_li304 = new_n1524_;
  assign n5564_li305_li305 = new_n2070_;
  assign n5573_li308_li308 = new_n1526_;
  assign n5576_li309_li309 = new_n2074_;
  assign n5609_li320_li320 = new_n1532_;
  assign n5612_li321_li321 = new_n2078_;
  assign n5621_li324_li324 = new_n1534_;
  assign n5624_li325_li325 = new_n2082_;
  assign n5633_li328_li328 = new_n1536_;
  assign n5636_li329_li329 = new_n2086_;
  assign n5645_li332_li332 = new_n1538_;
  assign n5648_li333_li333 = new_n2090_;
  assign n5657_li336_li336 = new_n1540_;
  assign n5660_li337_li337 = new_n2094_;
  assign n5669_li340_li340 = new_n1542_;
  assign n5672_li341_li341 = new_n2098_;
  assign n5675_li342_li342 = new_n2100_;
  assign n5678_li343_li343 = new_n4413_;
  assign n5681_li344_li344 = new_n1544_;
  assign n5684_li345_li345 = new_n2106_;
  assign n5693_li348_li348 = new_n1546_;
  assign n5696_li349_li349 = new_n2110_;
  assign n5729_li360_li360 = new_n1552_;
  assign n5732_li361_li361 = new_n2114_;
  assign n5741_li364_li364 = new_n1554_;
  assign n5744_li365_li365 = new_n2118_;
  assign n5753_li368_li368 = new_n1556_;
  assign n5756_li369_li369 = new_n2122_;
  assign n5765_li372_li372 = new_n1558_;
  assign n5768_li373_li373 = new_n2126_;
  assign n5777_li376_li376 = new_n1560_;
  assign n5780_li377_li377 = new_n2130_;
  assign n5789_li380_li380 = new_n1562_;
  assign n5792_li381_li381 = new_n2134_;
  assign n5795_li382_li382 = new_n2136_;
  assign n5798_li383_li383 = new_n4412_;
  assign n5801_li384_li384 = new_n1564_;
  assign n5804_li385_li385 = new_n2142_;
  assign n5813_li388_li388 = new_n1566_;
  assign n5816_li389_li389 = new_n2146_;
  assign n5849_li400_li400 = new_n1572_;
  assign n5852_li401_li401 = new_n2150_;
  assign n5861_li404_li404 = new_n1574_;
  assign n5864_li405_li405 = new_n2154_;
  assign n5873_li408_li408 = new_n1576_;
  assign n5876_li409_li409 = new_n2158_;
  assign n5885_li412_li412 = new_n1578_;
  assign n5888_li413_li413 = new_n2162_;
  assign n5897_li416_li416 = new_n1580_;
  assign n5900_li417_li417 = new_n2166_;
  assign n5909_li420_li420 = new_n1582_;
  assign n5912_li421_li421 = new_n2170_;
  assign n5915_li422_li422 = new_n2172_;
  assign n5918_li423_li423 = new_n4410_;
  assign n5921_li424_li424 = new_n1584_;
  assign n5924_li425_li425 = new_n2178_;
  assign n5933_li428_li428 = new_n1586_;
  assign n5936_li429_li429 = new_n2182_;
  assign n5969_li440_li440 = new_n1592_;
  assign n5972_li441_li441 = new_n2186_;
  assign n5981_li444_li444 = new_n1594_;
  assign n5984_li445_li445 = new_n2190_;
  assign n5993_li448_li448 = new_n1596_;
  assign n5996_li449_li449 = new_n2194_;
  assign n6005_li452_li452 = new_n1598_;
  assign n6008_li453_li453 = new_n2198_;
  assign n6017_li456_li456 = new_n1600_;
  assign n6020_li457_li457 = new_n2202_;
  assign n6023_li458_li458 = new_n2204_;
  assign n6026_li459_li459 = new_n2206_;
  assign n6029_li460_li460 = new_n1602_;
  assign n6032_li461_li461 = new_n2210_;
  assign n6035_li462_li462 = new_n2212_;
  assign n6038_li463_li463 = new_n2214_;
  assign n6041_li464_li464 = new_n1604_;
  assign n6053_li468_li468 = new_n1606_;
  assign n6056_li469_li469 = new_n2220_;
  assign n6059_li470_li470 = new_n2222_;
  assign n6062_li471_li471 = new_n4414_;
  assign n6065_li472_li472 = new_n1608_;
  assign n6068_li473_li473 = new_n2228_;
  assign n6071_li474_li474 = new_n2230_;
  assign n6074_li475_li475 = new_n2232_;
  assign n6077_li476_li476 = new_n1610_;
  assign n6089_li480_li480 = new_n1612_;
  assign n6092_li481_li481 = new_n2238_;
  assign n6095_li482_li482 = new_n2240_;
  assign n6098_li483_li483 = new_n2242_;
  assign n6101_li484_li484 = new_n1614_;
  assign n6104_li485_li485 = new_n2246_;
  assign n6107_li486_li486 = new_n2248_;
  assign n6110_li487_li487 = new_n2250_;
  assign n6113_li488_li488 = new_n1616_;
  assign n6116_li489_li489 = new_n2254_;
  assign n6119_li490_li490 = new_n2256_;
  assign n6122_li491_li491 = new_n2258_;
  assign n6125_li492_li492 = new_n1618_;
  assign n6128_li493_li493 = new_n2262_;
  assign n6131_li494_li494 = new_n2264_;
  assign n6134_li495_li495 = new_n2266_;
  assign n6137_li496_li496 = new_n1620_;
  assign n6140_li497_li497 = new_n2270_;
  assign n6149_li500_li500 = new_n1622_;
  assign n6152_li501_li501 = new_n2274_;
  assign n6158_li503_li503 = new_n4504_;
  assign n6161_li504_li504 = new_n1624_;
  assign n6173_li508_li508 = new_n1626_;
  assign n6176_li509_li509 = new_n2282_;
  assign n6185_li512_li512 = new_n1628_;
  assign n6188_li513_li513 = new_n2286_;
  assign n6194_li515_li515 = new_n4467_;
  assign n6197_li516_li516 = new_n1630_;
  assign n6200_li517_li517 = new_n2292_;
  assign n6203_li518_li518 = new_n2294_;
  assign n6209_li520_li520 = new_n1632_;
  assign n6212_li521_li521 = new_n2298_;
  assign n6215_li522_li522 = new_n2300_;
  assign n6221_li524_li524 = new_n1634_;
  assign n6224_li525_li525 = new_n2304_;
  assign n6227_li526_li526 = new_n2306_;
  assign n6230_li527_li527 = new_n4507_;
  assign n6233_li528_li528 = new_n1636_;
  assign n6236_li529_li529 = new_n2312_;
  assign n6239_li530_li530 = new_n2314_;
  assign n6245_li532_li532 = new_n1638_;
  assign n6248_li533_li533 = new_n2318_;
  assign n6251_li534_li534 = new_n2320_;
  assign n6254_li535_li535 = new_n4284_;
  assign n6257_li536_li536 = new_n1640_;
  assign n6260_li537_li537 = new_n2326_;
  assign n6263_li538_li538 = new_n2328_;
  assign n6266_li539_li539 = new_n4470_;
  assign n6269_li540_li540 = new_n1642_;
  assign n6272_li541_li541 = new_n2334_;
  assign n6278_li543_li543 = new_n4353_;
  assign n6281_li544_li544 = new_n1644_;
  assign n6284_li545_li545 = new_n2340_;
  assign n6287_li546_li546 = new_n2342_;
  assign n6290_li547_li547 = new_n2344_;
  assign n6293_li548_li548 = new_n1646_;
  assign n6296_li549_li549 = new_n2348_;
  assign n6302_li551_li551 = new_n4490_;
  assign n6305_li552_li552 = new_n1648_;
  assign n6308_li553_li553 = new_n2354_;
  assign n6314_li555_li555 = new_n4234_;
  assign n6317_li556_li556 = new_n1650_;
  assign n6320_li557_li557 = new_n2360_;
  assign n6326_li559_li559 = new_n4232_;
  assign n6329_li560_li560 = new_n1652_;
  assign n6332_li561_li561 = new_n2366_;
  assign n6335_li562_li562 = new_n2368_;
  assign n6338_li563_li563 = new_n4486_;
  assign n6341_li564_li564 = new_n1654_;
  assign n6344_li565_li565 = new_n2374_;
  assign n6347_li566_li566 = new_n2376_;
  assign n6350_li567_li567 = new_n4485_;
  assign n6353_li568_li568 = new_n1656_;
  assign n6356_li569_li569 = new_n2382_;
  assign n6359_li570_li570 = new_n2384_;
  assign n6362_li571_li571 = new_n4449_;
  assign n6365_li572_li572 = new_n1658_;
  assign n6368_li573_li573 = new_n2390_;
  assign n6371_li574_li574 = new_n2392_;
  assign n6374_li575_li575 = new_n4450_;
  assign n6389_li580_li580 = new_n1662_;
  assign n6401_li584_li584 = new_n1664_;
  assign n6404_li585_li585 = new_n2400_;
  assign n6407_li586_li586 = new_n2402_;
  assign n6410_li587_li587 = new_n2404_;
  assign n6413_li588_li588 = new_n1666_;
  assign n6416_li589_li589 = new_n2408_;
  assign n6425_li592_li592 = new_n1668_;
  assign n6428_li593_li593 = new_n2412_;
  assign n6437_li596_li596 = new_n1670_;
  assign n6440_li597_li597 = new_n2416_;
  assign n6443_li598_li598 = new_n2418_;
  assign n6449_li600_li600 = new_n1672_;
  assign n6452_li601_li601 = new_n2422_;
  assign n6455_li602_li602 = new_n2424_;
  assign n6461_li604_li604 = new_n1674_;
  assign n6464_li605_li605 = new_n2428_;
  assign n6473_li608_li608 = new_n1676_;
  assign n6476_li609_li609 = new_n2432_;
  assign n6485_li612_li612 = new_n1678_;
  assign n6488_li613_li613 = new_n2436_;
  assign n6491_li614_li614 = new_n2438_;
  assign n6497_li616_li616 = new_n1680_;
  assign n6500_li617_li617 = new_n2442_;
  assign n6503_li618_li618 = new_n2444_;
  assign n6509_li620_li620 = new_n1682_;
  assign n6512_li621_li621 = new_n2448_;
  assign n6515_li622_li622 = new_n2450_;
  assign n6521_li624_li624 = new_n1684_;
  assign n6524_li625_li625 = new_n2454_;
  assign n6527_li626_li626 = new_n2456_;
  assign n3603_i2 = new_n2512_;
  assign n3604_i2 = new_n2514_;
  assign n3618_i2 = new_n4324_;
  assign n3798_i2 = new_n4262_;
  assign n3846_i2 = new_n4302_;
  assign n4019_i2 = new_n4455_;
  assign n4017_i2 = new_n4359_;
  assign n2177_i2 = new_n4241_;
  assign n2150_i2 = new_n4464_;
  assign n2154_i2 = new_n4463_;
  assign n2184_i2 = new_n4240_;
  assign n2515_i2 = new_n4256_;
  assign n3837_i2 = new_n4575_;
  assign n2167_i2 = new_n4253_;
  assign n2118_i2 = new_n4488_;
  assign n2186_i2 = new_n4428_;
  assign n2174_i2 = new_n4252_;
  assign n3964_i2 = new_n4578_;
  assign n4005_i2 = new_n4389_;
  assign n4006_i2 = new_n4372_;
  assign n2195_i2 = new_n4495_;
  assign n2176_i2 = new_n4278_;
  assign n2227_i2 = new_n4313_;
  assign n2236_i2 = new_n4438_;
  assign n2245_i2 = new_n4311_;
  assign n2518_i2 = new_n4362_;
  assign n4023_i2 = new_n2786_;
  assign n4024_i2 = new_n2788_;
  assign n4038_i2 = new_n4376_;
  assign n4039_i2 = new_n4272_;
  assign n4040_i2 = new_n4273_;
  assign n2119_i2 = ~new_n4487_;
  assign n2275_i2 = new_n4404_;
  assign n2595_i2 = new_n4275_;
  assign n2594_i2 = new_n4274_;
  assign lo498_buf_i2 = new_n4588_;
  assign lo502_buf_i2 = new_n4549_;
  assign lo550_buf_i2 = new_n4544_;
  assign n2596_i2 = new_n4548_;
  assign n2593_i2 = ~new_n4457_;
  assign n2668_i2 = ~new_n4469_;
  assign lo542_buf_i2 = new_n4587_;
  assign n2667_i2 = new_n4468_;
  assign n2404_i2 = new_n4419_;
  assign n2410_i2 = new_n4444_;
  assign n2419_i2 = new_n4434_;
  assign n2392_i2 = new_n4447_;
  assign n2369_i2 = new_n4446_;
  assign n2397_i2 = new_n4448_;
  assign n2601_i2 = new_n4456_;
  assign n2658_i2 = ~new_n4484_;
  assign n2574_i2 = ~new_n4497_;
  assign n2205_i2 = new_n4589_;
  assign lo510_buf_i2 = new_n4584_;
  assign lo514_buf_i2 = new_n4586_;
  assign lo554_buf_i2 = new_n4583_;
  assign lo558_buf_i2 = new_n4585_;
  assign lo578_buf_i2 = new_n4593_;
  assign n2254_i2 = new_n4551_;
  assign n2421_i2 = new_n3167_;
  assign n2422_i2 = new_n3168_;
  assign n2130_i2 = new_n3169_;
  assign n2127_i2 = new_n3170_;
  assign n2131_i2 = new_n3171_;
  assign n2128_i2 = new_n3172_;
  assign n2264_i2 = new_n3173_;
  assign n2467_i2 = ~new_n3177_;
  assign n2471_i2 = new_n3178_;
  assign n2488_i2 = ~new_n3179_;
  assign n2478_i2 = ~new_n3183_;
  assign n2486_i2 = new_n3184_;
  assign n2485_i2 = new_n3188_;
  assign n2498_i2 = ~new_n3189_;
  assign n2495_i2 = new_n3193_;
  assign n2496_i2 = ~new_n3194_;
  assign n2458_i2 = new_n3195_;
  assign n2643_i2 = new_n3196_;
  assign n2462_i2 = new_n3200_;
  assign n2468_i2 = ~new_n3201_;
  assign n2639_i2 = new_n3202_;
  assign n2499_i2 = ~new_n3203_;
  assign n2472_i2 = new_n3204_;
  assign n2474_i2 = ~new_n3205_;
  assign n2489_i2 = new_n3206_;
  assign n2321_i2 = new_n3207_;
  assign n2322_i2 = new_n3208_;
  assign n2640_i2 = new_n3209_;
  assign n2642_i2 = new_n3210_;
  assign n2187_i2 = ~new_n4582_;
  assign n2373_i2 = new_n3214_;
  assign n2603_i2 = ~new_n3215_;
  assign n2388_i2 = new_n3218_;
  assign n2437_i2 = new_n3227_;
  assign n2356_i2 = new_n3232_;
  assign n2452_i2 = new_n3235_;
  assign n2347_i2 = new_n3238_;
  assign n2329_i2 = new_n3241_;
  assign n2669_i2 = ~new_n3242_;
  assign n2332_i2 = new_n3245_;
  assign n2664_i2 = new_n3248_;
  assign n2665_i2 = ~new_n3249_;
  assign n2653_i2 = new_n3252_;
  assign n2654_i2 = ~new_n3253_;
  assign n2636_i2 = ~new_n3270_;
  assign n2660_i2 = ~new_n3272_;
  assign n2318_i2 = ~new_n3288_;
  assign n2319_i2 = new_n3289_;
  assign n2586_i2 = ~new_n3293_;
  assign n2587_i2 = ~new_n3294_;
  assign n2288_i2 = new_n3309_;
  assign n2344_i2 = new_n3324_;
  assign n2530_i2 = new_n3333_;
  assign n2303_i2 = new_n3360_;
  assign n2566_i2 = new_n3367_;
  assign n2567_i2 = ~new_n3368_;
  assign n2554_i2 = new_n3395_;
  assign n2194_i2 = ~new_n4581_;
  assign lo582_buf_i2 = new_n4598_;
  assign lo030_buf_i2 = new_n1738_;
  assign lo174_buf_i2 = new_n1932_;
  assign lo178_buf_i2 = new_n1936_;
  assign lo186_buf_i2 = new_n1946_;
  assign lo266_buf_i2 = new_n2026_;
  assign lo306_buf_i2 = new_n2072_;
  assign lo346_buf_i2 = new_n2108_;
  assign lo386_buf_i2 = new_n2144_;
  assign lo426_buf_i2 = new_n2180_;
  assign lo590_buf_i2 = new_n2410_;
  assign lo594_buf_i2 = new_n2414_;
  assign lo606_buf_i2 = new_n2430_;
  assign lo610_buf_i2 = new_n2434_;
  assign n2238_i2 = new_n3403_;
  assign n2229_i2 = new_n3404_;
  assign n2242_i2 = new_n3405_;
  assign n2233_i2 = new_n3406_;
  assign n2168_i2 = new_n3407_;
  assign n2237_i2 = new_n3408_;
  assign n2228_i2 = new_n3409_;
  assign n2172_i2 = new_n3410_;
  assign n2223_i2 = new_n3411_;
  assign n2222_i2 = new_n3412_;
  assign n2170_i2 = new_n3414_;
  assign n2181_i2 = new_n3416_;
  assign n2510_i2 = new_n3420_;
  assign n2621_i2 = new_n3424_;
  assign lo466_buf_i2 = new_n4601_;
  assign lo478_buf_i2 = new_n2236_;
  assign n2149_i2 = new_n3427_;
  assign n2429_i2 = new_n3430_;
  assign n2444_i2 = new_n3433_;
  assign n2153_i2 = new_n3436_;
  assign n2433_i2 = new_n3439_;
  assign n2448_i2 = new_n3442_;
  assign n2367_i2 = new_n3451_;
  assign n2386_i2 = new_n3460_;
  assign n2539_i2 = new_n3469_;
  assign n2183_i2 = new_n3473_;
  assign n2220_i2 = new_n3482_;
  assign n2514_i2 = new_n3486_;
  assign n2196_i2 = ~new_n3487_;
  assign n2616_i2 = new_n3490_;
  assign n2612_i2 = new_n3493_;
  assign n2627_i2 = new_n3499_;
  assign n2140_i2 = ~new_n4604_;
  assign n2144_i2 = ~new_n4603_;
  assign lo149_buf_i2 = new_n1908_;
  assign lo197_buf_i2 = new_n1956_;
  assign lo118_buf_i2 = new_n1876_;
  assign lo158_buf_i2 = new_n1914_;
  assign lo166_buf_i2 = new_n1920_;
  assign lo242_buf_i2 = new_n2000_;
  assign lo286_buf_i2 = new_n2044_;
  assign lo506_buf_i2 = new_n2280_;
  assign n2198_i2 = new_n3508_;
  assign n2202_i2 = new_n3509_;
  assign n2197_i2 = new_n3510_;
  assign n2166_i2 = new_n3511_;
  assign n2146_i2 = ~new_n3512_;
  assign n2165_i2 = new_n3521_;
  assign lo312_buf_i2 = new_n1528_;
  assign lo316_buf_i2 = new_n1530_;
  assign lo352_buf_i2 = new_n1548_;
  assign lo356_buf_i2 = new_n1550_;
  assign lo392_buf_i2 = new_n1568_;
  assign lo396_buf_i2 = new_n1570_;
  assign lo432_buf_i2 = new_n1588_;
  assign lo436_buf_i2 = new_n1590_;
  assign lo576_buf_i2 = new_n1660_;
  assign new_n4161_ = new_n2245_;
  assign new_n4162_ = new_n2209_;
  assign new_n4163_ = new_n4162_;
  assign new_n4164_ = new_n4162_;
  assign new_n4165_ = new_n2840_;
  assign new_n4166_ = new_n4165_;
  assign new_n4167_ = new_n2844_;
  assign new_n4168_ = new_n2843_;
  assign new_n4169_ = new_n2253_;
  assign new_n4170_ = new_n4169_;
  assign new_n4171_ = new_n2848_;
  assign new_n4172_ = new_n4171_;
  assign new_n4173_ = new_n2855_;
  assign new_n4174_ = new_n2469_;
  assign new_n4175_ = new_n2260_;
  assign new_n4176_ = new_n4175_;
  assign new_n4177_ = new_n4175_;
  assign new_n4178_ = new_n2470_;
  assign new_n4179_ = new_n2261_;
  assign new_n4180_ = new_n4179_;
  assign new_n4181_ = new_n4179_;
  assign new_n4182_ = new_n2852_;
  assign new_n4183_ = new_n2226_;
  assign new_n4184_ = new_n2468_;
  assign new_n4185_ = new_n2591_;
  assign new_n4186_ = new_n4185_;
  assign new_n4187_ = new_n2657_;
  assign new_n4188_ = new_n2652_;
  assign new_n4189_ = new_n2656_;
  assign new_n4190_ = new_n2653_;
  assign new_n4191_ = new_n2680_;
  assign new_n4192_ = new_n2651_;
  assign new_n4193_ = new_n2681_;
  assign new_n4194_ = new_n2650_;
  assign new_n4195_ = new_n2482_;
  assign new_n4196_ = new_n1875_;
  assign new_n4197_ = new_n2590_;
  assign new_n4198_ = new_n2563_;
  assign new_n4199_ = new_n2562_;
  assign new_n4200_ = new_n2963_;
  assign new_n4201_ = new_n2964_;
  assign new_n4202_ = new_n2985_;
  assign new_n4203_ = new_n2992_;
  assign new_n4204_ = new_n2668_;
  assign new_n4205_ = new_n2994_;
  assign new_n4206_ = new_n2993_;
  assign new_n4207_ = new_n2884_;
  assign new_n4208_ = new_n2877_;
  assign new_n4209_ = new_n2899_;
  assign new_n4210_ = new_n2961_;
  assign new_n4211_ = new_n2981_;
  assign new_n4212_ = new_n2516_;
  assign new_n4213_ = new_n4212_;
  assign new_n4214_ = new_n4212_;
  assign new_n4215_ = new_n2517_;
  assign new_n4216_ = new_n4215_;
  assign new_n4217_ = new_n4215_;
  assign new_n4218_ = new_n2494_;
  assign new_n4219_ = new_n4218_;
  assign new_n4220_ = new_n4219_;
  assign new_n4221_ = new_n4219_;
  assign new_n4222_ = new_n4218_;
  assign new_n4223_ = new_n4222_;
  assign new_n4224_ = new_n4222_;
  assign new_n4225_ = new_n2495_;
  assign new_n4226_ = new_n4225_;
  assign new_n4227_ = new_n4226_;
  assign new_n4228_ = new_n4226_;
  assign new_n4229_ = new_n4225_;
  assign new_n4230_ = new_n4229_;
  assign new_n4231_ = new_n4229_;
  assign new_n4232_ = new_n2572_;
  assign new_n4233_ = new_n4232_;
  assign new_n4234_ = new_n2570_;
  assign new_n4235_ = new_n4234_;
  assign new_n4236_ = new_n2573_;
  assign new_n4237_ = new_n4236_;
  assign new_n4238_ = new_n2571_;
  assign new_n4239_ = new_n4238_;
  assign new_n4240_ = new_n3019_;
  assign new_n4241_ = new_n3013_;
  assign new_n4242_ = new_n2499_;
  assign new_n4243_ = new_n4242_;
  assign new_n4244_ = new_n4243_;
  assign new_n4245_ = new_n4243_;
  assign new_n4246_ = new_n4242_;
  assign new_n4247_ = new_n2498_;
  assign new_n4248_ = new_n4247_;
  assign new_n4249_ = new_n4248_;
  assign new_n4250_ = new_n4248_;
  assign new_n4251_ = new_n4247_;
  assign new_n4252_ = new_n3033_;
  assign new_n4253_ = new_n3023_;
  assign new_n4254_ = new_n2497_;
  assign new_n4255_ = new_n2496_;
  assign new_n4256_ = new_n3022_;
  assign new_n4257_ = new_n4256_;
  assign new_n4258_ = new_n2565_;
  assign new_n4259_ = new_n3021_;
  assign new_n4260_ = new_n2564_;
  assign new_n4261_ = new_n4260_;
  assign new_n4262_ = new_n4260_;
  assign new_n4263_ = new_n2379_;
  assign new_n4264_ = new_n2371_;
  assign new_n4265_ = new_n4264_;
  assign new_n4266_ = new_n2485_;
  assign new_n4267_ = new_n4266_;
  assign new_n4268_ = new_n4266_;
  assign new_n4269_ = new_n2484_;
  assign new_n4270_ = new_n4269_;
  assign new_n4271_ = new_n4269_;
  assign new_n4272_ = new_n2814_;
  assign new_n4273_ = new_n2816_;
  assign new_n4274_ = new_n3100_;
  assign new_n4275_ = new_n3098_;
  assign new_n4276_ = new_n3038_;
  assign new_n4277_ = new_n4276_;
  assign new_n4278_ = new_n4276_;
  assign new_n4279_ = new_n2697_;
  assign new_n4280_ = new_n3106_;
  assign new_n4281_ = new_n4280_;
  assign new_n4282_ = new_n4281_;
  assign new_n4283_ = new_n4280_;
  assign new_n4284_ = new_n2322_;
  assign new_n4285_ = new_n4284_;
  assign new_n4286_ = new_n3105_;
  assign new_n4287_ = new_n4286_;
  assign new_n4288_ = new_n4287_;
  assign new_n4289_ = new_n4286_;
  assign new_n4290_ = new_n3071_;
  assign new_n4291_ = new_n1768_;
  assign new_n4292_ = new_n4291_;
  assign new_n4293_ = new_n4292_;
  assign new_n4294_ = new_n4293_;
  assign new_n4295_ = new_n4292_;
  assign new_n4296_ = new_n4291_;
  assign new_n4297_ = new_n4296_;
  assign new_n4298_ = new_n4296_;
  assign new_n4299_ = new_n2576_;
  assign new_n4300_ = new_n4299_;
  assign new_n4301_ = new_n4300_;
  assign new_n4302_ = new_n4299_;
  assign new_n4303_ = new_n1769_;
  assign new_n4304_ = new_n4303_;
  assign new_n4305_ = new_n4304_;
  assign new_n4306_ = new_n4305_;
  assign new_n4307_ = new_n4304_;
  assign new_n4308_ = new_n4303_;
  assign new_n4309_ = new_n4308_;
  assign new_n4310_ = new_n4308_;
  assign new_n4311_ = new_n3072_;
  assign new_n4312_ = new_n4311_;
  assign new_n4313_ = new_n3047_;
  assign new_n4314_ = new_n4313_;
  assign new_n4315_ = new_n1834_;
  assign new_n4316_ = new_n4315_;
  assign new_n4317_ = new_n4316_;
  assign new_n4318_ = new_n4316_;
  assign new_n4319_ = new_n4315_;
  assign new_n4320_ = new_n4319_;
  assign new_n4321_ = new_n4319_;
  assign new_n4322_ = new_n2520_;
  assign new_n4323_ = new_n4322_;
  assign new_n4324_ = new_n4322_;
  assign new_n4325_ = new_n1835_;
  assign new_n4326_ = new_n4325_;
  assign new_n4327_ = new_n4326_;
  assign new_n4328_ = new_n4326_;
  assign new_n4329_ = new_n4325_;
  assign new_n4330_ = new_n4329_;
  assign new_n4331_ = new_n4329_;
  assign new_n4332_ = new_n2766_;
  assign new_n4333_ = new_n4332_;
  assign new_n4334_ = new_n2518_;
  assign new_n4335_ = new_n4334_;
  assign new_n4336_ = new_n2696_;
  assign new_n4337_ = new_n3127_;
  assign new_n4338_ = new_n4337_;
  assign new_n4339_ = new_n4337_;
  assign new_n4340_ = new_n2303_;
  assign new_n4341_ = new_n4340_;
  assign new_n4342_ = new_n4341_;
  assign new_n4343_ = new_n4340_;
  assign new_n4344_ = new_n3129_;
  assign new_n4345_ = new_n4344_;
  assign new_n4346_ = new_n4344_;
  assign new_n4347_ = new_n3137_;
  assign new_n4348_ = new_n4347_;
  assign new_n4349_ = new_n4347_;
  assign new_n4350_ = new_n3136_;
  assign new_n4351_ = new_n4350_;
  assign new_n4352_ = new_n2543_;
  assign new_n4353_ = new_n2542_;
  assign new_n4354_ = new_n4353_;
  assign new_n4355_ = new_n2774_;
  assign new_n4356_ = new_n4355_;
  assign new_n4357_ = new_n4356_;
  assign new_n4358_ = new_n4356_;
  assign new_n4359_ = new_n4355_;
  assign new_n4360_ = new_n2775_;
  assign new_n4361_ = new_n2577_;
  assign new_n4362_ = new_n3078_;
  assign new_n4363_ = new_n2752_;
  assign new_n4364_ = new_n4363_;
  assign new_n4365_ = new_n4364_;
  assign new_n4366_ = new_n4365_;
  assign new_n4367_ = new_n4365_;
  assign new_n4368_ = new_n4364_;
  assign new_n4369_ = new_n4368_;
  assign new_n4370_ = new_n4363_;
  assign new_n4371_ = new_n4370_;
  assign new_n4372_ = new_n4370_;
  assign new_n4373_ = new_n2812_;
  assign new_n4374_ = new_n4373_;
  assign new_n4375_ = new_n4374_;
  assign new_n4376_ = new_n4373_;
  assign new_n4377_ = new_n2753_;
  assign new_n4378_ = new_n4377_;
  assign new_n4379_ = new_n4378_;
  assign new_n4380_ = new_n4377_;
  assign new_n4381_ = new_n2750_;
  assign new_n4382_ = new_n4381_;
  assign new_n4383_ = new_n4382_;
  assign new_n4384_ = new_n4383_;
  assign new_n4385_ = new_n4383_;
  assign new_n4386_ = new_n4382_;
  assign new_n4387_ = new_n4381_;
  assign new_n4388_ = new_n4387_;
  assign new_n4389_ = new_n4387_;
  assign new_n4390_ = new_n2751_;
  assign new_n4391_ = new_n4390_;
  assign new_n4392_ = new_n4391_;
  assign new_n4393_ = new_n4392_;
  assign new_n4394_ = new_n4392_;
  assign new_n4395_ = new_n4391_;
  assign new_n4396_ = new_n4395_;
  assign new_n4397_ = new_n4395_;
  assign new_n4398_ = new_n4390_;
  assign new_n4399_ = new_n4398_;
  assign new_n4400_ = new_n4399_;
  assign new_n4401_ = new_n4399_;
  assign new_n4402_ = new_n4398_;
  assign new_n4403_ = new_n4402_;
  assign new_n4404_ = new_n3097_;
  assign new_n4405_ = new_n4404_;
  assign new_n4406_ = new_n2012_;
  assign new_n4407_ = new_n1884_;
  assign new_n4408_ = new_n1968_;
  assign new_n4409_ = new_n1926_;
  assign new_n4410_ = new_n2174_;
  assign new_n4411_ = new_n2066_;
  assign new_n4412_ = new_n2138_;
  assign new_n4413_ = new_n2102_;
  assign new_n4414_ = new_n2224_;
  assign new_n4415_ = new_n3176_;
  assign new_n4416_ = new_n2531_;
  assign new_n4417_ = new_n4416_;
  assign new_n4418_ = new_n4416_;
  assign new_n4419_ = new_n3111_;
  assign new_n4420_ = new_n2533_;
  assign new_n4421_ = new_n4420_;
  assign new_n4422_ = new_n3182_;
  assign new_n4423_ = new_n2567_;
  assign new_n4424_ = new_n4423_;
  assign new_n4425_ = new_n4423_;
  assign new_n4426_ = new_n3028_;
  assign new_n4427_ = new_n4426_;
  assign new_n4428_ = new_n4426_;
  assign new_n4429_ = new_n3187_;
  assign new_n4430_ = new_n2297_;
  assign new_n4431_ = new_n4430_;
  assign new_n4432_ = new_n4430_;
  assign new_n4433_ = new_n3192_;
  assign new_n4434_ = new_n3117_;
  assign new_n4435_ = new_n2309_;
  assign new_n4436_ = new_n4435_;
  assign new_n4437_ = new_n4435_;
  assign new_n4438_ = new_n3060_;
  assign new_n4439_ = new_n4438_;
  assign new_n4440_ = new_n3199_;
  assign new_n4441_ = new_n2317_;
  assign new_n4442_ = new_n4441_;
  assign new_n4443_ = new_n4441_;
  assign new_n4444_ = new_n3114_;
  assign new_n4445_ = new_n2323_;
  assign new_n4446_ = new_n3123_;
  assign new_n4447_ = new_n3120_;
  assign new_n4448_ = new_n3126_;
  assign new_n4449_ = new_n2386_;
  assign new_n4450_ = new_n2394_;
  assign new_n4451_ = new_n3059_;
  assign new_n4452_ = new_n3048_;
  assign new_n4453_ = new_n2778_;
  assign new_n4454_ = new_n4453_;
  assign new_n4455_ = new_n4453_;
  assign new_n4456_ = new_n3131_;
  assign new_n4457_ = new_n3104_;
  assign new_n4458_ = new_n2768_;
  assign new_n4459_ = new_n4458_;
  assign new_n4460_ = new_n3225_;
  assign new_n4461_ = new_n4460_;
  assign new_n4462_ = new_n4460_;
  assign new_n4463_ = new_n3017_;
  assign new_n4464_ = new_n3015_;
  assign new_n4465_ = new_n3230_;
  assign new_n4466_ = new_n4465_;
  assign new_n4467_ = new_n2568_;
  assign new_n4468_ = new_n3108_;
  assign new_n4469_ = new_n3107_;
  assign new_n4470_ = new_n2330_;
  assign new_n4471_ = new_n2331_;
  assign new_n4472_ = new_n2769_;
  assign new_n4473_ = new_n4472_;
  assign new_n4474_ = new_n3247_;
  assign new_n4475_ = new_n3246_;
  assign new_n4476_ = new_n2535_;
  assign new_n4477_ = new_n4476_;
  assign new_n4478_ = new_n3251_;
  assign new_n4479_ = new_n3250_;
  assign new_n4480_ = new_n3257_;
  assign new_n4481_ = new_n3254_;
  assign new_n4482_ = new_n2783_;
  assign new_n4483_ = new_n2781_;
  assign new_n4484_ = new_n3142_;
  assign new_n4485_ = new_n2378_;
  assign new_n4486_ = new_n2370_;
  assign new_n4487_ = new_n3079_;
  assign new_n4488_ = new_n3025_;
  assign new_n4489_ = new_n2459_;
  assign new_n4490_ = new_n2534_;
  assign new_n4491_ = new_n4490_;
  assign new_n4492_ = new_n2458_;
  assign new_n4493_ = new_n3287_;
  assign new_n4494_ = new_n3274_;
  assign new_n4495_ = new_n3036_;
  assign new_n4496_ = new_n3292_;
  assign new_n4497_ = new_n3151_;
  assign new_n4498_ = new_n4497_;
  assign new_n4499_ = new_n2447_;
  assign new_n4500_ = new_n2440_;
  assign new_n4501_ = new_n2446_;
  assign new_n4502_ = new_n2441_;
  assign new_n4503_ = new_n2530_;
  assign new_n4504_ = new_n2532_;
  assign new_n4505_ = new_n4504_;
  assign new_n4506_ = new_n2302_;
  assign new_n4507_ = new_n2308_;
  assign new_n4508_ = new_n4507_;
  assign new_n4509_ = new_n2453_;
  assign new_n4510_ = new_n2566_;
  assign new_n4511_ = new_n2452_;
  assign new_n4512_ = new_n2519_;
  assign new_n4513_ = new_n3229_;
  assign new_n4514_ = new_n2721_;
  assign new_n4515_ = new_n2718_;
  assign new_n4516_ = new_n2720_;
  assign new_n4517_ = new_n2719_;
  assign new_n4518_ = new_n2717_;
  assign new_n4519_ = new_n2714_;
  assign new_n4520_ = new_n2716_;
  assign new_n4521_ = new_n2715_;
  assign new_n4522_ = new_n3344_;
  assign new_n4523_ = new_n3338_;
  assign new_n4524_ = new_n3345_;
  assign new_n4525_ = new_n3339_;
  assign new_n4526_ = new_n2427_;
  assign new_n4527_ = new_n2420_;
  assign new_n4528_ = new_n2426_;
  assign new_n4529_ = new_n2421_;
  assign new_n4530_ = new_n3366_;
  assign new_n4531_ = new_n3363_;
  assign new_n4532_ = new_n2770_;
  assign new_n4533_ = new_n2771_;
  assign new_n4534_ = new_n2521_;
  assign new_n4535_ = new_n2767_;
  assign new_n4536_ = new_n3379_;
  assign new_n4537_ = new_n3373_;
  assign new_n4538_ = new_n3380_;
  assign new_n4539_ = new_n3374_;
  assign new_n4540_ = new_n3224_;
  assign new_n4541_ = new_n3103_;
  assign new_n4542_ = new_n4541_;
  assign new_n4543_ = new_n4541_;
  assign new_n4544_ = new_n2350_;
  assign new_n4545_ = new_n3102_;
  assign new_n4546_ = new_n4545_;
  assign new_n4547_ = new_n4546_;
  assign new_n4548_ = new_n4545_;
  assign new_n4549_ = new_n2276_;
  assign new_n4550_ = new_n3423_;
  assign new_n4551_ = new_n3166_;
  assign new_n4552_ = new_n4551_;
  assign new_n4553_ = new_n2575_;
  assign new_n4554_ = new_n4553_;
  assign new_n4555_ = new_n4554_;
  assign new_n4556_ = new_n4555_;
  assign new_n4557_ = new_n4555_;
  assign new_n4558_ = new_n4554_;
  assign new_n4559_ = new_n4558_;
  assign new_n4560_ = new_n4558_;
  assign new_n4561_ = new_n4553_;
  assign new_n4562_ = new_n4561_;
  assign new_n4563_ = new_n4561_;
  assign new_n4564_ = new_n2574_;
  assign new_n4565_ = new_n4564_;
  assign new_n4566_ = new_n4565_;
  assign new_n4567_ = new_n4566_;
  assign new_n4568_ = new_n4566_;
  assign new_n4569_ = new_n4565_;
  assign new_n4570_ = new_n4569_;
  assign new_n4571_ = new_n4569_;
  assign new_n4572_ = new_n4564_;
  assign new_n4573_ = new_n4572_;
  assign new_n4574_ = new_n4573_;
  assign new_n4575_ = new_n4572_;
  assign new_n4576_ = new_n2694_;
  assign new_n4577_ = new_n4576_;
  assign new_n4578_ = new_n4576_;
  assign new_n4579_ = new_n2695_;
  assign new_n4580_ = new_n4579_;
  assign new_n4581_ = new_n3402_;
  assign new_n4582_ = new_n3211_;
  assign new_n4583_ = new_n2356_;
  assign new_n4584_ = new_n2284_;
  assign new_n4585_ = new_n2362_;
  assign new_n4586_ = new_n2288_;
  assign new_n4587_ = new_n2336_;
  assign new_n4588_ = new_n2272_;
  assign new_n4589_ = new_n3157_;
  assign new_n4590_ = new_n2834_;
  assign new_n4591_ = new_n4590_;
  assign new_n4592_ = new_n4591_;
  assign new_n4593_ = new_n4590_;
  assign new_n4594_ = new_n2835_;
  assign new_n4595_ = new_n4594_;
  assign new_n4596_ = new_n4594_;
  assign new_n4597_ = new_n2399_;
  assign new_n4598_ = new_n2398_;
  assign new_n4599_ = new_n4598_;
  assign new_n4600_ = new_n2219_;
  assign new_n4601_ = new_n2218_;
  assign new_n4602_ = new_n4601_;
  assign new_n4603_ = new_n3507_;
  assign new_n4604_ = new_n3503_;
  assign new_n4605_ = new_n2269_;
  assign new_n4606_ = new_n2347_;
  assign new_n4607_ = new_n4606_;
  assign new_n4608_ = new_n2845_;
  assign new_n4609_ = new_n2861_;
  assign new_n4610_ = new_n2864_;
  assign new_n4611_ = new_n2869_;
  assign new_n4612_ = new_n2949_;
  assign new_n4613_ = new_n2975_;
  assign new_n4614_ = new_n3012_;
  assign new_n4615_ = 1'b0;
  always @ (posedge clock) begin
    n1416_lo <= n4649_li000_li000;
    n1419_lo <= n4652_li001_li001;
    n1422_lo <= n4655_li002_li002;
    n1425_lo <= n4658_li003_li003;
    n1428_lo <= n4661_li004_li004;
    n1431_lo <= n4664_li005_li005;
    n1434_lo <= n4667_li006_li006;
    n1437_lo <= n4670_li007_li007;
    n1440_lo <= n4673_li008_li008;
    n1443_lo <= n4676_li009_li009;
    n1446_lo <= n4679_li010_li010;
    n1449_lo <= n4682_li011_li011;
    n1452_lo <= n4685_li012_li012;
    n1455_lo <= n4688_li013_li013;
    n1458_lo <= n4691_li014_li014;
    n1464_lo <= n4697_li016_li016;
    n1467_lo <= n4700_li017_li017;
    n1470_lo <= n4703_li018_li018;
    n1476_lo <= n4709_li020_li020;
    n1479_lo <= n4712_li021_li021;
    n1482_lo <= n4715_li022_li022;
    n1488_lo <= n4721_li024_li024;
    n1491_lo <= n4724_li025_li025;
    n1494_lo <= n4727_li026_li026;
    n1497_lo <= n4730_li027_li027;
    n1500_lo <= n4733_li028_li028;
    n1503_lo <= n4736_li029_li029;
    n1512_lo <= n4745_li032_li032;
    n1515_lo <= n4748_li033_li033;
    n1518_lo <= n4751_li034_li034;
    n1521_lo <= n4754_li035_li035;
    n1524_lo <= n4757_li036_li036;
    n1527_lo <= n4760_li037_li037;
    n1530_lo <= n4763_li038_li038;
    n1533_lo <= n4766_li039_li039;
    n1536_lo <= n4769_li040_li040;
    n1539_lo <= n4772_li041_li041;
    n1542_lo <= n4775_li042_li042;
    n1545_lo <= n4778_li043_li043;
    n1548_lo <= n4781_li044_li044;
    n1551_lo <= n4784_li045_li045;
    n1554_lo <= n4787_li046_li046;
    n1560_lo <= n4793_li048_li048;
    n1563_lo <= n4796_li049_li049;
    n1566_lo <= n4799_li050_li050;
    n1572_lo <= n4805_li052_li052;
    n1575_lo <= n4808_li053_li053;
    n1578_lo <= n4811_li054_li054;
    n1584_lo <= n4817_li056_li056;
    n1587_lo <= n4820_li057_li057;
    n1590_lo <= n4823_li058_li058;
    n1596_lo <= n4829_li060_li060;
    n1599_lo <= n4832_li061_li061;
    n1602_lo <= n4835_li062_li062;
    n1608_lo <= n4841_li064_li064;
    n1611_lo <= n4844_li065_li065;
    n1614_lo <= n4847_li066_li066;
    n1620_lo <= n4853_li068_li068;
    n1623_lo <= n4856_li069_li069;
    n1626_lo <= n4859_li070_li070;
    n1632_lo <= n4865_li072_li072;
    n1635_lo <= n4868_li073_li073;
    n1638_lo <= n4871_li074_li074;
    n1644_lo <= n4877_li076_li076;
    n1647_lo <= n4880_li077_li077;
    n1650_lo <= n4883_li078_li078;
    n1656_lo <= n4889_li080_li080;
    n1659_lo <= n4892_li081_li081;
    n1662_lo <= n4895_li082_li082;
    n1668_lo <= n4901_li084_li084;
    n1671_lo <= n4904_li085_li085;
    n1674_lo <= n4907_li086_li086;
    n1680_lo <= n4913_li088_li088;
    n1683_lo <= n4916_li089_li089;
    n1686_lo <= n4919_li090_li090;
    n1692_lo <= n4925_li092_li092;
    n1695_lo <= n4928_li093_li093;
    n1698_lo <= n4931_li094_li094;
    n1704_lo <= n4937_li096_li096;
    n1707_lo <= n4940_li097_li097;
    n1710_lo <= n4943_li098_li098;
    n1716_lo <= n4949_li100_li100;
    n1719_lo <= n4952_li101_li101;
    n1722_lo <= n4955_li102_li102;
    n1728_lo <= n4961_li104_li104;
    n1731_lo <= n4964_li105_li105;
    n1734_lo <= n4967_li106_li106;
    n1740_lo <= n4973_li108_li108;
    n1743_lo <= n4976_li109_li109;
    n1746_lo <= n4979_li110_li110;
    n1749_lo <= n4982_li111_li111;
    n1752_lo <= n4985_li112_li112;
    n1755_lo <= n4988_li113_li113;
    n1758_lo <= n4991_li114_li114;
    n1761_lo <= n4994_li115_li115;
    n1764_lo <= n4997_li116_li116;
    n1776_lo <= n5009_li120_li120;
    n1788_lo <= n5021_li124_li124;
    n1791_lo <= n5024_li125_li125;
    n1794_lo <= n5027_li126_li126;
    n1797_lo <= n5030_li127_li127;
    n1800_lo <= n5033_li128_li128;
    n1803_lo <= n5036_li129_li129;
    n1812_lo <= n5045_li132_li132;
    n1815_lo <= n5048_li133_li133;
    n1824_lo <= n5057_li136_li136;
    n1827_lo <= n5060_li137_li137;
    n1836_lo <= n5069_li140_li140;
    n1839_lo <= n5072_li141_li141;
    n1848_lo <= n5081_li144_li144;
    n1851_lo <= n5084_li145_li145;
    n1860_lo <= n5093_li148_li148;
    n1872_lo <= n5105_li152_li152;
    n1875_lo <= n5108_li153_li153;
    n1884_lo <= n5117_li156_li156;
    n1896_lo <= n5129_li160_li160;
    n1899_lo <= n5132_li161_li161;
    n1908_lo <= n5141_li164_li164;
    n1920_lo <= n5153_li168_li168;
    n1923_lo <= n5156_li169_li169;
    n1926_lo <= n5159_li170_li170;
    n1929_lo <= n5162_li171_li171;
    n1932_lo <= n5165_li172_li172;
    n1935_lo <= n5168_li173_li173;
    n1944_lo <= n5177_li176_li176;
    n1947_lo <= n5180_li177_li177;
    n1956_lo <= n5189_li180_li180;
    n1959_lo <= n5192_li181_li181;
    n1962_lo <= n5195_li182_li182;
    n1968_lo <= n5201_li184_li184;
    n1971_lo <= n5204_li185_li185;
    n1980_lo <= n5213_li188_li188;
    n1983_lo <= n5216_li189_li189;
    n1992_lo <= n5225_li192_li192;
    n1995_lo <= n5228_li193_li193;
    n2004_lo <= n5237_li196_li196;
    n2016_lo <= n5249_li200_li200;
    n2019_lo <= n5252_li201_li201;
    n2028_lo <= n5261_li204_li204;
    n2040_lo <= n5273_li208_li208;
    n2043_lo <= n5276_li209_li209;
    n2046_lo <= n5279_li210_li210;
    n2049_lo <= n5282_li211_li211;
    n2052_lo <= n5285_li212_li212;
    n2055_lo <= n5288_li213_li213;
    n2064_lo <= n5297_li216_li216;
    n2067_lo <= n5300_li217_li217;
    n2076_lo <= n5309_li220_li220;
    n2079_lo <= n5312_li221_li221;
    n2088_lo <= n5321_li224_li224;
    n2091_lo <= n5324_li225_li225;
    n2100_lo <= n5333_li228_li228;
    n2103_lo <= n5336_li229_li229;
    n2112_lo <= n5345_li232_li232;
    n2115_lo <= n5348_li233_li233;
    n2124_lo <= n5357_li236_li236;
    n2127_lo <= n5360_li237_li237;
    n2136_lo <= n5369_li240_li240;
    n2148_lo <= n5381_li244_li244;
    n2151_lo <= n5384_li245_li245;
    n2160_lo <= n5393_li248_li248;
    n2172_lo <= n5405_li252_li252;
    n2175_lo <= n5408_li253_li253;
    n2178_lo <= n5411_li254_li254;
    n2181_lo <= n5414_li255_li255;
    n2184_lo <= n5417_li256_li256;
    n2187_lo <= n5420_li257_li257;
    n2196_lo <= n5429_li260_li260;
    n2199_lo <= n5432_li261_li261;
    n2208_lo <= n5441_li264_li264;
    n2211_lo <= n5444_li265_li265;
    n2220_lo <= n5453_li268_li268;
    n2223_lo <= n5456_li269_li269;
    n2232_lo <= n5465_li272_li272;
    n2235_lo <= n5468_li273_li273;
    n2244_lo <= n5477_li276_li276;
    n2247_lo <= n5480_li277_li277;
    n2256_lo <= n5489_li280_li280;
    n2259_lo <= n5492_li281_li281;
    n2268_lo <= n5501_li284_li284;
    n2280_lo <= n5513_li288_li288;
    n2283_lo <= n5516_li289_li289;
    n2292_lo <= n5525_li292_li292;
    n2295_lo <= n5528_li293_li293;
    n2298_lo <= n5531_li294_li294;
    n2301_lo <= n5534_li295_li295;
    n2304_lo <= n5537_li296_li296;
    n2307_lo <= n5540_li297_li297;
    n2316_lo <= n5549_li300_li300;
    n2319_lo <= n5552_li301_li301;
    n2322_lo <= n5555_li302_li302;
    n2325_lo <= n5558_li303_li303;
    n2328_lo <= n5561_li304_li304;
    n2331_lo <= n5564_li305_li305;
    n2340_lo <= n5573_li308_li308;
    n2343_lo <= n5576_li309_li309;
    n2376_lo <= n5609_li320_li320;
    n2379_lo <= n5612_li321_li321;
    n2388_lo <= n5621_li324_li324;
    n2391_lo <= n5624_li325_li325;
    n2400_lo <= n5633_li328_li328;
    n2403_lo <= n5636_li329_li329;
    n2412_lo <= n5645_li332_li332;
    n2415_lo <= n5648_li333_li333;
    n2424_lo <= n5657_li336_li336;
    n2427_lo <= n5660_li337_li337;
    n2436_lo <= n5669_li340_li340;
    n2439_lo <= n5672_li341_li341;
    n2442_lo <= n5675_li342_li342;
    n2445_lo <= n5678_li343_li343;
    n2448_lo <= n5681_li344_li344;
    n2451_lo <= n5684_li345_li345;
    n2460_lo <= n5693_li348_li348;
    n2463_lo <= n5696_li349_li349;
    n2496_lo <= n5729_li360_li360;
    n2499_lo <= n5732_li361_li361;
    n2508_lo <= n5741_li364_li364;
    n2511_lo <= n5744_li365_li365;
    n2520_lo <= n5753_li368_li368;
    n2523_lo <= n5756_li369_li369;
    n2532_lo <= n5765_li372_li372;
    n2535_lo <= n5768_li373_li373;
    n2544_lo <= n5777_li376_li376;
    n2547_lo <= n5780_li377_li377;
    n2556_lo <= n5789_li380_li380;
    n2559_lo <= n5792_li381_li381;
    n2562_lo <= n5795_li382_li382;
    n2565_lo <= n5798_li383_li383;
    n2568_lo <= n5801_li384_li384;
    n2571_lo <= n5804_li385_li385;
    n2580_lo <= n5813_li388_li388;
    n2583_lo <= n5816_li389_li389;
    n2616_lo <= n5849_li400_li400;
    n2619_lo <= n5852_li401_li401;
    n2628_lo <= n5861_li404_li404;
    n2631_lo <= n5864_li405_li405;
    n2640_lo <= n5873_li408_li408;
    n2643_lo <= n5876_li409_li409;
    n2652_lo <= n5885_li412_li412;
    n2655_lo <= n5888_li413_li413;
    n2664_lo <= n5897_li416_li416;
    n2667_lo <= n5900_li417_li417;
    n2676_lo <= n5909_li420_li420;
    n2679_lo <= n5912_li421_li421;
    n2682_lo <= n5915_li422_li422;
    n2685_lo <= n5918_li423_li423;
    n2688_lo <= n5921_li424_li424;
    n2691_lo <= n5924_li425_li425;
    n2700_lo <= n5933_li428_li428;
    n2703_lo <= n5936_li429_li429;
    n2736_lo <= n5969_li440_li440;
    n2739_lo <= n5972_li441_li441;
    n2748_lo <= n5981_li444_li444;
    n2751_lo <= n5984_li445_li445;
    n2760_lo <= n5993_li448_li448;
    n2763_lo <= n5996_li449_li449;
    n2772_lo <= n6005_li452_li452;
    n2775_lo <= n6008_li453_li453;
    n2784_lo <= n6017_li456_li456;
    n2787_lo <= n6020_li457_li457;
    n2790_lo <= n6023_li458_li458;
    n2793_lo <= n6026_li459_li459;
    n2796_lo <= n6029_li460_li460;
    n2799_lo <= n6032_li461_li461;
    n2802_lo <= n6035_li462_li462;
    n2805_lo <= n6038_li463_li463;
    n2808_lo <= n6041_li464_li464;
    n2820_lo <= n6053_li468_li468;
    n2823_lo <= n6056_li469_li469;
    n2826_lo <= n6059_li470_li470;
    n2829_lo <= n6062_li471_li471;
    n2832_lo <= n6065_li472_li472;
    n2835_lo <= n6068_li473_li473;
    n2838_lo <= n6071_li474_li474;
    n2841_lo <= n6074_li475_li475;
    n2844_lo <= n6077_li476_li476;
    n2856_lo <= n6089_li480_li480;
    n2859_lo <= n6092_li481_li481;
    n2862_lo <= n6095_li482_li482;
    n2865_lo <= n6098_li483_li483;
    n2868_lo <= n6101_li484_li484;
    n2871_lo <= n6104_li485_li485;
    n2874_lo <= n6107_li486_li486;
    n2877_lo <= n6110_li487_li487;
    n2880_lo <= n6113_li488_li488;
    n2883_lo <= n6116_li489_li489;
    n2886_lo <= n6119_li490_li490;
    n2889_lo <= n6122_li491_li491;
    n2892_lo <= n6125_li492_li492;
    n2895_lo <= n6128_li493_li493;
    n2898_lo <= n6131_li494_li494;
    n2901_lo <= n6134_li495_li495;
    n2904_lo <= n6137_li496_li496;
    n2907_lo <= n6140_li497_li497;
    n2916_lo <= n6149_li500_li500;
    n2919_lo <= n6152_li501_li501;
    n2925_lo <= n6158_li503_li503;
    n2928_lo <= n6161_li504_li504;
    n2940_lo <= n6173_li508_li508;
    n2943_lo <= n6176_li509_li509;
    n2952_lo <= n6185_li512_li512;
    n2955_lo <= n6188_li513_li513;
    n2961_lo <= n6194_li515_li515;
    n2964_lo <= n6197_li516_li516;
    n2967_lo <= n6200_li517_li517;
    n2970_lo <= n6203_li518_li518;
    n2976_lo <= n6209_li520_li520;
    n2979_lo <= n6212_li521_li521;
    n2982_lo <= n6215_li522_li522;
    n2988_lo <= n6221_li524_li524;
    n2991_lo <= n6224_li525_li525;
    n2994_lo <= n6227_li526_li526;
    n2997_lo <= n6230_li527_li527;
    n3000_lo <= n6233_li528_li528;
    n3003_lo <= n6236_li529_li529;
    n3006_lo <= n6239_li530_li530;
    n3012_lo <= n6245_li532_li532;
    n3015_lo <= n6248_li533_li533;
    n3018_lo <= n6251_li534_li534;
    n3021_lo <= n6254_li535_li535;
    n3024_lo <= n6257_li536_li536;
    n3027_lo <= n6260_li537_li537;
    n3030_lo <= n6263_li538_li538;
    n3033_lo <= n6266_li539_li539;
    n3036_lo <= n6269_li540_li540;
    n3039_lo <= n6272_li541_li541;
    n3045_lo <= n6278_li543_li543;
    n3048_lo <= n6281_li544_li544;
    n3051_lo <= n6284_li545_li545;
    n3054_lo <= n6287_li546_li546;
    n3057_lo <= n6290_li547_li547;
    n3060_lo <= n6293_li548_li548;
    n3063_lo <= n6296_li549_li549;
    n3069_lo <= n6302_li551_li551;
    n3072_lo <= n6305_li552_li552;
    n3075_lo <= n6308_li553_li553;
    n3081_lo <= n6314_li555_li555;
    n3084_lo <= n6317_li556_li556;
    n3087_lo <= n6320_li557_li557;
    n3093_lo <= n6326_li559_li559;
    n3096_lo <= n6329_li560_li560;
    n3099_lo <= n6332_li561_li561;
    n3102_lo <= n6335_li562_li562;
    n3105_lo <= n6338_li563_li563;
    n3108_lo <= n6341_li564_li564;
    n3111_lo <= n6344_li565_li565;
    n3114_lo <= n6347_li566_li566;
    n3117_lo <= n6350_li567_li567;
    n3120_lo <= n6353_li568_li568;
    n3123_lo <= n6356_li569_li569;
    n3126_lo <= n6359_li570_li570;
    n3129_lo <= n6362_li571_li571;
    n3132_lo <= n6365_li572_li572;
    n3135_lo <= n6368_li573_li573;
    n3138_lo <= n6371_li574_li574;
    n3141_lo <= n6374_li575_li575;
    n3156_lo <= n6389_li580_li580;
    n3168_lo <= n6401_li584_li584;
    n3171_lo <= n6404_li585_li585;
    n3174_lo <= n6407_li586_li586;
    n3177_lo <= n6410_li587_li587;
    n3180_lo <= n6413_li588_li588;
    n3183_lo <= n6416_li589_li589;
    n3192_lo <= n6425_li592_li592;
    n3195_lo <= n6428_li593_li593;
    n3204_lo <= n6437_li596_li596;
    n3207_lo <= n6440_li597_li597;
    n3210_lo <= n6443_li598_li598;
    n3216_lo <= n6449_li600_li600;
    n3219_lo <= n6452_li601_li601;
    n3222_lo <= n6455_li602_li602;
    n3228_lo <= n6461_li604_li604;
    n3231_lo <= n6464_li605_li605;
    n3240_lo <= n6473_li608_li608;
    n3243_lo <= n6476_li609_li609;
    n3252_lo <= n6485_li612_li612;
    n3255_lo <= n6488_li613_li613;
    n3258_lo <= n6491_li614_li614;
    n3264_lo <= n6497_li616_li616;
    n3267_lo <= n6500_li617_li617;
    n3270_lo <= n6503_li618_li618;
    n3276_lo <= n6509_li620_li620;
    n3279_lo <= n6512_li621_li621;
    n3282_lo <= n6515_li622_li622;
    n3288_lo <= n6521_li624_li624;
    n3291_lo <= n6524_li625_li625;
    n3294_lo <= n6527_li626_li626;
    n3603_o2 <= n3603_i2;
    n3604_o2 <= n3604_i2;
    n1391_inv <= n3618_i2;
    n3798_o2 <= n3798_i2;
    n3846_o2 <= n3846_i2;
    n4019_o2 <= n4019_i2;
    n4017_o2 <= n4017_i2;
    n2177_o2 <= n2177_i2;
    n2150_o2 <= n2150_i2;
    n2154_o2 <= n2154_i2;
    n2184_o2 <= n2184_i2;
    n2515_o2 <= n2515_i2;
    n3837_o2 <= n3837_i2;
    n2167_o2 <= n2167_i2;
    n2118_o2 <= n2118_i2;
    n2186_o2 <= n2186_i2;
    n2174_o2 <= n2174_i2;
    n3964_o2 <= n3964_i2;
    n4005_o2 <= n4005_i2;
    n4006_o2 <= n4006_i2;
    n1445_inv <= n2195_i2;
    n2176_o2 <= n2176_i2;
    n2227_o2 <= n2227_i2;
    n2236_o2 <= n2236_i2;
    n2245_o2 <= n2245_i2;
    n2518_o2 <= n2518_i2;
    n4023_o2 <= n4023_i2;
    n1466_inv <= n4024_i2;
    n4038_o2 <= n4038_i2;
    n4039_o2 <= n4039_i2;
    n1475_inv <= n4040_i2;
    n2119_o2 <= n2119_i2;
    n2275_o2 <= n2275_i2;
    n2595_o2 <= n2595_i2;
    n2594_o2 <= n2594_i2;
    lo498_buf_o2 <= lo498_buf_i2;
    lo502_buf_o2 <= lo502_buf_i2;
    lo550_buf_o2 <= lo550_buf_i2;
    n2596_o2 <= n2596_i2;
    n2593_o2 <= n2593_i2;
    n2668_o2 <= n2668_i2;
    lo542_buf_o2 <= lo542_buf_i2;
    n2667_o2 <= n2667_i2;
    n2404_o2 <= n2404_i2;
    n2410_o2 <= n2410_i2;
    n2419_o2 <= n2419_i2;
    n2392_o2 <= n2392_i2;
    n2369_o2 <= n2369_i2;
    n2397_o2 <= n2397_i2;
    n2601_o2 <= n2601_i2;
    n2658_o2 <= n2658_i2;
    n2574_o2 <= n2574_i2;
    n2205_o2 <= n2205_i2;
    lo510_buf_o2 <= lo510_buf_i2;
    lo514_buf_o2 <= lo514_buf_i2;
    lo554_buf_o2 <= lo554_buf_i2;
    lo558_buf_o2 <= lo558_buf_i2;
    lo578_buf_o2 <= lo578_buf_i2;
    n2254_o2 <= n2254_i2;
    n2421_o2 <= n2421_i2;
    n2422_o2 <= n2422_i2;
    n2130_o2 <= n2130_i2;
    n2127_o2 <= n2127_i2;
    n2131_o2 <= n2131_i2;
    n2128_o2 <= n2128_i2;
    n2264_o2 <= n2264_i2;
    n2467_o2 <= n2467_i2;
    n2471_o2 <= n2471_i2;
    n2488_o2 <= n2488_i2;
    n2478_o2 <= n2478_i2;
    n2486_o2 <= n2486_i2;
    n2485_o2 <= n2485_i2;
    n2498_o2 <= n2498_i2;
    n2495_o2 <= n2495_i2;
    n2496_o2 <= n2496_i2;
    n2458_o2 <= n2458_i2;
    n2643_o2 <= n2643_i2;
    n2462_o2 <= n2462_i2;
    n2468_o2 <= n2468_i2;
    n2639_o2 <= n2639_i2;
    n2499_o2 <= n2499_i2;
    n2472_o2 <= n2472_i2;
    n2474_o2 <= n2474_i2;
    n2489_o2 <= n2489_i2;
    n2321_o2 <= n2321_i2;
    n2322_o2 <= n2322_i2;
    n2640_o2 <= n2640_i2;
    n2642_o2 <= n2642_i2;
    n2187_o2 <= n2187_i2;
    n2373_o2 <= n2373_i2;
    n2603_o2 <= n2603_i2;
    n2388_o2 <= n2388_i2;
    n2437_o2 <= n2437_i2;
    n2356_o2 <= n2356_i2;
    n2452_o2 <= n2452_i2;
    n2347_o2 <= n2347_i2;
    n2329_o2 <= n2329_i2;
    n2669_o2 <= n2669_i2;
    n2332_o2 <= n2332_i2;
    n2664_o2 <= n2664_i2;
    n2665_o2 <= n2665_i2;
    n2653_o2 <= n2653_i2;
    n2654_o2 <= n2654_i2;
    n2636_o2 <= n2636_i2;
    n2660_o2 <= n2660_i2;
    n2318_o2 <= n2318_i2;
    n2319_o2 <= n2319_i2;
    n2586_o2 <= n2586_i2;
    n2587_o2 <= n2587_i2;
    n2288_o2 <= n2288_i2;
    n2344_o2 <= n2344_i2;
    n2530_o2 <= n2530_i2;
    n2303_o2 <= n2303_i2;
    n2566_o2 <= n2566_i2;
    n2567_o2 <= n2567_i2;
    n2554_o2 <= n2554_i2;
    n2194_o2 <= n2194_i2;
    lo582_buf_o2 <= lo582_buf_i2;
    lo030_buf_o2 <= lo030_buf_i2;
    lo174_buf_o2 <= lo174_buf_i2;
    lo178_buf_o2 <= lo178_buf_i2;
    lo186_buf_o2 <= lo186_buf_i2;
    lo266_buf_o2 <= lo266_buf_i2;
    lo306_buf_o2 <= lo306_buf_i2;
    lo346_buf_o2 <= lo346_buf_i2;
    lo386_buf_o2 <= lo386_buf_i2;
    lo426_buf_o2 <= lo426_buf_i2;
    lo590_buf_o2 <= lo590_buf_i2;
    lo594_buf_o2 <= lo594_buf_i2;
    lo606_buf_o2 <= lo606_buf_i2;
    lo610_buf_o2 <= lo610_buf_i2;
    n2238_o2 <= n2238_i2;
    n2229_o2 <= n2229_i2;
    n2242_o2 <= n2242_i2;
    n2233_o2 <= n2233_i2;
    n2168_o2 <= n2168_i2;
    n2237_o2 <= n2237_i2;
    n2228_o2 <= n2228_i2;
    n2172_o2 <= n2172_i2;
    n2223_o2 <= n2223_i2;
    n2222_o2 <= n2222_i2;
    n2170_o2 <= n2170_i2;
    n2181_o2 <= n2181_i2;
    n2510_o2 <= n2510_i2;
    n2621_o2 <= n2621_i2;
    lo466_buf_o2 <= lo466_buf_i2;
    lo478_buf_o2 <= lo478_buf_i2;
    n2149_o2 <= n2149_i2;
    n2429_o2 <= n2429_i2;
    n2444_o2 <= n2444_i2;
    n2153_o2 <= n2153_i2;
    n2433_o2 <= n2433_i2;
    n2448_o2 <= n2448_i2;
    n2367_o2 <= n2367_i2;
    n2386_o2 <= n2386_i2;
    n2539_o2 <= n2539_i2;
    n2183_o2 <= n2183_i2;
    n2220_o2 <= n2220_i2;
    n2514_o2 <= n2514_i2;
    n2196_o2 <= n2196_i2;
    n2616_o2 <= n2616_i2;
    n2612_o2 <= n2612_i2;
    n2627_o2 <= n2627_i2;
    n2140_o2 <= n2140_i2;
    n1877_inv <= n2144_i2;
    lo149_buf_o2 <= lo149_buf_i2;
    lo197_buf_o2 <= lo197_buf_i2;
    lo118_buf_o2 <= lo118_buf_i2;
    lo158_buf_o2 <= lo158_buf_i2;
    lo166_buf_o2 <= lo166_buf_i2;
    lo242_buf_o2 <= lo242_buf_i2;
    lo286_buf_o2 <= lo286_buf_i2;
    lo506_buf_o2 <= lo506_buf_i2;
    n2198_o2 <= n2198_i2;
    n2202_o2 <= n2202_i2;
    n2197_o2 <= n2197_i2;
    n1913_inv <= n2166_i2;
    n2146_o2 <= n2146_i2;
    n1919_inv <= n2165_i2;
    lo312_buf_o2 <= lo312_buf_i2;
    lo316_buf_o2 <= lo316_buf_i2;
    lo352_buf_o2 <= lo352_buf_i2;
    lo356_buf_o2 <= lo356_buf_i2;
    lo392_buf_o2 <= lo392_buf_i2;
    lo396_buf_o2 <= lo396_buf_i2;
    lo432_buf_o2 <= lo432_buf_i2;
    lo436_buf_o2 <= lo436_buf_i2;
    lo576_buf_o2 <= lo576_buf_i2;
  end
  initial begin
    n1416_lo <= 1'b0;
    n1419_lo <= 1'b0;
    n1422_lo <= 1'b0;
    n1425_lo <= 1'b0;
    n1428_lo <= 1'b0;
    n1431_lo <= 1'b0;
    n1434_lo <= 1'b0;
    n1437_lo <= 1'b0;
    n1440_lo <= 1'b0;
    n1443_lo <= 1'b0;
    n1446_lo <= 1'b0;
    n1449_lo <= 1'b0;
    n1452_lo <= 1'b0;
    n1455_lo <= 1'b0;
    n1458_lo <= 1'b0;
    n1464_lo <= 1'b0;
    n1467_lo <= 1'b0;
    n1470_lo <= 1'b0;
    n1476_lo <= 1'b0;
    n1479_lo <= 1'b0;
    n1482_lo <= 1'b0;
    n1488_lo <= 1'b0;
    n1491_lo <= 1'b0;
    n1494_lo <= 1'b0;
    n1497_lo <= 1'b0;
    n1500_lo <= 1'b0;
    n1503_lo <= 1'b0;
    n1512_lo <= 1'b0;
    n1515_lo <= 1'b0;
    n1518_lo <= 1'b0;
    n1521_lo <= 1'b0;
    n1524_lo <= 1'b0;
    n1527_lo <= 1'b0;
    n1530_lo <= 1'b0;
    n1533_lo <= 1'b0;
    n1536_lo <= 1'b0;
    n1539_lo <= 1'b0;
    n1542_lo <= 1'b0;
    n1545_lo <= 1'b0;
    n1548_lo <= 1'b0;
    n1551_lo <= 1'b0;
    n1554_lo <= 1'b0;
    n1560_lo <= 1'b0;
    n1563_lo <= 1'b0;
    n1566_lo <= 1'b0;
    n1572_lo <= 1'b0;
    n1575_lo <= 1'b0;
    n1578_lo <= 1'b0;
    n1584_lo <= 1'b0;
    n1587_lo <= 1'b0;
    n1590_lo <= 1'b0;
    n1596_lo <= 1'b0;
    n1599_lo <= 1'b0;
    n1602_lo <= 1'b0;
    n1608_lo <= 1'b0;
    n1611_lo <= 1'b0;
    n1614_lo <= 1'b0;
    n1620_lo <= 1'b0;
    n1623_lo <= 1'b0;
    n1626_lo <= 1'b0;
    n1632_lo <= 1'b0;
    n1635_lo <= 1'b0;
    n1638_lo <= 1'b0;
    n1644_lo <= 1'b0;
    n1647_lo <= 1'b0;
    n1650_lo <= 1'b0;
    n1656_lo <= 1'b0;
    n1659_lo <= 1'b0;
    n1662_lo <= 1'b0;
    n1668_lo <= 1'b0;
    n1671_lo <= 1'b0;
    n1674_lo <= 1'b0;
    n1680_lo <= 1'b0;
    n1683_lo <= 1'b0;
    n1686_lo <= 1'b0;
    n1692_lo <= 1'b0;
    n1695_lo <= 1'b0;
    n1698_lo <= 1'b0;
    n1704_lo <= 1'b0;
    n1707_lo <= 1'b0;
    n1710_lo <= 1'b0;
    n1716_lo <= 1'b0;
    n1719_lo <= 1'b0;
    n1722_lo <= 1'b0;
    n1728_lo <= 1'b0;
    n1731_lo <= 1'b0;
    n1734_lo <= 1'b0;
    n1740_lo <= 1'b0;
    n1743_lo <= 1'b0;
    n1746_lo <= 1'b0;
    n1749_lo <= 1'b0;
    n1752_lo <= 1'b0;
    n1755_lo <= 1'b0;
    n1758_lo <= 1'b0;
    n1761_lo <= 1'b0;
    n1764_lo <= 1'b0;
    n1776_lo <= 1'b0;
    n1788_lo <= 1'b0;
    n1791_lo <= 1'b0;
    n1794_lo <= 1'b0;
    n1797_lo <= 1'b0;
    n1800_lo <= 1'b0;
    n1803_lo <= 1'b0;
    n1812_lo <= 1'b0;
    n1815_lo <= 1'b0;
    n1824_lo <= 1'b0;
    n1827_lo <= 1'b0;
    n1836_lo <= 1'b0;
    n1839_lo <= 1'b0;
    n1848_lo <= 1'b0;
    n1851_lo <= 1'b0;
    n1860_lo <= 1'b0;
    n1872_lo <= 1'b0;
    n1875_lo <= 1'b0;
    n1884_lo <= 1'b0;
    n1896_lo <= 1'b0;
    n1899_lo <= 1'b0;
    n1908_lo <= 1'b0;
    n1920_lo <= 1'b0;
    n1923_lo <= 1'b0;
    n1926_lo <= 1'b0;
    n1929_lo <= 1'b0;
    n1932_lo <= 1'b0;
    n1935_lo <= 1'b0;
    n1944_lo <= 1'b0;
    n1947_lo <= 1'b0;
    n1956_lo <= 1'b0;
    n1959_lo <= 1'b0;
    n1962_lo <= 1'b0;
    n1968_lo <= 1'b0;
    n1971_lo <= 1'b0;
    n1980_lo <= 1'b0;
    n1983_lo <= 1'b0;
    n1992_lo <= 1'b0;
    n1995_lo <= 1'b0;
    n2004_lo <= 1'b0;
    n2016_lo <= 1'b0;
    n2019_lo <= 1'b0;
    n2028_lo <= 1'b0;
    n2040_lo <= 1'b0;
    n2043_lo <= 1'b0;
    n2046_lo <= 1'b0;
    n2049_lo <= 1'b0;
    n2052_lo <= 1'b0;
    n2055_lo <= 1'b0;
    n2064_lo <= 1'b0;
    n2067_lo <= 1'b0;
    n2076_lo <= 1'b0;
    n2079_lo <= 1'b0;
    n2088_lo <= 1'b0;
    n2091_lo <= 1'b0;
    n2100_lo <= 1'b0;
    n2103_lo <= 1'b0;
    n2112_lo <= 1'b0;
    n2115_lo <= 1'b0;
    n2124_lo <= 1'b0;
    n2127_lo <= 1'b0;
    n2136_lo <= 1'b0;
    n2148_lo <= 1'b0;
    n2151_lo <= 1'b0;
    n2160_lo <= 1'b0;
    n2172_lo <= 1'b0;
    n2175_lo <= 1'b0;
    n2178_lo <= 1'b0;
    n2181_lo <= 1'b0;
    n2184_lo <= 1'b0;
    n2187_lo <= 1'b0;
    n2196_lo <= 1'b0;
    n2199_lo <= 1'b0;
    n2208_lo <= 1'b0;
    n2211_lo <= 1'b0;
    n2220_lo <= 1'b0;
    n2223_lo <= 1'b0;
    n2232_lo <= 1'b0;
    n2235_lo <= 1'b0;
    n2244_lo <= 1'b0;
    n2247_lo <= 1'b0;
    n2256_lo <= 1'b0;
    n2259_lo <= 1'b0;
    n2268_lo <= 1'b0;
    n2280_lo <= 1'b0;
    n2283_lo <= 1'b0;
    n2292_lo <= 1'b0;
    n2295_lo <= 1'b0;
    n2298_lo <= 1'b0;
    n2301_lo <= 1'b0;
    n2304_lo <= 1'b0;
    n2307_lo <= 1'b0;
    n2316_lo <= 1'b0;
    n2319_lo <= 1'b0;
    n2322_lo <= 1'b0;
    n2325_lo <= 1'b0;
    n2328_lo <= 1'b0;
    n2331_lo <= 1'b0;
    n2340_lo <= 1'b0;
    n2343_lo <= 1'b0;
    n2376_lo <= 1'b0;
    n2379_lo <= 1'b0;
    n2388_lo <= 1'b0;
    n2391_lo <= 1'b0;
    n2400_lo <= 1'b0;
    n2403_lo <= 1'b0;
    n2412_lo <= 1'b0;
    n2415_lo <= 1'b0;
    n2424_lo <= 1'b0;
    n2427_lo <= 1'b0;
    n2436_lo <= 1'b0;
    n2439_lo <= 1'b0;
    n2442_lo <= 1'b0;
    n2445_lo <= 1'b0;
    n2448_lo <= 1'b0;
    n2451_lo <= 1'b0;
    n2460_lo <= 1'b0;
    n2463_lo <= 1'b0;
    n2496_lo <= 1'b0;
    n2499_lo <= 1'b0;
    n2508_lo <= 1'b0;
    n2511_lo <= 1'b0;
    n2520_lo <= 1'b0;
    n2523_lo <= 1'b0;
    n2532_lo <= 1'b0;
    n2535_lo <= 1'b0;
    n2544_lo <= 1'b0;
    n2547_lo <= 1'b0;
    n2556_lo <= 1'b0;
    n2559_lo <= 1'b0;
    n2562_lo <= 1'b0;
    n2565_lo <= 1'b0;
    n2568_lo <= 1'b0;
    n2571_lo <= 1'b0;
    n2580_lo <= 1'b0;
    n2583_lo <= 1'b0;
    n2616_lo <= 1'b0;
    n2619_lo <= 1'b0;
    n2628_lo <= 1'b0;
    n2631_lo <= 1'b0;
    n2640_lo <= 1'b0;
    n2643_lo <= 1'b0;
    n2652_lo <= 1'b0;
    n2655_lo <= 1'b0;
    n2664_lo <= 1'b0;
    n2667_lo <= 1'b0;
    n2676_lo <= 1'b0;
    n2679_lo <= 1'b0;
    n2682_lo <= 1'b0;
    n2685_lo <= 1'b0;
    n2688_lo <= 1'b0;
    n2691_lo <= 1'b0;
    n2700_lo <= 1'b0;
    n2703_lo <= 1'b0;
    n2736_lo <= 1'b0;
    n2739_lo <= 1'b0;
    n2748_lo <= 1'b0;
    n2751_lo <= 1'b0;
    n2760_lo <= 1'b0;
    n2763_lo <= 1'b0;
    n2772_lo <= 1'b0;
    n2775_lo <= 1'b0;
    n2784_lo <= 1'b0;
    n2787_lo <= 1'b0;
    n2790_lo <= 1'b0;
    n2793_lo <= 1'b0;
    n2796_lo <= 1'b0;
    n2799_lo <= 1'b0;
    n2802_lo <= 1'b0;
    n2805_lo <= 1'b0;
    n2808_lo <= 1'b0;
    n2820_lo <= 1'b0;
    n2823_lo <= 1'b0;
    n2826_lo <= 1'b0;
    n2829_lo <= 1'b0;
    n2832_lo <= 1'b0;
    n2835_lo <= 1'b0;
    n2838_lo <= 1'b0;
    n2841_lo <= 1'b0;
    n2844_lo <= 1'b0;
    n2856_lo <= 1'b0;
    n2859_lo <= 1'b0;
    n2862_lo <= 1'b0;
    n2865_lo <= 1'b0;
    n2868_lo <= 1'b0;
    n2871_lo <= 1'b0;
    n2874_lo <= 1'b0;
    n2877_lo <= 1'b0;
    n2880_lo <= 1'b0;
    n2883_lo <= 1'b0;
    n2886_lo <= 1'b0;
    n2889_lo <= 1'b0;
    n2892_lo <= 1'b0;
    n2895_lo <= 1'b0;
    n2898_lo <= 1'b0;
    n2901_lo <= 1'b0;
    n2904_lo <= 1'b0;
    n2907_lo <= 1'b0;
    n2916_lo <= 1'b0;
    n2919_lo <= 1'b0;
    n2925_lo <= 1'b0;
    n2928_lo <= 1'b0;
    n2940_lo <= 1'b0;
    n2943_lo <= 1'b0;
    n2952_lo <= 1'b0;
    n2955_lo <= 1'b0;
    n2961_lo <= 1'b0;
    n2964_lo <= 1'b0;
    n2967_lo <= 1'b0;
    n2970_lo <= 1'b0;
    n2976_lo <= 1'b0;
    n2979_lo <= 1'b0;
    n2982_lo <= 1'b0;
    n2988_lo <= 1'b0;
    n2991_lo <= 1'b0;
    n2994_lo <= 1'b0;
    n2997_lo <= 1'b0;
    n3000_lo <= 1'b0;
    n3003_lo <= 1'b0;
    n3006_lo <= 1'b0;
    n3012_lo <= 1'b0;
    n3015_lo <= 1'b0;
    n3018_lo <= 1'b0;
    n3021_lo <= 1'b0;
    n3024_lo <= 1'b0;
    n3027_lo <= 1'b0;
    n3030_lo <= 1'b0;
    n3033_lo <= 1'b0;
    n3036_lo <= 1'b0;
    n3039_lo <= 1'b0;
    n3045_lo <= 1'b0;
    n3048_lo <= 1'b0;
    n3051_lo <= 1'b0;
    n3054_lo <= 1'b0;
    n3057_lo <= 1'b0;
    n3060_lo <= 1'b0;
    n3063_lo <= 1'b0;
    n3069_lo <= 1'b0;
    n3072_lo <= 1'b0;
    n3075_lo <= 1'b0;
    n3081_lo <= 1'b0;
    n3084_lo <= 1'b0;
    n3087_lo <= 1'b0;
    n3093_lo <= 1'b0;
    n3096_lo <= 1'b0;
    n3099_lo <= 1'b0;
    n3102_lo <= 1'b0;
    n3105_lo <= 1'b0;
    n3108_lo <= 1'b0;
    n3111_lo <= 1'b0;
    n3114_lo <= 1'b0;
    n3117_lo <= 1'b0;
    n3120_lo <= 1'b0;
    n3123_lo <= 1'b0;
    n3126_lo <= 1'b0;
    n3129_lo <= 1'b0;
    n3132_lo <= 1'b0;
    n3135_lo <= 1'b0;
    n3138_lo <= 1'b0;
    n3141_lo <= 1'b0;
    n3156_lo <= 1'b0;
    n3168_lo <= 1'b0;
    n3171_lo <= 1'b0;
    n3174_lo <= 1'b0;
    n3177_lo <= 1'b0;
    n3180_lo <= 1'b0;
    n3183_lo <= 1'b0;
    n3192_lo <= 1'b0;
    n3195_lo <= 1'b0;
    n3204_lo <= 1'b0;
    n3207_lo <= 1'b0;
    n3210_lo <= 1'b0;
    n3216_lo <= 1'b0;
    n3219_lo <= 1'b0;
    n3222_lo <= 1'b0;
    n3228_lo <= 1'b0;
    n3231_lo <= 1'b0;
    n3240_lo <= 1'b0;
    n3243_lo <= 1'b0;
    n3252_lo <= 1'b0;
    n3255_lo <= 1'b0;
    n3258_lo <= 1'b0;
    n3264_lo <= 1'b0;
    n3267_lo <= 1'b0;
    n3270_lo <= 1'b0;
    n3276_lo <= 1'b0;
    n3279_lo <= 1'b0;
    n3282_lo <= 1'b0;
    n3288_lo <= 1'b0;
    n3291_lo <= 1'b0;
    n3294_lo <= 1'b0;
    n3603_o2 <= 1'b0;
    n3604_o2 <= 1'b0;
    n1391_inv <= 1'b0;
    n3798_o2 <= 1'b0;
    n3846_o2 <= 1'b0;
    n4019_o2 <= 1'b0;
    n4017_o2 <= 1'b0;
    n2177_o2 <= 1'b0;
    n2150_o2 <= 1'b0;
    n2154_o2 <= 1'b0;
    n2184_o2 <= 1'b0;
    n2515_o2 <= 1'b0;
    n3837_o2 <= 1'b0;
    n2167_o2 <= 1'b0;
    n2118_o2 <= 1'b0;
    n2186_o2 <= 1'b0;
    n2174_o2 <= 1'b0;
    n3964_o2 <= 1'b0;
    n4005_o2 <= 1'b0;
    n4006_o2 <= 1'b0;
    n1445_inv <= 1'b0;
    n2176_o2 <= 1'b0;
    n2227_o2 <= 1'b0;
    n2236_o2 <= 1'b0;
    n2245_o2 <= 1'b0;
    n2518_o2 <= 1'b0;
    n4023_o2 <= 1'b0;
    n1466_inv <= 1'b0;
    n4038_o2 <= 1'b0;
    n4039_o2 <= 1'b0;
    n1475_inv <= 1'b0;
    n2119_o2 <= 1'b0;
    n2275_o2 <= 1'b0;
    n2595_o2 <= 1'b0;
    n2594_o2 <= 1'b0;
    lo498_buf_o2 <= 1'b0;
    lo502_buf_o2 <= 1'b0;
    lo550_buf_o2 <= 1'b0;
    n2596_o2 <= 1'b0;
    n2593_o2 <= 1'b0;
    n2668_o2 <= 1'b0;
    lo542_buf_o2 <= 1'b0;
    n2667_o2 <= 1'b0;
    n2404_o2 <= 1'b0;
    n2410_o2 <= 1'b0;
    n2419_o2 <= 1'b0;
    n2392_o2 <= 1'b0;
    n2369_o2 <= 1'b0;
    n2397_o2 <= 1'b0;
    n2601_o2 <= 1'b0;
    n2658_o2 <= 1'b0;
    n2574_o2 <= 1'b0;
    n2205_o2 <= 1'b0;
    lo510_buf_o2 <= 1'b0;
    lo514_buf_o2 <= 1'b0;
    lo554_buf_o2 <= 1'b0;
    lo558_buf_o2 <= 1'b0;
    lo578_buf_o2 <= 1'b0;
    n2254_o2 <= 1'b0;
    n2421_o2 <= 1'b0;
    n2422_o2 <= 1'b0;
    n2130_o2 <= 1'b0;
    n2127_o2 <= 1'b0;
    n2131_o2 <= 1'b0;
    n2128_o2 <= 1'b0;
    n2264_o2 <= 1'b0;
    n2467_o2 <= 1'b0;
    n2471_o2 <= 1'b0;
    n2488_o2 <= 1'b0;
    n2478_o2 <= 1'b0;
    n2486_o2 <= 1'b0;
    n2485_o2 <= 1'b0;
    n2498_o2 <= 1'b0;
    n2495_o2 <= 1'b0;
    n2496_o2 <= 1'b0;
    n2458_o2 <= 1'b0;
    n2643_o2 <= 1'b0;
    n2462_o2 <= 1'b0;
    n2468_o2 <= 1'b0;
    n2639_o2 <= 1'b0;
    n2499_o2 <= 1'b0;
    n2472_o2 <= 1'b0;
    n2474_o2 <= 1'b0;
    n2489_o2 <= 1'b0;
    n2321_o2 <= 1'b0;
    n2322_o2 <= 1'b0;
    n2640_o2 <= 1'b0;
    n2642_o2 <= 1'b0;
    n2187_o2 <= 1'b0;
    n2373_o2 <= 1'b0;
    n2603_o2 <= 1'b0;
    n2388_o2 <= 1'b0;
    n2437_o2 <= 1'b0;
    n2356_o2 <= 1'b0;
    n2452_o2 <= 1'b0;
    n2347_o2 <= 1'b0;
    n2329_o2 <= 1'b0;
    n2669_o2 <= 1'b0;
    n2332_o2 <= 1'b0;
    n2664_o2 <= 1'b0;
    n2665_o2 <= 1'b0;
    n2653_o2 <= 1'b0;
    n2654_o2 <= 1'b0;
    n2636_o2 <= 1'b0;
    n2660_o2 <= 1'b0;
    n2318_o2 <= 1'b0;
    n2319_o2 <= 1'b0;
    n2586_o2 <= 1'b0;
    n2587_o2 <= 1'b0;
    n2288_o2 <= 1'b0;
    n2344_o2 <= 1'b0;
    n2530_o2 <= 1'b0;
    n2303_o2 <= 1'b0;
    n2566_o2 <= 1'b0;
    n2567_o2 <= 1'b0;
    n2554_o2 <= 1'b0;
    n2194_o2 <= 1'b0;
    lo582_buf_o2 <= 1'b0;
    lo030_buf_o2 <= 1'b0;
    lo174_buf_o2 <= 1'b0;
    lo178_buf_o2 <= 1'b0;
    lo186_buf_o2 <= 1'b0;
    lo266_buf_o2 <= 1'b0;
    lo306_buf_o2 <= 1'b0;
    lo346_buf_o2 <= 1'b0;
    lo386_buf_o2 <= 1'b0;
    lo426_buf_o2 <= 1'b0;
    lo590_buf_o2 <= 1'b0;
    lo594_buf_o2 <= 1'b0;
    lo606_buf_o2 <= 1'b0;
    lo610_buf_o2 <= 1'b0;
    n2238_o2 <= 1'b0;
    n2229_o2 <= 1'b0;
    n2242_o2 <= 1'b0;
    n2233_o2 <= 1'b0;
    n2168_o2 <= 1'b0;
    n2237_o2 <= 1'b0;
    n2228_o2 <= 1'b0;
    n2172_o2 <= 1'b0;
    n2223_o2 <= 1'b0;
    n2222_o2 <= 1'b0;
    n2170_o2 <= 1'b0;
    n2181_o2 <= 1'b0;
    n2510_o2 <= 1'b0;
    n2621_o2 <= 1'b0;
    lo466_buf_o2 <= 1'b0;
    lo478_buf_o2 <= 1'b0;
    n2149_o2 <= 1'b0;
    n2429_o2 <= 1'b0;
    n2444_o2 <= 1'b0;
    n2153_o2 <= 1'b0;
    n2433_o2 <= 1'b0;
    n2448_o2 <= 1'b0;
    n2367_o2 <= 1'b0;
    n2386_o2 <= 1'b0;
    n2539_o2 <= 1'b0;
    n2183_o2 <= 1'b0;
    n2220_o2 <= 1'b0;
    n2514_o2 <= 1'b0;
    n2196_o2 <= 1'b0;
    n2616_o2 <= 1'b0;
    n2612_o2 <= 1'b0;
    n2627_o2 <= 1'b0;
    n2140_o2 <= 1'b0;
    n1877_inv <= 1'b0;
    lo149_buf_o2 <= 1'b0;
    lo197_buf_o2 <= 1'b0;
    lo118_buf_o2 <= 1'b0;
    lo158_buf_o2 <= 1'b0;
    lo166_buf_o2 <= 1'b0;
    lo242_buf_o2 <= 1'b0;
    lo286_buf_o2 <= 1'b0;
    lo506_buf_o2 <= 1'b0;
    n2198_o2 <= 1'b0;
    n2202_o2 <= 1'b0;
    n2197_o2 <= 1'b0;
    n1913_inv <= 1'b0;
    n2146_o2 <= 1'b0;
    n1919_inv <= 1'b0;
    lo312_buf_o2 <= 1'b0;
    lo316_buf_o2 <= 1'b0;
    lo352_buf_o2 <= 1'b0;
    lo356_buf_o2 <= 1'b0;
    lo392_buf_o2 <= 1'b0;
    lo396_buf_o2 <= 1'b0;
    lo432_buf_o2 <= 1'b0;
    lo436_buf_o2 <= 1'b0;
    lo576_buf_o2 <= 1'b0;
  end
endmodule


