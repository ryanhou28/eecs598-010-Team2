
module mymod
(
  G1_p,
  G1_n,
  G2_p,
  G2_n,
  G3_p,
  G3_n,
  G4_p,
  G4_n,
  G5_p,
  G5_n,
  G6_p,
  G6_n,
  G7_p,
  G7_n,
  G8_p,
  G8_n,
  G9_p,
  G9_n,
  G10_p,
  G10_n,
  G11_p,
  G11_n,
  G12_p,
  G12_n,
  G13_p,
  G13_n,
  G14_p,
  G14_n,
  G15_p,
  G15_n,
  G16_p,
  G16_n,
  G17_p,
  G17_n,
  G18_p,
  G18_n,
  G19_p,
  G19_n,
  G20_p,
  G20_n,
  G21_p,
  G21_n,
  G22_p,
  G22_n,
  G23_p,
  G23_n,
  G24_p,
  G24_n,
  G25_p,
  G25_n,
  G26_p,
  G26_n,
  G27_p,
  G27_n,
  G28_p,
  G28_n,
  G29_p,
  G29_n,
  G30_p,
  G30_n,
  G31_p,
  G31_n,
  G32_p,
  G32_n,
  G33_p,
  G33_n,
  G1884_p,
  G1885_p,
  G1886_p,
  G1887_p,
  G1888_p,
  G1889_p,
  G1890_p,
  G1891_p,
  G1892_p,
  G1893_p,
  G1894_p,
  G1895_p,
  G1896_p,
  G1897_p,
  G1898_p,
  G1899_p,
  G1900_p,
  G1901_p,
  G1902_p,
  G1903_p,
  G1904_p,
  G1905_p,
  G1906_p,
  G1907_p,
  G1908_p
);

  input G1_p;input G1_n;input G2_p;input G2_n;input G3_p;input G3_n;input G4_p;input G4_n;input G5_p;input G5_n;input G6_p;input G6_n;input G7_p;input G7_n;input G8_p;input G8_n;input G9_p;input G9_n;input G10_p;input G10_n;input G11_p;input G11_n;input G12_p;input G12_n;input G13_p;input G13_n;input G14_p;input G14_n;input G15_p;input G15_n;input G16_p;input G16_n;input G17_p;input G17_n;input G18_p;input G18_n;input G19_p;input G19_n;input G20_p;input G20_n;input G21_p;input G21_n;input G22_p;input G22_n;input G23_p;input G23_n;input G24_p;input G24_n;input G25_p;input G25_n;input G26_p;input G26_n;input G27_p;input G27_n;input G28_p;input G28_n;input G29_p;input G29_n;input G30_p;input G30_n;input G31_p;input G31_n;input G32_p;input G32_n;input G33_p;input G33_n;
  output G1884_p;output G1885_p;output G1886_p;output G1887_p;output G1888_p;output G1889_p;output G1890_p;output G1891_p;output G1892_p;output G1893_p;output G1894_p;output G1895_p;output G1896_p;output G1897_p;output G1898_p;output G1899_p;output G1900_p;output G1901_p;output G1902_p;output G1903_p;output G1904_p;output G1905_p;output G1906_p;output G1907_p;output G1908_p;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire ffc_0_p;
  wire ffc_0_n;
  wire ffc_1_p;
  wire ffc_1_n;
  wire ffc_2_p;
  wire ffc_2_n;
  wire ffc_3_p;
  wire ffc_3_n;
  wire ffc_4_p;
  wire ffc_4_n;
  wire ffc_5_p;
  wire ffc_5_n;
  wire ffc_6_p;
  wire ffc_6_n;
  wire ffc_7_p;
  wire ffc_7_n;
  wire ffc_8_p;
  wire ffc_8_n;
  wire ffc_9_p;
  wire ffc_9_n;
  wire ffc_10_p;
  wire ffc_10_n;
  wire ffc_11_p;
  wire ffc_11_n;
  wire ffc_12_p;
  wire ffc_12_n;
  wire ffc_13_p;
  wire ffc_13_n;
  wire ffc_14_p;
  wire ffc_14_n;
  wire ffc_15_p;
  wire ffc_15_n;
  wire ffc_16_p;
  wire ffc_16_n;
  wire ffc_17_p;
  wire ffc_17_n;
  wire ffc_18_p;
  wire ffc_18_n;
  wire ffc_19_p;
  wire ffc_19_n;
  wire ffc_20_p;
  wire ffc_20_n;
  wire ffc_21_p;
  wire ffc_21_n;
  wire ffc_22_p;
  wire ffc_22_n;
  wire ffc_23_p;
  wire ffc_23_n;
  wire ffc_24_p;
  wire ffc_24_n;
  wire ffc_25_p;
  wire ffc_25_n;
  wire ffc_26_p;
  wire ffc_26_n;
  wire ffc_27_p;
  wire ffc_27_n;
  wire ffc_28_p;
  wire ffc_28_n;
  wire ffc_29_p;
  wire ffc_29_n;
  wire ffc_30_p;
  wire ffc_30_n;
  wire ffc_31_p;
  wire ffc_31_n;
  wire ffc_32_p;
  wire ffc_32_n;
  wire ffc_33_p;
  wire ffc_33_n;
  wire ffc_34_p;
  wire ffc_34_n;
  wire ffc_35_p;
  wire ffc_35_n;
  wire ffc_36_p;
  wire ffc_36_n;
  wire ffc_37_p;
  wire ffc_37_n;
  wire ffc_38_p;
  wire ffc_38_n;
  wire ffc_39_p;
  wire ffc_39_n;
  wire ffc_40_p;
  wire ffc_40_n;
  wire ffc_41_p;
  wire ffc_41_n;
  wire ffc_42_p;
  wire ffc_42_n;
  wire ffc_43_p;
  wire ffc_43_n;
  wire ffc_44_p;
  wire ffc_44_n;
  wire ffc_45_p;
  wire ffc_45_n;
  wire ffc_46_p;
  wire ffc_46_n;
  wire ffc_47_p;
  wire ffc_47_n;
  wire ffc_48_p;
  wire ffc_48_n;
  wire ffc_49_p;
  wire ffc_49_n;
  wire ffc_50_p;
  wire ffc_50_n;
  wire ffc_51_p;
  wire ffc_51_n;
  wire ffc_52_p;
  wire ffc_52_n;
  wire ffc_53_p;
  wire ffc_53_n;
  wire ffc_54_p;
  wire ffc_54_n;
  wire ffc_55_p;
  wire ffc_55_n;
  wire ffc_56_p;
  wire ffc_56_n;
  wire ffc_57_p;
  wire ffc_57_n;
  wire ffc_58_p;
  wire ffc_58_n;
  wire ffc_59_p;
  wire ffc_59_n;
  wire ffc_60_p;
  wire ffc_60_n;
  wire ffc_61_p;
  wire ffc_61_n;
  wire ffc_62_p;
  wire ffc_62_n;
  wire ffc_63_p;
  wire ffc_63_n;
  wire ffc_64_p;
  wire ffc_64_n;
  wire ffc_65_p;
  wire ffc_65_n;
  wire ffc_66_p;
  wire ffc_66_n;
  wire ffc_67_p;
  wire ffc_67_n;
  wire ffc_68_p;
  wire ffc_68_n;
  wire ffc_69_p;
  wire ffc_69_n;
  wire ffc_70_p;
  wire ffc_70_n;
  wire ffc_71_p;
  wire ffc_71_n;
  wire ffc_72_p;
  wire ffc_72_n;
  wire ffc_73_p;
  wire ffc_73_n;
  wire ffc_74_p;
  wire ffc_74_n;
  wire ffc_75_p;
  wire ffc_75_n;
  wire ffc_76_p;
  wire ffc_76_n;
  wire ffc_77_p;
  wire ffc_77_n;
  wire ffc_78_p;
  wire ffc_78_n;
  wire ffc_79_p;
  wire ffc_79_n;
  wire ffc_80_p;
  wire ffc_80_n;
  wire ffc_81_p;
  wire ffc_81_n;
  wire ffc_82_p;
  wire ffc_82_n;
  wire ffc_83_p;
  wire ffc_83_n;
  wire ffc_84_p;
  wire ffc_84_n;
  wire ffc_85_p;
  wire ffc_85_n;
  wire ffc_86_p;
  wire ffc_86_n;
  wire ffc_87_p;
  wire ffc_87_n;
  wire ffc_88_p;
  wire ffc_88_n;
  wire ffc_89_p;
  wire ffc_89_n;
  wire ffc_90_p;
  wire ffc_90_n;
  wire ffc_91_p;
  wire ffc_91_n;
  wire ffc_92_p;
  wire ffc_92_n;
  wire ffc_93_p;
  wire ffc_93_n;
  wire ffc_94_p;
  wire ffc_94_n;
  wire ffc_95_p;
  wire ffc_95_n;
  wire ffc_96_p;
  wire ffc_96_n;
  wire ffc_97_p;
  wire ffc_97_n;
  wire ffc_98_p;
  wire ffc_98_n;
  wire ffc_99_p;
  wire ffc_99_n;
  wire ffc_100_p;
  wire ffc_100_n;
  wire ffc_101_p;
  wire ffc_101_n;
  wire ffc_102_p;
  wire ffc_102_n;
  wire ffc_103_p;
  wire ffc_103_n;
  wire ffc_104_p;
  wire ffc_104_n;
  wire ffc_105_p;
  wire ffc_105_n;
  wire ffc_106_p;
  wire ffc_106_n;
  wire ffc_107_p;
  wire ffc_107_n;
  wire ffc_108_p;
  wire ffc_108_n;
  wire ffc_109_p;
  wire ffc_109_n;
  wire ffc_110_p;
  wire ffc_110_n;
  wire ffc_111_p;
  wire ffc_111_n;
  wire ffc_112_p;
  wire ffc_112_n;
  wire ffc_113_p;
  wire ffc_113_n;
  wire ffc_114_p;
  wire ffc_114_n;
  wire ffc_115_p;
  wire ffc_115_n;
  wire ffc_116_p;
  wire ffc_116_n;
  wire ffc_117_p;
  wire ffc_117_n;
  wire ffc_118_p;
  wire ffc_118_n;
  wire ffc_119_p;
  wire ffc_119_n;
  wire ffc_120_p;
  wire ffc_120_n;
  wire ffc_121_p;
  wire ffc_121_n;
  wire ffc_122_p;
  wire ffc_122_n;
  wire ffc_123_p;
  wire ffc_123_n;
  wire ffc_124_p;
  wire ffc_124_n;
  wire ffc_125_p;
  wire ffc_125_n;
  wire ffc_126_p;
  wire ffc_126_n;
  wire ffc_127_p;
  wire ffc_127_n;
  wire ffc_128_p;
  wire ffc_128_n;
  wire ffc_129_p;
  wire ffc_129_n;
  wire ffc_130_p;
  wire ffc_130_n;
  wire ffc_131_p;
  wire ffc_131_n;
  wire ffc_132_p;
  wire ffc_132_n;
  wire ffc_133_p;
  wire ffc_133_n;
  wire ffc_134_p;
  wire ffc_134_n;
  wire ffc_135_p;
  wire ffc_135_n;
  wire ffc_136_p;
  wire ffc_136_n;
  wire ffc_137_p;
  wire ffc_137_n;
  wire ffc_138_p;
  wire ffc_138_n;
  wire ffc_139_p;
  wire ffc_139_n;
  wire ffc_140_p;
  wire ffc_140_n;
  wire ffc_141_p;
  wire ffc_141_n;
  wire ffc_142_p;
  wire ffc_142_n;
  wire ffc_143_p;
  wire ffc_143_n;
  wire ffc_144_p;
  wire ffc_144_n;
  wire ffc_145_p;
  wire ffc_145_n;
  wire ffc_146_p;
  wire ffc_146_n;
  wire ffc_147_p;
  wire ffc_147_n;
  wire ffc_148_p;
  wire ffc_148_n;
  wire ffc_149_p;
  wire ffc_149_n;
  wire ffc_150_p;
  wire ffc_150_n;
  wire ffc_151_p;
  wire ffc_151_n;
  wire ffc_152_p;
  wire ffc_152_n;
  wire ffc_153_p;
  wire ffc_153_n;
  wire ffc_154_p;
  wire ffc_154_n;
  wire ffc_155_p;
  wire ffc_155_n;
  wire ffc_156_p;
  wire ffc_156_n;
  wire ffc_157_p;
  wire ffc_157_n;
  wire ffc_158_p;
  wire ffc_158_n;
  wire ffc_159_p;
  wire ffc_159_n;
  wire ffc_160_p;
  wire ffc_160_n;
  wire ffc_161_p;
  wire ffc_161_n;
  wire ffc_162_p;
  wire ffc_162_n;
  wire ffc_163_p;
  wire ffc_163_n;
  wire ffc_164_p;
  wire ffc_164_n;
  wire ffc_165_p;
  wire ffc_165_n;
  wire ffc_166_p;
  wire ffc_166_n;
  wire ffc_167_p;
  wire ffc_167_n;
  wire ffc_168_p;
  wire ffc_168_n;
  wire ffc_169_p;
  wire ffc_169_n;
  wire ffc_170_p;
  wire ffc_170_n;
  wire ffc_171_p;
  wire ffc_171_n;
  wire ffc_172_p;
  wire ffc_172_n;
  wire ffc_173_p;
  wire ffc_173_n;
  wire ffc_174_p;
  wire ffc_174_n;
  wire ffc_175_p;
  wire ffc_175_n;
  wire ffc_176_p;
  wire ffc_176_n;
  wire ffc_177_p;
  wire ffc_177_n;
  wire ffc_178_p;
  wire ffc_178_n;
  wire ffc_179_p;
  wire ffc_179_n;
  wire ffc_180_p;
  wire ffc_180_n;
  wire ffc_181_p;
  wire ffc_181_n;
  wire ffc_182_p;
  wire ffc_182_n;
  wire ffc_183_p;
  wire ffc_183_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire ffc_129_n_spl_;
  wire ffc_131_p_spl_;
  wire ffc_129_p_spl_;
  wire ffc_131_n_spl_;
  wire g218_n_spl_;
  wire g218_n_spl_0;
  wire g218_n_spl_00;
  wire g218_n_spl_01;
  wire g218_n_spl_1;
  wire g218_n_spl_10;
  wire g218_p_spl_;
  wire g218_p_spl_0;
  wire g218_p_spl_00;
  wire g218_p_spl_01;
  wire g218_p_spl_1;
  wire g218_p_spl_10;
  wire ffc_130_n_spl_;
  wire ffc_130_n_spl_0;
  wire ffc_130_p_spl_;
  wire ffc_130_p_spl_0;
  wire g231_n_spl_;
  wire g231_n_spl_0;
  wire g231_n_spl_00;
  wire g231_n_spl_01;
  wire g231_n_spl_1;
  wire g231_p_spl_;
  wire g231_p_spl_0;
  wire g231_p_spl_00;
  wire g231_p_spl_01;
  wire g231_p_spl_1;
  wire ffc_98_n_spl_;
  wire ffc_93_n_spl_;
  wire g242_p_spl_;
  wire g242_n_spl_;
  wire g243_n_spl_;
  wire g243_n_spl_0;
  wire g243_n_spl_1;
  wire g243_p_spl_;
  wire g243_p_spl_0;
  wire g243_p_spl_1;
  wire ffc_91_n_spl_;
  wire ffc_92_p_spl_;
  wire ffc_99_p_spl_;
  wire g263_n_spl_;
  wire g263_n_spl_0;
  wire g263_n_spl_1;
  wire g263_p_spl_;
  wire g263_p_spl_0;
  wire g263_p_spl_1;
  wire g276_n_spl_;
  wire g276_n_spl_0;
  wire g276_n_spl_00;
  wire g276_n_spl_01;
  wire g276_n_spl_1;
  wire ffc_58_p_spl_;
  wire ffc_58_p_spl_0;
  wire ffc_53_n_spl_;
  wire ffc_53_n_spl_0;
  wire ffc_53_n_spl_00;
  wire ffc_53_n_spl_1;
  wire ffc_53_p_spl_;
  wire ffc_53_p_spl_0;
  wire g276_p_spl_;
  wire g276_p_spl_0;
  wire ffc_97_p_spl_;
  wire ffc_97_p_spl_0;
  wire ffc_97_p_spl_00;
  wire ffc_97_p_spl_01;
  wire ffc_97_p_spl_1;
  wire ffc_58_n_spl_;
  wire g310_n_spl_;
  wire g310_p_spl_;
  wire g320_n_spl_;
  wire g320_p_spl_;
  wire ffc_142_n_spl_;
  wire ffc_102_n_spl_;
  wire ffc_102_p_spl_;
  wire ffc_102_p_spl_0;
  wire ffc_102_p_spl_1;
  wire ffc_152_p_spl_;
  wire g331_p_spl_;
  wire ffc_45_p_spl_;
  wire ffc_81_p_spl_;
  wire ffc_81_p_spl_0;
  wire ffc_81_p_spl_1;
  wire ffc_49_p_spl_;
  wire ffc_56_p_spl_;
  wire g332_n_spl_;
  wire ffc_32_p_spl_;
  wire ffc_141_p_spl_;
  wire ffc_140_p_spl_;
  wire g338_n_spl_;
  wire g345_p_spl_;
  wire g333_n_spl_;
  wire g337_p_spl_;
  wire g356_p_spl_;
  wire ffc_52_p_spl_;
  wire ffc_52_p_spl_0;
  wire ffc_52_p_spl_1;
  wire ffc_138_p_spl_;
  wire ffc_138_p_spl_0;
  wire ffc_162_n_spl_;
  wire ffc_163_p_spl_;
  wire ffc_162_p_spl_;
  wire ffc_163_n_spl_;
  wire ffc_161_p_spl_;
  wire ffc_119_n_spl_;
  wire ffc_119_n_spl_0;
  wire ffc_119_n_spl_1;
  wire ffc_119_p_spl_;
  wire ffc_119_p_spl_0;
  wire ffc_119_p_spl_00;
  wire ffc_119_p_spl_1;
  wire ffc_164_n_spl_;
  wire ffc_164_n_spl_0;
  wire ffc_164_n_spl_1;
  wire ffc_166_p_spl_;
  wire ffc_164_p_spl_;
  wire ffc_164_p_spl_0;
  wire ffc_164_p_spl_1;
  wire ffc_166_n_spl_;
  wire ffc_107_n_spl_;
  wire ffc_158_p_spl_;
  wire ffc_107_p_spl_;
  wire ffc_107_p_spl_0;
  wire ffc_158_n_spl_;
  wire ffc_165_p_spl_;
  wire ffc_165_p_spl_0;
  wire ffc_167_p_spl_;
  wire ffc_167_p_spl_0;
  wire ffc_167_p_spl_1;
  wire ffc_165_n_spl_;
  wire ffc_165_n_spl_0;
  wire ffc_167_n_spl_;
  wire ffc_167_n_spl_0;
  wire ffc_167_n_spl_1;
  wire ffc_116_n_spl_;
  wire ffc_135_p_spl_;
  wire ffc_135_p_spl_0;
  wire ffc_135_p_spl_00;
  wire ffc_135_p_spl_1;
  wire ffc_116_p_spl_;
  wire ffc_116_p_spl_0;
  wire ffc_135_n_spl_;
  wire ffc_135_n_spl_0;
  wire ffc_135_n_spl_1;
  wire g381_n_spl_;
  wire g384_p_spl_;
  wire g381_p_spl_;
  wire g384_n_spl_;
  wire g361_n_spl_;
  wire g391_p_spl_;
  wire g339_n_spl_;
  wire g392_n_spl_;
  wire g341_n_spl_;
  wire g394_n_spl_;
  wire g340_n_spl_;
  wire g358_n_spl_;
  wire g360_p_spl_;
  wire g399_p_spl_;
  wire g399_n_spl_;
  wire ffc_112_n_spl_;
  wire g403_n_spl_;
  wire ffc_112_p_spl_;
  wire ffc_112_p_spl_0;
  wire g403_p_spl_;
  wire ffc_134_p_spl_;
  wire ffc_134_p_spl_0;
  wire g410_p_spl_;
  wire ffc_134_n_spl_;
  wire g410_n_spl_;
  wire g357_p_spl_;
  wire g357_p_spl_0;
  wire g357_n_spl_;
  wire g357_n_spl_0;
  wire g357_n_spl_1;
  wire ffc_175_n_spl_;
  wire ffc_176_n_spl_;
  wire ffc_175_p_spl_;
  wire ffc_175_p_spl_0;
  wire ffc_176_p_spl_;
  wire ffc_176_p_spl_0;
  wire ffc_110_p_spl_;
  wire ffc_52_n_spl_;
  wire ffc_52_n_spl_0;
  wire g409_n_spl_;
  wire g419_n_spl_;
  wire g369_n_spl_;
  wire ffc_41_n_spl_;
  wire g426_p_spl_;
  wire g378_p_spl_;
  wire g390_p_spl_;
  wire g390_p_spl_0;
  wire g429_n_spl_;
  wire ffc_27_p_spl_;
  wire ffc_118_n_spl_;
  wire ffc_118_p_spl_;
  wire ffc_118_p_spl_0;
  wire g438_n_spl_;
  wire g441_p_spl_;
  wire ffc_154_p_spl_;
  wire ffc_117_p_spl_;
  wire ffc_117_p_spl_0;
  wire ffc_153_n_spl_;
  wire ffc_117_n_spl_;
  wire ffc_153_p_spl_;
  wire g444_p_spl_;
  wire g447_n_spl_;
  wire g444_n_spl_;
  wire g447_p_spl_;
  wire g387_p_spl_;
  wire ffc_178_p_spl_;
  wire ffc_178_p_spl_0;
  wire ffc_178_p_spl_00;
  wire ffc_178_p_spl_1;
  wire ffc_181_n_spl_;
  wire ffc_181_n_spl_0;
  wire ffc_178_n_spl_;
  wire ffc_178_n_spl_0;
  wire ffc_178_n_spl_1;
  wire ffc_181_p_spl_;
  wire ffc_181_p_spl_0;
  wire ffc_181_p_spl_1;
  wire ffc_19_p_spl_;
  wire ffc_19_p_spl_0;
  wire g456_n_spl_;
  wire ffc_19_n_spl_;
  wire g456_p_spl_;
  wire ffc_21_p_spl_;
  wire ffc_183_n_spl_;
  wire ffc_6_p_spl_;
  wire ffc_6_p_spl_0;
  wire ffc_174_n_spl_;
  wire ffc_174_n_spl_0;
  wire ffc_6_n_spl_;
  wire ffc_174_p_spl_;
  wire ffc_174_p_spl_0;
  wire ffc_174_p_spl_1;
  wire ffc_23_p_spl_;
  wire ffc_177_n_spl_;
  wire ffc_182_p_spl_;
  wire ffc_183_p_spl_;
  wire ffc_177_p_spl_;
  wire ffc_13_n_spl_;
  wire ffc_13_n_spl_0;
  wire g469_n_spl_;
  wire ffc_179_n_spl_;
  wire ffc_179_n_spl_0;
  wire ffc_179_p_spl_;
  wire ffc_179_p_spl_0;
  wire ffc_179_p_spl_1;
  wire ffc_172_p_spl_;
  wire ffc_172_p_spl_0;
  wire ffc_172_p_spl_00;
  wire ffc_172_p_spl_1;
  wire ffc_172_n_spl_;
  wire ffc_172_n_spl_0;
  wire ffc_172_n_spl_1;
  wire ffc_171_n_spl_;
  wire ffc_171_n_spl_0;
  wire ffc_171_p_spl_;
  wire ffc_171_p_spl_0;
  wire ffc_171_p_spl_1;
  wire g422_p_spl_;
  wire ffc_170_n_spl_;
  wire ffc_170_p_spl_;
  wire ffc_170_p_spl_0;
  wire ffc_0_p_spl_;
  wire ffc_173_p_spl_;
  wire ffc_173_p_spl_0;
  wire ffc_173_p_spl_00;
  wire ffc_173_p_spl_1;
  wire ffc_173_n_spl_;
  wire ffc_173_n_spl_0;
  wire ffc_173_n_spl_1;
  wire ffc_4_p_spl_;
  wire ffc_180_n_spl_;
  wire ffc_180_p_spl_;
  wire ffc_180_p_spl_0;
  wire ffc_13_p_spl_;
  wire g459_n_spl_;
  wire g459_n_spl_0;
  wire g507_n_spl_;

  andX
  g_g218_p
  (
    .dout(g218_p),
    .din1(ffc_129_n_spl_),
    .din2(ffc_131_p_spl_)
  );


  orX
  g_g218_n
  (
    .dout(g218_n),
    .din1(ffc_129_p_spl_),
    .din2(ffc_131_n_spl_)
  );


  andX
  g_g219_p
  (
    .dout(g219_p),
    .din1(ffc_1_n),
    .din2(g218_n_spl_00)
  );


  andX
  g_g220_p
  (
    .dout(g220_p),
    .din1(ffc_1_p),
    .din2(g218_p_spl_00)
  );


  orX
  g_g221_n
  (
    .dout(g221_n),
    .din1(g219_p),
    .din2(g220_p)
  );


  andX
  g_g222_p
  (
    .dout(g222_p),
    .din1(ffc_2_n),
    .din2(g218_n_spl_00)
  );


  andX
  g_g223_p
  (
    .dout(g223_p),
    .din1(ffc_2_p),
    .din2(g218_p_spl_00)
  );


  orX
  g_g224_n
  (
    .dout(g224_n),
    .din1(g222_p),
    .din2(g223_p)
  );


  andX
  g_g225_p
  (
    .dout(g225_p),
    .din1(ffc_3_n),
    .din2(g218_n_spl_01)
  );


  andX
  g_g226_p
  (
    .dout(g226_p),
    .din1(ffc_3_p),
    .din2(g218_p_spl_01)
  );


  orX
  g_g227_n
  (
    .dout(g227_n),
    .din1(g225_p),
    .din2(g226_p)
  );


  andX
  g_g228_p
  (
    .dout(g228_p),
    .din1(ffc_5_n),
    .din2(g218_n_spl_01)
  );


  andX
  g_g229_p
  (
    .dout(g229_p),
    .din1(ffc_5_p),
    .din2(g218_p_spl_01)
  );


  orX
  g_g230_n
  (
    .dout(g230_n),
    .din1(g228_p),
    .din2(g229_p)
  );


  andX
  g_g231_p
  (
    .dout(g231_p),
    .din1(ffc_130_n_spl_0),
    .din2(ffc_131_p_spl_)
  );


  orX
  g_g231_n
  (
    .dout(g231_n),
    .din1(ffc_130_p_spl_0),
    .din2(ffc_131_n_spl_)
  );


  andX
  g_g232_p
  (
    .dout(g232_p),
    .din1(ffc_12_n),
    .din2(g231_n_spl_00)
  );


  andX
  g_g233_p
  (
    .dout(g233_p),
    .din1(ffc_12_p),
    .din2(g231_p_spl_00)
  );


  orX
  g_g234_n
  (
    .dout(g234_n),
    .din1(g232_p),
    .din2(g233_p)
  );


  andX
  g_g235_p
  (
    .dout(g235_p),
    .din1(ffc_18_n),
    .din2(g231_n_spl_00)
  );


  andX
  g_g236_p
  (
    .dout(g236_p),
    .din1(ffc_18_p),
    .din2(g231_p_spl_00)
  );


  orX
  g_g237_n
  (
    .dout(g237_n),
    .din1(g235_p),
    .din2(g236_p)
  );


  andX
  g_g238_p
  (
    .dout(g238_p),
    .din1(ffc_20_n),
    .din2(g231_n_spl_01)
  );


  andX
  g_g239_p
  (
    .dout(g239_p),
    .din1(ffc_20_p),
    .din2(g231_p_spl_01)
  );


  orX
  g_g240_n
  (
    .dout(g240_n),
    .din1(g238_p),
    .din2(g239_p)
  );


  andX
  g_g241_p
  (
    .dout(g241_p),
    .din1(ffc_93_p),
    .din2(ffc_98_n_spl_)
  );


  orX
  g_g241_n
  (
    .dout(g241_n),
    .din1(ffc_93_n_spl_),
    .din2(ffc_98_p)
  );


  andX
  g_g242_p
  (
    .dout(g242_p),
    .din1(ffc_104_p),
    .din2(g241_p)
  );


  orX
  g_g242_n
  (
    .dout(g242_n),
    .din1(ffc_104_n),
    .din2(g241_n)
  );


  andX
  g_g243_p
  (
    .dout(g243_p),
    .din1(ffc_129_n_spl_),
    .din2(g242_p_spl_)
  );


  orX
  g_g243_n
  (
    .dout(g243_n),
    .din1(ffc_129_p_spl_),
    .din2(g242_n_spl_)
  );


  andX
  g_g244_p
  (
    .dout(g244_p),
    .din1(ffc_7_n),
    .din2(g243_n_spl_0)
  );


  andX
  g_g245_p
  (
    .dout(g245_p),
    .din1(ffc_7_p),
    .din2(g243_p_spl_0)
  );


  orX
  g_g246_n
  (
    .dout(g246_n),
    .din1(g244_p),
    .din2(g245_p)
  );


  andX
  g_g247_p
  (
    .dout(g247_p),
    .din1(ffc_8_n),
    .din2(g243_n_spl_0)
  );


  andX
  g_g248_p
  (
    .dout(g248_p),
    .din1(ffc_8_p),
    .din2(g243_p_spl_0)
  );


  orX
  g_g249_n
  (
    .dout(g249_n),
    .din1(g247_p),
    .din2(g248_p)
  );


  andX
  g_g250_p
  (
    .dout(g250_p),
    .din1(ffc_9_n),
    .din2(g243_n_spl_1)
  );


  andX
  g_g251_p
  (
    .dout(g251_p),
    .din1(ffc_9_p),
    .din2(g243_p_spl_1)
  );


  orX
  g_g252_n
  (
    .dout(g252_n),
    .din1(g250_p),
    .din2(g251_p)
  );


  andX
  g_g253_p
  (
    .dout(g253_p),
    .din1(ffc_10_n),
    .din2(g243_n_spl_1)
  );


  andX
  g_g254_p
  (
    .dout(g254_p),
    .din1(ffc_10_p),
    .din2(g243_p_spl_1)
  );


  orX
  g_g255_n
  (
    .dout(g255_n),
    .din1(g253_p),
    .din2(g254_p)
  );


  andX
  g_g256_p
  (
    .dout(g256_p),
    .din1(ffc_130_n_spl_0),
    .din2(g242_p_spl_)
  );


  orX
  g_g256_n
  (
    .dout(g256_n),
    .din1(ffc_130_p_spl_0),
    .din2(g242_n_spl_)
  );


  andX
  g_g257_p
  (
    .dout(g257_p),
    .din1(ffc_11_p),
    .din2(g256_p)
  );


  andX
  g_g258_p
  (
    .dout(g258_p),
    .din1(ffc_11_n),
    .din2(g256_n)
  );


  orX
  g_g259_n
  (
    .dout(g259_n),
    .din1(g257_p),
    .din2(g258_p)
  );


  andX
  g_g260_p
  (
    .dout(g260_p),
    .din1(ffc_91_p),
    .din2(ffc_130_n_spl_)
  );


  orX
  g_g260_n
  (
    .dout(g260_n),
    .din1(ffc_91_n_spl_),
    .din2(ffc_130_p_spl_)
  );


  andX
  g_g261_p
  (
    .dout(g261_p),
    .din1(ffc_92_p_spl_),
    .din2(g260_p)
  );


  orX
  g_g261_n
  (
    .dout(g261_n),
    .din1(ffc_92_n),
    .din2(g260_n)
  );


  andX
  g_g262_p
  (
    .dout(g262_p),
    .din1(ffc_103_n),
    .din2(g261_p)
  );


  orX
  g_g262_n
  (
    .dout(g262_n),
    .din1(ffc_103_p),
    .din2(g261_n)
  );


  andX
  g_g263_p
  (
    .dout(g263_p),
    .din1(ffc_99_p_spl_),
    .din2(g262_p)
  );


  orX
  g_g263_n
  (
    .dout(g263_n),
    .din1(ffc_99_n),
    .din2(g262_n)
  );


  andX
  g_g264_p
  (
    .dout(g264_p),
    .din1(ffc_14_n),
    .din2(g263_n_spl_0)
  );


  andX
  g_g265_p
  (
    .dout(g265_p),
    .din1(ffc_14_p),
    .din2(g263_p_spl_0)
  );


  orX
  g_g266_n
  (
    .dout(g266_n),
    .din1(g264_p),
    .din2(g265_p)
  );


  andX
  g_g267_p
  (
    .dout(g267_p),
    .din1(ffc_15_n),
    .din2(g263_n_spl_0)
  );


  andX
  g_g268_p
  (
    .dout(g268_p),
    .din1(ffc_15_p),
    .din2(g263_p_spl_0)
  );


  orX
  g_g269_n
  (
    .dout(g269_n),
    .din1(g267_p),
    .din2(g268_p)
  );


  andX
  g_g270_p
  (
    .dout(g270_p),
    .din1(ffc_16_n),
    .din2(g263_n_spl_1)
  );


  andX
  g_g271_p
  (
    .dout(g271_p),
    .din1(ffc_16_p),
    .din2(g263_p_spl_1)
  );


  orX
  g_g272_n
  (
    .dout(g272_n),
    .din1(g270_p),
    .din2(g271_p)
  );


  andX
  g_g273_p
  (
    .dout(g273_p),
    .din1(ffc_17_n),
    .din2(g263_n_spl_1)
  );


  andX
  g_g274_p
  (
    .dout(g274_p),
    .din1(ffc_17_p),
    .din2(g263_p_spl_1)
  );


  orX
  g_g275_n
  (
    .dout(g275_n),
    .din1(g273_p),
    .din2(g274_p)
  );


  andX
  g_g276_p
  (
    .dout(g276_p),
    .din1(g218_n_spl_10),
    .din2(g231_n_spl_01)
  );


  orX
  g_g276_n
  (
    .dout(g276_n),
    .din1(g218_p_spl_10),
    .din2(g231_p_spl_01)
  );


  andX
  g_g277_p
  (
    .dout(g277_p),
    .din1(ffc_57_p),
    .din2(g276_n_spl_00)
  );


  andX
  g_g278_p
  (
    .dout(g278_p),
    .din1(ffc_91_n_spl_),
    .din2(ffc_93_n_spl_)
  );


  andX
  g_g279_p
  (
    .dout(g279_p),
    .din1(ffc_98_n_spl_),
    .din2(g278_p)
  );


  andX
  g_g280_p
  (
    .dout(g280_p),
    .din1(ffc_92_p_spl_),
    .din2(g279_p)
  );


  andX
  g_g281_p
  (
    .dout(g281_p),
    .din1(ffc_99_p_spl_),
    .din2(g280_p)
  );


  orX
  g_g282_n
  (
    .dout(g282_n),
    .din1(ffc_58_p_spl_0),
    .din2(g281_p)
  );


  orX
  g_g283_n
  (
    .dout(g283_n),
    .din1(g277_p),
    .din2(g282_n)
  );


  andX
  g_g284_p
  (
    .dout(g284_p),
    .din1(ffc_53_n_spl_00),
    .din2(ffc_70_p)
  );


  orX
  g_g284_n
  (
    .dout(g284_n),
    .din1(ffc_53_p_spl_0),
    .din2(ffc_70_n)
  );


  andX
  g_g285_p
  (
    .dout(g285_p),
    .din1(g276_n_spl_00),
    .din2(g284_p)
  );


  orX
  g_g285_n
  (
    .dout(g285_n),
    .din1(g276_p_spl_0),
    .din2(g284_n)
  );


  andX
  g_g286_p
  (
    .dout(g286_p),
    .din1(ffc_65_n),
    .din2(g285_n)
  );


  andX
  g_g287_p
  (
    .dout(g287_p),
    .din1(ffc_65_p),
    .din2(g285_p)
  );


  orX
  g_g288_n
  (
    .dout(g288_n),
    .din1(g286_p),
    .din2(g287_p)
  );


  andX
  g_g289_p
  (
    .dout(g289_p),
    .din1(ffc_97_p_spl_00),
    .din2(g288_n)
  );


  andX
  g_g290_p
  (
    .dout(g290_p),
    .din1(ffc_33_p),
    .din2(ffc_53_n_spl_00)
  );


  orX
  g_g290_n
  (
    .dout(g290_n),
    .din1(ffc_33_n),
    .din2(ffc_53_p_spl_0)
  );


  andX
  g_g291_p
  (
    .dout(g291_p),
    .din1(g276_n_spl_01),
    .din2(g290_p)
  );


  orX
  g_g291_n
  (
    .dout(g291_n),
    .din1(g276_p_spl_0),
    .din2(g290_n)
  );


  andX
  g_g292_p
  (
    .dout(g292_p),
    .din1(ffc_73_p),
    .din2(g291_n)
  );


  andX
  g_g293_p
  (
    .dout(g293_p),
    .din1(ffc_73_n),
    .din2(g291_p)
  );


  orX
  g_g294_n
  (
    .dout(g294_n),
    .din1(g292_p),
    .din2(g293_p)
  );


  andX
  g_g295_p
  (
    .dout(g295_p),
    .din1(ffc_97_p_spl_00),
    .din2(g294_n)
  );


  andX
  g_g296_p
  (
    .dout(g296_p),
    .din1(ffc_39_p),
    .din2(ffc_53_n_spl_0)
  );


  andX
  g_g297_p
  (
    .dout(g297_p),
    .din1(g276_n_spl_01),
    .din2(g296_p)
  );


  orX
  g_g298_n
  (
    .dout(g298_n),
    .din1(ffc_64_n),
    .din2(g297_p)
  );


  andX
  g_g299_p
  (
    .dout(g299_p),
    .din1(ffc_97_p_spl_01),
    .din2(g298_n)
  );


  andX
  g_g300_p
  (
    .dout(g300_p),
    .din1(ffc_42_p),
    .din2(ffc_53_n_spl_1)
  );


  andX
  g_g301_p
  (
    .dout(g301_p),
    .din1(g276_n_spl_1),
    .din2(g300_p)
  );


  orX
  g_g302_n
  (
    .dout(g302_n),
    .din1(ffc_59_n),
    .din2(g301_p)
  );


  andX
  g_g303_p
  (
    .dout(g303_p),
    .din1(ffc_97_p_spl_01),
    .din2(g302_n)
  );


  andX
  g_g304_p
  (
    .dout(g304_p),
    .din1(ffc_53_n_spl_1),
    .din2(ffc_62_p)
  );


  andX
  g_g305_p
  (
    .dout(g305_p),
    .din1(g276_n_spl_1),
    .din2(g304_p)
  );


  orX
  g_g306_n
  (
    .dout(g306_n),
    .din1(ffc_61_p),
    .din2(g305_p)
  );


  andX
  g_g307_p
  (
    .dout(g307_p),
    .din1(ffc_97_p_spl_1),
    .din2(g306_n)
  );


  andX
  g_g308_p
  (
    .dout(g308_p),
    .din1(ffc_25_p),
    .din2(ffc_46_p)
  );


  orX
  g_g308_n
  (
    .dout(g308_n),
    .din1(ffc_25_n),
    .din2(ffc_46_n)
  );


  andX
  g_g309_p
  (
    .dout(g309_p),
    .din1(ffc_58_n_spl_),
    .din2(g308_n)
  );


  orX
  g_g309_n
  (
    .dout(g309_n),
    .din1(ffc_58_p_spl_0),
    .din2(g308_p)
  );


  andX
  g_g310_p
  (
    .dout(g310_p),
    .din1(ffc_60_p),
    .din2(ffc_95_p)
  );


  orX
  g_g310_n
  (
    .dout(g310_n),
    .din1(ffc_60_n),
    .din2(ffc_95_n)
  );


  andX
  g_g311_p
  (
    .dout(g311_p),
    .din1(g218_p_spl_10),
    .din2(g310_n_spl_)
  );


  orX
  g_g311_n
  (
    .dout(g311_n),
    .din1(g218_n_spl_10),
    .din2(g310_p_spl_)
  );


  andX
  g_g312_p
  (
    .dout(g312_p),
    .din1(g218_n_spl_1),
    .din2(g310_p_spl_)
  );


  orX
  g_g312_n
  (
    .dout(g312_n),
    .din1(g218_p_spl_1),
    .din2(g310_n_spl_)
  );


  andX
  g_g313_p
  (
    .dout(g313_p),
    .din1(g311_n),
    .din2(g312_n)
  );


  orX
  g_g313_n
  (
    .dout(g313_n),
    .din1(g311_p),
    .din2(g312_p)
  );


  andX
  g_g314_p
  (
    .dout(g314_p),
    .din1(g309_n),
    .din2(g313_n)
  );


  andX
  g_g315_p
  (
    .dout(g315_p),
    .din1(g309_p),
    .din2(g313_p)
  );


  orX
  g_g316_n
  (
    .dout(g316_n),
    .din1(g314_p),
    .din2(g315_p)
  );


  andX
  g_g317_p
  (
    .dout(g317_p),
    .din1(ffc_28_p),
    .din2(ffc_50_p)
  );


  orX
  g_g317_n
  (
    .dout(g317_n),
    .din1(ffc_28_n),
    .din2(ffc_50_n)
  );


  andX
  g_g318_p
  (
    .dout(g318_p),
    .din1(ffc_58_n_spl_),
    .din2(g317_n)
  );


  orX
  g_g318_n
  (
    .dout(g318_n),
    .din1(ffc_58_p_spl_),
    .din2(g317_p)
  );


  andX
  g_g319_p
  (
    .dout(g319_p),
    .din1(ffc_126_n),
    .din2(ffc_127_n)
  );


  orX
  g_g319_n
  (
    .dout(g319_n),
    .din1(ffc_126_p),
    .din2(ffc_127_p)
  );


  andX
  g_g320_p
  (
    .dout(g320_p),
    .din1(ffc_96_p),
    .din2(g319_n)
  );


  orX
  g_g320_n
  (
    .dout(g320_n),
    .din1(ffc_96_n),
    .din2(g319_p)
  );


  andX
  g_g321_p
  (
    .dout(g321_p),
    .din1(g231_p_spl_1),
    .din2(g320_n_spl_)
  );


  orX
  g_g321_n
  (
    .dout(g321_n),
    .din1(g231_n_spl_1),
    .din2(g320_p_spl_)
  );


  andX
  g_g322_p
  (
    .dout(g322_p),
    .din1(g231_n_spl_1),
    .din2(g320_p_spl_)
  );


  orX
  g_g322_n
  (
    .dout(g322_n),
    .din1(g231_p_spl_1),
    .din2(g320_n_spl_)
  );


  andX
  g_g323_p
  (
    .dout(g323_p),
    .din1(g321_n),
    .din2(g322_n)
  );


  orX
  g_g323_n
  (
    .dout(g323_n),
    .din1(g321_p),
    .din2(g322_p)
  );


  andX
  g_g324_p
  (
    .dout(g324_p),
    .din1(g318_n),
    .din2(g323_n)
  );


  andX
  g_g325_p
  (
    .dout(g325_p),
    .din1(g318_p),
    .din2(g323_p)
  );


  orX
  g_g326_n
  (
    .dout(g326_n),
    .din1(g324_p),
    .din2(g325_p)
  );


  orX
  g_g327_n
  (
    .dout(g327_n),
    .din1(ffc_36_n),
    .din2(ffc_53_p_spl_)
  );


  orX
  g_g328_n
  (
    .dout(g328_n),
    .din1(g276_p_spl_),
    .din2(g327_n)
  );


  andX
  g_g329_p
  (
    .dout(g329_p),
    .din1(ffc_63_n),
    .din2(g328_n)
  );


  andX
  g_g330_p
  (
    .dout(g330_p),
    .din1(ffc_97_p_spl_1),
    .din2(g329_p)
  );


  andX
  g_g331_p
  (
    .dout(g331_p),
    .din1(ffc_90_p),
    .din2(ffc_142_p)
  );


  orX
  g_g331_n
  (
    .dout(g331_n),
    .din1(ffc_90_n),
    .din2(ffc_142_n_spl_)
  );


  andX
  g_g332_p
  (
    .dout(g332_p),
    .din1(ffc_150_n),
    .din2(ffc_151_n)
  );


  orX
  g_g332_n
  (
    .dout(g332_n),
    .din1(ffc_150_p),
    .din2(ffc_151_p)
  );


  orX
  g_g333_n
  (
    .dout(g333_n),
    .din1(ffc_71_n),
    .din2(ffc_142_n_spl_)
  );


  andX
  g_g334_p
  (
    .dout(g334_p),
    .din1(ffc_102_n_spl_),
    .din2(ffc_152_n)
  );


  orX
  g_g334_n
  (
    .dout(g334_n),
    .din1(ffc_102_p_spl_0),
    .din2(ffc_152_p_spl_)
  );


  orX
  g_g335_n
  (
    .dout(g335_n),
    .din1(g331_p_spl_),
    .din2(g334_n)
  );


  orX
  g_g336_n
  (
    .dout(g336_n),
    .din1(g331_n),
    .din2(g334_p)
  );


  andX
  g_g337_p
  (
    .dout(g337_p),
    .din1(g335_n),
    .din2(g336_n)
  );


  orX
  g_g338_n
  (
    .dout(g338_n),
    .din1(ffc_87_n),
    .din2(ffc_111_n)
  );


  orX
  g_g339_n
  (
    .dout(g339_n),
    .din1(ffc_45_p_spl_),
    .din2(ffc_81_p_spl_0)
  );


  orX
  g_g340_n
  (
    .dout(g340_n),
    .din1(ffc_49_p_spl_),
    .din2(ffc_81_p_spl_0)
  );


  orX
  g_g341_n
  (
    .dout(g341_n),
    .din1(ffc_56_p_spl_),
    .din2(ffc_81_p_spl_1)
  );


  andX
  g_g342_p
  (
    .dout(g342_p),
    .din1(ffc_102_n_spl_),
    .din2(g332_n_spl_)
  );


  orX
  g_g342_n
  (
    .dout(g342_n),
    .din1(ffc_102_p_spl_0),
    .din2(g332_p)
  );


  orX
  g_g343_n
  (
    .dout(g343_n),
    .din1(ffc_32_p_spl_),
    .din2(g342_n)
  );


  orX
  g_g344_n
  (
    .dout(g344_n),
    .din1(ffc_32_n),
    .din2(g342_p)
  );


  andX
  g_g345_p
  (
    .dout(g345_p),
    .din1(g343_n),
    .din2(g344_n)
  );


  orX
  g_g346_n
  (
    .dout(g346_n),
    .din1(ffc_141_p_spl_),
    .din2(ffc_143_n)
  );


  andX
  g_g347_p
  (
    .dout(g347_p),
    .din1(ffc_146_n),
    .din2(ffc_147_n)
  );


  andX
  g_g348_p
  (
    .dout(g348_p),
    .din1(ffc_148_p),
    .din2(ffc_149_n)
  );


  andX
  g_g349_p
  (
    .dout(g349_p),
    .din1(g347_p),
    .din2(g348_p)
  );


  andX
  g_g350_p
  (
    .dout(g350_p),
    .din1(g346_n),
    .din2(g349_p)
  );


  orX
  g_g351_n
  (
    .dout(g351_n),
    .din1(ffc_140_n),
    .din2(ffc_144_n)
  );


  orX
  g_g352_n
  (
    .dout(g352_n),
    .din1(ffc_140_p_spl_),
    .din2(ffc_144_p)
  );


  orX
  g_g353_n
  (
    .dout(g353_n),
    .din1(ffc_141_n),
    .din2(ffc_143_p)
  );


  andX
  g_g354_p
  (
    .dout(g354_p),
    .din1(g352_n),
    .din2(g353_n)
  );


  andX
  g_g355_p
  (
    .dout(g355_p),
    .din1(g351_n),
    .din2(g354_p)
  );


  andX
  g_g356_p
  (
    .dout(g356_p),
    .din1(g350_p),
    .din2(g355_p)
  );


  andX
  g_g357_p
  (
    .dout(g357_p),
    .din1(ffc_168_n),
    .din2(ffc_169_n)
  );


  orX
  g_g357_n
  (
    .dout(g357_n),
    .din1(ffc_168_p),
    .din2(ffc_169_p)
  );


  orX
  g_g358_n
  (
    .dout(g358_n),
    .din1(g338_n_spl_),
    .din2(g345_p_spl_)
  );


  orX
  g_g359_n
  (
    .dout(g359_n),
    .din1(g333_n_spl_),
    .din2(g337_p_spl_)
  );


  andX
  g_g360_p
  (
    .dout(g360_p),
    .din1(g356_p_spl_),
    .din2(g359_n)
  );


  orX
  g_g361_n
  (
    .dout(g361_n),
    .din1(ffc_52_p_spl_0),
    .din2(ffc_138_p_spl_0)
  );


  andX
  g_g362_p
  (
    .dout(g362_p),
    .din1(ffc_162_n_spl_),
    .din2(ffc_163_p_spl_)
  );


  orX
  g_g362_n
  (
    .dout(g362_n),
    .din1(ffc_162_p_spl_),
    .din2(ffc_163_n_spl_)
  );


  andX
  g_g363_p
  (
    .dout(g363_p),
    .din1(ffc_162_p_spl_),
    .din2(ffc_163_n_spl_)
  );


  orX
  g_g363_n
  (
    .dout(g363_n),
    .din1(ffc_162_n_spl_),
    .din2(ffc_163_p_spl_)
  );


  andX
  g_g364_p
  (
    .dout(g364_p),
    .din1(g362_n),
    .din2(g363_n)
  );


  orX
  g_g364_n
  (
    .dout(g364_n),
    .din1(g362_p),
    .din2(g363_p)
  );


  andX
  g_g365_p
  (
    .dout(g365_p),
    .din1(ffc_138_n),
    .din2(ffc_161_p_spl_)
  );


  orX
  g_g365_n
  (
    .dout(g365_n),
    .din1(ffc_138_p_spl_0),
    .din2(ffc_161_n)
  );


  andX
  g_g366_p
  (
    .dout(g366_p),
    .din1(ffc_119_n_spl_0),
    .din2(g365_p)
  );


  orX
  g_g366_n
  (
    .dout(g366_n),
    .din1(ffc_119_p_spl_00),
    .din2(g365_n)
  );


  andX
  g_g367_p
  (
    .dout(g367_p),
    .din1(g364_n),
    .din2(g366_n)
  );


  andX
  g_g368_p
  (
    .dout(g368_p),
    .din1(g364_p),
    .din2(g366_p)
  );


  orX
  g_g369_n
  (
    .dout(g369_n),
    .din1(g367_p),
    .din2(g368_p)
  );


  andX
  g_g370_p
  (
    .dout(g370_p),
    .din1(ffc_164_n_spl_0),
    .din2(ffc_166_p_spl_)
  );


  orX
  g_g370_n
  (
    .dout(g370_n),
    .din1(ffc_164_p_spl_0),
    .din2(ffc_166_n_spl_)
  );


  andX
  g_g371_p
  (
    .dout(g371_p),
    .din1(ffc_164_p_spl_0),
    .din2(ffc_166_n_spl_)
  );


  orX
  g_g371_n
  (
    .dout(g371_n),
    .din1(ffc_164_n_spl_0),
    .din2(ffc_166_p_spl_)
  );


  andX
  g_g372_p
  (
    .dout(g372_p),
    .din1(g370_n),
    .din2(g371_n)
  );


  orX
  g_g372_n
  (
    .dout(g372_n),
    .din1(g370_p),
    .din2(g371_p)
  );


  andX
  g_g373_p
  (
    .dout(g373_p),
    .din1(ffc_107_n_spl_),
    .din2(ffc_158_p_spl_)
  );


  orX
  g_g373_n
  (
    .dout(g373_n),
    .din1(ffc_107_p_spl_0),
    .din2(ffc_158_n_spl_)
  );


  andX
  g_g374_p
  (
    .dout(g374_p),
    .din1(ffc_107_p_spl_0),
    .din2(ffc_158_n_spl_)
  );


  orX
  g_g374_n
  (
    .dout(g374_n),
    .din1(ffc_107_n_spl_),
    .din2(ffc_158_p_spl_)
  );


  andX
  g_g375_p
  (
    .dout(g375_p),
    .din1(g373_n),
    .din2(g374_n)
  );


  orX
  g_g375_n
  (
    .dout(g375_n),
    .din1(g373_p),
    .din2(g374_p)
  );


  orX
  g_g376_n
  (
    .dout(g376_n),
    .din1(g372_p),
    .din2(g375_p)
  );


  orX
  g_g377_n
  (
    .dout(g377_n),
    .din1(g372_n),
    .din2(g375_n)
  );


  andX
  g_g378_p
  (
    .dout(g378_p),
    .din1(g376_n),
    .din2(g377_n)
  );


  andX
  g_g379_p
  (
    .dout(g379_p),
    .din1(ffc_165_p_spl_0),
    .din2(ffc_167_p_spl_0)
  );


  orX
  g_g379_n
  (
    .dout(g379_n),
    .din1(ffc_165_n_spl_0),
    .din2(ffc_167_n_spl_0)
  );


  andX
  g_g380_p
  (
    .dout(g380_p),
    .din1(ffc_165_n_spl_0),
    .din2(ffc_167_n_spl_0)
  );


  orX
  g_g380_n
  (
    .dout(g380_n),
    .din1(ffc_165_p_spl_0),
    .din2(ffc_167_p_spl_0)
  );


  andX
  g_g381_p
  (
    .dout(g381_p),
    .din1(g379_n),
    .din2(g380_n)
  );


  orX
  g_g381_n
  (
    .dout(g381_n),
    .din1(g379_p),
    .din2(g380_p)
  );


  andX
  g_g382_p
  (
    .dout(g382_p),
    .din1(ffc_116_n_spl_),
    .din2(ffc_135_p_spl_00)
  );


  orX
  g_g382_n
  (
    .dout(g382_n),
    .din1(ffc_116_p_spl_0),
    .din2(ffc_135_n_spl_0)
  );


  andX
  g_g383_p
  (
    .dout(g383_p),
    .din1(ffc_116_p_spl_0),
    .din2(ffc_135_n_spl_0)
  );


  orX
  g_g383_n
  (
    .dout(g383_n),
    .din1(ffc_116_n_spl_),
    .din2(ffc_135_p_spl_00)
  );


  andX
  g_g384_p
  (
    .dout(g384_p),
    .din1(g382_n),
    .din2(g383_n)
  );


  orX
  g_g384_n
  (
    .dout(g384_n),
    .din1(g382_p),
    .din2(g383_p)
  );


  andX
  g_g385_p
  (
    .dout(g385_p),
    .din1(g381_n_spl_),
    .din2(g384_p_spl_)
  );


  orX
  g_g385_n
  (
    .dout(g385_n),
    .din1(g381_p_spl_),
    .din2(g384_n_spl_)
  );


  andX
  g_g386_p
  (
    .dout(g386_p),
    .din1(g381_p_spl_),
    .din2(g384_n_spl_)
  );


  orX
  g_g386_n
  (
    .dout(g386_n),
    .din1(g381_n_spl_),
    .din2(g384_p_spl_)
  );


  andX
  g_g387_p
  (
    .dout(g387_p),
    .din1(g385_n),
    .din2(g386_n)
  );


  orX
  g_g387_n
  (
    .dout(g387_n),
    .din1(g385_p),
    .din2(g386_p)
  );


  andX
  g_g388_p
  (
    .dout(g388_p),
    .din1(ffc_89_n),
    .din2(ffc_100_p)
  );


  andX
  g_g389_p
  (
    .dout(g389_p),
    .din1(ffc_89_p),
    .din2(ffc_100_n)
  );


  andX
  g_g390_p
  (
    .dout(g390_p),
    .din1(ffc_161_p_spl_),
    .din2(g361_n_spl_)
  );


  andX
  g_g391_p
  (
    .dout(g391_p),
    .din1(ffc_72_p),
    .din2(ffc_88_n)
  );


  orX
  g_g392_n
  (
    .dout(g392_n),
    .din1(ffc_102_p_spl_1),
    .din2(g391_p_spl_)
  );


  orX
  g_g393_n
  (
    .dout(g393_n),
    .din1(g339_n_spl_),
    .din2(g392_n_spl_)
  );


  orX
  g_g394_n
  (
    .dout(g394_n),
    .din1(g341_n_spl_),
    .din2(g391_p_spl_)
  );


  andX
  g_g395_p
  (
    .dout(g395_p),
    .din1(g393_n),
    .din2(g394_n_spl_)
  );


  orX
  g_g396_n
  (
    .dout(g396_n),
    .din1(g340_n_spl_),
    .din2(g392_n_spl_)
  );


  andX
  g_g397_p
  (
    .dout(g397_p),
    .din1(g394_n_spl_),
    .din2(g396_n)
  );


  andX
  g_g398_p
  (
    .dout(g398_p),
    .din1(g358_n_spl_),
    .din2(g360_p_spl_)
  );


  andX
  g_g399_p
  (
    .dout(g399_p),
    .din1(ffc_159_n),
    .din2(ffc_160_n)
  );


  orX
  g_g399_n
  (
    .dout(g399_n),
    .din1(ffc_159_p),
    .din2(ffc_160_p)
  );


  andX
  g_g400_p
  (
    .dout(g400_p),
    .din1(ffc_164_p_spl_1),
    .din2(g399_p_spl_)
  );


  orX
  g_g400_n
  (
    .dout(g400_n),
    .din1(ffc_164_n_spl_1),
    .din2(g399_n_spl_)
  );


  andX
  g_g401_p
  (
    .dout(g401_p),
    .din1(ffc_164_n_spl_1),
    .din2(g399_n_spl_)
  );


  orX
  g_g401_n
  (
    .dout(g401_n),
    .din1(ffc_164_p_spl_1),
    .din2(g399_p_spl_)
  );


  andX
  g_g402_p
  (
    .dout(g402_p),
    .din1(g400_n),
    .din2(g401_n)
  );


  orX
  g_g402_n
  (
    .dout(g402_n),
    .din1(g400_p),
    .din2(g401_p)
  );


  andX
  g_g403_p
  (
    .dout(g403_p),
    .din1(ffc_156_n),
    .din2(ffc_157_n)
  );


  orX
  g_g403_n
  (
    .dout(g403_n),
    .din1(ffc_156_p),
    .din2(ffc_157_p)
  );


  andX
  g_g404_p
  (
    .dout(g404_p),
    .din1(ffc_112_n_spl_),
    .din2(g403_n_spl_)
  );


  orX
  g_g404_n
  (
    .dout(g404_n),
    .din1(ffc_112_p_spl_0),
    .din2(g403_p_spl_)
  );


  andX
  g_g405_p
  (
    .dout(g405_p),
    .din1(ffc_112_p_spl_0),
    .din2(g403_p_spl_)
  );


  orX
  g_g405_n
  (
    .dout(g405_n),
    .din1(ffc_112_n_spl_),
    .din2(g403_n_spl_)
  );


  andX
  g_g406_p
  (
    .dout(g406_p),
    .din1(g404_n),
    .din2(g405_n)
  );


  orX
  g_g406_n
  (
    .dout(g406_n),
    .din1(g404_p),
    .din2(g405_p)
  );


  andX
  g_g407_p
  (
    .dout(g407_p),
    .din1(g402_n),
    .din2(g406_p)
  );


  andX
  g_g408_p
  (
    .dout(g408_p),
    .din1(g402_p),
    .din2(g406_n)
  );


  orX
  g_g409_n
  (
    .dout(g409_n),
    .din1(g407_p),
    .din2(g408_p)
  );


  andX
  g_g410_p
  (
    .dout(g410_p),
    .din1(ffc_119_n_spl_0),
    .din2(ffc_155_p)
  );


  orX
  g_g410_n
  (
    .dout(g410_n),
    .din1(ffc_119_p_spl_00),
    .din2(ffc_155_n)
  );


  andX
  g_g411_p
  (
    .dout(g411_p),
    .din1(ffc_134_p_spl_0),
    .din2(g410_p_spl_)
  );


  orX
  g_g411_n
  (
    .dout(g411_n),
    .din1(ffc_134_n_spl_),
    .din2(g410_n_spl_)
  );


  andX
  g_g412_p
  (
    .dout(g412_p),
    .din1(ffc_134_n_spl_),
    .din2(g410_n_spl_)
  );


  orX
  g_g412_n
  (
    .dout(g412_n),
    .din1(ffc_134_p_spl_0),
    .din2(g410_p_spl_)
  );


  andX
  g_g413_p
  (
    .dout(g413_p),
    .din1(g411_n),
    .din2(g412_n)
  );


  orX
  g_g413_n
  (
    .dout(g413_n),
    .din1(g411_p),
    .din2(g412_p)
  );


  andX
  g_g414_p
  (
    .dout(g414_p),
    .din1(ffc_167_p_spl_1),
    .din2(g357_p_spl_0)
  );


  orX
  g_g414_n
  (
    .dout(g414_n),
    .din1(ffc_167_n_spl_1),
    .din2(g357_n_spl_0)
  );


  andX
  g_g415_p
  (
    .dout(g415_p),
    .din1(ffc_167_n_spl_1),
    .din2(g357_n_spl_0)
  );


  orX
  g_g415_n
  (
    .dout(g415_n),
    .din1(ffc_167_p_spl_1),
    .din2(g357_p_spl_0)
  );


  andX
  g_g416_p
  (
    .dout(g416_p),
    .din1(g414_n),
    .din2(g415_n)
  );


  orX
  g_g416_n
  (
    .dout(g416_n),
    .din1(g414_p),
    .din2(g415_p)
  );


  andX
  g_g417_p
  (
    .dout(g417_p),
    .din1(g413_p),
    .din2(g416_n)
  );


  andX
  g_g418_p
  (
    .dout(g418_p),
    .din1(g413_n),
    .din2(g416_p)
  );


  orX
  g_g419_n
  (
    .dout(g419_n),
    .din1(g417_p),
    .din2(g418_p)
  );


  andX
  g_g420_p
  (
    .dout(g420_p),
    .din1(ffc_175_n_spl_),
    .din2(ffc_176_n_spl_)
  );


  orX
  g_g420_n
  (
    .dout(g420_n),
    .din1(ffc_175_p_spl_0),
    .din2(ffc_176_p_spl_0)
  );


  andX
  g_g421_p
  (
    .dout(g421_p),
    .din1(ffc_175_p_spl_0),
    .din2(ffc_176_p_spl_0)
  );


  orX
  g_g421_n
  (
    .dout(g421_n),
    .din1(ffc_175_n_spl_),
    .din2(ffc_176_n_spl_)
  );


  andX
  g_g422_p
  (
    .dout(g422_p),
    .din1(g420_n),
    .din2(g421_n)
  );


  orX
  g_g422_n
  (
    .dout(g422_n),
    .din1(g420_p),
    .din2(g421_p)
  );


  orX
  g_g423_n
  (
    .dout(g423_n),
    .din1(ffc_52_p_spl_0),
    .din2(ffc_110_p_spl_)
  );


  andX
  g_g424_p
  (
    .dout(g424_p),
    .din1(ffc_52_n_spl_0),
    .din2(g409_n_spl_)
  );


  andX
  g_g425_p
  (
    .dout(g425_p),
    .din1(ffc_52_n_spl_0),
    .din2(g419_n_spl_)
  );


  andX
  g_g426_p
  (
    .dout(g426_p),
    .din1(ffc_52_n_spl_),
    .din2(g369_n_spl_)
  );


  andX
  g_g427_p
  (
    .dout(g427_p),
    .din1(ffc_41_n_spl_),
    .din2(g426_p_spl_)
  );


  orX
  g_g428_n
  (
    .dout(g428_n),
    .din1(ffc_41_n_spl_),
    .din2(g426_p_spl_)
  );


  orX
  g_g429_n
  (
    .dout(g429_n),
    .din1(ffc_52_p_spl_1),
    .din2(g378_p_spl_)
  );


  orX
  g_g430_n
  (
    .dout(g430_n),
    .din1(g390_p_spl_0),
    .din2(g429_n_spl_)
  );


  andX
  g_g431_p
  (
    .dout(g431_p),
    .din1(g390_p_spl_0),
    .din2(g429_n_spl_)
  );


  andX
  g_g432_p
  (
    .dout(g432_p),
    .din1(ffc_27_p_spl_),
    .din2(ffc_119_n_spl_1)
  );


  orX
  g_g432_n
  (
    .dout(g432_n),
    .din1(ffc_27_n),
    .din2(ffc_119_p_spl_0)
  );


  andX
  g_g433_p
  (
    .dout(g433_p),
    .din1(ffc_118_n_spl_),
    .din2(ffc_135_n_spl_1)
  );


  orX
  g_g433_n
  (
    .dout(g433_n),
    .din1(ffc_118_p_spl_0),
    .din2(ffc_135_p_spl_0)
  );


  andX
  g_g434_p
  (
    .dout(g434_p),
    .din1(ffc_118_p_spl_0),
    .din2(ffc_135_p_spl_1)
  );


  orX
  g_g434_n
  (
    .dout(g434_n),
    .din1(ffc_118_n_spl_),
    .din2(ffc_135_n_spl_1)
  );


  andX
  g_g435_p
  (
    .dout(g435_p),
    .din1(g433_n),
    .din2(g434_n)
  );


  orX
  g_g435_n
  (
    .dout(g435_n),
    .din1(g433_p),
    .din2(g434_p)
  );


  andX
  g_g436_p
  (
    .dout(g436_p),
    .din1(g432_p),
    .din2(g435_n)
  );


  andX
  g_g437_p
  (
    .dout(g437_p),
    .din1(g432_n),
    .din2(g435_p)
  );


  orX
  g_g438_n
  (
    .dout(g438_n),
    .din1(g436_p),
    .din2(g437_p)
  );


  orX
  g_g439_n
  (
    .dout(g439_n),
    .din1(ffc_165_n_spl_),
    .din2(g357_n_spl_1)
  );


  orX
  g_g440_n
  (
    .dout(g440_n),
    .din1(ffc_165_p_spl_),
    .din2(g357_p_spl_)
  );


  andX
  g_g441_p
  (
    .dout(g441_p),
    .din1(g439_n),
    .din2(g440_n)
  );


  andX
  g_g442_p
  (
    .dout(g442_p),
    .din1(g438_n_spl_),
    .din2(g441_p_spl_)
  );


  orX
  g_g443_n
  (
    .dout(g443_n),
    .din1(g438_n_spl_),
    .din2(g441_p_spl_)
  );


  andX
  g_g444_p
  (
    .dout(g444_p),
    .din1(ffc_119_n_spl_1),
    .din2(ffc_154_p_spl_)
  );


  orX
  g_g444_n
  (
    .dout(g444_n),
    .din1(ffc_119_p_spl_1),
    .din2(ffc_154_n)
  );


  andX
  g_g445_p
  (
    .dout(g445_p),
    .din1(ffc_117_p_spl_0),
    .din2(ffc_153_n_spl_)
  );


  orX
  g_g445_n
  (
    .dout(g445_n),
    .din1(ffc_117_n_spl_),
    .din2(ffc_153_p_spl_)
  );


  andX
  g_g446_p
  (
    .dout(g446_p),
    .din1(ffc_117_n_spl_),
    .din2(ffc_153_p_spl_)
  );


  orX
  g_g446_n
  (
    .dout(g446_n),
    .din1(ffc_117_p_spl_0),
    .din2(ffc_153_n_spl_)
  );


  andX
  g_g447_p
  (
    .dout(g447_p),
    .din1(g445_n),
    .din2(g446_n)
  );


  orX
  g_g447_n
  (
    .dout(g447_n),
    .din1(g445_p),
    .din2(g446_p)
  );


  andX
  g_g448_p
  (
    .dout(g448_p),
    .din1(g444_p_spl_),
    .din2(g447_n_spl_)
  );


  orX
  g_g448_n
  (
    .dout(g448_n),
    .din1(g444_n_spl_),
    .din2(g447_p_spl_)
  );


  andX
  g_g449_p
  (
    .dout(g449_p),
    .din1(g444_n_spl_),
    .din2(g447_p_spl_)
  );


  orX
  g_g449_n
  (
    .dout(g449_n),
    .din1(g444_p_spl_),
    .din2(g447_n_spl_)
  );


  andX
  g_g450_p
  (
    .dout(g450_p),
    .din1(g448_n),
    .din2(g449_n)
  );


  orX
  g_g450_n
  (
    .dout(g450_n),
    .din1(g448_p),
    .din2(g449_p)
  );


  andX
  g_g451_p
  (
    .dout(g451_p),
    .din1(g387_n),
    .din2(g450_p)
  );


  andX
  g_g452_p
  (
    .dout(g452_p),
    .din1(g387_p_spl_),
    .din2(g450_n)
  );


  orX
  g_g453_n
  (
    .dout(g453_n),
    .din1(g451_p),
    .din2(g452_p)
  );


  andX
  g_g454_p
  (
    .dout(g454_p),
    .din1(ffc_178_p_spl_00),
    .din2(ffc_181_n_spl_0)
  );


  orX
  g_g454_n
  (
    .dout(g454_n),
    .din1(ffc_178_n_spl_0),
    .din2(ffc_181_p_spl_0)
  );


  andX
  g_g455_p
  (
    .dout(g455_p),
    .din1(ffc_178_n_spl_0),
    .din2(ffc_181_p_spl_0)
  );


  orX
  g_g455_n
  (
    .dout(g455_n),
    .din1(ffc_178_p_spl_00),
    .din2(ffc_181_n_spl_0)
  );


  andX
  g_g456_p
  (
    .dout(g456_p),
    .din1(g454_n),
    .din2(g455_n)
  );


  orX
  g_g456_n
  (
    .dout(g456_n),
    .din1(g454_p),
    .din2(g455_p)
  );


  andX
  g_g457_p
  (
    .dout(g457_p),
    .din1(ffc_19_p_spl_0),
    .din2(g456_n_spl_)
  );


  andX
  g_g458_p
  (
    .dout(g458_p),
    .din1(ffc_19_n_spl_),
    .din2(g456_p_spl_)
  );


  orX
  g_g459_n
  (
    .dout(g459_n),
    .din1(g457_p),
    .din2(g458_p)
  );


  andX
  g_g460_p
  (
    .dout(g460_p),
    .din1(ffc_21_p_spl_),
    .din2(ffc_183_n_spl_)
  );


  andX
  g_g461_p
  (
    .dout(g461_p),
    .din1(ffc_6_p_spl_0),
    .din2(ffc_174_n_spl_0)
  );


  andX
  g_g462_p
  (
    .dout(g462_p),
    .din1(ffc_6_n_spl_),
    .din2(ffc_174_p_spl_0)
  );


  andX
  g_g463_p
  (
    .dout(g463_p),
    .din1(ffc_23_p_spl_),
    .din2(ffc_29_n)
  );


  andX
  g_g464_p
  (
    .dout(g464_p),
    .din1(ffc_177_n_spl_),
    .din2(g463_p)
  );


  andX
  g_g465_p
  (
    .dout(g465_p),
    .din1(ffc_182_p_spl_),
    .din2(ffc_183_n_spl_)
  );


  orX
  g_g465_n
  (
    .dout(g465_n),
    .din1(ffc_182_n),
    .din2(ffc_183_p_spl_)
  );


  andX
  g_g466_p
  (
    .dout(g466_p),
    .din1(ffc_177_n_spl_),
    .din2(g465_p)
  );


  orX
  g_g466_n
  (
    .dout(g466_n),
    .din1(ffc_177_p_spl_),
    .din2(g465_n)
  );


  andX
  g_g467_p
  (
    .dout(g467_p),
    .din1(ffc_181_p_spl_1),
    .din2(g466_n)
  );


  andX
  g_g468_p
  (
    .dout(g468_p),
    .din1(ffc_181_n_spl_),
    .din2(g466_p)
  );


  orX
  g_g469_n
  (
    .dout(g469_n),
    .din1(g467_p),
    .din2(g468_p)
  );


  andX
  g_g470_p
  (
    .dout(g470_p),
    .din1(ffc_13_n_spl_0),
    .din2(g469_n_spl_)
  );


  orX
  g_g471_n
  (
    .dout(g471_n),
    .din1(ffc_13_n_spl_0),
    .din2(g469_n_spl_)
  );


  andX
  g_g472_p
  (
    .dout(g472_p),
    .din1(ffc_179_n_spl_0),
    .din2(g456_n_spl_)
  );


  andX
  g_g473_p
  (
    .dout(g473_p),
    .din1(ffc_179_p_spl_0),
    .din2(g456_p_spl_)
  );


  orX
  g_g474_n
  (
    .dout(g474_n),
    .din1(g472_p),
    .din2(g473_p)
  );


  andX
  g_g475_p
  (
    .dout(g475_p),
    .din1(ffc_172_p_spl_00),
    .din2(ffc_174_n_spl_0)
  );


  orX
  g_g475_n
  (
    .dout(g475_n),
    .din1(ffc_172_n_spl_0),
    .din2(ffc_174_p_spl_0)
  );


  andX
  g_g476_p
  (
    .dout(g476_p),
    .din1(ffc_172_n_spl_0),
    .din2(ffc_174_p_spl_1)
  );


  orX
  g_g476_n
  (
    .dout(g476_n),
    .din1(ffc_172_p_spl_00),
    .din2(ffc_174_n_spl_)
  );


  andX
  g_g477_p
  (
    .dout(g477_p),
    .din1(g475_n),
    .din2(g476_n)
  );


  orX
  g_g477_n
  (
    .dout(g477_n),
    .din1(g475_p),
    .din2(g476_p)
  );


  andX
  g_g478_p
  (
    .dout(g478_p),
    .din1(ffc_171_n_spl_0),
    .din2(g477_n)
  );


  andX
  g_g479_p
  (
    .dout(g479_p),
    .din1(ffc_171_p_spl_0),
    .din2(g477_p)
  );


  orX
  g_g480_n
  (
    .dout(g480_n),
    .din1(g478_p),
    .din2(g479_p)
  );


  andX
  g_g481_p
  (
    .dout(g481_p),
    .din1(ffc_19_p_spl_0),
    .din2(g422_n)
  );


  andX
  g_g482_p
  (
    .dout(g482_p),
    .din1(ffc_19_n_spl_),
    .din2(g422_p_spl_)
  );


  orX
  g_g483_n
  (
    .dout(g483_n),
    .din1(g481_p),
    .din2(g482_p)
  );


  andX
  g_g484_p
  (
    .dout(g484_p),
    .din1(ffc_170_n_spl_),
    .din2(ffc_171_n_spl_0)
  );


  orX
  g_g484_n
  (
    .dout(g484_n),
    .din1(ffc_170_p_spl_0),
    .din2(ffc_171_p_spl_0)
  );


  andX
  g_g485_p
  (
    .dout(g485_p),
    .din1(ffc_170_p_spl_0),
    .din2(ffc_171_p_spl_1)
  );


  orX
  g_g485_n
  (
    .dout(g485_n),
    .din1(ffc_170_n_spl_),
    .din2(ffc_171_n_spl_)
  );


  andX
  g_g486_p
  (
    .dout(g486_p),
    .din1(g484_n),
    .din2(g485_n)
  );


  orX
  g_g486_n
  (
    .dout(g486_n),
    .din1(g484_p),
    .din2(g485_p)
  );


  andX
  g_g487_p
  (
    .dout(g487_p),
    .din1(ffc_0_p_spl_),
    .din2(g486_n)
  );


  andX
  g_g488_p
  (
    .dout(g488_p),
    .din1(ffc_0_n),
    .din2(g486_p)
  );


  orX
  g_g489_n
  (
    .dout(g489_n),
    .din1(g487_p),
    .din2(g488_p)
  );


  andX
  g_g490_p
  (
    .dout(g490_p),
    .din1(ffc_173_p_spl_00),
    .din2(ffc_178_n_spl_1)
  );


  orX
  g_g490_n
  (
    .dout(g490_n),
    .din1(ffc_173_n_spl_0),
    .din2(ffc_178_p_spl_0)
  );


  andX
  g_g491_p
  (
    .dout(g491_p),
    .din1(ffc_173_n_spl_0),
    .din2(ffc_178_p_spl_1)
  );


  orX
  g_g491_n
  (
    .dout(g491_n),
    .din1(ffc_173_p_spl_00),
    .din2(ffc_178_n_spl_1)
  );


  andX
  g_g492_p
  (
    .dout(g492_p),
    .din1(g490_n),
    .din2(g491_n)
  );


  orX
  g_g492_n
  (
    .dout(g492_n),
    .din1(g490_p),
    .din2(g491_p)
  );


  andX
  g_g493_p
  (
    .dout(g493_p),
    .din1(ffc_4_n),
    .din2(g492_n)
  );


  andX
  g_g494_p
  (
    .dout(g494_p),
    .din1(ffc_4_p_spl_),
    .din2(g492_p)
  );


  orX
  g_g495_n
  (
    .dout(g495_n),
    .din1(g493_p),
    .din2(g494_p)
  );


  andX
  g_g496_p
  (
    .dout(g496_p),
    .din1(ffc_172_n_spl_1),
    .din2(ffc_173_n_spl_1)
  );


  orX
  g_g496_n
  (
    .dout(g496_n),
    .din1(ffc_172_p_spl_0),
    .din2(ffc_173_p_spl_0)
  );


  andX
  g_g497_p
  (
    .dout(g497_p),
    .din1(ffc_172_p_spl_1),
    .din2(ffc_173_p_spl_1)
  );


  orX
  g_g497_n
  (
    .dout(g497_n),
    .din1(ffc_172_n_spl_1),
    .din2(ffc_173_n_spl_1)
  );


  andX
  g_g498_p
  (
    .dout(g498_p),
    .din1(g496_n),
    .din2(g497_n)
  );


  orX
  g_g498_n
  (
    .dout(g498_n),
    .din1(g496_p),
    .din2(g497_p)
  );


  andX
  g_g499_p
  (
    .dout(g499_p),
    .din1(ffc_6_p_spl_0),
    .din2(g498_n)
  );


  andX
  g_g500_p
  (
    .dout(g500_p),
    .din1(ffc_6_n_spl_),
    .din2(g498_p)
  );


  orX
  g_g501_n
  (
    .dout(g501_n),
    .din1(g499_p),
    .din2(g500_p)
  );


  andX
  g_g502_p
  (
    .dout(g502_p),
    .din1(ffc_179_n_spl_0),
    .din2(ffc_180_n_spl_)
  );


  orX
  g_g502_n
  (
    .dout(g502_n),
    .din1(ffc_179_p_spl_0),
    .din2(ffc_180_p_spl_0)
  );


  andX
  g_g503_p
  (
    .dout(g503_p),
    .din1(ffc_179_p_spl_1),
    .din2(ffc_180_p_spl_0)
  );


  orX
  g_g503_n
  (
    .dout(g503_n),
    .din1(ffc_179_n_spl_),
    .din2(ffc_180_n_spl_)
  );


  andX
  g_g504_p
  (
    .dout(g504_p),
    .din1(g502_n),
    .din2(g503_n)
  );


  orX
  g_g504_n
  (
    .dout(g504_n),
    .din1(g502_p),
    .din2(g503_p)
  );


  andX
  g_g505_p
  (
    .dout(g505_p),
    .din1(ffc_13_p_spl_),
    .din2(g504_n)
  );


  andX
  g_g506_p
  (
    .dout(g506_p),
    .din1(ffc_13_n_spl_),
    .din2(g504_p)
  );


  orX
  g_g507_n
  (
    .dout(g507_n),
    .din1(g505_p),
    .din2(g506_p)
  );


  andX
  g_g508_p
  (
    .dout(g508_p),
    .din1(g459_n_spl_0),
    .din2(g507_n_spl_)
  );


  orX
  g_g509_n
  (
    .dout(g509_n),
    .din1(g459_n_spl_0),
    .din2(g507_n_spl_)
  );


  buf

  (
    G1884_p,
    g221_n
  );


  buf

  (
    G1885_p,
    g224_n
  );


  buf

  (
    G1886_p,
    g227_n
  );


  buf

  (
    G1887_p,
    g230_n
  );


  buf

  (
    G1888_p,
    g234_n
  );


  buf

  (
    G1889_p,
    g237_n
  );


  buf

  (
    G1890_p,
    g240_n
  );


  buf

  (
    G1891_p,
    g246_n
  );


  buf

  (
    G1892_p,
    g249_n
  );


  buf

  (
    G1893_p,
    g252_n
  );


  buf

  (
    G1894_p,
    g255_n
  );


  buf

  (
    G1895_p,
    g259_n
  );


  buf

  (
    G1896_p,
    g266_n
  );


  buf

  (
    G1897_p,
    g269_n
  );


  buf

  (
    G1898_p,
    g272_n
  );


  buf

  (
    G1899_p,
    g275_n
  );


  buf

  (
    G1900_p,
    g283_n
  );


  buf

  (
    G1901_p,
    g289_p
  );


  buf

  (
    G1902_p,
    g295_p
  );


  buf

  (
    G1903_p,
    g299_p
  );


  buf

  (
    G1904_p,
    g303_p
  );


  buf

  (
    G1905_p,
    g307_p
  );


  buf

  (
    G1906_p,
    g316_n
  );


  buf

  (
    G1907_p,
    g326_n
  );


  buf

  (
    G1908_p,
    g330_p
  );


  DROC
  ffc_0
  (
    .doutp(ffc_0_p),
    .doutn(ffc_0_n),
    .din(G1_p)
  );


  DROC
  ffc_1
  (
    .doutp(ffc_1_p),
    .doutn(ffc_1_n),
    .din(ffc_84_p)
  );


  DROC
  ffc_2
  (
    .doutp(ffc_2_p),
    .doutn(ffc_2_n),
    .din(ffc_74_p)
  );


  DROC
  ffc_3
  (
    .doutp(ffc_3_p),
    .doutn(ffc_3_n),
    .din(ffc_75_p)
  );


  DROC
  ffc_4
  (
    .doutp(ffc_4_p),
    .doutn(ffc_4_n),
    .din(G4_p)
  );


  DROC
  ffc_5
  (
    .doutp(ffc_5_p),
    .doutn(ffc_5_n),
    .din(ffc_85_p)
  );


  DROC
  ffc_6
  (
    .doutp(ffc_6_p),
    .doutn(ffc_6_n),
    .din(G5_p)
  );


  DROC
  ffc_7
  (
    .doutp(ffc_7_p),
    .doutn(ffc_7_n),
    .din(ffc_86_p)
  );


  DROC
  ffc_8
  (
    .doutp(ffc_8_p),
    .doutn(ffc_8_n),
    .din(ffc_76_p)
  );


  DROC
  ffc_9
  (
    .doutp(ffc_9_p),
    .doutn(ffc_9_n),
    .din(ffc_77_p)
  );


  DROC
  ffc_10
  (
    .doutp(ffc_10_p),
    .doutn(ffc_10_n),
    .din(ffc_78_p)
  );


  DROC
  ffc_11
  (
    .doutp(ffc_11_p),
    .doutn(ffc_11_n),
    .din(ffc_79_p)
  );


  DROC
  ffc_12
  (
    .doutp(ffc_12_p),
    .doutn(ffc_12_n),
    .din(ffc_66_p)
  );


  DROC
  ffc_13
  (
    .doutp(ffc_13_p),
    .doutn(ffc_13_n),
    .din(G11_p)
  );


  DROC
  ffc_14
  (
    .doutp(ffc_14_p),
    .doutn(ffc_14_n),
    .din(ffc_82_p)
  );


  DROC
  ffc_15
  (
    .doutp(ffc_15_p),
    .doutn(ffc_15_n),
    .din(ffc_67_p)
  );


  DROC
  ffc_16
  (
    .doutp(ffc_16_p),
    .doutn(ffc_16_n),
    .din(ffc_68_p)
  );


  DROC
  ffc_17
  (
    .doutp(ffc_17_p),
    .doutn(ffc_17_n),
    .din(ffc_80_p)
  );


  DROC
  ffc_18
  (
    .doutp(ffc_18_p),
    .doutn(ffc_18_n),
    .din(ffc_69_p)
  );


  DROC
  ffc_19
  (
    .doutp(ffc_19_p),
    .doutn(ffc_19_n),
    .din(G16_p)
  );


  DROC
  ffc_20
  (
    .doutp(ffc_20_p),
    .doutn(ffc_20_n),
    .din(ffc_83_p)
  );


  DROC
  ffc_21
  (
    .doutp(ffc_21_p),
    .doutn(ffc_21_n),
    .din(G17_p)
  );


  DROC
  ffc_22
  (
    .doutp(ffc_22_p),
    .doutn(ffc_22_n),
    .din(G19_p)
  );


  DROC
  ffc_23
  (
    .doutp(ffc_23_p),
    .doutn(ffc_23_n),
    .din(G20_p)
  );


  DROC
  ffc_24
  (
    .doutp(ffc_24_p),
    .doutn(ffc_24_n),
    .din(G21_p)
  );


  DROC
  ffc_25
  (
    .doutp(ffc_25_p),
    .doutn(ffc_25_n),
    .din(ffc_94_p)
  );


  DROC
  ffc_26
  (
    .doutp(ffc_26_p),
    .doutn(ffc_26_n),
    .din(G22_p)
  );


  DROC
  ffc_27
  (
    .doutp(ffc_27_p),
    .doutn(ffc_27_n),
    .din(ffc_26_p)
  );


  DROC
  ffc_28
  (
    .doutp(ffc_28_p),
    .doutn(ffc_28_n),
    .din(ffc_101_p)
  );


  DROC
  ffc_29
  (
    .doutp(ffc_29_p),
    .doutn(ffc_29_n),
    .din(G23_p)
  );


  DROC
  ffc_30
  (
    .doutp(ffc_30_p),
    .doutn(ffc_30_n),
    .din(G25_p)
  );


  DROC
  ffc_31
  (
    .doutp(ffc_31_p),
    .doutn(ffc_31_n),
    .din(ffc_30_p)
  );


  DROC
  ffc_32
  (
    .doutp(ffc_32_p),
    .doutn(ffc_32_n),
    .din(ffc_31_p)
  );


  DROC
  ffc_33
  (
    .doutp(ffc_33_p),
    .doutn(ffc_33_n),
    .din(ffc_32_p_spl_)
  );


  DROC
  ffc_34
  (
    .doutp(ffc_34_p),
    .doutn(ffc_34_n),
    .din(G26_p)
  );


  DROC
  ffc_35
  (
    .doutp(ffc_35_p),
    .doutn(ffc_35_n),
    .din(ffc_34_p)
  );


  DROC
  ffc_36
  (
    .doutp(ffc_36_p),
    .doutn(ffc_36_n),
    .din(ffc_140_p_spl_)
  );


  DROC
  ffc_37
  (
    .doutp(ffc_37_p),
    .doutn(ffc_37_n),
    .din(G27_p)
  );


  DROC
  ffc_38
  (
    .doutp(ffc_38_p),
    .doutn(ffc_38_n),
    .din(ffc_37_p)
  );


  DROC
  ffc_39
  (
    .doutp(ffc_39_p),
    .doutn(ffc_39_n),
    .din(ffc_141_p_spl_)
  );


  DROC
  ffc_40
  (
    .doutp(ffc_40_p),
    .doutn(ffc_40_n),
    .din(G28_p)
  );


  DROC
  ffc_41
  (
    .doutp(ffc_41_p),
    .doutn(ffc_41_n),
    .din(ffc_40_p)
  );


  DROC
  ffc_42
  (
    .doutp(ffc_42_p),
    .doutn(ffc_42_n),
    .din(ffc_125_p)
  );


  DROC
  ffc_43
  (
    .doutp(ffc_43_p),
    .doutn(ffc_43_n),
    .din(G29_p)
  );


  DROC
  ffc_44
  (
    .doutp(ffc_44_p),
    .doutn(ffc_44_n),
    .din(ffc_43_p)
  );


  DROC
  ffc_45
  (
    .doutp(ffc_45_p),
    .doutn(ffc_45_n),
    .din(ffc_44_p)
  );


  DROC
  ffc_46
  (
    .doutp(ffc_46_p),
    .doutn(ffc_46_n),
    .din(ffc_45_p_spl_)
  );


  DROC
  ffc_47
  (
    .doutp(ffc_47_p),
    .doutn(ffc_47_n),
    .din(G30_p)
  );


  DROC
  ffc_48
  (
    .doutp(ffc_48_p),
    .doutn(ffc_48_n),
    .din(ffc_47_p)
  );


  DROC
  ffc_49
  (
    .doutp(ffc_49_p),
    .doutn(ffc_49_n),
    .din(ffc_48_p)
  );


  DROC
  ffc_50
  (
    .doutp(ffc_50_p),
    .doutn(ffc_50_n),
    .din(ffc_49_p_spl_)
  );


  DROC
  ffc_51
  (
    .doutp(ffc_51_p),
    .doutn(ffc_51_n),
    .din(G31_p)
  );


  DROC
  ffc_52
  (
    .doutp(ffc_52_p),
    .doutn(ffc_52_n),
    .din(ffc_51_p)
  );


  DROC
  ffc_53
  (
    .doutp(ffc_53_p),
    .doutn(ffc_53_n),
    .din(ffc_102_p_spl_1)
  );


  DROC
  ffc_54
  (
    .doutp(ffc_54_p),
    .doutn(ffc_54_n),
    .din(G32_p)
  );


  DROC
  ffc_55
  (
    .doutp(ffc_55_p),
    .doutn(ffc_55_n),
    .din(ffc_54_p)
  );


  DROC
  ffc_56
  (
    .doutp(ffc_56_p),
    .doutn(ffc_56_n),
    .din(ffc_55_p)
  );


  DROC
  ffc_57
  (
    .doutp(ffc_57_p),
    .doutn(ffc_57_n),
    .din(ffc_56_p_spl_)
  );


  DROC
  ffc_58
  (
    .doutp(ffc_58_p),
    .doutn(ffc_58_n),
    .din(ffc_81_p_spl_1)
  );


  DROC
  ffc_59
  (
    .doutp(ffc_59_p),
    .doutn(ffc_59_n),
    .din(ffc_120_p)
  );


  DROC
  ffc_60
  (
    .doutp(ffc_60_p),
    .doutn(ffc_60_n),
    .din(ffc_122_p)
  );


  DROC
  ffc_61
  (
    .doutp(ffc_61_p),
    .doutn(ffc_61_n),
    .din(ffc_121_p)
  );


  DROC
  ffc_62
  (
    .doutp(ffc_62_p),
    .doutn(ffc_62_n),
    .din(ffc_128_p)
  );


  DROC
  ffc_63
  (
    .doutp(ffc_63_p),
    .doutn(ffc_63_n),
    .din(ffc_133_p)
  );


  DROC
  ffc_64
  (
    .doutp(ffc_64_p),
    .doutn(ffc_64_n),
    .din(ffc_132_p)
  );


  DROC
  ffc_65
  (
    .doutp(ffc_65_p),
    .doutn(ffc_65_n),
    .din(ffc_152_p_spl_)
  );


  DROC
  ffc_66
  (
    .doutp(ffc_66_p),
    .doutn(ffc_66_n),
    .din(ffc_105_p)
  );


  DROC
  ffc_67
  (
    .doutp(ffc_67_p),
    .doutn(ffc_67_n),
    .din(ffc_106_p)
  );


  DROC
  ffc_68
  (
    .doutp(ffc_68_p),
    .doutn(ffc_68_n),
    .din(ffc_107_p_spl_)
  );


  DROC
  ffc_69
  (
    .doutp(ffc_69_p),
    .doutn(ffc_69_n),
    .din(ffc_108_p)
  );


  DROC
  ffc_70
  (
    .doutp(ffc_70_p),
    .doutn(ffc_70_n),
    .din(g331_p_spl_)
  );


  DROC
  ffc_71
  (
    .doutp(ffc_71_p),
    .doutn(ffc_71_n),
    .din(ffc_109_p)
  );


  DROC
  ffc_72
  (
    .doutp(ffc_72_p),
    .doutn(ffc_72_n),
    .din(ffc_110_p_spl_)
  );


  DROC
  ffc_73
  (
    .doutp(ffc_73_p),
    .doutn(ffc_73_n),
    .din(g332_n_spl_)
  );


  DROC
  ffc_74
  (
    .doutp(ffc_74_p),
    .doutn(ffc_74_n),
    .din(ffc_112_p_spl_)
  );


  DROC
  ffc_75
  (
    .doutp(ffc_75_p),
    .doutn(ffc_75_n),
    .din(ffc_113_p)
  );


  DROC
  ffc_76
  (
    .doutp(ffc_76_p),
    .doutn(ffc_76_n),
    .din(ffc_114_p)
  );


  DROC
  ffc_77
  (
    .doutp(ffc_77_p),
    .doutn(ffc_77_n),
    .din(ffc_115_p)
  );


  DROC
  ffc_78
  (
    .doutp(ffc_78_p),
    .doutn(ffc_78_n),
    .din(ffc_116_p_spl_)
  );


  DROC
  ffc_79
  (
    .doutp(ffc_79_p),
    .doutn(ffc_79_n),
    .din(ffc_117_p_spl_)
  );


  DROC
  ffc_80
  (
    .doutp(ffc_80_p),
    .doutn(ffc_80_n),
    .din(ffc_118_p_spl_)
  );


  DROC
  ffc_81
  (
    .doutp(ffc_81_p),
    .doutn(ffc_81_n),
    .din(ffc_119_p_spl_1)
  );


  DROC
  ffc_82
  (
    .doutp(ffc_82_p),
    .doutn(ffc_82_n),
    .din(ffc_123_p)
  );


  DROC
  ffc_83
  (
    .doutp(ffc_83_p),
    .doutn(ffc_83_n),
    .din(ffc_124_p)
  );


  DROC
  ffc_84
  (
    .doutp(ffc_84_p),
    .doutn(ffc_84_n),
    .din(ffc_134_p_spl_)
  );


  DROC
  ffc_85
  (
    .doutp(ffc_85_p),
    .doutn(ffc_85_n),
    .din(ffc_135_p_spl_1)
  );


  DROC
  ffc_86
  (
    .doutp(ffc_86_p),
    .doutn(ffc_86_n),
    .din(ffc_136_p)
  );


  DROC
  ffc_87
  (
    .doutp(ffc_87_p),
    .doutn(ffc_87_n),
    .din(ffc_137_p)
  );


  DROC
  ffc_88
  (
    .doutp(ffc_88_p),
    .doutn(ffc_88_n),
    .din(ffc_138_p_spl_)
  );


  DROC
  ffc_89
  (
    .doutp(ffc_89_p),
    .doutn(ffc_89_n),
    .din(ffc_139_p)
  );


  DROC
  ffc_90
  (
    .doutp(ffc_90_p),
    .doutn(ffc_90_n),
    .din(ffc_145_p)
  );


  DROC
  ffc_91
  (
    .doutp(ffc_91_n),
    .doutn(ffc_91_p),
    .din(g333_n_spl_)
  );


  DROC
  ffc_92
  (
    .doutp(ffc_92_p),
    .doutn(ffc_92_n),
    .din(g337_p_spl_)
  );


  DROC
  ffc_93
  (
    .doutp(ffc_93_n),
    .doutn(ffc_93_p),
    .din(g338_n_spl_)
  );


  DROC
  ffc_94
  (
    .doutp(ffc_94_p),
    .doutn(ffc_94_n),
    .din(ffc_154_p_spl_)
  );


  DROC
  ffc_95
  (
    .doutp(ffc_95_p),
    .doutn(ffc_95_n),
    .din(g339_n_spl_)
  );


  DROC
  ffc_96
  (
    .doutp(ffc_96_p),
    .doutn(ffc_96_n),
    .din(g340_n_spl_)
  );


  DROC
  ffc_97
  (
    .doutp(ffc_97_p),
    .doutn(ffc_97_n),
    .din(g341_n_spl_)
  );


  DROC
  ffc_98
  (
    .doutp(ffc_98_n),
    .doutn(ffc_98_p),
    .din(g345_p_spl_)
  );


  DROC
  ffc_99
  (
    .doutp(ffc_99_p),
    .doutn(ffc_99_n),
    .din(g356_p_spl_)
  );


  DROC
  ffc_100
  (
    .doutp(ffc_100_p),
    .doutn(ffc_100_n),
    .din(g357_n_spl_1)
  );


  DROC
  ffc_101
  (
    .doutp(ffc_101_p),
    .doutn(ffc_101_n),
    .din(ffc_27_p_spl_)
  );


  DROC
  ffc_102
  (
    .doutp(ffc_102_p),
    .doutn(ffc_102_n),
    .din(ffc_52_p_spl_1)
  );


  DROC
  ffc_103
  (
    .doutp(ffc_103_n),
    .doutn(ffc_103_p),
    .din(g358_n_spl_)
  );


  DROC
  ffc_104
  (
    .doutp(ffc_104_p),
    .doutn(ffc_104_n),
    .din(g360_p_spl_)
  );


  DROC
  ffc_105
  (
    .doutp(ffc_105_p),
    .doutn(ffc_105_n),
    .din(ffc_178_p_spl_1)
  );


  DROC
  ffc_106
  (
    .doutp(ffc_106_p),
    .doutn(ffc_106_n),
    .din(ffc_179_p_spl_1)
  );


  DROC
  ffc_107
  (
    .doutp(ffc_107_p),
    .doutn(ffc_107_n),
    .din(ffc_180_p_spl_)
  );


  DROC
  ffc_108
  (
    .doutp(ffc_108_p),
    .doutn(ffc_108_n),
    .din(ffc_181_p_spl_1)
  );


  DROC
  ffc_109
  (
    .doutp(ffc_109_p),
    .doutn(ffc_109_n),
    .din(ffc_182_p_spl_)
  );


  DROC
  ffc_110
  (
    .doutp(ffc_110_p),
    .doutn(ffc_110_n),
    .din(ffc_183_p_spl_)
  );


  DROC
  ffc_111
  (
    .doutp(ffc_111_p),
    .doutn(ffc_111_n),
    .din(g361_n_spl_)
  );


  DROC
  ffc_112
  (
    .doutp(ffc_112_p),
    .doutn(ffc_112_n),
    .din(ffc_170_p_spl_)
  );


  DROC
  ffc_113
  (
    .doutp(ffc_113_p),
    .doutn(ffc_113_n),
    .din(ffc_171_p_spl_1)
  );


  DROC
  ffc_114
  (
    .doutp(ffc_114_p),
    .doutn(ffc_114_n),
    .din(ffc_172_p_spl_1)
  );


  DROC
  ffc_115
  (
    .doutp(ffc_115_p),
    .doutn(ffc_115_n),
    .din(ffc_173_p_spl_1)
  );


  DROC
  ffc_116
  (
    .doutp(ffc_116_p),
    .doutn(ffc_116_n),
    .din(ffc_174_p_spl_1)
  );


  DROC
  ffc_117
  (
    .doutp(ffc_117_p),
    .doutn(ffc_117_n),
    .din(ffc_175_p_spl_)
  );


  DROC
  ffc_118
  (
    .doutp(ffc_118_p),
    .doutn(ffc_118_n),
    .din(ffc_176_p_spl_)
  );


  DROC
  ffc_119
  (
    .doutp(ffc_119_p),
    .doutn(ffc_119_n),
    .din(ffc_177_p_spl_)
  );


  DROC
  ffc_120
  (
    .doutp(ffc_120_p),
    .doutn(ffc_120_n),
    .din(g369_n_spl_)
  );


  DROC
  ffc_121
  (
    .doutp(ffc_121_p),
    .doutn(ffc_121_n),
    .din(g378_p_spl_)
  );


  DROC
  ffc_122
  (
    .doutp(ffc_122_p),
    .doutn(ffc_122_n),
    .din(g387_p_spl_)
  );


  DROC
  ffc_123
  (
    .doutp(ffc_123_p),
    .doutn(ffc_123_n),
    .din(ffc_13_p_spl_)
  );


  DROC
  ffc_124
  (
    .doutp(ffc_124_p),
    .doutn(ffc_124_n),
    .din(ffc_19_p_spl_)
  );


  DROC
  ffc_125
  (
    .doutp(ffc_125_p),
    .doutn(ffc_125_n),
    .din(ffc_41_p)
  );


  DROC
  ffc_126
  (
    .doutp(ffc_126_p),
    .doutn(ffc_126_n),
    .din(g388_p)
  );


  DROC
  ffc_127
  (
    .doutp(ffc_127_p),
    .doutn(ffc_127_n),
    .din(g389_p)
  );


  DROC
  ffc_128
  (
    .doutp(ffc_128_p),
    .doutn(ffc_128_n),
    .din(g390_p_spl_)
  );


  DROC
  ffc_129
  (
    .doutp(ffc_129_p),
    .doutn(ffc_129_n),
    .din(g395_p)
  );


  DROC
  ffc_130
  (
    .doutp(ffc_130_p),
    .doutn(ffc_130_n),
    .din(g397_p)
  );


  DROC
  ffc_131
  (
    .doutp(ffc_131_p),
    .doutn(ffc_131_n),
    .din(g398_p)
  );


  DROC
  ffc_132
  (
    .doutp(ffc_132_p),
    .doutn(ffc_132_n),
    .din(g409_n_spl_)
  );


  DROC
  ffc_133
  (
    .doutp(ffc_133_n),
    .doutn(ffc_133_p),
    .din(g419_n_spl_)
  );


  DROC
  ffc_134
  (
    .doutp(ffc_134_p),
    .doutn(ffc_134_n),
    .din(ffc_0_p_spl_)
  );


  DROC
  ffc_135
  (
    .doutp(ffc_135_p),
    .doutn(ffc_135_n),
    .din(ffc_4_p_spl_)
  );


  DROC
  ffc_136
  (
    .doutp(ffc_136_p),
    .doutn(ffc_136_n),
    .din(ffc_6_p_spl_)
  );


  DROC
  ffc_137
  (
    .doutp(ffc_137_p),
    .doutn(ffc_137_n),
    .din(ffc_23_p_spl_)
  );


  DROC
  ffc_138
  (
    .doutp(ffc_138_p),
    .doutn(ffc_138_n),
    .din(ffc_29_p)
  );


  DROC
  ffc_139
  (
    .doutp(ffc_139_p),
    .doutn(ffc_139_n),
    .din(g422_p_spl_)
  );


  DROC
  ffc_140
  (
    .doutp(ffc_140_p),
    .doutn(ffc_140_n),
    .din(ffc_35_p)
  );


  DROC
  ffc_141
  (
    .doutp(ffc_141_p),
    .doutn(ffc_141_n),
    .din(ffc_38_p)
  );


  DROC
  ffc_142
  (
    .doutp(ffc_142_p),
    .doutn(ffc_142_n),
    .din(g423_n)
  );


  DROC
  ffc_143
  (
    .doutp(ffc_143_p),
    .doutn(ffc_143_n),
    .din(g424_p)
  );


  DROC
  ffc_144
  (
    .doutp(ffc_144_n),
    .doutn(ffc_144_p),
    .din(g425_p)
  );


  DROC
  ffc_145
  (
    .doutp(ffc_145_p),
    .doutn(ffc_145_n),
    .din(ffc_21_p_spl_)
  );


  DROC
  ffc_146
  (
    .doutp(ffc_146_p),
    .doutn(ffc_146_n),
    .din(g427_p)
  );


  DROC
  ffc_147
  (
    .doutp(ffc_147_n),
    .doutn(ffc_147_p),
    .din(g428_n)
  );


  DROC
  ffc_148
  (
    .doutp(ffc_148_p),
    .doutn(ffc_148_n),
    .din(g430_n)
  );


  DROC
  ffc_149
  (
    .doutp(ffc_149_p),
    .doutn(ffc_149_n),
    .din(g431_p)
  );


  DROC
  ffc_150
  (
    .doutp(ffc_150_p),
    .doutn(ffc_150_n),
    .din(g442_p)
  );


  DROC
  ffc_151
  (
    .doutp(ffc_151_n),
    .doutn(ffc_151_p),
    .din(g443_n)
  );


  DROC
  ffc_152
  (
    .doutp(ffc_152_p),
    .doutn(ffc_152_n),
    .din(g453_n)
  );


  DROC
  ffc_153
  (
    .doutp(ffc_153_n),
    .doutn(ffc_153_p),
    .din(g459_n_spl_)
  );


  DROC
  ffc_154
  (
    .doutp(ffc_154_p),
    .doutn(ffc_154_n),
    .din(ffc_24_p)
  );


  DROC
  ffc_155
  (
    .doutp(ffc_155_p),
    .doutn(ffc_155_n),
    .din(g460_p)
  );


  DROC
  ffc_156
  (
    .doutp(ffc_156_p),
    .doutn(ffc_156_n),
    .din(g461_p)
  );


  DROC
  ffc_157
  (
    .doutp(ffc_157_p),
    .doutn(ffc_157_n),
    .din(g462_p)
  );


  DROC
  ffc_158
  (
    .doutp(ffc_158_p),
    .doutn(ffc_158_n),
    .din(g464_p)
  );


  DROC
  ffc_159
  (
    .doutp(ffc_159_p),
    .doutn(ffc_159_n),
    .din(g470_p)
  );


  DROC
  ffc_160
  (
    .doutp(ffc_160_n),
    .doutn(ffc_160_p),
    .din(g471_n)
  );


  DROC
  ffc_161
  (
    .doutp(ffc_161_p),
    .doutn(ffc_161_n),
    .din(ffc_22_p)
  );


  DROC
  ffc_162
  (
    .doutp(ffc_162_p),
    .doutn(ffc_162_n),
    .din(g474_n)
  );


  DROC
  ffc_163
  (
    .doutp(ffc_163_p),
    .doutn(ffc_163_n),
    .din(g480_n)
  );


  DROC
  ffc_164
  (
    .doutp(ffc_164_p),
    .doutn(ffc_164_n),
    .din(g483_n)
  );


  DROC
  ffc_165
  (
    .doutp(ffc_165_p),
    .doutn(ffc_165_n),
    .din(g489_n)
  );


  DROC
  ffc_166
  (
    .doutp(ffc_166_p),
    .doutn(ffc_166_n),
    .din(g495_n)
  );


  DROC
  ffc_167
  (
    .doutp(ffc_167_p),
    .doutn(ffc_167_n),
    .din(g501_n)
  );


  DROC
  ffc_168
  (
    .doutp(ffc_168_p),
    .doutn(ffc_168_n),
    .din(g508_p)
  );


  DROC
  ffc_169
  (
    .doutp(ffc_169_n),
    .doutn(ffc_169_p),
    .din(g509_n)
  );


  DROC
  ffc_170
  (
    .doutp(ffc_170_p),
    .doutn(ffc_170_n),
    .din(G2_p)
  );


  DROC
  ffc_171
  (
    .doutp(ffc_171_p),
    .doutn(ffc_171_n),
    .din(G3_p)
  );


  DROC
  ffc_172
  (
    .doutp(ffc_172_p),
    .doutn(ffc_172_n),
    .din(G6_p)
  );


  DROC
  ffc_173
  (
    .doutp(ffc_173_p),
    .doutn(ffc_173_n),
    .din(G7_p)
  );


  DROC
  ffc_174
  (
    .doutp(ffc_174_p),
    .doutn(ffc_174_n),
    .din(G8_p)
  );


  DROC
  ffc_175
  (
    .doutp(ffc_175_p),
    .doutn(ffc_175_n),
    .din(G9_p)
  );


  DROC
  ffc_176
  (
    .doutp(ffc_176_p),
    .doutn(ffc_176_n),
    .din(G14_p)
  );


  DROC
  ffc_177
  (
    .doutp(ffc_177_p),
    .doutn(ffc_177_n),
    .din(G33_p)
  );


  DROC
  ffc_178
  (
    .doutp(ffc_178_p),
    .doutn(ffc_178_n),
    .din(G10_p)
  );


  DROC
  ffc_179
  (
    .doutp(ffc_179_p),
    .doutn(ffc_179_n),
    .din(G12_p)
  );


  DROC
  ffc_180
  (
    .doutp(ffc_180_p),
    .doutn(ffc_180_n),
    .din(G13_p)
  );


  DROC
  ffc_181
  (
    .doutp(ffc_181_p),
    .doutn(ffc_181_n),
    .din(G15_p)
  );


  DROC
  ffc_182
  (
    .doutp(ffc_182_p),
    .doutn(ffc_182_n),
    .din(G18_p)
  );


  DROC
  ffc_183
  (
    .doutp(ffc_183_p),
    .doutn(ffc_183_n),
    .din(G24_p)
  );


  buf

  (
    ffc_129_n_spl_,
    ffc_129_n
  );


  buf

  (
    ffc_131_p_spl_,
    ffc_131_p
  );


  buf

  (
    ffc_129_p_spl_,
    ffc_129_p
  );


  buf

  (
    ffc_131_n_spl_,
    ffc_131_n
  );


  buf

  (
    g218_n_spl_,
    g218_n
  );


  buf

  (
    g218_n_spl_0,
    g218_n_spl_
  );


  buf

  (
    g218_n_spl_00,
    g218_n_spl_0
  );


  buf

  (
    g218_n_spl_01,
    g218_n_spl_0
  );


  buf

  (
    g218_n_spl_1,
    g218_n_spl_
  );


  buf

  (
    g218_n_spl_10,
    g218_n_spl_1
  );


  buf

  (
    g218_p_spl_,
    g218_p
  );


  buf

  (
    g218_p_spl_0,
    g218_p_spl_
  );


  buf

  (
    g218_p_spl_00,
    g218_p_spl_0
  );


  buf

  (
    g218_p_spl_01,
    g218_p_spl_0
  );


  buf

  (
    g218_p_spl_1,
    g218_p_spl_
  );


  buf

  (
    g218_p_spl_10,
    g218_p_spl_1
  );


  buf

  (
    ffc_130_n_spl_,
    ffc_130_n
  );


  buf

  (
    ffc_130_n_spl_0,
    ffc_130_n_spl_
  );


  buf

  (
    ffc_130_p_spl_,
    ffc_130_p
  );


  buf

  (
    ffc_130_p_spl_0,
    ffc_130_p_spl_
  );


  buf

  (
    g231_n_spl_,
    g231_n
  );


  buf

  (
    g231_n_spl_0,
    g231_n_spl_
  );


  buf

  (
    g231_n_spl_00,
    g231_n_spl_0
  );


  buf

  (
    g231_n_spl_01,
    g231_n_spl_0
  );


  buf

  (
    g231_n_spl_1,
    g231_n_spl_
  );


  buf

  (
    g231_p_spl_,
    g231_p
  );


  buf

  (
    g231_p_spl_0,
    g231_p_spl_
  );


  buf

  (
    g231_p_spl_00,
    g231_p_spl_0
  );


  buf

  (
    g231_p_spl_01,
    g231_p_spl_0
  );


  buf

  (
    g231_p_spl_1,
    g231_p_spl_
  );


  buf

  (
    ffc_98_n_spl_,
    ffc_98_n
  );


  buf

  (
    ffc_93_n_spl_,
    ffc_93_n
  );


  buf

  (
    g242_p_spl_,
    g242_p
  );


  buf

  (
    g242_n_spl_,
    g242_n
  );


  buf

  (
    g243_n_spl_,
    g243_n
  );


  buf

  (
    g243_n_spl_0,
    g243_n_spl_
  );


  buf

  (
    g243_n_spl_1,
    g243_n_spl_
  );


  buf

  (
    g243_p_spl_,
    g243_p
  );


  buf

  (
    g243_p_spl_0,
    g243_p_spl_
  );


  buf

  (
    g243_p_spl_1,
    g243_p_spl_
  );


  buf

  (
    ffc_91_n_spl_,
    ffc_91_n
  );


  buf

  (
    ffc_92_p_spl_,
    ffc_92_p
  );


  buf

  (
    ffc_99_p_spl_,
    ffc_99_p
  );


  buf

  (
    g263_n_spl_,
    g263_n
  );


  buf

  (
    g263_n_spl_0,
    g263_n_spl_
  );


  buf

  (
    g263_n_spl_1,
    g263_n_spl_
  );


  buf

  (
    g263_p_spl_,
    g263_p
  );


  buf

  (
    g263_p_spl_0,
    g263_p_spl_
  );


  buf

  (
    g263_p_spl_1,
    g263_p_spl_
  );


  buf

  (
    g276_n_spl_,
    g276_n
  );


  buf

  (
    g276_n_spl_0,
    g276_n_spl_
  );


  buf

  (
    g276_n_spl_00,
    g276_n_spl_0
  );


  buf

  (
    g276_n_spl_01,
    g276_n_spl_0
  );


  buf

  (
    g276_n_spl_1,
    g276_n_spl_
  );


  buf

  (
    ffc_58_p_spl_,
    ffc_58_p
  );


  buf

  (
    ffc_58_p_spl_0,
    ffc_58_p_spl_
  );


  buf

  (
    ffc_53_n_spl_,
    ffc_53_n
  );


  buf

  (
    ffc_53_n_spl_0,
    ffc_53_n_spl_
  );


  buf

  (
    ffc_53_n_spl_00,
    ffc_53_n_spl_0
  );


  buf

  (
    ffc_53_n_spl_1,
    ffc_53_n_spl_
  );


  buf

  (
    ffc_53_p_spl_,
    ffc_53_p
  );


  buf

  (
    ffc_53_p_spl_0,
    ffc_53_p_spl_
  );


  buf

  (
    g276_p_spl_,
    g276_p
  );


  buf

  (
    g276_p_spl_0,
    g276_p_spl_
  );


  buf

  (
    ffc_97_p_spl_,
    ffc_97_p
  );


  buf

  (
    ffc_97_p_spl_0,
    ffc_97_p_spl_
  );


  buf

  (
    ffc_97_p_spl_00,
    ffc_97_p_spl_0
  );


  buf

  (
    ffc_97_p_spl_01,
    ffc_97_p_spl_0
  );


  buf

  (
    ffc_97_p_spl_1,
    ffc_97_p_spl_
  );


  buf

  (
    ffc_58_n_spl_,
    ffc_58_n
  );


  buf

  (
    g310_n_spl_,
    g310_n
  );


  buf

  (
    g310_p_spl_,
    g310_p
  );


  buf

  (
    g320_n_spl_,
    g320_n
  );


  buf

  (
    g320_p_spl_,
    g320_p
  );


  buf

  (
    ffc_142_n_spl_,
    ffc_142_n
  );


  buf

  (
    ffc_102_n_spl_,
    ffc_102_n
  );


  buf

  (
    ffc_102_p_spl_,
    ffc_102_p
  );


  buf

  (
    ffc_102_p_spl_0,
    ffc_102_p_spl_
  );


  buf

  (
    ffc_102_p_spl_1,
    ffc_102_p_spl_
  );


  buf

  (
    ffc_152_p_spl_,
    ffc_152_p
  );


  buf

  (
    g331_p_spl_,
    g331_p
  );


  buf

  (
    ffc_45_p_spl_,
    ffc_45_p
  );


  buf

  (
    ffc_81_p_spl_,
    ffc_81_p
  );


  buf

  (
    ffc_81_p_spl_0,
    ffc_81_p_spl_
  );


  buf

  (
    ffc_81_p_spl_1,
    ffc_81_p_spl_
  );


  buf

  (
    ffc_49_p_spl_,
    ffc_49_p
  );


  buf

  (
    ffc_56_p_spl_,
    ffc_56_p
  );


  buf

  (
    g332_n_spl_,
    g332_n
  );


  buf

  (
    ffc_32_p_spl_,
    ffc_32_p
  );


  buf

  (
    ffc_141_p_spl_,
    ffc_141_p
  );


  buf

  (
    ffc_140_p_spl_,
    ffc_140_p
  );


  buf

  (
    g338_n_spl_,
    g338_n
  );


  buf

  (
    g345_p_spl_,
    g345_p
  );


  buf

  (
    g333_n_spl_,
    g333_n
  );


  buf

  (
    g337_p_spl_,
    g337_p
  );


  buf

  (
    g356_p_spl_,
    g356_p
  );


  buf

  (
    ffc_52_p_spl_,
    ffc_52_p
  );


  buf

  (
    ffc_52_p_spl_0,
    ffc_52_p_spl_
  );


  buf

  (
    ffc_52_p_spl_1,
    ffc_52_p_spl_
  );


  buf

  (
    ffc_138_p_spl_,
    ffc_138_p
  );


  buf

  (
    ffc_138_p_spl_0,
    ffc_138_p_spl_
  );


  buf

  (
    ffc_162_n_spl_,
    ffc_162_n
  );


  buf

  (
    ffc_163_p_spl_,
    ffc_163_p
  );


  buf

  (
    ffc_162_p_spl_,
    ffc_162_p
  );


  buf

  (
    ffc_163_n_spl_,
    ffc_163_n
  );


  buf

  (
    ffc_161_p_spl_,
    ffc_161_p
  );


  buf

  (
    ffc_119_n_spl_,
    ffc_119_n
  );


  buf

  (
    ffc_119_n_spl_0,
    ffc_119_n_spl_
  );


  buf

  (
    ffc_119_n_spl_1,
    ffc_119_n_spl_
  );


  buf

  (
    ffc_119_p_spl_,
    ffc_119_p
  );


  buf

  (
    ffc_119_p_spl_0,
    ffc_119_p_spl_
  );


  buf

  (
    ffc_119_p_spl_00,
    ffc_119_p_spl_0
  );


  buf

  (
    ffc_119_p_spl_1,
    ffc_119_p_spl_
  );


  buf

  (
    ffc_164_n_spl_,
    ffc_164_n
  );


  buf

  (
    ffc_164_n_spl_0,
    ffc_164_n_spl_
  );


  buf

  (
    ffc_164_n_spl_1,
    ffc_164_n_spl_
  );


  buf

  (
    ffc_166_p_spl_,
    ffc_166_p
  );


  buf

  (
    ffc_164_p_spl_,
    ffc_164_p
  );


  buf

  (
    ffc_164_p_spl_0,
    ffc_164_p_spl_
  );


  buf

  (
    ffc_164_p_spl_1,
    ffc_164_p_spl_
  );


  buf

  (
    ffc_166_n_spl_,
    ffc_166_n
  );


  buf

  (
    ffc_107_n_spl_,
    ffc_107_n
  );


  buf

  (
    ffc_158_p_spl_,
    ffc_158_p
  );


  buf

  (
    ffc_107_p_spl_,
    ffc_107_p
  );


  buf

  (
    ffc_107_p_spl_0,
    ffc_107_p_spl_
  );


  buf

  (
    ffc_158_n_spl_,
    ffc_158_n
  );


  buf

  (
    ffc_165_p_spl_,
    ffc_165_p
  );


  buf

  (
    ffc_165_p_spl_0,
    ffc_165_p_spl_
  );


  buf

  (
    ffc_167_p_spl_,
    ffc_167_p
  );


  buf

  (
    ffc_167_p_spl_0,
    ffc_167_p_spl_
  );


  buf

  (
    ffc_167_p_spl_1,
    ffc_167_p_spl_
  );


  buf

  (
    ffc_165_n_spl_,
    ffc_165_n
  );


  buf

  (
    ffc_165_n_spl_0,
    ffc_165_n_spl_
  );


  buf

  (
    ffc_167_n_spl_,
    ffc_167_n
  );


  buf

  (
    ffc_167_n_spl_0,
    ffc_167_n_spl_
  );


  buf

  (
    ffc_167_n_spl_1,
    ffc_167_n_spl_
  );


  buf

  (
    ffc_116_n_spl_,
    ffc_116_n
  );


  buf

  (
    ffc_135_p_spl_,
    ffc_135_p
  );


  buf

  (
    ffc_135_p_spl_0,
    ffc_135_p_spl_
  );


  buf

  (
    ffc_135_p_spl_00,
    ffc_135_p_spl_0
  );


  buf

  (
    ffc_135_p_spl_1,
    ffc_135_p_spl_
  );


  buf

  (
    ffc_116_p_spl_,
    ffc_116_p
  );


  buf

  (
    ffc_116_p_spl_0,
    ffc_116_p_spl_
  );


  buf

  (
    ffc_135_n_spl_,
    ffc_135_n
  );


  buf

  (
    ffc_135_n_spl_0,
    ffc_135_n_spl_
  );


  buf

  (
    ffc_135_n_spl_1,
    ffc_135_n_spl_
  );


  buf

  (
    g381_n_spl_,
    g381_n
  );


  buf

  (
    g384_p_spl_,
    g384_p
  );


  buf

  (
    g381_p_spl_,
    g381_p
  );


  buf

  (
    g384_n_spl_,
    g384_n
  );


  buf

  (
    g361_n_spl_,
    g361_n
  );


  buf

  (
    g391_p_spl_,
    g391_p
  );


  buf

  (
    g339_n_spl_,
    g339_n
  );


  buf

  (
    g392_n_spl_,
    g392_n
  );


  buf

  (
    g341_n_spl_,
    g341_n
  );


  buf

  (
    g394_n_spl_,
    g394_n
  );


  buf

  (
    g340_n_spl_,
    g340_n
  );


  buf

  (
    g358_n_spl_,
    g358_n
  );


  buf

  (
    g360_p_spl_,
    g360_p
  );


  buf

  (
    g399_p_spl_,
    g399_p
  );


  buf

  (
    g399_n_spl_,
    g399_n
  );


  buf

  (
    ffc_112_n_spl_,
    ffc_112_n
  );


  buf

  (
    g403_n_spl_,
    g403_n
  );


  buf

  (
    ffc_112_p_spl_,
    ffc_112_p
  );


  buf

  (
    ffc_112_p_spl_0,
    ffc_112_p_spl_
  );


  buf

  (
    g403_p_spl_,
    g403_p
  );


  buf

  (
    ffc_134_p_spl_,
    ffc_134_p
  );


  buf

  (
    ffc_134_p_spl_0,
    ffc_134_p_spl_
  );


  buf

  (
    g410_p_spl_,
    g410_p
  );


  buf

  (
    ffc_134_n_spl_,
    ffc_134_n
  );


  buf

  (
    g410_n_spl_,
    g410_n
  );


  buf

  (
    g357_p_spl_,
    g357_p
  );


  buf

  (
    g357_p_spl_0,
    g357_p_spl_
  );


  buf

  (
    g357_n_spl_,
    g357_n
  );


  buf

  (
    g357_n_spl_0,
    g357_n_spl_
  );


  buf

  (
    g357_n_spl_1,
    g357_n_spl_
  );


  buf

  (
    ffc_175_n_spl_,
    ffc_175_n
  );


  buf

  (
    ffc_176_n_spl_,
    ffc_176_n
  );


  buf

  (
    ffc_175_p_spl_,
    ffc_175_p
  );


  buf

  (
    ffc_175_p_spl_0,
    ffc_175_p_spl_
  );


  buf

  (
    ffc_176_p_spl_,
    ffc_176_p
  );


  buf

  (
    ffc_176_p_spl_0,
    ffc_176_p_spl_
  );


  buf

  (
    ffc_110_p_spl_,
    ffc_110_p
  );


  buf

  (
    ffc_52_n_spl_,
    ffc_52_n
  );


  buf

  (
    ffc_52_n_spl_0,
    ffc_52_n_spl_
  );


  buf

  (
    g409_n_spl_,
    g409_n
  );


  buf

  (
    g419_n_spl_,
    g419_n
  );


  buf

  (
    g369_n_spl_,
    g369_n
  );


  buf

  (
    ffc_41_n_spl_,
    ffc_41_n
  );


  buf

  (
    g426_p_spl_,
    g426_p
  );


  buf

  (
    g378_p_spl_,
    g378_p
  );


  buf

  (
    g390_p_spl_,
    g390_p
  );


  buf

  (
    g390_p_spl_0,
    g390_p_spl_
  );


  buf

  (
    g429_n_spl_,
    g429_n
  );


  buf

  (
    ffc_27_p_spl_,
    ffc_27_p
  );


  buf

  (
    ffc_118_n_spl_,
    ffc_118_n
  );


  buf

  (
    ffc_118_p_spl_,
    ffc_118_p
  );


  buf

  (
    ffc_118_p_spl_0,
    ffc_118_p_spl_
  );


  buf

  (
    g438_n_spl_,
    g438_n
  );


  buf

  (
    g441_p_spl_,
    g441_p
  );


  buf

  (
    ffc_154_p_spl_,
    ffc_154_p
  );


  buf

  (
    ffc_117_p_spl_,
    ffc_117_p
  );


  buf

  (
    ffc_117_p_spl_0,
    ffc_117_p_spl_
  );


  buf

  (
    ffc_153_n_spl_,
    ffc_153_n
  );


  buf

  (
    ffc_117_n_spl_,
    ffc_117_n
  );


  buf

  (
    ffc_153_p_spl_,
    ffc_153_p
  );


  buf

  (
    g444_p_spl_,
    g444_p
  );


  buf

  (
    g447_n_spl_,
    g447_n
  );


  buf

  (
    g444_n_spl_,
    g444_n
  );


  buf

  (
    g447_p_spl_,
    g447_p
  );


  buf

  (
    g387_p_spl_,
    g387_p
  );


  buf

  (
    ffc_178_p_spl_,
    ffc_178_p
  );


  buf

  (
    ffc_178_p_spl_0,
    ffc_178_p_spl_
  );


  buf

  (
    ffc_178_p_spl_00,
    ffc_178_p_spl_0
  );


  buf

  (
    ffc_178_p_spl_1,
    ffc_178_p_spl_
  );


  buf

  (
    ffc_181_n_spl_,
    ffc_181_n
  );


  buf

  (
    ffc_181_n_spl_0,
    ffc_181_n_spl_
  );


  buf

  (
    ffc_178_n_spl_,
    ffc_178_n
  );


  buf

  (
    ffc_178_n_spl_0,
    ffc_178_n_spl_
  );


  buf

  (
    ffc_178_n_spl_1,
    ffc_178_n_spl_
  );


  buf

  (
    ffc_181_p_spl_,
    ffc_181_p
  );


  buf

  (
    ffc_181_p_spl_0,
    ffc_181_p_spl_
  );


  buf

  (
    ffc_181_p_spl_1,
    ffc_181_p_spl_
  );


  buf

  (
    ffc_19_p_spl_,
    ffc_19_p
  );


  buf

  (
    ffc_19_p_spl_0,
    ffc_19_p_spl_
  );


  buf

  (
    g456_n_spl_,
    g456_n
  );


  buf

  (
    ffc_19_n_spl_,
    ffc_19_n
  );


  buf

  (
    g456_p_spl_,
    g456_p
  );


  buf

  (
    ffc_21_p_spl_,
    ffc_21_p
  );


  buf

  (
    ffc_183_n_spl_,
    ffc_183_n
  );


  buf

  (
    ffc_6_p_spl_,
    ffc_6_p
  );


  buf

  (
    ffc_6_p_spl_0,
    ffc_6_p_spl_
  );


  buf

  (
    ffc_174_n_spl_,
    ffc_174_n
  );


  buf

  (
    ffc_174_n_spl_0,
    ffc_174_n_spl_
  );


  buf

  (
    ffc_6_n_spl_,
    ffc_6_n
  );


  buf

  (
    ffc_174_p_spl_,
    ffc_174_p
  );


  buf

  (
    ffc_174_p_spl_0,
    ffc_174_p_spl_
  );


  buf

  (
    ffc_174_p_spl_1,
    ffc_174_p_spl_
  );


  buf

  (
    ffc_23_p_spl_,
    ffc_23_p
  );


  buf

  (
    ffc_177_n_spl_,
    ffc_177_n
  );


  buf

  (
    ffc_182_p_spl_,
    ffc_182_p
  );


  buf

  (
    ffc_183_p_spl_,
    ffc_183_p
  );


  buf

  (
    ffc_177_p_spl_,
    ffc_177_p
  );


  buf

  (
    ffc_13_n_spl_,
    ffc_13_n
  );


  buf

  (
    ffc_13_n_spl_0,
    ffc_13_n_spl_
  );


  buf

  (
    g469_n_spl_,
    g469_n
  );


  buf

  (
    ffc_179_n_spl_,
    ffc_179_n
  );


  buf

  (
    ffc_179_n_spl_0,
    ffc_179_n_spl_
  );


  buf

  (
    ffc_179_p_spl_,
    ffc_179_p
  );


  buf

  (
    ffc_179_p_spl_0,
    ffc_179_p_spl_
  );


  buf

  (
    ffc_179_p_spl_1,
    ffc_179_p_spl_
  );


  buf

  (
    ffc_172_p_spl_,
    ffc_172_p
  );


  buf

  (
    ffc_172_p_spl_0,
    ffc_172_p_spl_
  );


  buf

  (
    ffc_172_p_spl_00,
    ffc_172_p_spl_0
  );


  buf

  (
    ffc_172_p_spl_1,
    ffc_172_p_spl_
  );


  buf

  (
    ffc_172_n_spl_,
    ffc_172_n
  );


  buf

  (
    ffc_172_n_spl_0,
    ffc_172_n_spl_
  );


  buf

  (
    ffc_172_n_spl_1,
    ffc_172_n_spl_
  );


  buf

  (
    ffc_171_n_spl_,
    ffc_171_n
  );


  buf

  (
    ffc_171_n_spl_0,
    ffc_171_n_spl_
  );


  buf

  (
    ffc_171_p_spl_,
    ffc_171_p
  );


  buf

  (
    ffc_171_p_spl_0,
    ffc_171_p_spl_
  );


  buf

  (
    ffc_171_p_spl_1,
    ffc_171_p_spl_
  );


  buf

  (
    g422_p_spl_,
    g422_p
  );


  buf

  (
    ffc_170_n_spl_,
    ffc_170_n
  );


  buf

  (
    ffc_170_p_spl_,
    ffc_170_p
  );


  buf

  (
    ffc_170_p_spl_0,
    ffc_170_p_spl_
  );


  buf

  (
    ffc_0_p_spl_,
    ffc_0_p
  );


  buf

  (
    ffc_173_p_spl_,
    ffc_173_p
  );


  buf

  (
    ffc_173_p_spl_0,
    ffc_173_p_spl_
  );


  buf

  (
    ffc_173_p_spl_00,
    ffc_173_p_spl_0
  );


  buf

  (
    ffc_173_p_spl_1,
    ffc_173_p_spl_
  );


  buf

  (
    ffc_173_n_spl_,
    ffc_173_n
  );


  buf

  (
    ffc_173_n_spl_0,
    ffc_173_n_spl_
  );


  buf

  (
    ffc_173_n_spl_1,
    ffc_173_n_spl_
  );


  buf

  (
    ffc_4_p_spl_,
    ffc_4_p
  );


  buf

  (
    ffc_180_n_spl_,
    ffc_180_n
  );


  buf

  (
    ffc_180_p_spl_,
    ffc_180_p
  );


  buf

  (
    ffc_180_p_spl_0,
    ffc_180_p_spl_
  );


  buf

  (
    ffc_13_p_spl_,
    ffc_13_p
  );


  buf

  (
    g459_n_spl_,
    g459_n
  );


  buf

  (
    g459_n_spl_0,
    g459_n_spl_
  );


  buf

  (
    g507_n_spl_,
    g507_n
  );


endmodule
