
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  G42,
  G43,
  G44,
  G45,
  G46,
  G47,
  G48,
  G49,
  G50,
  G51,
  G52,
  G53,
  G54,
  G55,
  G56,
  G57,
  G58,
  G59,
  G60,
  G61,
  G62,
  G63,
  G64,
  G65,
  G66,
  G67,
  G68,
  G69,
  G70,
  G71,
  G72,
  G73,
  G74,
  G75,
  G76,
  G77,
  G78,
  G79,
  G80,
  G81,
  G82,
  G83,
  G84,
  G85,
  G86,
  G87,
  G88,
  G89,
  G90,
  G91,
  G92,
  G93,
  G94,
  G95,
  G96,
  G97,
  G98,
  G99,
  G100,
  G101,
  G102,
  G103,
  G104,
  G105,
  G106,
  G107,
  G108,
  G109,
  G110,
  G111,
  G112,
  G113,
  G114,
  G115,
  G116,
  G117,
  G118,
  G119,
  G120,
  G121,
  G122,
  G123,
  G124,
  G125,
  G126,
  G127,
  G128,
  G129,
  G130,
  G131,
  G132,
  G133,
  G134,
  G135,
  G136,
  G137,
  G138,
  G139,
  G140,
  G141,
  G142,
  G143,
  G144,
  G145,
  G146,
  G147,
  G148,
  G149,
  G150,
  G151,
  G152,
  G153,
  G154,
  G155,
  G156,
  G157,
  G158,
  G159,
  G160,
  G161,
  G162,
  G163,
  G164,
  G165,
  G166,
  G167,
  G168,
  G169,
  G170,
  G171,
  G172,
  G173,
  G174,
  G175,
  G176,
  G177,
  G178,
  n2610_lo,
  n2613_lo,
  n2616_lo,
  n2619_lo,
  n2622_lo,
  n2625_lo,
  n2628_lo,
  n2634_lo,
  n2637_lo,
  n2640_lo,
  n2643_lo,
  n2646_lo,
  n2649_lo,
  n2652_lo,
  n2655_lo,
  n2658_lo,
  n2661_lo,
  n2664_lo,
  n2667_lo,
  n2670_lo,
  n2673_lo,
  n2676_lo,
  n2679_lo,
  n2682_lo,
  n2685_lo,
  n2688_lo,
  n2691_lo,
  n2694_lo,
  n2697_lo,
  n2700_lo,
  n2703_lo,
  n2706_lo,
  n2709_lo,
  n2712_lo,
  n2715_lo,
  n2718_lo,
  n2721_lo,
  n2724_lo,
  n2727_lo,
  n2730_lo,
  n2733_lo,
  n2736_lo,
  n2739_lo,
  n2742_lo,
  n2745_lo,
  n2748_lo,
  n2751_lo,
  n2754_lo,
  n2757_lo,
  n2760_lo,
  n2763_lo,
  n2766_lo,
  n2769_lo,
  n2772_lo,
  n2775_lo,
  n2778_lo,
  n2781_lo,
  n2784_lo,
  n2787_lo,
  n2790_lo,
  n2793_lo,
  n2796_lo,
  n2799_lo,
  n2802_lo,
  n2805_lo,
  n2808_lo,
  n2811_lo,
  n2814_lo,
  n2817_lo,
  n2820_lo,
  n2823_lo,
  n2826_lo,
  n2829_lo,
  n2832_lo,
  n2838_lo,
  n2841_lo,
  n2844_lo,
  n2847_lo,
  n2850_lo,
  n2853_lo,
  n2856_lo,
  n2862_lo,
  n2865_lo,
  n2868_lo,
  n2871_lo,
  n2874_lo,
  n2877_lo,
  n2880_lo,
  n2883_lo,
  n2886_lo,
  n2889_lo,
  n2892_lo,
  n2895_lo,
  n2898_lo,
  n2901_lo,
  n2904_lo,
  n2907_lo,
  n2910_lo,
  n2913_lo,
  n2916_lo,
  n2919_lo,
  n2922_lo,
  n2925_lo,
  n2928_lo,
  n2931_lo,
  n2934_lo,
  n2937_lo,
  n2940_lo,
  n2943_lo,
  n2946_lo,
  n2949_lo,
  n2952_lo,
  n2955_lo,
  n2958_lo,
  n2961_lo,
  n2964_lo,
  n2967_lo,
  n2970_lo,
  n2973_lo,
  n2976_lo,
  n2979_lo,
  n2982_lo,
  n2985_lo,
  n2988_lo,
  n2991_lo,
  n2994_lo,
  n2997_lo,
  n3000_lo,
  n3003_lo,
  n3006_lo,
  n3009_lo,
  n3012_lo,
  n3015_lo,
  n3018_lo,
  n3021_lo,
  n3024_lo,
  n3027_lo,
  n3030_lo,
  n3033_lo,
  n3036_lo,
  n3039_lo,
  n3042_lo,
  n3045_lo,
  n3048_lo,
  n3051_lo,
  n3054_lo,
  n3057_lo,
  n3060_lo,
  n3063_lo,
  n3066_lo,
  n3069_lo,
  n3072_lo,
  n3075_lo,
  n3078_lo,
  n3081_lo,
  n3084_lo,
  n3087_lo,
  n3090_lo,
  n3093_lo,
  n3096_lo,
  n3099_lo,
  n3102_lo,
  n3105_lo,
  n3108_lo,
  n3111_lo,
  n3114_lo,
  n3117_lo,
  n3120_lo,
  n3126_lo,
  n3129_lo,
  n3132_lo,
  n3138_lo,
  n3141_lo,
  n3144_lo,
  n3147_lo,
  n3150_lo,
  n3153_lo,
  n3156_lo,
  n3162_lo,
  n3165_lo,
  n3168_lo,
  n3174_lo,
  n3177_lo,
  n3180_lo,
  n3186_lo,
  n3189_lo,
  n3192_lo,
  n3195_lo,
  n3198_lo,
  n3201_lo,
  n3204_lo,
  n3210_lo,
  n3213_lo,
  n3216_lo,
  n3219_lo,
  n3222_lo,
  n3225_lo,
  n3228_lo,
  n3234_lo,
  n3237_lo,
  n3240_lo,
  n3243_lo,
  n3246_lo,
  n3249_lo,
  n3252_lo,
  n3255_lo,
  n3258_lo,
  n3261_lo,
  n3264_lo,
  n3267_lo,
  n3270_lo,
  n3273_lo,
  n3276_lo,
  n3279_lo,
  n3282_lo,
  n3285_lo,
  n3288_lo,
  n3294_lo,
  n3297_lo,
  n3300_lo,
  n3306_lo,
  n3309_lo,
  n3312_lo,
  n3318_lo,
  n3321_lo,
  n3324_lo,
  n3330_lo,
  n3333_lo,
  n3336_lo,
  n3339_lo,
  n3342_lo,
  n3345_lo,
  n3348_lo,
  n3351_lo,
  n3354_lo,
  n3357_lo,
  n3360_lo,
  n3363_lo,
  n3366_lo,
  n3369_lo,
  n3372_lo,
  n3375_lo,
  n3378_lo,
  n3381_lo,
  n3384_lo,
  n3387_lo,
  n3390_lo,
  n3393_lo,
  n3396_lo,
  n3399_lo,
  n3402_lo,
  n3405_lo,
  n3408_lo,
  n3411_lo,
  n3414_lo,
  n3417_lo,
  n3420_lo,
  n3423_lo,
  n3426_lo,
  n3429_lo,
  n3432_lo,
  n3435_lo,
  n3438_lo,
  n3441_lo,
  n3444_lo,
  n3447_lo,
  n3450_lo,
  n3453_lo,
  n3456_lo,
  n3459_lo,
  n3462_lo,
  n3465_lo,
  n3468_lo,
  n3471_lo,
  n3474_lo,
  n3477_lo,
  n3480_lo,
  n3483_lo,
  n3486_lo,
  n3489_lo,
  n3492_lo,
  n3495_lo,
  n3498_lo,
  n3501_lo,
  n3504_lo,
  n3507_lo,
  n3510_lo,
  n3513_lo,
  n3516_lo,
  n3519_lo,
  n3522_lo,
  n3525_lo,
  n3528_lo,
  n3531_lo,
  n3534_lo,
  n3537_lo,
  n3540_lo,
  n3543_lo,
  n3546_lo,
  n3549_lo,
  n3552_lo,
  n3555_lo,
  n3558_lo,
  n3561_lo,
  n3564_lo,
  n3567_lo,
  n3570_lo,
  n3573_lo,
  n3576_lo,
  n3579_lo,
  n3582_lo,
  n3585_lo,
  n3588_lo,
  n3591_lo,
  n3594_lo,
  n3597_lo,
  n3600_lo,
  n3603_lo,
  n3606_lo,
  n3609_lo,
  n3612_lo,
  n3615_lo,
  n3618_lo,
  n3621_lo,
  n3624_lo,
  n3627_lo,
  n3630_lo,
  n3633_lo,
  n3636_lo,
  n3639_lo,
  n3642_lo,
  n3645_lo,
  n3648_lo,
  n3651_lo,
  n3654_lo,
  n3666_lo,
  n3750_lo,
  n3762_lo,
  n3774_lo,
  n3786_lo,
  n3789_lo,
  n3792_lo,
  n3795_lo,
  n3798_lo,
  n3810_lo,
  n3822_lo,
  n3834_lo,
  n3846_lo,
  n3930_lo,
  n3933_lo,
  n3936_lo,
  n3942_lo,
  n3945_lo,
  n3948_lo,
  n3954_lo,
  n3957_lo,
  n3963_lo,
  n3966_lo,
  n3969_lo,
  n3975_lo,
  n3978_lo,
  n3990_lo,
  n4050_lo,
  n4062_lo,
  n4098_lo,
  n4107_lo,
  n4110_lo,
  n4122_lo,
  n4131_lo,
  n4155_lo,
  n4158_lo,
  n4170_lo,
  n4179_lo,
  n4182_lo,
  n4185_lo,
  n4188_lo,
  n4194_lo,
  n4197_lo,
  n4200_lo,
  n4206_lo,
  n4209_lo,
  n4212_lo,
  n4215_lo,
  n4230_lo,
  n4233_lo,
  n4236_lo,
  n4239_lo,
  n4242_lo,
  n4254_lo,
  n4290_lo,
  n4293_lo,
  n4302_lo,
  n4314_lo,
  n4350_lo,
  n4362_lo,
  n4374_lo,
  n4386_lo,
  n4398_lo,
  n4410_lo,
  n4413_lo,
  n4416_lo,
  n4419_lo,
  n4422_lo,
  n4425_lo,
  n4428_lo,
  n4431_lo,
  n4434_lo,
  n4437_lo,
  n4440_lo,
  n4443_lo,
  n4446_lo,
  n4449_lo,
  n4452_lo,
  n4455_lo,
  n4458_lo,
  n4461_lo,
  n4464_lo,
  n4467_lo,
  n4470_lo,
  n4473_lo,
  n4476_lo,
  n4479_lo,
  n4482_lo,
  n4485_lo,
  n4488_lo,
  n4494_lo,
  n4497_lo,
  n4500_lo,
  n4503_lo,
  n4506_lo,
  n4509_lo,
  n4512_lo,
  n4515_lo,
  n4518_lo,
  n4521_lo,
  n4524_lo,
  n4527_lo,
  n4530_lo,
  n4533_lo,
  n4536_lo,
  n4539_lo,
  n4542_lo,
  n4545_lo,
  n4554_lo,
  n4557_lo,
  n4560_lo,
  n4563_lo,
  n4566_lo,
  n4569_lo,
  n4572_lo,
  n4575_lo,
  n4578_lo,
  n4581_lo,
  n4584_lo,
  n4587_lo,
  n4590_lo,
  n4593_lo,
  n4596_lo,
  n4602_lo,
  n4605_lo,
  n4608_lo,
  n4614_lo,
  n4617_lo,
  n4620_lo,
  n4626_lo,
  n4629_lo,
  n4632_lo,
  n4638_lo,
  n4641_lo,
  n4644_lo,
  n4647_lo,
  n4650_lo,
  n4653_lo,
  n4656_lo,
  n4659_lo,
  n4662_lo,
  n4665_lo,
  n4668_lo,
  n4671_lo,
  n4674_lo,
  n4677_lo,
  n4680_lo,
  n4683_lo,
  n4686_lo,
  n4689_lo,
  n4692_lo,
  n4695_lo,
  n4698_lo,
  n4701_lo,
  n4704_lo,
  n4707_lo,
  n4710_lo,
  n4713_lo,
  n4716_lo,
  n4719_lo,
  n4722_lo,
  n4725_lo,
  n4728_lo,
  n4731_lo,
  n4734_lo,
  n4737_lo,
  n4740_lo,
  n4743_lo,
  n4970_o2,
  n4972_o2,
  n4989_o2,
  n5024_o2,
  n5025_o2,
  n5029_o2,
  n5042_o2,
  n5048_o2,
  n5093_o2,
  n5096_o2,
  n5193_o2,
  n5199_o2,
  n5203_o2,
  n5214_o2,
  n5221_o2,
  n5222_o2,
  n5273_o2,
  n5365_o2,
  n5385_o2,
  n5553_o2,
  n5636_o2,
  n5782_o2,
  n5778_o2,
  n5323_o2,
  n5325_o2,
  n5327_o2,
  n5329_o2,
  n5816_o2,
  n5817_o2,
  n5837_o2,
  n5844_o2,
  n5859_o2,
  n5857_o2,
  n5369_o2,
  n5371_o2,
  n5373_o2,
  n5400_o2,
  n5402_o2,
  n5404_o2,
  n5406_o2,
  n5407_o2,
  n5408_o2,
  n2722_o2,
  n1942_inv,
  n5412_o2,
  n1948_inv,
  n5557_o2,
  n5558_o2,
  n5559_o2,
  n5564_o2,
  n5565_o2,
  n1966_inv,
  n5568_o2,
  n5598_o2,
  n5600_o2,
  n5601_o2,
  n5602_o2,
  n5603_o2,
  n2853_o2,
  n5637_o2,
  n1993_inv,
  n1996_inv,
  n5635_o2,
  n5640_o2,
  n5641_o2,
  n5642_o2,
  n5650_o2,
  n5652_o2,
  n5653_o2,
  n5654_o2,
  n5655_o2,
  n5657_o2,
  n2029_inv,
  n5661_o2,
  n5656_o2,
  n5663_o2,
  n2041_inv,
  n5795_o2,
  n5796_o2,
  n5797_o2,
  n5739_o2,
  n5773_o2,
  n2059_inv,
  n5799_o2,
  n5802_o2,
  n2068_inv,
  n5831_o2,
  n5833_o2,
  n5820_o2,
  n5823_o2,
  n5824_o2,
  n5869_o2,
  n5848_o2,
  n5849_o2,
  n5856_o2,
  n5896_o2,
  n2754_o2,
  n2908_o2,
  n5892_o2,
  n5915_o2,
  n5919_o2,
  n5918_o2,
  n5920_o2,
  n5917_o2,
  lo586_buf_o2,
  n2818_o2,
  n2863_o2,
  n2134_inv,
  n2725_o2,
  n3016_o2,
  n3013_o2,
  n2655_o2,
  n2149_inv,
  lo562_buf_o2,
  n2155_inv,
  n2531_o2,
  n2700_o2,
  n5908_o2,
  n5910_o2,
  n5912_o2,
  n5914_o2,
  n2753_o2,
  n2878_o2,
  n2182_inv,
  n5934_o2,
  n5936_o2,
  n5938_o2,
  n2728_o2,
  lo358_buf_o2,
  lo418_buf_o2,
  lo474_buf_o2,
  lo554_buf_o2,
  lo558_buf_o2,
  lo574_buf_o2,
  n2215_inv,
  n2218_inv,
  n2221_inv,
  lo450_buf_o2,
  n2910_o2,
  n2683_o2,
  n2828_o2,
  n2582_o2,
  n2600_o2,
  n2542_o2,
  n2703_o2,
  lo510_buf_o2,
  lo514_buf_o2,
  lo538_buf_o2,
  lo578_buf_o2,
  n2260_inv,
  n2666_o2,
  n2667_o2,
  n2660_o2,
  n2272_inv,
  lo454_buf_o2,
  n3593_o2,
  n3048_o2,
  lo410_buf_o2,
  lo502_buf_o2,
  lo506_buf_o2,
  lo550_buf_o2,
  lo570_buf_o2,
  lo582_buf_o2,
  n2302_inv,
  n2305_inv,
  n3499_o2,
  n2311_inv,
  n2870_o2,
  n2317_inv,
  n2689_o2,
  n2323_inv,
  n2662_o2,
  lo350_buf_o2,
  lo498_buf_o2,
  lo518_buf_o2,
  lo522_buf_o2,
  lo598_buf_o2,
  n2344_inv,
  n2347_inv,
  n2350_inv,
  n2353_inv,
  n2356_inv,
  n2359_inv,
  n2872_o2,
  n3313_o2,
  n3273_o2,
  n2848_o2,
  n2893_o2,
  n3267_o2,
  n2925_o2,
  n2839_o2,
  n2831_o2,
  n2558_o2,
  n2562_o2,
  n2825_o2,
  n3263_o2,
  n3517_o2,
  n2873_o2,
  n2926_o2,
  n3261_o2,
  n3268_o2,
  n3274_o2,
  n3314_o2,
  n3571_o2,
  n2950_o2,
  n2951_o2,
  n3022_o2,
  n3023_o2,
  n3057_o2,
  n3058_o2,
  n2931_o2,
  n2911_o2,
  n2959_o2,
  n2960_o2,
  n2922_o2,
  n2888_o2,
  n2889_o2,
  n3051_o2,
  n3052_o2,
  n3063_o2,
  n2845_o2,
  n2476_inv,
  n3281_o2,
  n3294_o2,
  n2885_o2,
  n2786_o2,
  n2783_o2,
  n2801_o2,
  n2572_o2,
  n2628_o2,
  n2609_o2,
  n2618_o2,
  n2637_o2,
  n2525_o2,
  n2551_o2,
  n3759_o2,
  n2994_o2,
  n3040_o2,
  n2943_o2,
  n2991_o2,
  n3034_o2,
  n2881_o2,
  n3021_o2,
  n3062_o2,
  n2763_o2,
  n2764_o2,
  n2775_o2,
  n2776_o2,
  n2968_o2,
  n2969_o2,
  n2798_o2,
  n3661_o2,
  n2694_o2,
  n2572_inv,
  n2817_o2,
  n2514_o2,
  n2501_o2,
  n2584_inv,
  n2505_o2,
  n2492_o2,
  lo546_buf_o2,
  lo590_buf_o2,
  lo594_buf_o2,
  n2602_inv,
  n2605_inv,
  n2709_o2,
  n2611_inv,
  n2614_inv,
  n2617_inv,
  n2620_inv,
  n3590_o2,
  n3591_o2,
  n2629_inv,
  n3638_o2,
  n3639_o2,
  n2638_inv,
  n2641_inv,
  lo458_buf_o2,
  lo482_buf_o2,
  lo566_buf_o2,
  n2718_o2,
  n3707_o2,
  n3671_o2,
  n3680_o2,
  n3749_o2,
  n3716_o2,
  n3692_o2,
  n2591_o2,
  n3478_o2,
  n3610_o2,
  n3611_o2,
  n2686_inv,
  n2689_inv,
  n2738_o2,
  n3616_o2,
  n3617_o2,
  n3031_o2,
  n2704_inv,
  n3562_o2,
  n2502_o2,
  n3560_o2,
  n3554_o2,
  n3555_o2,
  n3536_o2,
  n3537_o2,
  n3508_o2,
  n3650_o2,
  n3740_o2,
  n3484_o2,
  n2740_inv,
  n2734_o2,
  n2735_o2,
  n2711_o2,
  lo585_buf_o2,
  n2719_o2,
  n2720_o2,
  n2723_o2,
  n2724_o2,
  n3624_o2,
  n3625_o2,
  n3015_o2,
  n3491_o2,
  n2779_inv,
  n2811_o2,
  n3010_o2,
  n3012_o2,
  lo382_buf_o2,
  lo386_buf_o2,
  lo390_buf_o2,
  lo398_buf_o2,
  lo402_buf_o2,
  lo406_buf_o2,
  n3492_o2,
  lo366_buf_o2,
  lo374_buf_o2,
  lo426_buf_o2,
  lo494_buf_o2,
  n2653_o2,
  n2654_o2,
  n2715_o2,
  n2740_o2,
  n2682_o2,
  n2736_o2,
  lo508_buf_o2,
  lo512_buf_o2,
  lo536_buf_o2,
  lo576_buf_o2,
  lo357_buf_o2,
  lo361_buf_o2,
  lo417_buf_o2,
  lo421_buf_o2,
  lo473_buf_o2,
  lo477_buf_o2,
  lo553_buf_o2,
  lo557_buf_o2,
  lo573_buf_o2,
  lo434_buf_o2,
  lo438_buf_o2,
  lo466_buf_o2,
  lo470_buf_o2,
  lo490_buf_o2,
  n2657_o2,
  n2658_o2,
  n2663_o2,
  n2664_o2,
  n2684_o2,
  n2685_o2,
  G5193,
  G5194,
  G5195,
  G5196,
  G5197,
  G5198,
  G5199,
  G5200,
  G5201,
  G5202,
  G5203,
  G5204,
  G5205,
  G5206,
  G5207,
  G5208,
  G5209,
  G5210,
  G5211,
  G5212,
  G5213,
  G5214,
  G5215,
  G5216,
  G5217,
  G5218,
  G5219,
  G5220,
  G5221,
  G5222,
  G5223,
  G5224,
  G5225,
  G5226,
  G5227,
  G5228,
  G5229,
  G5230,
  G5231,
  G5232,
  G5233,
  G5234,
  G5235,
  G5236,
  G5237,
  G5238,
  G5239,
  G5240,
  G5241,
  G5242,
  G5243,
  G5244,
  G5245,
  G5246,
  G5247,
  G5248,
  G5249,
  G5250,
  G5251,
  G5252,
  G5253,
  G5254,
  G5255,
  G5256,
  G5257,
  G5258,
  G5259,
  G5260,
  G5261,
  G5262,
  G5263,
  G5264,
  G5265,
  G5266,
  G5267,
  G5268,
  G5269,
  G5270,
  G5271,
  G5272,
  G5273,
  G5274,
  G5275,
  G5276,
  G5277,
  G5278,
  G5279,
  G5280,
  G5281,
  G5282,
  G5283,
  G5284,
  G5285,
  G5286,
  G5287,
  G5288,
  G5289,
  G5290,
  G5291,
  G5292,
  G5293,
  G5294,
  G5295,
  G5296,
  G5297,
  G5298,
  G5299,
  G5300,
  G5301,
  G5302,
  G5303,
  G5304,
  G5305,
  G5306,
  G5307,
  G5308,
  G5309,
  G5310,
  G5311,
  G5312,
  G5313,
  G5314,
  G5315,
  n7230_li000_li000,
  n7233_li001_li001,
  n7236_li002_li002,
  n7239_li003_li003,
  n7242_li004_li004,
  n7245_li005_li005,
  n7248_li006_li006,
  n7254_li008_li008,
  n7257_li009_li009,
  n7260_li010_li010,
  n7263_li011_li011,
  n7266_li012_li012,
  n7269_li013_li013,
  n7272_li014_li014,
  n7275_li015_li015,
  n7278_li016_li016,
  n7281_li017_li017,
  n7284_li018_li018,
  n7287_li019_li019,
  n7290_li020_li020,
  n7293_li021_li021,
  n7296_li022_li022,
  n7299_li023_li023,
  n7302_li024_li024,
  n7305_li025_li025,
  n7308_li026_li026,
  n7311_li027_li027,
  n7314_li028_li028,
  n7317_li029_li029,
  n7320_li030_li030,
  n7323_li031_li031,
  n7326_li032_li032,
  n7329_li033_li033,
  n7332_li034_li034,
  n7335_li035_li035,
  n7338_li036_li036,
  n7341_li037_li037,
  n7344_li038_li038,
  n7347_li039_li039,
  n7350_li040_li040,
  n7353_li041_li041,
  n7356_li042_li042,
  n7359_li043_li043,
  n7362_li044_li044,
  n7365_li045_li045,
  n7368_li046_li046,
  n7371_li047_li047,
  n7374_li048_li048,
  n7377_li049_li049,
  n7380_li050_li050,
  n7383_li051_li051,
  n7386_li052_li052,
  n7389_li053_li053,
  n7392_li054_li054,
  n7395_li055_li055,
  n7398_li056_li056,
  n7401_li057_li057,
  n7404_li058_li058,
  n7407_li059_li059,
  n7410_li060_li060,
  n7413_li061_li061,
  n7416_li062_li062,
  n7419_li063_li063,
  n7422_li064_li064,
  n7425_li065_li065,
  n7428_li066_li066,
  n7431_li067_li067,
  n7434_li068_li068,
  n7437_li069_li069,
  n7440_li070_li070,
  n7443_li071_li071,
  n7446_li072_li072,
  n7449_li073_li073,
  n7452_li074_li074,
  n7458_li076_li076,
  n7461_li077_li077,
  n7464_li078_li078,
  n7467_li079_li079,
  n7470_li080_li080,
  n7473_li081_li081,
  n7476_li082_li082,
  n7482_li084_li084,
  n7485_li085_li085,
  n7488_li086_li086,
  n7491_li087_li087,
  n7494_li088_li088,
  n7497_li089_li089,
  n7500_li090_li090,
  n7503_li091_li091,
  n7506_li092_li092,
  n7509_li093_li093,
  n7512_li094_li094,
  n7515_li095_li095,
  n7518_li096_li096,
  n7521_li097_li097,
  n7524_li098_li098,
  n7527_li099_li099,
  n7530_li100_li100,
  n7533_li101_li101,
  n7536_li102_li102,
  n7539_li103_li103,
  n7542_li104_li104,
  n7545_li105_li105,
  n7548_li106_li106,
  n7551_li107_li107,
  n7554_li108_li108,
  n7557_li109_li109,
  n7560_li110_li110,
  n7563_li111_li111,
  n7566_li112_li112,
  n7569_li113_li113,
  n7572_li114_li114,
  n7575_li115_li115,
  n7578_li116_li116,
  n7581_li117_li117,
  n7584_li118_li118,
  n7587_li119_li119,
  n7590_li120_li120,
  n7593_li121_li121,
  n7596_li122_li122,
  n7599_li123_li123,
  n7602_li124_li124,
  n7605_li125_li125,
  n7608_li126_li126,
  n7611_li127_li127,
  n7614_li128_li128,
  n7617_li129_li129,
  n7620_li130_li130,
  n7623_li131_li131,
  n7626_li132_li132,
  n7629_li133_li133,
  n7632_li134_li134,
  n7635_li135_li135,
  n7638_li136_li136,
  n7641_li137_li137,
  n7644_li138_li138,
  n7647_li139_li139,
  n7650_li140_li140,
  n7653_li141_li141,
  n7656_li142_li142,
  n7659_li143_li143,
  n7662_li144_li144,
  n7665_li145_li145,
  n7668_li146_li146,
  n7671_li147_li147,
  n7674_li148_li148,
  n7677_li149_li149,
  n7680_li150_li150,
  n7683_li151_li151,
  n7686_li152_li152,
  n7689_li153_li153,
  n7692_li154_li154,
  n7695_li155_li155,
  n7698_li156_li156,
  n7701_li157_li157,
  n7704_li158_li158,
  n7707_li159_li159,
  n7710_li160_li160,
  n7713_li161_li161,
  n7716_li162_li162,
  n7719_li163_li163,
  n7722_li164_li164,
  n7725_li165_li165,
  n7728_li166_li166,
  n7731_li167_li167,
  n7734_li168_li168,
  n7737_li169_li169,
  n7740_li170_li170,
  n7746_li172_li172,
  n7749_li173_li173,
  n7752_li174_li174,
  n7758_li176_li176,
  n7761_li177_li177,
  n7764_li178_li178,
  n7767_li179_li179,
  n7770_li180_li180,
  n7773_li181_li181,
  n7776_li182_li182,
  n7782_li184_li184,
  n7785_li185_li185,
  n7788_li186_li186,
  n7794_li188_li188,
  n7797_li189_li189,
  n7800_li190_li190,
  n7806_li192_li192,
  n7809_li193_li193,
  n7812_li194_li194,
  n7815_li195_li195,
  n7818_li196_li196,
  n7821_li197_li197,
  n7824_li198_li198,
  n7830_li200_li200,
  n7833_li201_li201,
  n7836_li202_li202,
  n7839_li203_li203,
  n7842_li204_li204,
  n7845_li205_li205,
  n7848_li206_li206,
  n7854_li208_li208,
  n7857_li209_li209,
  n7860_li210_li210,
  n7863_li211_li211,
  n7866_li212_li212,
  n7869_li213_li213,
  n7872_li214_li214,
  n7875_li215_li215,
  n7878_li216_li216,
  n7881_li217_li217,
  n7884_li218_li218,
  n7887_li219_li219,
  n7890_li220_li220,
  n7893_li221_li221,
  n7896_li222_li222,
  n7899_li223_li223,
  n7902_li224_li224,
  n7905_li225_li225,
  n7908_li226_li226,
  n7914_li228_li228,
  n7917_li229_li229,
  n7920_li230_li230,
  n7926_li232_li232,
  n7929_li233_li233,
  n7932_li234_li234,
  n7938_li236_li236,
  n7941_li237_li237,
  n7944_li238_li238,
  n7950_li240_li240,
  n7953_li241_li241,
  n7956_li242_li242,
  n7959_li243_li243,
  n7962_li244_li244,
  n7965_li245_li245,
  n7968_li246_li246,
  n7971_li247_li247,
  n7974_li248_li248,
  n7977_li249_li249,
  n7980_li250_li250,
  n7983_li251_li251,
  n7986_li252_li252,
  n7989_li253_li253,
  n7992_li254_li254,
  n7995_li255_li255,
  n7998_li256_li256,
  n8001_li257_li257,
  n8004_li258_li258,
  n8007_li259_li259,
  n8010_li260_li260,
  n8013_li261_li261,
  n8016_li262_li262,
  n8019_li263_li263,
  n8022_li264_li264,
  n8025_li265_li265,
  n8028_li266_li266,
  n8031_li267_li267,
  n8034_li268_li268,
  n8037_li269_li269,
  n8040_li270_li270,
  n8043_li271_li271,
  n8046_li272_li272,
  n8049_li273_li273,
  n8052_li274_li274,
  n8055_li275_li275,
  n8058_li276_li276,
  n8061_li277_li277,
  n8064_li278_li278,
  n8067_li279_li279,
  n8070_li280_li280,
  n8073_li281_li281,
  n8076_li282_li282,
  n8079_li283_li283,
  n8082_li284_li284,
  n8085_li285_li285,
  n8088_li286_li286,
  n8091_li287_li287,
  n8094_li288_li288,
  n8097_li289_li289,
  n8100_li290_li290,
  n8103_li291_li291,
  n8106_li292_li292,
  n8109_li293_li293,
  n8112_li294_li294,
  n8115_li295_li295,
  n8118_li296_li296,
  n8121_li297_li297,
  n8124_li298_li298,
  n8127_li299_li299,
  n8130_li300_li300,
  n8133_li301_li301,
  n8136_li302_li302,
  n8139_li303_li303,
  n8142_li304_li304,
  n8145_li305_li305,
  n8148_li306_li306,
  n8151_li307_li307,
  n8154_li308_li308,
  n8157_li309_li309,
  n8160_li310_li310,
  n8163_li311_li311,
  n8166_li312_li312,
  n8169_li313_li313,
  n8172_li314_li314,
  n8175_li315_li315,
  n8178_li316_li316,
  n8181_li317_li317,
  n8184_li318_li318,
  n8187_li319_li319,
  n8190_li320_li320,
  n8193_li321_li321,
  n8196_li322_li322,
  n8199_li323_li323,
  n8202_li324_li324,
  n8205_li325_li325,
  n8208_li326_li326,
  n8211_li327_li327,
  n8214_li328_li328,
  n8217_li329_li329,
  n8220_li330_li330,
  n8223_li331_li331,
  n8226_li332_li332,
  n8229_li333_li333,
  n8232_li334_li334,
  n8235_li335_li335,
  n8238_li336_li336,
  n8241_li337_li337,
  n8244_li338_li338,
  n8247_li339_li339,
  n8250_li340_li340,
  n8253_li341_li341,
  n8256_li342_li342,
  n8259_li343_li343,
  n8262_li344_li344,
  n8265_li345_li345,
  n8268_li346_li346,
  n8271_li347_li347,
  n8274_li348_li348,
  n8286_li352_li352,
  n8370_li380_li380,
  n8382_li384_li384,
  n8394_li388_li388,
  n8406_li392_li392,
  n8409_li393_li393,
  n8412_li394_li394,
  n8415_li395_li395,
  n8418_li396_li396,
  n8430_li400_li400,
  n8442_li404_li404,
  n8454_li408_li408,
  n8466_li412_li412,
  n8550_li440_li440,
  n8553_li441_li441,
  n8556_li442_li442,
  n8562_li444_li444,
  n8565_li445_li445,
  n8568_li446_li446,
  n8574_li448_li448,
  n8577_li449_li449,
  n8583_li451_li451,
  n8586_li452_li452,
  n8589_li453_li453,
  n8595_li455_li455,
  n8598_li456_li456,
  n8610_li460_li460,
  n8670_li480_li480,
  n8682_li484_li484,
  n8718_li496_li496,
  n8727_li499_li499,
  n8730_li500_li500,
  n8742_li504_li504,
  n8751_li507_li507,
  n8775_li515_li515,
  n8778_li516_li516,
  n8790_li520_li520,
  n8799_li523_li523,
  n8802_li524_li524,
  n8805_li525_li525,
  n8808_li526_li526,
  n8814_li528_li528,
  n8817_li529_li529,
  n8820_li530_li530,
  n8826_li532_li532,
  n8829_li533_li533,
  n8832_li534_li534,
  n8835_li535_li535,
  n8850_li540_li540,
  n8853_li541_li541,
  n8856_li542_li542,
  n8859_li543_li543,
  n8862_li544_li544,
  n8874_li548_li548,
  n8910_li560_li560,
  n8913_li561_li561,
  n8922_li564_li564,
  n8934_li568_li568,
  n8970_li580_li580,
  n8982_li584_li584,
  n8994_li588_li588,
  n9006_li592_li592,
  n9018_li596_li596,
  n9030_li600_li600,
  n9033_li601_li601,
  n9036_li602_li602,
  n9039_li603_li603,
  n9042_li604_li604,
  n9045_li605_li605,
  n9048_li606_li606,
  n9051_li607_li607,
  n9054_li608_li608,
  n9057_li609_li609,
  n9060_li610_li610,
  n9063_li611_li611,
  n9066_li612_li612,
  n9069_li613_li613,
  n9072_li614_li614,
  n9075_li615_li615,
  n9078_li616_li616,
  n9081_li617_li617,
  n9084_li618_li618,
  n9087_li619_li619,
  n9090_li620_li620,
  n9093_li621_li621,
  n9096_li622_li622,
  n9099_li623_li623,
  n9102_li624_li624,
  n9105_li625_li625,
  n9108_li626_li626,
  n9114_li628_li628,
  n9117_li629_li629,
  n9120_li630_li630,
  n9123_li631_li631,
  n9126_li632_li632,
  n9129_li633_li633,
  n9132_li634_li634,
  n9135_li635_li635,
  n9138_li636_li636,
  n9141_li637_li637,
  n9144_li638_li638,
  n9147_li639_li639,
  n9150_li640_li640,
  n9153_li641_li641,
  n9156_li642_li642,
  n9159_li643_li643,
  n9162_li644_li644,
  n9165_li645_li645,
  n9174_li648_li648,
  n9177_li649_li649,
  n9180_li650_li650,
  n9183_li651_li651,
  n9186_li652_li652,
  n9189_li653_li653,
  n9192_li654_li654,
  n9195_li655_li655,
  n9198_li656_li656,
  n9201_li657_li657,
  n9204_li658_li658,
  n9207_li659_li659,
  n9210_li660_li660,
  n9213_li661_li661,
  n9216_li662_li662,
  n9222_li664_li664,
  n9225_li665_li665,
  n9228_li666_li666,
  n9234_li668_li668,
  n9237_li669_li669,
  n9240_li670_li670,
  n9246_li672_li672,
  n9249_li673_li673,
  n9252_li674_li674,
  n9258_li676_li676,
  n9261_li677_li677,
  n9264_li678_li678,
  n9267_li679_li679,
  n9270_li680_li680,
  n9273_li681_li681,
  n9276_li682_li682,
  n9279_li683_li683,
  n9282_li684_li684,
  n9285_li685_li685,
  n9288_li686_li686,
  n9291_li687_li687,
  n9294_li688_li688,
  n9297_li689_li689,
  n9300_li690_li690,
  n9303_li691_li691,
  n9306_li692_li692,
  n9309_li693_li693,
  n9312_li694_li694,
  n9315_li695_li695,
  n9318_li696_li696,
  n9321_li697_li697,
  n9324_li698_li698,
  n9327_li699_li699,
  n9330_li700_li700,
  n9333_li701_li701,
  n9336_li702_li702,
  n9339_li703_li703,
  n9342_li704_li704,
  n9345_li705_li705,
  n9348_li706_li706,
  n9351_li707_li707,
  n9354_li708_li708,
  n9357_li709_li709,
  n9360_li710_li710,
  n9363_li711_li711,
  n4970_i2,
  n4972_i2,
  n4989_i2,
  n5024_i2,
  n5025_i2,
  n5029_i2,
  n5042_i2,
  n5048_i2,
  n5093_i2,
  n5096_i2,
  n5193_i2,
  n5199_i2,
  n5203_i2,
  n5214_i2,
  n5221_i2,
  n5222_i2,
  n5273_i2,
  n5365_i2,
  n5385_i2,
  n5553_i2,
  n5636_i2,
  n5782_i2,
  n5778_i2,
  n5323_i2,
  n5325_i2,
  n5327_i2,
  n5329_i2,
  n5816_i2,
  n5817_i2,
  n5837_i2,
  n5844_i2,
  n5859_i2,
  n5857_i2,
  n5369_i2,
  n5371_i2,
  n5373_i2,
  n5400_i2,
  n5402_i2,
  n5404_i2,
  n5406_i2,
  n5407_i2,
  n5408_i2,
  n2722_i2,
  n5411_i2,
  n5412_i2,
  n5413_i2,
  n5557_i2,
  n5558_i2,
  n5559_i2,
  n5564_i2,
  n5565_i2,
  n5561_i2,
  n5568_i2,
  n5598_i2,
  n5600_i2,
  n5601_i2,
  n5602_i2,
  n5603_i2,
  n2853_i2,
  n5637_i2,
  n5627_i2,
  n5628_i2,
  n5635_i2,
  n5640_i2,
  n5641_i2,
  n5642_i2,
  n5650_i2,
  n5652_i2,
  n5653_i2,
  n5654_i2,
  n5655_i2,
  n5657_i2,
  n5659_i2,
  n5661_i2,
  n5656_i2,
  n5663_i2,
  n5664_i2,
  n5795_i2,
  n5796_i2,
  n5797_i2,
  n5739_i2,
  n5773_i2,
  n5798_i2,
  n5799_i2,
  n5802_i2,
  n5803_i2,
  n5831_i2,
  n5833_i2,
  n5820_i2,
  n5823_i2,
  n5824_i2,
  n5869_i2,
  n5848_i2,
  n5849_i2,
  n5856_i2,
  n5896_i2,
  n2754_i2,
  n2908_i2,
  n5892_i2,
  n5915_i2,
  n5919_i2,
  n5918_i2,
  n5920_i2,
  n5917_i2,
  lo586_buf_i2,
  n2818_i2,
  n2863_i2,
  n2721_i2,
  n2725_i2,
  n3016_i2,
  n3013_i2,
  n2655_i2,
  n2741_i2,
  lo562_buf_i2,
  n2656_i2,
  n2531_i2,
  n2700_i2,
  n5908_i2,
  n5910_i2,
  n5912_i2,
  n5914_i2,
  n2753_i2,
  n2878_i2,
  n2836_i2,
  n5934_i2,
  n5936_i2,
  n5938_i2,
  n2728_i2,
  lo358_buf_i2,
  lo418_buf_i2,
  lo474_buf_i2,
  lo554_buf_i2,
  lo558_buf_i2,
  lo574_buf_i2,
  n2659_i2,
  n2665_i2,
  n2686_i2,
  lo450_buf_i2,
  n2910_i2,
  n2683_i2,
  n2828_i2,
  n2582_i2,
  n2600_i2,
  n2542_i2,
  n2703_i2,
  lo510_buf_i2,
  lo514_buf_i2,
  lo538_buf_i2,
  lo578_buf_i2,
  n2692_i2,
  n2666_i2,
  n2667_i2,
  n2660_i2,
  n2744_i2,
  lo454_buf_i2,
  n3593_i2,
  n3048_i2,
  lo410_buf_i2,
  lo502_buf_i2,
  lo506_buf_i2,
  lo550_buf_i2,
  lo570_buf_i2,
  lo582_buf_i2,
  n2646_i2,
  n2673_i2,
  n3499_i2,
  n2750_i2,
  n2870_i2,
  n2693_i2,
  n2689_i2,
  n2668_i2,
  n2662_i2,
  lo350_buf_i2,
  lo498_buf_i2,
  lo518_buf_i2,
  lo522_buf_i2,
  lo598_buf_i2,
  n2708_i2,
  n2674_i2,
  n2647_i2,
  n2751_i2,
  n2747_i2,
  n2669_i2,
  n2872_i2,
  n3313_i2,
  n3273_i2,
  n2848_i2,
  n2893_i2,
  n3267_i2,
  n2925_i2,
  n2839_i2,
  n2831_i2,
  n2558_i2,
  n2562_i2,
  n2825_i2,
  n3263_i2,
  n3517_i2,
  n2873_i2,
  n2926_i2,
  n3261_i2,
  n3268_i2,
  n3274_i2,
  n3314_i2,
  n3571_i2,
  n2950_i2,
  n2951_i2,
  n3022_i2,
  n3023_i2,
  n3057_i2,
  n3058_i2,
  n2931_i2,
  n2911_i2,
  n2959_i2,
  n2960_i2,
  n2922_i2,
  n2888_i2,
  n2889_i2,
  n3051_i2,
  n3052_i2,
  n3063_i2,
  n2845_i2,
  n2737_i2,
  n3281_i2,
  n3294_i2,
  n2885_i2,
  n2786_i2,
  n2783_i2,
  n2801_i2,
  n2572_i2,
  n2628_i2,
  n2609_i2,
  n2618_i2,
  n2637_i2,
  n2525_i2,
  n2551_i2,
  n3759_i2,
  n2994_i2,
  n3040_i2,
  n2943_i2,
  n2991_i2,
  n3034_i2,
  n2881_i2,
  n3021_i2,
  n3062_i2,
  n2763_i2,
  n2764_i2,
  n2775_i2,
  n2776_i2,
  n2968_i2,
  n2969_i2,
  n2798_i2,
  n3661_i2,
  n2694_i2,
  n2809_i2,
  n2817_i2,
  n2514_i2,
  n2501_i2,
  n2528_i2,
  n2505_i2,
  n2492_i2,
  lo546_buf_i2,
  lo590_buf_i2,
  lo594_buf_i2,
  n2679_i2,
  n2733_i2,
  n2709_i2,
  n2676_i2,
  n2649_i2,
  n2815_i2,
  n2704_i2,
  n3590_i2,
  n3591_i2,
  n2752_i2,
  n3638_i2,
  n3639_i2,
  n2695_i2,
  n3047_i2,
  lo458_buf_i2,
  lo482_buf_i2,
  lo566_buf_i2,
  n2718_i2,
  n3707_i2,
  n3671_i2,
  n3680_i2,
  n3749_i2,
  n3716_i2,
  n3692_i2,
  n2591_i2,
  n3478_i2,
  n3610_i2,
  n3611_i2,
  n2652_i2,
  n2714_i2,
  n2738_i2,
  n3616_i2,
  n3617_i2,
  n3031_i2,
  n2515_i2,
  n3562_i2,
  n2502_i2,
  n3560_i2,
  n3554_i2,
  n3555_i2,
  n3536_i2,
  n3537_i2,
  n3508_i2,
  n3650_i2,
  n3740_i2,
  n3484_i2,
  n2680_i2,
  n2734_i2,
  n2735_i2,
  n2711_i2,
  lo585_buf_i2,
  n2719_i2,
  n2720_i2,
  n2723_i2,
  n2724_i2,
  n3624_i2,
  n3625_i2,
  n3015_i2,
  n3491_i2,
  n2696_i2,
  n2811_i2,
  n3010_i2,
  n3012_i2,
  lo382_buf_i2,
  lo386_buf_i2,
  lo390_buf_i2,
  lo398_buf_i2,
  lo402_buf_i2,
  lo406_buf_i2,
  n3492_i2,
  lo366_buf_i2,
  lo374_buf_i2,
  lo426_buf_i2,
  lo494_buf_i2,
  n2653_i2,
  n2654_i2,
  n2715_i2,
  n2740_i2,
  n2682_i2,
  n2736_i2,
  lo508_buf_i2,
  lo512_buf_i2,
  lo536_buf_i2,
  lo576_buf_i2,
  lo357_buf_i2,
  lo361_buf_i2,
  lo417_buf_i2,
  lo421_buf_i2,
  lo473_buf_i2,
  lo477_buf_i2,
  lo553_buf_i2,
  lo557_buf_i2,
  lo573_buf_i2,
  lo434_buf_i2,
  lo438_buf_i2,
  lo466_buf_i2,
  lo470_buf_i2,
  lo490_buf_i2,
  n2657_i2,
  n2658_i2,
  n2663_i2,
  n2664_i2,
  n2684_i2,
  n2685_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input G42;input G43;input G44;input G45;input G46;input G47;input G48;input G49;input G50;input G51;input G52;input G53;input G54;input G55;input G56;input G57;input G58;input G59;input G60;input G61;input G62;input G63;input G64;input G65;input G66;input G67;input G68;input G69;input G70;input G71;input G72;input G73;input G74;input G75;input G76;input G77;input G78;input G79;input G80;input G81;input G82;input G83;input G84;input G85;input G86;input G87;input G88;input G89;input G90;input G91;input G92;input G93;input G94;input G95;input G96;input G97;input G98;input G99;input G100;input G101;input G102;input G103;input G104;input G105;input G106;input G107;input G108;input G109;input G110;input G111;input G112;input G113;input G114;input G115;input G116;input G117;input G118;input G119;input G120;input G121;input G122;input G123;input G124;input G125;input G126;input G127;input G128;input G129;input G130;input G131;input G132;input G133;input G134;input G135;input G136;input G137;input G138;input G139;input G140;input G141;input G142;input G143;input G144;input G145;input G146;input G147;input G148;input G149;input G150;input G151;input G152;input G153;input G154;input G155;input G156;input G157;input G158;input G159;input G160;input G161;input G162;input G163;input G164;input G165;input G166;input G167;input G168;input G169;input G170;input G171;input G172;input G173;input G174;input G175;input G176;input G177;input G178;input n2610_lo;input n2613_lo;input n2616_lo;input n2619_lo;input n2622_lo;input n2625_lo;input n2628_lo;input n2634_lo;input n2637_lo;input n2640_lo;input n2643_lo;input n2646_lo;input n2649_lo;input n2652_lo;input n2655_lo;input n2658_lo;input n2661_lo;input n2664_lo;input n2667_lo;input n2670_lo;input n2673_lo;input n2676_lo;input n2679_lo;input n2682_lo;input n2685_lo;input n2688_lo;input n2691_lo;input n2694_lo;input n2697_lo;input n2700_lo;input n2703_lo;input n2706_lo;input n2709_lo;input n2712_lo;input n2715_lo;input n2718_lo;input n2721_lo;input n2724_lo;input n2727_lo;input n2730_lo;input n2733_lo;input n2736_lo;input n2739_lo;input n2742_lo;input n2745_lo;input n2748_lo;input n2751_lo;input n2754_lo;input n2757_lo;input n2760_lo;input n2763_lo;input n2766_lo;input n2769_lo;input n2772_lo;input n2775_lo;input n2778_lo;input n2781_lo;input n2784_lo;input n2787_lo;input n2790_lo;input n2793_lo;input n2796_lo;input n2799_lo;input n2802_lo;input n2805_lo;input n2808_lo;input n2811_lo;input n2814_lo;input n2817_lo;input n2820_lo;input n2823_lo;input n2826_lo;input n2829_lo;input n2832_lo;input n2838_lo;input n2841_lo;input n2844_lo;input n2847_lo;input n2850_lo;input n2853_lo;input n2856_lo;input n2862_lo;input n2865_lo;input n2868_lo;input n2871_lo;input n2874_lo;input n2877_lo;input n2880_lo;input n2883_lo;input n2886_lo;input n2889_lo;input n2892_lo;input n2895_lo;input n2898_lo;input n2901_lo;input n2904_lo;input n2907_lo;input n2910_lo;input n2913_lo;input n2916_lo;input n2919_lo;input n2922_lo;input n2925_lo;input n2928_lo;input n2931_lo;input n2934_lo;input n2937_lo;input n2940_lo;input n2943_lo;input n2946_lo;input n2949_lo;input n2952_lo;input n2955_lo;input n2958_lo;input n2961_lo;input n2964_lo;input n2967_lo;input n2970_lo;input n2973_lo;input n2976_lo;input n2979_lo;input n2982_lo;input n2985_lo;input n2988_lo;input n2991_lo;input n2994_lo;input n2997_lo;input n3000_lo;input n3003_lo;input n3006_lo;input n3009_lo;input n3012_lo;input n3015_lo;input n3018_lo;input n3021_lo;input n3024_lo;input n3027_lo;input n3030_lo;input n3033_lo;input n3036_lo;input n3039_lo;input n3042_lo;input n3045_lo;input n3048_lo;input n3051_lo;input n3054_lo;input n3057_lo;input n3060_lo;input n3063_lo;input n3066_lo;input n3069_lo;input n3072_lo;input n3075_lo;input n3078_lo;input n3081_lo;input n3084_lo;input n3087_lo;input n3090_lo;input n3093_lo;input n3096_lo;input n3099_lo;input n3102_lo;input n3105_lo;input n3108_lo;input n3111_lo;input n3114_lo;input n3117_lo;input n3120_lo;input n3126_lo;input n3129_lo;input n3132_lo;input n3138_lo;input n3141_lo;input n3144_lo;input n3147_lo;input n3150_lo;input n3153_lo;input n3156_lo;input n3162_lo;input n3165_lo;input n3168_lo;input n3174_lo;input n3177_lo;input n3180_lo;input n3186_lo;input n3189_lo;input n3192_lo;input n3195_lo;input n3198_lo;input n3201_lo;input n3204_lo;input n3210_lo;input n3213_lo;input n3216_lo;input n3219_lo;input n3222_lo;input n3225_lo;input n3228_lo;input n3234_lo;input n3237_lo;input n3240_lo;input n3243_lo;input n3246_lo;input n3249_lo;input n3252_lo;input n3255_lo;input n3258_lo;input n3261_lo;input n3264_lo;input n3267_lo;input n3270_lo;input n3273_lo;input n3276_lo;input n3279_lo;input n3282_lo;input n3285_lo;input n3288_lo;input n3294_lo;input n3297_lo;input n3300_lo;input n3306_lo;input n3309_lo;input n3312_lo;input n3318_lo;input n3321_lo;input n3324_lo;input n3330_lo;input n3333_lo;input n3336_lo;input n3339_lo;input n3342_lo;input n3345_lo;input n3348_lo;input n3351_lo;input n3354_lo;input n3357_lo;input n3360_lo;input n3363_lo;input n3366_lo;input n3369_lo;input n3372_lo;input n3375_lo;input n3378_lo;input n3381_lo;input n3384_lo;input n3387_lo;input n3390_lo;input n3393_lo;input n3396_lo;input n3399_lo;input n3402_lo;input n3405_lo;input n3408_lo;input n3411_lo;input n3414_lo;input n3417_lo;input n3420_lo;input n3423_lo;input n3426_lo;input n3429_lo;input n3432_lo;input n3435_lo;input n3438_lo;input n3441_lo;input n3444_lo;input n3447_lo;input n3450_lo;input n3453_lo;input n3456_lo;input n3459_lo;input n3462_lo;input n3465_lo;input n3468_lo;input n3471_lo;input n3474_lo;input n3477_lo;input n3480_lo;input n3483_lo;input n3486_lo;input n3489_lo;input n3492_lo;input n3495_lo;input n3498_lo;input n3501_lo;input n3504_lo;input n3507_lo;input n3510_lo;input n3513_lo;input n3516_lo;input n3519_lo;input n3522_lo;input n3525_lo;input n3528_lo;input n3531_lo;input n3534_lo;input n3537_lo;input n3540_lo;input n3543_lo;input n3546_lo;input n3549_lo;input n3552_lo;input n3555_lo;input n3558_lo;input n3561_lo;input n3564_lo;input n3567_lo;input n3570_lo;input n3573_lo;input n3576_lo;input n3579_lo;input n3582_lo;input n3585_lo;input n3588_lo;input n3591_lo;input n3594_lo;input n3597_lo;input n3600_lo;input n3603_lo;input n3606_lo;input n3609_lo;input n3612_lo;input n3615_lo;input n3618_lo;input n3621_lo;input n3624_lo;input n3627_lo;input n3630_lo;input n3633_lo;input n3636_lo;input n3639_lo;input n3642_lo;input n3645_lo;input n3648_lo;input n3651_lo;input n3654_lo;input n3666_lo;input n3750_lo;input n3762_lo;input n3774_lo;input n3786_lo;input n3789_lo;input n3792_lo;input n3795_lo;input n3798_lo;input n3810_lo;input n3822_lo;input n3834_lo;input n3846_lo;input n3930_lo;input n3933_lo;input n3936_lo;input n3942_lo;input n3945_lo;input n3948_lo;input n3954_lo;input n3957_lo;input n3963_lo;input n3966_lo;input n3969_lo;input n3975_lo;input n3978_lo;input n3990_lo;input n4050_lo;input n4062_lo;input n4098_lo;input n4107_lo;input n4110_lo;input n4122_lo;input n4131_lo;input n4155_lo;input n4158_lo;input n4170_lo;input n4179_lo;input n4182_lo;input n4185_lo;input n4188_lo;input n4194_lo;input n4197_lo;input n4200_lo;input n4206_lo;input n4209_lo;input n4212_lo;input n4215_lo;input n4230_lo;input n4233_lo;input n4236_lo;input n4239_lo;input n4242_lo;input n4254_lo;input n4290_lo;input n4293_lo;input n4302_lo;input n4314_lo;input n4350_lo;input n4362_lo;input n4374_lo;input n4386_lo;input n4398_lo;input n4410_lo;input n4413_lo;input n4416_lo;input n4419_lo;input n4422_lo;input n4425_lo;input n4428_lo;input n4431_lo;input n4434_lo;input n4437_lo;input n4440_lo;input n4443_lo;input n4446_lo;input n4449_lo;input n4452_lo;input n4455_lo;input n4458_lo;input n4461_lo;input n4464_lo;input n4467_lo;input n4470_lo;input n4473_lo;input n4476_lo;input n4479_lo;input n4482_lo;input n4485_lo;input n4488_lo;input n4494_lo;input n4497_lo;input n4500_lo;input n4503_lo;input n4506_lo;input n4509_lo;input n4512_lo;input n4515_lo;input n4518_lo;input n4521_lo;input n4524_lo;input n4527_lo;input n4530_lo;input n4533_lo;input n4536_lo;input n4539_lo;input n4542_lo;input n4545_lo;input n4554_lo;input n4557_lo;input n4560_lo;input n4563_lo;input n4566_lo;input n4569_lo;input n4572_lo;input n4575_lo;input n4578_lo;input n4581_lo;input n4584_lo;input n4587_lo;input n4590_lo;input n4593_lo;input n4596_lo;input n4602_lo;input n4605_lo;input n4608_lo;input n4614_lo;input n4617_lo;input n4620_lo;input n4626_lo;input n4629_lo;input n4632_lo;input n4638_lo;input n4641_lo;input n4644_lo;input n4647_lo;input n4650_lo;input n4653_lo;input n4656_lo;input n4659_lo;input n4662_lo;input n4665_lo;input n4668_lo;input n4671_lo;input n4674_lo;input n4677_lo;input n4680_lo;input n4683_lo;input n4686_lo;input n4689_lo;input n4692_lo;input n4695_lo;input n4698_lo;input n4701_lo;input n4704_lo;input n4707_lo;input n4710_lo;input n4713_lo;input n4716_lo;input n4719_lo;input n4722_lo;input n4725_lo;input n4728_lo;input n4731_lo;input n4734_lo;input n4737_lo;input n4740_lo;input n4743_lo;input n4970_o2;input n4972_o2;input n4989_o2;input n5024_o2;input n5025_o2;input n5029_o2;input n5042_o2;input n5048_o2;input n5093_o2;input n5096_o2;input n5193_o2;input n5199_o2;input n5203_o2;input n5214_o2;input n5221_o2;input n5222_o2;input n5273_o2;input n5365_o2;input n5385_o2;input n5553_o2;input n5636_o2;input n5782_o2;input n5778_o2;input n5323_o2;input n5325_o2;input n5327_o2;input n5329_o2;input n5816_o2;input n5817_o2;input n5837_o2;input n5844_o2;input n5859_o2;input n5857_o2;input n5369_o2;input n5371_o2;input n5373_o2;input n5400_o2;input n5402_o2;input n5404_o2;input n5406_o2;input n5407_o2;input n5408_o2;input n2722_o2;input n1942_inv;input n5412_o2;input n1948_inv;input n5557_o2;input n5558_o2;input n5559_o2;input n5564_o2;input n5565_o2;input n1966_inv;input n5568_o2;input n5598_o2;input n5600_o2;input n5601_o2;input n5602_o2;input n5603_o2;input n2853_o2;input n5637_o2;input n1993_inv;input n1996_inv;input n5635_o2;input n5640_o2;input n5641_o2;input n5642_o2;input n5650_o2;input n5652_o2;input n5653_o2;input n5654_o2;input n5655_o2;input n5657_o2;input n2029_inv;input n5661_o2;input n5656_o2;input n5663_o2;input n2041_inv;input n5795_o2;input n5796_o2;input n5797_o2;input n5739_o2;input n5773_o2;input n2059_inv;input n5799_o2;input n5802_o2;input n2068_inv;input n5831_o2;input n5833_o2;input n5820_o2;input n5823_o2;input n5824_o2;input n5869_o2;input n5848_o2;input n5849_o2;input n5856_o2;input n5896_o2;input n2754_o2;input n2908_o2;input n5892_o2;input n5915_o2;input n5919_o2;input n5918_o2;input n5920_o2;input n5917_o2;input lo586_buf_o2;input n2818_o2;input n2863_o2;input n2134_inv;input n2725_o2;input n3016_o2;input n3013_o2;input n2655_o2;input n2149_inv;input lo562_buf_o2;input n2155_inv;input n2531_o2;input n2700_o2;input n5908_o2;input n5910_o2;input n5912_o2;input n5914_o2;input n2753_o2;input n2878_o2;input n2182_inv;input n5934_o2;input n5936_o2;input n5938_o2;input n2728_o2;input lo358_buf_o2;input lo418_buf_o2;input lo474_buf_o2;input lo554_buf_o2;input lo558_buf_o2;input lo574_buf_o2;input n2215_inv;input n2218_inv;input n2221_inv;input lo450_buf_o2;input n2910_o2;input n2683_o2;input n2828_o2;input n2582_o2;input n2600_o2;input n2542_o2;input n2703_o2;input lo510_buf_o2;input lo514_buf_o2;input lo538_buf_o2;input lo578_buf_o2;input n2260_inv;input n2666_o2;input n2667_o2;input n2660_o2;input n2272_inv;input lo454_buf_o2;input n3593_o2;input n3048_o2;input lo410_buf_o2;input lo502_buf_o2;input lo506_buf_o2;input lo550_buf_o2;input lo570_buf_o2;input lo582_buf_o2;input n2302_inv;input n2305_inv;input n3499_o2;input n2311_inv;input n2870_o2;input n2317_inv;input n2689_o2;input n2323_inv;input n2662_o2;input lo350_buf_o2;input lo498_buf_o2;input lo518_buf_o2;input lo522_buf_o2;input lo598_buf_o2;input n2344_inv;input n2347_inv;input n2350_inv;input n2353_inv;input n2356_inv;input n2359_inv;input n2872_o2;input n3313_o2;input n3273_o2;input n2848_o2;input n2893_o2;input n3267_o2;input n2925_o2;input n2839_o2;input n2831_o2;input n2558_o2;input n2562_o2;input n2825_o2;input n3263_o2;input n3517_o2;input n2873_o2;input n2926_o2;input n3261_o2;input n3268_o2;input n3274_o2;input n3314_o2;input n3571_o2;input n2950_o2;input n2951_o2;input n3022_o2;input n3023_o2;input n3057_o2;input n3058_o2;input n2931_o2;input n2911_o2;input n2959_o2;input n2960_o2;input n2922_o2;input n2888_o2;input n2889_o2;input n3051_o2;input n3052_o2;input n3063_o2;input n2845_o2;input n2476_inv;input n3281_o2;input n3294_o2;input n2885_o2;input n2786_o2;input n2783_o2;input n2801_o2;input n2572_o2;input n2628_o2;input n2609_o2;input n2618_o2;input n2637_o2;input n2525_o2;input n2551_o2;input n3759_o2;input n2994_o2;input n3040_o2;input n2943_o2;input n2991_o2;input n3034_o2;input n2881_o2;input n3021_o2;input n3062_o2;input n2763_o2;input n2764_o2;input n2775_o2;input n2776_o2;input n2968_o2;input n2969_o2;input n2798_o2;input n3661_o2;input n2694_o2;input n2572_inv;input n2817_o2;input n2514_o2;input n2501_o2;input n2584_inv;input n2505_o2;input n2492_o2;input lo546_buf_o2;input lo590_buf_o2;input lo594_buf_o2;input n2602_inv;input n2605_inv;input n2709_o2;input n2611_inv;input n2614_inv;input n2617_inv;input n2620_inv;input n3590_o2;input n3591_o2;input n2629_inv;input n3638_o2;input n3639_o2;input n2638_inv;input n2641_inv;input lo458_buf_o2;input lo482_buf_o2;input lo566_buf_o2;input n2718_o2;input n3707_o2;input n3671_o2;input n3680_o2;input n3749_o2;input n3716_o2;input n3692_o2;input n2591_o2;input n3478_o2;input n3610_o2;input n3611_o2;input n2686_inv;input n2689_inv;input n2738_o2;input n3616_o2;input n3617_o2;input n3031_o2;input n2704_inv;input n3562_o2;input n2502_o2;input n3560_o2;input n3554_o2;input n3555_o2;input n3536_o2;input n3537_o2;input n3508_o2;input n3650_o2;input n3740_o2;input n3484_o2;input n2740_inv;input n2734_o2;input n2735_o2;input n2711_o2;input lo585_buf_o2;input n2719_o2;input n2720_o2;input n2723_o2;input n2724_o2;input n3624_o2;input n3625_o2;input n3015_o2;input n3491_o2;input n2779_inv;input n2811_o2;input n3010_o2;input n3012_o2;input lo382_buf_o2;input lo386_buf_o2;input lo390_buf_o2;input lo398_buf_o2;input lo402_buf_o2;input lo406_buf_o2;input n3492_o2;input lo366_buf_o2;input lo374_buf_o2;input lo426_buf_o2;input lo494_buf_o2;input n2653_o2;input n2654_o2;input n2715_o2;input n2740_o2;input n2682_o2;input n2736_o2;input lo508_buf_o2;input lo512_buf_o2;input lo536_buf_o2;input lo576_buf_o2;input lo357_buf_o2;input lo361_buf_o2;input lo417_buf_o2;input lo421_buf_o2;input lo473_buf_o2;input lo477_buf_o2;input lo553_buf_o2;input lo557_buf_o2;input lo573_buf_o2;input lo434_buf_o2;input lo438_buf_o2;input lo466_buf_o2;input lo470_buf_o2;input lo490_buf_o2;input n2657_o2;input n2658_o2;input n2663_o2;input n2664_o2;input n2684_o2;input n2685_o2;
  output G5193;output G5194;output G5195;output G5196;output G5197;output G5198;output G5199;output G5200;output G5201;output G5202;output G5203;output G5204;output G5205;output G5206;output G5207;output G5208;output G5209;output G5210;output G5211;output G5212;output G5213;output G5214;output G5215;output G5216;output G5217;output G5218;output G5219;output G5220;output G5221;output G5222;output G5223;output G5224;output G5225;output G5226;output G5227;output G5228;output G5229;output G5230;output G5231;output G5232;output G5233;output G5234;output G5235;output G5236;output G5237;output G5238;output G5239;output G5240;output G5241;output G5242;output G5243;output G5244;output G5245;output G5246;output G5247;output G5248;output G5249;output G5250;output G5251;output G5252;output G5253;output G5254;output G5255;output G5256;output G5257;output G5258;output G5259;output G5260;output G5261;output G5262;output G5263;output G5264;output G5265;output G5266;output G5267;output G5268;output G5269;output G5270;output G5271;output G5272;output G5273;output G5274;output G5275;output G5276;output G5277;output G5278;output G5279;output G5280;output G5281;output G5282;output G5283;output G5284;output G5285;output G5286;output G5287;output G5288;output G5289;output G5290;output G5291;output G5292;output G5293;output G5294;output G5295;output G5296;output G5297;output G5298;output G5299;output G5300;output G5301;output G5302;output G5303;output G5304;output G5305;output G5306;output G5307;output G5308;output G5309;output G5310;output G5311;output G5312;output G5313;output G5314;output G5315;output n7230_li000_li000;output n7233_li001_li001;output n7236_li002_li002;output n7239_li003_li003;output n7242_li004_li004;output n7245_li005_li005;output n7248_li006_li006;output n7254_li008_li008;output n7257_li009_li009;output n7260_li010_li010;output n7263_li011_li011;output n7266_li012_li012;output n7269_li013_li013;output n7272_li014_li014;output n7275_li015_li015;output n7278_li016_li016;output n7281_li017_li017;output n7284_li018_li018;output n7287_li019_li019;output n7290_li020_li020;output n7293_li021_li021;output n7296_li022_li022;output n7299_li023_li023;output n7302_li024_li024;output n7305_li025_li025;output n7308_li026_li026;output n7311_li027_li027;output n7314_li028_li028;output n7317_li029_li029;output n7320_li030_li030;output n7323_li031_li031;output n7326_li032_li032;output n7329_li033_li033;output n7332_li034_li034;output n7335_li035_li035;output n7338_li036_li036;output n7341_li037_li037;output n7344_li038_li038;output n7347_li039_li039;output n7350_li040_li040;output n7353_li041_li041;output n7356_li042_li042;output n7359_li043_li043;output n7362_li044_li044;output n7365_li045_li045;output n7368_li046_li046;output n7371_li047_li047;output n7374_li048_li048;output n7377_li049_li049;output n7380_li050_li050;output n7383_li051_li051;output n7386_li052_li052;output n7389_li053_li053;output n7392_li054_li054;output n7395_li055_li055;output n7398_li056_li056;output n7401_li057_li057;output n7404_li058_li058;output n7407_li059_li059;output n7410_li060_li060;output n7413_li061_li061;output n7416_li062_li062;output n7419_li063_li063;output n7422_li064_li064;output n7425_li065_li065;output n7428_li066_li066;output n7431_li067_li067;output n7434_li068_li068;output n7437_li069_li069;output n7440_li070_li070;output n7443_li071_li071;output n7446_li072_li072;output n7449_li073_li073;output n7452_li074_li074;output n7458_li076_li076;output n7461_li077_li077;output n7464_li078_li078;output n7467_li079_li079;output n7470_li080_li080;output n7473_li081_li081;output n7476_li082_li082;output n7482_li084_li084;output n7485_li085_li085;output n7488_li086_li086;output n7491_li087_li087;output n7494_li088_li088;output n7497_li089_li089;output n7500_li090_li090;output n7503_li091_li091;output n7506_li092_li092;output n7509_li093_li093;output n7512_li094_li094;output n7515_li095_li095;output n7518_li096_li096;output n7521_li097_li097;output n7524_li098_li098;output n7527_li099_li099;output n7530_li100_li100;output n7533_li101_li101;output n7536_li102_li102;output n7539_li103_li103;output n7542_li104_li104;output n7545_li105_li105;output n7548_li106_li106;output n7551_li107_li107;output n7554_li108_li108;output n7557_li109_li109;output n7560_li110_li110;output n7563_li111_li111;output n7566_li112_li112;output n7569_li113_li113;output n7572_li114_li114;output n7575_li115_li115;output n7578_li116_li116;output n7581_li117_li117;output n7584_li118_li118;output n7587_li119_li119;output n7590_li120_li120;output n7593_li121_li121;output n7596_li122_li122;output n7599_li123_li123;output n7602_li124_li124;output n7605_li125_li125;output n7608_li126_li126;output n7611_li127_li127;output n7614_li128_li128;output n7617_li129_li129;output n7620_li130_li130;output n7623_li131_li131;output n7626_li132_li132;output n7629_li133_li133;output n7632_li134_li134;output n7635_li135_li135;output n7638_li136_li136;output n7641_li137_li137;output n7644_li138_li138;output n7647_li139_li139;output n7650_li140_li140;output n7653_li141_li141;output n7656_li142_li142;output n7659_li143_li143;output n7662_li144_li144;output n7665_li145_li145;output n7668_li146_li146;output n7671_li147_li147;output n7674_li148_li148;output n7677_li149_li149;output n7680_li150_li150;output n7683_li151_li151;output n7686_li152_li152;output n7689_li153_li153;output n7692_li154_li154;output n7695_li155_li155;output n7698_li156_li156;output n7701_li157_li157;output n7704_li158_li158;output n7707_li159_li159;output n7710_li160_li160;output n7713_li161_li161;output n7716_li162_li162;output n7719_li163_li163;output n7722_li164_li164;output n7725_li165_li165;output n7728_li166_li166;output n7731_li167_li167;output n7734_li168_li168;output n7737_li169_li169;output n7740_li170_li170;output n7746_li172_li172;output n7749_li173_li173;output n7752_li174_li174;output n7758_li176_li176;output n7761_li177_li177;output n7764_li178_li178;output n7767_li179_li179;output n7770_li180_li180;output n7773_li181_li181;output n7776_li182_li182;output n7782_li184_li184;output n7785_li185_li185;output n7788_li186_li186;output n7794_li188_li188;output n7797_li189_li189;output n7800_li190_li190;output n7806_li192_li192;output n7809_li193_li193;output n7812_li194_li194;output n7815_li195_li195;output n7818_li196_li196;output n7821_li197_li197;output n7824_li198_li198;output n7830_li200_li200;output n7833_li201_li201;output n7836_li202_li202;output n7839_li203_li203;output n7842_li204_li204;output n7845_li205_li205;output n7848_li206_li206;output n7854_li208_li208;output n7857_li209_li209;output n7860_li210_li210;output n7863_li211_li211;output n7866_li212_li212;output n7869_li213_li213;output n7872_li214_li214;output n7875_li215_li215;output n7878_li216_li216;output n7881_li217_li217;output n7884_li218_li218;output n7887_li219_li219;output n7890_li220_li220;output n7893_li221_li221;output n7896_li222_li222;output n7899_li223_li223;output n7902_li224_li224;output n7905_li225_li225;output n7908_li226_li226;output n7914_li228_li228;output n7917_li229_li229;output n7920_li230_li230;output n7926_li232_li232;output n7929_li233_li233;output n7932_li234_li234;output n7938_li236_li236;output n7941_li237_li237;output n7944_li238_li238;output n7950_li240_li240;output n7953_li241_li241;output n7956_li242_li242;output n7959_li243_li243;output n7962_li244_li244;output n7965_li245_li245;output n7968_li246_li246;output n7971_li247_li247;output n7974_li248_li248;output n7977_li249_li249;output n7980_li250_li250;output n7983_li251_li251;output n7986_li252_li252;output n7989_li253_li253;output n7992_li254_li254;output n7995_li255_li255;output n7998_li256_li256;output n8001_li257_li257;output n8004_li258_li258;output n8007_li259_li259;output n8010_li260_li260;output n8013_li261_li261;output n8016_li262_li262;output n8019_li263_li263;output n8022_li264_li264;output n8025_li265_li265;output n8028_li266_li266;output n8031_li267_li267;output n8034_li268_li268;output n8037_li269_li269;output n8040_li270_li270;output n8043_li271_li271;output n8046_li272_li272;output n8049_li273_li273;output n8052_li274_li274;output n8055_li275_li275;output n8058_li276_li276;output n8061_li277_li277;output n8064_li278_li278;output n8067_li279_li279;output n8070_li280_li280;output n8073_li281_li281;output n8076_li282_li282;output n8079_li283_li283;output n8082_li284_li284;output n8085_li285_li285;output n8088_li286_li286;output n8091_li287_li287;output n8094_li288_li288;output n8097_li289_li289;output n8100_li290_li290;output n8103_li291_li291;output n8106_li292_li292;output n8109_li293_li293;output n8112_li294_li294;output n8115_li295_li295;output n8118_li296_li296;output n8121_li297_li297;output n8124_li298_li298;output n8127_li299_li299;output n8130_li300_li300;output n8133_li301_li301;output n8136_li302_li302;output n8139_li303_li303;output n8142_li304_li304;output n8145_li305_li305;output n8148_li306_li306;output n8151_li307_li307;output n8154_li308_li308;output n8157_li309_li309;output n8160_li310_li310;output n8163_li311_li311;output n8166_li312_li312;output n8169_li313_li313;output n8172_li314_li314;output n8175_li315_li315;output n8178_li316_li316;output n8181_li317_li317;output n8184_li318_li318;output n8187_li319_li319;output n8190_li320_li320;output n8193_li321_li321;output n8196_li322_li322;output n8199_li323_li323;output n8202_li324_li324;output n8205_li325_li325;output n8208_li326_li326;output n8211_li327_li327;output n8214_li328_li328;output n8217_li329_li329;output n8220_li330_li330;output n8223_li331_li331;output n8226_li332_li332;output n8229_li333_li333;output n8232_li334_li334;output n8235_li335_li335;output n8238_li336_li336;output n8241_li337_li337;output n8244_li338_li338;output n8247_li339_li339;output n8250_li340_li340;output n8253_li341_li341;output n8256_li342_li342;output n8259_li343_li343;output n8262_li344_li344;output n8265_li345_li345;output n8268_li346_li346;output n8271_li347_li347;output n8274_li348_li348;output n8286_li352_li352;output n8370_li380_li380;output n8382_li384_li384;output n8394_li388_li388;output n8406_li392_li392;output n8409_li393_li393;output n8412_li394_li394;output n8415_li395_li395;output n8418_li396_li396;output n8430_li400_li400;output n8442_li404_li404;output n8454_li408_li408;output n8466_li412_li412;output n8550_li440_li440;output n8553_li441_li441;output n8556_li442_li442;output n8562_li444_li444;output n8565_li445_li445;output n8568_li446_li446;output n8574_li448_li448;output n8577_li449_li449;output n8583_li451_li451;output n8586_li452_li452;output n8589_li453_li453;output n8595_li455_li455;output n8598_li456_li456;output n8610_li460_li460;output n8670_li480_li480;output n8682_li484_li484;output n8718_li496_li496;output n8727_li499_li499;output n8730_li500_li500;output n8742_li504_li504;output n8751_li507_li507;output n8775_li515_li515;output n8778_li516_li516;output n8790_li520_li520;output n8799_li523_li523;output n8802_li524_li524;output n8805_li525_li525;output n8808_li526_li526;output n8814_li528_li528;output n8817_li529_li529;output n8820_li530_li530;output n8826_li532_li532;output n8829_li533_li533;output n8832_li534_li534;output n8835_li535_li535;output n8850_li540_li540;output n8853_li541_li541;output n8856_li542_li542;output n8859_li543_li543;output n8862_li544_li544;output n8874_li548_li548;output n8910_li560_li560;output n8913_li561_li561;output n8922_li564_li564;output n8934_li568_li568;output n8970_li580_li580;output n8982_li584_li584;output n8994_li588_li588;output n9006_li592_li592;output n9018_li596_li596;output n9030_li600_li600;output n9033_li601_li601;output n9036_li602_li602;output n9039_li603_li603;output n9042_li604_li604;output n9045_li605_li605;output n9048_li606_li606;output n9051_li607_li607;output n9054_li608_li608;output n9057_li609_li609;output n9060_li610_li610;output n9063_li611_li611;output n9066_li612_li612;output n9069_li613_li613;output n9072_li614_li614;output n9075_li615_li615;output n9078_li616_li616;output n9081_li617_li617;output n9084_li618_li618;output n9087_li619_li619;output n9090_li620_li620;output n9093_li621_li621;output n9096_li622_li622;output n9099_li623_li623;output n9102_li624_li624;output n9105_li625_li625;output n9108_li626_li626;output n9114_li628_li628;output n9117_li629_li629;output n9120_li630_li630;output n9123_li631_li631;output n9126_li632_li632;output n9129_li633_li633;output n9132_li634_li634;output n9135_li635_li635;output n9138_li636_li636;output n9141_li637_li637;output n9144_li638_li638;output n9147_li639_li639;output n9150_li640_li640;output n9153_li641_li641;output n9156_li642_li642;output n9159_li643_li643;output n9162_li644_li644;output n9165_li645_li645;output n9174_li648_li648;output n9177_li649_li649;output n9180_li650_li650;output n9183_li651_li651;output n9186_li652_li652;output n9189_li653_li653;output n9192_li654_li654;output n9195_li655_li655;output n9198_li656_li656;output n9201_li657_li657;output n9204_li658_li658;output n9207_li659_li659;output n9210_li660_li660;output n9213_li661_li661;output n9216_li662_li662;output n9222_li664_li664;output n9225_li665_li665;output n9228_li666_li666;output n9234_li668_li668;output n9237_li669_li669;output n9240_li670_li670;output n9246_li672_li672;output n9249_li673_li673;output n9252_li674_li674;output n9258_li676_li676;output n9261_li677_li677;output n9264_li678_li678;output n9267_li679_li679;output n9270_li680_li680;output n9273_li681_li681;output n9276_li682_li682;output n9279_li683_li683;output n9282_li684_li684;output n9285_li685_li685;output n9288_li686_li686;output n9291_li687_li687;output n9294_li688_li688;output n9297_li689_li689;output n9300_li690_li690;output n9303_li691_li691;output n9306_li692_li692;output n9309_li693_li693;output n9312_li694_li694;output n9315_li695_li695;output n9318_li696_li696;output n9321_li697_li697;output n9324_li698_li698;output n9327_li699_li699;output n9330_li700_li700;output n9333_li701_li701;output n9336_li702_li702;output n9339_li703_li703;output n9342_li704_li704;output n9345_li705_li705;output n9348_li706_li706;output n9351_li707_li707;output n9354_li708_li708;output n9357_li709_li709;output n9360_li710_li710;output n9363_li711_li711;output n4970_i2;output n4972_i2;output n4989_i2;output n5024_i2;output n5025_i2;output n5029_i2;output n5042_i2;output n5048_i2;output n5093_i2;output n5096_i2;output n5193_i2;output n5199_i2;output n5203_i2;output n5214_i2;output n5221_i2;output n5222_i2;output n5273_i2;output n5365_i2;output n5385_i2;output n5553_i2;output n5636_i2;output n5782_i2;output n5778_i2;output n5323_i2;output n5325_i2;output n5327_i2;output n5329_i2;output n5816_i2;output n5817_i2;output n5837_i2;output n5844_i2;output n5859_i2;output n5857_i2;output n5369_i2;output n5371_i2;output n5373_i2;output n5400_i2;output n5402_i2;output n5404_i2;output n5406_i2;output n5407_i2;output n5408_i2;output n2722_i2;output n5411_i2;output n5412_i2;output n5413_i2;output n5557_i2;output n5558_i2;output n5559_i2;output n5564_i2;output n5565_i2;output n5561_i2;output n5568_i2;output n5598_i2;output n5600_i2;output n5601_i2;output n5602_i2;output n5603_i2;output n2853_i2;output n5637_i2;output n5627_i2;output n5628_i2;output n5635_i2;output n5640_i2;output n5641_i2;output n5642_i2;output n5650_i2;output n5652_i2;output n5653_i2;output n5654_i2;output n5655_i2;output n5657_i2;output n5659_i2;output n5661_i2;output n5656_i2;output n5663_i2;output n5664_i2;output n5795_i2;output n5796_i2;output n5797_i2;output n5739_i2;output n5773_i2;output n5798_i2;output n5799_i2;output n5802_i2;output n5803_i2;output n5831_i2;output n5833_i2;output n5820_i2;output n5823_i2;output n5824_i2;output n5869_i2;output n5848_i2;output n5849_i2;output n5856_i2;output n5896_i2;output n2754_i2;output n2908_i2;output n5892_i2;output n5915_i2;output n5919_i2;output n5918_i2;output n5920_i2;output n5917_i2;output lo586_buf_i2;output n2818_i2;output n2863_i2;output n2721_i2;output n2725_i2;output n3016_i2;output n3013_i2;output n2655_i2;output n2741_i2;output lo562_buf_i2;output n2656_i2;output n2531_i2;output n2700_i2;output n5908_i2;output n5910_i2;output n5912_i2;output n5914_i2;output n2753_i2;output n2878_i2;output n2836_i2;output n5934_i2;output n5936_i2;output n5938_i2;output n2728_i2;output lo358_buf_i2;output lo418_buf_i2;output lo474_buf_i2;output lo554_buf_i2;output lo558_buf_i2;output lo574_buf_i2;output n2659_i2;output n2665_i2;output n2686_i2;output lo450_buf_i2;output n2910_i2;output n2683_i2;output n2828_i2;output n2582_i2;output n2600_i2;output n2542_i2;output n2703_i2;output lo510_buf_i2;output lo514_buf_i2;output lo538_buf_i2;output lo578_buf_i2;output n2692_i2;output n2666_i2;output n2667_i2;output n2660_i2;output n2744_i2;output lo454_buf_i2;output n3593_i2;output n3048_i2;output lo410_buf_i2;output lo502_buf_i2;output lo506_buf_i2;output lo550_buf_i2;output lo570_buf_i2;output lo582_buf_i2;output n2646_i2;output n2673_i2;output n3499_i2;output n2750_i2;output n2870_i2;output n2693_i2;output n2689_i2;output n2668_i2;output n2662_i2;output lo350_buf_i2;output lo498_buf_i2;output lo518_buf_i2;output lo522_buf_i2;output lo598_buf_i2;output n2708_i2;output n2674_i2;output n2647_i2;output n2751_i2;output n2747_i2;output n2669_i2;output n2872_i2;output n3313_i2;output n3273_i2;output n2848_i2;output n2893_i2;output n3267_i2;output n2925_i2;output n2839_i2;output n2831_i2;output n2558_i2;output n2562_i2;output n2825_i2;output n3263_i2;output n3517_i2;output n2873_i2;output n2926_i2;output n3261_i2;output n3268_i2;output n3274_i2;output n3314_i2;output n3571_i2;output n2950_i2;output n2951_i2;output n3022_i2;output n3023_i2;output n3057_i2;output n3058_i2;output n2931_i2;output n2911_i2;output n2959_i2;output n2960_i2;output n2922_i2;output n2888_i2;output n2889_i2;output n3051_i2;output n3052_i2;output n3063_i2;output n2845_i2;output n2737_i2;output n3281_i2;output n3294_i2;output n2885_i2;output n2786_i2;output n2783_i2;output n2801_i2;output n2572_i2;output n2628_i2;output n2609_i2;output n2618_i2;output n2637_i2;output n2525_i2;output n2551_i2;output n3759_i2;output n2994_i2;output n3040_i2;output n2943_i2;output n2991_i2;output n3034_i2;output n2881_i2;output n3021_i2;output n3062_i2;output n2763_i2;output n2764_i2;output n2775_i2;output n2776_i2;output n2968_i2;output n2969_i2;output n2798_i2;output n3661_i2;output n2694_i2;output n2809_i2;output n2817_i2;output n2514_i2;output n2501_i2;output n2528_i2;output n2505_i2;output n2492_i2;output lo546_buf_i2;output lo590_buf_i2;output lo594_buf_i2;output n2679_i2;output n2733_i2;output n2709_i2;output n2676_i2;output n2649_i2;output n2815_i2;output n2704_i2;output n3590_i2;output n3591_i2;output n2752_i2;output n3638_i2;output n3639_i2;output n2695_i2;output n3047_i2;output lo458_buf_i2;output lo482_buf_i2;output lo566_buf_i2;output n2718_i2;output n3707_i2;output n3671_i2;output n3680_i2;output n3749_i2;output n3716_i2;output n3692_i2;output n2591_i2;output n3478_i2;output n3610_i2;output n3611_i2;output n2652_i2;output n2714_i2;output n2738_i2;output n3616_i2;output n3617_i2;output n3031_i2;output n2515_i2;output n3562_i2;output n2502_i2;output n3560_i2;output n3554_i2;output n3555_i2;output n3536_i2;output n3537_i2;output n3508_i2;output n3650_i2;output n3740_i2;output n3484_i2;output n2680_i2;output n2734_i2;output n2735_i2;output n2711_i2;output lo585_buf_i2;output n2719_i2;output n2720_i2;output n2723_i2;output n2724_i2;output n3624_i2;output n3625_i2;output n3015_i2;output n3491_i2;output n2696_i2;output n2811_i2;output n3010_i2;output n3012_i2;output lo382_buf_i2;output lo386_buf_i2;output lo390_buf_i2;output lo398_buf_i2;output lo402_buf_i2;output lo406_buf_i2;output n3492_i2;output lo366_buf_i2;output lo374_buf_i2;output lo426_buf_i2;output lo494_buf_i2;output n2653_i2;output n2654_i2;output n2715_i2;output n2740_i2;output n2682_i2;output n2736_i2;output lo508_buf_i2;output lo512_buf_i2;output lo536_buf_i2;output lo576_buf_i2;output lo357_buf_i2;output lo361_buf_i2;output lo417_buf_i2;output lo421_buf_i2;output lo473_buf_i2;output lo477_buf_i2;output lo553_buf_i2;output lo557_buf_i2;output lo573_buf_i2;output lo434_buf_i2;output lo438_buf_i2;output lo466_buf_i2;output lo470_buf_i2;output lo490_buf_i2;output n2657_i2;output n2658_i2;output n2663_i2;output n2664_i2;output n2684_i2;output n2685_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire G51_p;
  wire G51_n;
  wire G52_p;
  wire G52_n;
  wire G53_p;
  wire G53_n;
  wire G54_p;
  wire G54_n;
  wire G55_p;
  wire G55_n;
  wire G56_p;
  wire G56_n;
  wire G57_p;
  wire G57_n;
  wire G58_p;
  wire G58_n;
  wire G59_p;
  wire G59_n;
  wire G60_p;
  wire G60_n;
  wire G61_p;
  wire G61_n;
  wire G62_p;
  wire G62_n;
  wire G63_p;
  wire G63_n;
  wire G64_p;
  wire G64_n;
  wire G65_p;
  wire G65_n;
  wire G66_p;
  wire G66_n;
  wire G67_p;
  wire G67_n;
  wire G68_p;
  wire G68_n;
  wire G69_p;
  wire G69_n;
  wire G70_p;
  wire G70_n;
  wire G71_p;
  wire G71_n;
  wire G72_p;
  wire G72_n;
  wire G73_p;
  wire G73_n;
  wire G74_p;
  wire G74_n;
  wire G75_p;
  wire G75_n;
  wire G76_p;
  wire G76_n;
  wire G77_p;
  wire G77_n;
  wire G78_p;
  wire G78_n;
  wire G79_p;
  wire G79_n;
  wire G80_p;
  wire G80_n;
  wire G81_p;
  wire G81_n;
  wire G82_p;
  wire G82_n;
  wire G83_p;
  wire G83_n;
  wire G84_p;
  wire G84_n;
  wire G85_p;
  wire G85_n;
  wire G86_p;
  wire G86_n;
  wire G87_p;
  wire G87_n;
  wire G88_p;
  wire G88_n;
  wire G89_p;
  wire G89_n;
  wire G90_p;
  wire G90_n;
  wire G91_p;
  wire G91_n;
  wire G92_p;
  wire G92_n;
  wire G93_p;
  wire G93_n;
  wire G94_p;
  wire G94_n;
  wire G95_p;
  wire G95_n;
  wire G96_p;
  wire G96_n;
  wire G97_p;
  wire G97_n;
  wire G98_p;
  wire G98_n;
  wire G99_p;
  wire G99_n;
  wire G100_p;
  wire G100_n;
  wire G101_p;
  wire G101_n;
  wire G102_p;
  wire G102_n;
  wire G103_p;
  wire G103_n;
  wire G104_p;
  wire G104_n;
  wire G105_p;
  wire G105_n;
  wire G106_p;
  wire G106_n;
  wire G107_p;
  wire G107_n;
  wire G108_p;
  wire G108_n;
  wire G109_p;
  wire G109_n;
  wire G110_p;
  wire G110_n;
  wire G111_p;
  wire G111_n;
  wire G112_p;
  wire G112_n;
  wire G113_p;
  wire G113_n;
  wire G114_p;
  wire G114_n;
  wire G115_p;
  wire G115_n;
  wire G116_p;
  wire G116_n;
  wire G117_p;
  wire G117_n;
  wire G118_p;
  wire G118_n;
  wire G119_p;
  wire G119_n;
  wire G120_p;
  wire G120_n;
  wire G121_p;
  wire G121_n;
  wire G122_p;
  wire G122_n;
  wire G123_p;
  wire G123_n;
  wire G124_p;
  wire G124_n;
  wire G125_p;
  wire G125_n;
  wire G126_p;
  wire G126_n;
  wire G127_p;
  wire G127_n;
  wire G128_p;
  wire G128_n;
  wire G129_p;
  wire G129_n;
  wire G130_p;
  wire G130_n;
  wire G131_p;
  wire G131_n;
  wire G132_p;
  wire G132_n;
  wire G133_p;
  wire G133_n;
  wire G134_p;
  wire G134_n;
  wire G135_p;
  wire G135_n;
  wire G136_p;
  wire G136_n;
  wire G137_p;
  wire G137_n;
  wire G138_p;
  wire G138_n;
  wire G139_p;
  wire G139_n;
  wire G140_p;
  wire G140_n;
  wire G141_p;
  wire G141_n;
  wire G142_p;
  wire G142_n;
  wire G143_p;
  wire G143_n;
  wire G144_p;
  wire G144_n;
  wire G145_p;
  wire G145_n;
  wire G146_p;
  wire G146_n;
  wire G147_p;
  wire G147_n;
  wire G148_p;
  wire G148_n;
  wire G149_p;
  wire G149_n;
  wire G150_p;
  wire G150_n;
  wire G151_p;
  wire G151_n;
  wire G152_p;
  wire G152_n;
  wire G153_p;
  wire G153_n;
  wire G154_p;
  wire G154_n;
  wire G155_p;
  wire G155_n;
  wire G156_p;
  wire G156_n;
  wire G157_p;
  wire G157_n;
  wire G158_p;
  wire G158_n;
  wire G159_p;
  wire G159_n;
  wire G160_p;
  wire G160_n;
  wire G161_p;
  wire G161_n;
  wire G162_p;
  wire G162_n;
  wire G163_p;
  wire G163_n;
  wire G164_p;
  wire G164_n;
  wire G165_p;
  wire G165_n;
  wire G166_p;
  wire G166_n;
  wire G167_p;
  wire G167_n;
  wire G168_p;
  wire G168_n;
  wire G169_p;
  wire G169_n;
  wire G170_p;
  wire G170_n;
  wire G171_p;
  wire G171_n;
  wire G172_p;
  wire G172_n;
  wire G173_p;
  wire G173_n;
  wire G174_p;
  wire G174_n;
  wire G175_p;
  wire G175_n;
  wire G176_p;
  wire G176_n;
  wire G177_p;
  wire G177_n;
  wire G178_p;
  wire G178_n;
  wire n2610_lo_p;
  wire n2610_lo_n;
  wire n2613_lo_p;
  wire n2613_lo_n;
  wire n2616_lo_p;
  wire n2616_lo_n;
  wire n2619_lo_p;
  wire n2619_lo_n;
  wire n2622_lo_p;
  wire n2622_lo_n;
  wire n2625_lo_p;
  wire n2625_lo_n;
  wire n2628_lo_p;
  wire n2628_lo_n;
  wire n2634_lo_p;
  wire n2634_lo_n;
  wire n2637_lo_p;
  wire n2637_lo_n;
  wire n2640_lo_p;
  wire n2640_lo_n;
  wire n2643_lo_p;
  wire n2643_lo_n;
  wire n2646_lo_p;
  wire n2646_lo_n;
  wire n2649_lo_p;
  wire n2649_lo_n;
  wire n2652_lo_p;
  wire n2652_lo_n;
  wire n2655_lo_p;
  wire n2655_lo_n;
  wire n2658_lo_p;
  wire n2658_lo_n;
  wire n2661_lo_p;
  wire n2661_lo_n;
  wire n2664_lo_p;
  wire n2664_lo_n;
  wire n2667_lo_p;
  wire n2667_lo_n;
  wire n2670_lo_p;
  wire n2670_lo_n;
  wire n2673_lo_p;
  wire n2673_lo_n;
  wire n2676_lo_p;
  wire n2676_lo_n;
  wire n2679_lo_p;
  wire n2679_lo_n;
  wire n2682_lo_p;
  wire n2682_lo_n;
  wire n2685_lo_p;
  wire n2685_lo_n;
  wire n2688_lo_p;
  wire n2688_lo_n;
  wire n2691_lo_p;
  wire n2691_lo_n;
  wire n2694_lo_p;
  wire n2694_lo_n;
  wire n2697_lo_p;
  wire n2697_lo_n;
  wire n2700_lo_p;
  wire n2700_lo_n;
  wire n2703_lo_p;
  wire n2703_lo_n;
  wire n2706_lo_p;
  wire n2706_lo_n;
  wire n2709_lo_p;
  wire n2709_lo_n;
  wire n2712_lo_p;
  wire n2712_lo_n;
  wire n2715_lo_p;
  wire n2715_lo_n;
  wire n2718_lo_p;
  wire n2718_lo_n;
  wire n2721_lo_p;
  wire n2721_lo_n;
  wire n2724_lo_p;
  wire n2724_lo_n;
  wire n2727_lo_p;
  wire n2727_lo_n;
  wire n2730_lo_p;
  wire n2730_lo_n;
  wire n2733_lo_p;
  wire n2733_lo_n;
  wire n2736_lo_p;
  wire n2736_lo_n;
  wire n2739_lo_p;
  wire n2739_lo_n;
  wire n2742_lo_p;
  wire n2742_lo_n;
  wire n2745_lo_p;
  wire n2745_lo_n;
  wire n2748_lo_p;
  wire n2748_lo_n;
  wire n2751_lo_p;
  wire n2751_lo_n;
  wire n2754_lo_p;
  wire n2754_lo_n;
  wire n2757_lo_p;
  wire n2757_lo_n;
  wire n2760_lo_p;
  wire n2760_lo_n;
  wire n2763_lo_p;
  wire n2763_lo_n;
  wire n2766_lo_p;
  wire n2766_lo_n;
  wire n2769_lo_p;
  wire n2769_lo_n;
  wire n2772_lo_p;
  wire n2772_lo_n;
  wire n2775_lo_p;
  wire n2775_lo_n;
  wire n2778_lo_p;
  wire n2778_lo_n;
  wire n2781_lo_p;
  wire n2781_lo_n;
  wire n2784_lo_p;
  wire n2784_lo_n;
  wire n2787_lo_p;
  wire n2787_lo_n;
  wire n2790_lo_p;
  wire n2790_lo_n;
  wire n2793_lo_p;
  wire n2793_lo_n;
  wire n2796_lo_p;
  wire n2796_lo_n;
  wire n2799_lo_p;
  wire n2799_lo_n;
  wire n2802_lo_p;
  wire n2802_lo_n;
  wire n2805_lo_p;
  wire n2805_lo_n;
  wire n2808_lo_p;
  wire n2808_lo_n;
  wire n2811_lo_p;
  wire n2811_lo_n;
  wire n2814_lo_p;
  wire n2814_lo_n;
  wire n2817_lo_p;
  wire n2817_lo_n;
  wire n2820_lo_p;
  wire n2820_lo_n;
  wire n2823_lo_p;
  wire n2823_lo_n;
  wire n2826_lo_p;
  wire n2826_lo_n;
  wire n2829_lo_p;
  wire n2829_lo_n;
  wire n2832_lo_p;
  wire n2832_lo_n;
  wire n2838_lo_p;
  wire n2838_lo_n;
  wire n2841_lo_p;
  wire n2841_lo_n;
  wire n2844_lo_p;
  wire n2844_lo_n;
  wire n2847_lo_p;
  wire n2847_lo_n;
  wire n2850_lo_p;
  wire n2850_lo_n;
  wire n2853_lo_p;
  wire n2853_lo_n;
  wire n2856_lo_p;
  wire n2856_lo_n;
  wire n2862_lo_p;
  wire n2862_lo_n;
  wire n2865_lo_p;
  wire n2865_lo_n;
  wire n2868_lo_p;
  wire n2868_lo_n;
  wire n2871_lo_p;
  wire n2871_lo_n;
  wire n2874_lo_p;
  wire n2874_lo_n;
  wire n2877_lo_p;
  wire n2877_lo_n;
  wire n2880_lo_p;
  wire n2880_lo_n;
  wire n2883_lo_p;
  wire n2883_lo_n;
  wire n2886_lo_p;
  wire n2886_lo_n;
  wire n2889_lo_p;
  wire n2889_lo_n;
  wire n2892_lo_p;
  wire n2892_lo_n;
  wire n2895_lo_p;
  wire n2895_lo_n;
  wire n2898_lo_p;
  wire n2898_lo_n;
  wire n2901_lo_p;
  wire n2901_lo_n;
  wire n2904_lo_p;
  wire n2904_lo_n;
  wire n2907_lo_p;
  wire n2907_lo_n;
  wire n2910_lo_p;
  wire n2910_lo_n;
  wire n2913_lo_p;
  wire n2913_lo_n;
  wire n2916_lo_p;
  wire n2916_lo_n;
  wire n2919_lo_p;
  wire n2919_lo_n;
  wire n2922_lo_p;
  wire n2922_lo_n;
  wire n2925_lo_p;
  wire n2925_lo_n;
  wire n2928_lo_p;
  wire n2928_lo_n;
  wire n2931_lo_p;
  wire n2931_lo_n;
  wire n2934_lo_p;
  wire n2934_lo_n;
  wire n2937_lo_p;
  wire n2937_lo_n;
  wire n2940_lo_p;
  wire n2940_lo_n;
  wire n2943_lo_p;
  wire n2943_lo_n;
  wire n2946_lo_p;
  wire n2946_lo_n;
  wire n2949_lo_p;
  wire n2949_lo_n;
  wire n2952_lo_p;
  wire n2952_lo_n;
  wire n2955_lo_p;
  wire n2955_lo_n;
  wire n2958_lo_p;
  wire n2958_lo_n;
  wire n2961_lo_p;
  wire n2961_lo_n;
  wire n2964_lo_p;
  wire n2964_lo_n;
  wire n2967_lo_p;
  wire n2967_lo_n;
  wire n2970_lo_p;
  wire n2970_lo_n;
  wire n2973_lo_p;
  wire n2973_lo_n;
  wire n2976_lo_p;
  wire n2976_lo_n;
  wire n2979_lo_p;
  wire n2979_lo_n;
  wire n2982_lo_p;
  wire n2982_lo_n;
  wire n2985_lo_p;
  wire n2985_lo_n;
  wire n2988_lo_p;
  wire n2988_lo_n;
  wire n2991_lo_p;
  wire n2991_lo_n;
  wire n2994_lo_p;
  wire n2994_lo_n;
  wire n2997_lo_p;
  wire n2997_lo_n;
  wire n3000_lo_p;
  wire n3000_lo_n;
  wire n3003_lo_p;
  wire n3003_lo_n;
  wire n3006_lo_p;
  wire n3006_lo_n;
  wire n3009_lo_p;
  wire n3009_lo_n;
  wire n3012_lo_p;
  wire n3012_lo_n;
  wire n3015_lo_p;
  wire n3015_lo_n;
  wire n3018_lo_p;
  wire n3018_lo_n;
  wire n3021_lo_p;
  wire n3021_lo_n;
  wire n3024_lo_p;
  wire n3024_lo_n;
  wire n3027_lo_p;
  wire n3027_lo_n;
  wire n3030_lo_p;
  wire n3030_lo_n;
  wire n3033_lo_p;
  wire n3033_lo_n;
  wire n3036_lo_p;
  wire n3036_lo_n;
  wire n3039_lo_p;
  wire n3039_lo_n;
  wire n3042_lo_p;
  wire n3042_lo_n;
  wire n3045_lo_p;
  wire n3045_lo_n;
  wire n3048_lo_p;
  wire n3048_lo_n;
  wire n3051_lo_p;
  wire n3051_lo_n;
  wire n3054_lo_p;
  wire n3054_lo_n;
  wire n3057_lo_p;
  wire n3057_lo_n;
  wire n3060_lo_p;
  wire n3060_lo_n;
  wire n3063_lo_p;
  wire n3063_lo_n;
  wire n3066_lo_p;
  wire n3066_lo_n;
  wire n3069_lo_p;
  wire n3069_lo_n;
  wire n3072_lo_p;
  wire n3072_lo_n;
  wire n3075_lo_p;
  wire n3075_lo_n;
  wire n3078_lo_p;
  wire n3078_lo_n;
  wire n3081_lo_p;
  wire n3081_lo_n;
  wire n3084_lo_p;
  wire n3084_lo_n;
  wire n3087_lo_p;
  wire n3087_lo_n;
  wire n3090_lo_p;
  wire n3090_lo_n;
  wire n3093_lo_p;
  wire n3093_lo_n;
  wire n3096_lo_p;
  wire n3096_lo_n;
  wire n3099_lo_p;
  wire n3099_lo_n;
  wire n3102_lo_p;
  wire n3102_lo_n;
  wire n3105_lo_p;
  wire n3105_lo_n;
  wire n3108_lo_p;
  wire n3108_lo_n;
  wire n3111_lo_p;
  wire n3111_lo_n;
  wire n3114_lo_p;
  wire n3114_lo_n;
  wire n3117_lo_p;
  wire n3117_lo_n;
  wire n3120_lo_p;
  wire n3120_lo_n;
  wire n3126_lo_p;
  wire n3126_lo_n;
  wire n3129_lo_p;
  wire n3129_lo_n;
  wire n3132_lo_p;
  wire n3132_lo_n;
  wire n3138_lo_p;
  wire n3138_lo_n;
  wire n3141_lo_p;
  wire n3141_lo_n;
  wire n3144_lo_p;
  wire n3144_lo_n;
  wire n3147_lo_p;
  wire n3147_lo_n;
  wire n3150_lo_p;
  wire n3150_lo_n;
  wire n3153_lo_p;
  wire n3153_lo_n;
  wire n3156_lo_p;
  wire n3156_lo_n;
  wire n3162_lo_p;
  wire n3162_lo_n;
  wire n3165_lo_p;
  wire n3165_lo_n;
  wire n3168_lo_p;
  wire n3168_lo_n;
  wire n3174_lo_p;
  wire n3174_lo_n;
  wire n3177_lo_p;
  wire n3177_lo_n;
  wire n3180_lo_p;
  wire n3180_lo_n;
  wire n3186_lo_p;
  wire n3186_lo_n;
  wire n3189_lo_p;
  wire n3189_lo_n;
  wire n3192_lo_p;
  wire n3192_lo_n;
  wire n3195_lo_p;
  wire n3195_lo_n;
  wire n3198_lo_p;
  wire n3198_lo_n;
  wire n3201_lo_p;
  wire n3201_lo_n;
  wire n3204_lo_p;
  wire n3204_lo_n;
  wire n3210_lo_p;
  wire n3210_lo_n;
  wire n3213_lo_p;
  wire n3213_lo_n;
  wire n3216_lo_p;
  wire n3216_lo_n;
  wire n3219_lo_p;
  wire n3219_lo_n;
  wire n3222_lo_p;
  wire n3222_lo_n;
  wire n3225_lo_p;
  wire n3225_lo_n;
  wire n3228_lo_p;
  wire n3228_lo_n;
  wire n3234_lo_p;
  wire n3234_lo_n;
  wire n3237_lo_p;
  wire n3237_lo_n;
  wire n3240_lo_p;
  wire n3240_lo_n;
  wire n3243_lo_p;
  wire n3243_lo_n;
  wire n3246_lo_p;
  wire n3246_lo_n;
  wire n3249_lo_p;
  wire n3249_lo_n;
  wire n3252_lo_p;
  wire n3252_lo_n;
  wire n3255_lo_p;
  wire n3255_lo_n;
  wire n3258_lo_p;
  wire n3258_lo_n;
  wire n3261_lo_p;
  wire n3261_lo_n;
  wire n3264_lo_p;
  wire n3264_lo_n;
  wire n3267_lo_p;
  wire n3267_lo_n;
  wire n3270_lo_p;
  wire n3270_lo_n;
  wire n3273_lo_p;
  wire n3273_lo_n;
  wire n3276_lo_p;
  wire n3276_lo_n;
  wire n3279_lo_p;
  wire n3279_lo_n;
  wire n3282_lo_p;
  wire n3282_lo_n;
  wire n3285_lo_p;
  wire n3285_lo_n;
  wire n3288_lo_p;
  wire n3288_lo_n;
  wire n3294_lo_p;
  wire n3294_lo_n;
  wire n3297_lo_p;
  wire n3297_lo_n;
  wire n3300_lo_p;
  wire n3300_lo_n;
  wire n3306_lo_p;
  wire n3306_lo_n;
  wire n3309_lo_p;
  wire n3309_lo_n;
  wire n3312_lo_p;
  wire n3312_lo_n;
  wire n3318_lo_p;
  wire n3318_lo_n;
  wire n3321_lo_p;
  wire n3321_lo_n;
  wire n3324_lo_p;
  wire n3324_lo_n;
  wire n3330_lo_p;
  wire n3330_lo_n;
  wire n3333_lo_p;
  wire n3333_lo_n;
  wire n3336_lo_p;
  wire n3336_lo_n;
  wire n3339_lo_p;
  wire n3339_lo_n;
  wire n3342_lo_p;
  wire n3342_lo_n;
  wire n3345_lo_p;
  wire n3345_lo_n;
  wire n3348_lo_p;
  wire n3348_lo_n;
  wire n3351_lo_p;
  wire n3351_lo_n;
  wire n3354_lo_p;
  wire n3354_lo_n;
  wire n3357_lo_p;
  wire n3357_lo_n;
  wire n3360_lo_p;
  wire n3360_lo_n;
  wire n3363_lo_p;
  wire n3363_lo_n;
  wire n3366_lo_p;
  wire n3366_lo_n;
  wire n3369_lo_p;
  wire n3369_lo_n;
  wire n3372_lo_p;
  wire n3372_lo_n;
  wire n3375_lo_p;
  wire n3375_lo_n;
  wire n3378_lo_p;
  wire n3378_lo_n;
  wire n3381_lo_p;
  wire n3381_lo_n;
  wire n3384_lo_p;
  wire n3384_lo_n;
  wire n3387_lo_p;
  wire n3387_lo_n;
  wire n3390_lo_p;
  wire n3390_lo_n;
  wire n3393_lo_p;
  wire n3393_lo_n;
  wire n3396_lo_p;
  wire n3396_lo_n;
  wire n3399_lo_p;
  wire n3399_lo_n;
  wire n3402_lo_p;
  wire n3402_lo_n;
  wire n3405_lo_p;
  wire n3405_lo_n;
  wire n3408_lo_p;
  wire n3408_lo_n;
  wire n3411_lo_p;
  wire n3411_lo_n;
  wire n3414_lo_p;
  wire n3414_lo_n;
  wire n3417_lo_p;
  wire n3417_lo_n;
  wire n3420_lo_p;
  wire n3420_lo_n;
  wire n3423_lo_p;
  wire n3423_lo_n;
  wire n3426_lo_p;
  wire n3426_lo_n;
  wire n3429_lo_p;
  wire n3429_lo_n;
  wire n3432_lo_p;
  wire n3432_lo_n;
  wire n3435_lo_p;
  wire n3435_lo_n;
  wire n3438_lo_p;
  wire n3438_lo_n;
  wire n3441_lo_p;
  wire n3441_lo_n;
  wire n3444_lo_p;
  wire n3444_lo_n;
  wire n3447_lo_p;
  wire n3447_lo_n;
  wire n3450_lo_p;
  wire n3450_lo_n;
  wire n3453_lo_p;
  wire n3453_lo_n;
  wire n3456_lo_p;
  wire n3456_lo_n;
  wire n3459_lo_p;
  wire n3459_lo_n;
  wire n3462_lo_p;
  wire n3462_lo_n;
  wire n3465_lo_p;
  wire n3465_lo_n;
  wire n3468_lo_p;
  wire n3468_lo_n;
  wire n3471_lo_p;
  wire n3471_lo_n;
  wire n3474_lo_p;
  wire n3474_lo_n;
  wire n3477_lo_p;
  wire n3477_lo_n;
  wire n3480_lo_p;
  wire n3480_lo_n;
  wire n3483_lo_p;
  wire n3483_lo_n;
  wire n3486_lo_p;
  wire n3486_lo_n;
  wire n3489_lo_p;
  wire n3489_lo_n;
  wire n3492_lo_p;
  wire n3492_lo_n;
  wire n3495_lo_p;
  wire n3495_lo_n;
  wire n3498_lo_p;
  wire n3498_lo_n;
  wire n3501_lo_p;
  wire n3501_lo_n;
  wire n3504_lo_p;
  wire n3504_lo_n;
  wire n3507_lo_p;
  wire n3507_lo_n;
  wire n3510_lo_p;
  wire n3510_lo_n;
  wire n3513_lo_p;
  wire n3513_lo_n;
  wire n3516_lo_p;
  wire n3516_lo_n;
  wire n3519_lo_p;
  wire n3519_lo_n;
  wire n3522_lo_p;
  wire n3522_lo_n;
  wire n3525_lo_p;
  wire n3525_lo_n;
  wire n3528_lo_p;
  wire n3528_lo_n;
  wire n3531_lo_p;
  wire n3531_lo_n;
  wire n3534_lo_p;
  wire n3534_lo_n;
  wire n3537_lo_p;
  wire n3537_lo_n;
  wire n3540_lo_p;
  wire n3540_lo_n;
  wire n3543_lo_p;
  wire n3543_lo_n;
  wire n3546_lo_p;
  wire n3546_lo_n;
  wire n3549_lo_p;
  wire n3549_lo_n;
  wire n3552_lo_p;
  wire n3552_lo_n;
  wire n3555_lo_p;
  wire n3555_lo_n;
  wire n3558_lo_p;
  wire n3558_lo_n;
  wire n3561_lo_p;
  wire n3561_lo_n;
  wire n3564_lo_p;
  wire n3564_lo_n;
  wire n3567_lo_p;
  wire n3567_lo_n;
  wire n3570_lo_p;
  wire n3570_lo_n;
  wire n3573_lo_p;
  wire n3573_lo_n;
  wire n3576_lo_p;
  wire n3576_lo_n;
  wire n3579_lo_p;
  wire n3579_lo_n;
  wire n3582_lo_p;
  wire n3582_lo_n;
  wire n3585_lo_p;
  wire n3585_lo_n;
  wire n3588_lo_p;
  wire n3588_lo_n;
  wire n3591_lo_p;
  wire n3591_lo_n;
  wire n3594_lo_p;
  wire n3594_lo_n;
  wire n3597_lo_p;
  wire n3597_lo_n;
  wire n3600_lo_p;
  wire n3600_lo_n;
  wire n3603_lo_p;
  wire n3603_lo_n;
  wire n3606_lo_p;
  wire n3606_lo_n;
  wire n3609_lo_p;
  wire n3609_lo_n;
  wire n3612_lo_p;
  wire n3612_lo_n;
  wire n3615_lo_p;
  wire n3615_lo_n;
  wire n3618_lo_p;
  wire n3618_lo_n;
  wire n3621_lo_p;
  wire n3621_lo_n;
  wire n3624_lo_p;
  wire n3624_lo_n;
  wire n3627_lo_p;
  wire n3627_lo_n;
  wire n3630_lo_p;
  wire n3630_lo_n;
  wire n3633_lo_p;
  wire n3633_lo_n;
  wire n3636_lo_p;
  wire n3636_lo_n;
  wire n3639_lo_p;
  wire n3639_lo_n;
  wire n3642_lo_p;
  wire n3642_lo_n;
  wire n3645_lo_p;
  wire n3645_lo_n;
  wire n3648_lo_p;
  wire n3648_lo_n;
  wire n3651_lo_p;
  wire n3651_lo_n;
  wire n3654_lo_p;
  wire n3654_lo_n;
  wire n3666_lo_p;
  wire n3666_lo_n;
  wire n3750_lo_p;
  wire n3750_lo_n;
  wire n3762_lo_p;
  wire n3762_lo_n;
  wire n3774_lo_p;
  wire n3774_lo_n;
  wire n3786_lo_p;
  wire n3786_lo_n;
  wire n3789_lo_p;
  wire n3789_lo_n;
  wire n3792_lo_p;
  wire n3792_lo_n;
  wire n3795_lo_p;
  wire n3795_lo_n;
  wire n3798_lo_p;
  wire n3798_lo_n;
  wire n3810_lo_p;
  wire n3810_lo_n;
  wire n3822_lo_p;
  wire n3822_lo_n;
  wire n3834_lo_p;
  wire n3834_lo_n;
  wire n3846_lo_p;
  wire n3846_lo_n;
  wire n3930_lo_p;
  wire n3930_lo_n;
  wire n3933_lo_p;
  wire n3933_lo_n;
  wire n3936_lo_p;
  wire n3936_lo_n;
  wire n3942_lo_p;
  wire n3942_lo_n;
  wire n3945_lo_p;
  wire n3945_lo_n;
  wire n3948_lo_p;
  wire n3948_lo_n;
  wire n3954_lo_p;
  wire n3954_lo_n;
  wire n3957_lo_p;
  wire n3957_lo_n;
  wire n3963_lo_p;
  wire n3963_lo_n;
  wire n3966_lo_p;
  wire n3966_lo_n;
  wire n3969_lo_p;
  wire n3969_lo_n;
  wire n3975_lo_p;
  wire n3975_lo_n;
  wire n3978_lo_p;
  wire n3978_lo_n;
  wire n3990_lo_p;
  wire n3990_lo_n;
  wire n4050_lo_p;
  wire n4050_lo_n;
  wire n4062_lo_p;
  wire n4062_lo_n;
  wire n4098_lo_p;
  wire n4098_lo_n;
  wire n4107_lo_p;
  wire n4107_lo_n;
  wire n4110_lo_p;
  wire n4110_lo_n;
  wire n4122_lo_p;
  wire n4122_lo_n;
  wire n4131_lo_p;
  wire n4131_lo_n;
  wire n4155_lo_p;
  wire n4155_lo_n;
  wire n4158_lo_p;
  wire n4158_lo_n;
  wire n4170_lo_p;
  wire n4170_lo_n;
  wire n4179_lo_p;
  wire n4179_lo_n;
  wire n4182_lo_p;
  wire n4182_lo_n;
  wire n4185_lo_p;
  wire n4185_lo_n;
  wire n4188_lo_p;
  wire n4188_lo_n;
  wire n4194_lo_p;
  wire n4194_lo_n;
  wire n4197_lo_p;
  wire n4197_lo_n;
  wire n4200_lo_p;
  wire n4200_lo_n;
  wire n4206_lo_p;
  wire n4206_lo_n;
  wire n4209_lo_p;
  wire n4209_lo_n;
  wire n4212_lo_p;
  wire n4212_lo_n;
  wire n4215_lo_p;
  wire n4215_lo_n;
  wire n4230_lo_p;
  wire n4230_lo_n;
  wire n4233_lo_p;
  wire n4233_lo_n;
  wire n4236_lo_p;
  wire n4236_lo_n;
  wire n4239_lo_p;
  wire n4239_lo_n;
  wire n4242_lo_p;
  wire n4242_lo_n;
  wire n4254_lo_p;
  wire n4254_lo_n;
  wire n4290_lo_p;
  wire n4290_lo_n;
  wire n4293_lo_p;
  wire n4293_lo_n;
  wire n4302_lo_p;
  wire n4302_lo_n;
  wire n4314_lo_p;
  wire n4314_lo_n;
  wire n4350_lo_p;
  wire n4350_lo_n;
  wire n4362_lo_p;
  wire n4362_lo_n;
  wire n4374_lo_p;
  wire n4374_lo_n;
  wire n4386_lo_p;
  wire n4386_lo_n;
  wire n4398_lo_p;
  wire n4398_lo_n;
  wire n4410_lo_p;
  wire n4410_lo_n;
  wire n4413_lo_p;
  wire n4413_lo_n;
  wire n4416_lo_p;
  wire n4416_lo_n;
  wire n4419_lo_p;
  wire n4419_lo_n;
  wire n4422_lo_p;
  wire n4422_lo_n;
  wire n4425_lo_p;
  wire n4425_lo_n;
  wire n4428_lo_p;
  wire n4428_lo_n;
  wire n4431_lo_p;
  wire n4431_lo_n;
  wire n4434_lo_p;
  wire n4434_lo_n;
  wire n4437_lo_p;
  wire n4437_lo_n;
  wire n4440_lo_p;
  wire n4440_lo_n;
  wire n4443_lo_p;
  wire n4443_lo_n;
  wire n4446_lo_p;
  wire n4446_lo_n;
  wire n4449_lo_p;
  wire n4449_lo_n;
  wire n4452_lo_p;
  wire n4452_lo_n;
  wire n4455_lo_p;
  wire n4455_lo_n;
  wire n4458_lo_p;
  wire n4458_lo_n;
  wire n4461_lo_p;
  wire n4461_lo_n;
  wire n4464_lo_p;
  wire n4464_lo_n;
  wire n4467_lo_p;
  wire n4467_lo_n;
  wire n4470_lo_p;
  wire n4470_lo_n;
  wire n4473_lo_p;
  wire n4473_lo_n;
  wire n4476_lo_p;
  wire n4476_lo_n;
  wire n4479_lo_p;
  wire n4479_lo_n;
  wire n4482_lo_p;
  wire n4482_lo_n;
  wire n4485_lo_p;
  wire n4485_lo_n;
  wire n4488_lo_p;
  wire n4488_lo_n;
  wire n4494_lo_p;
  wire n4494_lo_n;
  wire n4497_lo_p;
  wire n4497_lo_n;
  wire n4500_lo_p;
  wire n4500_lo_n;
  wire n4503_lo_p;
  wire n4503_lo_n;
  wire n4506_lo_p;
  wire n4506_lo_n;
  wire n4509_lo_p;
  wire n4509_lo_n;
  wire n4512_lo_p;
  wire n4512_lo_n;
  wire n4515_lo_p;
  wire n4515_lo_n;
  wire n4518_lo_p;
  wire n4518_lo_n;
  wire n4521_lo_p;
  wire n4521_lo_n;
  wire n4524_lo_p;
  wire n4524_lo_n;
  wire n4527_lo_p;
  wire n4527_lo_n;
  wire n4530_lo_p;
  wire n4530_lo_n;
  wire n4533_lo_p;
  wire n4533_lo_n;
  wire n4536_lo_p;
  wire n4536_lo_n;
  wire n4539_lo_p;
  wire n4539_lo_n;
  wire n4542_lo_p;
  wire n4542_lo_n;
  wire n4545_lo_p;
  wire n4545_lo_n;
  wire n4554_lo_p;
  wire n4554_lo_n;
  wire n4557_lo_p;
  wire n4557_lo_n;
  wire n4560_lo_p;
  wire n4560_lo_n;
  wire n4563_lo_p;
  wire n4563_lo_n;
  wire n4566_lo_p;
  wire n4566_lo_n;
  wire n4569_lo_p;
  wire n4569_lo_n;
  wire n4572_lo_p;
  wire n4572_lo_n;
  wire n4575_lo_p;
  wire n4575_lo_n;
  wire n4578_lo_p;
  wire n4578_lo_n;
  wire n4581_lo_p;
  wire n4581_lo_n;
  wire n4584_lo_p;
  wire n4584_lo_n;
  wire n4587_lo_p;
  wire n4587_lo_n;
  wire n4590_lo_p;
  wire n4590_lo_n;
  wire n4593_lo_p;
  wire n4593_lo_n;
  wire n4596_lo_p;
  wire n4596_lo_n;
  wire n4602_lo_p;
  wire n4602_lo_n;
  wire n4605_lo_p;
  wire n4605_lo_n;
  wire n4608_lo_p;
  wire n4608_lo_n;
  wire n4614_lo_p;
  wire n4614_lo_n;
  wire n4617_lo_p;
  wire n4617_lo_n;
  wire n4620_lo_p;
  wire n4620_lo_n;
  wire n4626_lo_p;
  wire n4626_lo_n;
  wire n4629_lo_p;
  wire n4629_lo_n;
  wire n4632_lo_p;
  wire n4632_lo_n;
  wire n4638_lo_p;
  wire n4638_lo_n;
  wire n4641_lo_p;
  wire n4641_lo_n;
  wire n4644_lo_p;
  wire n4644_lo_n;
  wire n4647_lo_p;
  wire n4647_lo_n;
  wire n4650_lo_p;
  wire n4650_lo_n;
  wire n4653_lo_p;
  wire n4653_lo_n;
  wire n4656_lo_p;
  wire n4656_lo_n;
  wire n4659_lo_p;
  wire n4659_lo_n;
  wire n4662_lo_p;
  wire n4662_lo_n;
  wire n4665_lo_p;
  wire n4665_lo_n;
  wire n4668_lo_p;
  wire n4668_lo_n;
  wire n4671_lo_p;
  wire n4671_lo_n;
  wire n4674_lo_p;
  wire n4674_lo_n;
  wire n4677_lo_p;
  wire n4677_lo_n;
  wire n4680_lo_p;
  wire n4680_lo_n;
  wire n4683_lo_p;
  wire n4683_lo_n;
  wire n4686_lo_p;
  wire n4686_lo_n;
  wire n4689_lo_p;
  wire n4689_lo_n;
  wire n4692_lo_p;
  wire n4692_lo_n;
  wire n4695_lo_p;
  wire n4695_lo_n;
  wire n4698_lo_p;
  wire n4698_lo_n;
  wire n4701_lo_p;
  wire n4701_lo_n;
  wire n4704_lo_p;
  wire n4704_lo_n;
  wire n4707_lo_p;
  wire n4707_lo_n;
  wire n4710_lo_p;
  wire n4710_lo_n;
  wire n4713_lo_p;
  wire n4713_lo_n;
  wire n4716_lo_p;
  wire n4716_lo_n;
  wire n4719_lo_p;
  wire n4719_lo_n;
  wire n4722_lo_p;
  wire n4722_lo_n;
  wire n4725_lo_p;
  wire n4725_lo_n;
  wire n4728_lo_p;
  wire n4728_lo_n;
  wire n4731_lo_p;
  wire n4731_lo_n;
  wire n4734_lo_p;
  wire n4734_lo_n;
  wire n4737_lo_p;
  wire n4737_lo_n;
  wire n4740_lo_p;
  wire n4740_lo_n;
  wire n4743_lo_p;
  wire n4743_lo_n;
  wire n4970_o2_p;
  wire n4970_o2_n;
  wire n4972_o2_p;
  wire n4972_o2_n;
  wire n4989_o2_p;
  wire n4989_o2_n;
  wire n5024_o2_p;
  wire n5024_o2_n;
  wire n5025_o2_p;
  wire n5025_o2_n;
  wire n5029_o2_p;
  wire n5029_o2_n;
  wire n5042_o2_p;
  wire n5042_o2_n;
  wire n5048_o2_p;
  wire n5048_o2_n;
  wire n5093_o2_p;
  wire n5093_o2_n;
  wire n5096_o2_p;
  wire n5096_o2_n;
  wire n5193_o2_p;
  wire n5193_o2_n;
  wire n5199_o2_p;
  wire n5199_o2_n;
  wire n5203_o2_p;
  wire n5203_o2_n;
  wire n5214_o2_p;
  wire n5214_o2_n;
  wire n5221_o2_p;
  wire n5221_o2_n;
  wire n5222_o2_p;
  wire n5222_o2_n;
  wire n5273_o2_p;
  wire n5273_o2_n;
  wire n5365_o2_p;
  wire n5365_o2_n;
  wire n5385_o2_p;
  wire n5385_o2_n;
  wire n5553_o2_p;
  wire n5553_o2_n;
  wire n5636_o2_p;
  wire n5636_o2_n;
  wire n5782_o2_p;
  wire n5782_o2_n;
  wire n5778_o2_p;
  wire n5778_o2_n;
  wire n5323_o2_p;
  wire n5323_o2_n;
  wire n5325_o2_p;
  wire n5325_o2_n;
  wire n5327_o2_p;
  wire n5327_o2_n;
  wire n5329_o2_p;
  wire n5329_o2_n;
  wire n5816_o2_p;
  wire n5816_o2_n;
  wire n5817_o2_p;
  wire n5817_o2_n;
  wire n5837_o2_p;
  wire n5837_o2_n;
  wire n5844_o2_p;
  wire n5844_o2_n;
  wire n5859_o2_p;
  wire n5859_o2_n;
  wire n5857_o2_p;
  wire n5857_o2_n;
  wire n5369_o2_p;
  wire n5369_o2_n;
  wire n5371_o2_p;
  wire n5371_o2_n;
  wire n5373_o2_p;
  wire n5373_o2_n;
  wire n5400_o2_p;
  wire n5400_o2_n;
  wire n5402_o2_p;
  wire n5402_o2_n;
  wire n5404_o2_p;
  wire n5404_o2_n;
  wire n5406_o2_p;
  wire n5406_o2_n;
  wire n5407_o2_p;
  wire n5407_o2_n;
  wire n5408_o2_p;
  wire n5408_o2_n;
  wire n2722_o2_p;
  wire n2722_o2_n;
  wire n1942_inv_p;
  wire n1942_inv_n;
  wire n5412_o2_p;
  wire n5412_o2_n;
  wire n1948_inv_p;
  wire n1948_inv_n;
  wire n5557_o2_p;
  wire n5557_o2_n;
  wire n5558_o2_p;
  wire n5558_o2_n;
  wire n5559_o2_p;
  wire n5559_o2_n;
  wire n5564_o2_p;
  wire n5564_o2_n;
  wire n5565_o2_p;
  wire n5565_o2_n;
  wire n1966_inv_p;
  wire n1966_inv_n;
  wire n5568_o2_p;
  wire n5568_o2_n;
  wire n5598_o2_p;
  wire n5598_o2_n;
  wire n5600_o2_p;
  wire n5600_o2_n;
  wire n5601_o2_p;
  wire n5601_o2_n;
  wire n5602_o2_p;
  wire n5602_o2_n;
  wire n5603_o2_p;
  wire n5603_o2_n;
  wire n2853_o2_p;
  wire n2853_o2_n;
  wire n5637_o2_p;
  wire n5637_o2_n;
  wire n1993_inv_p;
  wire n1993_inv_n;
  wire n1996_inv_p;
  wire n1996_inv_n;
  wire n5635_o2_p;
  wire n5635_o2_n;
  wire n5640_o2_p;
  wire n5640_o2_n;
  wire n5641_o2_p;
  wire n5641_o2_n;
  wire n5642_o2_p;
  wire n5642_o2_n;
  wire n5650_o2_p;
  wire n5650_o2_n;
  wire n5652_o2_p;
  wire n5652_o2_n;
  wire n5653_o2_p;
  wire n5653_o2_n;
  wire n5654_o2_p;
  wire n5654_o2_n;
  wire n5655_o2_p;
  wire n5655_o2_n;
  wire n5657_o2_p;
  wire n5657_o2_n;
  wire n2029_inv_p;
  wire n2029_inv_n;
  wire n5661_o2_p;
  wire n5661_o2_n;
  wire n5656_o2_p;
  wire n5656_o2_n;
  wire n5663_o2_p;
  wire n5663_o2_n;
  wire n2041_inv_p;
  wire n2041_inv_n;
  wire n5795_o2_p;
  wire n5795_o2_n;
  wire n5796_o2_p;
  wire n5796_o2_n;
  wire n5797_o2_p;
  wire n5797_o2_n;
  wire n5739_o2_p;
  wire n5739_o2_n;
  wire n5773_o2_p;
  wire n5773_o2_n;
  wire n2059_inv_p;
  wire n2059_inv_n;
  wire n5799_o2_p;
  wire n5799_o2_n;
  wire n5802_o2_p;
  wire n5802_o2_n;
  wire n2068_inv_p;
  wire n2068_inv_n;
  wire n5831_o2_p;
  wire n5831_o2_n;
  wire n5833_o2_p;
  wire n5833_o2_n;
  wire n5820_o2_p;
  wire n5820_o2_n;
  wire n5823_o2_p;
  wire n5823_o2_n;
  wire n5824_o2_p;
  wire n5824_o2_n;
  wire n5869_o2_p;
  wire n5869_o2_n;
  wire n5848_o2_p;
  wire n5848_o2_n;
  wire n5849_o2_p;
  wire n5849_o2_n;
  wire n5856_o2_p;
  wire n5856_o2_n;
  wire n5896_o2_p;
  wire n5896_o2_n;
  wire n2754_o2_p;
  wire n2754_o2_n;
  wire n2908_o2_p;
  wire n2908_o2_n;
  wire n5892_o2_p;
  wire n5892_o2_n;
  wire n5915_o2_p;
  wire n5915_o2_n;
  wire n5919_o2_p;
  wire n5919_o2_n;
  wire n5918_o2_p;
  wire n5918_o2_n;
  wire n5920_o2_p;
  wire n5920_o2_n;
  wire n5917_o2_p;
  wire n5917_o2_n;
  wire lo586_buf_o2_p;
  wire lo586_buf_o2_n;
  wire n2818_o2_p;
  wire n2818_o2_n;
  wire n2863_o2_p;
  wire n2863_o2_n;
  wire n2134_inv_p;
  wire n2134_inv_n;
  wire n2725_o2_p;
  wire n2725_o2_n;
  wire n3016_o2_p;
  wire n3016_o2_n;
  wire n3013_o2_p;
  wire n3013_o2_n;
  wire n2655_o2_p;
  wire n2655_o2_n;
  wire n2149_inv_p;
  wire n2149_inv_n;
  wire lo562_buf_o2_p;
  wire lo562_buf_o2_n;
  wire n2155_inv_p;
  wire n2155_inv_n;
  wire n2531_o2_p;
  wire n2531_o2_n;
  wire n2700_o2_p;
  wire n2700_o2_n;
  wire n5908_o2_p;
  wire n5908_o2_n;
  wire n5910_o2_p;
  wire n5910_o2_n;
  wire n5912_o2_p;
  wire n5912_o2_n;
  wire n5914_o2_p;
  wire n5914_o2_n;
  wire n2753_o2_p;
  wire n2753_o2_n;
  wire n2878_o2_p;
  wire n2878_o2_n;
  wire n2182_inv_p;
  wire n2182_inv_n;
  wire n5934_o2_p;
  wire n5934_o2_n;
  wire n5936_o2_p;
  wire n5936_o2_n;
  wire n5938_o2_p;
  wire n5938_o2_n;
  wire n2728_o2_p;
  wire n2728_o2_n;
  wire lo358_buf_o2_p;
  wire lo358_buf_o2_n;
  wire lo418_buf_o2_p;
  wire lo418_buf_o2_n;
  wire lo474_buf_o2_p;
  wire lo474_buf_o2_n;
  wire lo554_buf_o2_p;
  wire lo554_buf_o2_n;
  wire lo558_buf_o2_p;
  wire lo558_buf_o2_n;
  wire lo574_buf_o2_p;
  wire lo574_buf_o2_n;
  wire n2215_inv_p;
  wire n2215_inv_n;
  wire n2218_inv_p;
  wire n2218_inv_n;
  wire n2221_inv_p;
  wire n2221_inv_n;
  wire lo450_buf_o2_p;
  wire lo450_buf_o2_n;
  wire n2910_o2_p;
  wire n2910_o2_n;
  wire n2683_o2_p;
  wire n2683_o2_n;
  wire n2828_o2_p;
  wire n2828_o2_n;
  wire n2582_o2_p;
  wire n2582_o2_n;
  wire n2600_o2_p;
  wire n2600_o2_n;
  wire n2542_o2_p;
  wire n2542_o2_n;
  wire n2703_o2_p;
  wire n2703_o2_n;
  wire lo510_buf_o2_p;
  wire lo510_buf_o2_n;
  wire lo514_buf_o2_p;
  wire lo514_buf_o2_n;
  wire lo538_buf_o2_p;
  wire lo538_buf_o2_n;
  wire lo578_buf_o2_p;
  wire lo578_buf_o2_n;
  wire n2260_inv_p;
  wire n2260_inv_n;
  wire n2666_o2_p;
  wire n2666_o2_n;
  wire n2667_o2_p;
  wire n2667_o2_n;
  wire n2660_o2_p;
  wire n2660_o2_n;
  wire n2272_inv_p;
  wire n2272_inv_n;
  wire lo454_buf_o2_p;
  wire lo454_buf_o2_n;
  wire n3593_o2_p;
  wire n3593_o2_n;
  wire n3048_o2_p;
  wire n3048_o2_n;
  wire lo410_buf_o2_p;
  wire lo410_buf_o2_n;
  wire lo502_buf_o2_p;
  wire lo502_buf_o2_n;
  wire lo506_buf_o2_p;
  wire lo506_buf_o2_n;
  wire lo550_buf_o2_p;
  wire lo550_buf_o2_n;
  wire lo570_buf_o2_p;
  wire lo570_buf_o2_n;
  wire lo582_buf_o2_p;
  wire lo582_buf_o2_n;
  wire n2302_inv_p;
  wire n2302_inv_n;
  wire n2305_inv_p;
  wire n2305_inv_n;
  wire n3499_o2_p;
  wire n3499_o2_n;
  wire n2311_inv_p;
  wire n2311_inv_n;
  wire n2870_o2_p;
  wire n2870_o2_n;
  wire n2317_inv_p;
  wire n2317_inv_n;
  wire n2689_o2_p;
  wire n2689_o2_n;
  wire n2323_inv_p;
  wire n2323_inv_n;
  wire n2662_o2_p;
  wire n2662_o2_n;
  wire lo350_buf_o2_p;
  wire lo350_buf_o2_n;
  wire lo498_buf_o2_p;
  wire lo498_buf_o2_n;
  wire lo518_buf_o2_p;
  wire lo518_buf_o2_n;
  wire lo522_buf_o2_p;
  wire lo522_buf_o2_n;
  wire lo598_buf_o2_p;
  wire lo598_buf_o2_n;
  wire n2344_inv_p;
  wire n2344_inv_n;
  wire n2347_inv_p;
  wire n2347_inv_n;
  wire n2350_inv_p;
  wire n2350_inv_n;
  wire n2353_inv_p;
  wire n2353_inv_n;
  wire n2356_inv_p;
  wire n2356_inv_n;
  wire n2359_inv_p;
  wire n2359_inv_n;
  wire n2872_o2_p;
  wire n2872_o2_n;
  wire n3313_o2_p;
  wire n3313_o2_n;
  wire n3273_o2_p;
  wire n3273_o2_n;
  wire n2848_o2_p;
  wire n2848_o2_n;
  wire n2893_o2_p;
  wire n2893_o2_n;
  wire n3267_o2_p;
  wire n3267_o2_n;
  wire n2925_o2_p;
  wire n2925_o2_n;
  wire n2839_o2_p;
  wire n2839_o2_n;
  wire n2831_o2_p;
  wire n2831_o2_n;
  wire n2558_o2_p;
  wire n2558_o2_n;
  wire n2562_o2_p;
  wire n2562_o2_n;
  wire n2825_o2_p;
  wire n2825_o2_n;
  wire n3263_o2_p;
  wire n3263_o2_n;
  wire n3517_o2_p;
  wire n3517_o2_n;
  wire n2873_o2_p;
  wire n2873_o2_n;
  wire n2926_o2_p;
  wire n2926_o2_n;
  wire n3261_o2_p;
  wire n3261_o2_n;
  wire n3268_o2_p;
  wire n3268_o2_n;
  wire n3274_o2_p;
  wire n3274_o2_n;
  wire n3314_o2_p;
  wire n3314_o2_n;
  wire n3571_o2_p;
  wire n3571_o2_n;
  wire n2950_o2_p;
  wire n2950_o2_n;
  wire n2951_o2_p;
  wire n2951_o2_n;
  wire n3022_o2_p;
  wire n3022_o2_n;
  wire n3023_o2_p;
  wire n3023_o2_n;
  wire n3057_o2_p;
  wire n3057_o2_n;
  wire n3058_o2_p;
  wire n3058_o2_n;
  wire n2931_o2_p;
  wire n2931_o2_n;
  wire n2911_o2_p;
  wire n2911_o2_n;
  wire n2959_o2_p;
  wire n2959_o2_n;
  wire n2960_o2_p;
  wire n2960_o2_n;
  wire n2922_o2_p;
  wire n2922_o2_n;
  wire n2888_o2_p;
  wire n2888_o2_n;
  wire n2889_o2_p;
  wire n2889_o2_n;
  wire n3051_o2_p;
  wire n3051_o2_n;
  wire n3052_o2_p;
  wire n3052_o2_n;
  wire n3063_o2_p;
  wire n3063_o2_n;
  wire n2845_o2_p;
  wire n2845_o2_n;
  wire n2476_inv_p;
  wire n2476_inv_n;
  wire n3281_o2_p;
  wire n3281_o2_n;
  wire n3294_o2_p;
  wire n3294_o2_n;
  wire n2885_o2_p;
  wire n2885_o2_n;
  wire n2786_o2_p;
  wire n2786_o2_n;
  wire n2783_o2_p;
  wire n2783_o2_n;
  wire n2801_o2_p;
  wire n2801_o2_n;
  wire n2572_o2_p;
  wire n2572_o2_n;
  wire n2628_o2_p;
  wire n2628_o2_n;
  wire n2609_o2_p;
  wire n2609_o2_n;
  wire n2618_o2_p;
  wire n2618_o2_n;
  wire n2637_o2_p;
  wire n2637_o2_n;
  wire n2525_o2_p;
  wire n2525_o2_n;
  wire n2551_o2_p;
  wire n2551_o2_n;
  wire n3759_o2_p;
  wire n3759_o2_n;
  wire n2994_o2_p;
  wire n2994_o2_n;
  wire n3040_o2_p;
  wire n3040_o2_n;
  wire n2943_o2_p;
  wire n2943_o2_n;
  wire n2991_o2_p;
  wire n2991_o2_n;
  wire n3034_o2_p;
  wire n3034_o2_n;
  wire n2881_o2_p;
  wire n2881_o2_n;
  wire n3021_o2_p;
  wire n3021_o2_n;
  wire n3062_o2_p;
  wire n3062_o2_n;
  wire n2763_o2_p;
  wire n2763_o2_n;
  wire n2764_o2_p;
  wire n2764_o2_n;
  wire n2775_o2_p;
  wire n2775_o2_n;
  wire n2776_o2_p;
  wire n2776_o2_n;
  wire n2968_o2_p;
  wire n2968_o2_n;
  wire n2969_o2_p;
  wire n2969_o2_n;
  wire n2798_o2_p;
  wire n2798_o2_n;
  wire n3661_o2_p;
  wire n3661_o2_n;
  wire n2694_o2_p;
  wire n2694_o2_n;
  wire n2572_inv_p;
  wire n2572_inv_n;
  wire n2817_o2_p;
  wire n2817_o2_n;
  wire n2514_o2_p;
  wire n2514_o2_n;
  wire n2501_o2_p;
  wire n2501_o2_n;
  wire n2584_inv_p;
  wire n2584_inv_n;
  wire n2505_o2_p;
  wire n2505_o2_n;
  wire n2492_o2_p;
  wire n2492_o2_n;
  wire lo546_buf_o2_p;
  wire lo546_buf_o2_n;
  wire lo590_buf_o2_p;
  wire lo590_buf_o2_n;
  wire lo594_buf_o2_p;
  wire lo594_buf_o2_n;
  wire n2602_inv_p;
  wire n2602_inv_n;
  wire n2605_inv_p;
  wire n2605_inv_n;
  wire n2709_o2_p;
  wire n2709_o2_n;
  wire n2611_inv_p;
  wire n2611_inv_n;
  wire n2614_inv_p;
  wire n2614_inv_n;
  wire n2617_inv_p;
  wire n2617_inv_n;
  wire n2620_inv_p;
  wire n2620_inv_n;
  wire n3590_o2_p;
  wire n3590_o2_n;
  wire n3591_o2_p;
  wire n3591_o2_n;
  wire n2629_inv_p;
  wire n2629_inv_n;
  wire n3638_o2_p;
  wire n3638_o2_n;
  wire n3639_o2_p;
  wire n3639_o2_n;
  wire n2638_inv_p;
  wire n2638_inv_n;
  wire n2641_inv_p;
  wire n2641_inv_n;
  wire lo458_buf_o2_p;
  wire lo458_buf_o2_n;
  wire lo482_buf_o2_p;
  wire lo482_buf_o2_n;
  wire lo566_buf_o2_p;
  wire lo566_buf_o2_n;
  wire n2718_o2_p;
  wire n2718_o2_n;
  wire n3707_o2_p;
  wire n3707_o2_n;
  wire n3671_o2_p;
  wire n3671_o2_n;
  wire n3680_o2_p;
  wire n3680_o2_n;
  wire n3749_o2_p;
  wire n3749_o2_n;
  wire n3716_o2_p;
  wire n3716_o2_n;
  wire n3692_o2_p;
  wire n3692_o2_n;
  wire n2591_o2_p;
  wire n2591_o2_n;
  wire n3478_o2_p;
  wire n3478_o2_n;
  wire n3610_o2_p;
  wire n3610_o2_n;
  wire n3611_o2_p;
  wire n3611_o2_n;
  wire n2686_inv_p;
  wire n2686_inv_n;
  wire n2689_inv_p;
  wire n2689_inv_n;
  wire n2738_o2_p;
  wire n2738_o2_n;
  wire n3616_o2_p;
  wire n3616_o2_n;
  wire n3617_o2_p;
  wire n3617_o2_n;
  wire n3031_o2_p;
  wire n3031_o2_n;
  wire n2704_inv_p;
  wire n2704_inv_n;
  wire n3562_o2_p;
  wire n3562_o2_n;
  wire n2502_o2_p;
  wire n2502_o2_n;
  wire n3560_o2_p;
  wire n3560_o2_n;
  wire n3554_o2_p;
  wire n3554_o2_n;
  wire n3555_o2_p;
  wire n3555_o2_n;
  wire n3536_o2_p;
  wire n3536_o2_n;
  wire n3537_o2_p;
  wire n3537_o2_n;
  wire n3508_o2_p;
  wire n3508_o2_n;
  wire n3650_o2_p;
  wire n3650_o2_n;
  wire n3740_o2_p;
  wire n3740_o2_n;
  wire n3484_o2_p;
  wire n3484_o2_n;
  wire n2740_inv_p;
  wire n2740_inv_n;
  wire n2734_o2_p;
  wire n2734_o2_n;
  wire n2735_o2_p;
  wire n2735_o2_n;
  wire n2711_o2_p;
  wire n2711_o2_n;
  wire lo585_buf_o2_p;
  wire lo585_buf_o2_n;
  wire n2719_o2_p;
  wire n2719_o2_n;
  wire n2720_o2_p;
  wire n2720_o2_n;
  wire n2723_o2_p;
  wire n2723_o2_n;
  wire n2724_o2_p;
  wire n2724_o2_n;
  wire n3624_o2_p;
  wire n3624_o2_n;
  wire n3625_o2_p;
  wire n3625_o2_n;
  wire n3015_o2_p;
  wire n3015_o2_n;
  wire n3491_o2_p;
  wire n3491_o2_n;
  wire n2779_inv_p;
  wire n2779_inv_n;
  wire n2811_o2_p;
  wire n2811_o2_n;
  wire n3010_o2_p;
  wire n3010_o2_n;
  wire n3012_o2_p;
  wire n3012_o2_n;
  wire lo382_buf_o2_p;
  wire lo382_buf_o2_n;
  wire lo386_buf_o2_p;
  wire lo386_buf_o2_n;
  wire lo390_buf_o2_p;
  wire lo390_buf_o2_n;
  wire lo398_buf_o2_p;
  wire lo398_buf_o2_n;
  wire lo402_buf_o2_p;
  wire lo402_buf_o2_n;
  wire lo406_buf_o2_p;
  wire lo406_buf_o2_n;
  wire n3492_o2_p;
  wire n3492_o2_n;
  wire lo366_buf_o2_p;
  wire lo366_buf_o2_n;
  wire lo374_buf_o2_p;
  wire lo374_buf_o2_n;
  wire lo426_buf_o2_p;
  wire lo426_buf_o2_n;
  wire lo494_buf_o2_p;
  wire lo494_buf_o2_n;
  wire n2653_o2_p;
  wire n2653_o2_n;
  wire n2654_o2_p;
  wire n2654_o2_n;
  wire n2715_o2_p;
  wire n2715_o2_n;
  wire n2740_o2_p;
  wire n2740_o2_n;
  wire n2682_o2_p;
  wire n2682_o2_n;
  wire n2736_o2_p;
  wire n2736_o2_n;
  wire lo508_buf_o2_p;
  wire lo508_buf_o2_n;
  wire lo512_buf_o2_p;
  wire lo512_buf_o2_n;
  wire lo536_buf_o2_p;
  wire lo536_buf_o2_n;
  wire lo576_buf_o2_p;
  wire lo576_buf_o2_n;
  wire lo357_buf_o2_p;
  wire lo357_buf_o2_n;
  wire lo361_buf_o2_p;
  wire lo361_buf_o2_n;
  wire lo417_buf_o2_p;
  wire lo417_buf_o2_n;
  wire lo421_buf_o2_p;
  wire lo421_buf_o2_n;
  wire lo473_buf_o2_p;
  wire lo473_buf_o2_n;
  wire lo477_buf_o2_p;
  wire lo477_buf_o2_n;
  wire lo553_buf_o2_p;
  wire lo553_buf_o2_n;
  wire lo557_buf_o2_p;
  wire lo557_buf_o2_n;
  wire lo573_buf_o2_p;
  wire lo573_buf_o2_n;
  wire lo434_buf_o2_p;
  wire lo434_buf_o2_n;
  wire lo438_buf_o2_p;
  wire lo438_buf_o2_n;
  wire lo466_buf_o2_p;
  wire lo466_buf_o2_n;
  wire lo470_buf_o2_p;
  wire lo470_buf_o2_n;
  wire lo490_buf_o2_p;
  wire lo490_buf_o2_n;
  wire n2657_o2_p;
  wire n2657_o2_n;
  wire n2658_o2_p;
  wire n2658_o2_n;
  wire n2663_o2_p;
  wire n2663_o2_n;
  wire n2664_o2_p;
  wire n2664_o2_n;
  wire n2684_o2_p;
  wire n2684_o2_n;
  wire n2685_o2_p;
  wire n2685_o2_n;
  wire g1049_p;
  wire g1049_n;
  wire g1050_p;
  wire g1050_n;
  wire g1051_p;
  wire g1051_n;
  wire g1052_p;
  wire g1052_n;
  wire g1053_p;
  wire g1053_n;
  wire g1054_p;
  wire g1054_n;
  wire g1055_p;
  wire g1055_n;
  wire g1056_p;
  wire g1056_n;
  wire g1057_p;
  wire g1057_n;
  wire g1058_p;
  wire g1058_n;
  wire g1059_p;
  wire g1059_n;
  wire g1060_p;
  wire g1060_n;
  wire g1061_p;
  wire g1061_n;
  wire g1062_p;
  wire g1062_n;
  wire g1063_p;
  wire g1063_n;
  wire g1064_p;
  wire g1064_n;
  wire g1065_p;
  wire g1065_n;
  wire g1066_p;
  wire g1066_n;
  wire g1067_p;
  wire g1067_n;
  wire g1068_p;
  wire g1068_n;
  wire g1069_p;
  wire g1069_n;
  wire g1070_p;
  wire g1070_n;
  wire g1071_p;
  wire g1071_n;
  wire g1072_p;
  wire g1072_n;
  wire g1073_p;
  wire g1073_n;
  wire g1074_p;
  wire g1074_n;
  wire g1075_p;
  wire g1075_n;
  wire g1076_p;
  wire g1076_n;
  wire g1077_p;
  wire g1077_n;
  wire g1078_p;
  wire g1078_n;
  wire g1079_p;
  wire g1079_n;
  wire g1080_p;
  wire g1080_n;
  wire g1081_p;
  wire g1081_n;
  wire g1082_p;
  wire g1082_n;
  wire g1083_p;
  wire g1083_n;
  wire g1084_p;
  wire g1084_n;
  wire g1085_p;
  wire g1085_n;
  wire g1086_p;
  wire g1086_n;
  wire g1087_p;
  wire g1087_n;
  wire g1088_p;
  wire g1088_n;
  wire g1089_p;
  wire g1089_n;
  wire g1090_p;
  wire g1090_n;
  wire g1091_p;
  wire g1091_n;
  wire g1092_p;
  wire g1092_n;
  wire g1093_p;
  wire g1093_n;
  wire g1094_p;
  wire g1094_n;
  wire g1095_p;
  wire g1095_n;
  wire g1096_p;
  wire g1096_n;
  wire g1097_p;
  wire g1097_n;
  wire g1098_p;
  wire g1098_n;
  wire g1099_p;
  wire g1099_n;
  wire g1100_p;
  wire g1100_n;
  wire g1101_p;
  wire g1101_n;
  wire g1102_p;
  wire g1102_n;
  wire g1103_p;
  wire g1103_n;
  wire g1104_p;
  wire g1104_n;
  wire g1105_p;
  wire g1105_n;
  wire g1106_p;
  wire g1106_n;
  wire g1107_p;
  wire g1107_n;
  wire g1108_p;
  wire g1108_n;
  wire g1109_p;
  wire g1109_n;
  wire g1110_p;
  wire g1110_n;
  wire g1111_p;
  wire g1111_n;
  wire g1112_p;
  wire g1112_n;
  wire g1113_p;
  wire g1113_n;
  wire g1114_p;
  wire g1114_n;
  wire g1115_p;
  wire g1115_n;
  wire g1116_p;
  wire g1116_n;
  wire g1117_p;
  wire g1117_n;
  wire g1118_p;
  wire g1118_n;
  wire g1119_p;
  wire g1119_n;
  wire g1120_p;
  wire g1120_n;
  wire g1121_p;
  wire g1121_n;
  wire g1122_p;
  wire g1122_n;
  wire g1123_p;
  wire g1123_n;
  wire g1124_p;
  wire g1124_n;
  wire g1125_p;
  wire g1125_n;
  wire g1126_p;
  wire g1126_n;
  wire g1127_p;
  wire g1127_n;
  wire g1128_p;
  wire g1128_n;
  wire g1129_p;
  wire g1129_n;
  wire g1130_p;
  wire g1130_n;
  wire g1131_p;
  wire g1131_n;
  wire g1132_p;
  wire g1132_n;
  wire g1133_p;
  wire g1133_n;
  wire g1134_p;
  wire g1134_n;
  wire g1135_p;
  wire g1135_n;
  wire g1136_p;
  wire g1136_n;
  wire g1137_p;
  wire g1137_n;
  wire g1138_p;
  wire g1138_n;
  wire g1139_p;
  wire g1139_n;
  wire g1140_p;
  wire g1140_n;
  wire g1141_p;
  wire g1141_n;
  wire g1142_p;
  wire g1142_n;
  wire g1143_p;
  wire g1143_n;
  wire g1144_p;
  wire g1144_n;
  wire g1145_p;
  wire g1145_n;
  wire g1146_p;
  wire g1146_n;
  wire g1147_p;
  wire g1147_n;
  wire g1148_p;
  wire g1148_n;
  wire g1149_p;
  wire g1149_n;
  wire g1150_p;
  wire g1150_n;
  wire g1151_p;
  wire g1151_n;
  wire g1152_p;
  wire g1152_n;
  wire g1153_p;
  wire g1153_n;
  wire g1154_p;
  wire g1154_n;
  wire g1155_p;
  wire g1155_n;
  wire g1156_p;
  wire g1156_n;
  wire g1157_p;
  wire g1157_n;
  wire g1158_p;
  wire g1158_n;
  wire g1159_p;
  wire g1159_n;
  wire g1160_p;
  wire g1160_n;
  wire g1161_p;
  wire g1161_n;
  wire g1162_p;
  wire g1162_n;
  wire g1163_p;
  wire g1163_n;
  wire g1164_p;
  wire g1164_n;
  wire g1165_p;
  wire g1165_n;
  wire g1166_p;
  wire g1166_n;
  wire g1167_p;
  wire g1167_n;
  wire g1168_p;
  wire g1168_n;
  wire g1169_p;
  wire g1169_n;
  wire g1170_p;
  wire g1170_n;
  wire g1171_p;
  wire g1171_n;
  wire g1172_p;
  wire g1172_n;
  wire g1173_p;
  wire g1173_n;
  wire g1174_p;
  wire g1174_n;
  wire g1175_p;
  wire g1175_n;
  wire g1176_p;
  wire g1176_n;
  wire g1177_p;
  wire g1177_n;
  wire g1178_p;
  wire g1178_n;
  wire g1179_p;
  wire g1179_n;
  wire g1180_p;
  wire g1180_n;
  wire g1181_p;
  wire g1181_n;
  wire g1182_p;
  wire g1182_n;
  wire g1183_p;
  wire g1183_n;
  wire g1184_p;
  wire g1184_n;
  wire g1185_p;
  wire g1185_n;
  wire g1186_p;
  wire g1186_n;
  wire g1187_p;
  wire g1187_n;
  wire g1188_p;
  wire g1188_n;
  wire g1189_p;
  wire g1189_n;
  wire g1190_p;
  wire g1190_n;
  wire g1191_p;
  wire g1191_n;
  wire g1192_p;
  wire g1192_n;
  wire g1193_p;
  wire g1193_n;
  wire g1194_p;
  wire g1194_n;
  wire g1195_p;
  wire g1195_n;
  wire g1196_p;
  wire g1196_n;
  wire g1197_p;
  wire g1197_n;
  wire g1198_p;
  wire g1198_n;
  wire g1199_p;
  wire g1199_n;
  wire g1200_p;
  wire g1200_n;
  wire g1201_p;
  wire g1201_n;
  wire g1202_p;
  wire g1202_n;
  wire g1203_p;
  wire g1203_n;
  wire g1204_p;
  wire g1204_n;
  wire g1205_p;
  wire g1205_n;
  wire g1206_p;
  wire g1206_n;
  wire g1207_p;
  wire g1207_n;
  wire g1208_p;
  wire g1208_n;
  wire g1209_p;
  wire g1209_n;
  wire g1210_p;
  wire g1210_n;
  wire g1211_p;
  wire g1211_n;
  wire g1212_p;
  wire g1212_n;
  wire g1213_p;
  wire g1213_n;
  wire g1214_p;
  wire g1214_n;
  wire g1215_p;
  wire g1215_n;
  wire g1216_p;
  wire g1216_n;
  wire g1217_p;
  wire g1217_n;
  wire g1218_p;
  wire g1218_n;
  wire g1219_p;
  wire g1219_n;
  wire g1220_p;
  wire g1220_n;
  wire g1221_p;
  wire g1221_n;
  wire g1222_p;
  wire g1222_n;
  wire g1223_p;
  wire g1223_n;
  wire g1224_p;
  wire g1224_n;
  wire g1225_p;
  wire g1225_n;
  wire g1226_p;
  wire g1226_n;
  wire g1227_p;
  wire g1227_n;
  wire g1228_p;
  wire g1228_n;
  wire g1229_p;
  wire g1229_n;
  wire g1230_p;
  wire g1230_n;
  wire g1231_p;
  wire g1231_n;
  wire g1232_p;
  wire g1232_n;
  wire g1233_p;
  wire g1233_n;
  wire g1234_p;
  wire g1234_n;
  wire g1235_p;
  wire g1235_n;
  wire g1236_p;
  wire g1236_n;
  wire g1237_p;
  wire g1237_n;
  wire g1238_p;
  wire g1238_n;
  wire g1239_p;
  wire g1239_n;
  wire g1240_p;
  wire g1240_n;
  wire g1241_p;
  wire g1241_n;
  wire g1242_p;
  wire g1242_n;
  wire g1243_p;
  wire g1243_n;
  wire g1244_p;
  wire g1244_n;
  wire g1245_p;
  wire g1245_n;
  wire g1246_p;
  wire g1246_n;
  wire g1247_p;
  wire g1247_n;
  wire g1248_p;
  wire g1248_n;
  wire g1249_p;
  wire g1249_n;
  wire g1250_p;
  wire g1250_n;
  wire g1251_p;
  wire g1251_n;
  wire g1252_p;
  wire g1252_n;
  wire g1253_p;
  wire g1253_n;
  wire g1254_p;
  wire g1254_n;
  wire g1255_p;
  wire g1255_n;
  wire g1256_p;
  wire g1256_n;
  wire g1257_p;
  wire g1257_n;
  wire g1258_p;
  wire g1258_n;
  wire g1259_p;
  wire g1259_n;
  wire g1260_p;
  wire g1260_n;
  wire g1261_p;
  wire g1261_n;
  wire g1262_p;
  wire g1262_n;
  wire g1263_p;
  wire g1263_n;
  wire g1264_p;
  wire g1264_n;
  wire g1265_p;
  wire g1265_n;
  wire g1266_p;
  wire g1266_n;
  wire g1267_p;
  wire g1267_n;
  wire g1268_p;
  wire g1268_n;
  wire g1269_p;
  wire g1269_n;
  wire g1270_p;
  wire g1270_n;
  wire g1271_p;
  wire g1271_n;
  wire g1272_p;
  wire g1272_n;
  wire g1273_p;
  wire g1273_n;
  wire g1274_p;
  wire g1274_n;
  wire g1275_p;
  wire g1275_n;
  wire g1276_p;
  wire g1276_n;
  wire g1277_p;
  wire g1277_n;
  wire g1278_p;
  wire g1278_n;
  wire g1279_p;
  wire g1279_n;
  wire g1280_p;
  wire g1280_n;
  wire g1281_p;
  wire g1281_n;
  wire g1282_p;
  wire g1282_n;
  wire g1283_p;
  wire g1283_n;
  wire g1284_p;
  wire g1284_n;
  wire g1285_p;
  wire g1285_n;
  wire g1286_p;
  wire g1286_n;
  wire g1287_p;
  wire g1287_n;
  wire g1288_p;
  wire g1288_n;
  wire g1289_p;
  wire g1289_n;
  wire g1290_p;
  wire g1290_n;
  wire g1291_p;
  wire g1291_n;
  wire g1292_p;
  wire g1292_n;
  wire g1293_p;
  wire g1293_n;
  wire g1294_p;
  wire g1294_n;
  wire g1295_p;
  wire g1295_n;
  wire g1296_p;
  wire g1296_n;
  wire g1297_p;
  wire g1297_n;
  wire g1298_p;
  wire g1298_n;
  wire g1299_p;
  wire g1299_n;
  wire g1300_p;
  wire g1300_n;
  wire g1301_p;
  wire g1301_n;
  wire g1302_p;
  wire g1302_n;
  wire g1303_p;
  wire g1303_n;
  wire g1304_p;
  wire g1304_n;
  wire g1305_p;
  wire g1305_n;
  wire g1306_p;
  wire g1306_n;
  wire g1307_p;
  wire g1307_n;
  wire g1308_p;
  wire g1308_n;
  wire g1309_p;
  wire g1309_n;
  wire g1310_p;
  wire g1310_n;
  wire g1311_p;
  wire g1311_n;
  wire g1312_p;
  wire g1312_n;
  wire g1313_p;
  wire g1313_n;
  wire g1314_p;
  wire g1314_n;
  wire g1315_p;
  wire g1315_n;
  wire g1316_p;
  wire g1316_n;
  wire g1317_p;
  wire g1317_n;
  wire g1318_p;
  wire g1318_n;
  wire g1319_p;
  wire g1319_n;
  wire g1320_p;
  wire g1320_n;
  wire g1321_p;
  wire g1321_n;
  wire g1322_p;
  wire g1322_n;
  wire g1323_p;
  wire g1323_n;
  wire g1324_p;
  wire g1324_n;
  wire g1325_p;
  wire g1325_n;
  wire g1326_p;
  wire g1326_n;
  wire g1327_p;
  wire g1327_n;
  wire g1328_p;
  wire g1328_n;
  wire g1329_p;
  wire g1329_n;
  wire g1330_p;
  wire g1330_n;
  wire g1331_p;
  wire g1331_n;
  wire g1332_p;
  wire g1332_n;
  wire g1333_p;
  wire g1333_n;
  wire g1334_p;
  wire g1334_n;
  wire g1335_p;
  wire g1335_n;
  wire g1336_p;
  wire g1336_n;
  wire g1337_p;
  wire g1337_n;
  wire g1338_p;
  wire g1338_n;
  wire g1339_p;
  wire g1339_n;
  wire g1340_p;
  wire g1340_n;
  wire g1341_p;
  wire g1341_n;
  wire g1342_p;
  wire g1342_n;
  wire g1343_p;
  wire g1343_n;
  wire g1344_p;
  wire g1344_n;
  wire g1345_p;
  wire g1345_n;
  wire g1346_p;
  wire g1346_n;
  wire g1347_p;
  wire g1347_n;
  wire g1348_p;
  wire g1348_n;
  wire g1349_p;
  wire g1349_n;
  wire g1350_p;
  wire g1350_n;
  wire g1351_p;
  wire g1351_n;
  wire g1352_p;
  wire g1352_n;
  wire g1353_p;
  wire g1353_n;
  wire g1354_p;
  wire g1354_n;
  wire g1355_p;
  wire g1355_n;
  wire g1356_p;
  wire g1356_n;
  wire g1357_p;
  wire g1357_n;
  wire g1358_p;
  wire g1358_n;
  wire g1359_p;
  wire g1359_n;
  wire g1360_p;
  wire g1360_n;
  wire g1361_p;
  wire g1361_n;
  wire g1362_p;
  wire g1362_n;
  wire g1363_p;
  wire g1363_n;
  wire g1364_p;
  wire g1364_n;
  wire g1365_p;
  wire g1365_n;
  wire g1366_p;
  wire g1366_n;
  wire g1367_p;
  wire g1367_n;
  wire g1368_p;
  wire g1368_n;
  wire g1369_p;
  wire g1369_n;
  wire g1370_p;
  wire g1370_n;
  wire g1371_p;
  wire g1371_n;
  wire g1372_p;
  wire g1372_n;
  wire g1373_p;
  wire g1373_n;
  wire g1374_p;
  wire g1374_n;
  wire g1375_p;
  wire g1375_n;
  wire g1376_p;
  wire g1376_n;
  wire g1377_p;
  wire g1377_n;
  wire g1378_p;
  wire g1378_n;
  wire g1379_p;
  wire g1379_n;
  wire g1380_p;
  wire g1380_n;
  wire g1381_p;
  wire g1381_n;
  wire g1382_p;
  wire g1382_n;
  wire g1383_p;
  wire g1383_n;
  wire g1384_p;
  wire g1384_n;
  wire g1385_p;
  wire g1385_n;
  wire g1386_p;
  wire g1386_n;
  wire g1387_p;
  wire g1387_n;
  wire g1388_p;
  wire g1388_n;
  wire g1389_p;
  wire g1389_n;
  wire g1390_p;
  wire g1390_n;
  wire g1391_p;
  wire g1391_n;
  wire g1392_p;
  wire g1392_n;
  wire g1393_p;
  wire g1393_n;
  wire g1394_p;
  wire g1394_n;
  wire g1395_p;
  wire g1395_n;
  wire g1396_p;
  wire g1396_n;
  wire g1397_p;
  wire g1397_n;
  wire g1398_p;
  wire g1398_n;
  wire g1399_p;
  wire g1399_n;
  wire g1400_p;
  wire g1400_n;
  wire g1401_p;
  wire g1401_n;
  wire g1402_p;
  wire g1402_n;
  wire g1403_p;
  wire g1403_n;
  wire g1404_p;
  wire g1404_n;
  wire g1405_p;
  wire g1405_n;
  wire g1406_p;
  wire g1406_n;
  wire g1407_p;
  wire g1407_n;
  wire g1408_p;
  wire g1408_n;
  wire g1409_p;
  wire g1409_n;
  wire g1410_p;
  wire g1410_n;
  wire g1411_p;
  wire g1411_n;
  wire g1412_p;
  wire g1412_n;
  wire g1413_p;
  wire g1413_n;
  wire g1414_p;
  wire g1414_n;
  wire g1415_p;
  wire g1415_n;
  wire g1416_p;
  wire g1416_n;
  wire g1417_p;
  wire g1417_n;
  wire g1418_p;
  wire g1418_n;
  wire g1419_p;
  wire g1419_n;
  wire g1420_p;
  wire g1420_n;
  wire g1421_p;
  wire g1421_n;
  wire g1422_p;
  wire g1422_n;
  wire g1423_p;
  wire g1423_n;
  wire g1424_p;
  wire g1424_n;
  wire g1425_p;
  wire g1425_n;
  wire g1426_p;
  wire g1426_n;
  wire g1427_p;
  wire g1427_n;
  wire g1428_p;
  wire g1428_n;
  wire g1429_p;
  wire g1429_n;
  wire g1430_p;
  wire g1430_n;
  wire g1431_p;
  wire g1431_n;
  wire g1432_p;
  wire g1432_n;
  wire g1433_p;
  wire g1433_n;
  wire g1434_p;
  wire g1434_n;
  wire g1435_p;
  wire g1435_n;
  wire g1436_p;
  wire g1436_n;
  wire g1437_p;
  wire g1437_n;
  wire g1438_p;
  wire g1438_n;
  wire g1439_p;
  wire g1439_n;
  wire g1440_p;
  wire g1440_n;
  wire g1441_p;
  wire g1441_n;
  wire g1442_p;
  wire g1442_n;
  wire g1443_p;
  wire g1443_n;
  wire g1444_p;
  wire g1444_n;
  wire g1445_p;
  wire g1445_n;
  wire g1446_p;
  wire g1446_n;
  wire g1447_p;
  wire g1447_n;
  wire g1448_p;
  wire g1448_n;
  wire g1449_p;
  wire g1449_n;
  wire g1450_p;
  wire g1450_n;
  wire g1451_p;
  wire g1451_n;
  wire g1452_p;
  wire g1452_n;
  wire g1453_p;
  wire g1453_n;
  wire g1454_p;
  wire g1454_n;
  wire g1455_p;
  wire g1455_n;
  wire g1456_p;
  wire g1456_n;
  wire g1457_p;
  wire g1457_n;
  wire g1458_p;
  wire g1458_n;
  wire g1459_p;
  wire g1459_n;
  wire g1460_p;
  wire g1460_n;
  wire g1461_p;
  wire g1461_n;
  wire g1462_p;
  wire g1462_n;
  wire g1463_p;
  wire g1463_n;
  wire g1464_p;
  wire g1464_n;
  wire g1465_p;
  wire g1465_n;
  wire g1466_p;
  wire g1466_n;
  wire g1467_p;
  wire g1467_n;
  wire g1468_p;
  wire g1468_n;
  wire g1469_p;
  wire g1469_n;
  wire g1470_p;
  wire g1470_n;
  wire g1471_p;
  wire g1471_n;
  wire g1472_p;
  wire g1472_n;
  wire g1473_p;
  wire g1473_n;
  wire g1474_p;
  wire g1474_n;
  wire g1475_p;
  wire g1475_n;
  wire g1476_p;
  wire g1476_n;
  wire g1477_p;
  wire g1477_n;
  wire g1478_p;
  wire g1478_n;
  wire g1479_p;
  wire g1479_n;
  wire g1480_p;
  wire g1480_n;
  wire g1481_p;
  wire g1481_n;
  wire g1482_p;
  wire g1482_n;
  wire g1483_p;
  wire g1483_n;
  wire g1484_p;
  wire g1484_n;
  wire g1485_p;
  wire g1485_n;
  wire g1486_p;
  wire g1486_n;
  wire g1487_p;
  wire g1487_n;
  wire g1488_p;
  wire g1488_n;
  wire g1489_p;
  wire g1489_n;
  wire g1490_p;
  wire g1490_n;
  wire g1491_p;
  wire g1491_n;
  wire g1492_p;
  wire g1492_n;
  wire g1493_p;
  wire g1493_n;
  wire g1494_p;
  wire g1494_n;
  wire g1495_p;
  wire g1495_n;
  wire g1496_p;
  wire g1496_n;
  wire g1497_p;
  wire g1497_n;
  wire g1498_p;
  wire g1498_n;
  wire g1499_p;
  wire g1499_n;
  wire g1500_p;
  wire g1500_n;
  wire g1501_p;
  wire g1501_n;
  wire g1502_p;
  wire g1502_n;
  wire g1503_p;
  wire g1503_n;
  wire g1504_p;
  wire g1504_n;
  wire g1505_p;
  wire g1505_n;
  wire g1506_p;
  wire g1506_n;
  wire g1507_p;
  wire g1507_n;
  wire g1508_p;
  wire g1508_n;
  wire g1509_p;
  wire g1509_n;
  wire g1510_p;
  wire g1510_n;
  wire g1511_p;
  wire g1511_n;
  wire g1512_p;
  wire g1512_n;
  wire g1513_p;
  wire g1513_n;
  wire g1514_p;
  wire g1514_n;
  wire g1515_p;
  wire g1515_n;
  wire g1516_p;
  wire g1516_n;
  wire g1517_p;
  wire g1517_n;
  wire g1518_p;
  wire g1518_n;
  wire g1519_p;
  wire g1519_n;
  wire g1520_p;
  wire g1520_n;
  wire g1521_p;
  wire g1521_n;
  wire g1522_p;
  wire g1522_n;
  wire g1523_p;
  wire g1523_n;
  wire g1524_p;
  wire g1524_n;
  wire g1525_p;
  wire g1525_n;
  wire g1526_p;
  wire g1526_n;
  wire g1527_p;
  wire g1527_n;
  wire g1528_p;
  wire g1528_n;
  wire g1529_p;
  wire g1529_n;
  wire g1530_p;
  wire g1530_n;
  wire g1531_p;
  wire g1531_n;
  wire g1532_p;
  wire g1532_n;
  wire g1533_p;
  wire g1533_n;
  wire g1534_p;
  wire g1534_n;
  wire g1535_p;
  wire g1535_n;
  wire g1536_p;
  wire g1536_n;
  wire g1537_p;
  wire g1537_n;
  wire g1538_p;
  wire g1538_n;
  wire g1539_p;
  wire g1539_n;
  wire g1540_p;
  wire g1540_n;
  wire g1541_p;
  wire g1541_n;
  wire g1542_p;
  wire g1542_n;
  wire g1543_p;
  wire g1543_n;
  wire g1544_p;
  wire g1544_n;
  wire g1545_p;
  wire g1545_n;
  wire g1546_p;
  wire g1546_n;
  wire g1547_p;
  wire g1547_n;
  wire g1548_p;
  wire g1548_n;
  wire g1549_p;
  wire g1549_n;
  wire g1550_p;
  wire g1550_n;
  wire g1551_p;
  wire g1551_n;
  wire g1552_p;
  wire g1552_n;
  wire g1553_p;
  wire g1553_n;
  wire g1554_p;
  wire g1554_n;
  wire g1555_p;
  wire g1555_n;
  wire g1556_p;
  wire g1556_n;
  wire g1557_p;
  wire g1557_n;
  wire g1558_p;
  wire g1558_n;
  wire g1559_p;
  wire g1559_n;
  wire g1560_p;
  wire g1560_n;
  wire g1561_p;
  wire g1561_n;
  wire g1562_p;
  wire g1562_n;
  wire g1563_p;
  wire g1563_n;
  wire g1564_p;
  wire g1564_n;
  wire g1565_p;
  wire g1565_n;
  wire g1566_p;
  wire g1566_n;
  wire g1567_p;
  wire g1567_n;
  wire g1568_p;
  wire g1568_n;
  wire g1569_p;
  wire g1569_n;
  wire g1570_p;
  wire g1570_n;
  wire g1571_p;
  wire g1571_n;
  wire g1572_p;
  wire g1572_n;
  wire g1573_p;
  wire g1573_n;
  wire g1574_p;
  wire g1574_n;
  wire g1575_p;
  wire g1575_n;
  wire g1576_p;
  wire g1576_n;
  wire g1577_p;
  wire g1577_n;
  wire g1578_p;
  wire g1578_n;
  wire g1579_p;
  wire g1579_n;
  wire g1580_p;
  wire g1580_n;
  wire g1581_p;
  wire g1581_n;
  wire g1582_p;
  wire g1582_n;
  wire g1583_p;
  wire g1583_n;
  wire g1584_p;
  wire g1584_n;
  wire g1585_p;
  wire g1585_n;
  wire g1586_p;
  wire g1586_n;
  wire g1587_p;
  wire g1587_n;
  wire g1588_p;
  wire g1588_n;
  wire g1589_p;
  wire g1589_n;
  wire g1590_p;
  wire g1590_n;
  wire g1591_p;
  wire g1591_n;
  wire g1592_p;
  wire g1592_n;
  wire g1593_p;
  wire g1593_n;
  wire g1594_p;
  wire g1594_n;
  wire g1595_p;
  wire g1595_n;
  wire g1596_p;
  wire g1596_n;
  wire g1597_p;
  wire g1597_n;
  wire g1598_p;
  wire g1598_n;
  wire g1599_p;
  wire g1599_n;
  wire g1600_p;
  wire g1600_n;
  wire g1601_p;
  wire g1601_n;
  wire g1602_p;
  wire g1602_n;
  wire g1603_p;
  wire g1603_n;
  wire g1604_p;
  wire g1604_n;
  wire g1605_p;
  wire g1605_n;
  wire g1606_p;
  wire g1606_n;
  wire g1607_p;
  wire g1607_n;
  wire g1608_p;
  wire g1608_n;
  wire g1609_p;
  wire g1609_n;
  wire g1610_p;
  wire g1610_n;
  wire g1611_p;
  wire g1611_n;
  wire g1612_p;
  wire g1612_n;
  wire g1613_p;
  wire g1613_n;
  wire g1614_p;
  wire g1614_n;
  wire g1615_p;
  wire g1615_n;
  wire g1616_p;
  wire g1616_n;
  wire g1617_p;
  wire g1617_n;
  wire g1618_p;
  wire g1618_n;
  wire g1619_p;
  wire g1619_n;
  wire g1620_p;
  wire g1620_n;
  wire g1621_p;
  wire g1621_n;
  wire g1622_p;
  wire g1622_n;
  wire g1623_p;
  wire g1623_n;
  wire g1624_p;
  wire g1624_n;
  wire g1625_p;
  wire g1625_n;
  wire g1626_p;
  wire g1626_n;
  wire g1627_p;
  wire g1627_n;
  wire g1628_p;
  wire g1628_n;
  wire g1629_p;
  wire g1629_n;
  wire g1630_p;
  wire g1630_n;
  wire g1631_p;
  wire g1631_n;
  wire g1632_p;
  wire g1632_n;
  wire g1633_p;
  wire g1633_n;
  wire g1634_p;
  wire g1634_n;
  wire g1635_p;
  wire g1635_n;
  wire g1636_p;
  wire g1636_n;
  wire g1637_p;
  wire g1637_n;
  wire g1638_p;
  wire g1638_n;
  wire g1639_p;
  wire g1639_n;
  wire g1640_p;
  wire g1640_n;
  wire g1641_p;
  wire g1641_n;
  wire g1642_p;
  wire g1642_n;
  wire g1643_p;
  wire g1643_n;
  wire g1644_p;
  wire g1644_n;
  wire g1645_p;
  wire g1645_n;
  wire g1646_p;
  wire g1646_n;
  wire g1647_p;
  wire g1647_n;
  wire g1648_p;
  wire g1648_n;
  wire g1649_p;
  wire g1649_n;
  wire g1650_p;
  wire g1650_n;
  wire g1651_p;
  wire g1651_n;
  wire g1652_p;
  wire g1652_n;
  wire g1653_p;
  wire g1653_n;
  wire g1654_p;
  wire g1654_n;
  wire g1655_p;
  wire g1655_n;
  wire g1656_p;
  wire g1656_n;
  wire g1657_p;
  wire g1657_n;
  wire g1658_p;
  wire g1658_n;
  wire g1659_p;
  wire g1659_n;
  wire g1660_p;
  wire g1660_n;
  wire g1661_p;
  wire g1661_n;
  wire g1662_p;
  wire g1662_n;
  wire g1663_p;
  wire g1663_n;
  wire g1664_p;
  wire g1664_n;
  wire g1665_p;
  wire g1665_n;
  wire g1666_p;
  wire g1666_n;
  wire g1667_p;
  wire g1667_n;
  wire g1668_p;
  wire g1668_n;
  wire g1669_p;
  wire g1669_n;
  wire g1670_p;
  wire g1670_n;
  wire g1671_p;
  wire g1671_n;
  wire g1672_p;
  wire g1672_n;
  wire g1673_p;
  wire g1673_n;
  wire g1674_p;
  wire g1674_n;
  wire g1675_p;
  wire g1675_n;
  wire g1676_p;
  wire g1676_n;
  wire g1677_p;
  wire g1677_n;
  wire g1678_p;
  wire g1678_n;
  wire g1679_p;
  wire g1679_n;
  wire g1680_p;
  wire g1680_n;
  wire g1681_p;
  wire g1681_n;
  wire g1682_p;
  wire g1682_n;
  wire g1683_p;
  wire g1683_n;
  wire g1684_p;
  wire g1684_n;
  wire g1685_p;
  wire g1685_n;
  wire g1686_p;
  wire g1686_n;
  wire g1687_p;
  wire g1687_n;
  wire g1688_p;
  wire g1688_n;
  wire g1689_p;
  wire g1689_n;
  wire g1690_p;
  wire g1690_n;
  wire g1691_p;
  wire g1691_n;
  wire g1692_p;
  wire g1692_n;
  wire g1693_p;
  wire g1693_n;
  wire g1694_p;
  wire g1694_n;
  wire g1695_p;
  wire g1695_n;
  wire g1696_p;
  wire g1696_n;
  wire g1697_p;
  wire g1697_n;
  wire g1698_p;
  wire g1698_n;
  wire g1699_p;
  wire g1699_n;
  wire g1700_p;
  wire g1700_n;
  wire g1701_p;
  wire g1701_n;
  wire g1702_p;
  wire g1702_n;
  wire g1703_p;
  wire g1703_n;
  wire g1704_p;
  wire g1704_n;
  wire g1705_p;
  wire g1705_n;
  wire g1706_p;
  wire g1706_n;
  wire g1707_p;
  wire g1707_n;
  wire g1708_p;
  wire g1708_n;
  wire g1709_p;
  wire g1709_n;
  wire g1710_p;
  wire g1710_n;
  wire g1711_p;
  wire g1711_n;
  wire g1712_p;
  wire g1712_n;
  wire g1713_p;
  wire g1713_n;
  wire g1714_p;
  wire g1714_n;
  wire g1715_p;
  wire g1715_n;
  wire g1716_p;
  wire g1716_n;
  wire g1717_p;
  wire g1717_n;
  wire g1718_p;
  wire g1718_n;
  wire g1719_p;
  wire g1719_n;
  wire g1720_p;
  wire g1720_n;
  wire g1721_p;
  wire g1721_n;
  wire g1722_p;
  wire g1722_n;
  wire g1723_p;
  wire g1723_n;
  wire g1724_p;
  wire g1724_n;
  wire g1725_p;
  wire g1725_n;
  wire g1726_p;
  wire g1726_n;
  wire g1727_p;
  wire g1727_n;
  wire g1728_p;
  wire g1728_n;
  wire g1729_p;
  wire g1729_n;
  wire g1730_p;
  wire g1730_n;
  wire g1731_p;
  wire g1731_n;
  wire g1732_p;
  wire g1732_n;
  wire g1733_p;
  wire g1733_n;
  wire g1734_p;
  wire g1734_n;
  wire g1735_p;
  wire g1735_n;
  wire g1736_p;
  wire g1736_n;
  wire g1737_p;
  wire g1737_n;
  wire g1738_p;
  wire g1738_n;
  wire g1739_p;
  wire g1739_n;
  wire g1740_p;
  wire g1740_n;
  wire g1741_p;
  wire g1741_n;
  wire g1742_p;
  wire g1742_n;
  wire g1743_p;
  wire g1743_n;
  wire g1744_p;
  wire g1744_n;
  wire g1745_p;
  wire g1745_n;
  wire g1746_p;
  wire g1746_n;
  wire g1747_p;
  wire g1747_n;
  wire g1748_p;
  wire g1748_n;
  wire g1749_p;
  wire g1749_n;
  wire g1750_p;
  wire g1750_n;
  wire g1751_p;
  wire g1751_n;
  wire g1752_p;
  wire g1752_n;
  wire g1753_p;
  wire g1753_n;
  wire g1754_p;
  wire g1754_n;
  wire g1755_p;
  wire g1755_n;
  wire g1756_p;
  wire g1756_n;
  wire g1757_p;
  wire g1757_n;
  wire g1758_p;
  wire g1758_n;
  wire g1759_p;
  wire g1759_n;
  wire g1760_p;
  wire g1760_n;
  wire g1761_p;
  wire g1761_n;
  wire g1762_p;
  wire g1762_n;
  wire g1763_p;
  wire g1763_n;
  wire g1764_p;
  wire g1764_n;
  wire g1765_p;
  wire g1765_n;
  wire g1766_p;
  wire g1766_n;
  wire g1767_p;
  wire g1767_n;
  wire g1768_p;
  wire g1768_n;
  wire g1769_p;
  wire g1769_n;
  wire g1770_p;
  wire g1770_n;
  wire g1771_p;
  wire g1771_n;
  wire g1772_p;
  wire g1772_n;
  wire g1773_p;
  wire g1773_n;
  wire g1774_p;
  wire g1774_n;
  wire g1775_p;
  wire g1775_n;
  wire g1776_p;
  wire g1776_n;
  wire g1777_p;
  wire g1777_n;
  wire g1778_p;
  wire g1778_n;
  wire g1779_p;
  wire g1779_n;
  wire g1780_p;
  wire g1780_n;
  wire g1781_p;
  wire g1781_n;
  wire g1782_p;
  wire g1782_n;
  wire g1783_p;
  wire g1783_n;
  wire g1784_p;
  wire g1784_n;
  wire g1785_p;
  wire g1785_n;
  wire g1786_p;
  wire g1786_n;
  wire g1787_p;
  wire g1787_n;
  wire g1788_p;
  wire g1788_n;
  wire g1789_p;
  wire g1789_n;
  wire g1790_p;
  wire g1790_n;
  wire g1791_p;
  wire g1791_n;
  wire g1792_p;
  wire g1792_n;
  wire g1793_p;
  wire g1793_n;
  wire g1794_p;
  wire g1794_n;
  wire g1795_p;
  wire g1795_n;
  wire g1796_p;
  wire g1796_n;
  wire g1797_p;
  wire g1797_n;
  wire g1798_p;
  wire g1798_n;
  wire g1799_p;
  wire g1799_n;
  wire g1800_p;
  wire g1800_n;
  wire g1801_p;
  wire g1801_n;
  wire g1802_p;
  wire g1802_n;
  wire g1803_p;
  wire g1803_n;
  wire g1804_p;
  wire g1804_n;
  wire g1805_p;
  wire g1805_n;
  wire g1806_p;
  wire g1806_n;
  wire g1807_p;
  wire g1807_n;
  wire g1808_p;
  wire g1808_n;
  wire g1809_p;
  wire g1809_n;
  wire g1810_p;
  wire g1810_n;
  wire g1811_p;
  wire g1811_n;
  wire g1812_p;
  wire g1812_n;
  wire g1813_p;
  wire g1813_n;
  wire g1814_p;
  wire g1814_n;
  wire g1815_p;
  wire g1815_n;
  wire g1816_p;
  wire g1816_n;
  wire g1817_p;
  wire g1817_n;
  wire g1818_p;
  wire g1818_n;
  wire g1819_p;
  wire g1819_n;
  wire g1820_p;
  wire g1820_n;
  wire g1821_p;
  wire g1821_n;
  wire g1822_p;
  wire g1822_n;
  wire g1823_p;
  wire g1823_n;
  wire g1824_p;
  wire g1824_n;
  wire g1825_p;
  wire g1825_n;
  wire g1826_p;
  wire g1826_n;
  wire g1827_p;
  wire g1827_n;
  wire g1828_p;
  wire g1828_n;
  wire g1829_p;
  wire g1829_n;
  wire g1830_p;
  wire g1830_n;
  wire g1831_p;
  wire g1831_n;
  wire g1832_p;
  wire g1832_n;
  wire g1833_p;
  wire g1833_n;
  wire g1834_p;
  wire g1834_n;
  wire g1835_p;
  wire g1835_n;
  wire g1836_p;
  wire g1836_n;
  wire g1837_p;
  wire g1837_n;
  wire g1838_p;
  wire g1838_n;
  wire g1839_p;
  wire g1839_n;
  wire g1840_p;
  wire g1840_n;
  wire g1841_p;
  wire g1841_n;
  wire g1842_p;
  wire g1842_n;
  wire g1843_p;
  wire g1843_n;
  wire g1844_p;
  wire g1844_n;
  wire g1845_p;
  wire g1845_n;
  wire g1846_p;
  wire g1846_n;
  wire g1847_p;
  wire g1847_n;
  wire g1848_p;
  wire g1848_n;
  wire g1849_p;
  wire g1849_n;
  wire g1850_p;
  wire g1850_n;
  wire g1851_p;
  wire g1851_n;
  wire g1852_p;
  wire g1852_n;
  wire g1853_p;
  wire g1853_n;
  wire g1854_p;
  wire g1854_n;
  wire g1855_p;
  wire g1855_n;
  wire g1856_p;
  wire g1856_n;
  wire g1857_p;
  wire g1857_n;
  wire g1858_p;
  wire g1858_n;
  wire g1859_p;
  wire g1859_n;
  wire g1860_p;
  wire g1860_n;
  wire g1861_p;
  wire g1861_n;
  wire g1862_p;
  wire g1862_n;
  wire g1863_p;
  wire g1863_n;
  wire g1864_p;
  wire g1864_n;
  wire g1865_p;
  wire g1865_n;
  wire g1866_p;
  wire g1866_n;
  wire g1867_p;
  wire g1867_n;
  wire g1868_p;
  wire g1868_n;
  wire g1869_p;
  wire g1869_n;
  wire g1870_p;
  wire g1870_n;
  wire g1871_p;
  wire g1871_n;
  wire g1872_p;
  wire g1872_n;
  wire g1873_p;
  wire g1873_n;
  wire g1874_p;
  wire g1874_n;
  wire g1875_p;
  wire g1875_n;
  wire g1876_p;
  wire g1876_n;
  wire g1877_p;
  wire g1877_n;
  wire g1878_p;
  wire g1878_n;
  wire g1879_p;
  wire g1879_n;
  wire g1880_p;
  wire g1880_n;
  wire g1881_p;
  wire g1881_n;
  wire g1882_p;
  wire g1882_n;
  wire g1883_p;
  wire g1883_n;
  wire g1884_p;
  wire g1884_n;
  wire g1885_p;
  wire g1885_n;
  wire g1886_p;
  wire g1886_n;
  wire g1887_p;
  wire g1887_n;
  wire g1888_p;
  wire g1888_n;
  wire g1889_p;
  wire g1889_n;
  wire g1890_p;
  wire g1890_n;
  wire g1891_p;
  wire g1891_n;
  wire g1892_p;
  wire g1892_n;
  wire g1893_p;
  wire g1893_n;
  wire g1894_p;
  wire g1894_n;
  wire g1895_p;
  wire g1895_n;
  wire g1896_p;
  wire g1896_n;
  wire g1897_p;
  wire g1897_n;
  wire g1898_p;
  wire g1898_n;
  wire g1899_p;
  wire g1899_n;
  wire g1900_p;
  wire g1900_n;
  wire g1901_p;
  wire g1901_n;
  wire g1902_p;
  wire g1902_n;
  wire g1903_p;
  wire g1903_n;
  wire g1904_p;
  wire g1904_n;
  wire g1905_p;
  wire g1905_n;
  wire g1906_p;
  wire g1906_n;
  wire g1907_p;
  wire g1907_n;
  wire g1908_p;
  wire g1908_n;
  wire g1909_p;
  wire g1909_n;
  wire g1910_p;
  wire g1910_n;
  wire g1911_p;
  wire g1911_n;
  wire g1912_p;
  wire g1912_n;
  wire g1913_p;
  wire g1913_n;
  wire g1914_p;
  wire g1914_n;
  wire g1915_p;
  wire g1915_n;
  wire g1916_p;
  wire g1916_n;
  wire g1917_p;
  wire g1917_n;
  wire g1918_p;
  wire g1918_n;
  wire g1919_p;
  wire g1919_n;
  wire g1920_p;
  wire g1920_n;
  wire g1921_p;
  wire g1921_n;
  wire g1922_p;
  wire g1922_n;
  wire g1923_p;
  wire g1923_n;
  wire g1924_p;
  wire g1924_n;
  wire g1925_p;
  wire g1925_n;
  wire g1926_p;
  wire g1926_n;
  wire g1927_p;
  wire g1927_n;
  wire g1928_p;
  wire g1928_n;
  wire g1929_p;
  wire g1929_n;
  wire g1930_p;
  wire g1930_n;
  wire g1931_p;
  wire g1931_n;
  wire g1932_p;
  wire g1932_n;
  wire g1933_p;
  wire g1933_n;
  wire g1934_p;
  wire g1934_n;
  wire g1935_p;
  wire g1935_n;
  wire g1936_p;
  wire g1936_n;
  wire g1937_p;
  wire g1937_n;
  wire g1938_p;
  wire g1938_n;
  wire g1939_p;
  wire g1939_n;
  wire g1940_p;
  wire g1940_n;
  wire g1941_p;
  wire g1941_n;
  wire g1942_p;
  wire g1942_n;
  wire g1943_p;
  wire g1943_n;
  wire g1944_p;
  wire g1944_n;
  wire g1945_p;
  wire g1945_n;
  wire g1946_p;
  wire g1946_n;
  wire g1947_p;
  wire g1947_n;
  wire g1948_p;
  wire g1948_n;
  wire g1949_p;
  wire g1949_n;
  wire g1950_p;
  wire g1950_n;
  wire g1951_p;
  wire g1951_n;
  wire g1952_p;
  wire g1952_n;
  wire g1953_p;
  wire g1953_n;
  wire g1954_p;
  wire g1954_n;
  wire g1955_p;
  wire g1955_n;
  wire g1956_p;
  wire g1956_n;
  wire g1957_p;
  wire g1957_n;
  wire g1958_p;
  wire g1958_n;
  wire g1959_p;
  wire g1959_n;
  wire g1960_p;
  wire g1960_n;
  wire g1961_p;
  wire g1961_n;
  wire g1962_p;
  wire g1962_n;
  wire g1963_p;
  wire g1963_n;
  wire g1964_p;
  wire g1964_n;
  wire g1965_p;
  wire g1965_n;
  wire g1966_p;
  wire g1966_n;
  wire g1967_p;
  wire g1967_n;
  wire g1968_p;
  wire g1968_n;
  wire g1969_p;
  wire g1969_n;
  wire g1970_p;
  wire g1970_n;
  wire g1971_p;
  wire g1971_n;
  wire g1972_p;
  wire g1972_n;
  wire g1973_p;
  wire g1973_n;
  wire g1974_p;
  wire g1974_n;
  wire g1975_p;
  wire g1975_n;
  wire g1976_p;
  wire g1976_n;
  wire g1977_p;
  wire g1977_n;
  wire g1978_p;
  wire g1978_n;
  wire g1979_p;
  wire g1979_n;
  wire g1980_p;
  wire g1980_n;
  wire g1981_p;
  wire g1981_n;
  wire g1982_p;
  wire g1982_n;
  wire g1983_p;
  wire g1983_n;
  wire g1984_p;
  wire g1984_n;
  wire g1985_p;
  wire g1985_n;
  wire g1986_p;
  wire g1986_n;
  wire g1987_p;
  wire g1987_n;
  wire g1988_p;
  wire g1988_n;
  wire g1989_p;
  wire g1989_n;
  wire g1990_p;
  wire g1990_n;
  wire g1991_p;
  wire g1991_n;
  wire g1992_p;
  wire g1992_n;
  wire g1993_p;
  wire g1993_n;
  wire g1994_p;
  wire g1994_n;
  wire g1995_p;
  wire g1995_n;
  wire g1996_p;
  wire g1996_n;
  wire g1997_p;
  wire g1997_n;
  wire g1998_p;
  wire g1998_n;
  wire g1999_p;
  wire g1999_n;
  wire g2000_p;
  wire g2000_n;
  wire g2001_p;
  wire g2001_n;
  wire g2002_p;
  wire g2002_n;
  wire g2003_p;
  wire g2003_n;
  wire g2004_p;
  wire g2004_n;
  wire g2005_p;
  wire g2005_n;
  wire g2006_p;
  wire g2006_n;
  wire g2007_p;
  wire g2007_n;
  wire g2008_p;
  wire g2008_n;
  wire g2009_p;
  wire g2009_n;
  wire g2010_p;
  wire g2010_n;
  wire g2011_p;
  wire g2011_n;
  wire g2012_p;
  wire g2012_n;
  wire g2013_p;
  wire g2013_n;
  wire g2014_p;
  wire g2014_n;
  wire g2015_p;
  wire g2015_n;
  wire g2016_p;
  wire g2016_n;
  wire g2017_p;
  wire g2017_n;
  wire g2018_p;
  wire g2018_n;
  wire g2019_p;
  wire g2019_n;
  wire g2020_p;
  wire g2020_n;
  wire g2021_p;
  wire g2021_n;
  wire g2022_p;
  wire g2022_n;
  wire g2023_p;
  wire g2023_n;
  wire g2024_p;
  wire g2024_n;
  wire g2025_p;
  wire g2025_n;
  wire g2026_p;
  wire g2026_n;
  wire g2027_p;
  wire g2027_n;
  wire g2028_p;
  wire g2028_n;
  wire g2029_p;
  wire g2029_n;
  wire g2030_p;
  wire g2030_n;
  wire g2031_p;
  wire g2031_n;
  wire g2032_p;
  wire g2032_n;
  wire g2033_p;
  wire g2033_n;
  wire g2034_p;
  wire g2034_n;
  wire g2035_p;
  wire g2035_n;
  wire g2036_p;
  wire g2036_n;
  wire g2037_p;
  wire g2037_n;
  wire g2038_p;
  wire g2038_n;
  wire g2039_p;
  wire g2039_n;
  wire g2040_p;
  wire g2040_n;
  wire g2041_p;
  wire g2041_n;
  wire g2042_p;
  wire g2042_n;
  wire g2043_p;
  wire g2043_n;
  wire g2044_p;
  wire g2044_n;
  wire g2045_p;
  wire g2045_n;
  wire g2046_p;
  wire g2046_n;
  wire g2047_p;
  wire g2047_n;
  wire g2048_p;
  wire g2048_n;
  wire g2049_p;
  wire g2049_n;
  wire g2050_p;
  wire g2050_n;
  wire g2051_p;
  wire g2051_n;
  wire g2052_p;
  wire g2052_n;
  wire g2053_p;
  wire g2053_n;
  wire g2054_p;
  wire g2054_n;
  wire g2055_p;
  wire g2055_n;
  wire g2056_p;
  wire g2056_n;
  wire g2057_p;
  wire g2057_n;
  wire g2058_p;
  wire g2058_n;
  wire g2059_p;
  wire g2059_n;
  wire g2060_p;
  wire g2060_n;
  wire g2061_p;
  wire g2061_n;
  wire g2062_p;
  wire g2062_n;
  wire g2063_p;
  wire g2063_n;
  wire g2064_p;
  wire g2064_n;
  wire g2065_p;
  wire g2065_n;
  wire g2066_p;
  wire g2066_n;
  wire g2067_p;
  wire g2067_n;
  wire g2068_p;
  wire g2068_n;
  wire g2069_p;
  wire g2069_n;
  wire g2070_p;
  wire g2070_n;
  wire g2071_p;
  wire g2071_n;
  wire g2072_p;
  wire g2072_n;
  wire g2073_p;
  wire g2073_n;
  wire g2074_p;
  wire g2074_n;
  wire g2075_p;
  wire g2075_n;
  wire g2076_p;
  wire g2076_n;
  wire g2077_p;
  wire g2077_n;
  wire g2078_p;
  wire g2078_n;
  wire g2079_p;
  wire g2079_n;
  wire g2080_p;
  wire g2080_n;
  wire g2081_p;
  wire g2081_n;
  wire g2082_p;
  wire g2082_n;
  wire g2083_p;
  wire g2083_n;
  wire g2084_p;
  wire g2084_n;
  wire g2085_p;
  wire g2085_n;
  wire g2086_p;
  wire g2086_n;
  wire g2087_p;
  wire g2087_n;
  wire g2088_p;
  wire g2088_n;
  wire g2089_p;
  wire g2089_n;
  wire g2090_p;
  wire g2090_n;
  wire g2091_p;
  wire g2091_n;
  wire g2092_p;
  wire g2092_n;
  wire g2093_p;
  wire g2093_n;
  wire g2094_p;
  wire g2094_n;
  wire g2095_p;
  wire g2095_n;
  wire g2096_p;
  wire g2096_n;
  wire g2097_p;
  wire g2097_n;
  wire g2098_p;
  wire g2098_n;
  wire g2099_p;
  wire g2099_n;
  wire g2100_p;
  wire g2100_n;
  wire g2101_p;
  wire g2101_n;
  wire g2102_p;
  wire g2102_n;
  wire g2103_p;
  wire g2103_n;
  wire g2104_p;
  wire g2104_n;
  wire g2105_p;
  wire g2105_n;
  wire g2106_p;
  wire g2106_n;
  wire g2107_p;
  wire g2107_n;
  wire g2108_p;
  wire g2108_n;
  wire g2109_p;
  wire g2109_n;
  wire g2110_p;
  wire g2110_n;
  wire g2111_p;
  wire g2111_n;
  wire g2112_p;
  wire g2112_n;
  wire g2113_p;
  wire g2113_n;
  wire g2114_p;
  wire g2114_n;
  wire g2115_p;
  wire g2115_n;
  wire g2116_p;
  wire g2116_n;
  wire g2117_p;
  wire g2117_n;
  wire g2118_p;
  wire g2118_n;
  wire g2119_p;
  wire g2119_n;
  wire g2120_p;
  wire g2120_n;
  wire g2121_p;
  wire g2121_n;
  wire g2122_p;
  wire g2122_n;
  wire g2123_p;
  wire g2123_n;
  wire g2124_p;
  wire g2124_n;
  wire g2125_p;
  wire g2125_n;
  wire g2126_p;
  wire g2126_n;
  wire g2127_p;
  wire g2127_n;
  wire g2128_p;
  wire g2128_n;
  wire g2129_p;
  wire g2129_n;
  wire g2130_p;
  wire g2130_n;
  wire g2131_p;
  wire g2131_n;
  wire g2132_p;
  wire g2132_n;
  wire g2133_p;
  wire g2133_n;
  wire g2134_p;
  wire g2134_n;
  wire g2135_p;
  wire g2135_n;
  wire g2136_p;
  wire g2136_n;
  wire g2137_p;
  wire g2137_n;
  wire g2138_p;
  wire g2138_n;
  wire g2139_p;
  wire g2139_n;
  wire g2140_p;
  wire g2140_n;
  wire g2141_p;
  wire g2141_n;
  wire g2142_p;
  wire g2142_n;
  wire g2143_p;
  wire g2143_n;
  wire g2144_p;
  wire g2144_n;
  wire g2145_p;
  wire g2145_n;
  wire g2146_p;
  wire g2146_n;
  wire g2147_p;
  wire g2147_n;
  wire g2148_p;
  wire g2148_n;
  wire g2149_p;
  wire g2149_n;
  wire g2150_p;
  wire g2150_n;
  wire g2151_p;
  wire g2151_n;
  wire g2152_p;
  wire g2152_n;
  wire g2153_p;
  wire g2153_n;
  wire g2154_p;
  wire g2154_n;
  wire g2155_p;
  wire g2155_n;
  wire g2156_p;
  wire g2156_n;
  wire g2157_p;
  wire g2157_n;
  wire g2158_p;
  wire g2158_n;
  wire g2159_p;
  wire g2159_n;
  wire g2160_p;
  wire g2160_n;
  wire g2161_p;
  wire g2161_n;
  wire g2162_p;
  wire g2162_n;
  wire g2163_p;
  wire g2163_n;
  wire g2164_p;
  wire g2164_n;
  wire g2165_p;
  wire g2165_n;
  wire g2166_p;
  wire g2166_n;
  wire g2167_p;
  wire g2167_n;
  wire g2168_p;
  wire g2168_n;
  wire g2169_p;
  wire g2169_n;
  wire g2170_p;
  wire g2170_n;
  wire g2171_p;
  wire g2171_n;
  wire g2172_p;
  wire g2172_n;
  wire g2173_p;
  wire g2173_n;
  wire g2174_p;
  wire g2174_n;
  wire g2175_p;
  wire g2175_n;
  wire g2176_p;
  wire g2176_n;
  wire g2177_p;
  wire g2177_n;
  wire g2178_p;
  wire g2178_n;
  wire g2179_p;
  wire g2179_n;
  wire g2180_p;
  wire g2180_n;
  wire g2181_p;
  wire g2181_n;
  wire g2182_p;
  wire g2182_n;
  wire g2183_p;
  wire g2183_n;
  wire g2184_p;
  wire g2184_n;
  wire g2185_p;
  wire g2185_n;
  wire g2186_p;
  wire g2186_n;
  wire g2187_p;
  wire g2187_n;
  wire g2188_p;
  wire g2188_n;
  wire g2189_p;
  wire g2189_n;
  wire g2190_p;
  wire g2190_n;
  wire g2191_p;
  wire g2191_n;
  wire g2192_p;
  wire g2192_n;
  wire g2193_p;
  wire g2193_n;
  wire g2194_p;
  wire g2194_n;
  wire g2195_p;
  wire g2195_n;
  wire g2196_p;
  wire g2196_n;
  wire g2197_p;
  wire g2197_n;
  wire g2198_p;
  wire g2198_n;
  wire g2199_p;
  wire g2199_n;
  wire g2200_p;
  wire g2200_n;
  wire g2201_p;
  wire g2201_n;
  wire g2202_p;
  wire g2202_n;
  wire g2203_p;
  wire g2203_n;
  wire g2204_p;
  wire g2204_n;
  wire g2205_p;
  wire g2205_n;
  wire g2206_p;
  wire g2206_n;
  wire g2207_p;
  wire g2207_n;
  wire g2208_p;
  wire g2208_n;
  wire g2209_p;
  wire g2209_n;
  wire g2210_p;
  wire g2210_n;
  wire g2211_p;
  wire g2211_n;
  wire g2212_p;
  wire g2212_n;
  wire g2213_p;
  wire g2213_n;
  wire g2214_p;
  wire g2214_n;
  wire g2215_p;
  wire g2215_n;
  wire g2216_p;
  wire g2216_n;
  wire g2217_p;
  wire g2217_n;
  wire g2218_p;
  wire g2218_n;
  wire g2219_p;
  wire g2219_n;
  wire g2220_p;
  wire g2220_n;
  wire g2221_p;
  wire g2221_n;
  wire g2222_p;
  wire g2222_n;
  wire g2223_p;
  wire g2223_n;
  wire g2224_p;
  wire g2224_n;
  wire g2225_p;
  wire g2225_n;
  wire g2226_p;
  wire g2226_n;
  wire g2227_p;
  wire g2227_n;
  wire g2228_p;
  wire g2228_n;
  wire g2229_p;
  wire g2229_n;
  wire g2230_p;
  wire g2230_n;
  wire g2231_p;
  wire g2231_n;
  wire g2232_p;
  wire g2232_n;
  wire g2233_p;
  wire g2233_n;
  wire g2234_p;
  wire g2234_n;
  wire g2235_p;
  wire g2235_n;
  wire g2236_p;
  wire g2236_n;
  wire g2237_p;
  wire g2237_n;
  wire g2238_p;
  wire g2238_n;
  wire g2239_p;
  wire g2239_n;
  wire g2240_p;
  wire g2240_n;
  wire g2241_p;
  wire g2241_n;
  wire g2242_p;
  wire g2242_n;
  wire g2243_p;
  wire g2243_n;
  wire g2244_p;
  wire g2244_n;
  wire g2245_p;
  wire g2245_n;
  wire g2246_p;
  wire g2246_n;
  wire g2247_p;
  wire g2247_n;
  wire g2248_p;
  wire g2248_n;
  wire g2249_p;
  wire g2249_n;
  wire g2250_p;
  wire g2250_n;
  wire g2251_p;
  wire g2251_n;
  wire g2252_p;
  wire g2252_n;
  wire g2253_p;
  wire g2253_n;
  wire g2254_p;
  wire g2254_n;
  wire g2255_p;
  wire g2255_n;
  wire g2256_p;
  wire g2256_n;
  wire g2257_p;
  wire g2257_n;
  wire g2258_p;
  wire g2258_n;
  wire g2259_p;
  wire g2259_n;
  wire g2260_p;
  wire g2260_n;
  wire g2261_p;
  wire g2261_n;
  wire g2262_p;
  wire g2262_n;
  wire g2263_p;
  wire g2263_n;
  wire g2264_p;
  wire g2264_n;
  wire g2265_p;
  wire g2265_n;
  wire g2266_p;
  wire g2266_n;
  wire g2267_p;
  wire g2267_n;
  wire g2268_p;
  wire g2268_n;
  wire g2269_p;
  wire g2269_n;
  wire g2270_p;
  wire g2270_n;
  wire g2271_p;
  wire g2271_n;
  wire g2272_p;
  wire g2272_n;
  wire g2273_p;
  wire g2273_n;
  wire g2274_p;
  wire g2274_n;
  wire g2275_p;
  wire g2275_n;
  wire g2276_p;
  wire g2276_n;
  wire g2277_p;
  wire g2277_n;
  wire g2278_p;
  wire g2278_n;
  wire g2279_p;
  wire g2279_n;
  wire g2280_p;
  wire g2280_n;
  wire g2281_p;
  wire g2281_n;
  wire g2282_p;
  wire g2282_n;
  wire g2283_p;
  wire g2283_n;
  wire g2284_p;
  wire g2284_n;
  wire g2285_p;
  wire g2285_n;
  wire g2286_p;
  wire g2286_n;
  wire g2287_p;
  wire g2287_n;
  wire g2288_p;
  wire g2288_n;
  wire g2289_p;
  wire g2289_n;
  wire g2290_p;
  wire g2290_n;
  wire g2291_p;
  wire g2291_n;
  wire g2292_p;
  wire g2292_n;
  wire g2293_p;
  wire g2293_n;
  wire g2294_p;
  wire g2294_n;
  wire g2295_p;
  wire g2295_n;
  wire g2296_p;
  wire g2296_n;
  wire g2297_p;
  wire g2297_n;
  wire g2298_p;
  wire g2298_n;
  wire g2299_p;
  wire g2299_n;
  wire g2300_p;
  wire g2300_n;
  wire g2301_p;
  wire g2301_n;
  wire g2302_p;
  wire g2302_n;
  wire g2303_p;
  wire g2303_n;
  wire g2304_p;
  wire g2304_n;
  wire g2305_p;
  wire g2305_n;
  wire g2306_p;
  wire g2306_n;
  wire g2307_p;
  wire g2307_n;
  wire g2308_p;
  wire g2308_n;
  wire g2309_p;
  wire g2309_n;
  wire g2310_p;
  wire g2310_n;
  wire g2311_p;
  wire g2311_n;
  wire g2312_p;
  wire g2312_n;
  wire g2313_p;
  wire g2313_n;
  wire g2314_p;
  wire g2314_n;
  wire g2315_p;
  wire g2315_n;
  wire g2316_p;
  wire g2316_n;
  wire g2317_p;
  wire g2317_n;
  wire g2318_p;
  wire g2318_n;
  wire g2319_p;
  wire g2319_n;
  wire g2320_p;
  wire g2320_n;
  wire g2321_p;
  wire g2321_n;
  wire g2322_p;
  wire g2322_n;
  wire g2323_p;
  wire g2323_n;
  wire g2324_p;
  wire g2324_n;
  wire g2325_p;
  wire g2325_n;
  wire g2326_p;
  wire g2326_n;
  wire g2327_p;
  wire g2327_n;
  wire g2328_p;
  wire g2328_n;
  wire g2329_p;
  wire g2329_n;
  wire g2330_p;
  wire g2330_n;
  wire g2331_p;
  wire g2331_n;
  wire g2332_p;
  wire g2332_n;
  wire g2333_p;
  wire g2333_n;
  wire g2334_p;
  wire g2334_n;
  wire g2335_p;
  wire g2335_n;
  wire g2336_p;
  wire g2336_n;
  wire g2337_p;
  wire g2337_n;
  wire g2338_p;
  wire g2338_n;
  wire g2339_p;
  wire g2339_n;
  wire g2340_p;
  wire g2340_n;
  wire g2341_p;
  wire g2341_n;
  wire g2342_p;
  wire g2342_n;
  wire g2343_p;
  wire g2343_n;
  wire g2344_p;
  wire g2344_n;
  wire g2345_p;
  wire g2345_n;
  wire g2346_p;
  wire g2346_n;
  wire g2347_p;
  wire g2347_n;
  wire g2348_p;
  wire g2348_n;
  wire g2349_p;
  wire g2349_n;
  wire g2350_p;
  wire g2350_n;
  wire g2351_p;
  wire g2351_n;
  wire g2352_p;
  wire g2352_n;
  wire g2353_p;
  wire g2353_n;
  wire g2354_p;
  wire g2354_n;
  wire g2355_p;
  wire g2355_n;
  wire g2356_p;
  wire g2356_n;
  wire g2357_p;
  wire g2357_n;
  wire g2358_p;
  wire g2358_n;
  wire g2359_p;
  wire g2359_n;
  wire g2360_p;
  wire g2360_n;
  wire g2361_p;
  wire g2361_n;
  wire g2362_p;
  wire g2362_n;
  wire g2363_p;
  wire g2363_n;
  wire g2364_p;
  wire g2364_n;
  wire g2365_p;
  wire g2365_n;
  wire g2366_p;
  wire g2366_n;
  wire g2367_p;
  wire g2367_n;
  wire g2368_p;
  wire g2368_n;
  wire g2369_p;
  wire g2369_n;
  wire g2370_p;
  wire g2370_n;
  wire g2371_p;
  wire g2371_n;
  wire g2372_p;
  wire g2372_n;
  wire g2373_p;
  wire g2373_n;
  wire g2374_p;
  wire g2374_n;
  wire g2375_p;
  wire g2375_n;
  wire g2376_p;
  wire g2376_n;
  wire g2377_p;
  wire g2377_n;
  wire g2378_p;
  wire g2378_n;
  wire g2379_p;
  wire g2379_n;
  wire g2380_p;
  wire g2380_n;
  wire g2381_p;
  wire g2381_n;
  wire g2382_p;
  wire g2382_n;
  wire g2383_p;
  wire g2383_n;
  wire g2384_p;
  wire g2384_n;
  wire g2385_p;
  wire g2385_n;
  wire g2386_p;
  wire g2386_n;
  wire g2387_p;
  wire g2387_n;
  wire g2388_p;
  wire g2388_n;
  wire g2389_p;
  wire g2389_n;
  wire g2390_p;
  wire g2390_n;
  wire g2391_p;
  wire g2391_n;
  wire g2392_p;
  wire g2392_n;
  wire g2393_p;
  wire g2393_n;
  wire g2394_p;
  wire g2394_n;
  wire n4443_lo_n_spl_;
  wire n4479_lo_n_spl_;
  wire n3399_lo_p_spl_;
  wire n3399_lo_p_spl_0;
  wire n3399_lo_p_spl_00;
  wire n3399_lo_p_spl_01;
  wire n3399_lo_p_spl_1;
  wire n2619_lo_p_spl_;
  wire n4587_lo_n_spl_;
  wire n2739_lo_n_spl_;
  wire g1055_n_spl_;
  wire g1055_n_spl_0;
  wire g1055_n_spl_00;
  wire g1055_n_spl_000;
  wire g1055_n_spl_01;
  wire g1055_n_spl_1;
  wire g1055_n_spl_10;
  wire g1055_n_spl_11;
  wire n4563_lo_n_spl_;
  wire n4563_lo_n_spl_0;
  wire n4563_lo_n_spl_00;
  wire n4563_lo_n_spl_01;
  wire n4563_lo_n_spl_1;
  wire n4563_lo_p_spl_;
  wire n4563_lo_p_spl_0;
  wire n4563_lo_p_spl_00;
  wire n4563_lo_p_spl_01;
  wire n4563_lo_p_spl_1;
  wire n2551_o2_p_spl_;
  wire g1094_n_spl_;
  wire n5273_o2_n_spl_;
  wire g1101_n_spl_;
  wire n2786_o2_p_spl_;
  wire n2783_o2_p_spl_;
  wire n2786_o2_n_spl_;
  wire n2783_o2_n_spl_;
  wire n2801_o2_n_spl_;
  wire n2798_o2_n_spl_;
  wire n2801_o2_p_spl_;
  wire n2798_o2_p_spl_;
  wire n5837_o2_p_spl_;
  wire n5837_o2_p_spl_0;
  wire n2825_o2_p_spl_;
  wire n2825_o2_p_spl_0;
  wire n2825_o2_p_spl_00;
  wire n2825_o2_p_spl_000;
  wire n2825_o2_p_spl_001;
  wire n2825_o2_p_spl_01;
  wire n2825_o2_p_spl_010;
  wire n2825_o2_p_spl_011;
  wire n2825_o2_p_spl_1;
  wire n2825_o2_p_spl_10;
  wire n2825_o2_p_spl_100;
  wire n2825_o2_p_spl_101;
  wire n2825_o2_p_spl_11;
  wire n2825_o2_p_spl_110;
  wire n2825_o2_p_spl_111;
  wire n4731_lo_n_spl_;
  wire n4731_lo_n_spl_0;
  wire n4731_lo_n_spl_00;
  wire n4731_lo_n_spl_000;
  wire n4731_lo_n_spl_01;
  wire n4731_lo_n_spl_1;
  wire n4731_lo_n_spl_10;
  wire n4731_lo_n_spl_11;
  wire n4719_lo_p_spl_;
  wire n4719_lo_p_spl_0;
  wire n4719_lo_p_spl_00;
  wire n4719_lo_p_spl_000;
  wire n4719_lo_p_spl_001;
  wire n4719_lo_p_spl_01;
  wire n4719_lo_p_spl_010;
  wire n4719_lo_p_spl_011;
  wire n4719_lo_p_spl_1;
  wire n4719_lo_p_spl_10;
  wire n4719_lo_p_spl_100;
  wire n4719_lo_p_spl_101;
  wire n4719_lo_p_spl_11;
  wire n4719_lo_p_spl_110;
  wire n2825_o2_n_spl_;
  wire n4731_lo_p_spl_;
  wire n4731_lo_p_spl_0;
  wire n4731_lo_p_spl_00;
  wire n4731_lo_p_spl_000;
  wire n4731_lo_p_spl_01;
  wire n4731_lo_p_spl_1;
  wire n4731_lo_p_spl_10;
  wire n4731_lo_p_spl_11;
  wire n4719_lo_n_spl_;
  wire n4719_lo_n_spl_0;
  wire n4719_lo_n_spl_1;
  wire n2845_o2_p_spl_;
  wire n4683_lo_n_spl_;
  wire n4683_lo_n_spl_0;
  wire n4683_lo_n_spl_00;
  wire n4683_lo_n_spl_000;
  wire n4683_lo_n_spl_0000;
  wire n4683_lo_n_spl_0001;
  wire n4683_lo_n_spl_001;
  wire n4683_lo_n_spl_0010;
  wire n4683_lo_n_spl_0011;
  wire n4683_lo_n_spl_01;
  wire n4683_lo_n_spl_010;
  wire n4683_lo_n_spl_011;
  wire n4683_lo_n_spl_1;
  wire n4683_lo_n_spl_10;
  wire n4683_lo_n_spl_100;
  wire n4683_lo_n_spl_101;
  wire n4683_lo_n_spl_11;
  wire n4683_lo_n_spl_110;
  wire n4683_lo_n_spl_111;
  wire g1132_n_spl_;
  wire g1132_n_spl_0;
  wire g1132_n_spl_00;
  wire g1132_n_spl_1;
  wire n4683_lo_p_spl_;
  wire n4683_lo_p_spl_0;
  wire n4683_lo_p_spl_00;
  wire n4683_lo_p_spl_000;
  wire n4683_lo_p_spl_0000;
  wire n4683_lo_p_spl_0001;
  wire n4683_lo_p_spl_001;
  wire n4683_lo_p_spl_0010;
  wire n4683_lo_p_spl_0011;
  wire n4683_lo_p_spl_01;
  wire n4683_lo_p_spl_010;
  wire n4683_lo_p_spl_011;
  wire n4683_lo_p_spl_1;
  wire n4683_lo_p_spl_10;
  wire n4683_lo_p_spl_100;
  wire n4683_lo_p_spl_101;
  wire n4683_lo_p_spl_11;
  wire n4683_lo_p_spl_110;
  wire n4683_lo_p_spl_111;
  wire g1142_n_spl_;
  wire g1142_n_spl_0;
  wire g1142_n_spl_00;
  wire g1142_n_spl_1;
  wire n4671_lo_p_spl_;
  wire n4671_lo_p_spl_0;
  wire n4671_lo_p_spl_00;
  wire n4671_lo_p_spl_000;
  wire n4671_lo_p_spl_001;
  wire n4671_lo_p_spl_01;
  wire n4671_lo_p_spl_1;
  wire n4671_lo_p_spl_10;
  wire n4671_lo_p_spl_11;
  wire n2643_lo_p_spl_;
  wire n2871_lo_p_spl_;
  wire n4671_lo_n_spl_;
  wire n4671_lo_n_spl_0;
  wire n4671_lo_n_spl_00;
  wire n4671_lo_n_spl_000;
  wire n4671_lo_n_spl_001;
  wire n4671_lo_n_spl_01;
  wire n4671_lo_n_spl_1;
  wire n4671_lo_n_spl_10;
  wire n4671_lo_n_spl_11;
  wire n5636_o2_n_spl_;
  wire n2881_o2_n_spl_;
  wire g1159_n_spl_;
  wire n4695_lo_n_spl_;
  wire n4695_lo_n_spl_0;
  wire n4695_lo_n_spl_00;
  wire n4695_lo_n_spl_000;
  wire n4695_lo_n_spl_0000;
  wire n4695_lo_n_spl_0001;
  wire n4695_lo_n_spl_001;
  wire n4695_lo_n_spl_0010;
  wire n4695_lo_n_spl_0011;
  wire n4695_lo_n_spl_01;
  wire n4695_lo_n_spl_010;
  wire n4695_lo_n_spl_011;
  wire n4695_lo_n_spl_1;
  wire n4695_lo_n_spl_10;
  wire n4695_lo_n_spl_100;
  wire n4695_lo_n_spl_101;
  wire n4695_lo_n_spl_11;
  wire n4695_lo_n_spl_110;
  wire n4695_lo_n_spl_111;
  wire n4695_lo_p_spl_;
  wire n4695_lo_p_spl_0;
  wire n4695_lo_p_spl_00;
  wire n4695_lo_p_spl_000;
  wire n4695_lo_p_spl_0000;
  wire n4695_lo_p_spl_0001;
  wire n4695_lo_p_spl_001;
  wire n4695_lo_p_spl_0010;
  wire n4695_lo_p_spl_0011;
  wire n4695_lo_p_spl_01;
  wire n4695_lo_p_spl_010;
  wire n4695_lo_p_spl_011;
  wire n4695_lo_p_spl_1;
  wire n4695_lo_p_spl_10;
  wire n4695_lo_p_spl_100;
  wire n4695_lo_p_spl_101;
  wire n4695_lo_p_spl_11;
  wire n4695_lo_p_spl_110;
  wire n4695_lo_p_spl_111;
  wire n4707_lo_p_spl_;
  wire n4707_lo_p_spl_0;
  wire n4707_lo_p_spl_00;
  wire n4707_lo_p_spl_000;
  wire n4707_lo_p_spl_001;
  wire n4707_lo_p_spl_01;
  wire n4707_lo_p_spl_1;
  wire n4707_lo_p_spl_10;
  wire n4707_lo_p_spl_11;
  wire n4707_lo_n_spl_;
  wire n4707_lo_n_spl_0;
  wire n4707_lo_n_spl_00;
  wire n4707_lo_n_spl_000;
  wire n4707_lo_n_spl_001;
  wire n4707_lo_n_spl_01;
  wire n4707_lo_n_spl_1;
  wire n4707_lo_n_spl_10;
  wire n4707_lo_n_spl_11;
  wire g1176_n_spl_;
  wire g1183_n_spl_;
  wire g1188_n_spl_;
  wire n2853_o2_n_spl_;
  wire n2853_o2_n_spl_0;
  wire n2853_o2_n_spl_00;
  wire n2853_o2_n_spl_1;
  wire g1201_n_spl_;
  wire n2853_o2_p_spl_;
  wire n2853_o2_p_spl_0;
  wire n2853_o2_p_spl_1;
  wire g1201_p_spl_;
  wire g1205_p_spl_;
  wire g1206_n_spl_;
  wire g1205_n_spl_;
  wire g1206_p_spl_;
  wire n4972_o2_n_spl_;
  wire n4989_o2_p_spl_;
  wire n4972_o2_p_spl_;
  wire n4989_o2_n_spl_;
  wire n5025_o2_n_spl_;
  wire n5093_o2_p_spl_;
  wire n5025_o2_p_spl_;
  wire n5093_o2_n_spl_;
  wire g1215_n_spl_;
  wire g1218_p_spl_;
  wire g1215_p_spl_;
  wire g1218_n_spl_;
  wire n2994_o2_n_spl_;
  wire n2991_o2_p_spl_;
  wire n2994_o2_p_spl_;
  wire n2991_o2_n_spl_;
  wire n4970_o2_p_spl_;
  wire n5024_o2_n_spl_;
  wire n4970_o2_n_spl_;
  wire n5024_o2_p_spl_;
  wire g1224_n_spl_;
  wire g1227_p_spl_;
  wire g1224_p_spl_;
  wire g1227_n_spl_;
  wire g1234_n_spl_;
  wire n3021_o2_n_spl_;
  wire g1243_p_spl_;
  wire g1246_p_spl_;
  wire n3062_o2_p_spl_;
  wire g1250_p_spl_;
  wire g1249_p_spl_;
  wire n4503_lo_n_spl_;
  wire n4503_lo_n_spl_0;
  wire n4503_lo_n_spl_00;
  wire n4503_lo_n_spl_000;
  wire n4503_lo_n_spl_0000;
  wire n4503_lo_n_spl_0001;
  wire n4503_lo_n_spl_001;
  wire n4503_lo_n_spl_0010;
  wire n4503_lo_n_spl_0011;
  wire n4503_lo_n_spl_01;
  wire n4503_lo_n_spl_010;
  wire n4503_lo_n_spl_011;
  wire n4503_lo_n_spl_1;
  wire n4503_lo_n_spl_10;
  wire n4503_lo_n_spl_100;
  wire n4503_lo_n_spl_101;
  wire n4503_lo_n_spl_11;
  wire n4503_lo_n_spl_110;
  wire n4503_lo_n_spl_111;
  wire n4503_lo_p_spl_;
  wire n4503_lo_p_spl_0;
  wire n4503_lo_p_spl_00;
  wire n4503_lo_p_spl_000;
  wire n4503_lo_p_spl_0000;
  wire n4503_lo_p_spl_0001;
  wire n4503_lo_p_spl_001;
  wire n4503_lo_p_spl_0010;
  wire n4503_lo_p_spl_0011;
  wire n4503_lo_p_spl_01;
  wire n4503_lo_p_spl_010;
  wire n4503_lo_p_spl_011;
  wire n4503_lo_p_spl_1;
  wire n4503_lo_p_spl_10;
  wire n4503_lo_p_spl_100;
  wire n4503_lo_p_spl_101;
  wire n4503_lo_p_spl_11;
  wire n4503_lo_p_spl_110;
  wire n4503_lo_p_spl_111;
  wire n4515_lo_n_spl_;
  wire n4515_lo_n_spl_0;
  wire n4515_lo_n_spl_00;
  wire n4515_lo_n_spl_000;
  wire n4515_lo_n_spl_001;
  wire n4515_lo_n_spl_01;
  wire n4515_lo_n_spl_1;
  wire n4515_lo_n_spl_10;
  wire n4515_lo_n_spl_11;
  wire n3579_lo_p_spl_;
  wire n3567_lo_p_spl_;
  wire n4515_lo_p_spl_;
  wire n4515_lo_p_spl_0;
  wire n4515_lo_p_spl_00;
  wire n4515_lo_p_spl_000;
  wire n4515_lo_p_spl_001;
  wire n4515_lo_p_spl_01;
  wire n4515_lo_p_spl_1;
  wire n4515_lo_p_spl_10;
  wire n4515_lo_p_spl_11;
  wire n3375_lo_p_spl_;
  wire n3375_lo_p_spl_0;
  wire n3375_lo_p_spl_00;
  wire n3375_lo_p_spl_000;
  wire n3375_lo_p_spl_0000;
  wire n3375_lo_p_spl_001;
  wire n3375_lo_p_spl_01;
  wire n3375_lo_p_spl_010;
  wire n3375_lo_p_spl_011;
  wire n3375_lo_p_spl_1;
  wire n3375_lo_p_spl_10;
  wire n3375_lo_p_spl_100;
  wire n3375_lo_p_spl_101;
  wire n3375_lo_p_spl_11;
  wire n3375_lo_p_spl_110;
  wire n3375_lo_p_spl_111;
  wire n4527_lo_n_spl_;
  wire n4527_lo_n_spl_0;
  wire n4527_lo_n_spl_00;
  wire n4527_lo_n_spl_000;
  wire n4527_lo_n_spl_0000;
  wire n4527_lo_n_spl_0001;
  wire n4527_lo_n_spl_001;
  wire n4527_lo_n_spl_0010;
  wire n4527_lo_n_spl_0011;
  wire n4527_lo_n_spl_01;
  wire n4527_lo_n_spl_010;
  wire n4527_lo_n_spl_011;
  wire n4527_lo_n_spl_1;
  wire n4527_lo_n_spl_10;
  wire n4527_lo_n_spl_100;
  wire n4527_lo_n_spl_101;
  wire n4527_lo_n_spl_11;
  wire n4527_lo_n_spl_110;
  wire n4527_lo_n_spl_111;
  wire n4527_lo_p_spl_;
  wire n4527_lo_p_spl_0;
  wire n4527_lo_p_spl_00;
  wire n4527_lo_p_spl_000;
  wire n4527_lo_p_spl_0000;
  wire n4527_lo_p_spl_0001;
  wire n4527_lo_p_spl_001;
  wire n4527_lo_p_spl_0010;
  wire n4527_lo_p_spl_0011;
  wire n4527_lo_p_spl_01;
  wire n4527_lo_p_spl_010;
  wire n4527_lo_p_spl_011;
  wire n4527_lo_p_spl_1;
  wire n4527_lo_p_spl_10;
  wire n4527_lo_p_spl_100;
  wire n4527_lo_p_spl_101;
  wire n4527_lo_p_spl_11;
  wire n4527_lo_p_spl_110;
  wire n4527_lo_p_spl_111;
  wire n4539_lo_n_spl_;
  wire n4539_lo_n_spl_0;
  wire n4539_lo_n_spl_00;
  wire n4539_lo_n_spl_000;
  wire n4539_lo_n_spl_001;
  wire n4539_lo_n_spl_01;
  wire n4539_lo_n_spl_1;
  wire n4539_lo_n_spl_10;
  wire n4539_lo_n_spl_11;
  wire n4539_lo_p_spl_;
  wire n4539_lo_p_spl_0;
  wire n4539_lo_p_spl_00;
  wire n4539_lo_p_spl_000;
  wire n4539_lo_p_spl_001;
  wire n4539_lo_p_spl_01;
  wire n4539_lo_p_spl_1;
  wire n4539_lo_p_spl_10;
  wire n4539_lo_p_spl_11;
  wire n2775_lo_p_spl_;
  wire n2799_lo_p_spl_;
  wire g1182_n_spl_;
  wire g1182_n_spl_0;
  wire g1182_n_spl_00;
  wire g1182_n_spl_1;
  wire g1155_n_spl_;
  wire g1155_n_spl_0;
  wire g1155_n_spl_00;
  wire g1155_n_spl_1;
  wire n2679_lo_p_spl_;
  wire n2931_lo_p_spl_;
  wire g1187_n_spl_;
  wire g1187_n_spl_0;
  wire g1187_n_spl_00;
  wire g1187_n_spl_1;
  wire g1158_n_spl_;
  wire g1158_n_spl_0;
  wire g1158_n_spl_00;
  wire g1158_n_spl_1;
  wire n2667_lo_p_spl_;
  wire n2919_lo_p_spl_;
  wire g1194_n_spl_;
  wire g1194_n_spl_0;
  wire g1194_n_spl_00;
  wire g1194_n_spl_1;
  wire g1164_n_spl_;
  wire g1164_n_spl_0;
  wire g1164_n_spl_00;
  wire g1164_n_spl_1;
  wire n2907_lo_n_spl_;
  wire n2895_lo_n_spl_;
  wire g1200_p_spl_;
  wire g1200_p_spl_0;
  wire g1200_p_spl_00;
  wire g1200_p_spl_1;
  wire g1137_p_spl_;
  wire g1137_p_spl_0;
  wire g1137_p_spl_00;
  wire g1137_p_spl_1;
  wire n3519_lo_p_spl_;
  wire n3639_lo_p_spl_;
  wire n3471_lo_n_spl_;
  wire n3591_lo_n_spl_;
  wire n3375_lo_n_spl_;
  wire n3375_lo_n_spl_0;
  wire n3375_lo_n_spl_1;
  wire n3447_lo_p_spl_;
  wire n3459_lo_p_spl_;
  wire n3423_lo_p_spl_;
  wire n3435_lo_p_spl_;
  wire n4659_lo_n_spl_;
  wire n4659_lo_p_spl_;
  wire n3339_lo_n_spl_;
  wire n3339_lo_p_spl_;
  wire n5837_o2_n_spl_;
  wire g1437_n_spl_;
  wire n3795_lo_n_spl_;
  wire n4467_lo_n_spl_;
  wire g1049_n_spl_;
  wire g1054_n_spl_;
  wire g1111_n_spl_;
  wire g1120_n_spl_;
  wire g1212_n_spl_;
  wire g1233_n_spl_;
  wire n3099_lo_p_spl_;
  wire n3111_lo_p_spl_;
  wire g1470_n_spl_;
  wire g1470_n_spl_0;
  wire g1470_n_spl_00;
  wire g1470_n_spl_1;
  wire g1449_n_spl_;
  wire g1449_n_spl_0;
  wire g1449_n_spl_00;
  wire g1449_n_spl_1;
  wire n2823_lo_p_spl_;
  wire n2811_lo_p_spl_;
  wire g1476_n_spl_;
  wire g1476_n_spl_0;
  wire g1476_n_spl_00;
  wire g1476_n_spl_1;
  wire g1453_n_spl_;
  wire g1453_n_spl_0;
  wire g1453_n_spl_00;
  wire g1453_n_spl_1;
  wire n3087_lo_p_spl_;
  wire n3075_lo_p_spl_;
  wire g1482_n_spl_;
  wire g1482_n_spl_0;
  wire g1482_n_spl_00;
  wire g1482_n_spl_1;
  wire g1457_n_spl_;
  wire g1457_n_spl_0;
  wire g1457_n_spl_00;
  wire g1457_n_spl_1;
  wire n2787_lo_p_spl_;
  wire n3039_lo_p_spl_;
  wire g1486_n_spl_;
  wire g1486_n_spl_0;
  wire g1486_n_spl_00;
  wire g1486_n_spl_1;
  wire g1460_n_spl_;
  wire g1460_n_spl_0;
  wire g1460_n_spl_00;
  wire g1460_n_spl_1;
  wire n3531_lo_p_spl_;
  wire n3651_lo_p_spl_;
  wire n3507_lo_p_spl_;
  wire n3627_lo_p_spl_;
  wire n3495_lo_p_spl_;
  wire n3615_lo_p_spl_;
  wire n3483_lo_p_spl_;
  wire n3603_lo_p_spl_;
  wire g1640_n_spl_;
  wire g1639_n_spl_;
  wire g1645_n_spl_;
  wire n2883_lo_n_spl_;
  wire n2655_lo_n_spl_;
  wire g1653_p_spl_;
  wire g1653_p_spl_0;
  wire g1653_p_spl_1;
  wire g1656_p_spl_;
  wire g1656_p_spl_0;
  wire g1656_p_spl_1;
  wire n3555_lo_n_spl_;
  wire n3543_lo_n_spl_;
  wire n2134_inv_n_spl_;
  wire n2134_inv_n_spl_0;
  wire n2134_inv_n_spl_1;
  wire n2718_o2_n_spl_;
  wire n2134_inv_p_spl_;
  wire n2134_inv_p_spl_0;
  wire n2718_o2_p_spl_;
  wire n2718_o2_p_spl_0;
  wire g1690_n_spl_;
  wire n5663_o2_n_spl_;
  wire n5663_o2_n_spl_0;
  wire n5663_o2_n_spl_00;
  wire n5663_o2_n_spl_1;
  wire n2753_o2_n_spl_;
  wire n2628_lo_p_spl_;
  wire n2628_lo_p_spl_0;
  wire n2628_lo_p_spl_1;
  wire n5802_o2_p_spl_;
  wire g1695_n_spl_;
  wire n2715_o2_n_spl_;
  wire n2715_o2_p_spl_;
  wire n2715_o2_p_spl_0;
  wire n3010_o2_n_spl_;
  wire n3010_o2_p_spl_;
  wire n2653_o2_p_spl_;
  wire n2740_o2_p_spl_;
  wire n2740_o2_p_spl_0;
  wire n2736_o2_p_spl_;
  wire n2740_o2_n_spl_;
  wire n2614_inv_p_spl_;
  wire n2614_inv_p_spl_0;
  wire g1703_p_spl_;
  wire g1703_p_spl_0;
  wire n2614_inv_n_spl_;
  wire g1703_n_spl_;
  wire n4632_lo_n_spl_;
  wire n4632_lo_n_spl_0;
  wire n4632_lo_n_spl_00;
  wire n4632_lo_n_spl_000;
  wire n4632_lo_n_spl_001;
  wire n4632_lo_n_spl_01;
  wire n4632_lo_n_spl_010;
  wire n4632_lo_n_spl_011;
  wire n4632_lo_n_spl_1;
  wire n4632_lo_n_spl_10;
  wire n4632_lo_n_spl_11;
  wire n4596_lo_p_spl_;
  wire n4596_lo_p_spl_0;
  wire n4596_lo_p_spl_00;
  wire n4596_lo_p_spl_000;
  wire n4596_lo_p_spl_001;
  wire n4596_lo_p_spl_01;
  wire n4596_lo_p_spl_010;
  wire n4596_lo_p_spl_011;
  wire n4596_lo_p_spl_1;
  wire n4596_lo_p_spl_10;
  wire n4596_lo_p_spl_11;
  wire n5914_o2_p_spl_;
  wire n5914_o2_p_spl_0;
  wire lo382_buf_o2_p_spl_;
  wire lo382_buf_o2_p_spl_0;
  wire lo382_buf_o2_p_spl_00;
  wire lo382_buf_o2_p_spl_01;
  wire lo382_buf_o2_p_spl_1;
  wire n5914_o2_n_spl_;
  wire lo382_buf_o2_n_spl_;
  wire lo382_buf_o2_n_spl_0;
  wire lo382_buf_o2_n_spl_00;
  wire lo382_buf_o2_n_spl_1;
  wire n2629_inv_p_spl_;
  wire n2353_inv_p_spl_;
  wire g1698_n_spl_;
  wire g1698_n_spl_0;
  wire g1698_n_spl_1;
  wire g1698_p_spl_;
  wire g1698_p_spl_0;
  wire n2734_o2_n_spl_;
  wire n2734_o2_p_spl_;
  wire n2689_inv_p_spl_;
  wire n2689_inv_p_spl_0;
  wire n2689_inv_p_spl_1;
  wire n2711_o2_n_spl_;
  wire n2689_inv_n_spl_;
  wire n2689_inv_n_spl_0;
  wire n2711_o2_p_spl_;
  wire lo585_buf_o2_p_spl_;
  wire lo585_buf_o2_p_spl_0;
  wire lo585_buf_o2_p_spl_00;
  wire lo585_buf_o2_p_spl_1;
  wire g1700_n_spl_;
  wire g1700_n_spl_0;
  wire lo585_buf_o2_n_spl_;
  wire lo585_buf_o2_n_spl_0;
  wire lo585_buf_o2_n_spl_1;
  wire g1700_p_spl_;
  wire g1717_n_spl_;
  wire g1717_p_spl_;
  wire g1696_p_spl_;
  wire n5919_o2_p_spl_;
  wire g1723_n_spl_;
  wire n2611_inv_p_spl_;
  wire n2611_inv_p_spl_0;
  wire n2611_inv_p_spl_1;
  wire n2682_o2_p_spl_;
  wire n2682_o2_p_spl_0;
  wire n2682_o2_p_spl_1;
  wire n2611_inv_n_spl_;
  wire n2682_o2_n_spl_;
  wire n5849_o2_p_spl_;
  wire n5849_o2_p_spl_0;
  wire n5598_o2_n_spl_;
  wire n5598_o2_n_spl_0;
  wire n5598_o2_n_spl_1;
  wire n4620_lo_n_spl_;
  wire n4620_lo_n_spl_0;
  wire n4620_lo_n_spl_00;
  wire n4620_lo_n_spl_000;
  wire n4620_lo_n_spl_001;
  wire n4620_lo_n_spl_01;
  wire n4620_lo_n_spl_010;
  wire n4620_lo_n_spl_1;
  wire n4620_lo_n_spl_10;
  wire n4620_lo_n_spl_11;
  wire n5598_o2_p_spl_;
  wire n5598_o2_p_spl_0;
  wire n5598_o2_p_spl_1;
  wire n4608_lo_p_spl_;
  wire n4608_lo_p_spl_0;
  wire n4608_lo_p_spl_00;
  wire n4608_lo_p_spl_000;
  wire n4608_lo_p_spl_001;
  wire n4608_lo_p_spl_01;
  wire n4608_lo_p_spl_010;
  wire n4608_lo_p_spl_1;
  wire n4608_lo_p_spl_10;
  wire n4608_lo_p_spl_11;
  wire n5325_o2_n_spl_;
  wire n5325_o2_n_spl_0;
  wire n5325_o2_p_spl_;
  wire n5325_o2_p_spl_0;
  wire n5833_o2_n_spl_;
  wire n5833_o2_n_spl_0;
  wire n5833_o2_p_spl_;
  wire n5833_o2_p_spl_0;
  wire n4293_lo_p_spl_;
  wire n4293_lo_p_spl_0;
  wire n4293_lo_p_spl_00;
  wire n4293_lo_p_spl_1;
  wire g1711_n_spl_;
  wire g1711_n_spl_0;
  wire n4293_lo_n_spl_;
  wire n4293_lo_n_spl_0;
  wire n4293_lo_n_spl_1;
  wire g1711_p_spl_;
  wire g1756_p_spl_;
  wire lo494_buf_o2_p_spl_;
  wire lo494_buf_o2_p_spl_0;
  wire lo494_buf_o2_p_spl_00;
  wire lo494_buf_o2_p_spl_000;
  wire lo494_buf_o2_p_spl_001;
  wire lo494_buf_o2_p_spl_01;
  wire lo494_buf_o2_p_spl_1;
  wire lo494_buf_o2_p_spl_10;
  wire lo494_buf_o2_p_spl_11;
  wire lo434_buf_o2_p_spl_;
  wire lo494_buf_o2_n_spl_;
  wire lo494_buf_o2_n_spl_0;
  wire lo494_buf_o2_n_spl_00;
  wire lo494_buf_o2_n_spl_000;
  wire lo494_buf_o2_n_spl_01;
  wire lo494_buf_o2_n_spl_1;
  wire lo494_buf_o2_n_spl_10;
  wire lo494_buf_o2_n_spl_11;
  wire lo557_buf_o2_p_spl_;
  wire lo557_buf_o2_p_spl_0;
  wire g1721_n_spl_;
  wire g1721_n_spl_0;
  wire lo573_buf_o2_p_spl_;
  wire lo573_buf_o2_p_spl_0;
  wire g1720_n_spl_;
  wire g1720_n_spl_0;
  wire lo466_buf_o2_p_spl_;
  wire lo490_buf_o2_p_spl_;
  wire lo490_buf_o2_p_spl_0;
  wire lo490_buf_o2_p_spl_00;
  wire lo490_buf_o2_p_spl_000;
  wire lo490_buf_o2_p_spl_001;
  wire lo490_buf_o2_p_spl_01;
  wire lo490_buf_o2_p_spl_010;
  wire lo490_buf_o2_p_spl_011;
  wire lo490_buf_o2_p_spl_1;
  wire lo490_buf_o2_p_spl_10;
  wire lo490_buf_o2_p_spl_11;
  wire lo490_buf_o2_n_spl_;
  wire lo490_buf_o2_n_spl_0;
  wire lo490_buf_o2_n_spl_00;
  wire lo490_buf_o2_n_spl_000;
  wire lo490_buf_o2_n_spl_001;
  wire lo490_buf_o2_n_spl_01;
  wire lo490_buf_o2_n_spl_010;
  wire lo490_buf_o2_n_spl_1;
  wire lo490_buf_o2_n_spl_10;
  wire lo490_buf_o2_n_spl_11;
  wire g1704_p_spl_;
  wire g1719_p_spl_;
  wire g1719_p_spl_0;
  wire g1772_n_spl_;
  wire g1719_n_spl_;
  wire g1772_p_spl_;
  wire g1773_n_spl_;
  wire g1773_p_spl_;
  wire lo357_buf_o2_p_spl_;
  wire lo417_buf_o2_p_spl_;
  wire g1699_p_spl_;
  wire g1699_p_spl_0;
  wire g1781_p_spl_;
  wire g1699_n_spl_;
  wire g1699_n_spl_0;
  wire g1699_n_spl_1;
  wire g1781_n_spl_;
  wire g1712_p_spl_;
  wire g1712_p_spl_0;
  wire g1785_p_spl_;
  wire lo473_buf_o2_p_spl_;
  wire lo536_buf_o2_p_spl_;
  wire lo536_buf_o2_p_spl_0;
  wire g1761_n_spl_;
  wire g1761_n_spl_0;
  wire lo553_buf_o2_p_spl_;
  wire lo553_buf_o2_p_spl_0;
  wire g1722_n_spl_;
  wire g1722_n_spl_0;
  wire g1763_n_spl_;
  wire g1763_n_spl_0;
  wire g1763_n_spl_1;
  wire lo508_buf_o2_p_spl_;
  wire lo512_buf_o2_p_spl_;
  wire n4254_lo_p_spl_;
  wire n4254_lo_p_spl_0;
  wire g1780_n_spl_;
  wire g1780_n_spl_0;
  wire n4314_lo_p_spl_;
  wire n4314_lo_p_spl_0;
  wire g1777_n_spl_;
  wire g1777_n_spl_0;
  wire n4350_lo_p_spl_;
  wire n4350_lo_p_spl_0;
  wire g1790_n_spl_;
  wire g1790_n_spl_0;
  wire lo576_buf_o2_p_spl_;
  wire lo576_buf_o2_p_spl_0;
  wire g1767_n_spl_;
  wire g1767_n_spl_0;
  wire g1807_n_spl_;
  wire g1797_p_spl_;
  wire g1799_p_spl_;
  wire g1799_p_spl_0;
  wire n4728_lo_n_spl_;
  wire n4728_lo_n_spl_0;
  wire n4728_lo_n_spl_00;
  wire n4728_lo_n_spl_000;
  wire n4728_lo_n_spl_001;
  wire n4728_lo_n_spl_01;
  wire n4728_lo_n_spl_010;
  wire n4728_lo_n_spl_1;
  wire n4728_lo_n_spl_10;
  wire n4728_lo_n_spl_11;
  wire n4728_lo_p_spl_;
  wire n4728_lo_p_spl_0;
  wire n4728_lo_p_spl_00;
  wire n4728_lo_p_spl_000;
  wire n4728_lo_p_spl_001;
  wire n4728_lo_p_spl_01;
  wire n4728_lo_p_spl_010;
  wire n4728_lo_p_spl_011;
  wire n4728_lo_p_spl_1;
  wire n4728_lo_p_spl_10;
  wire n4728_lo_p_spl_100;
  wire n4728_lo_p_spl_101;
  wire n4728_lo_p_spl_11;
  wire n5327_o2_n_spl_;
  wire n5327_o2_n_spl_0;
  wire n5327_o2_p_spl_;
  wire n5327_o2_p_spl_0;
  wire n4716_lo_n_spl_;
  wire n4716_lo_n_spl_0;
  wire n3252_lo_p_spl_;
  wire n4716_lo_p_spl_;
  wire n4716_lo_p_spl_0;
  wire n5918_o2_n_spl_;
  wire n5918_o2_p_spl_;
  wire n5920_o2_p_spl_;
  wire n5920_o2_p_spl_0;
  wire n2149_inv_p_spl_;
  wire n3478_o2_p_spl_;
  wire n3484_o2_p_spl_;
  wire n3478_o2_n_spl_;
  wire n3484_o2_n_spl_;
  wire g1831_p_spl_;
  wire g1834_n_spl_;
  wire g1831_n_spl_;
  wire g1834_p_spl_;
  wire n5663_o2_p_spl_;
  wire g1692_p_spl_;
  wire g1692_p_spl_0;
  wire g1840_n_spl_;
  wire g1692_n_spl_;
  wire g1692_n_spl_0;
  wire g1840_p_spl_;
  wire g1755_n_spl_;
  wire g1737_n_spl_;
  wire g1746_n_spl_;
  wire g1854_p_spl_;
  wire g1855_n_spl_;
  wire g1854_n_spl_;
  wire g1855_p_spl_;
  wire n2502_o2_p_spl_;
  wire n2704_inv_p_spl_;
  wire g1859_p_spl_;
  wire g1860_p_spl_;
  wire g1859_n_spl_;
  wire g1860_n_spl_;
  wire n2620_inv_p_spl_;
  wire n2620_inv_p_spl_0;
  wire n2620_inv_p_spl_1;
  wire n2628_lo_n_spl_;
  wire n2620_inv_n_spl_;
  wire n2620_inv_n_spl_0;
  wire n2617_inv_n_spl_;
  wire n2617_inv_n_spl_0;
  wire n2617_inv_n_spl_1;
  wire n2617_inv_p_spl_;
  wire n2617_inv_p_spl_0;
  wire n2617_inv_p_spl_00;
  wire n2617_inv_p_spl_1;
  wire g1872_n_spl_;
  wire g1872_n_spl_0;
  wire g1872_n_spl_00;
  wire g1872_n_spl_1;
  wire g1872_p_spl_;
  wire g1872_p_spl_0;
  wire g1872_p_spl_00;
  wire g1872_p_spl_1;
  wire n3048_o2_p_spl_;
  wire n3048_o2_n_spl_;
  wire n3048_o2_n_spl_0;
  wire g1877_n_spl_;
  wire g1724_p_spl_;
  wire n4188_lo_p_spl_;
  wire n4188_lo_p_spl_0;
  wire g1884_n_spl_;
  wire n2863_o2_p_spl_;
  wire g1693_n_spl_;
  wire g1891_p_spl_;
  wire g1728_n_spl_;
  wire n5823_o2_p_spl_;
  wire g1895_n_spl_;
  wire n4098_lo_p_spl_;
  wire n2591_o2_n_spl_;
  wire n2591_o2_n_spl_0;
  wire g1708_n_spl_;
  wire n5400_o2_p_spl_;
  wire n5400_o2_p_spl_0;
  wire n5400_o2_n_spl_;
  wire n5400_o2_n_spl_0;
  wire n5323_o2_p_spl_;
  wire n5323_o2_p_spl_0;
  wire n5323_o2_n_spl_;
  wire n5323_o2_n_spl_0;
  wire n5402_o2_p_spl_;
  wire n5402_o2_p_spl_0;
  wire n5402_o2_n_spl_;
  wire n5402_o2_n_spl_0;
  wire n5369_o2_n_spl_;
  wire n5369_o2_n_spl_0;
  wire n5369_o2_n_spl_1;
  wire n5369_o2_p_spl_;
  wire n5369_o2_p_spl_0;
  wire n5369_o2_p_spl_1;
  wire n5896_o2_n_spl_;
  wire n5896_o2_n_spl_0;
  wire n5896_o2_n_spl_1;
  wire n5896_o2_p_spl_;
  wire n5896_o2_p_spl_0;
  wire n5896_o2_p_spl_1;
  wire n5600_o2_n_spl_;
  wire n5600_o2_n_spl_0;
  wire n5600_o2_p_spl_;
  wire n5600_o2_p_spl_0;
  wire n5557_o2_n_spl_;
  wire n5557_o2_n_spl_0;
  wire n5557_o2_p_spl_;
  wire n5557_o2_p_spl_0;
  wire n3671_o2_n_spl_;
  wire n3680_o2_p_spl_;
  wire n3671_o2_p_spl_;
  wire n3680_o2_n_spl_;
  wire n3692_o2_n_spl_;
  wire n3692_o2_p_spl_;
  wire n2591_o2_p_spl_;
  wire n2591_o2_p_spl_0;
  wire g1982_n_spl_;
  wire g1985_p_spl_;
  wire g1982_p_spl_;
  wire g1985_n_spl_;
  wire n3707_o2_n_spl_;
  wire n3716_o2_p_spl_;
  wire n3707_o2_p_spl_;
  wire n3716_o2_n_spl_;
  wire n3749_o2_n_spl_;
  wire n3740_o2_n_spl_;
  wire n3749_o2_p_spl_;
  wire n3740_o2_p_spl_;
  wire g1991_p_spl_;
  wire g1994_n_spl_;
  wire g1991_n_spl_;
  wire g1994_p_spl_;
  wire n3936_lo_p_spl_;
  wire n3936_lo_p_spl_0;
  wire n5329_o2_p_spl_;
  wire n3936_lo_n_spl_;
  wire n3936_lo_n_spl_0;
  wire n5329_o2_n_spl_;
  wire n2818_o2_p_spl_;
  wire n2655_o2_p_spl_;
  wire lo450_buf_o2_p_spl_;
  wire g2035_n_spl_;
  wire g2038_p_spl_;
  wire n4188_lo_n_spl_;
  wire n5653_o2_p_spl_;
  wire n5653_o2_n_spl_;
  wire g2046_n_spl_;
  wire g2049_p_spl_;
  wire g2054_n_spl_;
  wire g2057_n_spl_;
  wire g2069_p_spl_;
  wire g2070_n_spl_;
  wire g2069_n_spl_;
  wire g2070_p_spl_;
  wire n4488_lo_n_spl_;
  wire n4488_lo_n_spl_0;
  wire n4488_lo_n_spl_1;
  wire n4488_lo_p_spl_;
  wire n4488_lo_p_spl_0;
  wire n4488_lo_p_spl_1;
  wire g2075_p_spl_;
  wire g2076_p_spl_;
  wire g2075_n_spl_;
  wire g2076_n_spl_;
  wire g2082_n_spl_;
  wire g2082_p_spl_;
  wire g2085_p_spl_;
  wire g2085_n_spl_;
  wire g1793_p_spl_;
  wire g1796_p_spl_;
  wire g1796_p_spl_0;
  wire g1762_p_spl_;
  wire n5936_o2_n_spl_;
  wire lo398_buf_o2_n_spl_;
  wire lo398_buf_o2_n_spl_0;
  wire lo398_buf_o2_n_spl_00;
  wire lo398_buf_o2_n_spl_000;
  wire lo398_buf_o2_n_spl_001;
  wire lo398_buf_o2_n_spl_01;
  wire lo398_buf_o2_n_spl_010;
  wire lo398_buf_o2_n_spl_011;
  wire lo398_buf_o2_n_spl_1;
  wire lo398_buf_o2_n_spl_10;
  wire lo398_buf_o2_n_spl_100;
  wire lo398_buf_o2_n_spl_101;
  wire lo398_buf_o2_n_spl_11;
  wire lo398_buf_o2_n_spl_110;
  wire lo398_buf_o2_n_spl_111;
  wire n5936_o2_p_spl_;
  wire n5936_o2_p_spl_0;
  wire lo402_buf_o2_n_spl_;
  wire lo402_buf_o2_n_spl_0;
  wire lo402_buf_o2_n_spl_00;
  wire lo402_buf_o2_n_spl_000;
  wire lo402_buf_o2_n_spl_001;
  wire lo402_buf_o2_n_spl_01;
  wire lo402_buf_o2_n_spl_010;
  wire lo402_buf_o2_n_spl_011;
  wire lo402_buf_o2_n_spl_1;
  wire lo402_buf_o2_n_spl_10;
  wire lo402_buf_o2_n_spl_100;
  wire lo402_buf_o2_n_spl_101;
  wire lo402_buf_o2_n_spl_11;
  wire lo402_buf_o2_n_spl_110;
  wire lo406_buf_o2_p_spl_;
  wire lo406_buf_o2_p_spl_0;
  wire lo406_buf_o2_p_spl_00;
  wire lo406_buf_o2_p_spl_000;
  wire lo406_buf_o2_p_spl_001;
  wire lo406_buf_o2_p_spl_01;
  wire lo406_buf_o2_p_spl_010;
  wire lo406_buf_o2_p_spl_011;
  wire lo406_buf_o2_p_spl_1;
  wire lo406_buf_o2_p_spl_10;
  wire lo406_buf_o2_p_spl_100;
  wire lo406_buf_o2_p_spl_101;
  wire lo406_buf_o2_p_spl_11;
  wire lo390_buf_o2_p_spl_;
  wire lo390_buf_o2_p_spl_0;
  wire lo390_buf_o2_p_spl_00;
  wire lo390_buf_o2_p_spl_000;
  wire lo390_buf_o2_p_spl_001;
  wire lo390_buf_o2_p_spl_01;
  wire lo390_buf_o2_p_spl_010;
  wire lo390_buf_o2_p_spl_011;
  wire lo390_buf_o2_p_spl_1;
  wire lo390_buf_o2_p_spl_10;
  wire lo390_buf_o2_p_spl_100;
  wire lo390_buf_o2_p_spl_101;
  wire lo390_buf_o2_p_spl_11;
  wire lo390_buf_o2_p_spl_110;
  wire lo474_buf_o2_n_spl_;
  wire lo474_buf_o2_p_spl_;
  wire lo474_buf_o2_p_spl_0;
  wire lo518_buf_o2_p_spl_;
  wire lo458_buf_o2_p_spl_;
  wire n3957_lo_p_spl_;
  wire n3957_lo_p_spl_0;
  wire n3834_lo_p_spl_;
  wire n4110_lo_p_spl_;
  wire n4122_lo_p_spl_;
  wire n2811_o2_p_spl_;
  wire n2811_o2_p_spl_0;
  wire n2811_o2_p_spl_1;
  wire n2811_o2_n_spl_;
  wire n2811_o2_n_spl_0;
  wire n2811_o2_n_spl_1;
  wire n2740_inv_p_spl_;
  wire g1758_p_spl_;
  wire g1758_p_spl_0;
  wire g2139_n_spl_;
  wire g2139_n_spl_0;
  wire n2779_inv_n_spl_;
  wire n2779_inv_n_spl_0;
  wire n2779_inv_n_spl_1;
  wire g1725_n_spl_;
  wire g1758_n_spl_;
  wire g1758_n_spl_0;
  wire g1758_n_spl_1;
  wire g2142_n_spl_;
  wire n2317_inv_n_spl_;
  wire n2317_inv_p_spl_;
  wire n2317_inv_p_spl_0;
  wire n2572_inv_n_spl_;
  wire n2572_inv_n_spl_0;
  wire g2146_p_spl_;
  wire n2572_inv_p_spl_;
  wire n2572_inv_p_spl_0;
  wire n2572_inv_p_spl_1;
  wire g2146_n_spl_;
  wire n2689_o2_p_spl_;
  wire n2638_inv_p_spl_;
  wire n2779_inv_p_spl_;
  wire n2779_inv_p_spl_0;
  wire n2779_inv_p_spl_1;
  wire g2139_p_spl_;
  wire g2139_p_spl_0;
  wire g2151_n_spl_;
  wire g2151_n_spl_0;
  wire g2151_p_spl_;
  wire g2151_p_spl_0;
  wire g2157_n_spl_;
  wire g1702_n_spl_;
  wire g1702_n_spl_0;
  wire g2161_p_spl_;
  wire g1702_p_spl_;
  wire g2161_n_spl_;
  wire n2323_inv_n_spl_;
  wire n2323_inv_p_spl_;
  wire n2323_inv_p_spl_0;
  wire n2323_inv_p_spl_1;
  wire g2164_n_spl_;
  wire g2165_p_spl_;
  wire g1705_p_spl_;
  wire n2662_o2_p_spl_;
  wire n2662_o2_p_spl_0;
  wire g2169_n_spl_;
  wire n2662_o2_n_spl_;
  wire g2169_p_spl_;
  wire g2167_n_spl_;
  wire g2172_n_spl_;
  wire g2172_n_spl_0;
  wire g2096_n_spl_;
  wire g1805_p_spl_;
  wire g1808_p_spl_;
  wire n5938_o2_p_spl_;
  wire n3969_lo_p_spl_;
  wire n5912_o2_n_spl_;
  wire n5912_o2_p_spl_;
  wire n5912_o2_p_spl_0;
  wire lo554_buf_o2_p_spl_;
  wire n5910_o2_n_spl_;
  wire n5910_o2_p_spl_;
  wire n5910_o2_p_spl_0;
  wire lo558_buf_o2_p_spl_;
  wire n5908_o2_n_spl_;
  wire n5908_o2_p_spl_;
  wire n5908_o2_p_spl_0;
  wire lo574_buf_o2_p_spl_;
  wire n5934_o2_n_spl_;
  wire n5934_o2_p_spl_;
  wire n5934_o2_p_spl_0;
  wire lo538_buf_o2_p_spl_;
  wire lo418_buf_o2_n_spl_;
  wire lo418_buf_o2_p_spl_;
  wire lo418_buf_o2_p_spl_0;
  wire lo550_buf_o2_p_spl_;
  wire lo358_buf_o2_n_spl_;
  wire lo358_buf_o2_p_spl_;
  wire lo358_buf_o2_p_spl_0;
  wire lo570_buf_o2_p_spl_;
  wire lo350_buf_o2_n_spl_;
  wire lo350_buf_o2_p_spl_;
  wire lo350_buf_o2_p_spl_0;
  wire g1714_n_spl_;
  wire g1714_n_spl_0;
  wire g1714_p_spl_;
  wire n2694_o2_p_spl_;
  wire g2253_n_spl_;
  wire n2694_o2_n_spl_;
  wire g2253_p_spl_;
  wire g2250_p_spl_;
  wire g2259_n_spl_;
  wire n3654_lo_p_spl_;
  wire g1768_n_spl_;
  wire g2269_p_spl_;
  wire g2272_p_spl_;
  wire g1764_p_spl_;
  wire g1764_p_spl_0;
  wire g1809_p_spl_;
  wire g2099_p_spl_;
  wire g2099_p_spl_0;
  wire g2275_n_spl_;
  wire g2108_n_spl_;
  wire g2108_n_spl_0;
  wire g2123_n_spl_;
  wire g2123_n_spl_0;
  wire g2117_n_spl_;
  wire g2117_n_spl_0;
  wire g2126_p_spl_;
  wire g2126_p_spl_0;
  wire lo590_buf_o2_p_spl_;
  wire lo590_buf_o2_p_spl_0;
  wire lo590_buf_o2_n_spl_;
  wire lo398_buf_o2_p_spl_;
  wire lo398_buf_o2_p_spl_0;
  wire lo398_buf_o2_p_spl_00;
  wire lo398_buf_o2_p_spl_1;
  wire lo390_buf_o2_n_spl_;
  wire lo390_buf_o2_n_spl_0;
  wire lo390_buf_o2_n_spl_00;
  wire lo390_buf_o2_n_spl_1;
  wire lo482_buf_o2_n_spl_;
  wire lo482_buf_o2_n_spl_0;
  wire lo482_buf_o2_n_spl_1;
  wire lo482_buf_o2_p_spl_;
  wire lo482_buf_o2_p_spl_0;
  wire lo482_buf_o2_p_spl_00;
  wire lo482_buf_o2_p_spl_1;
  wire lo402_buf_o2_p_spl_;
  wire lo402_buf_o2_p_spl_0;
  wire lo402_buf_o2_p_spl_1;
  wire lo406_buf_o2_n_spl_;
  wire lo406_buf_o2_n_spl_0;
  wire lo406_buf_o2_n_spl_1;
  wire g2120_n_spl_;
  wire g2120_n_spl_0;
  wire g2295_n_spl_;
  wire lo510_buf_o2_n_spl_;
  wire lo510_buf_o2_p_spl_;
  wire lo510_buf_o2_p_spl_0;
  wire lo598_buf_o2_p_spl_;
  wire lo502_buf_o2_p_spl_;
  wire lo502_buf_o2_p_spl_0;
  wire lo502_buf_o2_n_spl_;
  wire lo594_buf_o2_p_spl_;
  wire g2306_n_spl_;
  wire g2315_p_spl_;
  wire n2641_inv_p_spl_;
  wire g1774_n_spl_;
  wire g1787_n_spl_;
  wire g1697_n_spl_;
  wire g1697_n_spl_0;
  wire g1701_p_spl_;
  wire g1697_p_spl_;
  wire g1701_n_spl_;
  wire g1701_n_spl_0;
  wire lo410_buf_o2_n_spl_;
  wire lo410_buf_o2_n_spl_0;
  wire lo410_buf_o2_n_spl_1;
  wire lo410_buf_o2_p_spl_;
  wire lo410_buf_o2_p_spl_0;
  wire lo410_buf_o2_p_spl_00;
  wire lo410_buf_o2_p_spl_1;
  wire lo546_buf_o2_p_spl_;
  wire lo546_buf_o2_p_spl_0;
  wire lo546_buf_o2_n_spl_;
  wire n4545_lo_n_spl_;
  wire n4545_lo_p_spl_;
  wire g1716_n_spl_;
  wire g1792_p_spl_;
  wire n4386_lo_p_spl_;
  wire g2132_n_spl_;
  wire n4398_lo_p_spl_;
  wire g1802_n_spl_;
  wire g2133_n_spl_;
  wire n3978_lo_p_spl_;
  wire n4050_lo_p_spl_;
  wire g2276_n_spl_;
  wire g2276_n_spl_0;
  wire g2137_p_spl_;
  wire g2137_p_spl_0;
  wire g2137_p_spl_1;
  wire g2160_n_spl_;
  wire g2160_n_spl_0;
  wire g2175_p_spl_;
  wire g2098_n_spl_;
  wire g2135_p_spl_;
  wire g1803_p_spl_;
  wire g1804_p_spl_;
  wire g2177_n_spl_;
  wire n4302_lo_p_spl_;
  wire n4302_lo_p_spl_0;
  wire g2264_n_spl_;
  wire g2264_n_spl_0;
  wire g2267_p_spl_;
  wire g2365_p_spl_;
  wire n4374_lo_p_spl_;
  wire g1898_n_spl_;
  wire g2268_n_spl_;
  wire n4242_lo_p_spl_;
  wire g2129_n_spl_;
  wire g2361_n_spl_;
  wire g2362_n_spl_;
  wire g2363_n_spl_;
  wire G92_p_spl_;
  wire G124_p_spl_;
  wire G124_p_spl_0;
  wire G124_p_spl_1;
  wire G124_n_spl_;
  wire G124_n_spl_0;
  wire G94_p_spl_;
  wire G107_p_spl_;
  wire n4419_lo_n_spl_;
  wire n4419_lo_n_spl_0;
  wire n4431_lo_p_spl_;
  wire n2619_lo_n_spl_;
  wire n2619_lo_n_spl_0;
  wire n2619_lo_n_spl_1;
  wire n3975_lo_n_spl_;
  wire g1064_n_spl_;
  wire g1102_n_spl_;
  wire g1106_p_spl_;
  wire g1126_p_spl_;
  wire g1127_n_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  buf

  (
    G42_p,
    G42
  );


  not

  (
    G42_n,
    G42
  );


  buf

  (
    G43_p,
    G43
  );


  not

  (
    G43_n,
    G43
  );


  buf

  (
    G44_p,
    G44
  );


  not

  (
    G44_n,
    G44
  );


  buf

  (
    G45_p,
    G45
  );


  not

  (
    G45_n,
    G45
  );


  buf

  (
    G46_p,
    G46
  );


  not

  (
    G46_n,
    G46
  );


  buf

  (
    G47_p,
    G47
  );


  not

  (
    G47_n,
    G47
  );


  buf

  (
    G48_p,
    G48
  );


  not

  (
    G48_n,
    G48
  );


  buf

  (
    G49_p,
    G49
  );


  not

  (
    G49_n,
    G49
  );


  buf

  (
    G50_p,
    G50
  );


  not

  (
    G50_n,
    G50
  );


  buf

  (
    G51_p,
    G51
  );


  not

  (
    G51_n,
    G51
  );


  buf

  (
    G52_p,
    G52
  );


  not

  (
    G52_n,
    G52
  );


  buf

  (
    G53_p,
    G53
  );


  not

  (
    G53_n,
    G53
  );


  buf

  (
    G54_p,
    G54
  );


  not

  (
    G54_n,
    G54
  );


  buf

  (
    G55_p,
    G55
  );


  not

  (
    G55_n,
    G55
  );


  buf

  (
    G56_p,
    G56
  );


  not

  (
    G56_n,
    G56
  );


  buf

  (
    G57_p,
    G57
  );


  not

  (
    G57_n,
    G57
  );


  buf

  (
    G58_p,
    G58
  );


  not

  (
    G58_n,
    G58
  );


  buf

  (
    G59_p,
    G59
  );


  not

  (
    G59_n,
    G59
  );


  buf

  (
    G60_p,
    G60
  );


  not

  (
    G60_n,
    G60
  );


  buf

  (
    G61_p,
    G61
  );


  not

  (
    G61_n,
    G61
  );


  buf

  (
    G62_p,
    G62
  );


  not

  (
    G62_n,
    G62
  );


  buf

  (
    G63_p,
    G63
  );


  not

  (
    G63_n,
    G63
  );


  buf

  (
    G64_p,
    G64
  );


  not

  (
    G64_n,
    G64
  );


  buf

  (
    G65_p,
    G65
  );


  not

  (
    G65_n,
    G65
  );


  buf

  (
    G66_p,
    G66
  );


  not

  (
    G66_n,
    G66
  );


  buf

  (
    G67_p,
    G67
  );


  not

  (
    G67_n,
    G67
  );


  buf

  (
    G68_p,
    G68
  );


  not

  (
    G68_n,
    G68
  );


  buf

  (
    G69_p,
    G69
  );


  not

  (
    G69_n,
    G69
  );


  buf

  (
    G70_p,
    G70
  );


  not

  (
    G70_n,
    G70
  );


  buf

  (
    G71_p,
    G71
  );


  not

  (
    G71_n,
    G71
  );


  buf

  (
    G72_p,
    G72
  );


  not

  (
    G72_n,
    G72
  );


  buf

  (
    G73_p,
    G73
  );


  not

  (
    G73_n,
    G73
  );


  buf

  (
    G74_p,
    G74
  );


  not

  (
    G74_n,
    G74
  );


  buf

  (
    G75_p,
    G75
  );


  not

  (
    G75_n,
    G75
  );


  buf

  (
    G76_p,
    G76
  );


  not

  (
    G76_n,
    G76
  );


  buf

  (
    G77_p,
    G77
  );


  not

  (
    G77_n,
    G77
  );


  buf

  (
    G78_p,
    G78
  );


  not

  (
    G78_n,
    G78
  );


  buf

  (
    G79_p,
    G79
  );


  not

  (
    G79_n,
    G79
  );


  buf

  (
    G80_p,
    G80
  );


  not

  (
    G80_n,
    G80
  );


  buf

  (
    G81_p,
    G81
  );


  not

  (
    G81_n,
    G81
  );


  buf

  (
    G82_p,
    G82
  );


  not

  (
    G82_n,
    G82
  );


  buf

  (
    G83_p,
    G83
  );


  not

  (
    G83_n,
    G83
  );


  buf

  (
    G84_p,
    G84
  );


  not

  (
    G84_n,
    G84
  );


  buf

  (
    G85_p,
    G85
  );


  not

  (
    G85_n,
    G85
  );


  buf

  (
    G86_p,
    G86
  );


  not

  (
    G86_n,
    G86
  );


  buf

  (
    G87_p,
    G87
  );


  not

  (
    G87_n,
    G87
  );


  buf

  (
    G88_p,
    G88
  );


  not

  (
    G88_n,
    G88
  );


  buf

  (
    G89_p,
    G89
  );


  not

  (
    G89_n,
    G89
  );


  buf

  (
    G90_p,
    G90
  );


  not

  (
    G90_n,
    G90
  );


  buf

  (
    G91_p,
    G91
  );


  not

  (
    G91_n,
    G91
  );


  buf

  (
    G92_p,
    G92
  );


  not

  (
    G92_n,
    G92
  );


  buf

  (
    G93_p,
    G93
  );


  not

  (
    G93_n,
    G93
  );


  buf

  (
    G94_p,
    G94
  );


  not

  (
    G94_n,
    G94
  );


  buf

  (
    G95_p,
    G95
  );


  not

  (
    G95_n,
    G95
  );


  buf

  (
    G96_p,
    G96
  );


  not

  (
    G96_n,
    G96
  );


  buf

  (
    G97_p,
    G97
  );


  not

  (
    G97_n,
    G97
  );


  buf

  (
    G98_p,
    G98
  );


  not

  (
    G98_n,
    G98
  );


  buf

  (
    G99_p,
    G99
  );


  not

  (
    G99_n,
    G99
  );


  buf

  (
    G100_p,
    G100
  );


  not

  (
    G100_n,
    G100
  );


  buf

  (
    G101_p,
    G101
  );


  not

  (
    G101_n,
    G101
  );


  buf

  (
    G102_p,
    G102
  );


  not

  (
    G102_n,
    G102
  );


  buf

  (
    G103_p,
    G103
  );


  not

  (
    G103_n,
    G103
  );


  buf

  (
    G104_p,
    G104
  );


  not

  (
    G104_n,
    G104
  );


  buf

  (
    G105_p,
    G105
  );


  not

  (
    G105_n,
    G105
  );


  buf

  (
    G106_p,
    G106
  );


  not

  (
    G106_n,
    G106
  );


  buf

  (
    G107_p,
    G107
  );


  not

  (
    G107_n,
    G107
  );


  buf

  (
    G108_p,
    G108
  );


  not

  (
    G108_n,
    G108
  );


  buf

  (
    G109_p,
    G109
  );


  not

  (
    G109_n,
    G109
  );


  buf

  (
    G110_p,
    G110
  );


  not

  (
    G110_n,
    G110
  );


  buf

  (
    G111_p,
    G111
  );


  not

  (
    G111_n,
    G111
  );


  buf

  (
    G112_p,
    G112
  );


  not

  (
    G112_n,
    G112
  );


  buf

  (
    G113_p,
    G113
  );


  not

  (
    G113_n,
    G113
  );


  buf

  (
    G114_p,
    G114
  );


  not

  (
    G114_n,
    G114
  );


  buf

  (
    G115_p,
    G115
  );


  not

  (
    G115_n,
    G115
  );


  buf

  (
    G116_p,
    G116
  );


  not

  (
    G116_n,
    G116
  );


  buf

  (
    G117_p,
    G117
  );


  not

  (
    G117_n,
    G117
  );


  buf

  (
    G118_p,
    G118
  );


  not

  (
    G118_n,
    G118
  );


  buf

  (
    G119_p,
    G119
  );


  not

  (
    G119_n,
    G119
  );


  buf

  (
    G120_p,
    G120
  );


  not

  (
    G120_n,
    G120
  );


  buf

  (
    G121_p,
    G121
  );


  not

  (
    G121_n,
    G121
  );


  buf

  (
    G122_p,
    G122
  );


  not

  (
    G122_n,
    G122
  );


  buf

  (
    G123_p,
    G123
  );


  not

  (
    G123_n,
    G123
  );


  buf

  (
    G124_p,
    G124
  );


  not

  (
    G124_n,
    G124
  );


  buf

  (
    G125_p,
    G125
  );


  not

  (
    G125_n,
    G125
  );


  buf

  (
    G126_p,
    G126
  );


  not

  (
    G126_n,
    G126
  );


  buf

  (
    G127_p,
    G127
  );


  not

  (
    G127_n,
    G127
  );


  buf

  (
    G128_p,
    G128
  );


  not

  (
    G128_n,
    G128
  );


  buf

  (
    G129_p,
    G129
  );


  not

  (
    G129_n,
    G129
  );


  buf

  (
    G130_p,
    G130
  );


  not

  (
    G130_n,
    G130
  );


  buf

  (
    G131_p,
    G131
  );


  not

  (
    G131_n,
    G131
  );


  buf

  (
    G132_p,
    G132
  );


  not

  (
    G132_n,
    G132
  );


  buf

  (
    G133_p,
    G133
  );


  not

  (
    G133_n,
    G133
  );


  buf

  (
    G134_p,
    G134
  );


  not

  (
    G134_n,
    G134
  );


  buf

  (
    G135_p,
    G135
  );


  not

  (
    G135_n,
    G135
  );


  buf

  (
    G136_p,
    G136
  );


  not

  (
    G136_n,
    G136
  );


  buf

  (
    G137_p,
    G137
  );


  not

  (
    G137_n,
    G137
  );


  buf

  (
    G138_p,
    G138
  );


  not

  (
    G138_n,
    G138
  );


  buf

  (
    G139_p,
    G139
  );


  not

  (
    G139_n,
    G139
  );


  buf

  (
    G140_p,
    G140
  );


  not

  (
    G140_n,
    G140
  );


  buf

  (
    G141_p,
    G141
  );


  not

  (
    G141_n,
    G141
  );


  buf

  (
    G142_p,
    G142
  );


  not

  (
    G142_n,
    G142
  );


  buf

  (
    G143_p,
    G143
  );


  not

  (
    G143_n,
    G143
  );


  buf

  (
    G144_p,
    G144
  );


  not

  (
    G144_n,
    G144
  );


  buf

  (
    G145_p,
    G145
  );


  not

  (
    G145_n,
    G145
  );


  buf

  (
    G146_p,
    G146
  );


  not

  (
    G146_n,
    G146
  );


  buf

  (
    G147_p,
    G147
  );


  not

  (
    G147_n,
    G147
  );


  buf

  (
    G148_p,
    G148
  );


  not

  (
    G148_n,
    G148
  );


  buf

  (
    G149_p,
    G149
  );


  not

  (
    G149_n,
    G149
  );


  buf

  (
    G150_p,
    G150
  );


  not

  (
    G150_n,
    G150
  );


  buf

  (
    G151_p,
    G151
  );


  not

  (
    G151_n,
    G151
  );


  buf

  (
    G152_p,
    G152
  );


  not

  (
    G152_n,
    G152
  );


  buf

  (
    G153_p,
    G153
  );


  not

  (
    G153_n,
    G153
  );


  buf

  (
    G154_p,
    G154
  );


  not

  (
    G154_n,
    G154
  );


  buf

  (
    G155_p,
    G155
  );


  not

  (
    G155_n,
    G155
  );


  buf

  (
    G156_p,
    G156
  );


  not

  (
    G156_n,
    G156
  );


  buf

  (
    G157_p,
    G157
  );


  not

  (
    G157_n,
    G157
  );


  buf

  (
    G158_p,
    G158
  );


  not

  (
    G158_n,
    G158
  );


  buf

  (
    G159_p,
    G159
  );


  not

  (
    G159_n,
    G159
  );


  buf

  (
    G160_p,
    G160
  );


  not

  (
    G160_n,
    G160
  );


  buf

  (
    G161_p,
    G161
  );


  not

  (
    G161_n,
    G161
  );


  buf

  (
    G162_p,
    G162
  );


  not

  (
    G162_n,
    G162
  );


  buf

  (
    G163_p,
    G163
  );


  not

  (
    G163_n,
    G163
  );


  buf

  (
    G164_p,
    G164
  );


  not

  (
    G164_n,
    G164
  );


  buf

  (
    G165_p,
    G165
  );


  not

  (
    G165_n,
    G165
  );


  buf

  (
    G166_p,
    G166
  );


  not

  (
    G166_n,
    G166
  );


  buf

  (
    G167_p,
    G167
  );


  not

  (
    G167_n,
    G167
  );


  buf

  (
    G168_p,
    G168
  );


  not

  (
    G168_n,
    G168
  );


  buf

  (
    G169_p,
    G169
  );


  not

  (
    G169_n,
    G169
  );


  buf

  (
    G170_p,
    G170
  );


  not

  (
    G170_n,
    G170
  );


  buf

  (
    G171_p,
    G171
  );


  not

  (
    G171_n,
    G171
  );


  buf

  (
    G172_p,
    G172
  );


  not

  (
    G172_n,
    G172
  );


  buf

  (
    G173_p,
    G173
  );


  not

  (
    G173_n,
    G173
  );


  buf

  (
    G174_p,
    G174
  );


  not

  (
    G174_n,
    G174
  );


  buf

  (
    G175_p,
    G175
  );


  not

  (
    G175_n,
    G175
  );


  buf

  (
    G176_p,
    G176
  );


  not

  (
    G176_n,
    G176
  );


  buf

  (
    G177_p,
    G177
  );


  not

  (
    G177_n,
    G177
  );


  buf

  (
    G178_p,
    G178
  );


  not

  (
    G178_n,
    G178
  );


  buf

  (
    n2610_lo_p,
    n2610_lo
  );


  not

  (
    n2610_lo_n,
    n2610_lo
  );


  buf

  (
    n2613_lo_p,
    n2613_lo
  );


  not

  (
    n2613_lo_n,
    n2613_lo
  );


  buf

  (
    n2616_lo_p,
    n2616_lo
  );


  not

  (
    n2616_lo_n,
    n2616_lo
  );


  buf

  (
    n2619_lo_p,
    n2619_lo
  );


  not

  (
    n2619_lo_n,
    n2619_lo
  );


  buf

  (
    n2622_lo_p,
    n2622_lo
  );


  not

  (
    n2622_lo_n,
    n2622_lo
  );


  buf

  (
    n2625_lo_p,
    n2625_lo
  );


  not

  (
    n2625_lo_n,
    n2625_lo
  );


  buf

  (
    n2628_lo_p,
    n2628_lo
  );


  not

  (
    n2628_lo_n,
    n2628_lo
  );


  buf

  (
    n2634_lo_p,
    n2634_lo
  );


  not

  (
    n2634_lo_n,
    n2634_lo
  );


  buf

  (
    n2637_lo_p,
    n2637_lo
  );


  not

  (
    n2637_lo_n,
    n2637_lo
  );


  buf

  (
    n2640_lo_p,
    n2640_lo
  );


  not

  (
    n2640_lo_n,
    n2640_lo
  );


  buf

  (
    n2643_lo_p,
    n2643_lo
  );


  not

  (
    n2643_lo_n,
    n2643_lo
  );


  buf

  (
    n2646_lo_p,
    n2646_lo
  );


  not

  (
    n2646_lo_n,
    n2646_lo
  );


  buf

  (
    n2649_lo_p,
    n2649_lo
  );


  not

  (
    n2649_lo_n,
    n2649_lo
  );


  buf

  (
    n2652_lo_p,
    n2652_lo
  );


  not

  (
    n2652_lo_n,
    n2652_lo
  );


  buf

  (
    n2655_lo_p,
    n2655_lo
  );


  not

  (
    n2655_lo_n,
    n2655_lo
  );


  buf

  (
    n2658_lo_p,
    n2658_lo
  );


  not

  (
    n2658_lo_n,
    n2658_lo
  );


  buf

  (
    n2661_lo_p,
    n2661_lo
  );


  not

  (
    n2661_lo_n,
    n2661_lo
  );


  buf

  (
    n2664_lo_p,
    n2664_lo
  );


  not

  (
    n2664_lo_n,
    n2664_lo
  );


  buf

  (
    n2667_lo_p,
    n2667_lo
  );


  not

  (
    n2667_lo_n,
    n2667_lo
  );


  buf

  (
    n2670_lo_p,
    n2670_lo
  );


  not

  (
    n2670_lo_n,
    n2670_lo
  );


  buf

  (
    n2673_lo_p,
    n2673_lo
  );


  not

  (
    n2673_lo_n,
    n2673_lo
  );


  buf

  (
    n2676_lo_p,
    n2676_lo
  );


  not

  (
    n2676_lo_n,
    n2676_lo
  );


  buf

  (
    n2679_lo_p,
    n2679_lo
  );


  not

  (
    n2679_lo_n,
    n2679_lo
  );


  buf

  (
    n2682_lo_p,
    n2682_lo
  );


  not

  (
    n2682_lo_n,
    n2682_lo
  );


  buf

  (
    n2685_lo_p,
    n2685_lo
  );


  not

  (
    n2685_lo_n,
    n2685_lo
  );


  buf

  (
    n2688_lo_p,
    n2688_lo
  );


  not

  (
    n2688_lo_n,
    n2688_lo
  );


  buf

  (
    n2691_lo_p,
    n2691_lo
  );


  not

  (
    n2691_lo_n,
    n2691_lo
  );


  buf

  (
    n2694_lo_p,
    n2694_lo
  );


  not

  (
    n2694_lo_n,
    n2694_lo
  );


  buf

  (
    n2697_lo_p,
    n2697_lo
  );


  not

  (
    n2697_lo_n,
    n2697_lo
  );


  buf

  (
    n2700_lo_p,
    n2700_lo
  );


  not

  (
    n2700_lo_n,
    n2700_lo
  );


  buf

  (
    n2703_lo_p,
    n2703_lo
  );


  not

  (
    n2703_lo_n,
    n2703_lo
  );


  buf

  (
    n2706_lo_p,
    n2706_lo
  );


  not

  (
    n2706_lo_n,
    n2706_lo
  );


  buf

  (
    n2709_lo_p,
    n2709_lo
  );


  not

  (
    n2709_lo_n,
    n2709_lo
  );


  buf

  (
    n2712_lo_p,
    n2712_lo
  );


  not

  (
    n2712_lo_n,
    n2712_lo
  );


  buf

  (
    n2715_lo_p,
    n2715_lo
  );


  not

  (
    n2715_lo_n,
    n2715_lo
  );


  buf

  (
    n2718_lo_p,
    n2718_lo
  );


  not

  (
    n2718_lo_n,
    n2718_lo
  );


  buf

  (
    n2721_lo_p,
    n2721_lo
  );


  not

  (
    n2721_lo_n,
    n2721_lo
  );


  buf

  (
    n2724_lo_p,
    n2724_lo
  );


  not

  (
    n2724_lo_n,
    n2724_lo
  );


  buf

  (
    n2727_lo_p,
    n2727_lo
  );


  not

  (
    n2727_lo_n,
    n2727_lo
  );


  buf

  (
    n2730_lo_p,
    n2730_lo
  );


  not

  (
    n2730_lo_n,
    n2730_lo
  );


  buf

  (
    n2733_lo_p,
    n2733_lo
  );


  not

  (
    n2733_lo_n,
    n2733_lo
  );


  buf

  (
    n2736_lo_p,
    n2736_lo
  );


  not

  (
    n2736_lo_n,
    n2736_lo
  );


  buf

  (
    n2739_lo_p,
    n2739_lo
  );


  not

  (
    n2739_lo_n,
    n2739_lo
  );


  buf

  (
    n2742_lo_p,
    n2742_lo
  );


  not

  (
    n2742_lo_n,
    n2742_lo
  );


  buf

  (
    n2745_lo_p,
    n2745_lo
  );


  not

  (
    n2745_lo_n,
    n2745_lo
  );


  buf

  (
    n2748_lo_p,
    n2748_lo
  );


  not

  (
    n2748_lo_n,
    n2748_lo
  );


  buf

  (
    n2751_lo_p,
    n2751_lo
  );


  not

  (
    n2751_lo_n,
    n2751_lo
  );


  buf

  (
    n2754_lo_p,
    n2754_lo
  );


  not

  (
    n2754_lo_n,
    n2754_lo
  );


  buf

  (
    n2757_lo_p,
    n2757_lo
  );


  not

  (
    n2757_lo_n,
    n2757_lo
  );


  buf

  (
    n2760_lo_p,
    n2760_lo
  );


  not

  (
    n2760_lo_n,
    n2760_lo
  );


  buf

  (
    n2763_lo_p,
    n2763_lo
  );


  not

  (
    n2763_lo_n,
    n2763_lo
  );


  buf

  (
    n2766_lo_p,
    n2766_lo
  );


  not

  (
    n2766_lo_n,
    n2766_lo
  );


  buf

  (
    n2769_lo_p,
    n2769_lo
  );


  not

  (
    n2769_lo_n,
    n2769_lo
  );


  buf

  (
    n2772_lo_p,
    n2772_lo
  );


  not

  (
    n2772_lo_n,
    n2772_lo
  );


  buf

  (
    n2775_lo_p,
    n2775_lo
  );


  not

  (
    n2775_lo_n,
    n2775_lo
  );


  buf

  (
    n2778_lo_p,
    n2778_lo
  );


  not

  (
    n2778_lo_n,
    n2778_lo
  );


  buf

  (
    n2781_lo_p,
    n2781_lo
  );


  not

  (
    n2781_lo_n,
    n2781_lo
  );


  buf

  (
    n2784_lo_p,
    n2784_lo
  );


  not

  (
    n2784_lo_n,
    n2784_lo
  );


  buf

  (
    n2787_lo_p,
    n2787_lo
  );


  not

  (
    n2787_lo_n,
    n2787_lo
  );


  buf

  (
    n2790_lo_p,
    n2790_lo
  );


  not

  (
    n2790_lo_n,
    n2790_lo
  );


  buf

  (
    n2793_lo_p,
    n2793_lo
  );


  not

  (
    n2793_lo_n,
    n2793_lo
  );


  buf

  (
    n2796_lo_p,
    n2796_lo
  );


  not

  (
    n2796_lo_n,
    n2796_lo
  );


  buf

  (
    n2799_lo_p,
    n2799_lo
  );


  not

  (
    n2799_lo_n,
    n2799_lo
  );


  buf

  (
    n2802_lo_p,
    n2802_lo
  );


  not

  (
    n2802_lo_n,
    n2802_lo
  );


  buf

  (
    n2805_lo_p,
    n2805_lo
  );


  not

  (
    n2805_lo_n,
    n2805_lo
  );


  buf

  (
    n2808_lo_p,
    n2808_lo
  );


  not

  (
    n2808_lo_n,
    n2808_lo
  );


  buf

  (
    n2811_lo_p,
    n2811_lo
  );


  not

  (
    n2811_lo_n,
    n2811_lo
  );


  buf

  (
    n2814_lo_p,
    n2814_lo
  );


  not

  (
    n2814_lo_n,
    n2814_lo
  );


  buf

  (
    n2817_lo_p,
    n2817_lo
  );


  not

  (
    n2817_lo_n,
    n2817_lo
  );


  buf

  (
    n2820_lo_p,
    n2820_lo
  );


  not

  (
    n2820_lo_n,
    n2820_lo
  );


  buf

  (
    n2823_lo_p,
    n2823_lo
  );


  not

  (
    n2823_lo_n,
    n2823_lo
  );


  buf

  (
    n2826_lo_p,
    n2826_lo
  );


  not

  (
    n2826_lo_n,
    n2826_lo
  );


  buf

  (
    n2829_lo_p,
    n2829_lo
  );


  not

  (
    n2829_lo_n,
    n2829_lo
  );


  buf

  (
    n2832_lo_p,
    n2832_lo
  );


  not

  (
    n2832_lo_n,
    n2832_lo
  );


  buf

  (
    n2838_lo_p,
    n2838_lo
  );


  not

  (
    n2838_lo_n,
    n2838_lo
  );


  buf

  (
    n2841_lo_p,
    n2841_lo
  );


  not

  (
    n2841_lo_n,
    n2841_lo
  );


  buf

  (
    n2844_lo_p,
    n2844_lo
  );


  not

  (
    n2844_lo_n,
    n2844_lo
  );


  buf

  (
    n2847_lo_p,
    n2847_lo
  );


  not

  (
    n2847_lo_n,
    n2847_lo
  );


  buf

  (
    n2850_lo_p,
    n2850_lo
  );


  not

  (
    n2850_lo_n,
    n2850_lo
  );


  buf

  (
    n2853_lo_p,
    n2853_lo
  );


  not

  (
    n2853_lo_n,
    n2853_lo
  );


  buf

  (
    n2856_lo_p,
    n2856_lo
  );


  not

  (
    n2856_lo_n,
    n2856_lo
  );


  buf

  (
    n2862_lo_p,
    n2862_lo
  );


  not

  (
    n2862_lo_n,
    n2862_lo
  );


  buf

  (
    n2865_lo_p,
    n2865_lo
  );


  not

  (
    n2865_lo_n,
    n2865_lo
  );


  buf

  (
    n2868_lo_p,
    n2868_lo
  );


  not

  (
    n2868_lo_n,
    n2868_lo
  );


  buf

  (
    n2871_lo_p,
    n2871_lo
  );


  not

  (
    n2871_lo_n,
    n2871_lo
  );


  buf

  (
    n2874_lo_p,
    n2874_lo
  );


  not

  (
    n2874_lo_n,
    n2874_lo
  );


  buf

  (
    n2877_lo_p,
    n2877_lo
  );


  not

  (
    n2877_lo_n,
    n2877_lo
  );


  buf

  (
    n2880_lo_p,
    n2880_lo
  );


  not

  (
    n2880_lo_n,
    n2880_lo
  );


  buf

  (
    n2883_lo_p,
    n2883_lo
  );


  not

  (
    n2883_lo_n,
    n2883_lo
  );


  buf

  (
    n2886_lo_p,
    n2886_lo
  );


  not

  (
    n2886_lo_n,
    n2886_lo
  );


  buf

  (
    n2889_lo_p,
    n2889_lo
  );


  not

  (
    n2889_lo_n,
    n2889_lo
  );


  buf

  (
    n2892_lo_p,
    n2892_lo
  );


  not

  (
    n2892_lo_n,
    n2892_lo
  );


  buf

  (
    n2895_lo_p,
    n2895_lo
  );


  not

  (
    n2895_lo_n,
    n2895_lo
  );


  buf

  (
    n2898_lo_p,
    n2898_lo
  );


  not

  (
    n2898_lo_n,
    n2898_lo
  );


  buf

  (
    n2901_lo_p,
    n2901_lo
  );


  not

  (
    n2901_lo_n,
    n2901_lo
  );


  buf

  (
    n2904_lo_p,
    n2904_lo
  );


  not

  (
    n2904_lo_n,
    n2904_lo
  );


  buf

  (
    n2907_lo_p,
    n2907_lo
  );


  not

  (
    n2907_lo_n,
    n2907_lo
  );


  buf

  (
    n2910_lo_p,
    n2910_lo
  );


  not

  (
    n2910_lo_n,
    n2910_lo
  );


  buf

  (
    n2913_lo_p,
    n2913_lo
  );


  not

  (
    n2913_lo_n,
    n2913_lo
  );


  buf

  (
    n2916_lo_p,
    n2916_lo
  );


  not

  (
    n2916_lo_n,
    n2916_lo
  );


  buf

  (
    n2919_lo_p,
    n2919_lo
  );


  not

  (
    n2919_lo_n,
    n2919_lo
  );


  buf

  (
    n2922_lo_p,
    n2922_lo
  );


  not

  (
    n2922_lo_n,
    n2922_lo
  );


  buf

  (
    n2925_lo_p,
    n2925_lo
  );


  not

  (
    n2925_lo_n,
    n2925_lo
  );


  buf

  (
    n2928_lo_p,
    n2928_lo
  );


  not

  (
    n2928_lo_n,
    n2928_lo
  );


  buf

  (
    n2931_lo_p,
    n2931_lo
  );


  not

  (
    n2931_lo_n,
    n2931_lo
  );


  buf

  (
    n2934_lo_p,
    n2934_lo
  );


  not

  (
    n2934_lo_n,
    n2934_lo
  );


  buf

  (
    n2937_lo_p,
    n2937_lo
  );


  not

  (
    n2937_lo_n,
    n2937_lo
  );


  buf

  (
    n2940_lo_p,
    n2940_lo
  );


  not

  (
    n2940_lo_n,
    n2940_lo
  );


  buf

  (
    n2943_lo_p,
    n2943_lo
  );


  not

  (
    n2943_lo_n,
    n2943_lo
  );


  buf

  (
    n2946_lo_p,
    n2946_lo
  );


  not

  (
    n2946_lo_n,
    n2946_lo
  );


  buf

  (
    n2949_lo_p,
    n2949_lo
  );


  not

  (
    n2949_lo_n,
    n2949_lo
  );


  buf

  (
    n2952_lo_p,
    n2952_lo
  );


  not

  (
    n2952_lo_n,
    n2952_lo
  );


  buf

  (
    n2955_lo_p,
    n2955_lo
  );


  not

  (
    n2955_lo_n,
    n2955_lo
  );


  buf

  (
    n2958_lo_p,
    n2958_lo
  );


  not

  (
    n2958_lo_n,
    n2958_lo
  );


  buf

  (
    n2961_lo_p,
    n2961_lo
  );


  not

  (
    n2961_lo_n,
    n2961_lo
  );


  buf

  (
    n2964_lo_p,
    n2964_lo
  );


  not

  (
    n2964_lo_n,
    n2964_lo
  );


  buf

  (
    n2967_lo_p,
    n2967_lo
  );


  not

  (
    n2967_lo_n,
    n2967_lo
  );


  buf

  (
    n2970_lo_p,
    n2970_lo
  );


  not

  (
    n2970_lo_n,
    n2970_lo
  );


  buf

  (
    n2973_lo_p,
    n2973_lo
  );


  not

  (
    n2973_lo_n,
    n2973_lo
  );


  buf

  (
    n2976_lo_p,
    n2976_lo
  );


  not

  (
    n2976_lo_n,
    n2976_lo
  );


  buf

  (
    n2979_lo_p,
    n2979_lo
  );


  not

  (
    n2979_lo_n,
    n2979_lo
  );


  buf

  (
    n2982_lo_p,
    n2982_lo
  );


  not

  (
    n2982_lo_n,
    n2982_lo
  );


  buf

  (
    n2985_lo_p,
    n2985_lo
  );


  not

  (
    n2985_lo_n,
    n2985_lo
  );


  buf

  (
    n2988_lo_p,
    n2988_lo
  );


  not

  (
    n2988_lo_n,
    n2988_lo
  );


  buf

  (
    n2991_lo_p,
    n2991_lo
  );


  not

  (
    n2991_lo_n,
    n2991_lo
  );


  buf

  (
    n2994_lo_p,
    n2994_lo
  );


  not

  (
    n2994_lo_n,
    n2994_lo
  );


  buf

  (
    n2997_lo_p,
    n2997_lo
  );


  not

  (
    n2997_lo_n,
    n2997_lo
  );


  buf

  (
    n3000_lo_p,
    n3000_lo
  );


  not

  (
    n3000_lo_n,
    n3000_lo
  );


  buf

  (
    n3003_lo_p,
    n3003_lo
  );


  not

  (
    n3003_lo_n,
    n3003_lo
  );


  buf

  (
    n3006_lo_p,
    n3006_lo
  );


  not

  (
    n3006_lo_n,
    n3006_lo
  );


  buf

  (
    n3009_lo_p,
    n3009_lo
  );


  not

  (
    n3009_lo_n,
    n3009_lo
  );


  buf

  (
    n3012_lo_p,
    n3012_lo
  );


  not

  (
    n3012_lo_n,
    n3012_lo
  );


  buf

  (
    n3015_lo_p,
    n3015_lo
  );


  not

  (
    n3015_lo_n,
    n3015_lo
  );


  buf

  (
    n3018_lo_p,
    n3018_lo
  );


  not

  (
    n3018_lo_n,
    n3018_lo
  );


  buf

  (
    n3021_lo_p,
    n3021_lo
  );


  not

  (
    n3021_lo_n,
    n3021_lo
  );


  buf

  (
    n3024_lo_p,
    n3024_lo
  );


  not

  (
    n3024_lo_n,
    n3024_lo
  );


  buf

  (
    n3027_lo_p,
    n3027_lo
  );


  not

  (
    n3027_lo_n,
    n3027_lo
  );


  buf

  (
    n3030_lo_p,
    n3030_lo
  );


  not

  (
    n3030_lo_n,
    n3030_lo
  );


  buf

  (
    n3033_lo_p,
    n3033_lo
  );


  not

  (
    n3033_lo_n,
    n3033_lo
  );


  buf

  (
    n3036_lo_p,
    n3036_lo
  );


  not

  (
    n3036_lo_n,
    n3036_lo
  );


  buf

  (
    n3039_lo_p,
    n3039_lo
  );


  not

  (
    n3039_lo_n,
    n3039_lo
  );


  buf

  (
    n3042_lo_p,
    n3042_lo
  );


  not

  (
    n3042_lo_n,
    n3042_lo
  );


  buf

  (
    n3045_lo_p,
    n3045_lo
  );


  not

  (
    n3045_lo_n,
    n3045_lo
  );


  buf

  (
    n3048_lo_p,
    n3048_lo
  );


  not

  (
    n3048_lo_n,
    n3048_lo
  );


  buf

  (
    n3051_lo_p,
    n3051_lo
  );


  not

  (
    n3051_lo_n,
    n3051_lo
  );


  buf

  (
    n3054_lo_p,
    n3054_lo
  );


  not

  (
    n3054_lo_n,
    n3054_lo
  );


  buf

  (
    n3057_lo_p,
    n3057_lo
  );


  not

  (
    n3057_lo_n,
    n3057_lo
  );


  buf

  (
    n3060_lo_p,
    n3060_lo
  );


  not

  (
    n3060_lo_n,
    n3060_lo
  );


  buf

  (
    n3063_lo_p,
    n3063_lo
  );


  not

  (
    n3063_lo_n,
    n3063_lo
  );


  buf

  (
    n3066_lo_p,
    n3066_lo
  );


  not

  (
    n3066_lo_n,
    n3066_lo
  );


  buf

  (
    n3069_lo_p,
    n3069_lo
  );


  not

  (
    n3069_lo_n,
    n3069_lo
  );


  buf

  (
    n3072_lo_p,
    n3072_lo
  );


  not

  (
    n3072_lo_n,
    n3072_lo
  );


  buf

  (
    n3075_lo_p,
    n3075_lo
  );


  not

  (
    n3075_lo_n,
    n3075_lo
  );


  buf

  (
    n3078_lo_p,
    n3078_lo
  );


  not

  (
    n3078_lo_n,
    n3078_lo
  );


  buf

  (
    n3081_lo_p,
    n3081_lo
  );


  not

  (
    n3081_lo_n,
    n3081_lo
  );


  buf

  (
    n3084_lo_p,
    n3084_lo
  );


  not

  (
    n3084_lo_n,
    n3084_lo
  );


  buf

  (
    n3087_lo_p,
    n3087_lo
  );


  not

  (
    n3087_lo_n,
    n3087_lo
  );


  buf

  (
    n3090_lo_p,
    n3090_lo
  );


  not

  (
    n3090_lo_n,
    n3090_lo
  );


  buf

  (
    n3093_lo_p,
    n3093_lo
  );


  not

  (
    n3093_lo_n,
    n3093_lo
  );


  buf

  (
    n3096_lo_p,
    n3096_lo
  );


  not

  (
    n3096_lo_n,
    n3096_lo
  );


  buf

  (
    n3099_lo_p,
    n3099_lo
  );


  not

  (
    n3099_lo_n,
    n3099_lo
  );


  buf

  (
    n3102_lo_p,
    n3102_lo
  );


  not

  (
    n3102_lo_n,
    n3102_lo
  );


  buf

  (
    n3105_lo_p,
    n3105_lo
  );


  not

  (
    n3105_lo_n,
    n3105_lo
  );


  buf

  (
    n3108_lo_p,
    n3108_lo
  );


  not

  (
    n3108_lo_n,
    n3108_lo
  );


  buf

  (
    n3111_lo_p,
    n3111_lo
  );


  not

  (
    n3111_lo_n,
    n3111_lo
  );


  buf

  (
    n3114_lo_p,
    n3114_lo
  );


  not

  (
    n3114_lo_n,
    n3114_lo
  );


  buf

  (
    n3117_lo_p,
    n3117_lo
  );


  not

  (
    n3117_lo_n,
    n3117_lo
  );


  buf

  (
    n3120_lo_p,
    n3120_lo
  );


  not

  (
    n3120_lo_n,
    n3120_lo
  );


  buf

  (
    n3126_lo_p,
    n3126_lo
  );


  not

  (
    n3126_lo_n,
    n3126_lo
  );


  buf

  (
    n3129_lo_p,
    n3129_lo
  );


  not

  (
    n3129_lo_n,
    n3129_lo
  );


  buf

  (
    n3132_lo_p,
    n3132_lo
  );


  not

  (
    n3132_lo_n,
    n3132_lo
  );


  buf

  (
    n3138_lo_p,
    n3138_lo
  );


  not

  (
    n3138_lo_n,
    n3138_lo
  );


  buf

  (
    n3141_lo_p,
    n3141_lo
  );


  not

  (
    n3141_lo_n,
    n3141_lo
  );


  buf

  (
    n3144_lo_p,
    n3144_lo
  );


  not

  (
    n3144_lo_n,
    n3144_lo
  );


  buf

  (
    n3147_lo_p,
    n3147_lo
  );


  not

  (
    n3147_lo_n,
    n3147_lo
  );


  buf

  (
    n3150_lo_p,
    n3150_lo
  );


  not

  (
    n3150_lo_n,
    n3150_lo
  );


  buf

  (
    n3153_lo_p,
    n3153_lo
  );


  not

  (
    n3153_lo_n,
    n3153_lo
  );


  buf

  (
    n3156_lo_p,
    n3156_lo
  );


  not

  (
    n3156_lo_n,
    n3156_lo
  );


  buf

  (
    n3162_lo_p,
    n3162_lo
  );


  not

  (
    n3162_lo_n,
    n3162_lo
  );


  buf

  (
    n3165_lo_p,
    n3165_lo
  );


  not

  (
    n3165_lo_n,
    n3165_lo
  );


  buf

  (
    n3168_lo_p,
    n3168_lo
  );


  not

  (
    n3168_lo_n,
    n3168_lo
  );


  buf

  (
    n3174_lo_p,
    n3174_lo
  );


  not

  (
    n3174_lo_n,
    n3174_lo
  );


  buf

  (
    n3177_lo_p,
    n3177_lo
  );


  not

  (
    n3177_lo_n,
    n3177_lo
  );


  buf

  (
    n3180_lo_p,
    n3180_lo
  );


  not

  (
    n3180_lo_n,
    n3180_lo
  );


  buf

  (
    n3186_lo_p,
    n3186_lo
  );


  not

  (
    n3186_lo_n,
    n3186_lo
  );


  buf

  (
    n3189_lo_p,
    n3189_lo
  );


  not

  (
    n3189_lo_n,
    n3189_lo
  );


  buf

  (
    n3192_lo_p,
    n3192_lo
  );


  not

  (
    n3192_lo_n,
    n3192_lo
  );


  buf

  (
    n3195_lo_p,
    n3195_lo
  );


  not

  (
    n3195_lo_n,
    n3195_lo
  );


  buf

  (
    n3198_lo_p,
    n3198_lo
  );


  not

  (
    n3198_lo_n,
    n3198_lo
  );


  buf

  (
    n3201_lo_p,
    n3201_lo
  );


  not

  (
    n3201_lo_n,
    n3201_lo
  );


  buf

  (
    n3204_lo_p,
    n3204_lo
  );


  not

  (
    n3204_lo_n,
    n3204_lo
  );


  buf

  (
    n3210_lo_p,
    n3210_lo
  );


  not

  (
    n3210_lo_n,
    n3210_lo
  );


  buf

  (
    n3213_lo_p,
    n3213_lo
  );


  not

  (
    n3213_lo_n,
    n3213_lo
  );


  buf

  (
    n3216_lo_p,
    n3216_lo
  );


  not

  (
    n3216_lo_n,
    n3216_lo
  );


  buf

  (
    n3219_lo_p,
    n3219_lo
  );


  not

  (
    n3219_lo_n,
    n3219_lo
  );


  buf

  (
    n3222_lo_p,
    n3222_lo
  );


  not

  (
    n3222_lo_n,
    n3222_lo
  );


  buf

  (
    n3225_lo_p,
    n3225_lo
  );


  not

  (
    n3225_lo_n,
    n3225_lo
  );


  buf

  (
    n3228_lo_p,
    n3228_lo
  );


  not

  (
    n3228_lo_n,
    n3228_lo
  );


  buf

  (
    n3234_lo_p,
    n3234_lo
  );


  not

  (
    n3234_lo_n,
    n3234_lo
  );


  buf

  (
    n3237_lo_p,
    n3237_lo
  );


  not

  (
    n3237_lo_n,
    n3237_lo
  );


  buf

  (
    n3240_lo_p,
    n3240_lo
  );


  not

  (
    n3240_lo_n,
    n3240_lo
  );


  buf

  (
    n3243_lo_p,
    n3243_lo
  );


  not

  (
    n3243_lo_n,
    n3243_lo
  );


  buf

  (
    n3246_lo_p,
    n3246_lo
  );


  not

  (
    n3246_lo_n,
    n3246_lo
  );


  buf

  (
    n3249_lo_p,
    n3249_lo
  );


  not

  (
    n3249_lo_n,
    n3249_lo
  );


  buf

  (
    n3252_lo_p,
    n3252_lo
  );


  not

  (
    n3252_lo_n,
    n3252_lo
  );


  buf

  (
    n3255_lo_p,
    n3255_lo
  );


  not

  (
    n3255_lo_n,
    n3255_lo
  );


  buf

  (
    n3258_lo_p,
    n3258_lo
  );


  not

  (
    n3258_lo_n,
    n3258_lo
  );


  buf

  (
    n3261_lo_p,
    n3261_lo
  );


  not

  (
    n3261_lo_n,
    n3261_lo
  );


  buf

  (
    n3264_lo_p,
    n3264_lo
  );


  not

  (
    n3264_lo_n,
    n3264_lo
  );


  buf

  (
    n3267_lo_p,
    n3267_lo
  );


  not

  (
    n3267_lo_n,
    n3267_lo
  );


  buf

  (
    n3270_lo_p,
    n3270_lo
  );


  not

  (
    n3270_lo_n,
    n3270_lo
  );


  buf

  (
    n3273_lo_p,
    n3273_lo
  );


  not

  (
    n3273_lo_n,
    n3273_lo
  );


  buf

  (
    n3276_lo_p,
    n3276_lo
  );


  not

  (
    n3276_lo_n,
    n3276_lo
  );


  buf

  (
    n3279_lo_p,
    n3279_lo
  );


  not

  (
    n3279_lo_n,
    n3279_lo
  );


  buf

  (
    n3282_lo_p,
    n3282_lo
  );


  not

  (
    n3282_lo_n,
    n3282_lo
  );


  buf

  (
    n3285_lo_p,
    n3285_lo
  );


  not

  (
    n3285_lo_n,
    n3285_lo
  );


  buf

  (
    n3288_lo_p,
    n3288_lo
  );


  not

  (
    n3288_lo_n,
    n3288_lo
  );


  buf

  (
    n3294_lo_p,
    n3294_lo
  );


  not

  (
    n3294_lo_n,
    n3294_lo
  );


  buf

  (
    n3297_lo_p,
    n3297_lo
  );


  not

  (
    n3297_lo_n,
    n3297_lo
  );


  buf

  (
    n3300_lo_p,
    n3300_lo
  );


  not

  (
    n3300_lo_n,
    n3300_lo
  );


  buf

  (
    n3306_lo_p,
    n3306_lo
  );


  not

  (
    n3306_lo_n,
    n3306_lo
  );


  buf

  (
    n3309_lo_p,
    n3309_lo
  );


  not

  (
    n3309_lo_n,
    n3309_lo
  );


  buf

  (
    n3312_lo_p,
    n3312_lo
  );


  not

  (
    n3312_lo_n,
    n3312_lo
  );


  buf

  (
    n3318_lo_p,
    n3318_lo
  );


  not

  (
    n3318_lo_n,
    n3318_lo
  );


  buf

  (
    n3321_lo_p,
    n3321_lo
  );


  not

  (
    n3321_lo_n,
    n3321_lo
  );


  buf

  (
    n3324_lo_p,
    n3324_lo
  );


  not

  (
    n3324_lo_n,
    n3324_lo
  );


  buf

  (
    n3330_lo_p,
    n3330_lo
  );


  not

  (
    n3330_lo_n,
    n3330_lo
  );


  buf

  (
    n3333_lo_p,
    n3333_lo
  );


  not

  (
    n3333_lo_n,
    n3333_lo
  );


  buf

  (
    n3336_lo_p,
    n3336_lo
  );


  not

  (
    n3336_lo_n,
    n3336_lo
  );


  buf

  (
    n3339_lo_p,
    n3339_lo
  );


  not

  (
    n3339_lo_n,
    n3339_lo
  );


  buf

  (
    n3342_lo_p,
    n3342_lo
  );


  not

  (
    n3342_lo_n,
    n3342_lo
  );


  buf

  (
    n3345_lo_p,
    n3345_lo
  );


  not

  (
    n3345_lo_n,
    n3345_lo
  );


  buf

  (
    n3348_lo_p,
    n3348_lo
  );


  not

  (
    n3348_lo_n,
    n3348_lo
  );


  buf

  (
    n3351_lo_p,
    n3351_lo
  );


  not

  (
    n3351_lo_n,
    n3351_lo
  );


  buf

  (
    n3354_lo_p,
    n3354_lo
  );


  not

  (
    n3354_lo_n,
    n3354_lo
  );


  buf

  (
    n3357_lo_p,
    n3357_lo
  );


  not

  (
    n3357_lo_n,
    n3357_lo
  );


  buf

  (
    n3360_lo_p,
    n3360_lo
  );


  not

  (
    n3360_lo_n,
    n3360_lo
  );


  buf

  (
    n3363_lo_p,
    n3363_lo
  );


  not

  (
    n3363_lo_n,
    n3363_lo
  );


  buf

  (
    n3366_lo_p,
    n3366_lo
  );


  not

  (
    n3366_lo_n,
    n3366_lo
  );


  buf

  (
    n3369_lo_p,
    n3369_lo
  );


  not

  (
    n3369_lo_n,
    n3369_lo
  );


  buf

  (
    n3372_lo_p,
    n3372_lo
  );


  not

  (
    n3372_lo_n,
    n3372_lo
  );


  buf

  (
    n3375_lo_p,
    n3375_lo
  );


  not

  (
    n3375_lo_n,
    n3375_lo
  );


  buf

  (
    n3378_lo_p,
    n3378_lo
  );


  not

  (
    n3378_lo_n,
    n3378_lo
  );


  buf

  (
    n3381_lo_p,
    n3381_lo
  );


  not

  (
    n3381_lo_n,
    n3381_lo
  );


  buf

  (
    n3384_lo_p,
    n3384_lo
  );


  not

  (
    n3384_lo_n,
    n3384_lo
  );


  buf

  (
    n3387_lo_p,
    n3387_lo
  );


  not

  (
    n3387_lo_n,
    n3387_lo
  );


  buf

  (
    n3390_lo_p,
    n3390_lo
  );


  not

  (
    n3390_lo_n,
    n3390_lo
  );


  buf

  (
    n3393_lo_p,
    n3393_lo
  );


  not

  (
    n3393_lo_n,
    n3393_lo
  );


  buf

  (
    n3396_lo_p,
    n3396_lo
  );


  not

  (
    n3396_lo_n,
    n3396_lo
  );


  buf

  (
    n3399_lo_p,
    n3399_lo
  );


  not

  (
    n3399_lo_n,
    n3399_lo
  );


  buf

  (
    n3402_lo_p,
    n3402_lo
  );


  not

  (
    n3402_lo_n,
    n3402_lo
  );


  buf

  (
    n3405_lo_p,
    n3405_lo
  );


  not

  (
    n3405_lo_n,
    n3405_lo
  );


  buf

  (
    n3408_lo_p,
    n3408_lo
  );


  not

  (
    n3408_lo_n,
    n3408_lo
  );


  buf

  (
    n3411_lo_p,
    n3411_lo
  );


  not

  (
    n3411_lo_n,
    n3411_lo
  );


  buf

  (
    n3414_lo_p,
    n3414_lo
  );


  not

  (
    n3414_lo_n,
    n3414_lo
  );


  buf

  (
    n3417_lo_p,
    n3417_lo
  );


  not

  (
    n3417_lo_n,
    n3417_lo
  );


  buf

  (
    n3420_lo_p,
    n3420_lo
  );


  not

  (
    n3420_lo_n,
    n3420_lo
  );


  buf

  (
    n3423_lo_p,
    n3423_lo
  );


  not

  (
    n3423_lo_n,
    n3423_lo
  );


  buf

  (
    n3426_lo_p,
    n3426_lo
  );


  not

  (
    n3426_lo_n,
    n3426_lo
  );


  buf

  (
    n3429_lo_p,
    n3429_lo
  );


  not

  (
    n3429_lo_n,
    n3429_lo
  );


  buf

  (
    n3432_lo_p,
    n3432_lo
  );


  not

  (
    n3432_lo_n,
    n3432_lo
  );


  buf

  (
    n3435_lo_p,
    n3435_lo
  );


  not

  (
    n3435_lo_n,
    n3435_lo
  );


  buf

  (
    n3438_lo_p,
    n3438_lo
  );


  not

  (
    n3438_lo_n,
    n3438_lo
  );


  buf

  (
    n3441_lo_p,
    n3441_lo
  );


  not

  (
    n3441_lo_n,
    n3441_lo
  );


  buf

  (
    n3444_lo_p,
    n3444_lo
  );


  not

  (
    n3444_lo_n,
    n3444_lo
  );


  buf

  (
    n3447_lo_p,
    n3447_lo
  );


  not

  (
    n3447_lo_n,
    n3447_lo
  );


  buf

  (
    n3450_lo_p,
    n3450_lo
  );


  not

  (
    n3450_lo_n,
    n3450_lo
  );


  buf

  (
    n3453_lo_p,
    n3453_lo
  );


  not

  (
    n3453_lo_n,
    n3453_lo
  );


  buf

  (
    n3456_lo_p,
    n3456_lo
  );


  not

  (
    n3456_lo_n,
    n3456_lo
  );


  buf

  (
    n3459_lo_p,
    n3459_lo
  );


  not

  (
    n3459_lo_n,
    n3459_lo
  );


  buf

  (
    n3462_lo_p,
    n3462_lo
  );


  not

  (
    n3462_lo_n,
    n3462_lo
  );


  buf

  (
    n3465_lo_p,
    n3465_lo
  );


  not

  (
    n3465_lo_n,
    n3465_lo
  );


  buf

  (
    n3468_lo_p,
    n3468_lo
  );


  not

  (
    n3468_lo_n,
    n3468_lo
  );


  buf

  (
    n3471_lo_p,
    n3471_lo
  );


  not

  (
    n3471_lo_n,
    n3471_lo
  );


  buf

  (
    n3474_lo_p,
    n3474_lo
  );


  not

  (
    n3474_lo_n,
    n3474_lo
  );


  buf

  (
    n3477_lo_p,
    n3477_lo
  );


  not

  (
    n3477_lo_n,
    n3477_lo
  );


  buf

  (
    n3480_lo_p,
    n3480_lo
  );


  not

  (
    n3480_lo_n,
    n3480_lo
  );


  buf

  (
    n3483_lo_p,
    n3483_lo
  );


  not

  (
    n3483_lo_n,
    n3483_lo
  );


  buf

  (
    n3486_lo_p,
    n3486_lo
  );


  not

  (
    n3486_lo_n,
    n3486_lo
  );


  buf

  (
    n3489_lo_p,
    n3489_lo
  );


  not

  (
    n3489_lo_n,
    n3489_lo
  );


  buf

  (
    n3492_lo_p,
    n3492_lo
  );


  not

  (
    n3492_lo_n,
    n3492_lo
  );


  buf

  (
    n3495_lo_p,
    n3495_lo
  );


  not

  (
    n3495_lo_n,
    n3495_lo
  );


  buf

  (
    n3498_lo_p,
    n3498_lo
  );


  not

  (
    n3498_lo_n,
    n3498_lo
  );


  buf

  (
    n3501_lo_p,
    n3501_lo
  );


  not

  (
    n3501_lo_n,
    n3501_lo
  );


  buf

  (
    n3504_lo_p,
    n3504_lo
  );


  not

  (
    n3504_lo_n,
    n3504_lo
  );


  buf

  (
    n3507_lo_p,
    n3507_lo
  );


  not

  (
    n3507_lo_n,
    n3507_lo
  );


  buf

  (
    n3510_lo_p,
    n3510_lo
  );


  not

  (
    n3510_lo_n,
    n3510_lo
  );


  buf

  (
    n3513_lo_p,
    n3513_lo
  );


  not

  (
    n3513_lo_n,
    n3513_lo
  );


  buf

  (
    n3516_lo_p,
    n3516_lo
  );


  not

  (
    n3516_lo_n,
    n3516_lo
  );


  buf

  (
    n3519_lo_p,
    n3519_lo
  );


  not

  (
    n3519_lo_n,
    n3519_lo
  );


  buf

  (
    n3522_lo_p,
    n3522_lo
  );


  not

  (
    n3522_lo_n,
    n3522_lo
  );


  buf

  (
    n3525_lo_p,
    n3525_lo
  );


  not

  (
    n3525_lo_n,
    n3525_lo
  );


  buf

  (
    n3528_lo_p,
    n3528_lo
  );


  not

  (
    n3528_lo_n,
    n3528_lo
  );


  buf

  (
    n3531_lo_p,
    n3531_lo
  );


  not

  (
    n3531_lo_n,
    n3531_lo
  );


  buf

  (
    n3534_lo_p,
    n3534_lo
  );


  not

  (
    n3534_lo_n,
    n3534_lo
  );


  buf

  (
    n3537_lo_p,
    n3537_lo
  );


  not

  (
    n3537_lo_n,
    n3537_lo
  );


  buf

  (
    n3540_lo_p,
    n3540_lo
  );


  not

  (
    n3540_lo_n,
    n3540_lo
  );


  buf

  (
    n3543_lo_p,
    n3543_lo
  );


  not

  (
    n3543_lo_n,
    n3543_lo
  );


  buf

  (
    n3546_lo_p,
    n3546_lo
  );


  not

  (
    n3546_lo_n,
    n3546_lo
  );


  buf

  (
    n3549_lo_p,
    n3549_lo
  );


  not

  (
    n3549_lo_n,
    n3549_lo
  );


  buf

  (
    n3552_lo_p,
    n3552_lo
  );


  not

  (
    n3552_lo_n,
    n3552_lo
  );


  buf

  (
    n3555_lo_p,
    n3555_lo
  );


  not

  (
    n3555_lo_n,
    n3555_lo
  );


  buf

  (
    n3558_lo_p,
    n3558_lo
  );


  not

  (
    n3558_lo_n,
    n3558_lo
  );


  buf

  (
    n3561_lo_p,
    n3561_lo
  );


  not

  (
    n3561_lo_n,
    n3561_lo
  );


  buf

  (
    n3564_lo_p,
    n3564_lo
  );


  not

  (
    n3564_lo_n,
    n3564_lo
  );


  buf

  (
    n3567_lo_p,
    n3567_lo
  );


  not

  (
    n3567_lo_n,
    n3567_lo
  );


  buf

  (
    n3570_lo_p,
    n3570_lo
  );


  not

  (
    n3570_lo_n,
    n3570_lo
  );


  buf

  (
    n3573_lo_p,
    n3573_lo
  );


  not

  (
    n3573_lo_n,
    n3573_lo
  );


  buf

  (
    n3576_lo_p,
    n3576_lo
  );


  not

  (
    n3576_lo_n,
    n3576_lo
  );


  buf

  (
    n3579_lo_p,
    n3579_lo
  );


  not

  (
    n3579_lo_n,
    n3579_lo
  );


  buf

  (
    n3582_lo_p,
    n3582_lo
  );


  not

  (
    n3582_lo_n,
    n3582_lo
  );


  buf

  (
    n3585_lo_p,
    n3585_lo
  );


  not

  (
    n3585_lo_n,
    n3585_lo
  );


  buf

  (
    n3588_lo_p,
    n3588_lo
  );


  not

  (
    n3588_lo_n,
    n3588_lo
  );


  buf

  (
    n3591_lo_p,
    n3591_lo
  );


  not

  (
    n3591_lo_n,
    n3591_lo
  );


  buf

  (
    n3594_lo_p,
    n3594_lo
  );


  not

  (
    n3594_lo_n,
    n3594_lo
  );


  buf

  (
    n3597_lo_p,
    n3597_lo
  );


  not

  (
    n3597_lo_n,
    n3597_lo
  );


  buf

  (
    n3600_lo_p,
    n3600_lo
  );


  not

  (
    n3600_lo_n,
    n3600_lo
  );


  buf

  (
    n3603_lo_p,
    n3603_lo
  );


  not

  (
    n3603_lo_n,
    n3603_lo
  );


  buf

  (
    n3606_lo_p,
    n3606_lo
  );


  not

  (
    n3606_lo_n,
    n3606_lo
  );


  buf

  (
    n3609_lo_p,
    n3609_lo
  );


  not

  (
    n3609_lo_n,
    n3609_lo
  );


  buf

  (
    n3612_lo_p,
    n3612_lo
  );


  not

  (
    n3612_lo_n,
    n3612_lo
  );


  buf

  (
    n3615_lo_p,
    n3615_lo
  );


  not

  (
    n3615_lo_n,
    n3615_lo
  );


  buf

  (
    n3618_lo_p,
    n3618_lo
  );


  not

  (
    n3618_lo_n,
    n3618_lo
  );


  buf

  (
    n3621_lo_p,
    n3621_lo
  );


  not

  (
    n3621_lo_n,
    n3621_lo
  );


  buf

  (
    n3624_lo_p,
    n3624_lo
  );


  not

  (
    n3624_lo_n,
    n3624_lo
  );


  buf

  (
    n3627_lo_p,
    n3627_lo
  );


  not

  (
    n3627_lo_n,
    n3627_lo
  );


  buf

  (
    n3630_lo_p,
    n3630_lo
  );


  not

  (
    n3630_lo_n,
    n3630_lo
  );


  buf

  (
    n3633_lo_p,
    n3633_lo
  );


  not

  (
    n3633_lo_n,
    n3633_lo
  );


  buf

  (
    n3636_lo_p,
    n3636_lo
  );


  not

  (
    n3636_lo_n,
    n3636_lo
  );


  buf

  (
    n3639_lo_p,
    n3639_lo
  );


  not

  (
    n3639_lo_n,
    n3639_lo
  );


  buf

  (
    n3642_lo_p,
    n3642_lo
  );


  not

  (
    n3642_lo_n,
    n3642_lo
  );


  buf

  (
    n3645_lo_p,
    n3645_lo
  );


  not

  (
    n3645_lo_n,
    n3645_lo
  );


  buf

  (
    n3648_lo_p,
    n3648_lo
  );


  not

  (
    n3648_lo_n,
    n3648_lo
  );


  buf

  (
    n3651_lo_p,
    n3651_lo
  );


  not

  (
    n3651_lo_n,
    n3651_lo
  );


  buf

  (
    n3654_lo_p,
    n3654_lo
  );


  not

  (
    n3654_lo_n,
    n3654_lo
  );


  buf

  (
    n3666_lo_p,
    n3666_lo
  );


  not

  (
    n3666_lo_n,
    n3666_lo
  );


  buf

  (
    n3750_lo_p,
    n3750_lo
  );


  not

  (
    n3750_lo_n,
    n3750_lo
  );


  buf

  (
    n3762_lo_p,
    n3762_lo
  );


  not

  (
    n3762_lo_n,
    n3762_lo
  );


  buf

  (
    n3774_lo_p,
    n3774_lo
  );


  not

  (
    n3774_lo_n,
    n3774_lo
  );


  buf

  (
    n3786_lo_p,
    n3786_lo
  );


  not

  (
    n3786_lo_n,
    n3786_lo
  );


  buf

  (
    n3789_lo_p,
    n3789_lo
  );


  not

  (
    n3789_lo_n,
    n3789_lo
  );


  buf

  (
    n3792_lo_p,
    n3792_lo
  );


  not

  (
    n3792_lo_n,
    n3792_lo
  );


  buf

  (
    n3795_lo_p,
    n3795_lo
  );


  not

  (
    n3795_lo_n,
    n3795_lo
  );


  buf

  (
    n3798_lo_p,
    n3798_lo
  );


  not

  (
    n3798_lo_n,
    n3798_lo
  );


  buf

  (
    n3810_lo_p,
    n3810_lo
  );


  not

  (
    n3810_lo_n,
    n3810_lo
  );


  buf

  (
    n3822_lo_p,
    n3822_lo
  );


  not

  (
    n3822_lo_n,
    n3822_lo
  );


  buf

  (
    n3834_lo_p,
    n3834_lo
  );


  not

  (
    n3834_lo_n,
    n3834_lo
  );


  buf

  (
    n3846_lo_p,
    n3846_lo
  );


  not

  (
    n3846_lo_n,
    n3846_lo
  );


  buf

  (
    n3930_lo_p,
    n3930_lo
  );


  not

  (
    n3930_lo_n,
    n3930_lo
  );


  buf

  (
    n3933_lo_p,
    n3933_lo
  );


  not

  (
    n3933_lo_n,
    n3933_lo
  );


  buf

  (
    n3936_lo_p,
    n3936_lo
  );


  not

  (
    n3936_lo_n,
    n3936_lo
  );


  buf

  (
    n3942_lo_p,
    n3942_lo
  );


  not

  (
    n3942_lo_n,
    n3942_lo
  );


  buf

  (
    n3945_lo_p,
    n3945_lo
  );


  not

  (
    n3945_lo_n,
    n3945_lo
  );


  buf

  (
    n3948_lo_p,
    n3948_lo
  );


  not

  (
    n3948_lo_n,
    n3948_lo
  );


  buf

  (
    n3954_lo_p,
    n3954_lo
  );


  not

  (
    n3954_lo_n,
    n3954_lo
  );


  buf

  (
    n3957_lo_p,
    n3957_lo
  );


  not

  (
    n3957_lo_n,
    n3957_lo
  );


  buf

  (
    n3963_lo_p,
    n3963_lo
  );


  not

  (
    n3963_lo_n,
    n3963_lo
  );


  buf

  (
    n3966_lo_p,
    n3966_lo
  );


  not

  (
    n3966_lo_n,
    n3966_lo
  );


  buf

  (
    n3969_lo_p,
    n3969_lo
  );


  not

  (
    n3969_lo_n,
    n3969_lo
  );


  buf

  (
    n3975_lo_p,
    n3975_lo
  );


  not

  (
    n3975_lo_n,
    n3975_lo
  );


  buf

  (
    n3978_lo_p,
    n3978_lo
  );


  not

  (
    n3978_lo_n,
    n3978_lo
  );


  buf

  (
    n3990_lo_p,
    n3990_lo
  );


  not

  (
    n3990_lo_n,
    n3990_lo
  );


  buf

  (
    n4050_lo_p,
    n4050_lo
  );


  not

  (
    n4050_lo_n,
    n4050_lo
  );


  buf

  (
    n4062_lo_p,
    n4062_lo
  );


  not

  (
    n4062_lo_n,
    n4062_lo
  );


  buf

  (
    n4098_lo_p,
    n4098_lo
  );


  not

  (
    n4098_lo_n,
    n4098_lo
  );


  buf

  (
    n4107_lo_p,
    n4107_lo
  );


  not

  (
    n4107_lo_n,
    n4107_lo
  );


  buf

  (
    n4110_lo_p,
    n4110_lo
  );


  not

  (
    n4110_lo_n,
    n4110_lo
  );


  buf

  (
    n4122_lo_p,
    n4122_lo
  );


  not

  (
    n4122_lo_n,
    n4122_lo
  );


  buf

  (
    n4131_lo_p,
    n4131_lo
  );


  not

  (
    n4131_lo_n,
    n4131_lo
  );


  buf

  (
    n4155_lo_p,
    n4155_lo
  );


  not

  (
    n4155_lo_n,
    n4155_lo
  );


  buf

  (
    n4158_lo_p,
    n4158_lo
  );


  not

  (
    n4158_lo_n,
    n4158_lo
  );


  buf

  (
    n4170_lo_p,
    n4170_lo
  );


  not

  (
    n4170_lo_n,
    n4170_lo
  );


  buf

  (
    n4179_lo_p,
    n4179_lo
  );


  not

  (
    n4179_lo_n,
    n4179_lo
  );


  buf

  (
    n4182_lo_p,
    n4182_lo
  );


  not

  (
    n4182_lo_n,
    n4182_lo
  );


  buf

  (
    n4185_lo_p,
    n4185_lo
  );


  not

  (
    n4185_lo_n,
    n4185_lo
  );


  buf

  (
    n4188_lo_p,
    n4188_lo
  );


  not

  (
    n4188_lo_n,
    n4188_lo
  );


  buf

  (
    n4194_lo_p,
    n4194_lo
  );


  not

  (
    n4194_lo_n,
    n4194_lo
  );


  buf

  (
    n4197_lo_p,
    n4197_lo
  );


  not

  (
    n4197_lo_n,
    n4197_lo
  );


  buf

  (
    n4200_lo_p,
    n4200_lo
  );


  not

  (
    n4200_lo_n,
    n4200_lo
  );


  buf

  (
    n4206_lo_p,
    n4206_lo
  );


  not

  (
    n4206_lo_n,
    n4206_lo
  );


  buf

  (
    n4209_lo_p,
    n4209_lo
  );


  not

  (
    n4209_lo_n,
    n4209_lo
  );


  buf

  (
    n4212_lo_p,
    n4212_lo
  );


  not

  (
    n4212_lo_n,
    n4212_lo
  );


  buf

  (
    n4215_lo_p,
    n4215_lo
  );


  not

  (
    n4215_lo_n,
    n4215_lo
  );


  buf

  (
    n4230_lo_p,
    n4230_lo
  );


  not

  (
    n4230_lo_n,
    n4230_lo
  );


  buf

  (
    n4233_lo_p,
    n4233_lo
  );


  not

  (
    n4233_lo_n,
    n4233_lo
  );


  buf

  (
    n4236_lo_p,
    n4236_lo
  );


  not

  (
    n4236_lo_n,
    n4236_lo
  );


  buf

  (
    n4239_lo_p,
    n4239_lo
  );


  not

  (
    n4239_lo_n,
    n4239_lo
  );


  buf

  (
    n4242_lo_p,
    n4242_lo
  );


  not

  (
    n4242_lo_n,
    n4242_lo
  );


  buf

  (
    n4254_lo_p,
    n4254_lo
  );


  not

  (
    n4254_lo_n,
    n4254_lo
  );


  buf

  (
    n4290_lo_p,
    n4290_lo
  );


  not

  (
    n4290_lo_n,
    n4290_lo
  );


  buf

  (
    n4293_lo_p,
    n4293_lo
  );


  not

  (
    n4293_lo_n,
    n4293_lo
  );


  buf

  (
    n4302_lo_p,
    n4302_lo
  );


  not

  (
    n4302_lo_n,
    n4302_lo
  );


  buf

  (
    n4314_lo_p,
    n4314_lo
  );


  not

  (
    n4314_lo_n,
    n4314_lo
  );


  buf

  (
    n4350_lo_p,
    n4350_lo
  );


  not

  (
    n4350_lo_n,
    n4350_lo
  );


  buf

  (
    n4362_lo_p,
    n4362_lo
  );


  not

  (
    n4362_lo_n,
    n4362_lo
  );


  buf

  (
    n4374_lo_p,
    n4374_lo
  );


  not

  (
    n4374_lo_n,
    n4374_lo
  );


  buf

  (
    n4386_lo_p,
    n4386_lo
  );


  not

  (
    n4386_lo_n,
    n4386_lo
  );


  buf

  (
    n4398_lo_p,
    n4398_lo
  );


  not

  (
    n4398_lo_n,
    n4398_lo
  );


  buf

  (
    n4410_lo_p,
    n4410_lo
  );


  not

  (
    n4410_lo_n,
    n4410_lo
  );


  buf

  (
    n4413_lo_p,
    n4413_lo
  );


  not

  (
    n4413_lo_n,
    n4413_lo
  );


  buf

  (
    n4416_lo_p,
    n4416_lo
  );


  not

  (
    n4416_lo_n,
    n4416_lo
  );


  buf

  (
    n4419_lo_p,
    n4419_lo
  );


  not

  (
    n4419_lo_n,
    n4419_lo
  );


  buf

  (
    n4422_lo_p,
    n4422_lo
  );


  not

  (
    n4422_lo_n,
    n4422_lo
  );


  buf

  (
    n4425_lo_p,
    n4425_lo
  );


  not

  (
    n4425_lo_n,
    n4425_lo
  );


  buf

  (
    n4428_lo_p,
    n4428_lo
  );


  not

  (
    n4428_lo_n,
    n4428_lo
  );


  buf

  (
    n4431_lo_p,
    n4431_lo
  );


  not

  (
    n4431_lo_n,
    n4431_lo
  );


  buf

  (
    n4434_lo_p,
    n4434_lo
  );


  not

  (
    n4434_lo_n,
    n4434_lo
  );


  buf

  (
    n4437_lo_p,
    n4437_lo
  );


  not

  (
    n4437_lo_n,
    n4437_lo
  );


  buf

  (
    n4440_lo_p,
    n4440_lo
  );


  not

  (
    n4440_lo_n,
    n4440_lo
  );


  buf

  (
    n4443_lo_p,
    n4443_lo
  );


  not

  (
    n4443_lo_n,
    n4443_lo
  );


  buf

  (
    n4446_lo_p,
    n4446_lo
  );


  not

  (
    n4446_lo_n,
    n4446_lo
  );


  buf

  (
    n4449_lo_p,
    n4449_lo
  );


  not

  (
    n4449_lo_n,
    n4449_lo
  );


  buf

  (
    n4452_lo_p,
    n4452_lo
  );


  not

  (
    n4452_lo_n,
    n4452_lo
  );


  buf

  (
    n4455_lo_p,
    n4455_lo
  );


  not

  (
    n4455_lo_n,
    n4455_lo
  );


  buf

  (
    n4458_lo_p,
    n4458_lo
  );


  not

  (
    n4458_lo_n,
    n4458_lo
  );


  buf

  (
    n4461_lo_p,
    n4461_lo
  );


  not

  (
    n4461_lo_n,
    n4461_lo
  );


  buf

  (
    n4464_lo_p,
    n4464_lo
  );


  not

  (
    n4464_lo_n,
    n4464_lo
  );


  buf

  (
    n4467_lo_p,
    n4467_lo
  );


  not

  (
    n4467_lo_n,
    n4467_lo
  );


  buf

  (
    n4470_lo_p,
    n4470_lo
  );


  not

  (
    n4470_lo_n,
    n4470_lo
  );


  buf

  (
    n4473_lo_p,
    n4473_lo
  );


  not

  (
    n4473_lo_n,
    n4473_lo
  );


  buf

  (
    n4476_lo_p,
    n4476_lo
  );


  not

  (
    n4476_lo_n,
    n4476_lo
  );


  buf

  (
    n4479_lo_p,
    n4479_lo
  );


  not

  (
    n4479_lo_n,
    n4479_lo
  );


  buf

  (
    n4482_lo_p,
    n4482_lo
  );


  not

  (
    n4482_lo_n,
    n4482_lo
  );


  buf

  (
    n4485_lo_p,
    n4485_lo
  );


  not

  (
    n4485_lo_n,
    n4485_lo
  );


  buf

  (
    n4488_lo_p,
    n4488_lo
  );


  not

  (
    n4488_lo_n,
    n4488_lo
  );


  buf

  (
    n4494_lo_p,
    n4494_lo
  );


  not

  (
    n4494_lo_n,
    n4494_lo
  );


  buf

  (
    n4497_lo_p,
    n4497_lo
  );


  not

  (
    n4497_lo_n,
    n4497_lo
  );


  buf

  (
    n4500_lo_p,
    n4500_lo
  );


  not

  (
    n4500_lo_n,
    n4500_lo
  );


  buf

  (
    n4503_lo_p,
    n4503_lo
  );


  not

  (
    n4503_lo_n,
    n4503_lo
  );


  buf

  (
    n4506_lo_p,
    n4506_lo
  );


  not

  (
    n4506_lo_n,
    n4506_lo
  );


  buf

  (
    n4509_lo_p,
    n4509_lo
  );


  not

  (
    n4509_lo_n,
    n4509_lo
  );


  buf

  (
    n4512_lo_p,
    n4512_lo
  );


  not

  (
    n4512_lo_n,
    n4512_lo
  );


  buf

  (
    n4515_lo_p,
    n4515_lo
  );


  not

  (
    n4515_lo_n,
    n4515_lo
  );


  buf

  (
    n4518_lo_p,
    n4518_lo
  );


  not

  (
    n4518_lo_n,
    n4518_lo
  );


  buf

  (
    n4521_lo_p,
    n4521_lo
  );


  not

  (
    n4521_lo_n,
    n4521_lo
  );


  buf

  (
    n4524_lo_p,
    n4524_lo
  );


  not

  (
    n4524_lo_n,
    n4524_lo
  );


  buf

  (
    n4527_lo_p,
    n4527_lo
  );


  not

  (
    n4527_lo_n,
    n4527_lo
  );


  buf

  (
    n4530_lo_p,
    n4530_lo
  );


  not

  (
    n4530_lo_n,
    n4530_lo
  );


  buf

  (
    n4533_lo_p,
    n4533_lo
  );


  not

  (
    n4533_lo_n,
    n4533_lo
  );


  buf

  (
    n4536_lo_p,
    n4536_lo
  );


  not

  (
    n4536_lo_n,
    n4536_lo
  );


  buf

  (
    n4539_lo_p,
    n4539_lo
  );


  not

  (
    n4539_lo_n,
    n4539_lo
  );


  buf

  (
    n4542_lo_p,
    n4542_lo
  );


  not

  (
    n4542_lo_n,
    n4542_lo
  );


  buf

  (
    n4545_lo_p,
    n4545_lo
  );


  not

  (
    n4545_lo_n,
    n4545_lo
  );


  buf

  (
    n4554_lo_p,
    n4554_lo
  );


  not

  (
    n4554_lo_n,
    n4554_lo
  );


  buf

  (
    n4557_lo_p,
    n4557_lo
  );


  not

  (
    n4557_lo_n,
    n4557_lo
  );


  buf

  (
    n4560_lo_p,
    n4560_lo
  );


  not

  (
    n4560_lo_n,
    n4560_lo
  );


  buf

  (
    n4563_lo_p,
    n4563_lo
  );


  not

  (
    n4563_lo_n,
    n4563_lo
  );


  buf

  (
    n4566_lo_p,
    n4566_lo
  );


  not

  (
    n4566_lo_n,
    n4566_lo
  );


  buf

  (
    n4569_lo_p,
    n4569_lo
  );


  not

  (
    n4569_lo_n,
    n4569_lo
  );


  buf

  (
    n4572_lo_p,
    n4572_lo
  );


  not

  (
    n4572_lo_n,
    n4572_lo
  );


  buf

  (
    n4575_lo_p,
    n4575_lo
  );


  not

  (
    n4575_lo_n,
    n4575_lo
  );


  buf

  (
    n4578_lo_p,
    n4578_lo
  );


  not

  (
    n4578_lo_n,
    n4578_lo
  );


  buf

  (
    n4581_lo_p,
    n4581_lo
  );


  not

  (
    n4581_lo_n,
    n4581_lo
  );


  buf

  (
    n4584_lo_p,
    n4584_lo
  );


  not

  (
    n4584_lo_n,
    n4584_lo
  );


  buf

  (
    n4587_lo_p,
    n4587_lo
  );


  not

  (
    n4587_lo_n,
    n4587_lo
  );


  buf

  (
    n4590_lo_p,
    n4590_lo
  );


  not

  (
    n4590_lo_n,
    n4590_lo
  );


  buf

  (
    n4593_lo_p,
    n4593_lo
  );


  not

  (
    n4593_lo_n,
    n4593_lo
  );


  buf

  (
    n4596_lo_p,
    n4596_lo
  );


  not

  (
    n4596_lo_n,
    n4596_lo
  );


  buf

  (
    n4602_lo_p,
    n4602_lo
  );


  not

  (
    n4602_lo_n,
    n4602_lo
  );


  buf

  (
    n4605_lo_p,
    n4605_lo
  );


  not

  (
    n4605_lo_n,
    n4605_lo
  );


  buf

  (
    n4608_lo_p,
    n4608_lo
  );


  not

  (
    n4608_lo_n,
    n4608_lo
  );


  buf

  (
    n4614_lo_p,
    n4614_lo
  );


  not

  (
    n4614_lo_n,
    n4614_lo
  );


  buf

  (
    n4617_lo_p,
    n4617_lo
  );


  not

  (
    n4617_lo_n,
    n4617_lo
  );


  buf

  (
    n4620_lo_p,
    n4620_lo
  );


  not

  (
    n4620_lo_n,
    n4620_lo
  );


  buf

  (
    n4626_lo_p,
    n4626_lo
  );


  not

  (
    n4626_lo_n,
    n4626_lo
  );


  buf

  (
    n4629_lo_p,
    n4629_lo
  );


  not

  (
    n4629_lo_n,
    n4629_lo
  );


  buf

  (
    n4632_lo_p,
    n4632_lo
  );


  not

  (
    n4632_lo_n,
    n4632_lo
  );


  buf

  (
    n4638_lo_p,
    n4638_lo
  );


  not

  (
    n4638_lo_n,
    n4638_lo
  );


  buf

  (
    n4641_lo_p,
    n4641_lo
  );


  not

  (
    n4641_lo_n,
    n4641_lo
  );


  buf

  (
    n4644_lo_p,
    n4644_lo
  );


  not

  (
    n4644_lo_n,
    n4644_lo
  );


  buf

  (
    n4647_lo_p,
    n4647_lo
  );


  not

  (
    n4647_lo_n,
    n4647_lo
  );


  buf

  (
    n4650_lo_p,
    n4650_lo
  );


  not

  (
    n4650_lo_n,
    n4650_lo
  );


  buf

  (
    n4653_lo_p,
    n4653_lo
  );


  not

  (
    n4653_lo_n,
    n4653_lo
  );


  buf

  (
    n4656_lo_p,
    n4656_lo
  );


  not

  (
    n4656_lo_n,
    n4656_lo
  );


  buf

  (
    n4659_lo_p,
    n4659_lo
  );


  not

  (
    n4659_lo_n,
    n4659_lo
  );


  buf

  (
    n4662_lo_p,
    n4662_lo
  );


  not

  (
    n4662_lo_n,
    n4662_lo
  );


  buf

  (
    n4665_lo_p,
    n4665_lo
  );


  not

  (
    n4665_lo_n,
    n4665_lo
  );


  buf

  (
    n4668_lo_p,
    n4668_lo
  );


  not

  (
    n4668_lo_n,
    n4668_lo
  );


  buf

  (
    n4671_lo_p,
    n4671_lo
  );


  not

  (
    n4671_lo_n,
    n4671_lo
  );


  buf

  (
    n4674_lo_p,
    n4674_lo
  );


  not

  (
    n4674_lo_n,
    n4674_lo
  );


  buf

  (
    n4677_lo_p,
    n4677_lo
  );


  not

  (
    n4677_lo_n,
    n4677_lo
  );


  buf

  (
    n4680_lo_p,
    n4680_lo
  );


  not

  (
    n4680_lo_n,
    n4680_lo
  );


  buf

  (
    n4683_lo_p,
    n4683_lo
  );


  not

  (
    n4683_lo_n,
    n4683_lo
  );


  buf

  (
    n4686_lo_p,
    n4686_lo
  );


  not

  (
    n4686_lo_n,
    n4686_lo
  );


  buf

  (
    n4689_lo_p,
    n4689_lo
  );


  not

  (
    n4689_lo_n,
    n4689_lo
  );


  buf

  (
    n4692_lo_p,
    n4692_lo
  );


  not

  (
    n4692_lo_n,
    n4692_lo
  );


  buf

  (
    n4695_lo_p,
    n4695_lo
  );


  not

  (
    n4695_lo_n,
    n4695_lo
  );


  buf

  (
    n4698_lo_p,
    n4698_lo
  );


  not

  (
    n4698_lo_n,
    n4698_lo
  );


  buf

  (
    n4701_lo_p,
    n4701_lo
  );


  not

  (
    n4701_lo_n,
    n4701_lo
  );


  buf

  (
    n4704_lo_p,
    n4704_lo
  );


  not

  (
    n4704_lo_n,
    n4704_lo
  );


  buf

  (
    n4707_lo_p,
    n4707_lo
  );


  not

  (
    n4707_lo_n,
    n4707_lo
  );


  buf

  (
    n4710_lo_p,
    n4710_lo
  );


  not

  (
    n4710_lo_n,
    n4710_lo
  );


  buf

  (
    n4713_lo_p,
    n4713_lo
  );


  not

  (
    n4713_lo_n,
    n4713_lo
  );


  buf

  (
    n4716_lo_p,
    n4716_lo
  );


  not

  (
    n4716_lo_n,
    n4716_lo
  );


  buf

  (
    n4719_lo_p,
    n4719_lo
  );


  not

  (
    n4719_lo_n,
    n4719_lo
  );


  buf

  (
    n4722_lo_p,
    n4722_lo
  );


  not

  (
    n4722_lo_n,
    n4722_lo
  );


  buf

  (
    n4725_lo_p,
    n4725_lo
  );


  not

  (
    n4725_lo_n,
    n4725_lo
  );


  buf

  (
    n4728_lo_p,
    n4728_lo
  );


  not

  (
    n4728_lo_n,
    n4728_lo
  );


  buf

  (
    n4731_lo_p,
    n4731_lo
  );


  not

  (
    n4731_lo_n,
    n4731_lo
  );


  buf

  (
    n4734_lo_p,
    n4734_lo
  );


  not

  (
    n4734_lo_n,
    n4734_lo
  );


  buf

  (
    n4737_lo_p,
    n4737_lo
  );


  not

  (
    n4737_lo_n,
    n4737_lo
  );


  buf

  (
    n4740_lo_p,
    n4740_lo
  );


  not

  (
    n4740_lo_n,
    n4740_lo
  );


  buf

  (
    n4743_lo_p,
    n4743_lo
  );


  not

  (
    n4743_lo_n,
    n4743_lo
  );


  buf

  (
    n4970_o2_p,
    n4970_o2
  );


  not

  (
    n4970_o2_n,
    n4970_o2
  );


  buf

  (
    n4972_o2_p,
    n4972_o2
  );


  not

  (
    n4972_o2_n,
    n4972_o2
  );


  buf

  (
    n4989_o2_p,
    n4989_o2
  );


  not

  (
    n4989_o2_n,
    n4989_o2
  );


  buf

  (
    n5024_o2_p,
    n5024_o2
  );


  not

  (
    n5024_o2_n,
    n5024_o2
  );


  buf

  (
    n5025_o2_p,
    n5025_o2
  );


  not

  (
    n5025_o2_n,
    n5025_o2
  );


  buf

  (
    n5029_o2_p,
    n5029_o2
  );


  not

  (
    n5029_o2_n,
    n5029_o2
  );


  buf

  (
    n5042_o2_p,
    n5042_o2
  );


  not

  (
    n5042_o2_n,
    n5042_o2
  );


  buf

  (
    n5048_o2_p,
    n5048_o2
  );


  not

  (
    n5048_o2_n,
    n5048_o2
  );


  buf

  (
    n5093_o2_p,
    n5093_o2
  );


  not

  (
    n5093_o2_n,
    n5093_o2
  );


  buf

  (
    n5096_o2_p,
    n5096_o2
  );


  not

  (
    n5096_o2_n,
    n5096_o2
  );


  buf

  (
    n5193_o2_p,
    n5193_o2
  );


  not

  (
    n5193_o2_n,
    n5193_o2
  );


  buf

  (
    n5199_o2_p,
    n5199_o2
  );


  not

  (
    n5199_o2_n,
    n5199_o2
  );


  buf

  (
    n5203_o2_p,
    n5203_o2
  );


  not

  (
    n5203_o2_n,
    n5203_o2
  );


  buf

  (
    n5214_o2_p,
    n5214_o2
  );


  not

  (
    n5214_o2_n,
    n5214_o2
  );


  buf

  (
    n5221_o2_p,
    n5221_o2
  );


  not

  (
    n5221_o2_n,
    n5221_o2
  );


  buf

  (
    n5222_o2_p,
    n5222_o2
  );


  not

  (
    n5222_o2_n,
    n5222_o2
  );


  buf

  (
    n5273_o2_p,
    n5273_o2
  );


  not

  (
    n5273_o2_n,
    n5273_o2
  );


  buf

  (
    n5365_o2_p,
    n5365_o2
  );


  not

  (
    n5365_o2_n,
    n5365_o2
  );


  buf

  (
    n5385_o2_p,
    n5385_o2
  );


  not

  (
    n5385_o2_n,
    n5385_o2
  );


  buf

  (
    n5553_o2_p,
    n5553_o2
  );


  not

  (
    n5553_o2_n,
    n5553_o2
  );


  buf

  (
    n5636_o2_p,
    n5636_o2
  );


  not

  (
    n5636_o2_n,
    n5636_o2
  );


  buf

  (
    n5782_o2_p,
    n5782_o2
  );


  not

  (
    n5782_o2_n,
    n5782_o2
  );


  buf

  (
    n5778_o2_p,
    n5778_o2
  );


  not

  (
    n5778_o2_n,
    n5778_o2
  );


  buf

  (
    n5323_o2_p,
    n5323_o2
  );


  not

  (
    n5323_o2_n,
    n5323_o2
  );


  buf

  (
    n5325_o2_p,
    n5325_o2
  );


  not

  (
    n5325_o2_n,
    n5325_o2
  );


  buf

  (
    n5327_o2_p,
    n5327_o2
  );


  not

  (
    n5327_o2_n,
    n5327_o2
  );


  buf

  (
    n5329_o2_p,
    n5329_o2
  );


  not

  (
    n5329_o2_n,
    n5329_o2
  );


  buf

  (
    n5816_o2_p,
    n5816_o2
  );


  not

  (
    n5816_o2_n,
    n5816_o2
  );


  buf

  (
    n5817_o2_p,
    n5817_o2
  );


  not

  (
    n5817_o2_n,
    n5817_o2
  );


  buf

  (
    n5837_o2_p,
    n5837_o2
  );


  not

  (
    n5837_o2_n,
    n5837_o2
  );


  buf

  (
    n5844_o2_p,
    n5844_o2
  );


  not

  (
    n5844_o2_n,
    n5844_o2
  );


  buf

  (
    n5859_o2_p,
    n5859_o2
  );


  not

  (
    n5859_o2_n,
    n5859_o2
  );


  buf

  (
    n5857_o2_p,
    n5857_o2
  );


  not

  (
    n5857_o2_n,
    n5857_o2
  );


  buf

  (
    n5369_o2_p,
    n5369_o2
  );


  not

  (
    n5369_o2_n,
    n5369_o2
  );


  buf

  (
    n5371_o2_p,
    n5371_o2
  );


  not

  (
    n5371_o2_n,
    n5371_o2
  );


  buf

  (
    n5373_o2_p,
    n5373_o2
  );


  not

  (
    n5373_o2_n,
    n5373_o2
  );


  buf

  (
    n5400_o2_p,
    n5400_o2
  );


  not

  (
    n5400_o2_n,
    n5400_o2
  );


  buf

  (
    n5402_o2_p,
    n5402_o2
  );


  not

  (
    n5402_o2_n,
    n5402_o2
  );


  buf

  (
    n5404_o2_p,
    n5404_o2
  );


  not

  (
    n5404_o2_n,
    n5404_o2
  );


  buf

  (
    n5406_o2_p,
    n5406_o2
  );


  not

  (
    n5406_o2_n,
    n5406_o2
  );


  buf

  (
    n5407_o2_p,
    n5407_o2
  );


  not

  (
    n5407_o2_n,
    n5407_o2
  );


  buf

  (
    n5408_o2_p,
    n5408_o2
  );


  not

  (
    n5408_o2_n,
    n5408_o2
  );


  buf

  (
    n2722_o2_p,
    n2722_o2
  );


  not

  (
    n2722_o2_n,
    n2722_o2
  );


  buf

  (
    n1942_inv_p,
    n1942_inv
  );


  not

  (
    n1942_inv_n,
    n1942_inv
  );


  buf

  (
    n5412_o2_p,
    n5412_o2
  );


  not

  (
    n5412_o2_n,
    n5412_o2
  );


  buf

  (
    n1948_inv_p,
    n1948_inv
  );


  not

  (
    n1948_inv_n,
    n1948_inv
  );


  buf

  (
    n5557_o2_p,
    n5557_o2
  );


  not

  (
    n5557_o2_n,
    n5557_o2
  );


  buf

  (
    n5558_o2_p,
    n5558_o2
  );


  not

  (
    n5558_o2_n,
    n5558_o2
  );


  buf

  (
    n5559_o2_p,
    n5559_o2
  );


  not

  (
    n5559_o2_n,
    n5559_o2
  );


  buf

  (
    n5564_o2_p,
    n5564_o2
  );


  not

  (
    n5564_o2_n,
    n5564_o2
  );


  buf

  (
    n5565_o2_p,
    n5565_o2
  );


  not

  (
    n5565_o2_n,
    n5565_o2
  );


  buf

  (
    n1966_inv_p,
    n1966_inv
  );


  not

  (
    n1966_inv_n,
    n1966_inv
  );


  buf

  (
    n5568_o2_p,
    n5568_o2
  );


  not

  (
    n5568_o2_n,
    n5568_o2
  );


  buf

  (
    n5598_o2_p,
    n5598_o2
  );


  not

  (
    n5598_o2_n,
    n5598_o2
  );


  buf

  (
    n5600_o2_p,
    n5600_o2
  );


  not

  (
    n5600_o2_n,
    n5600_o2
  );


  buf

  (
    n5601_o2_p,
    n5601_o2
  );


  not

  (
    n5601_o2_n,
    n5601_o2
  );


  buf

  (
    n5602_o2_p,
    n5602_o2
  );


  not

  (
    n5602_o2_n,
    n5602_o2
  );


  buf

  (
    n5603_o2_p,
    n5603_o2
  );


  not

  (
    n5603_o2_n,
    n5603_o2
  );


  buf

  (
    n2853_o2_p,
    n2853_o2
  );


  not

  (
    n2853_o2_n,
    n2853_o2
  );


  buf

  (
    n5637_o2_p,
    n5637_o2
  );


  not

  (
    n5637_o2_n,
    n5637_o2
  );


  buf

  (
    n1993_inv_p,
    n1993_inv
  );


  not

  (
    n1993_inv_n,
    n1993_inv
  );


  buf

  (
    n1996_inv_p,
    n1996_inv
  );


  not

  (
    n1996_inv_n,
    n1996_inv
  );


  buf

  (
    n5635_o2_p,
    n5635_o2
  );


  not

  (
    n5635_o2_n,
    n5635_o2
  );


  buf

  (
    n5640_o2_p,
    n5640_o2
  );


  not

  (
    n5640_o2_n,
    n5640_o2
  );


  buf

  (
    n5641_o2_p,
    n5641_o2
  );


  not

  (
    n5641_o2_n,
    n5641_o2
  );


  buf

  (
    n5642_o2_p,
    n5642_o2
  );


  not

  (
    n5642_o2_n,
    n5642_o2
  );


  buf

  (
    n5650_o2_p,
    n5650_o2
  );


  not

  (
    n5650_o2_n,
    n5650_o2
  );


  buf

  (
    n5652_o2_p,
    n5652_o2
  );


  not

  (
    n5652_o2_n,
    n5652_o2
  );


  buf

  (
    n5653_o2_p,
    n5653_o2
  );


  not

  (
    n5653_o2_n,
    n5653_o2
  );


  buf

  (
    n5654_o2_p,
    n5654_o2
  );


  not

  (
    n5654_o2_n,
    n5654_o2
  );


  buf

  (
    n5655_o2_p,
    n5655_o2
  );


  not

  (
    n5655_o2_n,
    n5655_o2
  );


  buf

  (
    n5657_o2_p,
    n5657_o2
  );


  not

  (
    n5657_o2_n,
    n5657_o2
  );


  buf

  (
    n2029_inv_p,
    n2029_inv
  );


  not

  (
    n2029_inv_n,
    n2029_inv
  );


  buf

  (
    n5661_o2_p,
    n5661_o2
  );


  not

  (
    n5661_o2_n,
    n5661_o2
  );


  buf

  (
    n5656_o2_p,
    n5656_o2
  );


  not

  (
    n5656_o2_n,
    n5656_o2
  );


  buf

  (
    n5663_o2_p,
    n5663_o2
  );


  not

  (
    n5663_o2_n,
    n5663_o2
  );


  buf

  (
    n2041_inv_p,
    n2041_inv
  );


  not

  (
    n2041_inv_n,
    n2041_inv
  );


  buf

  (
    n5795_o2_p,
    n5795_o2
  );


  not

  (
    n5795_o2_n,
    n5795_o2
  );


  buf

  (
    n5796_o2_p,
    n5796_o2
  );


  not

  (
    n5796_o2_n,
    n5796_o2
  );


  buf

  (
    n5797_o2_p,
    n5797_o2
  );


  not

  (
    n5797_o2_n,
    n5797_o2
  );


  buf

  (
    n5739_o2_p,
    n5739_o2
  );


  not

  (
    n5739_o2_n,
    n5739_o2
  );


  buf

  (
    n5773_o2_p,
    n5773_o2
  );


  not

  (
    n5773_o2_n,
    n5773_o2
  );


  buf

  (
    n2059_inv_p,
    n2059_inv
  );


  not

  (
    n2059_inv_n,
    n2059_inv
  );


  buf

  (
    n5799_o2_p,
    n5799_o2
  );


  not

  (
    n5799_o2_n,
    n5799_o2
  );


  buf

  (
    n5802_o2_p,
    n5802_o2
  );


  not

  (
    n5802_o2_n,
    n5802_o2
  );


  buf

  (
    n2068_inv_p,
    n2068_inv
  );


  not

  (
    n2068_inv_n,
    n2068_inv
  );


  buf

  (
    n5831_o2_p,
    n5831_o2
  );


  not

  (
    n5831_o2_n,
    n5831_o2
  );


  buf

  (
    n5833_o2_p,
    n5833_o2
  );


  not

  (
    n5833_o2_n,
    n5833_o2
  );


  buf

  (
    n5820_o2_p,
    n5820_o2
  );


  not

  (
    n5820_o2_n,
    n5820_o2
  );


  buf

  (
    n5823_o2_p,
    n5823_o2
  );


  not

  (
    n5823_o2_n,
    n5823_o2
  );


  buf

  (
    n5824_o2_p,
    n5824_o2
  );


  not

  (
    n5824_o2_n,
    n5824_o2
  );


  buf

  (
    n5869_o2_p,
    n5869_o2
  );


  not

  (
    n5869_o2_n,
    n5869_o2
  );


  buf

  (
    n5848_o2_p,
    n5848_o2
  );


  not

  (
    n5848_o2_n,
    n5848_o2
  );


  buf

  (
    n5849_o2_p,
    n5849_o2
  );


  not

  (
    n5849_o2_n,
    n5849_o2
  );


  buf

  (
    n5856_o2_p,
    n5856_o2
  );


  not

  (
    n5856_o2_n,
    n5856_o2
  );


  buf

  (
    n5896_o2_p,
    n5896_o2
  );


  not

  (
    n5896_o2_n,
    n5896_o2
  );


  buf

  (
    n2754_o2_p,
    n2754_o2
  );


  not

  (
    n2754_o2_n,
    n2754_o2
  );


  buf

  (
    n2908_o2_p,
    n2908_o2
  );


  not

  (
    n2908_o2_n,
    n2908_o2
  );


  buf

  (
    n5892_o2_p,
    n5892_o2
  );


  not

  (
    n5892_o2_n,
    n5892_o2
  );


  buf

  (
    n5915_o2_p,
    n5915_o2
  );


  not

  (
    n5915_o2_n,
    n5915_o2
  );


  buf

  (
    n5919_o2_p,
    n5919_o2
  );


  not

  (
    n5919_o2_n,
    n5919_o2
  );


  buf

  (
    n5918_o2_p,
    n5918_o2
  );


  not

  (
    n5918_o2_n,
    n5918_o2
  );


  buf

  (
    n5920_o2_p,
    n5920_o2
  );


  not

  (
    n5920_o2_n,
    n5920_o2
  );


  buf

  (
    n5917_o2_p,
    n5917_o2
  );


  not

  (
    n5917_o2_n,
    n5917_o2
  );


  buf

  (
    lo586_buf_o2_p,
    lo586_buf_o2
  );


  not

  (
    lo586_buf_o2_n,
    lo586_buf_o2
  );


  buf

  (
    n2818_o2_p,
    n2818_o2
  );


  not

  (
    n2818_o2_n,
    n2818_o2
  );


  buf

  (
    n2863_o2_p,
    n2863_o2
  );


  not

  (
    n2863_o2_n,
    n2863_o2
  );


  buf

  (
    n2134_inv_p,
    n2134_inv
  );


  not

  (
    n2134_inv_n,
    n2134_inv
  );


  buf

  (
    n2725_o2_p,
    n2725_o2
  );


  not

  (
    n2725_o2_n,
    n2725_o2
  );


  buf

  (
    n3016_o2_p,
    n3016_o2
  );


  not

  (
    n3016_o2_n,
    n3016_o2
  );


  buf

  (
    n3013_o2_p,
    n3013_o2
  );


  not

  (
    n3013_o2_n,
    n3013_o2
  );


  buf

  (
    n2655_o2_p,
    n2655_o2
  );


  not

  (
    n2655_o2_n,
    n2655_o2
  );


  buf

  (
    n2149_inv_p,
    n2149_inv
  );


  not

  (
    n2149_inv_n,
    n2149_inv
  );


  buf

  (
    lo562_buf_o2_p,
    lo562_buf_o2
  );


  not

  (
    lo562_buf_o2_n,
    lo562_buf_o2
  );


  buf

  (
    n2155_inv_p,
    n2155_inv
  );


  not

  (
    n2155_inv_n,
    n2155_inv
  );


  buf

  (
    n2531_o2_p,
    n2531_o2
  );


  not

  (
    n2531_o2_n,
    n2531_o2
  );


  buf

  (
    n2700_o2_p,
    n2700_o2
  );


  not

  (
    n2700_o2_n,
    n2700_o2
  );


  buf

  (
    n5908_o2_p,
    n5908_o2
  );


  not

  (
    n5908_o2_n,
    n5908_o2
  );


  buf

  (
    n5910_o2_p,
    n5910_o2
  );


  not

  (
    n5910_o2_n,
    n5910_o2
  );


  buf

  (
    n5912_o2_p,
    n5912_o2
  );


  not

  (
    n5912_o2_n,
    n5912_o2
  );


  buf

  (
    n5914_o2_p,
    n5914_o2
  );


  not

  (
    n5914_o2_n,
    n5914_o2
  );


  buf

  (
    n2753_o2_p,
    n2753_o2
  );


  not

  (
    n2753_o2_n,
    n2753_o2
  );


  buf

  (
    n2878_o2_p,
    n2878_o2
  );


  not

  (
    n2878_o2_n,
    n2878_o2
  );


  buf

  (
    n2182_inv_p,
    n2182_inv
  );


  not

  (
    n2182_inv_n,
    n2182_inv
  );


  buf

  (
    n5934_o2_p,
    n5934_o2
  );


  not

  (
    n5934_o2_n,
    n5934_o2
  );


  buf

  (
    n5936_o2_p,
    n5936_o2
  );


  not

  (
    n5936_o2_n,
    n5936_o2
  );


  buf

  (
    n5938_o2_p,
    n5938_o2
  );


  not

  (
    n5938_o2_n,
    n5938_o2
  );


  buf

  (
    n2728_o2_p,
    n2728_o2
  );


  not

  (
    n2728_o2_n,
    n2728_o2
  );


  buf

  (
    lo358_buf_o2_p,
    lo358_buf_o2
  );


  not

  (
    lo358_buf_o2_n,
    lo358_buf_o2
  );


  buf

  (
    lo418_buf_o2_p,
    lo418_buf_o2
  );


  not

  (
    lo418_buf_o2_n,
    lo418_buf_o2
  );


  buf

  (
    lo474_buf_o2_p,
    lo474_buf_o2
  );


  not

  (
    lo474_buf_o2_n,
    lo474_buf_o2
  );


  buf

  (
    lo554_buf_o2_p,
    lo554_buf_o2
  );


  not

  (
    lo554_buf_o2_n,
    lo554_buf_o2
  );


  buf

  (
    lo558_buf_o2_p,
    lo558_buf_o2
  );


  not

  (
    lo558_buf_o2_n,
    lo558_buf_o2
  );


  buf

  (
    lo574_buf_o2_p,
    lo574_buf_o2
  );


  not

  (
    lo574_buf_o2_n,
    lo574_buf_o2
  );


  buf

  (
    n2215_inv_p,
    n2215_inv
  );


  not

  (
    n2215_inv_n,
    n2215_inv
  );


  buf

  (
    n2218_inv_p,
    n2218_inv
  );


  not

  (
    n2218_inv_n,
    n2218_inv
  );


  buf

  (
    n2221_inv_p,
    n2221_inv
  );


  not

  (
    n2221_inv_n,
    n2221_inv
  );


  buf

  (
    lo450_buf_o2_p,
    lo450_buf_o2
  );


  not

  (
    lo450_buf_o2_n,
    lo450_buf_o2
  );


  buf

  (
    n2910_o2_p,
    n2910_o2
  );


  not

  (
    n2910_o2_n,
    n2910_o2
  );


  buf

  (
    n2683_o2_p,
    n2683_o2
  );


  not

  (
    n2683_o2_n,
    n2683_o2
  );


  buf

  (
    n2828_o2_p,
    n2828_o2
  );


  not

  (
    n2828_o2_n,
    n2828_o2
  );


  buf

  (
    n2582_o2_p,
    n2582_o2
  );


  not

  (
    n2582_o2_n,
    n2582_o2
  );


  buf

  (
    n2600_o2_p,
    n2600_o2
  );


  not

  (
    n2600_o2_n,
    n2600_o2
  );


  buf

  (
    n2542_o2_p,
    n2542_o2
  );


  not

  (
    n2542_o2_n,
    n2542_o2
  );


  buf

  (
    n2703_o2_p,
    n2703_o2
  );


  not

  (
    n2703_o2_n,
    n2703_o2
  );


  buf

  (
    lo510_buf_o2_p,
    lo510_buf_o2
  );


  not

  (
    lo510_buf_o2_n,
    lo510_buf_o2
  );


  buf

  (
    lo514_buf_o2_p,
    lo514_buf_o2
  );


  not

  (
    lo514_buf_o2_n,
    lo514_buf_o2
  );


  buf

  (
    lo538_buf_o2_p,
    lo538_buf_o2
  );


  not

  (
    lo538_buf_o2_n,
    lo538_buf_o2
  );


  buf

  (
    lo578_buf_o2_p,
    lo578_buf_o2
  );


  not

  (
    lo578_buf_o2_n,
    lo578_buf_o2
  );


  buf

  (
    n2260_inv_p,
    n2260_inv
  );


  not

  (
    n2260_inv_n,
    n2260_inv
  );


  buf

  (
    n2666_o2_p,
    n2666_o2
  );


  not

  (
    n2666_o2_n,
    n2666_o2
  );


  buf

  (
    n2667_o2_p,
    n2667_o2
  );


  not

  (
    n2667_o2_n,
    n2667_o2
  );


  buf

  (
    n2660_o2_p,
    n2660_o2
  );


  not

  (
    n2660_o2_n,
    n2660_o2
  );


  buf

  (
    n2272_inv_p,
    n2272_inv
  );


  not

  (
    n2272_inv_n,
    n2272_inv
  );


  buf

  (
    lo454_buf_o2_p,
    lo454_buf_o2
  );


  not

  (
    lo454_buf_o2_n,
    lo454_buf_o2
  );


  buf

  (
    n3593_o2_p,
    n3593_o2
  );


  not

  (
    n3593_o2_n,
    n3593_o2
  );


  buf

  (
    n3048_o2_p,
    n3048_o2
  );


  not

  (
    n3048_o2_n,
    n3048_o2
  );


  buf

  (
    lo410_buf_o2_p,
    lo410_buf_o2
  );


  not

  (
    lo410_buf_o2_n,
    lo410_buf_o2
  );


  buf

  (
    lo502_buf_o2_p,
    lo502_buf_o2
  );


  not

  (
    lo502_buf_o2_n,
    lo502_buf_o2
  );


  buf

  (
    lo506_buf_o2_p,
    lo506_buf_o2
  );


  not

  (
    lo506_buf_o2_n,
    lo506_buf_o2
  );


  buf

  (
    lo550_buf_o2_p,
    lo550_buf_o2
  );


  not

  (
    lo550_buf_o2_n,
    lo550_buf_o2
  );


  buf

  (
    lo570_buf_o2_p,
    lo570_buf_o2
  );


  not

  (
    lo570_buf_o2_n,
    lo570_buf_o2
  );


  buf

  (
    lo582_buf_o2_p,
    lo582_buf_o2
  );


  not

  (
    lo582_buf_o2_n,
    lo582_buf_o2
  );


  buf

  (
    n2302_inv_p,
    n2302_inv
  );


  not

  (
    n2302_inv_n,
    n2302_inv
  );


  buf

  (
    n2305_inv_p,
    n2305_inv
  );


  not

  (
    n2305_inv_n,
    n2305_inv
  );


  buf

  (
    n3499_o2_p,
    n3499_o2
  );


  not

  (
    n3499_o2_n,
    n3499_o2
  );


  buf

  (
    n2311_inv_p,
    n2311_inv
  );


  not

  (
    n2311_inv_n,
    n2311_inv
  );


  buf

  (
    n2870_o2_p,
    n2870_o2
  );


  not

  (
    n2870_o2_n,
    n2870_o2
  );


  buf

  (
    n2317_inv_p,
    n2317_inv
  );


  not

  (
    n2317_inv_n,
    n2317_inv
  );


  buf

  (
    n2689_o2_p,
    n2689_o2
  );


  not

  (
    n2689_o2_n,
    n2689_o2
  );


  buf

  (
    n2323_inv_p,
    n2323_inv
  );


  not

  (
    n2323_inv_n,
    n2323_inv
  );


  buf

  (
    n2662_o2_p,
    n2662_o2
  );


  not

  (
    n2662_o2_n,
    n2662_o2
  );


  buf

  (
    lo350_buf_o2_p,
    lo350_buf_o2
  );


  not

  (
    lo350_buf_o2_n,
    lo350_buf_o2
  );


  buf

  (
    lo498_buf_o2_p,
    lo498_buf_o2
  );


  not

  (
    lo498_buf_o2_n,
    lo498_buf_o2
  );


  buf

  (
    lo518_buf_o2_p,
    lo518_buf_o2
  );


  not

  (
    lo518_buf_o2_n,
    lo518_buf_o2
  );


  buf

  (
    lo522_buf_o2_p,
    lo522_buf_o2
  );


  not

  (
    lo522_buf_o2_n,
    lo522_buf_o2
  );


  buf

  (
    lo598_buf_o2_p,
    lo598_buf_o2
  );


  not

  (
    lo598_buf_o2_n,
    lo598_buf_o2
  );


  buf

  (
    n2344_inv_p,
    n2344_inv
  );


  not

  (
    n2344_inv_n,
    n2344_inv
  );


  buf

  (
    n2347_inv_p,
    n2347_inv
  );


  not

  (
    n2347_inv_n,
    n2347_inv
  );


  buf

  (
    n2350_inv_p,
    n2350_inv
  );


  not

  (
    n2350_inv_n,
    n2350_inv
  );


  buf

  (
    n2353_inv_p,
    n2353_inv
  );


  not

  (
    n2353_inv_n,
    n2353_inv
  );


  buf

  (
    n2356_inv_p,
    n2356_inv
  );


  not

  (
    n2356_inv_n,
    n2356_inv
  );


  buf

  (
    n2359_inv_p,
    n2359_inv
  );


  not

  (
    n2359_inv_n,
    n2359_inv
  );


  buf

  (
    n2872_o2_p,
    n2872_o2
  );


  not

  (
    n2872_o2_n,
    n2872_o2
  );


  buf

  (
    n3313_o2_p,
    n3313_o2
  );


  not

  (
    n3313_o2_n,
    n3313_o2
  );


  buf

  (
    n3273_o2_p,
    n3273_o2
  );


  not

  (
    n3273_o2_n,
    n3273_o2
  );


  buf

  (
    n2848_o2_p,
    n2848_o2
  );


  not

  (
    n2848_o2_n,
    n2848_o2
  );


  buf

  (
    n2893_o2_p,
    n2893_o2
  );


  not

  (
    n2893_o2_n,
    n2893_o2
  );


  buf

  (
    n3267_o2_p,
    n3267_o2
  );


  not

  (
    n3267_o2_n,
    n3267_o2
  );


  buf

  (
    n2925_o2_p,
    n2925_o2
  );


  not

  (
    n2925_o2_n,
    n2925_o2
  );


  buf

  (
    n2839_o2_p,
    n2839_o2
  );


  not

  (
    n2839_o2_n,
    n2839_o2
  );


  buf

  (
    n2831_o2_p,
    n2831_o2
  );


  not

  (
    n2831_o2_n,
    n2831_o2
  );


  buf

  (
    n2558_o2_p,
    n2558_o2
  );


  not

  (
    n2558_o2_n,
    n2558_o2
  );


  buf

  (
    n2562_o2_p,
    n2562_o2
  );


  not

  (
    n2562_o2_n,
    n2562_o2
  );


  buf

  (
    n2825_o2_p,
    n2825_o2
  );


  not

  (
    n2825_o2_n,
    n2825_o2
  );


  buf

  (
    n3263_o2_p,
    n3263_o2
  );


  not

  (
    n3263_o2_n,
    n3263_o2
  );


  buf

  (
    n3517_o2_p,
    n3517_o2
  );


  not

  (
    n3517_o2_n,
    n3517_o2
  );


  buf

  (
    n2873_o2_p,
    n2873_o2
  );


  not

  (
    n2873_o2_n,
    n2873_o2
  );


  buf

  (
    n2926_o2_p,
    n2926_o2
  );


  not

  (
    n2926_o2_n,
    n2926_o2
  );


  buf

  (
    n3261_o2_p,
    n3261_o2
  );


  not

  (
    n3261_o2_n,
    n3261_o2
  );


  buf

  (
    n3268_o2_p,
    n3268_o2
  );


  not

  (
    n3268_o2_n,
    n3268_o2
  );


  buf

  (
    n3274_o2_p,
    n3274_o2
  );


  not

  (
    n3274_o2_n,
    n3274_o2
  );


  buf

  (
    n3314_o2_p,
    n3314_o2
  );


  not

  (
    n3314_o2_n,
    n3314_o2
  );


  buf

  (
    n3571_o2_p,
    n3571_o2
  );


  not

  (
    n3571_o2_n,
    n3571_o2
  );


  buf

  (
    n2950_o2_p,
    n2950_o2
  );


  not

  (
    n2950_o2_n,
    n2950_o2
  );


  buf

  (
    n2951_o2_p,
    n2951_o2
  );


  not

  (
    n2951_o2_n,
    n2951_o2
  );


  buf

  (
    n3022_o2_p,
    n3022_o2
  );


  not

  (
    n3022_o2_n,
    n3022_o2
  );


  buf

  (
    n3023_o2_p,
    n3023_o2
  );


  not

  (
    n3023_o2_n,
    n3023_o2
  );


  buf

  (
    n3057_o2_p,
    n3057_o2
  );


  not

  (
    n3057_o2_n,
    n3057_o2
  );


  buf

  (
    n3058_o2_p,
    n3058_o2
  );


  not

  (
    n3058_o2_n,
    n3058_o2
  );


  buf

  (
    n2931_o2_p,
    n2931_o2
  );


  not

  (
    n2931_o2_n,
    n2931_o2
  );


  buf

  (
    n2911_o2_p,
    n2911_o2
  );


  not

  (
    n2911_o2_n,
    n2911_o2
  );


  buf

  (
    n2959_o2_p,
    n2959_o2
  );


  not

  (
    n2959_o2_n,
    n2959_o2
  );


  buf

  (
    n2960_o2_p,
    n2960_o2
  );


  not

  (
    n2960_o2_n,
    n2960_o2
  );


  buf

  (
    n2922_o2_p,
    n2922_o2
  );


  not

  (
    n2922_o2_n,
    n2922_o2
  );


  buf

  (
    n2888_o2_p,
    n2888_o2
  );


  not

  (
    n2888_o2_n,
    n2888_o2
  );


  buf

  (
    n2889_o2_p,
    n2889_o2
  );


  not

  (
    n2889_o2_n,
    n2889_o2
  );


  buf

  (
    n3051_o2_p,
    n3051_o2
  );


  not

  (
    n3051_o2_n,
    n3051_o2
  );


  buf

  (
    n3052_o2_p,
    n3052_o2
  );


  not

  (
    n3052_o2_n,
    n3052_o2
  );


  buf

  (
    n3063_o2_p,
    n3063_o2
  );


  not

  (
    n3063_o2_n,
    n3063_o2
  );


  buf

  (
    n2845_o2_p,
    n2845_o2
  );


  not

  (
    n2845_o2_n,
    n2845_o2
  );


  buf

  (
    n2476_inv_p,
    n2476_inv
  );


  not

  (
    n2476_inv_n,
    n2476_inv
  );


  buf

  (
    n3281_o2_p,
    n3281_o2
  );


  not

  (
    n3281_o2_n,
    n3281_o2
  );


  buf

  (
    n3294_o2_p,
    n3294_o2
  );


  not

  (
    n3294_o2_n,
    n3294_o2
  );


  buf

  (
    n2885_o2_p,
    n2885_o2
  );


  not

  (
    n2885_o2_n,
    n2885_o2
  );


  buf

  (
    n2786_o2_p,
    n2786_o2
  );


  not

  (
    n2786_o2_n,
    n2786_o2
  );


  buf

  (
    n2783_o2_p,
    n2783_o2
  );


  not

  (
    n2783_o2_n,
    n2783_o2
  );


  buf

  (
    n2801_o2_p,
    n2801_o2
  );


  not

  (
    n2801_o2_n,
    n2801_o2
  );


  buf

  (
    n2572_o2_p,
    n2572_o2
  );


  not

  (
    n2572_o2_n,
    n2572_o2
  );


  buf

  (
    n2628_o2_p,
    n2628_o2
  );


  not

  (
    n2628_o2_n,
    n2628_o2
  );


  buf

  (
    n2609_o2_p,
    n2609_o2
  );


  not

  (
    n2609_o2_n,
    n2609_o2
  );


  buf

  (
    n2618_o2_p,
    n2618_o2
  );


  not

  (
    n2618_o2_n,
    n2618_o2
  );


  buf

  (
    n2637_o2_p,
    n2637_o2
  );


  not

  (
    n2637_o2_n,
    n2637_o2
  );


  buf

  (
    n2525_o2_p,
    n2525_o2
  );


  not

  (
    n2525_o2_n,
    n2525_o2
  );


  buf

  (
    n2551_o2_p,
    n2551_o2
  );


  not

  (
    n2551_o2_n,
    n2551_o2
  );


  buf

  (
    n3759_o2_p,
    n3759_o2
  );


  not

  (
    n3759_o2_n,
    n3759_o2
  );


  buf

  (
    n2994_o2_p,
    n2994_o2
  );


  not

  (
    n2994_o2_n,
    n2994_o2
  );


  buf

  (
    n3040_o2_p,
    n3040_o2
  );


  not

  (
    n3040_o2_n,
    n3040_o2
  );


  buf

  (
    n2943_o2_p,
    n2943_o2
  );


  not

  (
    n2943_o2_n,
    n2943_o2
  );


  buf

  (
    n2991_o2_p,
    n2991_o2
  );


  not

  (
    n2991_o2_n,
    n2991_o2
  );


  buf

  (
    n3034_o2_p,
    n3034_o2
  );


  not

  (
    n3034_o2_n,
    n3034_o2
  );


  buf

  (
    n2881_o2_p,
    n2881_o2
  );


  not

  (
    n2881_o2_n,
    n2881_o2
  );


  buf

  (
    n3021_o2_p,
    n3021_o2
  );


  not

  (
    n3021_o2_n,
    n3021_o2
  );


  buf

  (
    n3062_o2_p,
    n3062_o2
  );


  not

  (
    n3062_o2_n,
    n3062_o2
  );


  buf

  (
    n2763_o2_p,
    n2763_o2
  );


  not

  (
    n2763_o2_n,
    n2763_o2
  );


  buf

  (
    n2764_o2_p,
    n2764_o2
  );


  not

  (
    n2764_o2_n,
    n2764_o2
  );


  buf

  (
    n2775_o2_p,
    n2775_o2
  );


  not

  (
    n2775_o2_n,
    n2775_o2
  );


  buf

  (
    n2776_o2_p,
    n2776_o2
  );


  not

  (
    n2776_o2_n,
    n2776_o2
  );


  buf

  (
    n2968_o2_p,
    n2968_o2
  );


  not

  (
    n2968_o2_n,
    n2968_o2
  );


  buf

  (
    n2969_o2_p,
    n2969_o2
  );


  not

  (
    n2969_o2_n,
    n2969_o2
  );


  buf

  (
    n2798_o2_p,
    n2798_o2
  );


  not

  (
    n2798_o2_n,
    n2798_o2
  );


  buf

  (
    n3661_o2_p,
    n3661_o2
  );


  not

  (
    n3661_o2_n,
    n3661_o2
  );


  buf

  (
    n2694_o2_p,
    n2694_o2
  );


  not

  (
    n2694_o2_n,
    n2694_o2
  );


  buf

  (
    n2572_inv_p,
    n2572_inv
  );


  not

  (
    n2572_inv_n,
    n2572_inv
  );


  buf

  (
    n2817_o2_p,
    n2817_o2
  );


  not

  (
    n2817_o2_n,
    n2817_o2
  );


  buf

  (
    n2514_o2_p,
    n2514_o2
  );


  not

  (
    n2514_o2_n,
    n2514_o2
  );


  buf

  (
    n2501_o2_p,
    n2501_o2
  );


  not

  (
    n2501_o2_n,
    n2501_o2
  );


  buf

  (
    n2584_inv_p,
    n2584_inv
  );


  not

  (
    n2584_inv_n,
    n2584_inv
  );


  buf

  (
    n2505_o2_p,
    n2505_o2
  );


  not

  (
    n2505_o2_n,
    n2505_o2
  );


  buf

  (
    n2492_o2_p,
    n2492_o2
  );


  not

  (
    n2492_o2_n,
    n2492_o2
  );


  buf

  (
    lo546_buf_o2_p,
    lo546_buf_o2
  );


  not

  (
    lo546_buf_o2_n,
    lo546_buf_o2
  );


  buf

  (
    lo590_buf_o2_p,
    lo590_buf_o2
  );


  not

  (
    lo590_buf_o2_n,
    lo590_buf_o2
  );


  buf

  (
    lo594_buf_o2_p,
    lo594_buf_o2
  );


  not

  (
    lo594_buf_o2_n,
    lo594_buf_o2
  );


  buf

  (
    n2602_inv_p,
    n2602_inv
  );


  not

  (
    n2602_inv_n,
    n2602_inv
  );


  buf

  (
    n2605_inv_p,
    n2605_inv
  );


  not

  (
    n2605_inv_n,
    n2605_inv
  );


  buf

  (
    n2709_o2_p,
    n2709_o2
  );


  not

  (
    n2709_o2_n,
    n2709_o2
  );


  buf

  (
    n2611_inv_p,
    n2611_inv
  );


  not

  (
    n2611_inv_n,
    n2611_inv
  );


  buf

  (
    n2614_inv_p,
    n2614_inv
  );


  not

  (
    n2614_inv_n,
    n2614_inv
  );


  buf

  (
    n2617_inv_p,
    n2617_inv
  );


  not

  (
    n2617_inv_n,
    n2617_inv
  );


  buf

  (
    n2620_inv_p,
    n2620_inv
  );


  not

  (
    n2620_inv_n,
    n2620_inv
  );


  buf

  (
    n3590_o2_p,
    n3590_o2
  );


  not

  (
    n3590_o2_n,
    n3590_o2
  );


  buf

  (
    n3591_o2_p,
    n3591_o2
  );


  not

  (
    n3591_o2_n,
    n3591_o2
  );


  buf

  (
    n2629_inv_p,
    n2629_inv
  );


  not

  (
    n2629_inv_n,
    n2629_inv
  );


  buf

  (
    n3638_o2_p,
    n3638_o2
  );


  not

  (
    n3638_o2_n,
    n3638_o2
  );


  buf

  (
    n3639_o2_p,
    n3639_o2
  );


  not

  (
    n3639_o2_n,
    n3639_o2
  );


  buf

  (
    n2638_inv_p,
    n2638_inv
  );


  not

  (
    n2638_inv_n,
    n2638_inv
  );


  buf

  (
    n2641_inv_p,
    n2641_inv
  );


  not

  (
    n2641_inv_n,
    n2641_inv
  );


  buf

  (
    lo458_buf_o2_p,
    lo458_buf_o2
  );


  not

  (
    lo458_buf_o2_n,
    lo458_buf_o2
  );


  buf

  (
    lo482_buf_o2_p,
    lo482_buf_o2
  );


  not

  (
    lo482_buf_o2_n,
    lo482_buf_o2
  );


  buf

  (
    lo566_buf_o2_p,
    lo566_buf_o2
  );


  not

  (
    lo566_buf_o2_n,
    lo566_buf_o2
  );


  buf

  (
    n2718_o2_p,
    n2718_o2
  );


  not

  (
    n2718_o2_n,
    n2718_o2
  );


  buf

  (
    n3707_o2_p,
    n3707_o2
  );


  not

  (
    n3707_o2_n,
    n3707_o2
  );


  buf

  (
    n3671_o2_p,
    n3671_o2
  );


  not

  (
    n3671_o2_n,
    n3671_o2
  );


  buf

  (
    n3680_o2_p,
    n3680_o2
  );


  not

  (
    n3680_o2_n,
    n3680_o2
  );


  buf

  (
    n3749_o2_p,
    n3749_o2
  );


  not

  (
    n3749_o2_n,
    n3749_o2
  );


  buf

  (
    n3716_o2_p,
    n3716_o2
  );


  not

  (
    n3716_o2_n,
    n3716_o2
  );


  buf

  (
    n3692_o2_p,
    n3692_o2
  );


  not

  (
    n3692_o2_n,
    n3692_o2
  );


  buf

  (
    n2591_o2_p,
    n2591_o2
  );


  not

  (
    n2591_o2_n,
    n2591_o2
  );


  buf

  (
    n3478_o2_p,
    n3478_o2
  );


  not

  (
    n3478_o2_n,
    n3478_o2
  );


  buf

  (
    n3610_o2_p,
    n3610_o2
  );


  not

  (
    n3610_o2_n,
    n3610_o2
  );


  buf

  (
    n3611_o2_p,
    n3611_o2
  );


  not

  (
    n3611_o2_n,
    n3611_o2
  );


  buf

  (
    n2686_inv_p,
    n2686_inv
  );


  not

  (
    n2686_inv_n,
    n2686_inv
  );


  buf

  (
    n2689_inv_p,
    n2689_inv
  );


  not

  (
    n2689_inv_n,
    n2689_inv
  );


  buf

  (
    n2738_o2_p,
    n2738_o2
  );


  not

  (
    n2738_o2_n,
    n2738_o2
  );


  buf

  (
    n3616_o2_p,
    n3616_o2
  );


  not

  (
    n3616_o2_n,
    n3616_o2
  );


  buf

  (
    n3617_o2_p,
    n3617_o2
  );


  not

  (
    n3617_o2_n,
    n3617_o2
  );


  buf

  (
    n3031_o2_p,
    n3031_o2
  );


  not

  (
    n3031_o2_n,
    n3031_o2
  );


  buf

  (
    n2704_inv_p,
    n2704_inv
  );


  not

  (
    n2704_inv_n,
    n2704_inv
  );


  buf

  (
    n3562_o2_p,
    n3562_o2
  );


  not

  (
    n3562_o2_n,
    n3562_o2
  );


  buf

  (
    n2502_o2_p,
    n2502_o2
  );


  not

  (
    n2502_o2_n,
    n2502_o2
  );


  buf

  (
    n3560_o2_p,
    n3560_o2
  );


  not

  (
    n3560_o2_n,
    n3560_o2
  );


  buf

  (
    n3554_o2_p,
    n3554_o2
  );


  not

  (
    n3554_o2_n,
    n3554_o2
  );


  buf

  (
    n3555_o2_p,
    n3555_o2
  );


  not

  (
    n3555_o2_n,
    n3555_o2
  );


  buf

  (
    n3536_o2_p,
    n3536_o2
  );


  not

  (
    n3536_o2_n,
    n3536_o2
  );


  buf

  (
    n3537_o2_p,
    n3537_o2
  );


  not

  (
    n3537_o2_n,
    n3537_o2
  );


  buf

  (
    n3508_o2_p,
    n3508_o2
  );


  not

  (
    n3508_o2_n,
    n3508_o2
  );


  buf

  (
    n3650_o2_p,
    n3650_o2
  );


  not

  (
    n3650_o2_n,
    n3650_o2
  );


  buf

  (
    n3740_o2_p,
    n3740_o2
  );


  not

  (
    n3740_o2_n,
    n3740_o2
  );


  buf

  (
    n3484_o2_p,
    n3484_o2
  );


  not

  (
    n3484_o2_n,
    n3484_o2
  );


  buf

  (
    n2740_inv_p,
    n2740_inv
  );


  not

  (
    n2740_inv_n,
    n2740_inv
  );


  buf

  (
    n2734_o2_p,
    n2734_o2
  );


  not

  (
    n2734_o2_n,
    n2734_o2
  );


  buf

  (
    n2735_o2_p,
    n2735_o2
  );


  not

  (
    n2735_o2_n,
    n2735_o2
  );


  buf

  (
    n2711_o2_p,
    n2711_o2
  );


  not

  (
    n2711_o2_n,
    n2711_o2
  );


  buf

  (
    lo585_buf_o2_p,
    lo585_buf_o2
  );


  not

  (
    lo585_buf_o2_n,
    lo585_buf_o2
  );


  buf

  (
    n2719_o2_p,
    n2719_o2
  );


  not

  (
    n2719_o2_n,
    n2719_o2
  );


  buf

  (
    n2720_o2_p,
    n2720_o2
  );


  not

  (
    n2720_o2_n,
    n2720_o2
  );


  buf

  (
    n2723_o2_p,
    n2723_o2
  );


  not

  (
    n2723_o2_n,
    n2723_o2
  );


  buf

  (
    n2724_o2_p,
    n2724_o2
  );


  not

  (
    n2724_o2_n,
    n2724_o2
  );


  buf

  (
    n3624_o2_p,
    n3624_o2
  );


  not

  (
    n3624_o2_n,
    n3624_o2
  );


  buf

  (
    n3625_o2_p,
    n3625_o2
  );


  not

  (
    n3625_o2_n,
    n3625_o2
  );


  buf

  (
    n3015_o2_p,
    n3015_o2
  );


  not

  (
    n3015_o2_n,
    n3015_o2
  );


  buf

  (
    n3491_o2_p,
    n3491_o2
  );


  not

  (
    n3491_o2_n,
    n3491_o2
  );


  buf

  (
    n2779_inv_p,
    n2779_inv
  );


  not

  (
    n2779_inv_n,
    n2779_inv
  );


  buf

  (
    n2811_o2_p,
    n2811_o2
  );


  not

  (
    n2811_o2_n,
    n2811_o2
  );


  buf

  (
    n3010_o2_p,
    n3010_o2
  );


  not

  (
    n3010_o2_n,
    n3010_o2
  );


  buf

  (
    n3012_o2_p,
    n3012_o2
  );


  not

  (
    n3012_o2_n,
    n3012_o2
  );


  buf

  (
    lo382_buf_o2_p,
    lo382_buf_o2
  );


  not

  (
    lo382_buf_o2_n,
    lo382_buf_o2
  );


  buf

  (
    lo386_buf_o2_p,
    lo386_buf_o2
  );


  not

  (
    lo386_buf_o2_n,
    lo386_buf_o2
  );


  buf

  (
    lo390_buf_o2_p,
    lo390_buf_o2
  );


  not

  (
    lo390_buf_o2_n,
    lo390_buf_o2
  );


  buf

  (
    lo398_buf_o2_p,
    lo398_buf_o2
  );


  not

  (
    lo398_buf_o2_n,
    lo398_buf_o2
  );


  buf

  (
    lo402_buf_o2_p,
    lo402_buf_o2
  );


  not

  (
    lo402_buf_o2_n,
    lo402_buf_o2
  );


  buf

  (
    lo406_buf_o2_p,
    lo406_buf_o2
  );


  not

  (
    lo406_buf_o2_n,
    lo406_buf_o2
  );


  buf

  (
    n3492_o2_p,
    n3492_o2
  );


  not

  (
    n3492_o2_n,
    n3492_o2
  );


  buf

  (
    lo366_buf_o2_p,
    lo366_buf_o2
  );


  not

  (
    lo366_buf_o2_n,
    lo366_buf_o2
  );


  buf

  (
    lo374_buf_o2_p,
    lo374_buf_o2
  );


  not

  (
    lo374_buf_o2_n,
    lo374_buf_o2
  );


  buf

  (
    lo426_buf_o2_p,
    lo426_buf_o2
  );


  not

  (
    lo426_buf_o2_n,
    lo426_buf_o2
  );


  buf

  (
    lo494_buf_o2_p,
    lo494_buf_o2
  );


  not

  (
    lo494_buf_o2_n,
    lo494_buf_o2
  );


  buf

  (
    n2653_o2_p,
    n2653_o2
  );


  not

  (
    n2653_o2_n,
    n2653_o2
  );


  buf

  (
    n2654_o2_p,
    n2654_o2
  );


  not

  (
    n2654_o2_n,
    n2654_o2
  );


  buf

  (
    n2715_o2_p,
    n2715_o2
  );


  not

  (
    n2715_o2_n,
    n2715_o2
  );


  buf

  (
    n2740_o2_p,
    n2740_o2
  );


  not

  (
    n2740_o2_n,
    n2740_o2
  );


  buf

  (
    n2682_o2_p,
    n2682_o2
  );


  not

  (
    n2682_o2_n,
    n2682_o2
  );


  buf

  (
    n2736_o2_p,
    n2736_o2
  );


  not

  (
    n2736_o2_n,
    n2736_o2
  );


  buf

  (
    lo508_buf_o2_p,
    lo508_buf_o2
  );


  not

  (
    lo508_buf_o2_n,
    lo508_buf_o2
  );


  buf

  (
    lo512_buf_o2_p,
    lo512_buf_o2
  );


  not

  (
    lo512_buf_o2_n,
    lo512_buf_o2
  );


  buf

  (
    lo536_buf_o2_p,
    lo536_buf_o2
  );


  not

  (
    lo536_buf_o2_n,
    lo536_buf_o2
  );


  buf

  (
    lo576_buf_o2_p,
    lo576_buf_o2
  );


  not

  (
    lo576_buf_o2_n,
    lo576_buf_o2
  );


  buf

  (
    lo357_buf_o2_p,
    lo357_buf_o2
  );


  not

  (
    lo357_buf_o2_n,
    lo357_buf_o2
  );


  buf

  (
    lo361_buf_o2_p,
    lo361_buf_o2
  );


  not

  (
    lo361_buf_o2_n,
    lo361_buf_o2
  );


  buf

  (
    lo417_buf_o2_p,
    lo417_buf_o2
  );


  not

  (
    lo417_buf_o2_n,
    lo417_buf_o2
  );


  buf

  (
    lo421_buf_o2_p,
    lo421_buf_o2
  );


  not

  (
    lo421_buf_o2_n,
    lo421_buf_o2
  );


  buf

  (
    lo473_buf_o2_p,
    lo473_buf_o2
  );


  not

  (
    lo473_buf_o2_n,
    lo473_buf_o2
  );


  buf

  (
    lo477_buf_o2_p,
    lo477_buf_o2
  );


  not

  (
    lo477_buf_o2_n,
    lo477_buf_o2
  );


  buf

  (
    lo553_buf_o2_p,
    lo553_buf_o2
  );


  not

  (
    lo553_buf_o2_n,
    lo553_buf_o2
  );


  buf

  (
    lo557_buf_o2_p,
    lo557_buf_o2
  );


  not

  (
    lo557_buf_o2_n,
    lo557_buf_o2
  );


  buf

  (
    lo573_buf_o2_p,
    lo573_buf_o2
  );


  not

  (
    lo573_buf_o2_n,
    lo573_buf_o2
  );


  buf

  (
    lo434_buf_o2_p,
    lo434_buf_o2
  );


  not

  (
    lo434_buf_o2_n,
    lo434_buf_o2
  );


  buf

  (
    lo438_buf_o2_p,
    lo438_buf_o2
  );


  not

  (
    lo438_buf_o2_n,
    lo438_buf_o2
  );


  buf

  (
    lo466_buf_o2_p,
    lo466_buf_o2
  );


  not

  (
    lo466_buf_o2_n,
    lo466_buf_o2
  );


  buf

  (
    lo470_buf_o2_p,
    lo470_buf_o2
  );


  not

  (
    lo470_buf_o2_n,
    lo470_buf_o2
  );


  buf

  (
    lo490_buf_o2_p,
    lo490_buf_o2
  );


  not

  (
    lo490_buf_o2_n,
    lo490_buf_o2
  );


  buf

  (
    n2657_o2_p,
    n2657_o2
  );


  not

  (
    n2657_o2_n,
    n2657_o2
  );


  buf

  (
    n2658_o2_p,
    n2658_o2
  );


  not

  (
    n2658_o2_n,
    n2658_o2
  );


  buf

  (
    n2663_o2_p,
    n2663_o2
  );


  not

  (
    n2663_o2_n,
    n2663_o2
  );


  buf

  (
    n2664_o2_p,
    n2664_o2
  );


  not

  (
    n2664_o2_n,
    n2664_o2
  );


  buf

  (
    n2684_o2_p,
    n2684_o2
  );


  not

  (
    n2684_o2_n,
    n2684_o2
  );


  buf

  (
    n2685_o2_p,
    n2685_o2
  );


  not

  (
    n2685_o2_n,
    n2685_o2
  );


  or

  (
    g1049_n,
    n4443_lo_n_spl_,
    n4479_lo_n_spl_
  );


  and

  (
    g1050_p,
    n3399_lo_p_spl_00,
    n3411_lo_p
  );


  and

  (
    g1051_p,
    n2619_lo_p_spl_,
    n4215_lo_p
  );


  and

  (
    g1052_p,
    n3363_lo_p,
    n4587_lo_n_spl_
  );


  or

  (
    g1053_n,
    n2739_lo_n_spl_,
    n4575_lo_p
  );


  or

  (
    g1054_n,
    n4239_lo_n,
    n4455_lo_n
  );


  or

  (
    g1055_n,
    n2739_lo_n_spl_,
    n2751_lo_n
  );


  or

  (
    g1056_n,
    n3387_lo_n,
    g1055_n_spl_000
  );


  or

  (
    g1057_n,
    n3015_lo_n,
    n4563_lo_n_spl_00
  );


  or

  (
    g1058_n,
    n3003_lo_n,
    n4563_lo_p_spl_00
  );


  and

  (
    g1059_p,
    g1057_n,
    g1058_n
  );


  or

  (
    g1060_n,
    g1055_n_spl_000,
    g1059_p
  );


  or

  (
    g1061_n,
    n2763_lo_n,
    n4563_lo_n_spl_00
  );


  or

  (
    g1062_n,
    n3027_lo_n,
    n4563_lo_p_spl_00
  );


  and

  (
    g1063_p,
    g1061_n,
    g1062_n
  );


  or

  (
    g1064_n,
    g1055_n_spl_00,
    g1063_p
  );


  or

  (
    g1065_n,
    n2991_lo_n,
    g1055_n_spl_01
  );


  and

  (
    g1066_p,
    n2715_lo_p,
    n4563_lo_n_spl_01
  );


  and

  (
    g1067_p,
    n2703_lo_p,
    n4563_lo_p_spl_01
  );


  or

  (
    g1068_n,
    g1055_n_spl_01,
    g1067_p
  );


  or

  (
    g1069_n,
    g1066_p,
    g1068_n
  );


  and

  (
    g1070_p,
    n3399_lo_p_spl_00,
    g1069_n
  );


  and

  (
    g1071_p,
    n2967_lo_p,
    n4563_lo_n_spl_01
  );


  and

  (
    g1072_p,
    n2727_lo_p,
    n4563_lo_p_spl_01
  );


  or

  (
    g1073_n,
    g1055_n_spl_10,
    g1072_p
  );


  or

  (
    g1074_n,
    g1071_p,
    g1073_n
  );


  and

  (
    g1075_p,
    n3399_lo_p_spl_01,
    g1074_n
  );


  and

  (
    g1076_p,
    n2691_lo_p,
    n4563_lo_n_spl_1
  );


  and

  (
    g1077_p,
    n2943_lo_p,
    n4563_lo_p_spl_1
  );


  or

  (
    g1078_n,
    g1055_n_spl_10,
    g1077_p
  );


  or

  (
    g1079_n,
    g1076_p,
    g1078_n
  );


  and

  (
    g1080_p,
    n3399_lo_p_spl_01,
    g1079_n
  );


  and

  (
    g1081_p,
    n2955_lo_p,
    n4563_lo_n_spl_1
  );


  and

  (
    g1082_p,
    n2979_lo_p,
    n4563_lo_p_spl_1
  );


  or

  (
    g1083_n,
    g1055_n_spl_11,
    g1082_p
  );


  or

  (
    g1084_n,
    g1081_p,
    g1083_n
  );


  and

  (
    g1085_p,
    n3399_lo_p_spl_1,
    g1084_n
  );


  and

  (
    g1086_p,
    n5859_o2_p,
    n5857_o2_p
  );


  and

  (
    g1087_p,
    n5778_o2_n,
    n2531_o2_p
  );


  and

  (
    g1088_p,
    n2525_o2_p,
    g1087_p
  );


  and

  (
    g1089_p,
    n2542_o2_p,
    n2551_o2_p_spl_
  );


  and

  (
    g1090_p,
    g1088_p,
    g1089_p
  );


  and

  (
    g1091_p,
    g1086_p,
    g1090_p
  );


  and

  (
    g1092_p,
    n2609_o2_p,
    n2618_o2_p
  );


  and

  (
    g1093_p,
    n2628_o2_p,
    g1092_p
  );


  or

  (
    g1094_n,
    n2558_o2_p,
    n2562_o2_p
  );


  and

  (
    g1095_p,
    n2572_o2_p,
    g1094_n_spl_
  );


  and

  (
    g1096_p,
    n5844_o2_p,
    n2582_o2_p
  );


  and

  (
    g1097_p,
    n2600_o2_p,
    n2637_o2_p
  );


  and

  (
    g1098_p,
    g1096_p,
    g1097_p
  );


  and

  (
    g1099_p,
    g1095_p,
    g1098_p
  );


  and

  (
    g1100_p,
    g1093_p,
    g1099_p
  );


  or

  (
    g1101_n,
    n5048_o2_n,
    n5273_o2_n_spl_
  );


  or

  (
    g1102_n,
    n5817_o2_n,
    g1101_n_spl_
  );


  and

  (
    g1103_p,
    n5385_o2_p,
    n2722_o2_n
  );


  and

  (
    g1104_p,
    n5199_o2_p,
    g1103_p
  );


  and

  (
    g1105_p,
    n5222_o2_p,
    n2754_o2_p
  );


  and

  (
    g1106_p,
    g1104_p,
    g1105_p
  );


  and

  (
    g1107_p,
    n2763_o2_n,
    n2764_o2_n
  );


  or

  (
    g1107_n,
    n2763_o2_p,
    n2764_o2_p
  );


  and

  (
    g1108_p,
    n2775_o2_n,
    n2776_o2_n
  );


  or

  (
    g1108_n,
    n2775_o2_p,
    n2776_o2_p
  );


  and

  (
    g1109_p,
    g1107_n,
    g1108_p
  );


  and

  (
    g1110_p,
    g1107_p,
    g1108_n
  );


  or

  (
    g1111_n,
    g1109_p,
    g1110_p
  );


  and

  (
    g1112_p,
    n2786_o2_p_spl_,
    n2783_o2_p_spl_
  );


  or

  (
    g1112_n,
    n2786_o2_n_spl_,
    n2783_o2_n_spl_
  );


  and

  (
    g1113_p,
    n2786_o2_n_spl_,
    n2783_o2_n_spl_
  );


  or

  (
    g1113_n,
    n2786_o2_p_spl_,
    n2783_o2_p_spl_
  );


  and

  (
    g1114_p,
    g1112_n,
    g1113_n
  );


  or

  (
    g1114_n,
    g1112_p,
    g1113_p
  );


  and

  (
    g1115_p,
    n2801_o2_n_spl_,
    n2798_o2_n_spl_
  );


  or

  (
    g1115_n,
    n2801_o2_p_spl_,
    n2798_o2_p_spl_
  );


  and

  (
    g1116_p,
    n2801_o2_p_spl_,
    n2798_o2_p_spl_
  );


  or

  (
    g1116_n,
    n2801_o2_n_spl_,
    n2798_o2_n_spl_
  );


  and

  (
    g1117_p,
    g1115_n,
    g1116_n
  );


  or

  (
    g1117_n,
    g1115_p,
    g1116_p
  );


  and

  (
    g1118_p,
    g1114_n,
    g1117_p
  );


  and

  (
    g1119_p,
    g1114_p,
    g1117_n
  );


  or

  (
    g1120_n,
    g1118_p,
    g1119_p
  );


  or

  (
    g1121_n,
    n5816_o2_n,
    g1101_n_spl_
  );


  or

  (
    g1122_n,
    n5203_o2_n,
    n5273_o2_n_spl_
  );


  or

  (
    g1123_n,
    n5042_o2_n,
    n5221_o2_n
  );


  and

  (
    g1124_p,
    n5193_o2_n,
    g1123_n
  );


  and

  (
    g1125_p,
    g1122_n,
    g1124_p
  );


  and

  (
    g1126_p,
    g1121_n,
    g1125_p
  );


  or

  (
    g1127_n,
    n5214_o2_n,
    n5837_o2_p_spl_0
  );


  and

  (
    g1128_p,
    n2828_o2_n,
    n2825_o2_p_spl_000
  );


  or

  (
    g1129_n,
    n4731_lo_n_spl_000,
    n5778_o2_p
  );


  and

  (
    g1130_p,
    n4719_lo_p_spl_000,
    n2831_o2_p
  );


  and

  (
    g1131_p,
    g1129_n,
    g1130_p
  );


  or

  (
    g1132_n,
    g1128_p,
    g1131_p
  );


  or

  (
    g1133_n,
    n5365_o2_n,
    n2825_o2_n_spl_
  );


  and

  (
    g1134_p,
    n4731_lo_p_spl_000,
    n2551_o2_p_spl_
  );


  or

  (
    g1135_n,
    n4719_lo_n_spl_0,
    n2839_o2_n
  );


  or

  (
    g1136_n,
    g1134_p,
    g1135_n
  );


  and

  (
    g1137_p,
    g1133_n,
    g1136_n
  );


  and

  (
    g1138_p,
    n2825_o2_p_spl_000,
    n2845_o2_p_spl_
  );


  or

  (
    g1139_n,
    n4731_lo_n_spl_000,
    n2572_o2_n
  );


  and

  (
    g1140_p,
    n4719_lo_p_spl_000,
    n2848_o2_p
  );


  and

  (
    g1141_p,
    g1139_n,
    g1140_p
  );


  or

  (
    g1142_n,
    g1138_p,
    g1141_p
  );


  or

  (
    g1143_n,
    n4683_lo_n_spl_0000,
    g1132_n_spl_00
  );


  or

  (
    g1144_n,
    n4683_lo_p_spl_0000,
    g1142_n_spl_00
  );


  and

  (
    g1145_p,
    g1143_n,
    g1144_n
  );


  and

  (
    g1146_p,
    n4671_lo_p_spl_000,
    g1145_p
  );


  or

  (
    g1147_n,
    n2643_lo_p_spl_,
    n4683_lo_n_spl_0000
  );


  or

  (
    g1148_n,
    n2871_lo_p_spl_,
    n4683_lo_p_spl_0000
  );


  and

  (
    g1149_p,
    g1147_n,
    g1148_n
  );


  and

  (
    g1150_p,
    n4671_lo_n_spl_000,
    g1149_p
  );


  or

  (
    g1151_n,
    g1146_p,
    g1150_p
  );


  and

  (
    g1152_p,
    n5636_o2_n_spl_,
    n2825_o2_p_spl_001
  );


  or

  (
    g1153_n,
    n2872_o2_p,
    n2873_o2_p
  );


  and

  (
    g1154_p,
    n4719_lo_p_spl_001,
    g1153_n
  );


  or

  (
    g1155_n,
    g1152_p,
    g1154_p
  );


  and

  (
    g1156_p,
    n2825_o2_p_spl_001,
    n2881_o2_n_spl_
  );


  and

  (
    g1157_p,
    n4719_lo_p_spl_001,
    n2885_o2_p
  );


  or

  (
    g1158_n,
    g1156_p,
    g1157_p
  );


  or

  (
    g1159_n,
    n2888_o2_p,
    n2889_o2_n
  );


  and

  (
    g1160_p,
    n2825_o2_p_spl_010,
    g1159_n_spl_
  );


  or

  (
    g1161_n,
    n4731_lo_n_spl_00,
    n2525_o2_n
  );


  and

  (
    g1162_p,
    n4719_lo_p_spl_010,
    n2893_o2_p
  );


  and

  (
    g1163_p,
    g1161_n,
    g1162_p
  );


  or

  (
    g1164_n,
    g1160_p,
    g1163_p
  );


  or

  (
    g1165_n,
    n4695_lo_n_spl_0000,
    g1132_n_spl_00
  );


  or

  (
    g1166_n,
    n4695_lo_p_spl_0000,
    g1142_n_spl_00
  );


  and

  (
    g1167_p,
    g1165_n,
    g1166_n
  );


  and

  (
    g1168_p,
    n4707_lo_p_spl_000,
    g1167_p
  );


  or

  (
    g1169_n,
    n2643_lo_p_spl_,
    n4695_lo_n_spl_0000
  );


  or

  (
    g1170_n,
    n2871_lo_p_spl_,
    n4695_lo_p_spl_0000
  );


  and

  (
    g1171_p,
    g1169_n,
    g1170_n
  );


  and

  (
    g1172_p,
    n4707_lo_n_spl_000,
    g1171_p
  );


  or

  (
    g1173_n,
    g1168_p,
    g1172_p
  );


  and

  (
    g1174_p,
    n5553_o2_n,
    n2911_o2_n
  );


  and

  (
    g1175_p,
    n5553_o2_p,
    n2911_o2_p
  );


  or

  (
    g1176_n,
    g1174_p,
    g1175_p
  );


  and

  (
    g1177_p,
    n2825_o2_p_spl_010,
    g1176_n_spl_
  );


  and

  (
    g1178_p,
    n3243_lo_p,
    n4731_lo_n_spl_01
  );


  and

  (
    g1179_p,
    n4731_lo_p_spl_000,
    n2609_o2_n
  );


  or

  (
    g1180_n,
    g1178_p,
    g1179_p
  );


  and

  (
    g1181_p,
    n4719_lo_p_spl_010,
    g1180_n
  );


  or

  (
    g1182_n,
    g1177_p,
    g1181_p
  );


  or

  (
    g1183_n,
    n2910_o2_p,
    n2922_o2_n
  );


  and

  (
    g1184_p,
    n2825_o2_p_spl_011,
    g1183_n_spl_
  );


  or

  (
    g1185_n,
    n2925_o2_p,
    n2926_o2_p
  );


  and

  (
    g1186_p,
    n4719_lo_p_spl_011,
    g1185_n
  );


  or

  (
    g1187_n,
    g1184_p,
    g1186_p
  );


  or

  (
    g1188_n,
    n2908_o2_p,
    n2931_o2_n
  );


  and

  (
    g1189_p,
    n2825_o2_p_spl_011,
    g1188_n_spl_
  );


  and

  (
    g1190_p,
    n3279_lo_p,
    n4731_lo_n_spl_01
  );


  and

  (
    g1191_p,
    n4731_lo_p_spl_00,
    n2628_o2_n
  );


  or

  (
    g1192_n,
    g1190_p,
    g1191_p
  );


  and

  (
    g1193_p,
    n4719_lo_p_spl_011,
    g1192_n
  );


  or

  (
    g1194_n,
    g1189_p,
    g1193_p
  );


  or

  (
    g1195_n,
    n2825_o2_n_spl_,
    n2943_o2_p
  );


  and

  (
    g1196_p,
    n4731_lo_p_spl_01,
    g1094_n_spl_
  );


  and

  (
    g1197_p,
    n3267_lo_n,
    n4731_lo_n_spl_10
  );


  or

  (
    g1198_n,
    n4719_lo_n_spl_0,
    g1197_p
  );


  or

  (
    g1199_n,
    g1196_p,
    g1198_n
  );


  and

  (
    g1200_p,
    g1195_n,
    g1199_n
  );


  and

  (
    g1201_p,
    n2950_o2_n,
    n2951_o2_n
  );


  or

  (
    g1201_n,
    n2950_o2_p,
    n2951_o2_p
  );


  and

  (
    g1202_p,
    n2853_o2_n_spl_00,
    g1201_n_spl_
  );


  or

  (
    g1202_n,
    n2853_o2_p_spl_0,
    g1201_p_spl_
  );


  and

  (
    g1203_p,
    n2853_o2_p_spl_0,
    g1201_p_spl_
  );


  or

  (
    g1203_n,
    n2853_o2_n_spl_00,
    g1201_n_spl_
  );


  and

  (
    g1204_p,
    g1202_n,
    g1203_n
  );


  or

  (
    g1204_n,
    g1202_p,
    g1203_p
  );


  and

  (
    g1205_p,
    n2959_o2_p,
    n2960_o2_n
  );


  or

  (
    g1205_n,
    n2959_o2_n,
    n2960_o2_p
  );


  and

  (
    g1206_p,
    n2968_o2_p,
    n2969_o2_n
  );


  or

  (
    g1206_n,
    n2968_o2_n,
    n2969_o2_p
  );


  and

  (
    g1207_p,
    g1205_p_spl_,
    g1206_n_spl_
  );


  or

  (
    g1207_n,
    g1205_n_spl_,
    g1206_p_spl_
  );


  and

  (
    g1208_p,
    g1205_n_spl_,
    g1206_p_spl_
  );


  or

  (
    g1208_n,
    g1205_p_spl_,
    g1206_n_spl_
  );


  and

  (
    g1209_p,
    g1207_n,
    g1208_n
  );


  or

  (
    g1209_n,
    g1207_p,
    g1208_p
  );


  and

  (
    g1210_p,
    g1204_n,
    g1209_p
  );


  and

  (
    g1211_p,
    g1204_p,
    g1209_n
  );


  or

  (
    g1212_n,
    g1210_p,
    g1211_p
  );


  and

  (
    g1213_p,
    n4972_o2_n_spl_,
    n4989_o2_p_spl_
  );


  or

  (
    g1213_n,
    n4972_o2_p_spl_,
    n4989_o2_n_spl_
  );


  and

  (
    g1214_p,
    n4972_o2_p_spl_,
    n4989_o2_n_spl_
  );


  or

  (
    g1214_n,
    n4972_o2_n_spl_,
    n4989_o2_p_spl_
  );


  and

  (
    g1215_p,
    g1213_n,
    g1214_n
  );


  or

  (
    g1215_n,
    g1213_p,
    g1214_p
  );


  and

  (
    g1216_p,
    n5025_o2_n_spl_,
    n5093_o2_p_spl_
  );


  or

  (
    g1216_n,
    n5025_o2_p_spl_,
    n5093_o2_n_spl_
  );


  and

  (
    g1217_p,
    n5025_o2_p_spl_,
    n5093_o2_n_spl_
  );


  or

  (
    g1217_n,
    n5025_o2_n_spl_,
    n5093_o2_p_spl_
  );


  and

  (
    g1218_p,
    g1216_n,
    g1217_n
  );


  or

  (
    g1218_n,
    g1216_p,
    g1217_p
  );


  and

  (
    g1219_p,
    g1215_n_spl_,
    g1218_p_spl_
  );


  or

  (
    g1219_n,
    g1215_p_spl_,
    g1218_n_spl_
  );


  and

  (
    g1220_p,
    g1215_p_spl_,
    g1218_n_spl_
  );


  or

  (
    g1220_n,
    g1215_n_spl_,
    g1218_p_spl_
  );


  and

  (
    g1221_p,
    g1219_n,
    g1220_n
  );


  or

  (
    g1221_n,
    g1219_p,
    g1220_p
  );


  and

  (
    g1222_p,
    n2994_o2_n_spl_,
    n2991_o2_p_spl_
  );


  or

  (
    g1222_n,
    n2994_o2_p_spl_,
    n2991_o2_n_spl_
  );


  and

  (
    g1223_p,
    n2994_o2_p_spl_,
    n2991_o2_n_spl_
  );


  or

  (
    g1223_n,
    n2994_o2_n_spl_,
    n2991_o2_p_spl_
  );


  and

  (
    g1224_p,
    g1222_n,
    g1223_n
  );


  or

  (
    g1224_n,
    g1222_p,
    g1223_p
  );


  and

  (
    g1225_p,
    n4970_o2_p_spl_,
    n5024_o2_n_spl_
  );


  or

  (
    g1225_n,
    n4970_o2_n_spl_,
    n5024_o2_p_spl_
  );


  and

  (
    g1226_p,
    n4970_o2_n_spl_,
    n5024_o2_p_spl_
  );


  or

  (
    g1226_n,
    n4970_o2_p_spl_,
    n5024_o2_n_spl_
  );


  and

  (
    g1227_p,
    g1225_n,
    g1226_n
  );


  or

  (
    g1227_n,
    g1225_p,
    g1226_p
  );


  and

  (
    g1228_p,
    g1224_n_spl_,
    g1227_p_spl_
  );


  or

  (
    g1228_n,
    g1224_p_spl_,
    g1227_n_spl_
  );


  and

  (
    g1229_p,
    g1224_p_spl_,
    g1227_n_spl_
  );


  or

  (
    g1229_n,
    g1224_n_spl_,
    g1227_p_spl_
  );


  and

  (
    g1230_p,
    g1228_n,
    g1229_n
  );


  or

  (
    g1230_n,
    g1228_p,
    g1229_p
  );


  and

  (
    g1231_p,
    g1221_n,
    g1230_p
  );


  and

  (
    g1232_p,
    g1221_p,
    g1230_n
  );


  or

  (
    g1233_n,
    g1231_p,
    g1232_p
  );


  or

  (
    g1234_n,
    n3022_o2_p,
    n3023_o2_p
  );


  or

  (
    g1235_n,
    n2845_o2_p_spl_,
    n2943_o2_n
  );


  or

  (
    g1236_n,
    g1188_n_spl_,
    g1235_n
  );


  or

  (
    g1237_n,
    g1183_n_spl_,
    g1236_n
  );


  or

  (
    g1238_n,
    g1176_n_spl_,
    g1237_n
  );


  or

  (
    g1239_n,
    g1234_n_spl_,
    g1238_n
  );


  or

  (
    g1240_n,
    n3021_o2_n_spl_,
    g1239_n
  );


  or

  (
    g1241_n,
    n5096_o2_n,
    n3034_o2_p
  );


  or

  (
    g1242_n,
    n5096_o2_p,
    n3034_o2_n
  );


  and

  (
    g1243_p,
    g1241_n,
    g1242_n
  );


  or

  (
    g1244_n,
    n5029_o2_n,
    n3040_o2_n
  );


  or

  (
    g1245_n,
    n5029_o2_p,
    n3040_o2_p
  );


  and

  (
    g1246_p,
    g1244_n,
    g1245_n
  );


  or

  (
    g1247_n,
    g1243_p_spl_,
    g1246_p_spl_
  );


  or

  (
    g1248_n,
    g1240_n,
    g1247_n
  );


  and

  (
    g1249_p,
    n3051_o2_p,
    n3052_o2_n
  );


  and

  (
    g1250_p,
    n3057_o2_n,
    n3058_o2_p
  );


  or

  (
    g1251_n,
    n5365_o2_p,
    n3063_o2_n
  );


  or

  (
    g1252_n,
    g1159_n_spl_,
    g1251_n
  );


  or

  (
    g1253_n,
    n5636_o2_n_spl_,
    g1252_n
  );


  or

  (
    g1254_n,
    n2881_o2_n_spl_,
    g1253_n
  );


  or

  (
    g1255_n,
    n3062_o2_p_spl_,
    g1254_n
  );


  or

  (
    g1256_n,
    g1250_p_spl_,
    g1255_n
  );


  or

  (
    g1257_n,
    g1249_p_spl_,
    g1256_n
  );


  and

  (
    g1258_p,
    n4503_lo_n_spl_0000,
    g1142_n_spl_0
  );


  and

  (
    g1259_p,
    n4503_lo_p_spl_0000,
    g1132_n_spl_0
  );


  or

  (
    g1260_n,
    n4515_lo_n_spl_000,
    g1259_p
  );


  or

  (
    g1261_n,
    g1258_p,
    g1260_n
  );


  and

  (
    g1262_p,
    n3579_lo_p_spl_,
    n4503_lo_n_spl_0000
  );


  and

  (
    g1263_p,
    n3567_lo_p_spl_,
    n4503_lo_p_spl_0000
  );


  or

  (
    g1264_n,
    n4515_lo_p_spl_000,
    g1263_p
  );


  or

  (
    g1265_n,
    g1262_p,
    g1264_n
  );


  and

  (
    g1266_p,
    n3375_lo_p_spl_0000,
    g1265_n
  );


  and

  (
    g1267_p,
    g1261_n,
    g1266_p
  );


  and

  (
    g1268_p,
    n4527_lo_n_spl_0000,
    g1142_n_spl_1
  );


  and

  (
    g1269_p,
    n4527_lo_p_spl_0000,
    g1132_n_spl_1
  );


  or

  (
    g1270_n,
    n4539_lo_n_spl_000,
    g1269_p
  );


  or

  (
    g1271_n,
    g1268_p,
    g1270_n
  );


  and

  (
    g1272_p,
    n3579_lo_p_spl_,
    n4527_lo_n_spl_0000
  );


  and

  (
    g1273_p,
    n3567_lo_p_spl_,
    n4527_lo_p_spl_0000
  );


  or

  (
    g1274_n,
    n4539_lo_p_spl_000,
    g1273_p
  );


  or

  (
    g1275_n,
    g1272_p,
    g1274_n
  );


  and

  (
    g1276_p,
    n3375_lo_p_spl_0000,
    g1275_n
  );


  and

  (
    g1277_p,
    g1271_n,
    g1276_p
  );


  or

  (
    g1278_n,
    n2775_lo_p_spl_,
    n4683_lo_p_spl_0001
  );


  or

  (
    g1279_n,
    n2799_lo_p_spl_,
    n4683_lo_n_spl_0001
  );


  and

  (
    g1280_p,
    g1278_n,
    g1279_n
  );


  or

  (
    g1281_n,
    n4671_lo_p_spl_000,
    g1280_p
  );


  and

  (
    g1282_p,
    n4683_lo_n_spl_0001,
    g1182_n_spl_00
  );


  and

  (
    g1283_p,
    n4683_lo_p_spl_0001,
    g1155_n_spl_00
  );


  or

  (
    g1284_n,
    n4671_lo_n_spl_000,
    g1283_p
  );


  or

  (
    g1285_n,
    g1282_p,
    g1284_n
  );


  and

  (
    g1286_p,
    g1281_n,
    g1285_n
  );


  or

  (
    g1287_n,
    n2679_lo_p_spl_,
    n4683_lo_p_spl_0010
  );


  or

  (
    g1288_n,
    n2931_lo_p_spl_,
    n4683_lo_n_spl_0010
  );


  and

  (
    g1289_p,
    g1287_n,
    g1288_n
  );


  or

  (
    g1290_n,
    n4671_lo_p_spl_001,
    g1289_p
  );


  and

  (
    g1291_p,
    n4683_lo_n_spl_0010,
    g1187_n_spl_00
  );


  and

  (
    g1292_p,
    n4683_lo_p_spl_0010,
    g1158_n_spl_00
  );


  or

  (
    g1293_n,
    n4671_lo_n_spl_001,
    g1292_p
  );


  or

  (
    g1294_n,
    g1291_p,
    g1293_n
  );


  and

  (
    g1295_p,
    g1290_n,
    g1294_n
  );


  or

  (
    g1296_n,
    n2667_lo_p_spl_,
    n4683_lo_p_spl_0011
  );


  or

  (
    g1297_n,
    n2919_lo_p_spl_,
    n4683_lo_n_spl_0011
  );


  and

  (
    g1298_p,
    g1296_n,
    g1297_n
  );


  or

  (
    g1299_n,
    n4671_lo_p_spl_001,
    g1298_p
  );


  and

  (
    g1300_p,
    n4683_lo_n_spl_0011,
    g1194_n_spl_00
  );


  and

  (
    g1301_p,
    n4683_lo_p_spl_0011,
    g1164_n_spl_00
  );


  or

  (
    g1302_n,
    n4671_lo_n_spl_001,
    g1301_p
  );


  or

  (
    g1303_n,
    g1300_p,
    g1302_n
  );


  and

  (
    g1304_p,
    g1299_n,
    g1303_n
  );


  or

  (
    g1305_n,
    n2907_lo_n_spl_,
    n4683_lo_p_spl_010
  );


  or

  (
    g1306_n,
    n2895_lo_n_spl_,
    n4683_lo_n_spl_010
  );


  and

  (
    g1307_p,
    g1305_n,
    g1306_n
  );


  or

  (
    g1308_n,
    n4671_lo_p_spl_01,
    g1307_p
  );


  and

  (
    g1309_p,
    n4683_lo_n_spl_010,
    g1200_p_spl_00
  );


  and

  (
    g1310_p,
    n4683_lo_p_spl_010,
    g1137_p_spl_00
  );


  or

  (
    g1311_n,
    n4671_lo_n_spl_01,
    g1310_p
  );


  or

  (
    g1312_n,
    g1309_p,
    g1311_n
  );


  and

  (
    g1313_p,
    g1308_n,
    g1312_n
  );


  or

  (
    g1314_n,
    n2775_lo_p_spl_,
    n4695_lo_p_spl_0001
  );


  or

  (
    g1315_n,
    n2799_lo_p_spl_,
    n4695_lo_n_spl_0001
  );


  and

  (
    g1316_p,
    g1314_n,
    g1315_n
  );


  or

  (
    g1317_n,
    n4707_lo_p_spl_000,
    g1316_p
  );


  and

  (
    g1318_p,
    n4695_lo_n_spl_0001,
    g1182_n_spl_00
  );


  and

  (
    g1319_p,
    n4695_lo_p_spl_0001,
    g1155_n_spl_00
  );


  or

  (
    g1320_n,
    n4707_lo_n_spl_000,
    g1319_p
  );


  or

  (
    g1321_n,
    g1318_p,
    g1320_n
  );


  and

  (
    g1322_p,
    g1317_n,
    g1321_n
  );


  or

  (
    g1323_n,
    n2679_lo_p_spl_,
    n4695_lo_p_spl_0010
  );


  or

  (
    g1324_n,
    n2931_lo_p_spl_,
    n4695_lo_n_spl_0010
  );


  and

  (
    g1325_p,
    g1323_n,
    g1324_n
  );


  or

  (
    g1326_n,
    n4707_lo_p_spl_001,
    g1325_p
  );


  and

  (
    g1327_p,
    n4695_lo_n_spl_0010,
    g1187_n_spl_00
  );


  and

  (
    g1328_p,
    n4695_lo_p_spl_0010,
    g1158_n_spl_00
  );


  or

  (
    g1329_n,
    n4707_lo_n_spl_001,
    g1328_p
  );


  or

  (
    g1330_n,
    g1327_p,
    g1329_n
  );


  and

  (
    g1331_p,
    g1326_n,
    g1330_n
  );


  or

  (
    g1332_n,
    n2667_lo_p_spl_,
    n4695_lo_p_spl_0011
  );


  or

  (
    g1333_n,
    n2919_lo_p_spl_,
    n4695_lo_n_spl_0011
  );


  and

  (
    g1334_p,
    g1332_n,
    g1333_n
  );


  or

  (
    g1335_n,
    n4707_lo_p_spl_001,
    g1334_p
  );


  and

  (
    g1336_p,
    n4695_lo_n_spl_0011,
    g1194_n_spl_00
  );


  and

  (
    g1337_p,
    n4695_lo_p_spl_0011,
    g1164_n_spl_00
  );


  or

  (
    g1338_n,
    n4707_lo_n_spl_001,
    g1337_p
  );


  or

  (
    g1339_n,
    g1336_p,
    g1338_n
  );


  and

  (
    g1340_p,
    g1335_n,
    g1339_n
  );


  or

  (
    g1341_n,
    n2907_lo_n_spl_,
    n4695_lo_p_spl_010
  );


  or

  (
    g1342_n,
    n2895_lo_n_spl_,
    n4695_lo_n_spl_010
  );


  and

  (
    g1343_p,
    g1341_n,
    g1342_n
  );


  or

  (
    g1344_n,
    n4707_lo_p_spl_01,
    g1343_p
  );


  and

  (
    g1345_p,
    n4695_lo_n_spl_010,
    g1200_p_spl_00
  );


  and

  (
    g1346_p,
    n4695_lo_p_spl_010,
    g1137_p_spl_00
  );


  or

  (
    g1347_n,
    n4707_lo_n_spl_01,
    g1346_p
  );


  or

  (
    g1348_n,
    g1345_p,
    g1347_n
  );


  and

  (
    g1349_p,
    g1344_n,
    g1348_n
  );


  and

  (
    g1350_p,
    n4503_lo_n_spl_0001,
    g1182_n_spl_0
  );


  and

  (
    g1351_p,
    n4503_lo_p_spl_0001,
    g1155_n_spl_0
  );


  or

  (
    g1352_n,
    n4515_lo_n_spl_000,
    g1351_p
  );


  or

  (
    g1353_n,
    g1350_p,
    g1352_n
  );


  and

  (
    g1354_p,
    n3519_lo_p_spl_,
    n4503_lo_n_spl_0001
  );


  and

  (
    g1355_p,
    n3639_lo_p_spl_,
    n4503_lo_p_spl_0001
  );


  or

  (
    g1356_n,
    n4515_lo_p_spl_000,
    g1355_p
  );


  or

  (
    g1357_n,
    g1354_p,
    g1356_n
  );


  and

  (
    g1358_p,
    n3375_lo_p_spl_000,
    g1357_n
  );


  and

  (
    g1359_p,
    g1353_n,
    g1358_p
  );


  or

  (
    g1360_n,
    n4503_lo_p_spl_0010,
    g1200_p_spl_0
  );


  or

  (
    g1361_n,
    n4503_lo_n_spl_0010,
    g1137_p_spl_0
  );


  and

  (
    g1362_p,
    n4515_lo_p_spl_001,
    g1361_n
  );


  and

  (
    g1363_p,
    g1360_n,
    g1362_p
  );


  or

  (
    g1364_n,
    n3471_lo_n_spl_,
    n4503_lo_p_spl_0010
  );


  or

  (
    g1365_n,
    n3591_lo_n_spl_,
    n4503_lo_n_spl_0010
  );


  and

  (
    g1366_p,
    n4515_lo_n_spl_001,
    g1365_n
  );


  and

  (
    g1367_p,
    g1364_n,
    g1366_p
  );


  or

  (
    g1368_n,
    n3375_lo_n_spl_0,
    g1367_p
  );


  or

  (
    g1369_n,
    g1363_p,
    g1368_n
  );


  and

  (
    g1370_p,
    n4503_lo_n_spl_0011,
    g1194_n_spl_0
  );


  and

  (
    g1371_p,
    n4503_lo_p_spl_0011,
    g1164_n_spl_0
  );


  or

  (
    g1372_n,
    n4515_lo_n_spl_001,
    g1371_p
  );


  or

  (
    g1373_n,
    g1370_p,
    g1372_n
  );


  and

  (
    g1374_p,
    n3447_lo_p_spl_,
    n4503_lo_n_spl_0011
  );


  and

  (
    g1375_p,
    n3459_lo_p_spl_,
    n4503_lo_p_spl_0011
  );


  or

  (
    g1376_n,
    n4515_lo_p_spl_001,
    g1375_p
  );


  or

  (
    g1377_n,
    g1374_p,
    g1376_n
  );


  and

  (
    g1378_p,
    n3375_lo_p_spl_001,
    g1377_n
  );


  and

  (
    g1379_p,
    g1373_n,
    g1378_p
  );


  and

  (
    g1380_p,
    n4503_lo_n_spl_010,
    g1187_n_spl_0
  );


  and

  (
    g1381_p,
    n4503_lo_p_spl_010,
    g1158_n_spl_0
  );


  or

  (
    g1382_n,
    n4515_lo_n_spl_01,
    g1381_p
  );


  or

  (
    g1383_n,
    g1380_p,
    g1382_n
  );


  and

  (
    g1384_p,
    n3423_lo_p_spl_,
    n4503_lo_n_spl_010
  );


  and

  (
    g1385_p,
    n3435_lo_p_spl_,
    n4503_lo_p_spl_010
  );


  or

  (
    g1386_n,
    n4515_lo_p_spl_01,
    g1385_p
  );


  or

  (
    g1387_n,
    g1384_p,
    g1386_n
  );


  and

  (
    g1388_p,
    n3375_lo_p_spl_001,
    g1387_n
  );


  and

  (
    g1389_p,
    g1383_n,
    g1388_p
  );


  and

  (
    g1390_p,
    n4527_lo_n_spl_0001,
    g1182_n_spl_1
  );


  and

  (
    g1391_p,
    n4527_lo_p_spl_0001,
    g1155_n_spl_1
  );


  or

  (
    g1392_n,
    n4539_lo_n_spl_000,
    g1391_p
  );


  or

  (
    g1393_n,
    g1390_p,
    g1392_n
  );


  and

  (
    g1394_p,
    n3519_lo_p_spl_,
    n4527_lo_n_spl_0001
  );


  and

  (
    g1395_p,
    n3639_lo_p_spl_,
    n4527_lo_p_spl_0001
  );


  or

  (
    g1396_n,
    n4539_lo_p_spl_000,
    g1395_p
  );


  or

  (
    g1397_n,
    g1394_p,
    g1396_n
  );


  and

  (
    g1398_p,
    n3375_lo_p_spl_010,
    g1397_n
  );


  and

  (
    g1399_p,
    g1393_n,
    g1398_p
  );


  or

  (
    g1400_n,
    n4527_lo_p_spl_0010,
    g1200_p_spl_1
  );


  or

  (
    g1401_n,
    n4527_lo_n_spl_0010,
    g1137_p_spl_1
  );


  and

  (
    g1402_p,
    n4539_lo_p_spl_001,
    g1401_n
  );


  and

  (
    g1403_p,
    g1400_n,
    g1402_p
  );


  or

  (
    g1404_n,
    n3471_lo_n_spl_,
    n4527_lo_p_spl_0010
  );


  or

  (
    g1405_n,
    n3591_lo_n_spl_,
    n4527_lo_n_spl_0010
  );


  and

  (
    g1406_p,
    n4539_lo_n_spl_001,
    g1405_n
  );


  and

  (
    g1407_p,
    g1404_n,
    g1406_p
  );


  or

  (
    g1408_n,
    n3375_lo_n_spl_0,
    g1407_p
  );


  or

  (
    g1409_n,
    g1403_p,
    g1408_n
  );


  and

  (
    g1410_p,
    n4527_lo_n_spl_0011,
    g1194_n_spl_1
  );


  and

  (
    g1411_p,
    n4527_lo_p_spl_0011,
    g1164_n_spl_1
  );


  or

  (
    g1412_n,
    n4539_lo_n_spl_001,
    g1411_p
  );


  or

  (
    g1413_n,
    g1410_p,
    g1412_n
  );


  and

  (
    g1414_p,
    n3447_lo_p_spl_,
    n4527_lo_n_spl_0011
  );


  and

  (
    g1415_p,
    n3459_lo_p_spl_,
    n4527_lo_p_spl_0011
  );


  or

  (
    g1416_n,
    n4539_lo_p_spl_001,
    g1415_p
  );


  or

  (
    g1417_n,
    g1414_p,
    g1416_n
  );


  and

  (
    g1418_p,
    n3375_lo_p_spl_010,
    g1417_n
  );


  and

  (
    g1419_p,
    g1413_n,
    g1418_p
  );


  and

  (
    g1420_p,
    n3423_lo_p_spl_,
    n4527_lo_n_spl_010
  );


  and

  (
    g1421_p,
    n3435_lo_p_spl_,
    n4527_lo_p_spl_010
  );


  or

  (
    g1422_n,
    g1420_p,
    g1421_p
  );


  and

  (
    g1423_p,
    n4539_lo_n_spl_01,
    g1422_n
  );


  or

  (
    g1424_n,
    n4527_lo_p_spl_010,
    g1187_n_spl_1
  );


  or

  (
    g1425_n,
    n4527_lo_n_spl_010,
    g1158_n_spl_1
  );


  and

  (
    g1426_p,
    n4539_lo_p_spl_01,
    g1425_n
  );


  and

  (
    g1427_p,
    g1424_n,
    g1426_p
  );


  or

  (
    g1428_n,
    g1423_p,
    g1427_p
  );


  and

  (
    g1429_p,
    n3375_lo_p_spl_011,
    g1428_n
  );


  or

  (
    g1430_n,
    n3351_lo_n,
    n4743_lo_n
  );


  and

  (
    g1431_p,
    n3255_lo_p,
    n4659_lo_n_spl_
  );


  and

  (
    g1432_p,
    n4659_lo_p_spl_,
    n2853_o2_n_spl_0
  );


  or

  (
    g1433_n,
    g1431_p,
    g1432_p
  );


  and

  (
    g1434_p,
    n4647_lo_p,
    g1433_n
  );


  and

  (
    g1435_p,
    n3339_lo_n_spl_,
    n5837_o2_p_spl_0
  );


  or

  (
    g1435_n,
    n3339_lo_p_spl_,
    n5837_o2_n_spl_
  );


  and

  (
    g1436_p,
    n3339_lo_p_spl_,
    n5837_o2_n_spl_
  );


  or

  (
    g1436_n,
    n3339_lo_n_spl_,
    n5837_o2_p_spl_
  );


  and

  (
    g1437_p,
    g1435_n,
    g1436_n
  );


  or

  (
    g1437_n,
    g1435_p,
    g1436_p
  );


  and

  (
    g1438_p,
    n4659_lo_p_spl_,
    g1437_n_spl_
  );


  and

  (
    g1439_p,
    n4659_lo_n_spl_,
    n5782_o2_p
  );


  or

  (
    g1440_n,
    g1438_p,
    g1439_p
  );


  and

  (
    g1441_p,
    n4647_lo_n,
    g1440_n
  );


  or

  (
    g1442_n,
    g1434_p,
    g1441_p
  );


  and

  (
    g1443_p,
    g1430_n,
    g1442_n
  );


  or

  (
    g1444_n,
    n2853_o2_p_spl_1,
    g1437_p
  );


  or

  (
    g1445_n,
    n2853_o2_n_spl_1,
    g1437_n_spl_
  );


  and

  (
    g1446_p,
    g1444_n,
    g1445_n
  );


  and

  (
    g1447_p,
    n2853_o2_n_spl_1,
    n2825_o2_p_spl_100
  );


  and

  (
    g1448_p,
    n3263_o2_p,
    n3261_o2_n
  );


  or

  (
    g1449_n,
    g1447_p,
    g1448_p
  );


  and

  (
    g1450_p,
    n2825_o2_p_spl_100,
    g1249_p_spl_
  );


  or

  (
    g1451_n,
    n3267_o2_p,
    n3268_o2_p
  );


  and

  (
    g1452_p,
    n4719_lo_p_spl_100,
    g1451_n
  );


  or

  (
    g1453_n,
    g1450_p,
    g1452_p
  );


  and

  (
    g1454_p,
    n2825_o2_p_spl_101,
    g1250_p_spl_
  );


  or

  (
    g1455_n,
    n3273_o2_p,
    n3274_o2_p
  );


  and

  (
    g1456_p,
    n4719_lo_p_spl_100,
    g1455_n
  );


  or

  (
    g1457_n,
    g1454_p,
    g1456_p
  );


  and

  (
    g1458_p,
    n2825_o2_p_spl_101,
    n3062_o2_p_spl_
  );


  and

  (
    g1459_p,
    n4719_lo_p_spl_101,
    n3281_o2_p
  );


  or

  (
    g1460_n,
    g1458_p,
    g1459_p
  );


  or

  (
    g1461_n,
    n3795_lo_n_spl_,
    n4467_lo_n_spl_
  );


  or

  (
    g1462_n,
    g1049_n_spl_,
    g1461_n
  );


  or

  (
    g1463_n,
    g1054_n_spl_,
    g1462_n
  );


  or

  (
    g1464_n,
    g1111_n_spl_,
    g1463_n
  );


  or

  (
    g1465_n,
    g1120_n_spl_,
    g1464_n
  );


  or

  (
    g1466_n,
    g1212_n_spl_,
    g1465_n
  );


  or

  (
    g1467_n,
    g1233_n_spl_,
    g1466_n
  );


  and

  (
    g1468_p,
    n2825_o2_p_spl_110,
    n3021_o2_n_spl_
  );


  and

  (
    g1469_p,
    n4719_lo_p_spl_101,
    n3294_o2_p
  );


  or

  (
    g1470_n,
    g1468_p,
    g1469_p
  );


  and

  (
    g1471_p,
    n2825_o2_p_spl_110,
    g1243_p_spl_
  );


  and

  (
    g1472_p,
    n3147_lo_p,
    n4731_lo_n_spl_10
  );


  and

  (
    g1473_p,
    n4731_lo_p_spl_01,
    n2618_o2_n
  );


  or

  (
    g1474_n,
    g1472_p,
    g1473_p
  );


  and

  (
    g1475_p,
    n4719_lo_p_spl_110,
    g1474_n
  );


  or

  (
    g1476_n,
    g1471_p,
    g1475_p
  );


  and

  (
    g1477_p,
    n2825_o2_p_spl_111,
    g1246_p_spl_
  );


  and

  (
    g1478_p,
    n2847_lo_p,
    n4731_lo_n_spl_11
  );


  and

  (
    g1479_p,
    n4731_lo_p_spl_10,
    n2637_o2_n
  );


  or

  (
    g1480_n,
    g1478_p,
    g1479_p
  );


  and

  (
    g1481_p,
    n4719_lo_p_spl_110,
    g1480_n
  );


  or

  (
    g1482_n,
    g1477_p,
    g1481_p
  );


  and

  (
    g1483_p,
    n2825_o2_p_spl_111,
    g1234_n_spl_
  );


  or

  (
    g1484_n,
    n3313_o2_p,
    n3314_o2_p
  );


  and

  (
    g1485_p,
    n4719_lo_p_spl_11,
    g1484_n
  );


  or

  (
    g1486_n,
    g1483_p,
    g1485_p
  );


  and

  (
    g1487_p,
    n3099_lo_p_spl_,
    n4695_lo_n_spl_011
  );


  and

  (
    g1488_p,
    n3111_lo_p_spl_,
    n4695_lo_p_spl_011
  );


  or

  (
    g1489_n,
    g1487_p,
    g1488_p
  );


  and

  (
    g1490_p,
    n4707_lo_n_spl_01,
    g1489_n
  );


  and

  (
    g1491_p,
    n4695_lo_n_spl_011,
    g1470_n_spl_00
  );


  and

  (
    g1492_p,
    n4695_lo_p_spl_011,
    g1449_n_spl_00
  );


  or

  (
    g1493_n,
    g1491_p,
    g1492_p
  );


  and

  (
    g1494_p,
    n4707_lo_p_spl_01,
    g1493_n
  );


  or

  (
    g1495_n,
    g1490_p,
    g1494_p
  );


  and

  (
    g1496_p,
    n4683_lo_n_spl_011,
    g1470_n_spl_00
  );


  and

  (
    g1497_p,
    n4683_lo_p_spl_011,
    g1449_n_spl_00
  );


  or

  (
    g1498_n,
    n4671_lo_n_spl_01,
    g1497_p
  );


  or

  (
    g1499_n,
    g1496_p,
    g1498_n
  );


  or

  (
    g1500_n,
    n3099_lo_p_spl_,
    n4683_lo_p_spl_011
  );


  or

  (
    g1501_n,
    n3111_lo_p_spl_,
    n4683_lo_n_spl_011
  );


  and

  (
    g1502_p,
    g1500_n,
    g1501_n
  );


  or

  (
    g1503_n,
    n4671_lo_p_spl_01,
    g1502_p
  );


  and

  (
    g1504_p,
    g1499_n,
    g1503_n
  );


  or

  (
    g1505_n,
    n2823_lo_p_spl_,
    n4683_lo_p_spl_100
  );


  or

  (
    g1506_n,
    n2811_lo_p_spl_,
    n4683_lo_n_spl_100
  );


  and

  (
    g1507_p,
    g1505_n,
    g1506_n
  );


  or

  (
    g1508_n,
    n4671_lo_p_spl_10,
    g1507_p
  );


  and

  (
    g1509_p,
    n4683_lo_n_spl_100,
    g1476_n_spl_00
  );


  and

  (
    g1510_p,
    n4683_lo_p_spl_100,
    g1453_n_spl_00
  );


  or

  (
    g1511_n,
    n4671_lo_n_spl_10,
    g1510_p
  );


  or

  (
    g1512_n,
    g1509_p,
    g1511_n
  );


  and

  (
    g1513_p,
    g1508_n,
    g1512_n
  );


  or

  (
    g1514_n,
    n3087_lo_p_spl_,
    n4683_lo_p_spl_101
  );


  or

  (
    g1515_n,
    n3075_lo_p_spl_,
    n4683_lo_n_spl_101
  );


  and

  (
    g1516_p,
    g1514_n,
    g1515_n
  );


  or

  (
    g1517_n,
    n4671_lo_p_spl_10,
    g1516_p
  );


  and

  (
    g1518_p,
    n4683_lo_n_spl_101,
    g1482_n_spl_00
  );


  and

  (
    g1519_p,
    n4683_lo_p_spl_101,
    g1457_n_spl_00
  );


  or

  (
    g1520_n,
    n4671_lo_n_spl_10,
    g1519_p
  );


  or

  (
    g1521_n,
    g1518_p,
    g1520_n
  );


  and

  (
    g1522_p,
    g1517_n,
    g1521_n
  );


  or

  (
    g1523_n,
    n2787_lo_p_spl_,
    n4683_lo_p_spl_110
  );


  or

  (
    g1524_n,
    n3039_lo_p_spl_,
    n4683_lo_n_spl_110
  );


  and

  (
    g1525_p,
    g1523_n,
    g1524_n
  );


  or

  (
    g1526_n,
    n4671_lo_p_spl_11,
    g1525_p
  );


  and

  (
    g1527_p,
    n4683_lo_n_spl_110,
    g1486_n_spl_00
  );


  and

  (
    g1528_p,
    n4683_lo_p_spl_110,
    g1460_n_spl_00
  );


  or

  (
    g1529_n,
    n4671_lo_n_spl_11,
    g1528_p
  );


  or

  (
    g1530_n,
    g1527_p,
    g1529_n
  );


  and

  (
    g1531_p,
    g1526_n,
    g1530_n
  );


  or

  (
    g1532_n,
    n2823_lo_p_spl_,
    n4695_lo_p_spl_100
  );


  or

  (
    g1533_n,
    n2811_lo_p_spl_,
    n4695_lo_n_spl_100
  );


  and

  (
    g1534_p,
    g1532_n,
    g1533_n
  );


  or

  (
    g1535_n,
    n4707_lo_p_spl_10,
    g1534_p
  );


  and

  (
    g1536_p,
    n4695_lo_n_spl_100,
    g1476_n_spl_00
  );


  and

  (
    g1537_p,
    n4695_lo_p_spl_100,
    g1453_n_spl_00
  );


  or

  (
    g1538_n,
    n4707_lo_n_spl_10,
    g1537_p
  );


  or

  (
    g1539_n,
    g1536_p,
    g1538_n
  );


  and

  (
    g1540_p,
    g1535_n,
    g1539_n
  );


  or

  (
    g1541_n,
    n3087_lo_p_spl_,
    n4695_lo_p_spl_101
  );


  or

  (
    g1542_n,
    n3075_lo_p_spl_,
    n4695_lo_n_spl_101
  );


  and

  (
    g1543_p,
    g1541_n,
    g1542_n
  );


  or

  (
    g1544_n,
    n4707_lo_p_spl_10,
    g1543_p
  );


  and

  (
    g1545_p,
    n4695_lo_n_spl_101,
    g1482_n_spl_00
  );


  and

  (
    g1546_p,
    n4695_lo_p_spl_101,
    g1457_n_spl_00
  );


  or

  (
    g1547_n,
    n4707_lo_n_spl_10,
    g1546_p
  );


  or

  (
    g1548_n,
    g1545_p,
    g1547_n
  );


  and

  (
    g1549_p,
    g1544_n,
    g1548_n
  );


  or

  (
    g1550_n,
    n2787_lo_p_spl_,
    n4695_lo_p_spl_110
  );


  or

  (
    g1551_n,
    n3039_lo_p_spl_,
    n4695_lo_n_spl_110
  );


  and

  (
    g1552_p,
    g1550_n,
    g1551_n
  );


  or

  (
    g1553_n,
    n4707_lo_p_spl_11,
    g1552_p
  );


  and

  (
    g1554_p,
    n4695_lo_n_spl_110,
    g1486_n_spl_00
  );


  and

  (
    g1555_p,
    n4695_lo_p_spl_110,
    g1460_n_spl_00
  );


  or

  (
    g1556_n,
    n4707_lo_n_spl_11,
    g1555_p
  );


  or

  (
    g1557_n,
    g1554_p,
    g1556_n
  );


  and

  (
    g1558_p,
    g1553_n,
    g1557_n
  );


  and

  (
    g1559_p,
    n4503_lo_n_spl_011,
    g1486_n_spl_0
  );


  and

  (
    g1560_p,
    n4503_lo_p_spl_011,
    g1460_n_spl_0
  );


  or

  (
    g1561_n,
    n4515_lo_n_spl_01,
    g1560_p
  );


  or

  (
    g1562_n,
    g1559_p,
    g1561_n
  );


  and

  (
    g1563_p,
    n3531_lo_p_spl_,
    n4503_lo_n_spl_011
  );


  and

  (
    g1564_p,
    n3651_lo_p_spl_,
    n4503_lo_p_spl_011
  );


  or

  (
    g1565_n,
    n4515_lo_p_spl_01,
    g1564_p
  );


  or

  (
    g1566_n,
    g1563_p,
    g1565_n
  );


  and

  (
    g1567_p,
    n3375_lo_p_spl_011,
    g1566_n
  );


  and

  (
    g1568_p,
    g1562_n,
    g1567_p
  );


  and

  (
    g1569_p,
    n4503_lo_n_spl_100,
    g1482_n_spl_0
  );


  and

  (
    g1570_p,
    n4503_lo_p_spl_100,
    g1457_n_spl_0
  );


  or

  (
    g1571_n,
    n4515_lo_n_spl_10,
    g1570_p
  );


  or

  (
    g1572_n,
    g1569_p,
    g1571_n
  );


  and

  (
    g1573_p,
    n3507_lo_p_spl_,
    n4503_lo_n_spl_100
  );


  and

  (
    g1574_p,
    n3627_lo_p_spl_,
    n4503_lo_p_spl_100
  );


  or

  (
    g1575_n,
    n4515_lo_p_spl_10,
    g1574_p
  );


  or

  (
    g1576_n,
    g1573_p,
    g1575_n
  );


  and

  (
    g1577_p,
    n3375_lo_p_spl_100,
    g1576_n
  );


  and

  (
    g1578_p,
    g1572_n,
    g1577_p
  );


  and

  (
    g1579_p,
    n4503_lo_n_spl_101,
    g1476_n_spl_0
  );


  and

  (
    g1580_p,
    n4503_lo_p_spl_101,
    g1453_n_spl_0
  );


  or

  (
    g1581_n,
    n4515_lo_n_spl_10,
    g1580_p
  );


  or

  (
    g1582_n,
    g1579_p,
    g1581_n
  );


  and

  (
    g1583_p,
    n3495_lo_p_spl_,
    n4503_lo_n_spl_101
  );


  and

  (
    g1584_p,
    n3615_lo_p_spl_,
    n4503_lo_p_spl_101
  );


  or

  (
    g1585_n,
    n4515_lo_p_spl_10,
    g1584_p
  );


  or

  (
    g1586_n,
    g1583_p,
    g1585_n
  );


  and

  (
    g1587_p,
    n3375_lo_p_spl_100,
    g1586_n
  );


  and

  (
    g1588_p,
    g1582_n,
    g1587_p
  );


  and

  (
    g1589_p,
    n3483_lo_p_spl_,
    n4503_lo_n_spl_110
  );


  and

  (
    g1590_p,
    n3603_lo_p_spl_,
    n4503_lo_p_spl_110
  );


  or

  (
    g1591_n,
    g1589_p,
    g1590_p
  );


  and

  (
    g1592_p,
    n4515_lo_n_spl_11,
    g1591_n
  );


  and

  (
    g1593_p,
    n4503_lo_n_spl_110,
    g1470_n_spl_0
  );


  and

  (
    g1594_p,
    n4503_lo_p_spl_110,
    g1449_n_spl_0
  );


  or

  (
    g1595_n,
    g1593_p,
    g1594_p
  );


  and

  (
    g1596_p,
    n4515_lo_p_spl_11,
    g1595_n
  );


  or

  (
    g1597_n,
    g1592_p,
    g1596_p
  );


  and

  (
    g1598_p,
    n3375_lo_p_spl_101,
    g1597_n
  );


  and

  (
    g1599_p,
    n3531_lo_p_spl_,
    n4527_lo_n_spl_011
  );


  and

  (
    g1600_p,
    n3651_lo_p_spl_,
    n4527_lo_p_spl_011
  );


  or

  (
    g1601_n,
    g1599_p,
    g1600_p
  );


  and

  (
    g1602_p,
    n4539_lo_n_spl_01,
    g1601_n
  );


  or

  (
    g1603_n,
    n4527_lo_p_spl_011,
    g1486_n_spl_1
  );


  or

  (
    g1604_n,
    n4527_lo_n_spl_011,
    g1460_n_spl_1
  );


  and

  (
    g1605_p,
    n4539_lo_p_spl_01,
    g1604_n
  );


  and

  (
    g1606_p,
    g1603_n,
    g1605_p
  );


  or

  (
    g1607_n,
    g1602_p,
    g1606_p
  );


  and

  (
    g1608_p,
    n3375_lo_p_spl_101,
    g1607_n
  );


  and

  (
    g1609_p,
    n4527_lo_n_spl_100,
    g1482_n_spl_1
  );


  and

  (
    g1610_p,
    n4527_lo_p_spl_100,
    g1457_n_spl_1
  );


  or

  (
    g1611_n,
    n4539_lo_n_spl_10,
    g1610_p
  );


  or

  (
    g1612_n,
    g1609_p,
    g1611_n
  );


  and

  (
    g1613_p,
    n3507_lo_p_spl_,
    n4527_lo_n_spl_100
  );


  and

  (
    g1614_p,
    n3627_lo_p_spl_,
    n4527_lo_p_spl_100
  );


  or

  (
    g1615_n,
    n4539_lo_p_spl_10,
    g1614_p
  );


  or

  (
    g1616_n,
    g1613_p,
    g1615_n
  );


  and

  (
    g1617_p,
    n3375_lo_p_spl_110,
    g1616_n
  );


  and

  (
    g1618_p,
    g1612_n,
    g1617_p
  );


  and

  (
    g1619_p,
    n4527_lo_n_spl_101,
    g1476_n_spl_1
  );


  and

  (
    g1620_p,
    n4527_lo_p_spl_101,
    g1453_n_spl_1
  );


  or

  (
    g1621_n,
    n4539_lo_n_spl_10,
    g1620_p
  );


  or

  (
    g1622_n,
    g1619_p,
    g1621_n
  );


  and

  (
    g1623_p,
    n3495_lo_p_spl_,
    n4527_lo_n_spl_101
  );


  and

  (
    g1624_p,
    n3615_lo_p_spl_,
    n4527_lo_p_spl_101
  );


  or

  (
    g1625_n,
    n4539_lo_p_spl_10,
    g1624_p
  );


  or

  (
    g1626_n,
    g1623_p,
    g1625_n
  );


  and

  (
    g1627_p,
    n3375_lo_p_spl_110,
    g1626_n
  );


  and

  (
    g1628_p,
    g1622_n,
    g1627_p
  );


  and

  (
    g1629_p,
    n4527_lo_n_spl_110,
    g1470_n_spl_1
  );


  and

  (
    g1630_p,
    n4527_lo_p_spl_110,
    g1449_n_spl_1
  );


  or

  (
    g1631_n,
    n4539_lo_n_spl_11,
    g1630_p
  );


  or

  (
    g1632_n,
    g1629_p,
    g1631_n
  );


  and

  (
    g1633_p,
    n3483_lo_p_spl_,
    n4527_lo_n_spl_110
  );


  and

  (
    g1634_p,
    n3603_lo_p_spl_,
    n4527_lo_p_spl_110
  );


  or

  (
    g1635_n,
    n4539_lo_p_spl_11,
    g1634_p
  );


  or

  (
    g1636_n,
    g1633_p,
    g1635_n
  );


  and

  (
    g1637_p,
    n3375_lo_p_spl_111,
    g1636_n
  );


  and

  (
    g1638_p,
    g1632_n,
    g1637_p
  );


  or

  (
    g1639_n,
    n3517_o2_p,
    n3571_o2_n
  );


  or

  (
    g1640_n,
    n4719_lo_n_spl_1,
    n4731_lo_p_spl_10
  );


  or

  (
    g1641_n,
    n3219_lo_p,
    g1640_n_spl_
  );


  and

  (
    g1642_p,
    g1639_n_spl_,
    g1641_n
  );


  and

  (
    g1643_p,
    n4719_lo_n_spl_1,
    n3661_o2_n
  );


  or

  (
    g1644_n,
    n4731_lo_n_spl_11,
    n3759_o2_p
  );


  or

  (
    g1645_n,
    g1643_p,
    g1644_n
  );


  or

  (
    g1646_n,
    n3195_lo_p,
    g1640_n_spl_
  );


  and

  (
    g1647_p,
    g1645_n_spl_,
    g1646_n
  );


  and

  (
    g1648_p,
    n2883_lo_n_spl_,
    n4683_lo_n_spl_111
  );


  and

  (
    g1649_p,
    n2655_lo_n_spl_,
    n4683_lo_p_spl_111
  );


  or

  (
    g1650_n,
    g1648_p,
    g1649_p
  );


  and

  (
    g1651_p,
    n4671_lo_n_spl_11,
    g1650_n
  );


  or

  (
    g1652_n,
    n3063_lo_n,
    n4731_lo_p_spl_11
  );


  and

  (
    g1653_p,
    g1645_n_spl_,
    g1652_n
  );


  or

  (
    g1654_n,
    n4683_lo_p_spl_111,
    g1653_p_spl_0
  );


  or

  (
    g1655_n,
    n3051_lo_n,
    n4731_lo_p_spl_11
  );


  and

  (
    g1656_p,
    g1639_n_spl_,
    g1655_n
  );


  or

  (
    g1657_n,
    n4683_lo_n_spl_111,
    g1656_p_spl_0
  );


  and

  (
    g1658_p,
    n4671_lo_p_spl_11,
    g1657_n
  );


  and

  (
    g1659_p,
    g1654_n,
    g1658_p
  );


  or

  (
    g1660_n,
    g1651_p,
    g1659_p
  );


  and

  (
    g1661_p,
    n2883_lo_n_spl_,
    n4695_lo_n_spl_111
  );


  and

  (
    g1662_p,
    n2655_lo_n_spl_,
    n4695_lo_p_spl_111
  );


  or

  (
    g1663_n,
    g1661_p,
    g1662_p
  );


  and

  (
    g1664_p,
    n4707_lo_n_spl_11,
    g1663_n
  );


  or

  (
    g1665_n,
    n4695_lo_p_spl_111,
    g1653_p_spl_0
  );


  or

  (
    g1666_n,
    n4695_lo_n_spl_111,
    g1656_p_spl_0
  );


  and

  (
    g1667_p,
    n4707_lo_p_spl_11,
    g1666_n
  );


  and

  (
    g1668_p,
    g1665_n,
    g1667_p
  );


  or

  (
    g1669_n,
    g1664_p,
    g1668_p
  );


  or

  (
    g1670_n,
    n4503_lo_p_spl_111,
    g1653_p_spl_1
  );


  or

  (
    g1671_n,
    n4503_lo_n_spl_111,
    g1656_p_spl_1
  );


  and

  (
    g1672_p,
    n4515_lo_p_spl_11,
    g1671_n
  );


  and

  (
    g1673_p,
    g1670_n,
    g1672_p
  );


  or

  (
    g1674_n,
    n3555_lo_n_spl_,
    n4503_lo_p_spl_111
  );


  or

  (
    g1675_n,
    n3543_lo_n_spl_,
    n4503_lo_n_spl_111
  );


  and

  (
    g1676_p,
    n4515_lo_n_spl_11,
    g1675_n
  );


  and

  (
    g1677_p,
    g1674_n,
    g1676_p
  );


  or

  (
    g1678_n,
    n3375_lo_n_spl_1,
    g1677_p
  );


  or

  (
    g1679_n,
    g1673_p,
    g1678_n
  );


  or

  (
    g1680_n,
    n3555_lo_n_spl_,
    n4527_lo_p_spl_111
  );


  or

  (
    g1681_n,
    n3543_lo_n_spl_,
    n4527_lo_n_spl_111
  );


  and

  (
    g1682_p,
    g1680_n,
    g1681_n
  );


  or

  (
    g1683_n,
    n4539_lo_p_spl_11,
    g1682_p
  );


  and

  (
    g1684_p,
    n4527_lo_n_spl_111,
    g1653_p_spl_1
  );


  and

  (
    g1685_p,
    n4527_lo_p_spl_111,
    g1656_p_spl_1
  );


  or

  (
    g1686_n,
    n4539_lo_n_spl_11,
    g1685_p
  );


  or

  (
    g1687_n,
    g1684_p,
    g1686_n
  );


  and

  (
    g1688_p,
    g1683_n,
    g1687_n
  );


  or

  (
    g1689_n,
    n3375_lo_n_spl_1,
    g1688_p
  );


  and

  (
    g1690_p,
    n2134_inv_n_spl_0,
    n2718_o2_n_spl_
  );


  or

  (
    g1690_n,
    n2134_inv_p_spl_0,
    n2718_o2_p_spl_0
  );


  and

  (
    g1691_p,
    n2134_inv_p_spl_0,
    n2718_o2_p_spl_0
  );


  or

  (
    g1691_n,
    n2134_inv_n_spl_0,
    n2718_o2_n_spl_
  );


  and

  (
    g1692_p,
    g1690_n_spl_,
    g1691_n
  );


  or

  (
    g1692_n,
    g1690_p,
    g1691_p
  );


  or

  (
    g1693_n,
    n5663_o2_n_spl_00,
    n2753_o2_n_spl_
  );


  and

  (
    g1694_p,
    n2628_lo_p_spl_0,
    n5892_o2_p
  );


  or

  (
    g1695_n,
    n5773_o2_p,
    g1694_p
  );


  and

  (
    g1696_p,
    n5802_o2_p_spl_,
    g1695_n_spl_
  );


  and

  (
    g1697_p,
    n2660_o2_n,
    n2817_o2_n
  );


  or

  (
    g1697_n,
    n2660_o2_p,
    n2817_o2_p
  );


  and

  (
    g1698_p,
    n2709_o2_n,
    n2715_o2_n_spl_
  );


  or

  (
    g1698_n,
    n2709_o2_p,
    n2715_o2_p_spl_0
  );


  and

  (
    g1699_p,
    n2719_o2_n,
    n2720_o2_n
  );


  or

  (
    g1699_n,
    n2719_o2_p,
    n2720_o2_p
  );


  and

  (
    g1700_p,
    n2723_o2_n,
    n2724_o2_n
  );


  or

  (
    g1700_n,
    n2723_o2_p,
    n2724_o2_p
  );


  and

  (
    g1701_p,
    n3015_o2_n,
    n3010_o2_n_spl_
  );


  or

  (
    g1701_n,
    n3015_o2_p,
    n3010_o2_p_spl_
  );


  and

  (
    g1702_p,
    n3010_o2_n_spl_,
    n3012_o2_n
  );


  or

  (
    g1702_n,
    n3010_o2_p_spl_,
    n3012_o2_p
  );


  and

  (
    g1703_p,
    n2653_o2_n,
    n2654_o2_p
  );


  or

  (
    g1703_n,
    n2653_o2_p_spl_,
    n2654_o2_n
  );


  and

  (
    g1704_p,
    n2740_o2_p_spl_0,
    n2736_o2_p_spl_
  );


  or

  (
    g1704_n,
    n2740_o2_n_spl_,
    n2736_o2_n
  );


  and

  (
    g1705_p,
    n2614_inv_p_spl_0,
    g1703_p_spl_0
  );


  or

  (
    g1705_n,
    n2614_inv_n_spl_,
    g1703_n_spl_
  );


  and

  (
    g1706_p,
    n4632_lo_n_spl_000,
    n5796_o2_p
  );


  and

  (
    g1707_p,
    n4596_lo_p_spl_000,
    n5796_o2_n
  );


  or

  (
    g1708_n,
    g1706_p,
    g1707_p
  );


  and

  (
    g1709_p,
    n5914_o2_p_spl_0,
    lo382_buf_o2_p_spl_00
  );


  or

  (
    g1709_n,
    n5914_o2_n_spl_,
    lo382_buf_o2_n_spl_00
  );


  and

  (
    g1710_p,
    n5914_o2_n_spl_,
    lo386_buf_o2_p
  );


  or

  (
    g1710_n,
    n5914_o2_p_spl_0,
    lo386_buf_o2_n
  );


  and

  (
    g1711_p,
    g1709_n,
    g1710_n
  );


  or

  (
    g1711_n,
    g1709_p,
    g1710_p
  );


  and

  (
    g1712_p,
    n2353_inv_n,
    n2629_inv_p_spl_
  );


  or

  (
    g1712_n,
    n2353_inv_p_spl_,
    n2629_inv_n
  );


  and

  (
    g1713_p,
    n2735_o2_p,
    g1698_n_spl_0
  );


  or

  (
    g1713_n,
    n2735_o2_n,
    g1698_p_spl_0
  );


  and

  (
    g1714_p,
    n2734_o2_n_spl_,
    g1713_n
  );


  or

  (
    g1714_n,
    n2734_o2_p_spl_,
    g1713_p
  );


  and

  (
    g1715_p,
    n2689_inv_p_spl_0,
    n2711_o2_n_spl_
  );


  or

  (
    g1715_n,
    n2689_inv_n_spl_0,
    n2711_o2_p_spl_
  );


  and

  (
    g1716_p,
    n2715_o2_n_spl_,
    g1715_n
  );


  or

  (
    g1716_n,
    n2715_o2_p_spl_0,
    g1715_p
  );


  and

  (
    g1717_p,
    lo585_buf_o2_p_spl_00,
    g1700_n_spl_0
  );


  or

  (
    g1717_n,
    lo585_buf_o2_n_spl_0,
    g1700_p_spl_
  );


  and

  (
    g1718_p,
    lo585_buf_o2_n_spl_0,
    g1700_p_spl_
  );


  or

  (
    g1718_n,
    lo585_buf_o2_p_spl_00,
    g1700_n_spl_0
  );


  and

  (
    g1719_p,
    g1717_n_spl_,
    g1718_n
  );


  or

  (
    g1719_n,
    g1717_p_spl_,
    g1718_p
  );


  and

  (
    g1720_p,
    n2657_o2_n,
    n2658_o2_n
  );


  or

  (
    g1720_n,
    n2657_o2_p,
    n2658_o2_p
  );


  and

  (
    g1721_p,
    n2663_o2_n,
    n2664_o2_n
  );


  or

  (
    g1721_n,
    n2663_o2_p,
    n2664_o2_p
  );


  and

  (
    g1722_p,
    n2684_o2_n,
    n2685_o2_n
  );


  or

  (
    g1722_n,
    n2684_o2_p,
    n2685_o2_p
  );


  or

  (
    g1723_n,
    n5657_o2_p,
    g1696_p_spl_
  );


  and

  (
    g1724_p,
    n5919_o2_p_spl_,
    g1723_n_spl_
  );


  and

  (
    g1725_p,
    n2611_inv_p_spl_0,
    n2682_o2_p_spl_0
  );


  or

  (
    g1725_n,
    n2611_inv_n_spl_,
    n2682_o2_n_spl_
  );


  and

  (
    g1726_p,
    n2856_lo_p,
    n5849_o2_p_spl_0
  );


  and

  (
    g1727_p,
    n2856_lo_n,
    n5849_o2_n
  );


  or

  (
    g1728_n,
    g1726_p,
    g1727_p
  );


  and

  (
    g1729_p,
    n4632_lo_n_spl_000,
    n5598_o2_n_spl_0
  );


  and

  (
    g1730_p,
    n4620_lo_n_spl_000,
    n5598_o2_p_spl_0
  );


  or

  (
    g1731_n,
    g1729_p,
    g1730_p
  );


  and

  (
    g1732_p,
    n5795_o2_p,
    g1731_n
  );


  and

  (
    g1733_p,
    n4608_lo_p_spl_000,
    n5598_o2_p_spl_0
  );


  and

  (
    g1734_p,
    n4596_lo_p_spl_000,
    n5598_o2_n_spl_0
  );


  or

  (
    g1735_n,
    g1733_p,
    g1734_p
  );


  and

  (
    g1736_p,
    n5795_o2_n,
    g1735_n
  );


  or

  (
    g1737_n,
    g1732_p,
    g1736_p
  );


  and

  (
    g1738_p,
    n4632_lo_n_spl_001,
    n5325_o2_n_spl_0
  );


  and

  (
    g1739_p,
    n4620_lo_n_spl_000,
    n5325_o2_p_spl_0
  );


  or

  (
    g1740_n,
    g1738_p,
    g1739_p
  );


  and

  (
    g1741_p,
    n5407_o2_p,
    g1740_n
  );


  and

  (
    g1742_p,
    n4608_lo_p_spl_000,
    n5325_o2_p_spl_0
  );


  and

  (
    g1743_p,
    n4596_lo_p_spl_001,
    n5325_o2_n_spl_0
  );


  or

  (
    g1744_n,
    g1742_p,
    g1743_p
  );


  and

  (
    g1745_p,
    n5407_o2_n,
    g1744_n
  );


  or

  (
    g1746_n,
    g1741_p,
    g1745_p
  );


  and

  (
    g1747_p,
    n4632_lo_n_spl_001,
    n5833_o2_n_spl_0
  );


  and

  (
    g1748_p,
    n4620_lo_n_spl_001,
    n5833_o2_p_spl_0
  );


  or

  (
    g1749_n,
    g1747_p,
    g1748_p
  );


  and

  (
    g1750_p,
    lo586_buf_o2_p,
    g1749_n
  );


  and

  (
    g1751_p,
    n4608_lo_p_spl_001,
    n5833_o2_p_spl_0
  );


  and

  (
    g1752_p,
    n4596_lo_p_spl_001,
    n5833_o2_n_spl_0
  );


  or

  (
    g1753_n,
    g1751_p,
    g1752_p
  );


  and

  (
    g1754_p,
    lo586_buf_o2_n,
    g1753_n
  );


  or

  (
    g1755_n,
    g1750_p,
    g1754_p
  );


  and

  (
    g1756_p,
    n4293_lo_p_spl_00,
    g1711_n_spl_0
  );


  or

  (
    g1756_n,
    n4293_lo_n_spl_0,
    g1711_p_spl_
  );


  and

  (
    g1757_p,
    n4293_lo_n_spl_0,
    g1711_p_spl_
  );


  or

  (
    g1757_n,
    n4293_lo_p_spl_00,
    g1711_n_spl_0
  );


  and

  (
    g1758_p,
    g1756_n,
    g1757_n
  );


  or

  (
    g1758_n,
    g1756_p_spl_,
    g1757_p
  );


  and

  (
    g1759_p,
    lo494_buf_o2_p_spl_000,
    lo434_buf_o2_p_spl_
  );


  or

  (
    g1759_n,
    lo494_buf_o2_n_spl_000,
    lo434_buf_o2_n
  );


  and

  (
    g1760_p,
    lo494_buf_o2_n_spl_000,
    lo438_buf_o2_p
  );


  or

  (
    g1760_n,
    lo494_buf_o2_p_spl_000,
    lo438_buf_o2_n
  );


  and

  (
    g1761_p,
    g1759_n,
    g1760_n
  );


  or

  (
    g1761_n,
    g1759_p,
    g1760_p
  );


  and

  (
    g1762_p,
    lo557_buf_o2_p_spl_0,
    g1721_n_spl_0
  );


  or

  (
    g1762_n,
    lo557_buf_o2_n,
    g1721_p
  );


  or

  (
    g1763_n,
    lo557_buf_o2_p_spl_0,
    g1721_n_spl_0
  );


  and

  (
    g1764_p,
    lo573_buf_o2_p_spl_0,
    g1720_n_spl_0
  );


  or

  (
    g1764_n,
    lo573_buf_o2_n,
    g1720_p
  );


  and

  (
    g1765_p,
    lo466_buf_o2_p_spl_,
    lo490_buf_o2_p_spl_000
  );


  or

  (
    g1765_n,
    lo466_buf_o2_n,
    lo490_buf_o2_n_spl_000
  );


  and

  (
    g1766_p,
    lo470_buf_o2_p,
    lo490_buf_o2_n_spl_000
  );


  or

  (
    g1766_n,
    lo470_buf_o2_n,
    lo490_buf_o2_p_spl_000
  );


  and

  (
    g1767_p,
    g1765_n,
    g1766_n
  );


  or

  (
    g1767_n,
    g1765_p,
    g1766_p
  );


  or

  (
    g1768_n,
    n2611_inv_p_spl_0,
    n2682_o2_p_spl_0
  );


  and

  (
    g1769_p,
    g1698_n_spl_0,
    g1704_p_spl_
  );


  or

  (
    g1769_n,
    g1698_p_spl_0,
    g1704_n
  );


  and

  (
    g1770_p,
    n2734_o2_p_spl_,
    n2740_o2_p_spl_0
  );


  or

  (
    g1770_n,
    n2734_o2_n_spl_,
    n2740_o2_n_spl_
  );


  and

  (
    g1771_p,
    n2738_o2_n,
    g1770_n
  );


  or

  (
    g1771_n,
    n2738_o2_p,
    g1770_p
  );


  and

  (
    g1772_p,
    g1769_n,
    g1771_p
  );


  or

  (
    g1772_n,
    g1769_p,
    g1771_n
  );


  and

  (
    g1773_p,
    g1719_p_spl_0,
    g1772_n_spl_
  );


  or

  (
    g1773_n,
    g1719_n_spl_,
    g1772_p_spl_
  );


  and

  (
    g1774_p,
    g1717_n_spl_,
    g1773_n_spl_
  );


  or

  (
    g1774_n,
    g1717_p_spl_,
    g1773_p_spl_
  );


  and

  (
    g1775_p,
    lo494_buf_o2_p_spl_001,
    lo357_buf_o2_p_spl_
  );


  or

  (
    g1775_n,
    lo494_buf_o2_n_spl_00,
    lo357_buf_o2_n
  );


  and

  (
    g1776_p,
    lo494_buf_o2_n_spl_01,
    lo361_buf_o2_p
  );


  or

  (
    g1776_n,
    lo494_buf_o2_p_spl_001,
    lo361_buf_o2_n
  );


  and

  (
    g1777_p,
    g1775_n,
    g1776_n
  );


  or

  (
    g1777_n,
    g1775_p,
    g1776_p
  );


  and

  (
    g1778_p,
    lo494_buf_o2_p_spl_01,
    lo417_buf_o2_p_spl_
  );


  or

  (
    g1778_n,
    lo494_buf_o2_n_spl_01,
    lo417_buf_o2_n
  );


  and

  (
    g1779_p,
    lo494_buf_o2_n_spl_10,
    lo421_buf_o2_p
  );


  or

  (
    g1779_n,
    lo494_buf_o2_p_spl_01,
    lo421_buf_o2_n
  );


  and

  (
    g1780_p,
    g1778_n,
    g1779_n
  );


  or

  (
    g1780_n,
    g1778_p,
    g1779_p
  );


  and

  (
    g1781_p,
    n3491_o2_n,
    n3492_o2_p
  );


  or

  (
    g1781_n,
    n3491_o2_p,
    n3492_o2_n
  );


  and

  (
    g1782_p,
    g1699_p_spl_0,
    g1781_p_spl_
  );


  or

  (
    g1782_n,
    g1699_n_spl_0,
    g1781_n_spl_
  );


  and

  (
    g1783_p,
    g1699_n_spl_0,
    g1781_n_spl_
  );


  or

  (
    g1783_n,
    g1699_p_spl_0,
    g1781_p_spl_
  );


  and

  (
    g1784_p,
    g1782_n,
    g1783_n
  );


  or

  (
    g1784_n,
    g1782_p,
    g1783_p
  );


  and

  (
    g1785_p,
    g1712_n,
    g1784_p
  );


  and

  (
    g1786_p,
    g1712_p_spl_0,
    g1784_n
  );


  or

  (
    g1787_n,
    g1785_p_spl_,
    g1786_p
  );


  and

  (
    g1788_p,
    lo473_buf_o2_p_spl_,
    lo490_buf_o2_p_spl_001
  );


  and

  (
    g1789_p,
    lo477_buf_o2_p,
    lo490_buf_o2_n_spl_001
  );


  or

  (
    g1790_n,
    g1788_p,
    g1789_p
  );


  and

  (
    g1791_p,
    g1719_n_spl_,
    g1772_p_spl_
  );


  or

  (
    g1791_n,
    g1719_p_spl_0,
    g1772_n_spl_
  );


  and

  (
    g1792_p,
    g1773_n_spl_,
    g1791_n
  );


  or

  (
    g1792_n,
    g1773_p_spl_,
    g1791_p
  );


  and

  (
    g1793_p,
    lo536_buf_o2_p_spl_0,
    g1761_n_spl_0
  );


  or

  (
    g1793_n,
    lo536_buf_o2_n,
    g1761_p
  );


  and

  (
    g1794_p,
    lo553_buf_o2_p_spl_0,
    g1722_n_spl_0
  );


  or

  (
    g1794_n,
    lo553_buf_o2_n,
    g1722_p
  );


  or

  (
    g1795_n,
    lo553_buf_o2_p_spl_0,
    g1722_n_spl_0
  );


  and

  (
    g1796_p,
    g1794_n,
    g1795_n
  );


  and

  (
    g1797_p,
    g1762_n,
    g1763_n_spl_0
  );


  or

  (
    g1798_n,
    lo573_buf_o2_p_spl_0,
    g1720_n_spl_0
  );


  and

  (
    g1799_p,
    g1764_n,
    g1798_n
  );


  and

  (
    g1800_p,
    lo508_buf_o2_p_spl_,
    lo490_buf_o2_p_spl_001
  );


  or

  (
    g1800_n,
    lo508_buf_o2_n,
    lo490_buf_o2_n_spl_001
  );


  and

  (
    g1801_p,
    lo512_buf_o2_p_spl_,
    lo490_buf_o2_n_spl_010
  );


  or

  (
    g1801_n,
    lo512_buf_o2_n,
    lo490_buf_o2_p_spl_010
  );


  and

  (
    g1802_p,
    g1800_n,
    g1801_n
  );


  or

  (
    g1802_n,
    g1800_p,
    g1801_p
  );


  and

  (
    g1803_p,
    n4254_lo_p_spl_0,
    g1780_n_spl_0
  );


  or

  (
    g1803_n,
    n4254_lo_n,
    g1780_p
  );


  and

  (
    g1804_p,
    n4314_lo_p_spl_0,
    g1777_n_spl_0
  );


  or

  (
    g1804_n,
    n4314_lo_n,
    g1777_p
  );


  and

  (
    g1805_p,
    n4350_lo_p_spl_0,
    g1790_n_spl_0
  );


  and

  (
    g1806_p,
    lo576_buf_o2_p_spl_0,
    g1767_n_spl_0
  );


  or

  (
    g1806_n,
    lo576_buf_o2_n,
    g1767_p
  );


  or

  (
    g1807_n,
    lo576_buf_o2_p_spl_0,
    g1767_n_spl_0
  );


  and

  (
    g1808_p,
    g1806_n,
    g1807_n_spl_
  );


  and

  (
    g1809_p,
    g1797_p_spl_,
    g1799_p_spl_0
  );


  and

  (
    g1810_p,
    n2832_lo_p,
    n4728_lo_n_spl_000
  );


  and

  (
    g1811_p,
    n3132_lo_p,
    n4728_lo_n_spl_000
  );


  and

  (
    g1812_p,
    n3168_lo_p,
    n4728_lo_n_spl_001
  );


  or

  (
    g1813_n,
    n3180_lo_p,
    n4728_lo_p_spl_000
  );


  or

  (
    g1814_n,
    n3204_lo_p,
    n4728_lo_p_spl_000
  );


  and

  (
    g1815_p,
    n3228_lo_p,
    n4728_lo_n_spl_001
  );


  and

  (
    g1816_p,
    n3288_lo_p,
    n4728_lo_n_spl_010
  );


  or

  (
    g1817_n,
    n3300_lo_p,
    n4728_lo_p_spl_001
  );


  or

  (
    g1818_n,
    n3324_lo_p,
    n4728_lo_p_spl_001
  );


  and

  (
    g1819_p,
    n4632_lo_n_spl_010,
    n5327_o2_n_spl_0
  );


  and

  (
    g1820_p,
    n4620_lo_n_spl_001,
    n5327_o2_p_spl_0
  );


  or

  (
    g1821_n,
    g1819_p,
    g1820_p
  );


  and

  (
    g1822_p,
    n5406_o2_p,
    g1821_n
  );


  and

  (
    g1823_p,
    n4608_lo_p_spl_001,
    n5327_o2_p_spl_0
  );


  and

  (
    g1824_p,
    n4596_lo_p_spl_010,
    n5327_o2_n_spl_0
  );


  or

  (
    g1825_n,
    g1823_p,
    g1824_p
  );


  and

  (
    g1826_p,
    n5406_o2_n,
    g1825_n
  );


  and

  (
    g1827_p,
    n4716_lo_n_spl_0,
    n4728_lo_p_spl_010
  );


  or

  (
    g1828_n,
    n3252_lo_p_spl_,
    n4728_lo_p_spl_010
  );


  and

  (
    g1829_p,
    n4716_lo_p_spl_0,
    g1828_n
  );


  and

  (
    g1830_p,
    n5918_o2_n_spl_,
    n5920_o2_n
  );


  or

  (
    g1830_n,
    n5918_o2_p_spl_,
    n5920_o2_p_spl_0
  );


  and

  (
    g1831_p,
    n2149_inv_n,
    g1830_n
  );


  or

  (
    g1831_n,
    n2149_inv_p_spl_,
    g1830_p
  );


  and

  (
    g1832_p,
    n3478_o2_p_spl_,
    n3484_o2_p_spl_
  );


  or

  (
    g1832_n,
    n3478_o2_n_spl_,
    n3484_o2_n_spl_
  );


  and

  (
    g1833_p,
    n3478_o2_n_spl_,
    n3484_o2_n_spl_
  );


  or

  (
    g1833_n,
    n3478_o2_p_spl_,
    n3484_o2_p_spl_
  );


  and

  (
    g1834_p,
    g1832_n,
    g1833_n
  );


  or

  (
    g1834_n,
    g1832_p,
    g1833_p
  );


  and

  (
    g1835_p,
    g1831_p_spl_,
    g1834_n_spl_
  );


  or

  (
    g1835_n,
    g1831_n_spl_,
    g1834_p_spl_
  );


  and

  (
    g1836_p,
    g1831_n_spl_,
    g1834_p_spl_
  );


  or

  (
    g1836_n,
    g1831_p_spl_,
    g1834_n_spl_
  );


  and

  (
    g1837_p,
    g1835_n,
    g1836_n
  );


  or

  (
    g1837_n,
    g1835_p,
    g1836_p
  );


  and

  (
    g1838_p,
    n5663_o2_p_spl_,
    n3499_o2_p
  );


  or

  (
    g1838_n,
    n5663_o2_n_spl_00,
    n3499_o2_n
  );


  and

  (
    g1839_p,
    n5663_o2_n_spl_0,
    n3508_o2_n
  );


  or

  (
    g1839_n,
    n5663_o2_p_spl_,
    n3508_o2_p
  );


  and

  (
    g1840_p,
    g1838_n,
    g1839_n
  );


  or

  (
    g1840_n,
    g1838_p,
    g1839_p
  );


  and

  (
    g1841_p,
    g1692_p_spl_0,
    g1840_n_spl_
  );


  or

  (
    g1841_n,
    g1692_n_spl_0,
    g1840_p_spl_
  );


  and

  (
    g1842_p,
    g1692_n_spl_0,
    g1840_p_spl_
  );


  or

  (
    g1842_n,
    g1692_p_spl_0,
    g1840_n_spl_
  );


  and

  (
    g1843_p,
    g1841_n,
    g1842_n
  );


  or

  (
    g1843_n,
    g1841_p,
    g1842_p
  );


  and

  (
    g1844_p,
    g1837_n,
    g1843_p
  );


  and

  (
    g1845_p,
    g1837_p,
    g1843_n
  );


  or

  (
    g1846_n,
    g1844_p,
    g1845_p
  );


  and

  (
    g1847_p,
    n4716_lo_n_spl_0,
    g1846_n
  );


  or

  (
    g1848_n,
    n4728_lo_n_spl_010,
    g1755_n_spl_
  );


  or

  (
    g1849_n,
    n4728_lo_n_spl_01,
    g1737_n_spl_
  );


  and

  (
    g1850_p,
    n4728_lo_p_spl_011,
    n2492_o2_n
  );


  and

  (
    g1851_p,
    n4728_lo_p_spl_011,
    n2505_o2_p
  );


  and

  (
    g1852_p,
    n4728_lo_p_spl_100,
    n2514_o2_n
  );


  or

  (
    g1853_n,
    n4728_lo_n_spl_10,
    g1746_n_spl_
  );


  and

  (
    g1854_p,
    n3536_o2_n,
    n3537_o2_n
  );


  or

  (
    g1854_n,
    n3536_o2_p,
    n3537_o2_p
  );


  and

  (
    g1855_p,
    n3554_o2_n,
    n3555_o2_n
  );


  or

  (
    g1855_n,
    n3554_o2_p,
    n3555_o2_p
  );


  and

  (
    g1856_p,
    g1854_p_spl_,
    g1855_n_spl_
  );


  or

  (
    g1856_n,
    g1854_n_spl_,
    g1855_p_spl_
  );


  and

  (
    g1857_p,
    g1854_n_spl_,
    g1855_p_spl_
  );


  or

  (
    g1857_n,
    g1854_p_spl_,
    g1855_n_spl_
  );


  and

  (
    g1858_p,
    g1856_n,
    g1857_n
  );


  or

  (
    g1858_n,
    g1856_p,
    g1857_p
  );


  and

  (
    g1859_p,
    n2502_o2_n,
    n3560_o2_p
  );


  or

  (
    g1859_n,
    n2502_o2_p_spl_,
    n3560_o2_n
  );


  and

  (
    g1860_p,
    n2704_inv_n,
    n3562_o2_n
  );


  or

  (
    g1860_n,
    n2704_inv_p_spl_,
    n3562_o2_p
  );


  and

  (
    g1861_p,
    g1859_p_spl_,
    g1860_p_spl_
  );


  or

  (
    g1861_n,
    g1859_n_spl_,
    g1860_n_spl_
  );


  and

  (
    g1862_p,
    g1859_n_spl_,
    g1860_n_spl_
  );


  or

  (
    g1862_n,
    g1859_p_spl_,
    g1860_p_spl_
  );


  and

  (
    g1863_p,
    g1861_n,
    g1862_n
  );


  or

  (
    g1863_n,
    g1861_p,
    g1862_p
  );


  and

  (
    g1864_p,
    g1858_p,
    g1863_p
  );


  and

  (
    g1865_p,
    g1858_n,
    g1863_n
  );


  or

  (
    g1866_n,
    n4716_lo_n_spl_,
    g1865_p
  );


  or

  (
    g1867_n,
    g1864_p,
    g1866_n
  );


  and

  (
    g1868_p,
    n4728_lo_p_spl_100,
    g1867_n
  );


  and

  (
    g1869_p,
    n5568_o2_n,
    n5635_o2_p
  );


  and

  (
    g1870_p,
    n5568_o2_p,
    n5635_o2_n
  );


  and

  (
    g1871_p,
    n2628_lo_p_spl_0,
    n2620_inv_p_spl_0
  );


  or

  (
    g1871_n,
    n2628_lo_n_spl_,
    n2620_inv_n_spl_0
  );


  and

  (
    g1872_p,
    n2617_inv_n_spl_0,
    g1871_n
  );


  or

  (
    g1872_n,
    n2617_inv_p_spl_00,
    g1871_p
  );


  and

  (
    g1873_p,
    n5641_o2_n,
    g1872_n_spl_00
  );


  and

  (
    g1874_p,
    n5641_o2_p,
    g1872_p_spl_00
  );


  and

  (
    g1875_p,
    n5820_o2_p,
    n3048_o2_p_spl_
  );


  and

  (
    g1876_p,
    n5661_o2_n,
    n3048_o2_n_spl_0
  );


  or

  (
    g1877_n,
    g1875_p,
    g1876_p
  );


  or

  (
    g1878_n,
    n5663_o2_n_spl_1,
    g1877_n_spl_
  );


  and

  (
    g1879_p,
    n5663_o2_n_spl_1,
    g1877_n_spl_
  );


  or

  (
    g1880_n,
    n5802_o2_p_spl_,
    g1695_n_spl_
  );


  or

  (
    g1881_n,
    n5869_o2_p,
    g1724_p_spl_
  );


  and

  (
    g1882_p,
    n4188_lo_p_spl_0,
    n5373_o2_p
  );


  and

  (
    g1883_p,
    n4200_lo_p,
    n5373_o2_n
  );


  or

  (
    g1884_n,
    g1882_p,
    g1883_p
  );


  or

  (
    g1885_n,
    n5849_o2_p_spl_0,
    g1884_n_spl_
  );


  and

  (
    g1886_p,
    n5849_o2_p_spl_,
    g1884_n_spl_
  );


  or

  (
    g1887_n,
    n5919_o2_p_spl_,
    g1723_n_spl_
  );


  and

  (
    g1888_p,
    n5920_o2_p_spl_0,
    n2863_o2_p_spl_
  );


  or

  (
    g1889_n,
    n5920_o2_p_spl_,
    n2863_o2_p_spl_
  );


  or

  (
    g1890_n,
    n3048_o2_n_spl_0,
    g1693_n_spl_
  );


  and

  (
    g1891_p,
    n5824_o2_n,
    g1890_n
  );


  and

  (
    g1892_p,
    n2134_inv_n_spl_1,
    g1891_p_spl_
  );


  or

  (
    g1893_n,
    n2134_inv_n_spl_1,
    g1891_p_spl_
  );


  or

  (
    g1894_n,
    g1692_n_spl_,
    g1728_n_spl_
  );


  and

  (
    g1895_p,
    n2628_lo_p_spl_1,
    n5823_o2_p_spl_
  );


  or

  (
    g1895_n,
    n2628_lo_n_spl_,
    n5823_o2_n
  );


  or

  (
    g1896_n,
    n2628_lo_p_spl_1,
    n5823_o2_p_spl_
  );


  and

  (
    g1897_p,
    g1895_n_spl_,
    g1896_n
  );


  and

  (
    g1898_p,
    n4098_lo_n,
    lo490_buf_o2_n_spl_010
  );


  or

  (
    g1898_n,
    n4098_lo_p_spl_,
    lo490_buf_o2_p_spl_010
  );


  and

  (
    g1899_p,
    n3120_lo_p,
    n4728_lo_n_spl_10
  );


  and

  (
    g1900_p,
    n4728_lo_p_spl_101,
    n2501_o2_n
  );


  or

  (
    g1901_n,
    g1899_p,
    g1900_p
  );


  and

  (
    g1902_p,
    n3156_lo_p,
    n4728_lo_n_spl_11
  );


  and

  (
    g1903_p,
    n4728_lo_p_spl_101,
    n2591_o2_n_spl_0
  );


  or

  (
    g1904_n,
    g1902_p,
    g1903_p
  );


  or

  (
    g1905_n,
    n3312_lo_n,
    n4728_lo_p_spl_11
  );


  or

  (
    g1906_n,
    n4728_lo_n_spl_11,
    g1708_n_spl_
  );


  and

  (
    g1907_p,
    g1905_n,
    g1906_n
  );


  or

  (
    g1908_n,
    n5400_o2_p_spl_0,
    n5650_o2_p
  );


  or

  (
    g1909_n,
    n5400_o2_n_spl_0,
    n5650_o2_n
  );


  and

  (
    g1910_p,
    g1908_n,
    g1909_n
  );


  and

  (
    g1911_p,
    n5323_o2_p_spl_0,
    n5325_o2_n_spl_
  );


  and

  (
    g1912_p,
    n5323_o2_n_spl_0,
    n5325_o2_p_spl_
  );


  or

  (
    g1913_n,
    g1911_p,
    g1912_p
  );


  and

  (
    g1914_p,
    n5327_o2_n_spl_,
    n5402_o2_p_spl_0
  );


  and

  (
    g1915_p,
    n5327_o2_p_spl_,
    n5402_o2_n_spl_0
  );


  or

  (
    g1916_n,
    g1914_p,
    g1915_p
  );


  and

  (
    g1917_p,
    n4632_lo_n_spl_010,
    n5369_o2_n_spl_0
  );


  and

  (
    g1918_p,
    n4620_lo_n_spl_010,
    n5369_o2_p_spl_0
  );


  or

  (
    g1919_n,
    g1917_p,
    g1918_p
  );


  and

  (
    g1920_p,
    n5559_o2_p,
    g1919_n
  );


  and

  (
    g1921_p,
    n4608_lo_p_spl_010,
    n5369_o2_p_spl_0
  );


  and

  (
    g1922_p,
    n4596_lo_p_spl_010,
    n5369_o2_n_spl_0
  );


  or

  (
    g1923_n,
    g1921_p,
    g1922_p
  );


  and

  (
    g1924_p,
    n5559_o2_n,
    g1923_n
  );


  or

  (
    g1925_n,
    g1920_p,
    g1924_p
  );


  and

  (
    g1926_p,
    n4632_lo_n_spl_011,
    n5402_o2_n_spl_0
  );


  and

  (
    g1927_p,
    n4620_lo_n_spl_010,
    n5402_o2_p_spl_0
  );


  or

  (
    g1928_n,
    g1926_p,
    g1927_p
  );


  and

  (
    g1929_p,
    n5602_o2_p,
    g1928_n
  );


  and

  (
    g1930_p,
    n4608_lo_p_spl_010,
    n5402_o2_p_spl_
  );


  and

  (
    g1931_p,
    n4596_lo_p_spl_011,
    n5402_o2_n_spl_
  );


  or

  (
    g1932_n,
    g1930_p,
    g1931_p
  );


  and

  (
    g1933_p,
    n5602_o2_n,
    g1932_n
  );


  or

  (
    g1934_n,
    g1929_p,
    g1933_p
  );


  and

  (
    g1935_p,
    n4632_lo_n_spl_011,
    n5896_o2_n_spl_0
  );


  and

  (
    g1936_p,
    n4620_lo_n_spl_01,
    n5896_o2_p_spl_0
  );


  or

  (
    g1937_n,
    g1935_p,
    g1936_p
  );


  and

  (
    g1938_p,
    lo562_buf_o2_p,
    g1937_n
  );


  and

  (
    g1939_p,
    n4608_lo_p_spl_01,
    n5896_o2_p_spl_0
  );


  and

  (
    g1940_p,
    n4596_lo_p_spl_011,
    n5896_o2_n_spl_0
  );


  or

  (
    g1941_n,
    g1939_p,
    g1940_p
  );


  and

  (
    g1942_p,
    lo562_buf_o2_n,
    g1941_n
  );


  or

  (
    g1943_n,
    g1938_p,
    g1942_p
  );


  and

  (
    g1944_p,
    n4632_lo_n_spl_10,
    n5400_o2_n_spl_0
  );


  and

  (
    g1945_p,
    n4620_lo_n_spl_10,
    n5400_o2_p_spl_0
  );


  or

  (
    g1946_n,
    g1944_p,
    g1945_p
  );


  and

  (
    g1947_p,
    n5603_o2_p,
    g1946_n
  );


  and

  (
    g1948_p,
    n4608_lo_p_spl_10,
    n5400_o2_p_spl_
  );


  and

  (
    g1949_p,
    n4596_lo_p_spl_10,
    n5400_o2_n_spl_
  );


  or

  (
    g1950_n,
    g1948_p,
    g1949_p
  );


  and

  (
    g1951_p,
    n5603_o2_n,
    g1950_n
  );


  or

  (
    g1952_n,
    g1947_p,
    g1951_p
  );


  and

  (
    g1953_p,
    n4632_lo_n_spl_10,
    n5323_o2_n_spl_0
  );


  and

  (
    g1954_p,
    n4620_lo_n_spl_10,
    n5323_o2_p_spl_0
  );


  or

  (
    g1955_n,
    g1953_p,
    g1954_p
  );


  and

  (
    g1956_p,
    n5408_o2_p,
    g1955_n
  );


  and

  (
    g1957_p,
    n4608_lo_p_spl_10,
    n5323_o2_p_spl_
  );


  and

  (
    g1958_p,
    n4596_lo_p_spl_10,
    n5323_o2_n_spl_
  );


  or

  (
    g1959_n,
    g1957_p,
    g1958_p
  );


  and

  (
    g1960_p,
    n5408_o2_n,
    g1959_n
  );


  or

  (
    g1961_n,
    g1956_p,
    g1960_p
  );


  and

  (
    g1962_p,
    n4632_lo_n_spl_11,
    n5600_o2_n_spl_0
  );


  and

  (
    g1963_p,
    n4620_lo_n_spl_11,
    n5600_o2_p_spl_0
  );


  or

  (
    g1964_n,
    g1962_p,
    g1963_p
  );


  and

  (
    g1965_p,
    n5797_o2_p,
    g1964_n
  );


  and

  (
    g1966_p,
    n4608_lo_p_spl_11,
    n5600_o2_p_spl_0
  );


  and

  (
    g1967_p,
    n4596_lo_p_spl_11,
    n5600_o2_n_spl_0
  );


  or

  (
    g1968_n,
    g1966_p,
    g1967_p
  );


  and

  (
    g1969_p,
    n5797_o2_n,
    g1968_n
  );


  or

  (
    g1970_n,
    g1965_p,
    g1969_p
  );


  and

  (
    g1971_p,
    n4632_lo_n_spl_11,
    n5557_o2_n_spl_0
  );


  and

  (
    g1972_p,
    n4620_lo_n_spl_11,
    n5557_o2_p_spl_0
  );


  or

  (
    g1973_n,
    g1971_p,
    g1972_p
  );


  and

  (
    g1974_p,
    n5655_o2_p,
    g1973_n
  );


  and

  (
    g1975_p,
    n4608_lo_p_spl_11,
    n5557_o2_p_spl_0
  );


  and

  (
    g1976_p,
    n4596_lo_p_spl_11,
    n5557_o2_n_spl_0
  );


  or

  (
    g1977_n,
    g1975_p,
    g1976_p
  );


  and

  (
    g1978_p,
    n5655_o2_n,
    g1977_n
  );


  or

  (
    g1979_n,
    g1974_p,
    g1978_p
  );


  and

  (
    g1980_p,
    n3671_o2_n_spl_,
    n3680_o2_p_spl_
  );


  or

  (
    g1980_n,
    n3671_o2_p_spl_,
    n3680_o2_n_spl_
  );


  and

  (
    g1981_p,
    n3671_o2_p_spl_,
    n3680_o2_n_spl_
  );


  or

  (
    g1981_n,
    n3671_o2_n_spl_,
    n3680_o2_p_spl_
  );


  and

  (
    g1982_p,
    g1980_n,
    g1981_n
  );


  or

  (
    g1982_n,
    g1980_p,
    g1981_p
  );


  and

  (
    g1983_p,
    n3692_o2_n_spl_,
    n2591_o2_n_spl_0
  );


  or

  (
    g1983_n,
    n3692_o2_p_spl_,
    n2591_o2_p_spl_0
  );


  and

  (
    g1984_p,
    n3692_o2_p_spl_,
    n2591_o2_p_spl_0
  );


  or

  (
    g1984_n,
    n3692_o2_n_spl_,
    n2591_o2_n_spl_
  );


  and

  (
    g1985_p,
    g1983_n,
    g1984_n
  );


  or

  (
    g1985_n,
    g1983_p,
    g1984_p
  );


  and

  (
    g1986_p,
    g1982_n_spl_,
    g1985_p_spl_
  );


  or

  (
    g1986_n,
    g1982_p_spl_,
    g1985_n_spl_
  );


  and

  (
    g1987_p,
    g1982_p_spl_,
    g1985_n_spl_
  );


  or

  (
    g1987_n,
    g1982_n_spl_,
    g1985_p_spl_
  );


  and

  (
    g1988_p,
    g1986_n,
    g1987_n
  );


  or

  (
    g1988_n,
    g1986_p,
    g1987_p
  );


  and

  (
    g1989_p,
    n3707_o2_n_spl_,
    n3716_o2_p_spl_
  );


  or

  (
    g1989_n,
    n3707_o2_p_spl_,
    n3716_o2_n_spl_
  );


  and

  (
    g1990_p,
    n3707_o2_p_spl_,
    n3716_o2_n_spl_
  );


  or

  (
    g1990_n,
    n3707_o2_n_spl_,
    n3716_o2_p_spl_
  );


  and

  (
    g1991_p,
    g1989_n,
    g1990_n
  );


  or

  (
    g1991_n,
    g1989_p,
    g1990_p
  );


  and

  (
    g1992_p,
    n3749_o2_n_spl_,
    n3740_o2_n_spl_
  );


  or

  (
    g1992_n,
    n3749_o2_p_spl_,
    n3740_o2_p_spl_
  );


  and

  (
    g1993_p,
    n3749_o2_p_spl_,
    n3740_o2_p_spl_
  );


  or

  (
    g1993_n,
    n3749_o2_n_spl_,
    n3740_o2_n_spl_
  );


  and

  (
    g1994_p,
    g1992_n,
    g1993_n
  );


  or

  (
    g1994_n,
    g1992_p,
    g1993_p
  );


  and

  (
    g1995_p,
    g1991_p_spl_,
    g1994_n_spl_
  );


  or

  (
    g1995_n,
    g1991_n_spl_,
    g1994_p_spl_
  );


  and

  (
    g1996_p,
    g1991_n_spl_,
    g1994_p_spl_
  );


  or

  (
    g1996_n,
    g1991_p_spl_,
    g1994_n_spl_
  );


  and

  (
    g1997_p,
    g1995_n,
    g1996_n
  );


  or

  (
    g1997_n,
    g1995_p,
    g1996_p
  );


  or

  (
    g1998_n,
    g1988_p,
    g1997_n
  );


  or

  (
    g1999_n,
    g1988_n,
    g1997_p
  );


  and

  (
    g2000_p,
    n4716_lo_p_spl_0,
    g1999_n
  );


  and

  (
    g2001_p,
    g1998_n,
    g2000_p
  );


  and

  (
    g2002_p,
    n5412_o2_n,
    n2700_o2_p
  );


  and

  (
    g2003_p,
    n5412_o2_p,
    n2700_o2_n
  );


  or

  (
    g2004_n,
    g2002_p,
    g2003_p
  );


  or

  (
    g2005_n,
    n5565_o2_n,
    g1872_p_spl_00
  );


  or

  (
    g2006_n,
    n5564_o2_p,
    g1872_n_spl_00
  );


  and

  (
    g2007_p,
    g2005_n,
    g2006_n
  );


  and

  (
    g2008_p,
    n5637_o2_n,
    g1895_n_spl_
  );


  or

  (
    g2008_n,
    n5637_o2_p,
    g1895_p
  );


  or

  (
    g2009_n,
    n5640_o2_p,
    g2008_n
  );


  or

  (
    g2010_n,
    n5640_o2_n,
    g2008_p
  );


  and

  (
    g2011_p,
    g2009_n,
    g2010_n
  );


  and

  (
    g2012_p,
    n3936_lo_p_spl_0,
    n5329_o2_p_spl_
  );


  or

  (
    g2012_n,
    n3936_lo_n_spl_0,
    n5329_o2_n_spl_
  );


  and

  (
    g2013_p,
    n3948_lo_p,
    n5329_o2_n_spl_
  );


  or

  (
    g2013_n,
    n3948_lo_n,
    n5329_o2_p_spl_
  );


  and

  (
    g2014_p,
    g2012_n,
    g2013_n
  );


  or

  (
    g2014_n,
    g2012_p,
    g2013_p
  );


  or

  (
    g2015_n,
    n5848_o2_p,
    g2014_n
  );


  or

  (
    g2016_n,
    n5848_o2_n,
    g2014_p
  );


  and

  (
    g2017_p,
    g2015_n,
    g2016_n
  );


  and

  (
    g2018_p,
    n5856_o2_p,
    g1872_n_spl_0
  );


  and

  (
    g2019_p,
    n2818_o2_p_spl_,
    g1872_p_spl_0
  );


  or

  (
    g2020_n,
    g2018_p,
    g2019_p
  );


  or

  (
    g2021_n,
    n5918_o2_n_spl_,
    n2878_o2_n
  );


  or

  (
    g2022_n,
    n5918_o2_p_spl_,
    n2878_o2_p
  );


  and

  (
    g2023_p,
    g2021_n,
    g2022_n
  );


  and

  (
    g2024_p,
    n3013_o2_p,
    g1872_n_spl_1
  );


  or

  (
    g2024_n,
    n3013_o2_n,
    g1872_p_spl_1
  );


  and

  (
    g2025_p,
    n3016_o2_p,
    g1872_p_spl_1
  );


  or

  (
    g2025_n,
    n3016_o2_n,
    g1872_n_spl_1
  );


  and

  (
    g2026_p,
    g2024_n,
    g2025_n
  );


  or

  (
    g2026_n,
    g2024_p,
    g2025_p
  );


  and

  (
    g2027_p,
    n2655_o2_p_spl_,
    g2026_p
  );


  and

  (
    g2028_p,
    n2655_o2_n,
    g2026_n
  );


  or

  (
    g2029_n,
    g2027_p,
    g2028_p
  );


  and

  (
    g2030_p,
    n2753_o2_n_spl_,
    n3048_o2_p_spl_
  );


  and

  (
    g2031_p,
    n2753_o2_p,
    n3048_o2_n_spl_
  );


  or

  (
    g2032_n,
    g2030_p,
    g2031_p
  );


  and

  (
    g2033_p,
    n5371_o2_p,
    n5404_o2_n
  );


  and

  (
    g2034_p,
    n5371_o2_n,
    n5404_o2_p
  );


  or

  (
    g2035_n,
    g2033_p,
    g2034_p
  );


  or

  (
    g2036_n,
    n5831_o2_p,
    lo450_buf_o2_n
  );


  or

  (
    g2037_n,
    n5831_o2_n,
    lo450_buf_o2_p_spl_
  );


  and

  (
    g2038_p,
    g2036_n,
    g2037_n
  );


  and

  (
    g2039_p,
    g2035_n_spl_,
    g2038_p_spl_
  );


  or

  (
    g2040_n,
    g2035_n_spl_,
    g2038_p_spl_
  );


  and

  (
    g2041_p,
    n4188_lo_n_spl_,
    n5653_o2_p_spl_
  );


  or

  (
    g2041_n,
    n4188_lo_p_spl_0,
    n5653_o2_n_spl_
  );


  and

  (
    g2042_p,
    n4188_lo_p_spl_,
    n5653_o2_n_spl_
  );


  or

  (
    g2042_n,
    n4188_lo_n_spl_,
    n5653_o2_p_spl_
  );


  and

  (
    g2043_p,
    g2041_n,
    g2042_n
  );


  or

  (
    g2043_n,
    g2041_p,
    g2042_p
  );


  and

  (
    g2044_p,
    n5833_o2_p_spl_,
    g2043_p
  );


  and

  (
    g2045_p,
    n5833_o2_n_spl_,
    g2043_n
  );


  or

  (
    g2046_n,
    g2044_p,
    g2045_p
  );


  or

  (
    g2047_n,
    n5557_o2_p_spl_,
    n5600_o2_n_spl_
  );


  or

  (
    g2048_n,
    n5557_o2_n_spl_,
    n5600_o2_p_spl_
  );


  and

  (
    g2049_p,
    g2047_n,
    g2048_n
  );


  and

  (
    g2050_p,
    g2046_n_spl_,
    g2049_p_spl_
  );


  or

  (
    g2051_n,
    g2046_n_spl_,
    g2049_p_spl_
  );


  and

  (
    g2052_p,
    n5739_o2_n,
    n2725_o2_p
  );


  and

  (
    g2053_p,
    n5739_o2_p,
    n2725_o2_n
  );


  or

  (
    g2054_n,
    g2052_p,
    g2053_p
  );


  and

  (
    g2055_p,
    n5656_o2_n,
    n5799_o2_p
  );


  and

  (
    g2056_p,
    n5656_o2_p,
    n5799_o2_n
  );


  or

  (
    g2057_n,
    g2055_p,
    g2056_p
  );


  or

  (
    g2058_n,
    g2054_n_spl_,
    g2057_n_spl_
  );


  and

  (
    g2059_p,
    g2054_n_spl_,
    g2057_n_spl_
  );


  and

  (
    g2060_p,
    n5598_o2_n_spl_1,
    n5896_o2_p_spl_1
  );


  or

  (
    g2060_n,
    n5598_o2_p_spl_1,
    n5896_o2_n_spl_1
  );


  and

  (
    g2061_p,
    n5598_o2_p_spl_1,
    n5896_o2_n_spl_1
  );


  or

  (
    g2061_n,
    n5598_o2_n_spl_1,
    n5896_o2_p_spl_1
  );


  and

  (
    g2062_p,
    g2060_n,
    g2061_n
  );


  or

  (
    g2062_n,
    g2060_p,
    g2061_p
  );


  and

  (
    g2063_p,
    n3936_lo_n_spl_0,
    n5369_o2_p_spl_1
  );


  or

  (
    g2063_n,
    n3936_lo_p_spl_0,
    n5369_o2_n_spl_1
  );


  and

  (
    g2064_p,
    n3936_lo_p_spl_,
    n5369_o2_n_spl_1
  );


  or

  (
    g2064_n,
    n3936_lo_n_spl_,
    n5369_o2_p_spl_1
  );


  and

  (
    g2065_p,
    g2063_n,
    g2064_n
  );


  or

  (
    g2065_n,
    g2063_p,
    g2064_p
  );


  or

  (
    g2066_n,
    g2062_n,
    g2065_n
  );


  or

  (
    g2067_n,
    g2062_p,
    g2065_p
  );


  and

  (
    g2068_p,
    g2066_n,
    g2067_n
  );


  and

  (
    g2069_p,
    n3590_o2_p,
    n3591_o2_n
  );


  or

  (
    g2069_n,
    n3590_o2_n,
    n3591_o2_p
  );


  and

  (
    g2070_p,
    n2683_o2_n,
    n3593_o2_p
  );


  or

  (
    g2070_n,
    n2683_o2_p,
    n3593_o2_n
  );


  and

  (
    g2071_p,
    g2069_p_spl_,
    g2070_n_spl_
  );


  or

  (
    g2071_n,
    g2069_n_spl_,
    g2070_p_spl_
  );


  and

  (
    g2072_p,
    g2069_n_spl_,
    g2070_p_spl_
  );


  or

  (
    g2072_n,
    g2069_p_spl_,
    g2070_n_spl_
  );


  and

  (
    g2073_p,
    g2071_n,
    g2072_n
  );


  or

  (
    g2073_n,
    g2071_p,
    g2072_p
  );


  and

  (
    g2074_p,
    n4488_lo_n_spl_0,
    g2073_n
  );


  or

  (
    g2074_n,
    n4488_lo_p_spl_0,
    g2073_p
  );


  and

  (
    g2075_p,
    n3610_o2_n,
    n3611_o2_p
  );


  or

  (
    g2075_n,
    n3610_o2_p,
    n3611_o2_n
  );


  and

  (
    g2076_p,
    n3616_o2_p,
    n3617_o2_n
  );


  or

  (
    g2076_n,
    n3616_o2_n,
    n3617_o2_p
  );


  and

  (
    g2077_p,
    g2075_p_spl_,
    g2076_p_spl_
  );


  or

  (
    g2077_n,
    g2075_n_spl_,
    g2076_n_spl_
  );


  and

  (
    g2078_p,
    g2075_n_spl_,
    g2076_n_spl_
  );


  or

  (
    g2078_n,
    g2075_p_spl_,
    g2076_p_spl_
  );


  and

  (
    g2079_p,
    g2077_n,
    g2078_n
  );


  or

  (
    g2079_n,
    g2077_p,
    g2078_p
  );


  and

  (
    g2080_p,
    n4488_lo_p_spl_0,
    g2079_p
  );


  or

  (
    g2080_n,
    n4488_lo_n_spl_0,
    g2079_n
  );


  and

  (
    g2081_p,
    g2074_n,
    g2080_n
  );


  or

  (
    g2081_n,
    g2074_p,
    g2080_p
  );


  and

  (
    g2082_p,
    n3638_o2_n,
    n3639_o2_p
  );


  or

  (
    g2082_n,
    n3638_o2_p,
    n3639_o2_n
  );


  and

  (
    g2083_p,
    n2617_inv_n_spl_0,
    n2620_inv_n_spl_0
  );


  or

  (
    g2083_n,
    n2617_inv_p_spl_00,
    n2620_inv_p_spl_0
  );


  and

  (
    g2084_p,
    g2082_n_spl_,
    g2083_n
  );


  or

  (
    g2084_n,
    g2082_p_spl_,
    g2083_p
  );


  and

  (
    g2085_p,
    n2617_inv_n_spl_1,
    n3650_o2_n
  );


  or

  (
    g2085_n,
    n2617_inv_p_spl_0,
    n3650_o2_p
  );


  and

  (
    g2086_p,
    n2620_inv_n_spl_,
    g2085_p_spl_
  );


  or

  (
    g2086_n,
    n2620_inv_p_spl_1,
    g2085_n_spl_
  );


  and

  (
    g2087_p,
    g2084_n,
    g2086_n
  );


  or

  (
    g2087_n,
    g2084_p,
    g2086_p
  );


  and

  (
    g2088_p,
    n4488_lo_p_spl_1,
    g2087_n
  );


  or

  (
    g2088_n,
    n4488_lo_n_spl_1,
    g2087_p
  );


  and

  (
    g2089_p,
    n2617_inv_p_spl_1,
    g2082_n_spl_
  );


  or

  (
    g2089_n,
    n2617_inv_n_spl_1,
    g2082_p_spl_
  );


  and

  (
    g2090_p,
    g2085_n_spl_,
    g2089_n
  );


  or

  (
    g2090_n,
    g2085_p_spl_,
    g2089_p
  );


  and

  (
    g2091_p,
    n4488_lo_n_spl_1,
    g2090_n
  );


  or

  (
    g2091_n,
    n4488_lo_p_spl_1,
    g2090_p
  );


  and

  (
    g2092_p,
    g2088_n,
    g2091_n
  );


  or

  (
    g2092_n,
    g2088_p,
    g2091_p
  );


  or

  (
    g2093_n,
    g2081_p,
    g2092_n
  );


  or

  (
    g2094_n,
    g2081_n,
    g2092_p
  );


  and

  (
    g2095_p,
    g2093_n,
    g2094_n
  );


  or

  (
    g2096_n,
    lo536_buf_o2_p_spl_0,
    g1761_n_spl_0
  );


  and

  (
    g2097_p,
    g1793_p_spl_,
    g1796_p_spl_0
  );


  or

  (
    g2098_n,
    g1794_p,
    g2097_p
  );


  and

  (
    g2099_p,
    g1762_p_spl_,
    g1799_p_spl_0
  );


  and

  (
    g2100_p,
    n5936_o2_n_spl_,
    lo398_buf_o2_n_spl_000
  );


  and

  (
    g2101_p,
    n5936_o2_p_spl_0,
    lo402_buf_o2_n_spl_000
  );


  or

  (
    g2102_n,
    g2100_p,
    g2101_p
  );


  and

  (
    g2103_p,
    lo578_buf_o2_p,
    g2102_n
  );


  and

  (
    g2104_p,
    n5936_o2_p_spl_0,
    lo406_buf_o2_p_spl_000
  );


  and

  (
    g2105_p,
    n5936_o2_n_spl_,
    lo390_buf_o2_p_spl_000
  );


  or

  (
    g2106_n,
    g2104_p,
    g2105_p
  );


  and

  (
    g2107_p,
    lo578_buf_o2_n,
    g2106_n
  );


  or

  (
    g2108_n,
    g2103_p,
    g2107_p
  );


  and

  (
    g2109_p,
    lo474_buf_o2_n_spl_,
    lo398_buf_o2_n_spl_000
  );


  and

  (
    g2110_p,
    lo474_buf_o2_p_spl_0,
    lo402_buf_o2_n_spl_000
  );


  or

  (
    g2111_n,
    g2109_p,
    g2110_p
  );


  and

  (
    g2112_p,
    lo582_buf_o2_p,
    g2111_n
  );


  and

  (
    g2113_p,
    lo474_buf_o2_p_spl_0,
    lo406_buf_o2_p_spl_000
  );


  and

  (
    g2114_p,
    lo474_buf_o2_n_spl_,
    lo390_buf_o2_p_spl_000
  );


  or

  (
    g2115_n,
    g2113_p,
    g2114_p
  );


  and

  (
    g2116_p,
    lo582_buf_o2_n,
    g2115_n
  );


  or

  (
    g2117_n,
    g2112_p,
    g2116_p
  );


  and

  (
    g2118_p,
    lo518_buf_o2_n,
    lo398_buf_o2_n_spl_001
  );


  and

  (
    g2119_p,
    lo518_buf_o2_p_spl_,
    lo402_buf_o2_n_spl_001
  );


  or

  (
    g2120_n,
    g2118_p,
    g2119_p
  );


  and

  (
    g2121_p,
    lo458_buf_o2_n,
    lo398_buf_o2_n_spl_001
  );


  and

  (
    g2122_p,
    lo458_buf_o2_p_spl_,
    lo402_buf_o2_n_spl_001
  );


  or

  (
    g2123_n,
    g2121_p,
    g2122_p
  );


  or

  (
    g2124_n,
    n3957_lo_p_spl_0,
    lo390_buf_o2_p_spl_001
  );


  or

  (
    g2125_n,
    n3957_lo_n,
    lo406_buf_o2_p_spl_001
  );


  and

  (
    g2126_p,
    g2124_n,
    g2125_n
  );


  and

  (
    g2127_p,
    n3834_lo_p_spl_,
    lo494_buf_o2_p_spl_10
  );


  or

  (
    g2127_n,
    n3834_lo_n,
    lo494_buf_o2_n_spl_10
  );


  and

  (
    g2128_p,
    n3846_lo_p,
    lo494_buf_o2_n_spl_11
  );


  or

  (
    g2128_n,
    n3846_lo_n,
    lo494_buf_o2_p_spl_10
  );


  and

  (
    g2129_p,
    g2127_n,
    g2128_n
  );


  or

  (
    g2129_n,
    g2127_p,
    g2128_p
  );


  and

  (
    g2130_p,
    n4110_lo_p_spl_,
    lo490_buf_o2_p_spl_011
  );


  or

  (
    g2130_n,
    n4110_lo_n,
    lo490_buf_o2_n_spl_01
  );


  and

  (
    g2131_p,
    n4122_lo_p_spl_,
    lo490_buf_o2_n_spl_10
  );


  or

  (
    g2131_n,
    n4122_lo_n,
    lo490_buf_o2_p_spl_011
  );


  and

  (
    g2132_p,
    g2130_n,
    g2131_n
  );


  or

  (
    g2132_n,
    g2130_p,
    g2131_p
  );


  or

  (
    g2133_n,
    n4398_lo_n,
    g1802_p
  );


  or

  (
    g2134_n,
    n4254_lo_p_spl_0,
    g1780_n_spl_0
  );


  and

  (
    g2135_p,
    g1803_n,
    g2134_n
  );


  or

  (
    g2136_n,
    n4314_lo_p_spl_0,
    g1777_n_spl_0
  );


  and

  (
    g2137_p,
    g1804_n,
    g2136_n
  );


  and

  (
    g2138_p,
    n2811_o2_p_spl_0,
    n2682_o2_p_spl_1
  );


  or

  (
    g2138_n,
    n2811_o2_n_spl_0,
    n2682_o2_n_spl_
  );


  and

  (
    g2139_p,
    n2740_inv_n,
    g2138_n
  );


  or

  (
    g2139_n,
    n2740_inv_p_spl_,
    g2138_p
  );


  and

  (
    g2140_p,
    g1758_p_spl_0,
    g2139_n_spl_0
  );


  or

  (
    g2141_n,
    g1756_p_spl_,
    g2140_p
  );


  or

  (
    g2142_n,
    n2779_inv_n_spl_0,
    g1725_n_spl_
  );


  or

  (
    g2143_n,
    g1758_n_spl_0,
    g2142_n_spl_
  );


  and

  (
    g2144_p,
    n2317_inv_n_spl_,
    n2811_o2_p_spl_0
  );


  or

  (
    g2144_n,
    n2317_inv_p_spl_0,
    n2811_o2_n_spl_0
  );


  and

  (
    g2145_p,
    n2317_inv_p_spl_0,
    n2811_o2_n_spl_1
  );


  or

  (
    g2145_n,
    n2317_inv_n_spl_,
    n2811_o2_p_spl_1
  );


  and

  (
    g2146_p,
    g2144_n,
    g2145_n
  );


  or

  (
    g2146_n,
    g2144_p,
    g2145_p
  );


  and

  (
    g2147_p,
    n2572_inv_n_spl_0,
    g2146_p_spl_
  );


  or

  (
    g2147_n,
    n2572_inv_p_spl_0,
    g2146_n_spl_
  );


  and

  (
    g2148_p,
    n2572_inv_p_spl_0,
    g2146_n_spl_
  );


  or

  (
    g2148_n,
    n2572_inv_n_spl_0,
    g2146_p_spl_
  );


  and

  (
    g2149_p,
    g2147_n,
    g2148_n
  );


  or

  (
    g2149_n,
    g2147_p,
    g2148_p
  );


  and

  (
    g2150_p,
    n2689_o2_n,
    n2638_inv_n
  );


  or

  (
    g2150_n,
    n2689_o2_p_spl_,
    n2638_inv_p_spl_
  );


  and

  (
    g2151_p,
    n2779_inv_n_spl_0,
    g2150_n
  );


  or

  (
    g2151_n,
    n2779_inv_p_spl_0,
    g2150_p
  );


  and

  (
    g2152_p,
    g2139_p_spl_0,
    g2151_n_spl_0
  );


  or

  (
    g2152_n,
    g2139_n_spl_0,
    g2151_p_spl_0
  );


  and

  (
    g2153_p,
    g2139_n_spl_,
    g2151_p_spl_0
  );


  or

  (
    g2153_n,
    g2139_p_spl_0,
    g2151_n_spl_0
  );


  and

  (
    g2154_p,
    g2152_n,
    g2153_n
  );


  or

  (
    g2154_n,
    g2152_p,
    g2153_p
  );


  and

  (
    g2155_p,
    g2149_n,
    g2154_n
  );


  and

  (
    g2156_p,
    g2149_p,
    g2154_p
  );


  or

  (
    g2157_n,
    g2155_p,
    g2156_p
  );


  and

  (
    g2158_p,
    g1758_n_spl_0,
    g2157_n_spl_
  );


  or

  (
    g2159_n,
    g1758_n_spl_1,
    g2157_n_spl_
  );


  or

  (
    g2160_n,
    n4350_lo_p_spl_0,
    g1790_n_spl_0
  );


  and

  (
    g2161_p,
    n3624_o2_n,
    n3625_o2_p
  );


  or

  (
    g2161_n,
    n3624_o2_p,
    n3625_o2_n
  );


  and

  (
    g2162_p,
    g1702_n_spl_0,
    g2161_p_spl_
  );


  or

  (
    g2162_n,
    g1702_p_spl_,
    g2161_n_spl_
  );


  and

  (
    g2163_p,
    g1702_p_spl_,
    g2161_n_spl_
  );


  or

  (
    g2163_n,
    g1702_n_spl_0,
    g2161_p_spl_
  );


  and

  (
    g2164_p,
    g2162_n,
    g2163_n
  );


  or

  (
    g2164_n,
    g2162_p,
    g2163_p
  );


  and

  (
    g2165_p,
    n2323_inv_n_spl_,
    g2164_p
  );


  or

  (
    g2165_n,
    n2323_inv_p_spl_0,
    g2164_n_spl_
  );


  and

  (
    g2166_p,
    n2323_inv_p_spl_0,
    g2164_n_spl_
  );


  or

  (
    g2167_n,
    g2165_p_spl_,
    g2166_p
  );


  and

  (
    g2168_p,
    n2614_inv_n_spl_,
    g1703_n_spl_
  );


  or

  (
    g2168_n,
    n2614_inv_p_spl_0,
    g1703_p_spl_0
  );


  and

  (
    g2169_p,
    g1705_n,
    g2168_n
  );


  or

  (
    g2169_n,
    g1705_p_spl_,
    g2168_p
  );


  and

  (
    g2170_p,
    n2662_o2_p_spl_0,
    g2169_n_spl_
  );


  or

  (
    g2170_n,
    n2662_o2_n_spl_,
    g2169_p_spl_
  );


  and

  (
    g2171_p,
    n2662_o2_n_spl_,
    g2169_p_spl_
  );


  or

  (
    g2171_n,
    n2662_o2_p_spl_0,
    g2169_n_spl_
  );


  and

  (
    g2172_p,
    g2170_n,
    g2171_n
  );


  or

  (
    g2172_n,
    g2170_p,
    g2171_p
  );


  and

  (
    g2173_p,
    g2167_n_spl_,
    g2172_n_spl_0
  );


  or

  (
    g2174_n,
    g2167_n_spl_,
    g2172_n_spl_0
  );


  and

  (
    g2175_p,
    g1793_n,
    g2096_n_spl_
  );


  and

  (
    g2176_p,
    g1805_p_spl_,
    g1808_p_spl_
  );


  or

  (
    g2177_n,
    g1806_p,
    g2176_p
  );


  and

  (
    g2178_p,
    n3957_lo_p_spl_0,
    n5938_o2_p_spl_
  );


  and

  (
    g2179_p,
    n3969_lo_p_spl_,
    n5938_o2_n
  );


  or

  (
    g2180_n,
    g2178_p,
    g2179_p
  );


  and

  (
    g2181_p,
    n5912_o2_n_spl_,
    lo398_buf_o2_n_spl_010
  );


  and

  (
    g2182_p,
    n5912_o2_p_spl_0,
    lo402_buf_o2_n_spl_010
  );


  or

  (
    g2183_n,
    g2181_p,
    g2182_p
  );


  and

  (
    g2184_p,
    lo554_buf_o2_p_spl_,
    g2183_n
  );


  and

  (
    g2185_p,
    n5912_o2_p_spl_0,
    lo406_buf_o2_p_spl_001
  );


  and

  (
    g2186_p,
    n5912_o2_n_spl_,
    lo390_buf_o2_p_spl_001
  );


  or

  (
    g2187_n,
    g2185_p,
    g2186_p
  );


  and

  (
    g2188_p,
    lo554_buf_o2_n,
    g2187_n
  );


  or

  (
    g2189_n,
    g2184_p,
    g2188_p
  );


  and

  (
    g2190_p,
    n5910_o2_n_spl_,
    lo398_buf_o2_n_spl_010
  );


  and

  (
    g2191_p,
    n5910_o2_p_spl_0,
    lo402_buf_o2_n_spl_010
  );


  or

  (
    g2192_n,
    g2190_p,
    g2191_p
  );


  and

  (
    g2193_p,
    lo558_buf_o2_p_spl_,
    g2192_n
  );


  and

  (
    g2194_p,
    n5910_o2_p_spl_0,
    lo406_buf_o2_p_spl_010
  );


  and

  (
    g2195_p,
    n5910_o2_n_spl_,
    lo390_buf_o2_p_spl_010
  );


  or

  (
    g2196_n,
    g2194_p,
    g2195_p
  );


  and

  (
    g2197_p,
    lo558_buf_o2_n,
    g2196_n
  );


  or

  (
    g2198_n,
    g2193_p,
    g2197_p
  );


  and

  (
    g2199_p,
    n5908_o2_n_spl_,
    lo398_buf_o2_n_spl_011
  );


  and

  (
    g2200_p,
    n5908_o2_p_spl_0,
    lo402_buf_o2_n_spl_011
  );


  or

  (
    g2201_n,
    g2199_p,
    g2200_p
  );


  and

  (
    g2202_p,
    lo574_buf_o2_p_spl_,
    g2201_n
  );


  and

  (
    g2203_p,
    n5908_o2_p_spl_0,
    lo406_buf_o2_p_spl_010
  );


  and

  (
    g2204_p,
    n5908_o2_n_spl_,
    lo390_buf_o2_p_spl_010
  );


  or

  (
    g2205_n,
    g2203_p,
    g2204_p
  );


  and

  (
    g2206_p,
    lo574_buf_o2_n,
    g2205_n
  );


  or

  (
    g2207_n,
    g2202_p,
    g2206_p
  );


  and

  (
    g2208_p,
    n5934_o2_n_spl_,
    lo398_buf_o2_n_spl_011
  );


  and

  (
    g2209_p,
    n5934_o2_p_spl_0,
    lo402_buf_o2_n_spl_011
  );


  or

  (
    g2210_n,
    g2208_p,
    g2209_p
  );


  and

  (
    g2211_p,
    lo538_buf_o2_p_spl_,
    g2210_n
  );


  and

  (
    g2212_p,
    n5934_o2_p_spl_0,
    lo406_buf_o2_p_spl_011
  );


  and

  (
    g2213_p,
    n5934_o2_n_spl_,
    lo390_buf_o2_p_spl_011
  );


  or

  (
    g2214_n,
    g2212_p,
    g2213_p
  );


  and

  (
    g2215_p,
    lo538_buf_o2_n,
    g2214_n
  );


  or

  (
    g2216_n,
    g2211_p,
    g2215_p
  );


  and

  (
    g2217_p,
    lo418_buf_o2_n_spl_,
    lo398_buf_o2_n_spl_100
  );


  and

  (
    g2218_p,
    lo418_buf_o2_p_spl_0,
    lo402_buf_o2_n_spl_100
  );


  or

  (
    g2219_n,
    g2217_p,
    g2218_p
  );


  and

  (
    g2220_p,
    lo550_buf_o2_p_spl_,
    g2219_n
  );


  and

  (
    g2221_p,
    lo418_buf_o2_p_spl_0,
    lo406_buf_o2_p_spl_011
  );


  and

  (
    g2222_p,
    lo418_buf_o2_n_spl_,
    lo390_buf_o2_p_spl_011
  );


  or

  (
    g2223_n,
    g2221_p,
    g2222_p
  );


  and

  (
    g2224_p,
    lo550_buf_o2_n,
    g2223_n
  );


  or

  (
    g2225_n,
    g2220_p,
    g2224_p
  );


  and

  (
    g2226_p,
    lo358_buf_o2_n_spl_,
    lo398_buf_o2_n_spl_100
  );


  and

  (
    g2227_p,
    lo358_buf_o2_p_spl_0,
    lo402_buf_o2_n_spl_100
  );


  or

  (
    g2228_n,
    g2226_p,
    g2227_p
  );


  and

  (
    g2229_p,
    lo570_buf_o2_p_spl_,
    g2228_n
  );


  and

  (
    g2230_p,
    lo358_buf_o2_p_spl_0,
    lo406_buf_o2_p_spl_100
  );


  and

  (
    g2231_p,
    lo358_buf_o2_n_spl_,
    lo390_buf_o2_p_spl_100
  );


  or

  (
    g2232_n,
    g2230_p,
    g2231_p
  );


  and

  (
    g2233_p,
    lo570_buf_o2_n,
    g2232_n
  );


  or

  (
    g2234_n,
    g2229_p,
    g2233_p
  );


  and

  (
    g2235_p,
    lo350_buf_o2_n_spl_,
    lo402_buf_o2_n_spl_101
  );


  and

  (
    g2236_p,
    lo350_buf_o2_p_spl_0,
    lo398_buf_o2_n_spl_101
  );


  or

  (
    g2237_n,
    g2235_p,
    g2236_p
  );


  and

  (
    g2238_p,
    lo566_buf_o2_p,
    g2237_n
  );


  and

  (
    g2239_p,
    lo350_buf_o2_n_spl_,
    lo406_buf_o2_p_spl_100
  );


  and

  (
    g2240_p,
    lo350_buf_o2_p_spl_0,
    lo390_buf_o2_p_spl_100
  );


  or

  (
    g2241_n,
    g2239_p,
    g2240_p
  );


  and

  (
    g2242_p,
    lo566_buf_o2_n,
    g2241_n
  );


  or

  (
    g2243_n,
    g2238_p,
    g2242_p
  );


  and

  (
    g2244_p,
    n2689_inv_n_spl_0,
    g1714_n_spl_0
  );


  or

  (
    g2244_n,
    n2689_inv_p_spl_0,
    g1714_p_spl_
  );


  and

  (
    g2245_p,
    n2689_inv_p_spl_1,
    g1714_p_spl_
  );


  or

  (
    g2245_n,
    n2689_inv_n_spl_,
    g1714_n_spl_0
  );


  and

  (
    g2246_p,
    g2244_n,
    g2245_n
  );


  or

  (
    g2246_n,
    g2244_p,
    g2245_p
  );


  and

  (
    g2247_p,
    g1698_p_spl_,
    g2246_n
  );


  and

  (
    g2248_p,
    g1698_n_spl_1,
    g2246_p
  );


  or

  (
    g2249_n,
    g2247_p,
    g2248_p
  );


  and

  (
    g2250_p,
    g2139_p_spl_,
    g2142_n_spl_
  );


  and

  (
    g2251_p,
    n2572_inv_n_spl_,
    n2779_inv_n_spl_1
  );


  or

  (
    g2251_n,
    n2572_inv_p_spl_1,
    n2779_inv_p_spl_0
  );


  and

  (
    g2252_p,
    n2611_inv_p_spl_1,
    n2779_inv_p_spl_1
  );


  or

  (
    g2252_n,
    n2611_inv_n_spl_,
    n2779_inv_n_spl_1
  );


  and

  (
    g2253_p,
    n2811_o2_n_spl_1,
    g2252_n
  );


  or

  (
    g2253_n,
    n2811_o2_p_spl_1,
    g2252_p
  );


  and

  (
    g2254_p,
    n2694_o2_p_spl_,
    g2253_n_spl_
  );


  or

  (
    g2254_n,
    n2694_o2_n_spl_,
    g2253_p_spl_
  );


  and

  (
    g2255_p,
    n2694_o2_n_spl_,
    g2253_p_spl_
  );


  or

  (
    g2255_n,
    n2694_o2_p_spl_,
    g2253_n_spl_
  );


  and

  (
    g2256_p,
    g2254_n,
    g2255_n
  );


  or

  (
    g2256_n,
    g2254_p,
    g2255_p
  );


  and

  (
    g2257_p,
    g2251_n,
    g2256_p
  );


  and

  (
    g2258_p,
    g2251_p,
    g2256_n
  );


  or

  (
    g2259_n,
    g2257_p,
    g2258_p
  );


  or

  (
    g2260_n,
    g2250_p_spl_,
    g2259_n_spl_
  );


  and

  (
    g2261_p,
    g2250_p_spl_,
    g2259_n_spl_
  );


  and

  (
    g2262_p,
    n3654_lo_p_spl_,
    lo494_buf_o2_p_spl_11
  );


  and

  (
    g2263_p,
    n3666_lo_p,
    lo494_buf_o2_n_spl_11
  );


  or

  (
    g2264_n,
    g2262_p,
    g2263_p
  );


  or

  (
    g2265_n,
    n4158_lo_n,
    lo490_buf_o2_n_spl_10
  );


  or

  (
    g2266_n,
    n4170_lo_n,
    lo490_buf_o2_p_spl_10
  );


  and

  (
    g2267_p,
    g2265_n,
    g2266_n
  );


  or

  (
    g2268_n,
    n4374_lo_n,
    g1898_p
  );


  and

  (
    g2269_p,
    g1725_n_spl_,
    g1768_n_spl_
  );


  or

  (
    g2270_n,
    g1758_p_spl_0,
    g2151_p_spl_
  );


  or

  (
    g2271_n,
    g1758_n_spl_1,
    g2151_n_spl_
  );


  and

  (
    g2272_p,
    g2270_n,
    g2271_n
  );


  or

  (
    g2273_n,
    g2269_p_spl_,
    g2272_p_spl_
  );


  and

  (
    g2274_p,
    g2269_p_spl_,
    g2272_p_spl_
  );


  or

  (
    g2275_n,
    g1764_p_spl_0,
    g1809_p_spl_
  );


  or

  (
    g2276_n,
    g2099_p_spl_0,
    g2275_n_spl_
  );


  and

  (
    g2277_p,
    g2108_n_spl_0,
    g2123_n_spl_0
  );


  or

  (
    g2278_n,
    g2108_n_spl_0,
    g2123_n_spl_0
  );


  and

  (
    g2279_p,
    g2117_n_spl_0,
    g2126_p_spl_0
  );


  or

  (
    g2280_n,
    g2117_n_spl_0,
    g2126_p_spl_0
  );


  and

  (
    g2281_p,
    lo590_buf_o2_p_spl_0,
    lo398_buf_o2_n_spl_101
  );


  or

  (
    g2281_n,
    lo590_buf_o2_n_spl_,
    lo398_buf_o2_p_spl_00
  );


  and

  (
    g2282_p,
    lo590_buf_o2_n_spl_,
    lo390_buf_o2_p_spl_101
  );


  or

  (
    g2282_n,
    lo590_buf_o2_p_spl_0,
    lo390_buf_o2_n_spl_00
  );


  and

  (
    g2283_p,
    g2281_n,
    g2282_n
  );


  or

  (
    g2283_n,
    g2281_p,
    g2282_p
  );


  and

  (
    g2284_p,
    lo482_buf_o2_n_spl_0,
    lo398_buf_o2_n_spl_110
  );


  or

  (
    g2284_n,
    lo482_buf_o2_p_spl_00,
    lo398_buf_o2_p_spl_00
  );


  and

  (
    g2285_p,
    lo482_buf_o2_p_spl_00,
    lo402_buf_o2_n_spl_101
  );


  or

  (
    g2285_n,
    lo482_buf_o2_n_spl_0,
    lo402_buf_o2_p_spl_0
  );


  and

  (
    g2286_p,
    g2284_n,
    g2285_n
  );


  or

  (
    g2286_n,
    g2284_p,
    g2285_p
  );


  and

  (
    g2287_p,
    lo585_buf_o2_p_spl_0,
    g2286_n
  );


  or

  (
    g2287_n,
    lo585_buf_o2_n_spl_1,
    g2286_p
  );


  and

  (
    g2288_p,
    lo482_buf_o2_p_spl_0,
    lo406_buf_o2_p_spl_101
  );


  or

  (
    g2288_n,
    lo482_buf_o2_n_spl_1,
    lo406_buf_o2_n_spl_0
  );


  and

  (
    g2289_p,
    lo482_buf_o2_n_spl_1,
    lo390_buf_o2_p_spl_101
  );


  or

  (
    g2289_n,
    lo482_buf_o2_p_spl_1,
    lo390_buf_o2_n_spl_00
  );


  and

  (
    g2290_p,
    g2288_n,
    g2289_n
  );


  or

  (
    g2290_n,
    g2288_p,
    g2289_p
  );


  and

  (
    g2291_p,
    lo585_buf_o2_n_spl_1,
    g2290_n
  );


  or

  (
    g2291_n,
    lo585_buf_o2_p_spl_1,
    g2290_p
  );


  and

  (
    g2292_p,
    g2287_n,
    g2291_n
  );


  or

  (
    g2292_n,
    g2287_p,
    g2291_p
  );


  and

  (
    g2293_p,
    g2283_p,
    g2292_n
  );


  and

  (
    g2294_p,
    g2283_n,
    g2292_p
  );


  or

  (
    g2295_n,
    g2293_p,
    g2294_p
  );


  or

  (
    g2296_n,
    g2120_n_spl_0,
    g2295_n_spl_
  );


  and

  (
    g2297_p,
    g2120_n_spl_0,
    g2295_n_spl_
  );


  and

  (
    g2298_p,
    lo510_buf_o2_n_spl_,
    lo398_buf_o2_n_spl_110
  );


  and

  (
    g2299_p,
    lo510_buf_o2_p_spl_0,
    lo402_buf_o2_n_spl_110
  );


  or

  (
    g2300_n,
    g2298_p,
    g2299_p
  );


  and

  (
    g2301_p,
    lo598_buf_o2_p_spl_,
    g2300_n
  );


  and

  (
    g2302_p,
    lo510_buf_o2_p_spl_0,
    lo406_buf_o2_p_spl_101
  );


  and

  (
    g2303_p,
    lo510_buf_o2_n_spl_,
    lo390_buf_o2_p_spl_110
  );


  or

  (
    g2304_n,
    g2302_p,
    g2303_p
  );


  and

  (
    g2305_p,
    lo598_buf_o2_n,
    g2304_n
  );


  or

  (
    g2306_n,
    g2301_p,
    g2305_p
  );


  or

  (
    g2307_n,
    lo502_buf_o2_p_spl_0,
    lo398_buf_o2_p_spl_0
  );


  or

  (
    g2308_n,
    lo502_buf_o2_n_spl_,
    lo402_buf_o2_p_spl_0
  );


  and

  (
    g2309_p,
    g2307_n,
    g2308_n
  );


  or

  (
    g2310_n,
    lo594_buf_o2_n,
    g2309_p
  );


  or

  (
    g2311_n,
    lo502_buf_o2_n_spl_,
    lo406_buf_o2_n_spl_0
  );


  or

  (
    g2312_n,
    lo502_buf_o2_p_spl_0,
    lo390_buf_o2_n_spl_0
  );


  and

  (
    g2313_p,
    g2311_n,
    g2312_n
  );


  or

  (
    g2314_n,
    lo594_buf_o2_p_spl_,
    g2313_p
  );


  and

  (
    g2315_p,
    g2310_n,
    g2314_n
  );


  or

  (
    g2316_n,
    g2306_n_spl_,
    g2315_p_spl_
  );


  and

  (
    g2317_p,
    g2306_n_spl_,
    g2315_p_spl_
  );


  and

  (
    g2318_p,
    n2641_inv_n,
    g1699_n_spl_1
  );


  and

  (
    g2319_p,
    n2641_inv_p_spl_,
    g1699_p_spl_
  );


  or

  (
    g2320_n,
    g2318_p,
    g2319_p
  );


  and

  (
    g2321_p,
    g1712_p_spl_0,
    g2320_n
  );


  or

  (
    g2322_n,
    g1785_p_spl_,
    g2321_p
  );


  and

  (
    g2323_p,
    g1774_p,
    g2322_n
  );


  and

  (
    g2324_p,
    g1774_n_spl_,
    g1787_n_spl_
  );


  or

  (
    g2325_n,
    g2323_p,
    g2324_p
  );


  and

  (
    g2326_p,
    g1697_n_spl_0,
    g1701_p_spl_
  );


  or

  (
    g2326_n,
    g1697_p_spl_,
    g1701_n_spl_0
  );


  and

  (
    g2327_p,
    g1697_p_spl_,
    g1701_n_spl_0
  );


  or

  (
    g2327_n,
    g1697_n_spl_0,
    g1701_p_spl_
  );


  and

  (
    g2328_p,
    n2323_inv_p_spl_1,
    g2327_n
  );


  or

  (
    g2328_n,
    n2323_inv_n_spl_,
    g2327_p
  );


  and

  (
    g2329_p,
    g2326_n,
    g2328_p
  );


  or

  (
    g2329_n,
    g2326_p,
    g2328_n
  );


  and

  (
    g2330_p,
    g2165_n,
    g2329_n
  );


  or

  (
    g2330_n,
    g2165_p_spl_,
    g2329_p
  );


  or

  (
    g2331_n,
    g2172_p,
    g2330_p
  );


  or

  (
    g2332_n,
    g2172_n_spl_,
    g2330_n
  );


  and

  (
    g2333_p,
    g2331_n,
    g2332_n
  );


  and

  (
    g2334_p,
    lo410_buf_o2_n_spl_0,
    lo398_buf_o2_n_spl_111
  );


  or

  (
    g2334_n,
    lo410_buf_o2_p_spl_00,
    lo398_buf_o2_p_spl_1
  );


  and

  (
    g2335_p,
    lo410_buf_o2_p_spl_00,
    lo402_buf_o2_n_spl_110
  );


  or

  (
    g2335_n,
    lo410_buf_o2_n_spl_0,
    lo402_buf_o2_p_spl_1
  );


  and

  (
    g2336_p,
    g2334_n,
    g2335_n
  );


  or

  (
    g2336_n,
    g2334_p,
    g2335_p
  );


  and

  (
    g2337_p,
    lo546_buf_o2_p_spl_0,
    g2336_n
  );


  or

  (
    g2337_n,
    lo546_buf_o2_n_spl_,
    g2336_p
  );


  and

  (
    g2338_p,
    lo410_buf_o2_p_spl_0,
    lo406_buf_o2_p_spl_11
  );


  or

  (
    g2338_n,
    lo410_buf_o2_n_spl_1,
    lo406_buf_o2_n_spl_1
  );


  and

  (
    g2339_p,
    lo410_buf_o2_n_spl_1,
    lo390_buf_o2_p_spl_110
  );


  or

  (
    g2339_n,
    lo410_buf_o2_p_spl_1,
    lo390_buf_o2_n_spl_1
  );


  and

  (
    g2340_p,
    g2338_n,
    g2339_n
  );


  or

  (
    g2340_n,
    g2338_p,
    g2339_p
  );


  and

  (
    g2341_p,
    lo546_buf_o2_n_spl_,
    g2340_n
  );


  or

  (
    g2341_n,
    lo546_buf_o2_p_spl_0,
    g2340_p
  );


  and

  (
    g2342_p,
    g2337_n,
    g2341_n
  );


  or

  (
    g2342_n,
    g2337_p,
    g2341_p
  );


  and

  (
    g2343_p,
    lo382_buf_o2_n_spl_00,
    lo398_buf_o2_n_spl_111
  );


  or

  (
    g2343_n,
    lo382_buf_o2_p_spl_00,
    lo398_buf_o2_p_spl_1
  );


  and

  (
    g2344_p,
    lo382_buf_o2_p_spl_01,
    lo402_buf_o2_n_spl_11
  );


  or

  (
    g2344_n,
    lo382_buf_o2_n_spl_0,
    lo402_buf_o2_p_spl_1
  );


  and

  (
    g2345_p,
    g2343_n,
    g2344_n
  );


  or

  (
    g2345_n,
    g2343_p,
    g2344_p
  );


  and

  (
    g2346_p,
    n4293_lo_p_spl_0,
    g2345_n
  );


  or

  (
    g2346_n,
    n4293_lo_n_spl_1,
    g2345_p
  );


  and

  (
    g2347_p,
    lo382_buf_o2_p_spl_01,
    lo406_buf_o2_p_spl_11
  );


  or

  (
    g2347_n,
    lo382_buf_o2_n_spl_1,
    lo406_buf_o2_n_spl_1
  );


  and

  (
    g2348_p,
    lo382_buf_o2_n_spl_1,
    lo390_buf_o2_p_spl_11
  );


  or

  (
    g2348_n,
    lo382_buf_o2_p_spl_1,
    lo390_buf_o2_n_spl_1
  );


  and

  (
    g2349_p,
    g2347_n,
    g2348_n
  );


  or

  (
    g2349_n,
    g2347_p,
    g2348_p
  );


  and

  (
    g2350_p,
    n4293_lo_n_spl_1,
    g2349_n
  );


  or

  (
    g2350_n,
    n4293_lo_p_spl_1,
    g2349_p
  );


  and

  (
    g2351_p,
    g2346_n,
    g2350_n
  );


  or

  (
    g2351_n,
    g2346_p,
    g2350_p
  );


  and

  (
    g2352_p,
    g2342_p,
    g2351_n
  );


  and

  (
    g2353_p,
    g2342_n,
    g2351_p
  );


  or

  (
    g2354_n,
    g2352_p,
    g2353_p
  );


  and

  (
    g2355_p,
    n4545_lo_n_spl_,
    g1716_p
  );


  or

  (
    g2355_n,
    n4545_lo_p_spl_,
    g1716_n_spl_
  );


  and

  (
    g2356_p,
    n4545_lo_p_spl_,
    n2711_o2_n_spl_
  );


  or

  (
    g2356_n,
    n4545_lo_n_spl_,
    n2711_o2_p_spl_
  );


  and

  (
    g2357_p,
    g2355_n,
    g2356_n
  );


  or

  (
    g2357_n,
    g2355_p,
    g2356_p
  );


  and

  (
    g2358_p,
    g1792_p_spl_,
    g2357_n
  );


  and

  (
    g2359_p,
    g1792_n,
    g2357_p
  );


  or

  (
    g2360_n,
    g2358_p,
    g2359_p
  );


  or

  (
    g2361_n,
    n4242_lo_n,
    g2129_p
  );


  or

  (
    g2362_n,
    n4386_lo_n,
    g2132_p
  );


  or

  (
    g2363_n,
    n4386_lo_p_spl_,
    g2132_n_spl_
  );


  or

  (
    g2364_n,
    n4398_lo_p_spl_,
    g1802_n_spl_
  );


  and

  (
    g2365_p,
    g2133_n_spl_,
    g2364_n
  );


  and

  (
    g2366_p,
    n3978_lo_p_spl_,
    lo490_buf_o2_p_spl_10
  );


  and

  (
    g2367_p,
    n3990_lo_p,
    lo490_buf_o2_n_spl_11
  );


  and

  (
    g2368_p,
    n4050_lo_p_spl_,
    lo490_buf_o2_p_spl_11
  );


  and

  (
    g2369_p,
    n4062_lo_p,
    lo490_buf_o2_n_spl_11
  );


  and

  (
    g2370_p,
    g1763_n_spl_0,
    g2276_n_spl_0
  );


  or

  (
    g2371_n,
    g1763_n_spl_1,
    g2276_n_spl_0
  );


  and

  (
    g2372_p,
    g1764_p_spl_0,
    g2137_p_spl_0
  );


  and

  (
    g2373_p,
    g1807_n_spl_,
    g2160_n_spl_0
  );


  and

  (
    g2374_p,
    g1796_p_spl_0,
    g2175_p_spl_
  );


  and

  (
    g2375_p,
    g2098_n_spl_,
    g2135_p_spl_
  );


  or

  (
    g2376_n,
    g1803_p_spl_,
    g2375_p
  );


  and

  (
    g2377_p,
    g2099_p_spl_0,
    g2137_p_spl_0
  );


  or

  (
    g2378_n,
    g1804_p_spl_,
    g2377_p
  );


  and

  (
    g2379_p,
    g2137_p_spl_1,
    g2275_n_spl_
  );


  or

  (
    g2380_n,
    g2160_n_spl_0,
    g2177_n_spl_
  );


  and

  (
    g2381_p,
    n4302_lo_p_spl_0,
    g2264_n_spl_0
  );


  or

  (
    g2382_n,
    n4302_lo_p_spl_0,
    g2264_n_spl_0
  );


  and

  (
    g2383_p,
    g2267_p_spl_,
    g2365_p_spl_
  );


  or

  (
    g2384_n,
    n4374_lo_p_spl_,
    g1898_n_spl_
  );


  and

  (
    g2385_p,
    g2268_n_spl_,
    g2384_n
  );


  or

  (
    g2386_n,
    n4242_lo_p_spl_,
    g2129_n_spl_
  );


  and

  (
    g2387_p,
    g2361_n_spl_,
    g2386_n
  );


  and

  (
    g2388_p,
    g2362_n_spl_,
    g2363_n_spl_
  );


  and

  (
    g2389_p,
    G92_p_spl_,
    G124_p_spl_0
  );


  and

  (
    g2390_p,
    G93_p,
    G124_n_spl_0
  );


  and

  (
    g2391_p,
    G94_p_spl_,
    G124_p_spl_0
  );


  and

  (
    g2392_p,
    G95_p,
    G124_n_spl_0
  );


  and

  (
    g2393_p,
    G107_p_spl_,
    G124_p_spl_1
  );


  and

  (
    g2394_p,
    G108_p,
    G124_n_spl_
  );


  buf

  (
    G5193,
    n3399_lo_n
  );


  buf

  (
    G5194,
    n3963_lo_n
  );


  buf

  (
    G5195,
    n4587_lo_n_spl_
  );


  buf

  (
    G5196,
    n4419_lo_n_spl_0
  );


  buf

  (
    G5197,
    n4131_lo_n
  );


  buf

  (
    G5198,
    n4179_lo_n
  );


  not

  (
    G5199,
    g1049_n_spl_
  );


  buf

  (
    G5200,
    n4431_lo_n
  );


  buf

  (
    G5201,
    n4419_lo_n_spl_0
  );


  buf

  (
    G5202,
    n4419_lo_n_spl_
  );


  buf

  (
    G5203,
    n4107_lo_n
  );


  buf

  (
    G5204,
    n4155_lo_n
  );


  buf

  (
    G5205,
    g1050_p
  );


  buf

  (
    G5206,
    n3795_lo_n_spl_
  );


  buf

  (
    G5207,
    n4443_lo_n_spl_
  );


  buf

  (
    G5208,
    n4479_lo_n_spl_
  );


  buf

  (
    G5209,
    n4467_lo_n_spl_
  );


  buf

  (
    G5210,
    g1051_p
  );


  buf

  (
    G5211,
    g1052_p
  );


  buf

  (
    G5212,
    g1053_n
  );


  buf

  (
    G5213,
    g1054_n_spl_
  );


  buf

  (
    G5214,
    n3375_lo_p_spl_111
  );


  buf

  (
    G5215,
    n3399_lo_p_spl_1
  );


  buf

  (
    G5216,
    n2619_lo_p_spl_
  );


  buf

  (
    G5217,
    n4431_lo_p_spl_
  );


  buf

  (
    G5218,
    n3975_lo_p
  );


  buf

  (
    G5219,
    n4431_lo_p_spl_
  );


  buf

  (
    G5220,
    g1056_n
  );


  buf

  (
    G5221,
    g1055_n_spl_11
  );


  buf

  (
    G5222,
    n2619_lo_n_spl_0
  );


  buf

  (
    G5223,
    n2619_lo_n_spl_0
  );


  buf

  (
    G5224,
    n2619_lo_n_spl_1
  );


  buf

  (
    G5225,
    n2619_lo_n_spl_1
  );


  buf

  (
    G5226,
    n3975_lo_n_spl_
  );


  buf

  (
    G5227,
    n3975_lo_n_spl_
  );


  buf

  (
    G5228,
    g1060_n
  );


  buf

  (
    G5229,
    g1064_n_spl_
  );


  buf

  (
    G5230,
    g1064_n_spl_
  );


  buf

  (
    G5231,
    g1065_n
  );


  buf

  (
    G5232,
    g1070_p
  );


  buf

  (
    G5233,
    g1075_p
  );


  buf

  (
    G5234,
    g1080_p
  );


  buf

  (
    G5235,
    g1085_p
  );


  buf

  (
    G5236,
    g1091_p
  );


  buf

  (
    G5237,
    g1100_p
  );


  not

  (
    G5238,
    g1102_n_spl_
  );


  buf

  (
    G5239,
    g1106_p_spl_
  );


  buf

  (
    G5240,
    g1106_p_spl_
  );


  not

  (
    G5241,
    g1102_n_spl_
  );


  not

  (
    G5242,
    g1111_n_spl_
  );


  not

  (
    G5243,
    g1120_n_spl_
  );


  not

  (
    G5244,
    g1126_p_spl_
  );


  buf

  (
    G5245,
    g1127_n_spl_
  );


  not

  (
    G5246,
    g1126_p_spl_
  );


  buf

  (
    G5247,
    g1127_n_spl_
  );


  not

  (
    G5248,
    g1132_n_spl_1
  );


  buf

  (
    G5249,
    g1137_p_spl_1
  );


  not

  (
    G5250,
    g1142_n_spl_1
  );


  buf

  (
    G5251,
    n2853_o2_p_spl_1
  );


  buf

  (
    G5252,
    g1151_n
  );


  not

  (
    G5253,
    g1155_n_spl_1
  );


  not

  (
    G5254,
    g1158_n_spl_1
  );


  not

  (
    G5255,
    g1164_n_spl_1
  );


  buf

  (
    G5256,
    g1173_n
  );


  not

  (
    G5257,
    g1182_n_spl_1
  );


  not

  (
    G5258,
    g1187_n_spl_1
  );


  not

  (
    G5259,
    g1194_n_spl_1
  );


  buf

  (
    G5260,
    g1200_p_spl_1
  );


  not

  (
    G5261,
    g1212_n_spl_
  );


  not

  (
    G5262,
    g1233_n_spl_
  );


  not

  (
    G5263,
    g1248_n
  );


  not

  (
    G5264,
    g1257_n
  );


  buf

  (
    G5265,
    g1267_p
  );


  buf

  (
    G5266,
    g1277_p
  );


  buf

  (
    G5267,
    g1286_p
  );


  buf

  (
    G5268,
    g1295_p
  );


  buf

  (
    G5269,
    g1304_p
  );


  not

  (
    G5270,
    g1313_p
  );


  buf

  (
    G5271,
    g1322_p
  );


  buf

  (
    G5272,
    g1331_p
  );


  buf

  (
    G5273,
    g1340_p
  );


  not

  (
    G5274,
    g1349_p
  );


  buf

  (
    G5275,
    g1359_p
  );


  not

  (
    G5276,
    g1369_n
  );


  buf

  (
    G5277,
    g1379_p
  );


  buf

  (
    G5278,
    g1389_p
  );


  buf

  (
    G5279,
    g1399_p
  );


  not

  (
    G5280,
    g1409_n
  );


  buf

  (
    G5281,
    g1419_p
  );


  buf

  (
    G5282,
    g1429_p
  );


  buf

  (
    G5283,
    g1443_p
  );


  buf

  (
    G5284,
    g1446_p
  );


  not

  (
    G5285,
    g1449_n_spl_1
  );


  not

  (
    G5286,
    g1453_n_spl_1
  );


  not

  (
    G5287,
    g1457_n_spl_1
  );


  not

  (
    G5288,
    g1460_n_spl_1
  );


  not

  (
    G5289,
    g1467_n
  );


  not

  (
    G5290,
    g1470_n_spl_1
  );


  not

  (
    G5291,
    g1476_n_spl_1
  );


  not

  (
    G5292,
    g1482_n_spl_1
  );


  not

  (
    G5293,
    g1486_n_spl_1
  );


  buf

  (
    G5294,
    g1495_n
  );


  buf

  (
    G5295,
    g1504_p
  );


  buf

  (
    G5296,
    g1513_p
  );


  buf

  (
    G5297,
    g1522_p
  );


  buf

  (
    G5298,
    g1531_p
  );


  buf

  (
    G5299,
    g1540_p
  );


  buf

  (
    G5300,
    g1549_p
  );


  buf

  (
    G5301,
    g1558_p
  );


  buf

  (
    G5302,
    g1568_p
  );


  buf

  (
    G5303,
    g1578_p
  );


  buf

  (
    G5304,
    g1588_p
  );


  buf

  (
    G5305,
    g1598_p
  );


  buf

  (
    G5306,
    g1608_p
  );


  buf

  (
    G5307,
    g1618_p
  );


  buf

  (
    G5308,
    g1628_p
  );


  buf

  (
    G5309,
    g1638_p
  );


  buf

  (
    G5310,
    g1642_p
  );


  buf

  (
    G5311,
    g1647_p
  );


  not

  (
    G5312,
    g1660_n
  );


  not

  (
    G5313,
    g1669_n
  );


  buf

  (
    G5314,
    g1679_n
  );


  buf

  (
    G5315,
    g1689_n
  );


  buf

  (
    n7230_li000_li000,
    G1_p
  );


  buf

  (
    n7233_li001_li001,
    n2610_lo_p
  );


  buf

  (
    n7236_li002_li002,
    n2613_lo_p
  );


  buf

  (
    n7239_li003_li003,
    n2616_lo_p
  );


  buf

  (
    n7242_li004_li004,
    G2_p
  );


  buf

  (
    n7245_li005_li005,
    n2622_lo_p
  );


  buf

  (
    n7248_li006_li006,
    n2625_lo_p
  );


  buf

  (
    n7254_li008_li008,
    G3_p
  );


  buf

  (
    n7257_li009_li009,
    n2634_lo_p
  );


  buf

  (
    n7260_li010_li010,
    n2637_lo_p
  );


  buf

  (
    n7263_li011_li011,
    n2640_lo_p
  );


  buf

  (
    n7266_li012_li012,
    G4_p
  );


  buf

  (
    n7269_li013_li013,
    n2646_lo_p
  );


  buf

  (
    n7272_li014_li014,
    n2649_lo_p
  );


  buf

  (
    n7275_li015_li015,
    n2652_lo_p
  );


  buf

  (
    n7278_li016_li016,
    G5_p
  );


  buf

  (
    n7281_li017_li017,
    n2658_lo_p
  );


  buf

  (
    n7284_li018_li018,
    n2661_lo_p
  );


  buf

  (
    n7287_li019_li019,
    n2664_lo_p
  );


  buf

  (
    n7290_li020_li020,
    G6_p
  );


  buf

  (
    n7293_li021_li021,
    n2670_lo_p
  );


  buf

  (
    n7296_li022_li022,
    n2673_lo_p
  );


  buf

  (
    n7299_li023_li023,
    n2676_lo_p
  );


  buf

  (
    n7302_li024_li024,
    G7_p
  );


  buf

  (
    n7305_li025_li025,
    n2682_lo_p
  );


  buf

  (
    n7308_li026_li026,
    n2685_lo_p
  );


  buf

  (
    n7311_li027_li027,
    n2688_lo_p
  );


  buf

  (
    n7314_li028_li028,
    G8_p
  );


  buf

  (
    n7317_li029_li029,
    n2694_lo_p
  );


  buf

  (
    n7320_li030_li030,
    n2697_lo_p
  );


  buf

  (
    n7323_li031_li031,
    n2700_lo_p
  );


  buf

  (
    n7326_li032_li032,
    G9_p
  );


  buf

  (
    n7329_li033_li033,
    n2706_lo_p
  );


  buf

  (
    n7332_li034_li034,
    n2709_lo_p
  );


  buf

  (
    n7335_li035_li035,
    n2712_lo_p
  );


  buf

  (
    n7338_li036_li036,
    G10_p
  );


  buf

  (
    n7341_li037_li037,
    n2718_lo_p
  );


  buf

  (
    n7344_li038_li038,
    n2721_lo_p
  );


  buf

  (
    n7347_li039_li039,
    n2724_lo_p
  );


  buf

  (
    n7350_li040_li040,
    G11_p
  );


  buf

  (
    n7353_li041_li041,
    n2730_lo_p
  );


  buf

  (
    n7356_li042_li042,
    n2733_lo_p
  );


  buf

  (
    n7359_li043_li043,
    n2736_lo_p
  );


  buf

  (
    n7362_li044_li044,
    G12_p
  );


  buf

  (
    n7365_li045_li045,
    n2742_lo_p
  );


  buf

  (
    n7368_li046_li046,
    n2745_lo_p
  );


  buf

  (
    n7371_li047_li047,
    n2748_lo_p
  );


  buf

  (
    n7374_li048_li048,
    G13_p
  );


  buf

  (
    n7377_li049_li049,
    n2754_lo_p
  );


  buf

  (
    n7380_li050_li050,
    n2757_lo_p
  );


  buf

  (
    n7383_li051_li051,
    n2760_lo_p
  );


  buf

  (
    n7386_li052_li052,
    G14_p
  );


  buf

  (
    n7389_li053_li053,
    n2766_lo_p
  );


  buf

  (
    n7392_li054_li054,
    n2769_lo_p
  );


  buf

  (
    n7395_li055_li055,
    n2772_lo_p
  );


  buf

  (
    n7398_li056_li056,
    G15_p
  );


  buf

  (
    n7401_li057_li057,
    n2778_lo_p
  );


  buf

  (
    n7404_li058_li058,
    n2781_lo_p
  );


  buf

  (
    n7407_li059_li059,
    n2784_lo_p
  );


  buf

  (
    n7410_li060_li060,
    G16_p
  );


  buf

  (
    n7413_li061_li061,
    n2790_lo_p
  );


  buf

  (
    n7416_li062_li062,
    n2793_lo_p
  );


  buf

  (
    n7419_li063_li063,
    n2796_lo_p
  );


  buf

  (
    n7422_li064_li064,
    G17_p
  );


  buf

  (
    n7425_li065_li065,
    n2802_lo_p
  );


  buf

  (
    n7428_li066_li066,
    n2805_lo_p
  );


  buf

  (
    n7431_li067_li067,
    n2808_lo_p
  );


  buf

  (
    n7434_li068_li068,
    G18_p
  );


  buf

  (
    n7437_li069_li069,
    n2814_lo_p
  );


  buf

  (
    n7440_li070_li070,
    n2817_lo_p
  );


  buf

  (
    n7443_li071_li071,
    n2820_lo_p
  );


  buf

  (
    n7446_li072_li072,
    G19_p
  );


  buf

  (
    n7449_li073_li073,
    n2826_lo_p
  );


  buf

  (
    n7452_li074_li074,
    n2829_lo_p
  );


  buf

  (
    n7458_li076_li076,
    G20_p
  );


  buf

  (
    n7461_li077_li077,
    n2838_lo_p
  );


  buf

  (
    n7464_li078_li078,
    n2841_lo_p
  );


  buf

  (
    n7467_li079_li079,
    n2844_lo_p
  );


  buf

  (
    n7470_li080_li080,
    G21_p
  );


  buf

  (
    n7473_li081_li081,
    n2850_lo_p
  );


  buf

  (
    n7476_li082_li082,
    n2853_lo_p
  );


  buf

  (
    n7482_li084_li084,
    G22_p
  );


  buf

  (
    n7485_li085_li085,
    n2862_lo_p
  );


  buf

  (
    n7488_li086_li086,
    n2865_lo_p
  );


  buf

  (
    n7491_li087_li087,
    n2868_lo_p
  );


  buf

  (
    n7494_li088_li088,
    G23_p
  );


  buf

  (
    n7497_li089_li089,
    n2874_lo_p
  );


  buf

  (
    n7500_li090_li090,
    n2877_lo_p
  );


  buf

  (
    n7503_li091_li091,
    n2880_lo_p
  );


  buf

  (
    n7506_li092_li092,
    G24_p
  );


  buf

  (
    n7509_li093_li093,
    n2886_lo_p
  );


  buf

  (
    n7512_li094_li094,
    n2889_lo_p
  );


  buf

  (
    n7515_li095_li095,
    n2892_lo_p
  );


  buf

  (
    n7518_li096_li096,
    G25_p
  );


  buf

  (
    n7521_li097_li097,
    n2898_lo_p
  );


  buf

  (
    n7524_li098_li098,
    n2901_lo_p
  );


  buf

  (
    n7527_li099_li099,
    n2904_lo_p
  );


  buf

  (
    n7530_li100_li100,
    G26_p
  );


  buf

  (
    n7533_li101_li101,
    n2910_lo_p
  );


  buf

  (
    n7536_li102_li102,
    n2913_lo_p
  );


  buf

  (
    n7539_li103_li103,
    n2916_lo_p
  );


  buf

  (
    n7542_li104_li104,
    G27_p
  );


  buf

  (
    n7545_li105_li105,
    n2922_lo_p
  );


  buf

  (
    n7548_li106_li106,
    n2925_lo_p
  );


  buf

  (
    n7551_li107_li107,
    n2928_lo_p
  );


  buf

  (
    n7554_li108_li108,
    G28_p
  );


  buf

  (
    n7557_li109_li109,
    n2934_lo_p
  );


  buf

  (
    n7560_li110_li110,
    n2937_lo_p
  );


  buf

  (
    n7563_li111_li111,
    n2940_lo_p
  );


  buf

  (
    n7566_li112_li112,
    G29_p
  );


  buf

  (
    n7569_li113_li113,
    n2946_lo_p
  );


  buf

  (
    n7572_li114_li114,
    n2949_lo_p
  );


  buf

  (
    n7575_li115_li115,
    n2952_lo_p
  );


  buf

  (
    n7578_li116_li116,
    G30_p
  );


  buf

  (
    n7581_li117_li117,
    n2958_lo_p
  );


  buf

  (
    n7584_li118_li118,
    n2961_lo_p
  );


  buf

  (
    n7587_li119_li119,
    n2964_lo_p
  );


  buf

  (
    n7590_li120_li120,
    G31_p
  );


  buf

  (
    n7593_li121_li121,
    n2970_lo_p
  );


  buf

  (
    n7596_li122_li122,
    n2973_lo_p
  );


  buf

  (
    n7599_li123_li123,
    n2976_lo_p
  );


  buf

  (
    n7602_li124_li124,
    G32_p
  );


  buf

  (
    n7605_li125_li125,
    n2982_lo_p
  );


  buf

  (
    n7608_li126_li126,
    n2985_lo_p
  );


  buf

  (
    n7611_li127_li127,
    n2988_lo_p
  );


  buf

  (
    n7614_li128_li128,
    G33_p
  );


  buf

  (
    n7617_li129_li129,
    n2994_lo_p
  );


  buf

  (
    n7620_li130_li130,
    n2997_lo_p
  );


  buf

  (
    n7623_li131_li131,
    n3000_lo_p
  );


  buf

  (
    n7626_li132_li132,
    G34_p
  );


  buf

  (
    n7629_li133_li133,
    n3006_lo_p
  );


  buf

  (
    n7632_li134_li134,
    n3009_lo_p
  );


  buf

  (
    n7635_li135_li135,
    n3012_lo_p
  );


  buf

  (
    n7638_li136_li136,
    G35_p
  );


  buf

  (
    n7641_li137_li137,
    n3018_lo_p
  );


  buf

  (
    n7644_li138_li138,
    n3021_lo_p
  );


  buf

  (
    n7647_li139_li139,
    n3024_lo_p
  );


  buf

  (
    n7650_li140_li140,
    G36_p
  );


  buf

  (
    n7653_li141_li141,
    n3030_lo_p
  );


  buf

  (
    n7656_li142_li142,
    n3033_lo_p
  );


  buf

  (
    n7659_li143_li143,
    n3036_lo_p
  );


  buf

  (
    n7662_li144_li144,
    G37_p
  );


  buf

  (
    n7665_li145_li145,
    n3042_lo_p
  );


  buf

  (
    n7668_li146_li146,
    n3045_lo_p
  );


  buf

  (
    n7671_li147_li147,
    n3048_lo_p
  );


  buf

  (
    n7674_li148_li148,
    G38_p
  );


  buf

  (
    n7677_li149_li149,
    n3054_lo_p
  );


  buf

  (
    n7680_li150_li150,
    n3057_lo_p
  );


  buf

  (
    n7683_li151_li151,
    n3060_lo_p
  );


  buf

  (
    n7686_li152_li152,
    G39_p
  );


  buf

  (
    n7689_li153_li153,
    n3066_lo_p
  );


  buf

  (
    n7692_li154_li154,
    n3069_lo_p
  );


  buf

  (
    n7695_li155_li155,
    n3072_lo_p
  );


  buf

  (
    n7698_li156_li156,
    G40_p
  );


  buf

  (
    n7701_li157_li157,
    n3078_lo_p
  );


  buf

  (
    n7704_li158_li158,
    n3081_lo_p
  );


  buf

  (
    n7707_li159_li159,
    n3084_lo_p
  );


  buf

  (
    n7710_li160_li160,
    G41_p
  );


  buf

  (
    n7713_li161_li161,
    n3090_lo_p
  );


  buf

  (
    n7716_li162_li162,
    n3093_lo_p
  );


  buf

  (
    n7719_li163_li163,
    n3096_lo_p
  );


  buf

  (
    n7722_li164_li164,
    G42_p
  );


  buf

  (
    n7725_li165_li165,
    n3102_lo_p
  );


  buf

  (
    n7728_li166_li166,
    n3105_lo_p
  );


  buf

  (
    n7731_li167_li167,
    n3108_lo_p
  );


  buf

  (
    n7734_li168_li168,
    G43_p
  );


  buf

  (
    n7737_li169_li169,
    n3114_lo_p
  );


  buf

  (
    n7740_li170_li170,
    n3117_lo_p
  );


  buf

  (
    n7746_li172_li172,
    G44_p
  );


  buf

  (
    n7749_li173_li173,
    n3126_lo_p
  );


  buf

  (
    n7752_li174_li174,
    n3129_lo_p
  );


  buf

  (
    n7758_li176_li176,
    G45_p
  );


  buf

  (
    n7761_li177_li177,
    n3138_lo_p
  );


  buf

  (
    n7764_li178_li178,
    n3141_lo_p
  );


  buf

  (
    n7767_li179_li179,
    n3144_lo_p
  );


  buf

  (
    n7770_li180_li180,
    G46_p
  );


  buf

  (
    n7773_li181_li181,
    n3150_lo_p
  );


  buf

  (
    n7776_li182_li182,
    n3153_lo_p
  );


  buf

  (
    n7782_li184_li184,
    G47_p
  );


  buf

  (
    n7785_li185_li185,
    n3162_lo_p
  );


  buf

  (
    n7788_li186_li186,
    n3165_lo_p
  );


  buf

  (
    n7794_li188_li188,
    G48_p
  );


  buf

  (
    n7797_li189_li189,
    n3174_lo_p
  );


  buf

  (
    n7800_li190_li190,
    n3177_lo_p
  );


  buf

  (
    n7806_li192_li192,
    G49_p
  );


  buf

  (
    n7809_li193_li193,
    n3186_lo_p
  );


  buf

  (
    n7812_li194_li194,
    n3189_lo_p
  );


  buf

  (
    n7815_li195_li195,
    n3192_lo_p
  );


  buf

  (
    n7818_li196_li196,
    G50_p
  );


  buf

  (
    n7821_li197_li197,
    n3198_lo_p
  );


  buf

  (
    n7824_li198_li198,
    n3201_lo_p
  );


  buf

  (
    n7830_li200_li200,
    G51_p
  );


  buf

  (
    n7833_li201_li201,
    n3210_lo_p
  );


  buf

  (
    n7836_li202_li202,
    n3213_lo_p
  );


  buf

  (
    n7839_li203_li203,
    n3216_lo_p
  );


  buf

  (
    n7842_li204_li204,
    G52_p
  );


  buf

  (
    n7845_li205_li205,
    n3222_lo_p
  );


  buf

  (
    n7848_li206_li206,
    n3225_lo_p
  );


  buf

  (
    n7854_li208_li208,
    G53_p
  );


  buf

  (
    n7857_li209_li209,
    n3234_lo_p
  );


  buf

  (
    n7860_li210_li210,
    n3237_lo_p
  );


  buf

  (
    n7863_li211_li211,
    n3240_lo_p
  );


  buf

  (
    n7866_li212_li212,
    G54_p
  );


  buf

  (
    n7869_li213_li213,
    n3246_lo_p
  );


  buf

  (
    n7872_li214_li214,
    n3249_lo_p
  );


  buf

  (
    n7875_li215_li215,
    n3252_lo_p_spl_
  );


  buf

  (
    n7878_li216_li216,
    G55_p
  );


  buf

  (
    n7881_li217_li217,
    n3258_lo_p
  );


  buf

  (
    n7884_li218_li218,
    n3261_lo_p
  );


  buf

  (
    n7887_li219_li219,
    n3264_lo_p
  );


  buf

  (
    n7890_li220_li220,
    G56_p
  );


  buf

  (
    n7893_li221_li221,
    n3270_lo_p
  );


  buf

  (
    n7896_li222_li222,
    n3273_lo_p
  );


  buf

  (
    n7899_li223_li223,
    n3276_lo_p
  );


  buf

  (
    n7902_li224_li224,
    G57_p
  );


  buf

  (
    n7905_li225_li225,
    n3282_lo_p
  );


  buf

  (
    n7908_li226_li226,
    n3285_lo_p
  );


  buf

  (
    n7914_li228_li228,
    G58_p
  );


  buf

  (
    n7917_li229_li229,
    n3294_lo_p
  );


  buf

  (
    n7920_li230_li230,
    n3297_lo_p
  );


  buf

  (
    n7926_li232_li232,
    G59_p
  );


  buf

  (
    n7929_li233_li233,
    n3306_lo_p
  );


  buf

  (
    n7932_li234_li234,
    n3309_lo_p
  );


  buf

  (
    n7938_li236_li236,
    G60_p
  );


  buf

  (
    n7941_li237_li237,
    n3318_lo_p
  );


  buf

  (
    n7944_li238_li238,
    n3321_lo_p
  );


  buf

  (
    n7950_li240_li240,
    G61_p
  );


  buf

  (
    n7953_li241_li241,
    n3330_lo_p
  );


  buf

  (
    n7956_li242_li242,
    n3333_lo_p
  );


  buf

  (
    n7959_li243_li243,
    n3336_lo_p
  );


  buf

  (
    n7962_li244_li244,
    G62_p
  );


  buf

  (
    n7965_li245_li245,
    n3342_lo_p
  );


  buf

  (
    n7968_li246_li246,
    n3345_lo_p
  );


  buf

  (
    n7971_li247_li247,
    n3348_lo_p
  );


  buf

  (
    n7974_li248_li248,
    G63_p
  );


  buf

  (
    n7977_li249_li249,
    n3354_lo_p
  );


  buf

  (
    n7980_li250_li250,
    n3357_lo_p
  );


  buf

  (
    n7983_li251_li251,
    n3360_lo_p
  );


  buf

  (
    n7986_li252_li252,
    G64_p
  );


  buf

  (
    n7989_li253_li253,
    n3366_lo_p
  );


  buf

  (
    n7992_li254_li254,
    n3369_lo_p
  );


  buf

  (
    n7995_li255_li255,
    n3372_lo_p
  );


  buf

  (
    n7998_li256_li256,
    G65_p
  );


  buf

  (
    n8001_li257_li257,
    n3378_lo_p
  );


  buf

  (
    n8004_li258_li258,
    n3381_lo_p
  );


  buf

  (
    n8007_li259_li259,
    n3384_lo_p
  );


  buf

  (
    n8010_li260_li260,
    G66_p
  );


  buf

  (
    n8013_li261_li261,
    n3390_lo_p
  );


  buf

  (
    n8016_li262_li262,
    n3393_lo_p
  );


  buf

  (
    n8019_li263_li263,
    n3396_lo_p
  );


  buf

  (
    n8022_li264_li264,
    G67_p
  );


  buf

  (
    n8025_li265_li265,
    n3402_lo_p
  );


  buf

  (
    n8028_li266_li266,
    n3405_lo_p
  );


  buf

  (
    n8031_li267_li267,
    n3408_lo_p
  );


  buf

  (
    n8034_li268_li268,
    G68_p
  );


  buf

  (
    n8037_li269_li269,
    n3414_lo_p
  );


  buf

  (
    n8040_li270_li270,
    n3417_lo_p
  );


  buf

  (
    n8043_li271_li271,
    n3420_lo_p
  );


  buf

  (
    n8046_li272_li272,
    G69_p
  );


  buf

  (
    n8049_li273_li273,
    n3426_lo_p
  );


  buf

  (
    n8052_li274_li274,
    n3429_lo_p
  );


  buf

  (
    n8055_li275_li275,
    n3432_lo_p
  );


  buf

  (
    n8058_li276_li276,
    G70_p
  );


  buf

  (
    n8061_li277_li277,
    n3438_lo_p
  );


  buf

  (
    n8064_li278_li278,
    n3441_lo_p
  );


  buf

  (
    n8067_li279_li279,
    n3444_lo_p
  );


  buf

  (
    n8070_li280_li280,
    G71_p
  );


  buf

  (
    n8073_li281_li281,
    n3450_lo_p
  );


  buf

  (
    n8076_li282_li282,
    n3453_lo_p
  );


  buf

  (
    n8079_li283_li283,
    n3456_lo_p
  );


  buf

  (
    n8082_li284_li284,
    G72_p
  );


  buf

  (
    n8085_li285_li285,
    n3462_lo_p
  );


  buf

  (
    n8088_li286_li286,
    n3465_lo_p
  );


  buf

  (
    n8091_li287_li287,
    n3468_lo_p
  );


  buf

  (
    n8094_li288_li288,
    G73_p
  );


  buf

  (
    n8097_li289_li289,
    n3474_lo_p
  );


  buf

  (
    n8100_li290_li290,
    n3477_lo_p
  );


  buf

  (
    n8103_li291_li291,
    n3480_lo_p
  );


  buf

  (
    n8106_li292_li292,
    G74_p
  );


  buf

  (
    n8109_li293_li293,
    n3486_lo_p
  );


  buf

  (
    n8112_li294_li294,
    n3489_lo_p
  );


  buf

  (
    n8115_li295_li295,
    n3492_lo_p
  );


  buf

  (
    n8118_li296_li296,
    G75_p
  );


  buf

  (
    n8121_li297_li297,
    n3498_lo_p
  );


  buf

  (
    n8124_li298_li298,
    n3501_lo_p
  );


  buf

  (
    n8127_li299_li299,
    n3504_lo_p
  );


  buf

  (
    n8130_li300_li300,
    G76_p
  );


  buf

  (
    n8133_li301_li301,
    n3510_lo_p
  );


  buf

  (
    n8136_li302_li302,
    n3513_lo_p
  );


  buf

  (
    n8139_li303_li303,
    n3516_lo_p
  );


  buf

  (
    n8142_li304_li304,
    G77_p
  );


  buf

  (
    n8145_li305_li305,
    n3522_lo_p
  );


  buf

  (
    n8148_li306_li306,
    n3525_lo_p
  );


  buf

  (
    n8151_li307_li307,
    n3528_lo_p
  );


  buf

  (
    n8154_li308_li308,
    G78_p
  );


  buf

  (
    n8157_li309_li309,
    n3534_lo_p
  );


  buf

  (
    n8160_li310_li310,
    n3537_lo_p
  );


  buf

  (
    n8163_li311_li311,
    n3540_lo_p
  );


  buf

  (
    n8166_li312_li312,
    G79_p
  );


  buf

  (
    n8169_li313_li313,
    n3546_lo_p
  );


  buf

  (
    n8172_li314_li314,
    n3549_lo_p
  );


  buf

  (
    n8175_li315_li315,
    n3552_lo_p
  );


  buf

  (
    n8178_li316_li316,
    G80_p
  );


  buf

  (
    n8181_li317_li317,
    n3558_lo_p
  );


  buf

  (
    n8184_li318_li318,
    n3561_lo_p
  );


  buf

  (
    n8187_li319_li319,
    n3564_lo_p
  );


  buf

  (
    n8190_li320_li320,
    G81_p
  );


  buf

  (
    n8193_li321_li321,
    n3570_lo_p
  );


  buf

  (
    n8196_li322_li322,
    n3573_lo_p
  );


  buf

  (
    n8199_li323_li323,
    n3576_lo_p
  );


  buf

  (
    n8202_li324_li324,
    G82_p
  );


  buf

  (
    n8205_li325_li325,
    n3582_lo_p
  );


  buf

  (
    n8208_li326_li326,
    n3585_lo_p
  );


  buf

  (
    n8211_li327_li327,
    n3588_lo_p
  );


  buf

  (
    n8214_li328_li328,
    G83_p
  );


  buf

  (
    n8217_li329_li329,
    n3594_lo_p
  );


  buf

  (
    n8220_li330_li330,
    n3597_lo_p
  );


  buf

  (
    n8223_li331_li331,
    n3600_lo_p
  );


  buf

  (
    n8226_li332_li332,
    G84_p
  );


  buf

  (
    n8229_li333_li333,
    n3606_lo_p
  );


  buf

  (
    n8232_li334_li334,
    n3609_lo_p
  );


  buf

  (
    n8235_li335_li335,
    n3612_lo_p
  );


  buf

  (
    n8238_li336_li336,
    G85_p
  );


  buf

  (
    n8241_li337_li337,
    n3618_lo_p
  );


  buf

  (
    n8244_li338_li338,
    n3621_lo_p
  );


  buf

  (
    n8247_li339_li339,
    n3624_lo_p
  );


  buf

  (
    n8250_li340_li340,
    G86_p
  );


  buf

  (
    n8253_li341_li341,
    n3630_lo_p
  );


  buf

  (
    n8256_li342_li342,
    n3633_lo_p
  );


  buf

  (
    n8259_li343_li343,
    n3636_lo_p
  );


  buf

  (
    n8262_li344_li344,
    G87_p
  );


  buf

  (
    n8265_li345_li345,
    n3642_lo_p
  );


  buf

  (
    n8268_li346_li346,
    n3645_lo_p
  );


  buf

  (
    n8271_li347_li347,
    n3648_lo_p
  );


  buf

  (
    n8274_li348_li348,
    G88_p
  );


  buf

  (
    n8286_li352_li352,
    G89_p
  );


  buf

  (
    n8370_li380_li380,
    G96_p
  );


  buf

  (
    n8382_li384_li384,
    G97_p
  );


  buf

  (
    n8394_li388_li388,
    G98_p
  );


  buf

  (
    n8406_li392_li392,
    G99_p
  );


  buf

  (
    n8409_li393_li393,
    n3786_lo_p
  );


  buf

  (
    n8412_li394_li394,
    n3789_lo_p
  );


  buf

  (
    n8415_li395_li395,
    n3792_lo_p
  );


  buf

  (
    n8418_li396_li396,
    G100_p
  );


  buf

  (
    n8430_li400_li400,
    G101_p
  );


  buf

  (
    n8442_li404_li404,
    G102_p
  );


  buf

  (
    n8454_li408_li408,
    G103_p
  );


  buf

  (
    n8466_li412_li412,
    G104_p
  );


  buf

  (
    n8550_li440_li440,
    G111_p
  );


  buf

  (
    n8553_li441_li441,
    n3930_lo_p
  );


  buf

  (
    n8556_li442_li442,
    n3933_lo_p
  );


  buf

  (
    n8562_li444_li444,
    G112_p
  );


  buf

  (
    n8565_li445_li445,
    n3942_lo_p
  );


  buf

  (
    n8568_li446_li446,
    n3945_lo_p
  );


  buf

  (
    n8574_li448_li448,
    G113_p
  );


  buf

  (
    n8577_li449_li449,
    n3954_lo_p
  );


  buf

  (
    n8583_li451_li451,
    lo450_buf_o2_p_spl_
  );


  buf

  (
    n8586_li452_li452,
    G114_p
  );


  buf

  (
    n8589_li453_li453,
    n3966_lo_p
  );


  buf

  (
    n8595_li455_li455,
    lo454_buf_o2_p
  );


  buf

  (
    n8598_li456_li456,
    G115_p
  );


  buf

  (
    n8610_li460_li460,
    G116_p
  );


  buf

  (
    n8670_li480_li480,
    G121_p
  );


  buf

  (
    n8682_li484_li484,
    G122_p
  );


  buf

  (
    n8718_li496_li496,
    G125_p
  );


  buf

  (
    n8727_li499_li499,
    n5652_o2_p
  );


  buf

  (
    n8730_li500_li500,
    G126_p
  );


  buf

  (
    n8742_li504_li504,
    G127_p
  );


  buf

  (
    n8751_li507_li507,
    n5601_o2_p
  );


  buf

  (
    n8775_li515_li515,
    n5558_o2_p
  );


  buf

  (
    n8778_li516_li516,
    G130_p
  );


  buf

  (
    n8790_li520_li520,
    G131_p
  );


  buf

  (
    n8799_li523_li523,
    n5654_o2_p
  );


  buf

  (
    n8802_li524_li524,
    G132_p
  );


  buf

  (
    n8805_li525_li525,
    n4182_lo_p
  );


  buf

  (
    n8808_li526_li526,
    n4185_lo_p
  );


  buf

  (
    n8814_li528_li528,
    G133_p
  );


  buf

  (
    n8817_li529_li529,
    n4194_lo_p
  );


  buf

  (
    n8820_li530_li530,
    n4197_lo_p
  );


  buf

  (
    n8826_li532_li532,
    G134_p
  );


  buf

  (
    n8829_li533_li533,
    n4206_lo_p
  );


  buf

  (
    n8832_li534_li534,
    n4209_lo_p
  );


  buf

  (
    n8835_li535_li535,
    n4212_lo_p
  );


  buf

  (
    n8850_li540_li540,
    G136_p
  );


  buf

  (
    n8853_li541_li541,
    n4230_lo_p
  );


  buf

  (
    n8856_li542_li542,
    n4233_lo_p
  );


  buf

  (
    n8859_li543_li543,
    n4236_lo_p
  );


  buf

  (
    n8862_li544_li544,
    G137_p
  );


  buf

  (
    n8874_li548_li548,
    G138_p
  );


  buf

  (
    n8910_li560_li560,
    G141_p
  );


  buf

  (
    n8913_li561_li561,
    n4290_lo_p
  );


  buf

  (
    n8922_li564_li564,
    G142_p
  );


  buf

  (
    n8934_li568_li568,
    G143_p
  );


  buf

  (
    n8970_li580_li580,
    G146_p
  );


  buf

  (
    n8982_li584_li584,
    G147_p
  );


  buf

  (
    n8994_li588_li588,
    G148_p
  );


  buf

  (
    n9006_li592_li592,
    G149_p
  );


  buf

  (
    n9018_li596_li596,
    G150_p
  );


  buf

  (
    n9030_li600_li600,
    G151_p
  );


  buf

  (
    n9033_li601_li601,
    n4410_lo_p
  );


  buf

  (
    n9036_li602_li602,
    n4413_lo_p
  );


  buf

  (
    n9039_li603_li603,
    n4416_lo_p
  );


  buf

  (
    n9042_li604_li604,
    G152_p
  );


  buf

  (
    n9045_li605_li605,
    n4422_lo_p
  );


  buf

  (
    n9048_li606_li606,
    n4425_lo_p
  );


  buf

  (
    n9051_li607_li607,
    n4428_lo_p
  );


  buf

  (
    n9054_li608_li608,
    G153_p
  );


  buf

  (
    n9057_li609_li609,
    n4434_lo_p
  );


  buf

  (
    n9060_li610_li610,
    n4437_lo_p
  );


  buf

  (
    n9063_li611_li611,
    n4440_lo_p
  );


  buf

  (
    n9066_li612_li612,
    G154_p
  );


  buf

  (
    n9069_li613_li613,
    n4446_lo_p
  );


  buf

  (
    n9072_li614_li614,
    n4449_lo_p
  );


  buf

  (
    n9075_li615_li615,
    n4452_lo_p
  );


  buf

  (
    n9078_li616_li616,
    G155_p
  );


  buf

  (
    n9081_li617_li617,
    n4458_lo_p
  );


  buf

  (
    n9084_li618_li618,
    n4461_lo_p
  );


  buf

  (
    n9087_li619_li619,
    n4464_lo_p
  );


  buf

  (
    n9090_li620_li620,
    G156_p
  );


  buf

  (
    n9093_li621_li621,
    n4470_lo_p
  );


  buf

  (
    n9096_li622_li622,
    n4473_lo_p
  );


  buf

  (
    n9099_li623_li623,
    n4476_lo_p
  );


  buf

  (
    n9102_li624_li624,
    G157_p
  );


  buf

  (
    n9105_li625_li625,
    n4482_lo_p
  );


  buf

  (
    n9108_li626_li626,
    n4485_lo_p
  );


  buf

  (
    n9114_li628_li628,
    G158_p
  );


  buf

  (
    n9117_li629_li629,
    n4494_lo_p
  );


  buf

  (
    n9120_li630_li630,
    n4497_lo_p
  );


  buf

  (
    n9123_li631_li631,
    n4500_lo_p
  );


  buf

  (
    n9126_li632_li632,
    G159_p
  );


  buf

  (
    n9129_li633_li633,
    n4506_lo_p
  );


  buf

  (
    n9132_li634_li634,
    n4509_lo_p
  );


  buf

  (
    n9135_li635_li635,
    n4512_lo_p
  );


  buf

  (
    n9138_li636_li636,
    G160_p
  );


  buf

  (
    n9141_li637_li637,
    n4518_lo_p
  );


  buf

  (
    n9144_li638_li638,
    n4521_lo_p
  );


  buf

  (
    n9147_li639_li639,
    n4524_lo_p
  );


  buf

  (
    n9150_li640_li640,
    G161_p
  );


  buf

  (
    n9153_li641_li641,
    n4530_lo_p
  );


  buf

  (
    n9156_li642_li642,
    n4533_lo_p
  );


  buf

  (
    n9159_li643_li643,
    n4536_lo_p
  );


  buf

  (
    n9162_li644_li644,
    G162_p
  );


  buf

  (
    n9165_li645_li645,
    n4542_lo_p
  );


  buf

  (
    n9174_li648_li648,
    G163_p
  );


  buf

  (
    n9177_li649_li649,
    n4554_lo_p
  );


  buf

  (
    n9180_li650_li650,
    n4557_lo_p
  );


  buf

  (
    n9183_li651_li651,
    n4560_lo_p
  );


  buf

  (
    n9186_li652_li652,
    G164_p
  );


  buf

  (
    n9189_li653_li653,
    n4566_lo_p
  );


  buf

  (
    n9192_li654_li654,
    n4569_lo_p
  );


  buf

  (
    n9195_li655_li655,
    n4572_lo_p
  );


  buf

  (
    n9198_li656_li656,
    G165_p
  );


  buf

  (
    n9201_li657_li657,
    n4578_lo_p
  );


  buf

  (
    n9204_li658_li658,
    n4581_lo_p
  );


  buf

  (
    n9207_li659_li659,
    n4584_lo_p
  );


  buf

  (
    n9210_li660_li660,
    G166_p
  );


  buf

  (
    n9213_li661_li661,
    n4590_lo_p
  );


  buf

  (
    n9216_li662_li662,
    n4593_lo_p
  );


  buf

  (
    n9222_li664_li664,
    G167_p
  );


  buf

  (
    n9225_li665_li665,
    n4602_lo_p
  );


  buf

  (
    n9228_li666_li666,
    n4605_lo_p
  );


  buf

  (
    n9234_li668_li668,
    G168_p
  );


  buf

  (
    n9237_li669_li669,
    n4614_lo_p
  );


  buf

  (
    n9240_li670_li670,
    n4617_lo_p
  );


  buf

  (
    n9246_li672_li672,
    G169_p
  );


  buf

  (
    n9249_li673_li673,
    n4626_lo_p
  );


  buf

  (
    n9252_li674_li674,
    n4629_lo_p
  );


  buf

  (
    n9258_li676_li676,
    G170_p
  );


  buf

  (
    n9261_li677_li677,
    n4638_lo_p
  );


  buf

  (
    n9264_li678_li678,
    n4641_lo_p
  );


  buf

  (
    n9267_li679_li679,
    n4644_lo_p
  );


  buf

  (
    n9270_li680_li680,
    G171_p
  );


  buf

  (
    n9273_li681_li681,
    n4650_lo_p
  );


  buf

  (
    n9276_li682_li682,
    n4653_lo_p
  );


  buf

  (
    n9279_li683_li683,
    n4656_lo_p
  );


  buf

  (
    n9282_li684_li684,
    G172_p
  );


  buf

  (
    n9285_li685_li685,
    n4662_lo_p
  );


  buf

  (
    n9288_li686_li686,
    n4665_lo_p
  );


  buf

  (
    n9291_li687_li687,
    n4668_lo_p
  );


  buf

  (
    n9294_li688_li688,
    G173_p
  );


  buf

  (
    n9297_li689_li689,
    n4674_lo_p
  );


  buf

  (
    n9300_li690_li690,
    n4677_lo_p
  );


  buf

  (
    n9303_li691_li691,
    n4680_lo_p
  );


  buf

  (
    n9306_li692_li692,
    G174_p
  );


  buf

  (
    n9309_li693_li693,
    n4686_lo_p
  );


  buf

  (
    n9312_li694_li694,
    n4689_lo_p
  );


  buf

  (
    n9315_li695_li695,
    n4692_lo_p
  );


  buf

  (
    n9318_li696_li696,
    G175_p
  );


  buf

  (
    n9321_li697_li697,
    n4698_lo_p
  );


  buf

  (
    n9324_li698_li698,
    n4701_lo_p
  );


  buf

  (
    n9327_li699_li699,
    n4704_lo_p
  );


  buf

  (
    n9330_li700_li700,
    G176_p
  );


  buf

  (
    n9333_li701_li701,
    n4710_lo_p
  );


  buf

  (
    n9336_li702_li702,
    n4713_lo_p
  );


  buf

  (
    n9339_li703_li703,
    n4716_lo_p_spl_
  );


  buf

  (
    n9342_li704_li704,
    G177_p
  );


  buf

  (
    n9345_li705_li705,
    n4722_lo_p
  );


  buf

  (
    n9348_li706_li706,
    n4725_lo_p
  );


  buf

  (
    n9351_li707_li707,
    n4728_lo_p_spl_11
  );


  buf

  (
    n9354_li708_li708,
    G178_p
  );


  buf

  (
    n9357_li709_li709,
    n4734_lo_p
  );


  buf

  (
    n9360_li710_li710,
    n4737_lo_p
  );


  buf

  (
    n9363_li711_li711,
    n4740_lo_p
  );


  buf

  (
    n4970_i2,
    n1942_inv_p
  );


  buf

  (
    n4972_i2,
    n1948_inv_p
  );


  buf

  (
    n4989_i2,
    n1966_inv_p
  );


  buf

  (
    n5024_i2,
    n1993_inv_p
  );


  buf

  (
    n5025_i2,
    n1996_inv_p
  );


  buf

  (
    n5029_i2,
    n5642_o2_p
  );


  buf

  (
    n5042_i2,
    n2029_inv_p
  );


  buf

  (
    n5048_i2,
    n2041_inv_p
  );


  buf

  (
    n5093_i2,
    n2059_inv_p
  );


  buf

  (
    n5096_i2,
    n2068_inv_p
  );


  buf

  (
    n5193_i2,
    n5915_o2_p
  );


  buf

  (
    n5199_i2,
    n5917_o2_p
  );


  buf

  (
    n5203_i2,
    n2818_o2_p_spl_
  );


  buf

  (
    n5214_i2,
    n2134_inv_p_spl_
  );


  buf

  (
    n5221_i2,
    n2655_o2_p_spl_
  );


  buf

  (
    n5222_i2,
    n2149_inv_p_spl_
  );


  buf

  (
    n5273_i2,
    n2155_inv_p
  );


  buf

  (
    n5365_i2,
    n2182_inv_p
  );


  buf

  (
    n5385_i2,
    n2728_o2_p
  );


  buf

  (
    n5553_i2,
    n2703_o2_p
  );


  buf

  (
    n5636_i2,
    n2870_o2_p
  );


  buf

  (
    n5782_i2,
    n2492_o2_p
  );


  buf

  (
    n5778_i2,
    n2584_inv_p
  );


  buf

  (
    n5323_i2,
    n5908_o2_p_spl_
  );


  buf

  (
    n5325_i2,
    n5910_o2_p_spl_
  );


  buf

  (
    n5327_i2,
    n5912_o2_p_spl_
  );


  buf

  (
    n5329_i2,
    n5914_o2_p_spl_
  );


  buf

  (
    n5816_i2,
    n2617_inv_p_spl_1
  );


  buf

  (
    n5817_i2,
    n2620_inv_p_spl_1
  );


  buf

  (
    n5837_i2,
    n2718_o2_p_spl_
  );


  buf

  (
    n5844_i2,
    n2591_o2_p_spl_
  );


  buf

  (
    n5859_i2,
    n2502_o2_p_spl_
  );


  buf

  (
    n5857_i2,
    n2704_inv_p_spl_
  );


  buf

  (
    n5369_i2,
    n5934_o2_p_spl_
  );


  buf

  (
    n5371_i2,
    n5936_o2_p_spl_
  );


  buf

  (
    n5373_i2,
    n5938_o2_p_spl_
  );


  buf

  (
    n5400_i2,
    lo358_buf_o2_p_spl_
  );


  buf

  (
    n5402_i2,
    lo418_buf_o2_p_spl_
  );


  buf

  (
    n5404_i2,
    lo474_buf_o2_p_spl_
  );


  buf

  (
    n5406_i2,
    lo554_buf_o2_p_spl_
  );


  buf

  (
    n5407_i2,
    lo558_buf_o2_p_spl_
  );


  buf

  (
    n5408_i2,
    lo574_buf_o2_p_spl_
  );


  buf

  (
    n2722_i2,
    g1690_n_spl_
  );


  buf

  (
    n5411_i2,
    n2215_inv_p
  );


  buf

  (
    n5412_i2,
    n2218_inv_p
  );


  buf

  (
    n5413_i2,
    n2221_inv_p
  );


  buf

  (
    n5557_i2,
    lo510_buf_o2_p_spl_
  );


  buf

  (
    n5558_i2,
    lo514_buf_o2_p
  );


  buf

  (
    n5559_i2,
    lo538_buf_o2_p_spl_
  );


  buf

  (
    n5564_i2,
    n2666_o2_p
  );


  buf

  (
    n5565_i2,
    n2667_o2_p
  );


  buf

  (
    n5561_i2,
    n2260_inv_p
  );


  buf

  (
    n5568_i2,
    n2272_inv_p
  );


  buf

  (
    n5598_i2,
    lo410_buf_o2_p_spl_1
  );


  buf

  (
    n5600_i2,
    lo502_buf_o2_p_spl_
  );


  buf

  (
    n5601_i2,
    lo506_buf_o2_p
  );


  buf

  (
    n5602_i2,
    lo550_buf_o2_p_spl_
  );


  buf

  (
    n5603_i2,
    lo570_buf_o2_p_spl_
  );


  buf

  (
    n2853_i2,
    g1692_p_spl_
  );


  buf

  (
    n5637_i2,
    n2317_inv_p_spl_
  );


  buf

  (
    n5627_i2,
    n2302_inv_p
  );


  buf

  (
    n5628_i2,
    n2305_inv_p
  );


  buf

  (
    n5635_i2,
    n2311_inv_p
  );


  buf

  (
    n5640_i2,
    n2689_o2_p_spl_
  );


  buf

  (
    n5641_i2,
    n2323_inv_p_spl_1
  );


  buf

  (
    n5642_i2,
    n2662_o2_p_spl_
  );


  buf

  (
    n5650_i2,
    lo350_buf_o2_p_spl_
  );


  buf

  (
    n5652_i2,
    lo498_buf_o2_p
  );


  buf

  (
    n5653_i2,
    lo518_buf_o2_p_spl_
  );


  buf

  (
    n5654_i2,
    lo522_buf_o2_p
  );


  buf

  (
    n5655_i2,
    lo598_buf_o2_p_spl_
  );


  buf

  (
    n5657_i2,
    n2347_inv_p
  );


  buf

  (
    n5659_i2,
    n2350_inv_p
  );


  buf

  (
    n5661_i2,
    n2353_inv_p_spl_
  );


  buf

  (
    n5656_i2,
    n2344_inv_p
  );


  buf

  (
    n5663_i2,
    n2356_inv_p
  );


  buf

  (
    n5664_i2,
    n2359_inv_p
  );


  buf

  (
    n5795_i2,
    lo546_buf_o2_p_spl_
  );


  buf

  (
    n5796_i2,
    lo590_buf_o2_p_spl_
  );


  buf

  (
    n5797_i2,
    lo594_buf_o2_p_spl_
  );


  buf

  (
    n5739_i2,
    n2476_inv_p
  );


  buf

  (
    n5773_i2,
    n2572_inv_p_spl_1
  );


  buf

  (
    n5798_i2,
    n2602_inv_p
  );


  buf

  (
    n5799_i2,
    n2605_inv_p
  );


  buf

  (
    n5802_i2,
    n2611_inv_p_spl_1
  );


  buf

  (
    n5803_i2,
    n2614_inv_p_spl_
  );


  buf

  (
    n5831_i2,
    lo458_buf_o2_p_spl_
  );


  buf

  (
    n5833_i2,
    lo482_buf_o2_p_spl_1
  );


  buf

  (
    n5820_i2,
    n2629_inv_p_spl_
  );


  buf

  (
    n5823_i2,
    n2638_inv_p_spl_
  );


  buf

  (
    n5824_i2,
    n2641_inv_p_spl_
  );


  buf

  (
    n5869_i2,
    n2740_inv_p_spl_
  );


  buf

  (
    n5848_i2,
    n2686_inv_p
  );


  buf

  (
    n5849_i2,
    n2689_inv_p_spl_1
  );


  buf

  (
    n5856_i2,
    n3031_o2_p
  );


  buf

  (
    n5896_i2,
    lo382_buf_o2_p_spl_1
  );


  not

  (
    n2754_i2,
    g1693_n_spl_
  );


  buf

  (
    n2908_i2,
    g1696_p_spl_
  );


  buf

  (
    n5892_i2,
    n2779_inv_p_spl_1
  );


  buf

  (
    n5915_i2,
    n2653_o2_p_spl_
  );


  buf

  (
    n5919_i2,
    n2682_o2_p_spl_1
  );


  buf

  (
    n5918_i2,
    n2740_o2_p_spl_
  );


  buf

  (
    n5920_i2,
    n2736_o2_p_spl_
  );


  buf

  (
    n5917_i2,
    n2715_o2_p_spl_
  );


  buf

  (
    lo586_buf_i2,
    lo585_buf_o2_p_spl_1
  );


  buf

  (
    n2818_i2,
    g1697_n_spl_
  );


  buf

  (
    n2863_i2,
    g1698_n_spl_1
  );


  buf

  (
    n2721_i2,
    g1699_n_spl_1
  );


  buf

  (
    n2725_i2,
    g1700_n_spl_
  );


  buf

  (
    n3016_i2,
    g1701_n_spl_
  );


  buf

  (
    n3013_i2,
    g1702_n_spl_
  );


  buf

  (
    n2655_i2,
    g1703_p_spl_
  );


  buf

  (
    n2741_i2,
    g1704_p_spl_
  );


  buf

  (
    lo562_buf_i2,
    n4293_lo_p_spl_1
  );


  buf

  (
    n2656_i2,
    g1705_p_spl_
  );


  buf

  (
    n2531_i2,
    g1708_n_spl_
  );


  buf

  (
    n2700_i2,
    g1711_n_spl_
  );


  buf

  (
    n5908_i2,
    lo366_buf_o2_p
  );


  buf

  (
    n5910_i2,
    lo374_buf_o2_p
  );


  buf

  (
    n5912_i2,
    lo426_buf_o2_p
  );


  buf

  (
    n5914_i2,
    lo494_buf_o2_p_spl_11
  );


  buf

  (
    n2753_i2,
    g1712_p_spl_
  );


  buf

  (
    n2878_i2,
    g1714_n_spl_
  );


  buf

  (
    n2836_i2,
    g1716_n_spl_
  );


  buf

  (
    n5934_i2,
    lo434_buf_o2_p_spl_
  );


  buf

  (
    n5936_i2,
    lo466_buf_o2_p_spl_
  );


  buf

  (
    n5938_i2,
    lo490_buf_o2_p_spl_11
  );


  buf

  (
    n2728_i2,
    g1719_p_spl_
  );


  buf

  (
    lo358_buf_i2,
    lo357_buf_o2_p_spl_
  );


  buf

  (
    lo418_buf_i2,
    lo417_buf_o2_p_spl_
  );


  buf

  (
    lo474_buf_i2,
    lo473_buf_o2_p_spl_
  );


  buf

  (
    lo554_buf_i2,
    lo553_buf_o2_p_spl_
  );


  buf

  (
    lo558_buf_i2,
    lo557_buf_o2_p_spl_
  );


  buf

  (
    lo574_buf_i2,
    lo573_buf_o2_p_spl_
  );


  buf

  (
    n2659_i2,
    g1720_n_spl_
  );


  buf

  (
    n2665_i2,
    g1721_n_spl_
  );


  buf

  (
    n2686_i2,
    g1722_n_spl_
  );


  buf

  (
    lo450_buf_i2,
    n3957_lo_p_spl_
  );


  buf

  (
    n2910_i2,
    g1724_p_spl_
  );


  buf

  (
    n2683_i2,
    g1725_p
  );


  not

  (
    n2828_i2,
    g1728_n_spl_
  );


  buf

  (
    n2582_i2,
    g1737_n_spl_
  );


  buf

  (
    n2600_i2,
    g1746_n_spl_
  );


  buf

  (
    n2542_i2,
    g1755_n_spl_
  );


  buf

  (
    n2703_i2,
    g1758_p_spl_
  );


  buf

  (
    lo510_buf_i2,
    lo508_buf_o2_p_spl_
  );


  buf

  (
    lo514_buf_i2,
    lo512_buf_o2_p_spl_
  );


  buf

  (
    lo538_buf_i2,
    lo536_buf_o2_p_spl_
  );


  buf

  (
    lo578_buf_i2,
    lo576_buf_o2_p_spl_
  );


  buf

  (
    n2692_i2,
    g1761_n_spl_
  );


  buf

  (
    n2666_i2,
    g1762_p_spl_
  );


  buf

  (
    n2667_i2,
    g1763_n_spl_1
  );


  buf

  (
    n2660_i2,
    g1764_p_spl_
  );


  buf

  (
    n2744_i2,
    g1767_n_spl_
  );


  buf

  (
    lo454_buf_i2,
    n3969_lo_p_spl_
  );


  buf

  (
    n3593_i2,
    g1768_n_spl_
  );


  buf

  (
    n3048_i2,
    g1774_n_spl_
  );


  buf

  (
    lo410_buf_i2,
    n3834_lo_p_spl_
  );


  buf

  (
    lo502_buf_i2,
    n4110_lo_p_spl_
  );


  buf

  (
    lo506_buf_i2,
    n4122_lo_p_spl_
  );


  buf

  (
    lo550_buf_i2,
    n4254_lo_p_spl_
  );


  buf

  (
    lo570_buf_i2,
    n4314_lo_p_spl_
  );


  buf

  (
    lo582_buf_i2,
    n4350_lo_p_spl_
  );


  buf

  (
    n2646_i2,
    g1777_n_spl_
  );


  buf

  (
    n2673_i2,
    g1780_n_spl_
  );


  not

  (
    n3499_i2,
    g1787_n_spl_
  );


  buf

  (
    n2750_i2,
    g1790_n_spl_
  );


  buf

  (
    n2870_i2,
    g1792_p_spl_
  );


  buf

  (
    n2693_i2,
    g1793_p_spl_
  );


  buf

  (
    n2689_i2,
    g1796_p_spl_
  );


  buf

  (
    n2668_i2,
    g1797_p_spl_
  );


  buf

  (
    n2662_i2,
    g1799_p_spl_
  );


  buf

  (
    lo350_buf_i2,
    n3654_lo_p_spl_
  );


  buf

  (
    lo498_buf_i2,
    n4098_lo_p_spl_
  );


  buf

  (
    lo518_buf_i2,
    n4158_lo_p
  );


  buf

  (
    lo522_buf_i2,
    n4170_lo_p
  );


  buf

  (
    lo598_buf_i2,
    n4398_lo_p_spl_
  );


  buf

  (
    n2708_i2,
    g1802_n_spl_
  );


  buf

  (
    n2674_i2,
    g1803_p_spl_
  );


  buf

  (
    n2647_i2,
    g1804_p_spl_
  );


  buf

  (
    n2751_i2,
    g1805_p_spl_
  );


  buf

  (
    n2747_i2,
    g1808_p_spl_
  );


  buf

  (
    n2669_i2,
    g1809_p_spl_
  );


  buf

  (
    n2872_i2,
    g1810_p
  );


  buf

  (
    n3313_i2,
    g1811_p
  );


  buf

  (
    n3273_i2,
    g1812_p
  );


  buf

  (
    n2848_i2,
    g1813_n
  );


  buf

  (
    n2893_i2,
    g1814_n
  );


  buf

  (
    n3267_i2,
    g1815_p
  );


  buf

  (
    n2925_i2,
    g1816_p
  );


  buf

  (
    n2839_i2,
    g1817_n
  );


  buf

  (
    n2831_i2,
    g1818_n
  );


  buf

  (
    n2558_i2,
    g1822_p
  );


  buf

  (
    n2562_i2,
    g1826_p
  );


  buf

  (
    n2825_i2,
    g1827_p
  );


  buf

  (
    n3263_i2,
    g1829_p
  );


  buf

  (
    n3517_i2,
    g1847_p
  );


  not

  (
    n2873_i2,
    g1848_n
  );


  not

  (
    n2926_i2,
    g1849_n
  );


  buf

  (
    n3261_i2,
    g1850_p
  );


  buf

  (
    n3268_i2,
    g1851_p
  );


  buf

  (
    n3274_i2,
    g1852_p
  );


  not

  (
    n3314_i2,
    g1853_n
  );


  buf

  (
    n3571_i2,
    g1868_p
  );


  buf

  (
    n2950_i2,
    g1869_p
  );


  buf

  (
    n2951_i2,
    g1870_p
  );


  buf

  (
    n3022_i2,
    g1873_p
  );


  buf

  (
    n3023_i2,
    g1874_p
  );


  not

  (
    n3057_i2,
    g1878_n
  );


  not

  (
    n3058_i2,
    g1879_p
  );


  buf

  (
    n2931_i2,
    g1880_n
  );


  buf

  (
    n2911_i2,
    g1881_n
  );


  buf

  (
    n2959_i2,
    g1885_n
  );


  buf

  (
    n2960_i2,
    g1886_p
  );


  buf

  (
    n2922_i2,
    g1887_n
  );


  buf

  (
    n2888_i2,
    g1888_p
  );


  buf

  (
    n2889_i2,
    g1889_n
  );


  not

  (
    n3051_i2,
    g1892_p
  );


  not

  (
    n3052_i2,
    g1893_n
  );


  not

  (
    n3063_i2,
    g1894_n
  );


  buf

  (
    n2845_i2,
    g1897_p
  );


  buf

  (
    n2737_i2,
    g1898_n_spl_
  );


  buf

  (
    n3281_i2,
    g1901_n
  );


  buf

  (
    n3294_i2,
    g1904_n
  );


  not

  (
    n2885_i2,
    g1907_p
  );


  buf

  (
    n2786_i2,
    g1910_p
  );


  buf

  (
    n2783_i2,
    g1913_n
  );


  buf

  (
    n2801_i2,
    g1916_n
  );


  buf

  (
    n2572_i2,
    g1925_n
  );


  buf

  (
    n2628_i2,
    g1934_n
  );


  buf

  (
    n2609_i2,
    g1943_n
  );


  buf

  (
    n2618_i2,
    g1952_n
  );


  buf

  (
    n2637_i2,
    g1961_n
  );


  buf

  (
    n2525_i2,
    g1970_n
  );


  buf

  (
    n2551_i2,
    g1979_n
  );


  buf

  (
    n3759_i2,
    g2001_p
  );


  buf

  (
    n2994_i2,
    g2004_n
  );


  buf

  (
    n3040_i2,
    g2007_p
  );


  buf

  (
    n2943_i2,
    g2011_p
  );


  buf

  (
    n2991_i2,
    g2017_p
  );


  buf

  (
    n3034_i2,
    g2020_n
  );


  buf

  (
    n2881_i2,
    g2023_p
  );


  buf

  (
    n3021_i2,
    g2029_n
  );


  buf

  (
    n3062_i2,
    g2032_n
  );


  buf

  (
    n2763_i2,
    g2039_p
  );


  not

  (
    n2764_i2,
    g2040_n
  );


  buf

  (
    n2775_i2,
    g2050_p
  );


  not

  (
    n2776_i2,
    g2051_n
  );


  buf

  (
    n2968_i2,
    g2058_n
  );


  buf

  (
    n2969_i2,
    g2059_p
  );


  buf

  (
    n2798_i2,
    g2068_p
  );


  buf

  (
    n3661_i2,
    g2095_p
  );


  buf

  (
    n2694_i2,
    g2096_n_spl_
  );


  buf

  (
    n2809_i2,
    g2098_n_spl_
  );


  buf

  (
    n2817_i2,
    g2099_p_spl_
  );


  buf

  (
    n2514_i2,
    g2108_n_spl_
  );


  buf

  (
    n2501_i2,
    g2117_n_spl_
  );


  not

  (
    n2528_i2,
    g2120_n_spl_
  );


  not

  (
    n2505_i2,
    g2123_n_spl_
  );


  buf

  (
    n2492_i2,
    g2126_p_spl_
  );


  buf

  (
    lo546_buf_i2,
    n4242_lo_p_spl_
  );


  buf

  (
    lo590_buf_i2,
    n4374_lo_p_spl_
  );


  buf

  (
    lo594_buf_i2,
    n4386_lo_p_spl_
  );


  buf

  (
    n2679_i2,
    g2129_n_spl_
  );


  buf

  (
    n2733_i2,
    g2132_n_spl_
  );


  not

  (
    n2709_i2,
    g2133_n_spl_
  );


  buf

  (
    n2676_i2,
    g2135_p_spl_
  );


  buf

  (
    n2649_i2,
    g2137_p_spl_1
  );


  buf

  (
    n2815_i2,
    g2141_n
  );


  not

  (
    n2704_i2,
    g2143_n
  );


  not

  (
    n3590_i2,
    g2158_p
  );


  not

  (
    n3591_i2,
    g2159_n
  );


  buf

  (
    n2752_i2,
    g2160_n_spl_
  );


  buf

  (
    n3638_i2,
    g2173_p
  );


  buf

  (
    n3639_i2,
    g2174_n
  );


  buf

  (
    n2695_i2,
    g2175_p_spl_
  );


  buf

  (
    n3047_i2,
    g2177_n_spl_
  );


  buf

  (
    lo458_buf_i2,
    n3978_lo_p_spl_
  );


  buf

  (
    lo482_buf_i2,
    n4050_lo_p_spl_
  );


  buf

  (
    lo566_buf_i2,
    n4302_lo_p_spl_
  );


  buf

  (
    n2718_i2,
    g2180_n
  );


  buf

  (
    n3707_i2,
    g2189_n
  );


  buf

  (
    n3671_i2,
    g2198_n
  );


  buf

  (
    n3680_i2,
    g2207_n
  );


  buf

  (
    n3749_i2,
    g2216_n
  );


  buf

  (
    n3716_i2,
    g2225_n
  );


  buf

  (
    n3692_i2,
    g2234_n
  );


  buf

  (
    n2591_i2,
    g2243_n
  );


  buf

  (
    n3478_i2,
    g2249_n
  );


  not

  (
    n3610_i2,
    g2260_n
  );


  not

  (
    n3611_i2,
    g2261_p
  );


  buf

  (
    n2652_i2,
    g2264_n_spl_
  );


  not

  (
    n2714_i2,
    g2267_p_spl_
  );


  not

  (
    n2738_i2,
    g2268_n_spl_
  );


  buf

  (
    n3616_i2,
    g2273_n
  );


  buf

  (
    n3617_i2,
    g2274_p
  );


  buf

  (
    n3031_i2,
    g2276_n_spl_
  );


  buf

  (
    n2515_i2,
    g2277_p
  );


  not

  (
    n3562_i2,
    g2278_n
  );


  buf

  (
    n2502_i2,
    g2279_p
  );


  buf

  (
    n3560_i2,
    g2280_n
  );


  not

  (
    n3554_i2,
    g2296_n
  );


  buf

  (
    n3555_i2,
    g2297_p
  );


  not

  (
    n3536_i2,
    g2316_n
  );


  buf

  (
    n3537_i2,
    g2317_p
  );


  not

  (
    n3508_i2,
    g2325_n
  );


  buf

  (
    n3650_i2,
    g2333_p
  );


  buf

  (
    n3740_i2,
    g2354_n
  );


  buf

  (
    n3484_i2,
    g2360_n
  );


  not

  (
    n2680_i2,
    g2361_n_spl_
  );


  not

  (
    n2734_i2,
    g2362_n_spl_
  );


  buf

  (
    n2735_i2,
    g2363_n_spl_
  );


  buf

  (
    n2711_i2,
    g2365_p_spl_
  );


  buf

  (
    lo585_buf_i2,
    n4362_lo_p
  );


  buf

  (
    n2719_i2,
    g2366_p
  );


  buf

  (
    n2720_i2,
    g2367_p
  );


  buf

  (
    n2723_i2,
    g2368_p
  );


  buf

  (
    n2724_i2,
    g2369_p
  );


  buf

  (
    n3624_i2,
    g2370_p
  );


  buf

  (
    n3625_i2,
    g2371_n
  );


  buf

  (
    n3015_i2,
    g2372_p
  );


  buf

  (
    n3491_i2,
    g2373_p
  );


  buf

  (
    n2696_i2,
    g2374_p
  );


  buf

  (
    n2811_i2,
    g2376_n
  );


  buf

  (
    n3010_i2,
    g2378_n
  );


  buf

  (
    n3012_i2,
    g2379_p
  );


  buf

  (
    lo382_buf_i2,
    n3750_lo_p
  );


  buf

  (
    lo386_buf_i2,
    n3762_lo_p
  );


  buf

  (
    lo390_buf_i2,
    n3774_lo_p
  );


  buf

  (
    lo398_buf_i2,
    n3798_lo_p
  );


  buf

  (
    lo402_buf_i2,
    n3810_lo_p
  );


  buf

  (
    lo406_buf_i2,
    n3822_lo_p
  );


  buf

  (
    n3492_i2,
    g2380_n
  );


  buf

  (
    lo366_buf_i2,
    G92_p_spl_
  );


  buf

  (
    lo374_buf_i2,
    G94_p_spl_
  );


  buf

  (
    lo426_buf_i2,
    G107_p_spl_
  );


  buf

  (
    lo494_buf_i2,
    G124_p_spl_1
  );


  buf

  (
    n2653_i2,
    g2381_p
  );


  buf

  (
    n2654_i2,
    g2382_n
  );


  buf

  (
    n2715_i2,
    g2383_p
  );


  buf

  (
    n2740_i2,
    g2385_p
  );


  buf

  (
    n2682_i2,
    g2387_p
  );


  buf

  (
    n2736_i2,
    g2388_p
  );


  buf

  (
    lo508_buf_i2,
    G128_p
  );


  buf

  (
    lo512_buf_i2,
    G129_p
  );


  buf

  (
    lo536_buf_i2,
    G135_p
  );


  buf

  (
    lo576_buf_i2,
    G145_p
  );


  buf

  (
    lo357_buf_i2,
    G90_p
  );


  buf

  (
    lo361_buf_i2,
    G91_p
  );


  buf

  (
    lo417_buf_i2,
    G105_p
  );


  buf

  (
    lo421_buf_i2,
    G106_p
  );


  buf

  (
    lo473_buf_i2,
    G119_p
  );


  buf

  (
    lo477_buf_i2,
    G120_p
  );


  buf

  (
    lo553_buf_i2,
    G139_p
  );


  buf

  (
    lo557_buf_i2,
    G140_p
  );


  buf

  (
    lo573_buf_i2,
    G144_p
  );


  buf

  (
    lo434_buf_i2,
    G109_p
  );


  buf

  (
    lo438_buf_i2,
    G110_p
  );


  buf

  (
    lo466_buf_i2,
    G117_p
  );


  buf

  (
    lo470_buf_i2,
    G118_p
  );


  buf

  (
    lo490_buf_i2,
    G123_p
  );


  buf

  (
    n2657_i2,
    g2389_p
  );


  buf

  (
    n2658_i2,
    g2390_p
  );


  buf

  (
    n2663_i2,
    g2391_p
  );


  buf

  (
    n2664_i2,
    g2392_p
  );


  buf

  (
    n2684_i2,
    g2393_p
  );


  buf

  (
    n2685_i2,
    g2394_p
  );


  buf

  (
    n4443_lo_n_spl_,
    n4443_lo_n
  );


  buf

  (
    n4479_lo_n_spl_,
    n4479_lo_n
  );


  buf

  (
    n3399_lo_p_spl_,
    n3399_lo_p
  );


  buf

  (
    n3399_lo_p_spl_0,
    n3399_lo_p_spl_
  );


  buf

  (
    n3399_lo_p_spl_00,
    n3399_lo_p_spl_0
  );


  buf

  (
    n3399_lo_p_spl_01,
    n3399_lo_p_spl_0
  );


  buf

  (
    n3399_lo_p_spl_1,
    n3399_lo_p_spl_
  );


  buf

  (
    n2619_lo_p_spl_,
    n2619_lo_p
  );


  buf

  (
    n4587_lo_n_spl_,
    n4587_lo_n
  );


  buf

  (
    n2739_lo_n_spl_,
    n2739_lo_n
  );


  buf

  (
    g1055_n_spl_,
    g1055_n
  );


  buf

  (
    g1055_n_spl_0,
    g1055_n_spl_
  );


  buf

  (
    g1055_n_spl_00,
    g1055_n_spl_0
  );


  buf

  (
    g1055_n_spl_000,
    g1055_n_spl_00
  );


  buf

  (
    g1055_n_spl_01,
    g1055_n_spl_0
  );


  buf

  (
    g1055_n_spl_1,
    g1055_n_spl_
  );


  buf

  (
    g1055_n_spl_10,
    g1055_n_spl_1
  );


  buf

  (
    g1055_n_spl_11,
    g1055_n_spl_1
  );


  buf

  (
    n4563_lo_n_spl_,
    n4563_lo_n
  );


  buf

  (
    n4563_lo_n_spl_0,
    n4563_lo_n_spl_
  );


  buf

  (
    n4563_lo_n_spl_00,
    n4563_lo_n_spl_0
  );


  buf

  (
    n4563_lo_n_spl_01,
    n4563_lo_n_spl_0
  );


  buf

  (
    n4563_lo_n_spl_1,
    n4563_lo_n_spl_
  );


  buf

  (
    n4563_lo_p_spl_,
    n4563_lo_p
  );


  buf

  (
    n4563_lo_p_spl_0,
    n4563_lo_p_spl_
  );


  buf

  (
    n4563_lo_p_spl_00,
    n4563_lo_p_spl_0
  );


  buf

  (
    n4563_lo_p_spl_01,
    n4563_lo_p_spl_0
  );


  buf

  (
    n4563_lo_p_spl_1,
    n4563_lo_p_spl_
  );


  buf

  (
    n2551_o2_p_spl_,
    n2551_o2_p
  );


  buf

  (
    g1094_n_spl_,
    g1094_n
  );


  buf

  (
    n5273_o2_n_spl_,
    n5273_o2_n
  );


  buf

  (
    g1101_n_spl_,
    g1101_n
  );


  buf

  (
    n2786_o2_p_spl_,
    n2786_o2_p
  );


  buf

  (
    n2783_o2_p_spl_,
    n2783_o2_p
  );


  buf

  (
    n2786_o2_n_spl_,
    n2786_o2_n
  );


  buf

  (
    n2783_o2_n_spl_,
    n2783_o2_n
  );


  buf

  (
    n2801_o2_n_spl_,
    n2801_o2_n
  );


  buf

  (
    n2798_o2_n_spl_,
    n2798_o2_n
  );


  buf

  (
    n2801_o2_p_spl_,
    n2801_o2_p
  );


  buf

  (
    n2798_o2_p_spl_,
    n2798_o2_p
  );


  buf

  (
    n5837_o2_p_spl_,
    n5837_o2_p
  );


  buf

  (
    n5837_o2_p_spl_0,
    n5837_o2_p_spl_
  );


  buf

  (
    n2825_o2_p_spl_,
    n2825_o2_p
  );


  buf

  (
    n2825_o2_p_spl_0,
    n2825_o2_p_spl_
  );


  buf

  (
    n2825_o2_p_spl_00,
    n2825_o2_p_spl_0
  );


  buf

  (
    n2825_o2_p_spl_000,
    n2825_o2_p_spl_00
  );


  buf

  (
    n2825_o2_p_spl_001,
    n2825_o2_p_spl_00
  );


  buf

  (
    n2825_o2_p_spl_01,
    n2825_o2_p_spl_0
  );


  buf

  (
    n2825_o2_p_spl_010,
    n2825_o2_p_spl_01
  );


  buf

  (
    n2825_o2_p_spl_011,
    n2825_o2_p_spl_01
  );


  buf

  (
    n2825_o2_p_spl_1,
    n2825_o2_p_spl_
  );


  buf

  (
    n2825_o2_p_spl_10,
    n2825_o2_p_spl_1
  );


  buf

  (
    n2825_o2_p_spl_100,
    n2825_o2_p_spl_10
  );


  buf

  (
    n2825_o2_p_spl_101,
    n2825_o2_p_spl_10
  );


  buf

  (
    n2825_o2_p_spl_11,
    n2825_o2_p_spl_1
  );


  buf

  (
    n2825_o2_p_spl_110,
    n2825_o2_p_spl_11
  );


  buf

  (
    n2825_o2_p_spl_111,
    n2825_o2_p_spl_11
  );


  buf

  (
    n4731_lo_n_spl_,
    n4731_lo_n
  );


  buf

  (
    n4731_lo_n_spl_0,
    n4731_lo_n_spl_
  );


  buf

  (
    n4731_lo_n_spl_00,
    n4731_lo_n_spl_0
  );


  buf

  (
    n4731_lo_n_spl_000,
    n4731_lo_n_spl_00
  );


  buf

  (
    n4731_lo_n_spl_01,
    n4731_lo_n_spl_0
  );


  buf

  (
    n4731_lo_n_spl_1,
    n4731_lo_n_spl_
  );


  buf

  (
    n4731_lo_n_spl_10,
    n4731_lo_n_spl_1
  );


  buf

  (
    n4731_lo_n_spl_11,
    n4731_lo_n_spl_1
  );


  buf

  (
    n4719_lo_p_spl_,
    n4719_lo_p
  );


  buf

  (
    n4719_lo_p_spl_0,
    n4719_lo_p_spl_
  );


  buf

  (
    n4719_lo_p_spl_00,
    n4719_lo_p_spl_0
  );


  buf

  (
    n4719_lo_p_spl_000,
    n4719_lo_p_spl_00
  );


  buf

  (
    n4719_lo_p_spl_001,
    n4719_lo_p_spl_00
  );


  buf

  (
    n4719_lo_p_spl_01,
    n4719_lo_p_spl_0
  );


  buf

  (
    n4719_lo_p_spl_010,
    n4719_lo_p_spl_01
  );


  buf

  (
    n4719_lo_p_spl_011,
    n4719_lo_p_spl_01
  );


  buf

  (
    n4719_lo_p_spl_1,
    n4719_lo_p_spl_
  );


  buf

  (
    n4719_lo_p_spl_10,
    n4719_lo_p_spl_1
  );


  buf

  (
    n4719_lo_p_spl_100,
    n4719_lo_p_spl_10
  );


  buf

  (
    n4719_lo_p_spl_101,
    n4719_lo_p_spl_10
  );


  buf

  (
    n4719_lo_p_spl_11,
    n4719_lo_p_spl_1
  );


  buf

  (
    n4719_lo_p_spl_110,
    n4719_lo_p_spl_11
  );


  buf

  (
    n2825_o2_n_spl_,
    n2825_o2_n
  );


  buf

  (
    n4731_lo_p_spl_,
    n4731_lo_p
  );


  buf

  (
    n4731_lo_p_spl_0,
    n4731_lo_p_spl_
  );


  buf

  (
    n4731_lo_p_spl_00,
    n4731_lo_p_spl_0
  );


  buf

  (
    n4731_lo_p_spl_000,
    n4731_lo_p_spl_00
  );


  buf

  (
    n4731_lo_p_spl_01,
    n4731_lo_p_spl_0
  );


  buf

  (
    n4731_lo_p_spl_1,
    n4731_lo_p_spl_
  );


  buf

  (
    n4731_lo_p_spl_10,
    n4731_lo_p_spl_1
  );


  buf

  (
    n4731_lo_p_spl_11,
    n4731_lo_p_spl_1
  );


  buf

  (
    n4719_lo_n_spl_,
    n4719_lo_n
  );


  buf

  (
    n4719_lo_n_spl_0,
    n4719_lo_n_spl_
  );


  buf

  (
    n4719_lo_n_spl_1,
    n4719_lo_n_spl_
  );


  buf

  (
    n2845_o2_p_spl_,
    n2845_o2_p
  );


  buf

  (
    n4683_lo_n_spl_,
    n4683_lo_n
  );


  buf

  (
    n4683_lo_n_spl_0,
    n4683_lo_n_spl_
  );


  buf

  (
    n4683_lo_n_spl_00,
    n4683_lo_n_spl_0
  );


  buf

  (
    n4683_lo_n_spl_000,
    n4683_lo_n_spl_00
  );


  buf

  (
    n4683_lo_n_spl_0000,
    n4683_lo_n_spl_000
  );


  buf

  (
    n4683_lo_n_spl_0001,
    n4683_lo_n_spl_000
  );


  buf

  (
    n4683_lo_n_spl_001,
    n4683_lo_n_spl_00
  );


  buf

  (
    n4683_lo_n_spl_0010,
    n4683_lo_n_spl_001
  );


  buf

  (
    n4683_lo_n_spl_0011,
    n4683_lo_n_spl_001
  );


  buf

  (
    n4683_lo_n_spl_01,
    n4683_lo_n_spl_0
  );


  buf

  (
    n4683_lo_n_spl_010,
    n4683_lo_n_spl_01
  );


  buf

  (
    n4683_lo_n_spl_011,
    n4683_lo_n_spl_01
  );


  buf

  (
    n4683_lo_n_spl_1,
    n4683_lo_n_spl_
  );


  buf

  (
    n4683_lo_n_spl_10,
    n4683_lo_n_spl_1
  );


  buf

  (
    n4683_lo_n_spl_100,
    n4683_lo_n_spl_10
  );


  buf

  (
    n4683_lo_n_spl_101,
    n4683_lo_n_spl_10
  );


  buf

  (
    n4683_lo_n_spl_11,
    n4683_lo_n_spl_1
  );


  buf

  (
    n4683_lo_n_spl_110,
    n4683_lo_n_spl_11
  );


  buf

  (
    n4683_lo_n_spl_111,
    n4683_lo_n_spl_11
  );


  buf

  (
    g1132_n_spl_,
    g1132_n
  );


  buf

  (
    g1132_n_spl_0,
    g1132_n_spl_
  );


  buf

  (
    g1132_n_spl_00,
    g1132_n_spl_0
  );


  buf

  (
    g1132_n_spl_1,
    g1132_n_spl_
  );


  buf

  (
    n4683_lo_p_spl_,
    n4683_lo_p
  );


  buf

  (
    n4683_lo_p_spl_0,
    n4683_lo_p_spl_
  );


  buf

  (
    n4683_lo_p_spl_00,
    n4683_lo_p_spl_0
  );


  buf

  (
    n4683_lo_p_spl_000,
    n4683_lo_p_spl_00
  );


  buf

  (
    n4683_lo_p_spl_0000,
    n4683_lo_p_spl_000
  );


  buf

  (
    n4683_lo_p_spl_0001,
    n4683_lo_p_spl_000
  );


  buf

  (
    n4683_lo_p_spl_001,
    n4683_lo_p_spl_00
  );


  buf

  (
    n4683_lo_p_spl_0010,
    n4683_lo_p_spl_001
  );


  buf

  (
    n4683_lo_p_spl_0011,
    n4683_lo_p_spl_001
  );


  buf

  (
    n4683_lo_p_spl_01,
    n4683_lo_p_spl_0
  );


  buf

  (
    n4683_lo_p_spl_010,
    n4683_lo_p_spl_01
  );


  buf

  (
    n4683_lo_p_spl_011,
    n4683_lo_p_spl_01
  );


  buf

  (
    n4683_lo_p_spl_1,
    n4683_lo_p_spl_
  );


  buf

  (
    n4683_lo_p_spl_10,
    n4683_lo_p_spl_1
  );


  buf

  (
    n4683_lo_p_spl_100,
    n4683_lo_p_spl_10
  );


  buf

  (
    n4683_lo_p_spl_101,
    n4683_lo_p_spl_10
  );


  buf

  (
    n4683_lo_p_spl_11,
    n4683_lo_p_spl_1
  );


  buf

  (
    n4683_lo_p_spl_110,
    n4683_lo_p_spl_11
  );


  buf

  (
    n4683_lo_p_spl_111,
    n4683_lo_p_spl_11
  );


  buf

  (
    g1142_n_spl_,
    g1142_n
  );


  buf

  (
    g1142_n_spl_0,
    g1142_n_spl_
  );


  buf

  (
    g1142_n_spl_00,
    g1142_n_spl_0
  );


  buf

  (
    g1142_n_spl_1,
    g1142_n_spl_
  );


  buf

  (
    n4671_lo_p_spl_,
    n4671_lo_p
  );


  buf

  (
    n4671_lo_p_spl_0,
    n4671_lo_p_spl_
  );


  buf

  (
    n4671_lo_p_spl_00,
    n4671_lo_p_spl_0
  );


  buf

  (
    n4671_lo_p_spl_000,
    n4671_lo_p_spl_00
  );


  buf

  (
    n4671_lo_p_spl_001,
    n4671_lo_p_spl_00
  );


  buf

  (
    n4671_lo_p_spl_01,
    n4671_lo_p_spl_0
  );


  buf

  (
    n4671_lo_p_spl_1,
    n4671_lo_p_spl_
  );


  buf

  (
    n4671_lo_p_spl_10,
    n4671_lo_p_spl_1
  );


  buf

  (
    n4671_lo_p_spl_11,
    n4671_lo_p_spl_1
  );


  buf

  (
    n2643_lo_p_spl_,
    n2643_lo_p
  );


  buf

  (
    n2871_lo_p_spl_,
    n2871_lo_p
  );


  buf

  (
    n4671_lo_n_spl_,
    n4671_lo_n
  );


  buf

  (
    n4671_lo_n_spl_0,
    n4671_lo_n_spl_
  );


  buf

  (
    n4671_lo_n_spl_00,
    n4671_lo_n_spl_0
  );


  buf

  (
    n4671_lo_n_spl_000,
    n4671_lo_n_spl_00
  );


  buf

  (
    n4671_lo_n_spl_001,
    n4671_lo_n_spl_00
  );


  buf

  (
    n4671_lo_n_spl_01,
    n4671_lo_n_spl_0
  );


  buf

  (
    n4671_lo_n_spl_1,
    n4671_lo_n_spl_
  );


  buf

  (
    n4671_lo_n_spl_10,
    n4671_lo_n_spl_1
  );


  buf

  (
    n4671_lo_n_spl_11,
    n4671_lo_n_spl_1
  );


  buf

  (
    n5636_o2_n_spl_,
    n5636_o2_n
  );


  buf

  (
    n2881_o2_n_spl_,
    n2881_o2_n
  );


  buf

  (
    g1159_n_spl_,
    g1159_n
  );


  buf

  (
    n4695_lo_n_spl_,
    n4695_lo_n
  );


  buf

  (
    n4695_lo_n_spl_0,
    n4695_lo_n_spl_
  );


  buf

  (
    n4695_lo_n_spl_00,
    n4695_lo_n_spl_0
  );


  buf

  (
    n4695_lo_n_spl_000,
    n4695_lo_n_spl_00
  );


  buf

  (
    n4695_lo_n_spl_0000,
    n4695_lo_n_spl_000
  );


  buf

  (
    n4695_lo_n_spl_0001,
    n4695_lo_n_spl_000
  );


  buf

  (
    n4695_lo_n_spl_001,
    n4695_lo_n_spl_00
  );


  buf

  (
    n4695_lo_n_spl_0010,
    n4695_lo_n_spl_001
  );


  buf

  (
    n4695_lo_n_spl_0011,
    n4695_lo_n_spl_001
  );


  buf

  (
    n4695_lo_n_spl_01,
    n4695_lo_n_spl_0
  );


  buf

  (
    n4695_lo_n_spl_010,
    n4695_lo_n_spl_01
  );


  buf

  (
    n4695_lo_n_spl_011,
    n4695_lo_n_spl_01
  );


  buf

  (
    n4695_lo_n_spl_1,
    n4695_lo_n_spl_
  );


  buf

  (
    n4695_lo_n_spl_10,
    n4695_lo_n_spl_1
  );


  buf

  (
    n4695_lo_n_spl_100,
    n4695_lo_n_spl_10
  );


  buf

  (
    n4695_lo_n_spl_101,
    n4695_lo_n_spl_10
  );


  buf

  (
    n4695_lo_n_spl_11,
    n4695_lo_n_spl_1
  );


  buf

  (
    n4695_lo_n_spl_110,
    n4695_lo_n_spl_11
  );


  buf

  (
    n4695_lo_n_spl_111,
    n4695_lo_n_spl_11
  );


  buf

  (
    n4695_lo_p_spl_,
    n4695_lo_p
  );


  buf

  (
    n4695_lo_p_spl_0,
    n4695_lo_p_spl_
  );


  buf

  (
    n4695_lo_p_spl_00,
    n4695_lo_p_spl_0
  );


  buf

  (
    n4695_lo_p_spl_000,
    n4695_lo_p_spl_00
  );


  buf

  (
    n4695_lo_p_spl_0000,
    n4695_lo_p_spl_000
  );


  buf

  (
    n4695_lo_p_spl_0001,
    n4695_lo_p_spl_000
  );


  buf

  (
    n4695_lo_p_spl_001,
    n4695_lo_p_spl_00
  );


  buf

  (
    n4695_lo_p_spl_0010,
    n4695_lo_p_spl_001
  );


  buf

  (
    n4695_lo_p_spl_0011,
    n4695_lo_p_spl_001
  );


  buf

  (
    n4695_lo_p_spl_01,
    n4695_lo_p_spl_0
  );


  buf

  (
    n4695_lo_p_spl_010,
    n4695_lo_p_spl_01
  );


  buf

  (
    n4695_lo_p_spl_011,
    n4695_lo_p_spl_01
  );


  buf

  (
    n4695_lo_p_spl_1,
    n4695_lo_p_spl_
  );


  buf

  (
    n4695_lo_p_spl_10,
    n4695_lo_p_spl_1
  );


  buf

  (
    n4695_lo_p_spl_100,
    n4695_lo_p_spl_10
  );


  buf

  (
    n4695_lo_p_spl_101,
    n4695_lo_p_spl_10
  );


  buf

  (
    n4695_lo_p_spl_11,
    n4695_lo_p_spl_1
  );


  buf

  (
    n4695_lo_p_spl_110,
    n4695_lo_p_spl_11
  );


  buf

  (
    n4695_lo_p_spl_111,
    n4695_lo_p_spl_11
  );


  buf

  (
    n4707_lo_p_spl_,
    n4707_lo_p
  );


  buf

  (
    n4707_lo_p_spl_0,
    n4707_lo_p_spl_
  );


  buf

  (
    n4707_lo_p_spl_00,
    n4707_lo_p_spl_0
  );


  buf

  (
    n4707_lo_p_spl_000,
    n4707_lo_p_spl_00
  );


  buf

  (
    n4707_lo_p_spl_001,
    n4707_lo_p_spl_00
  );


  buf

  (
    n4707_lo_p_spl_01,
    n4707_lo_p_spl_0
  );


  buf

  (
    n4707_lo_p_spl_1,
    n4707_lo_p_spl_
  );


  buf

  (
    n4707_lo_p_spl_10,
    n4707_lo_p_spl_1
  );


  buf

  (
    n4707_lo_p_spl_11,
    n4707_lo_p_spl_1
  );


  buf

  (
    n4707_lo_n_spl_,
    n4707_lo_n
  );


  buf

  (
    n4707_lo_n_spl_0,
    n4707_lo_n_spl_
  );


  buf

  (
    n4707_lo_n_spl_00,
    n4707_lo_n_spl_0
  );


  buf

  (
    n4707_lo_n_spl_000,
    n4707_lo_n_spl_00
  );


  buf

  (
    n4707_lo_n_spl_001,
    n4707_lo_n_spl_00
  );


  buf

  (
    n4707_lo_n_spl_01,
    n4707_lo_n_spl_0
  );


  buf

  (
    n4707_lo_n_spl_1,
    n4707_lo_n_spl_
  );


  buf

  (
    n4707_lo_n_spl_10,
    n4707_lo_n_spl_1
  );


  buf

  (
    n4707_lo_n_spl_11,
    n4707_lo_n_spl_1
  );


  buf

  (
    g1176_n_spl_,
    g1176_n
  );


  buf

  (
    g1183_n_spl_,
    g1183_n
  );


  buf

  (
    g1188_n_spl_,
    g1188_n
  );


  buf

  (
    n2853_o2_n_spl_,
    n2853_o2_n
  );


  buf

  (
    n2853_o2_n_spl_0,
    n2853_o2_n_spl_
  );


  buf

  (
    n2853_o2_n_spl_00,
    n2853_o2_n_spl_0
  );


  buf

  (
    n2853_o2_n_spl_1,
    n2853_o2_n_spl_
  );


  buf

  (
    g1201_n_spl_,
    g1201_n
  );


  buf

  (
    n2853_o2_p_spl_,
    n2853_o2_p
  );


  buf

  (
    n2853_o2_p_spl_0,
    n2853_o2_p_spl_
  );


  buf

  (
    n2853_o2_p_spl_1,
    n2853_o2_p_spl_
  );


  buf

  (
    g1201_p_spl_,
    g1201_p
  );


  buf

  (
    g1205_p_spl_,
    g1205_p
  );


  buf

  (
    g1206_n_spl_,
    g1206_n
  );


  buf

  (
    g1205_n_spl_,
    g1205_n
  );


  buf

  (
    g1206_p_spl_,
    g1206_p
  );


  buf

  (
    n4972_o2_n_spl_,
    n4972_o2_n
  );


  buf

  (
    n4989_o2_p_spl_,
    n4989_o2_p
  );


  buf

  (
    n4972_o2_p_spl_,
    n4972_o2_p
  );


  buf

  (
    n4989_o2_n_spl_,
    n4989_o2_n
  );


  buf

  (
    n5025_o2_n_spl_,
    n5025_o2_n
  );


  buf

  (
    n5093_o2_p_spl_,
    n5093_o2_p
  );


  buf

  (
    n5025_o2_p_spl_,
    n5025_o2_p
  );


  buf

  (
    n5093_o2_n_spl_,
    n5093_o2_n
  );


  buf

  (
    g1215_n_spl_,
    g1215_n
  );


  buf

  (
    g1218_p_spl_,
    g1218_p
  );


  buf

  (
    g1215_p_spl_,
    g1215_p
  );


  buf

  (
    g1218_n_spl_,
    g1218_n
  );


  buf

  (
    n2994_o2_n_spl_,
    n2994_o2_n
  );


  buf

  (
    n2991_o2_p_spl_,
    n2991_o2_p
  );


  buf

  (
    n2994_o2_p_spl_,
    n2994_o2_p
  );


  buf

  (
    n2991_o2_n_spl_,
    n2991_o2_n
  );


  buf

  (
    n4970_o2_p_spl_,
    n4970_o2_p
  );


  buf

  (
    n5024_o2_n_spl_,
    n5024_o2_n
  );


  buf

  (
    n4970_o2_n_spl_,
    n4970_o2_n
  );


  buf

  (
    n5024_o2_p_spl_,
    n5024_o2_p
  );


  buf

  (
    g1224_n_spl_,
    g1224_n
  );


  buf

  (
    g1227_p_spl_,
    g1227_p
  );


  buf

  (
    g1224_p_spl_,
    g1224_p
  );


  buf

  (
    g1227_n_spl_,
    g1227_n
  );


  buf

  (
    g1234_n_spl_,
    g1234_n
  );


  buf

  (
    n3021_o2_n_spl_,
    n3021_o2_n
  );


  buf

  (
    g1243_p_spl_,
    g1243_p
  );


  buf

  (
    g1246_p_spl_,
    g1246_p
  );


  buf

  (
    n3062_o2_p_spl_,
    n3062_o2_p
  );


  buf

  (
    g1250_p_spl_,
    g1250_p
  );


  buf

  (
    g1249_p_spl_,
    g1249_p
  );


  buf

  (
    n4503_lo_n_spl_,
    n4503_lo_n
  );


  buf

  (
    n4503_lo_n_spl_0,
    n4503_lo_n_spl_
  );


  buf

  (
    n4503_lo_n_spl_00,
    n4503_lo_n_spl_0
  );


  buf

  (
    n4503_lo_n_spl_000,
    n4503_lo_n_spl_00
  );


  buf

  (
    n4503_lo_n_spl_0000,
    n4503_lo_n_spl_000
  );


  buf

  (
    n4503_lo_n_spl_0001,
    n4503_lo_n_spl_000
  );


  buf

  (
    n4503_lo_n_spl_001,
    n4503_lo_n_spl_00
  );


  buf

  (
    n4503_lo_n_spl_0010,
    n4503_lo_n_spl_001
  );


  buf

  (
    n4503_lo_n_spl_0011,
    n4503_lo_n_spl_001
  );


  buf

  (
    n4503_lo_n_spl_01,
    n4503_lo_n_spl_0
  );


  buf

  (
    n4503_lo_n_spl_010,
    n4503_lo_n_spl_01
  );


  buf

  (
    n4503_lo_n_spl_011,
    n4503_lo_n_spl_01
  );


  buf

  (
    n4503_lo_n_spl_1,
    n4503_lo_n_spl_
  );


  buf

  (
    n4503_lo_n_spl_10,
    n4503_lo_n_spl_1
  );


  buf

  (
    n4503_lo_n_spl_100,
    n4503_lo_n_spl_10
  );


  buf

  (
    n4503_lo_n_spl_101,
    n4503_lo_n_spl_10
  );


  buf

  (
    n4503_lo_n_spl_11,
    n4503_lo_n_spl_1
  );


  buf

  (
    n4503_lo_n_spl_110,
    n4503_lo_n_spl_11
  );


  buf

  (
    n4503_lo_n_spl_111,
    n4503_lo_n_spl_11
  );


  buf

  (
    n4503_lo_p_spl_,
    n4503_lo_p
  );


  buf

  (
    n4503_lo_p_spl_0,
    n4503_lo_p_spl_
  );


  buf

  (
    n4503_lo_p_spl_00,
    n4503_lo_p_spl_0
  );


  buf

  (
    n4503_lo_p_spl_000,
    n4503_lo_p_spl_00
  );


  buf

  (
    n4503_lo_p_spl_0000,
    n4503_lo_p_spl_000
  );


  buf

  (
    n4503_lo_p_spl_0001,
    n4503_lo_p_spl_000
  );


  buf

  (
    n4503_lo_p_spl_001,
    n4503_lo_p_spl_00
  );


  buf

  (
    n4503_lo_p_spl_0010,
    n4503_lo_p_spl_001
  );


  buf

  (
    n4503_lo_p_spl_0011,
    n4503_lo_p_spl_001
  );


  buf

  (
    n4503_lo_p_spl_01,
    n4503_lo_p_spl_0
  );


  buf

  (
    n4503_lo_p_spl_010,
    n4503_lo_p_spl_01
  );


  buf

  (
    n4503_lo_p_spl_011,
    n4503_lo_p_spl_01
  );


  buf

  (
    n4503_lo_p_spl_1,
    n4503_lo_p_spl_
  );


  buf

  (
    n4503_lo_p_spl_10,
    n4503_lo_p_spl_1
  );


  buf

  (
    n4503_lo_p_spl_100,
    n4503_lo_p_spl_10
  );


  buf

  (
    n4503_lo_p_spl_101,
    n4503_lo_p_spl_10
  );


  buf

  (
    n4503_lo_p_spl_11,
    n4503_lo_p_spl_1
  );


  buf

  (
    n4503_lo_p_spl_110,
    n4503_lo_p_spl_11
  );


  buf

  (
    n4503_lo_p_spl_111,
    n4503_lo_p_spl_11
  );


  buf

  (
    n4515_lo_n_spl_,
    n4515_lo_n
  );


  buf

  (
    n4515_lo_n_spl_0,
    n4515_lo_n_spl_
  );


  buf

  (
    n4515_lo_n_spl_00,
    n4515_lo_n_spl_0
  );


  buf

  (
    n4515_lo_n_spl_000,
    n4515_lo_n_spl_00
  );


  buf

  (
    n4515_lo_n_spl_001,
    n4515_lo_n_spl_00
  );


  buf

  (
    n4515_lo_n_spl_01,
    n4515_lo_n_spl_0
  );


  buf

  (
    n4515_lo_n_spl_1,
    n4515_lo_n_spl_
  );


  buf

  (
    n4515_lo_n_spl_10,
    n4515_lo_n_spl_1
  );


  buf

  (
    n4515_lo_n_spl_11,
    n4515_lo_n_spl_1
  );


  buf

  (
    n3579_lo_p_spl_,
    n3579_lo_p
  );


  buf

  (
    n3567_lo_p_spl_,
    n3567_lo_p
  );


  buf

  (
    n4515_lo_p_spl_,
    n4515_lo_p
  );


  buf

  (
    n4515_lo_p_spl_0,
    n4515_lo_p_spl_
  );


  buf

  (
    n4515_lo_p_spl_00,
    n4515_lo_p_spl_0
  );


  buf

  (
    n4515_lo_p_spl_000,
    n4515_lo_p_spl_00
  );


  buf

  (
    n4515_lo_p_spl_001,
    n4515_lo_p_spl_00
  );


  buf

  (
    n4515_lo_p_spl_01,
    n4515_lo_p_spl_0
  );


  buf

  (
    n4515_lo_p_spl_1,
    n4515_lo_p_spl_
  );


  buf

  (
    n4515_lo_p_spl_10,
    n4515_lo_p_spl_1
  );


  buf

  (
    n4515_lo_p_spl_11,
    n4515_lo_p_spl_1
  );


  buf

  (
    n3375_lo_p_spl_,
    n3375_lo_p
  );


  buf

  (
    n3375_lo_p_spl_0,
    n3375_lo_p_spl_
  );


  buf

  (
    n3375_lo_p_spl_00,
    n3375_lo_p_spl_0
  );


  buf

  (
    n3375_lo_p_spl_000,
    n3375_lo_p_spl_00
  );


  buf

  (
    n3375_lo_p_spl_0000,
    n3375_lo_p_spl_000
  );


  buf

  (
    n3375_lo_p_spl_001,
    n3375_lo_p_spl_00
  );


  buf

  (
    n3375_lo_p_spl_01,
    n3375_lo_p_spl_0
  );


  buf

  (
    n3375_lo_p_spl_010,
    n3375_lo_p_spl_01
  );


  buf

  (
    n3375_lo_p_spl_011,
    n3375_lo_p_spl_01
  );


  buf

  (
    n3375_lo_p_spl_1,
    n3375_lo_p_spl_
  );


  buf

  (
    n3375_lo_p_spl_10,
    n3375_lo_p_spl_1
  );


  buf

  (
    n3375_lo_p_spl_100,
    n3375_lo_p_spl_10
  );


  buf

  (
    n3375_lo_p_spl_101,
    n3375_lo_p_spl_10
  );


  buf

  (
    n3375_lo_p_spl_11,
    n3375_lo_p_spl_1
  );


  buf

  (
    n3375_lo_p_spl_110,
    n3375_lo_p_spl_11
  );


  buf

  (
    n3375_lo_p_spl_111,
    n3375_lo_p_spl_11
  );


  buf

  (
    n4527_lo_n_spl_,
    n4527_lo_n
  );


  buf

  (
    n4527_lo_n_spl_0,
    n4527_lo_n_spl_
  );


  buf

  (
    n4527_lo_n_spl_00,
    n4527_lo_n_spl_0
  );


  buf

  (
    n4527_lo_n_spl_000,
    n4527_lo_n_spl_00
  );


  buf

  (
    n4527_lo_n_spl_0000,
    n4527_lo_n_spl_000
  );


  buf

  (
    n4527_lo_n_spl_0001,
    n4527_lo_n_spl_000
  );


  buf

  (
    n4527_lo_n_spl_001,
    n4527_lo_n_spl_00
  );


  buf

  (
    n4527_lo_n_spl_0010,
    n4527_lo_n_spl_001
  );


  buf

  (
    n4527_lo_n_spl_0011,
    n4527_lo_n_spl_001
  );


  buf

  (
    n4527_lo_n_spl_01,
    n4527_lo_n_spl_0
  );


  buf

  (
    n4527_lo_n_spl_010,
    n4527_lo_n_spl_01
  );


  buf

  (
    n4527_lo_n_spl_011,
    n4527_lo_n_spl_01
  );


  buf

  (
    n4527_lo_n_spl_1,
    n4527_lo_n_spl_
  );


  buf

  (
    n4527_lo_n_spl_10,
    n4527_lo_n_spl_1
  );


  buf

  (
    n4527_lo_n_spl_100,
    n4527_lo_n_spl_10
  );


  buf

  (
    n4527_lo_n_spl_101,
    n4527_lo_n_spl_10
  );


  buf

  (
    n4527_lo_n_spl_11,
    n4527_lo_n_spl_1
  );


  buf

  (
    n4527_lo_n_spl_110,
    n4527_lo_n_spl_11
  );


  buf

  (
    n4527_lo_n_spl_111,
    n4527_lo_n_spl_11
  );


  buf

  (
    n4527_lo_p_spl_,
    n4527_lo_p
  );


  buf

  (
    n4527_lo_p_spl_0,
    n4527_lo_p_spl_
  );


  buf

  (
    n4527_lo_p_spl_00,
    n4527_lo_p_spl_0
  );


  buf

  (
    n4527_lo_p_spl_000,
    n4527_lo_p_spl_00
  );


  buf

  (
    n4527_lo_p_spl_0000,
    n4527_lo_p_spl_000
  );


  buf

  (
    n4527_lo_p_spl_0001,
    n4527_lo_p_spl_000
  );


  buf

  (
    n4527_lo_p_spl_001,
    n4527_lo_p_spl_00
  );


  buf

  (
    n4527_lo_p_spl_0010,
    n4527_lo_p_spl_001
  );


  buf

  (
    n4527_lo_p_spl_0011,
    n4527_lo_p_spl_001
  );


  buf

  (
    n4527_lo_p_spl_01,
    n4527_lo_p_spl_0
  );


  buf

  (
    n4527_lo_p_spl_010,
    n4527_lo_p_spl_01
  );


  buf

  (
    n4527_lo_p_spl_011,
    n4527_lo_p_spl_01
  );


  buf

  (
    n4527_lo_p_spl_1,
    n4527_lo_p_spl_
  );


  buf

  (
    n4527_lo_p_spl_10,
    n4527_lo_p_spl_1
  );


  buf

  (
    n4527_lo_p_spl_100,
    n4527_lo_p_spl_10
  );


  buf

  (
    n4527_lo_p_spl_101,
    n4527_lo_p_spl_10
  );


  buf

  (
    n4527_lo_p_spl_11,
    n4527_lo_p_spl_1
  );


  buf

  (
    n4527_lo_p_spl_110,
    n4527_lo_p_spl_11
  );


  buf

  (
    n4527_lo_p_spl_111,
    n4527_lo_p_spl_11
  );


  buf

  (
    n4539_lo_n_spl_,
    n4539_lo_n
  );


  buf

  (
    n4539_lo_n_spl_0,
    n4539_lo_n_spl_
  );


  buf

  (
    n4539_lo_n_spl_00,
    n4539_lo_n_spl_0
  );


  buf

  (
    n4539_lo_n_spl_000,
    n4539_lo_n_spl_00
  );


  buf

  (
    n4539_lo_n_spl_001,
    n4539_lo_n_spl_00
  );


  buf

  (
    n4539_lo_n_spl_01,
    n4539_lo_n_spl_0
  );


  buf

  (
    n4539_lo_n_spl_1,
    n4539_lo_n_spl_
  );


  buf

  (
    n4539_lo_n_spl_10,
    n4539_lo_n_spl_1
  );


  buf

  (
    n4539_lo_n_spl_11,
    n4539_lo_n_spl_1
  );


  buf

  (
    n4539_lo_p_spl_,
    n4539_lo_p
  );


  buf

  (
    n4539_lo_p_spl_0,
    n4539_lo_p_spl_
  );


  buf

  (
    n4539_lo_p_spl_00,
    n4539_lo_p_spl_0
  );


  buf

  (
    n4539_lo_p_spl_000,
    n4539_lo_p_spl_00
  );


  buf

  (
    n4539_lo_p_spl_001,
    n4539_lo_p_spl_00
  );


  buf

  (
    n4539_lo_p_spl_01,
    n4539_lo_p_spl_0
  );


  buf

  (
    n4539_lo_p_spl_1,
    n4539_lo_p_spl_
  );


  buf

  (
    n4539_lo_p_spl_10,
    n4539_lo_p_spl_1
  );


  buf

  (
    n4539_lo_p_spl_11,
    n4539_lo_p_spl_1
  );


  buf

  (
    n2775_lo_p_spl_,
    n2775_lo_p
  );


  buf

  (
    n2799_lo_p_spl_,
    n2799_lo_p
  );


  buf

  (
    g1182_n_spl_,
    g1182_n
  );


  buf

  (
    g1182_n_spl_0,
    g1182_n_spl_
  );


  buf

  (
    g1182_n_spl_00,
    g1182_n_spl_0
  );


  buf

  (
    g1182_n_spl_1,
    g1182_n_spl_
  );


  buf

  (
    g1155_n_spl_,
    g1155_n
  );


  buf

  (
    g1155_n_spl_0,
    g1155_n_spl_
  );


  buf

  (
    g1155_n_spl_00,
    g1155_n_spl_0
  );


  buf

  (
    g1155_n_spl_1,
    g1155_n_spl_
  );


  buf

  (
    n2679_lo_p_spl_,
    n2679_lo_p
  );


  buf

  (
    n2931_lo_p_spl_,
    n2931_lo_p
  );


  buf

  (
    g1187_n_spl_,
    g1187_n
  );


  buf

  (
    g1187_n_spl_0,
    g1187_n_spl_
  );


  buf

  (
    g1187_n_spl_00,
    g1187_n_spl_0
  );


  buf

  (
    g1187_n_spl_1,
    g1187_n_spl_
  );


  buf

  (
    g1158_n_spl_,
    g1158_n
  );


  buf

  (
    g1158_n_spl_0,
    g1158_n_spl_
  );


  buf

  (
    g1158_n_spl_00,
    g1158_n_spl_0
  );


  buf

  (
    g1158_n_spl_1,
    g1158_n_spl_
  );


  buf

  (
    n2667_lo_p_spl_,
    n2667_lo_p
  );


  buf

  (
    n2919_lo_p_spl_,
    n2919_lo_p
  );


  buf

  (
    g1194_n_spl_,
    g1194_n
  );


  buf

  (
    g1194_n_spl_0,
    g1194_n_spl_
  );


  buf

  (
    g1194_n_spl_00,
    g1194_n_spl_0
  );


  buf

  (
    g1194_n_spl_1,
    g1194_n_spl_
  );


  buf

  (
    g1164_n_spl_,
    g1164_n
  );


  buf

  (
    g1164_n_spl_0,
    g1164_n_spl_
  );


  buf

  (
    g1164_n_spl_00,
    g1164_n_spl_0
  );


  buf

  (
    g1164_n_spl_1,
    g1164_n_spl_
  );


  buf

  (
    n2907_lo_n_spl_,
    n2907_lo_n
  );


  buf

  (
    n2895_lo_n_spl_,
    n2895_lo_n
  );


  buf

  (
    g1200_p_spl_,
    g1200_p
  );


  buf

  (
    g1200_p_spl_0,
    g1200_p_spl_
  );


  buf

  (
    g1200_p_spl_00,
    g1200_p_spl_0
  );


  buf

  (
    g1200_p_spl_1,
    g1200_p_spl_
  );


  buf

  (
    g1137_p_spl_,
    g1137_p
  );


  buf

  (
    g1137_p_spl_0,
    g1137_p_spl_
  );


  buf

  (
    g1137_p_spl_00,
    g1137_p_spl_0
  );


  buf

  (
    g1137_p_spl_1,
    g1137_p_spl_
  );


  buf

  (
    n3519_lo_p_spl_,
    n3519_lo_p
  );


  buf

  (
    n3639_lo_p_spl_,
    n3639_lo_p
  );


  buf

  (
    n3471_lo_n_spl_,
    n3471_lo_n
  );


  buf

  (
    n3591_lo_n_spl_,
    n3591_lo_n
  );


  buf

  (
    n3375_lo_n_spl_,
    n3375_lo_n
  );


  buf

  (
    n3375_lo_n_spl_0,
    n3375_lo_n_spl_
  );


  buf

  (
    n3375_lo_n_spl_1,
    n3375_lo_n_spl_
  );


  buf

  (
    n3447_lo_p_spl_,
    n3447_lo_p
  );


  buf

  (
    n3459_lo_p_spl_,
    n3459_lo_p
  );


  buf

  (
    n3423_lo_p_spl_,
    n3423_lo_p
  );


  buf

  (
    n3435_lo_p_spl_,
    n3435_lo_p
  );


  buf

  (
    n4659_lo_n_spl_,
    n4659_lo_n
  );


  buf

  (
    n4659_lo_p_spl_,
    n4659_lo_p
  );


  buf

  (
    n3339_lo_n_spl_,
    n3339_lo_n
  );


  buf

  (
    n3339_lo_p_spl_,
    n3339_lo_p
  );


  buf

  (
    n5837_o2_n_spl_,
    n5837_o2_n
  );


  buf

  (
    g1437_n_spl_,
    g1437_n
  );


  buf

  (
    n3795_lo_n_spl_,
    n3795_lo_n
  );


  buf

  (
    n4467_lo_n_spl_,
    n4467_lo_n
  );


  buf

  (
    g1049_n_spl_,
    g1049_n
  );


  buf

  (
    g1054_n_spl_,
    g1054_n
  );


  buf

  (
    g1111_n_spl_,
    g1111_n
  );


  buf

  (
    g1120_n_spl_,
    g1120_n
  );


  buf

  (
    g1212_n_spl_,
    g1212_n
  );


  buf

  (
    g1233_n_spl_,
    g1233_n
  );


  buf

  (
    n3099_lo_p_spl_,
    n3099_lo_p
  );


  buf

  (
    n3111_lo_p_spl_,
    n3111_lo_p
  );


  buf

  (
    g1470_n_spl_,
    g1470_n
  );


  buf

  (
    g1470_n_spl_0,
    g1470_n_spl_
  );


  buf

  (
    g1470_n_spl_00,
    g1470_n_spl_0
  );


  buf

  (
    g1470_n_spl_1,
    g1470_n_spl_
  );


  buf

  (
    g1449_n_spl_,
    g1449_n
  );


  buf

  (
    g1449_n_spl_0,
    g1449_n_spl_
  );


  buf

  (
    g1449_n_spl_00,
    g1449_n_spl_0
  );


  buf

  (
    g1449_n_spl_1,
    g1449_n_spl_
  );


  buf

  (
    n2823_lo_p_spl_,
    n2823_lo_p
  );


  buf

  (
    n2811_lo_p_spl_,
    n2811_lo_p
  );


  buf

  (
    g1476_n_spl_,
    g1476_n
  );


  buf

  (
    g1476_n_spl_0,
    g1476_n_spl_
  );


  buf

  (
    g1476_n_spl_00,
    g1476_n_spl_0
  );


  buf

  (
    g1476_n_spl_1,
    g1476_n_spl_
  );


  buf

  (
    g1453_n_spl_,
    g1453_n
  );


  buf

  (
    g1453_n_spl_0,
    g1453_n_spl_
  );


  buf

  (
    g1453_n_spl_00,
    g1453_n_spl_0
  );


  buf

  (
    g1453_n_spl_1,
    g1453_n_spl_
  );


  buf

  (
    n3087_lo_p_spl_,
    n3087_lo_p
  );


  buf

  (
    n3075_lo_p_spl_,
    n3075_lo_p
  );


  buf

  (
    g1482_n_spl_,
    g1482_n
  );


  buf

  (
    g1482_n_spl_0,
    g1482_n_spl_
  );


  buf

  (
    g1482_n_spl_00,
    g1482_n_spl_0
  );


  buf

  (
    g1482_n_spl_1,
    g1482_n_spl_
  );


  buf

  (
    g1457_n_spl_,
    g1457_n
  );


  buf

  (
    g1457_n_spl_0,
    g1457_n_spl_
  );


  buf

  (
    g1457_n_spl_00,
    g1457_n_spl_0
  );


  buf

  (
    g1457_n_spl_1,
    g1457_n_spl_
  );


  buf

  (
    n2787_lo_p_spl_,
    n2787_lo_p
  );


  buf

  (
    n3039_lo_p_spl_,
    n3039_lo_p
  );


  buf

  (
    g1486_n_spl_,
    g1486_n
  );


  buf

  (
    g1486_n_spl_0,
    g1486_n_spl_
  );


  buf

  (
    g1486_n_spl_00,
    g1486_n_spl_0
  );


  buf

  (
    g1486_n_spl_1,
    g1486_n_spl_
  );


  buf

  (
    g1460_n_spl_,
    g1460_n
  );


  buf

  (
    g1460_n_spl_0,
    g1460_n_spl_
  );


  buf

  (
    g1460_n_spl_00,
    g1460_n_spl_0
  );


  buf

  (
    g1460_n_spl_1,
    g1460_n_spl_
  );


  buf

  (
    n3531_lo_p_spl_,
    n3531_lo_p
  );


  buf

  (
    n3651_lo_p_spl_,
    n3651_lo_p
  );


  buf

  (
    n3507_lo_p_spl_,
    n3507_lo_p
  );


  buf

  (
    n3627_lo_p_spl_,
    n3627_lo_p
  );


  buf

  (
    n3495_lo_p_spl_,
    n3495_lo_p
  );


  buf

  (
    n3615_lo_p_spl_,
    n3615_lo_p
  );


  buf

  (
    n3483_lo_p_spl_,
    n3483_lo_p
  );


  buf

  (
    n3603_lo_p_spl_,
    n3603_lo_p
  );


  buf

  (
    g1640_n_spl_,
    g1640_n
  );


  buf

  (
    g1639_n_spl_,
    g1639_n
  );


  buf

  (
    g1645_n_spl_,
    g1645_n
  );


  buf

  (
    n2883_lo_n_spl_,
    n2883_lo_n
  );


  buf

  (
    n2655_lo_n_spl_,
    n2655_lo_n
  );


  buf

  (
    g1653_p_spl_,
    g1653_p
  );


  buf

  (
    g1653_p_spl_0,
    g1653_p_spl_
  );


  buf

  (
    g1653_p_spl_1,
    g1653_p_spl_
  );


  buf

  (
    g1656_p_spl_,
    g1656_p
  );


  buf

  (
    g1656_p_spl_0,
    g1656_p_spl_
  );


  buf

  (
    g1656_p_spl_1,
    g1656_p_spl_
  );


  buf

  (
    n3555_lo_n_spl_,
    n3555_lo_n
  );


  buf

  (
    n3543_lo_n_spl_,
    n3543_lo_n
  );


  buf

  (
    n2134_inv_n_spl_,
    n2134_inv_n
  );


  buf

  (
    n2134_inv_n_spl_0,
    n2134_inv_n_spl_
  );


  buf

  (
    n2134_inv_n_spl_1,
    n2134_inv_n_spl_
  );


  buf

  (
    n2718_o2_n_spl_,
    n2718_o2_n
  );


  buf

  (
    n2134_inv_p_spl_,
    n2134_inv_p
  );


  buf

  (
    n2134_inv_p_spl_0,
    n2134_inv_p_spl_
  );


  buf

  (
    n2718_o2_p_spl_,
    n2718_o2_p
  );


  buf

  (
    n2718_o2_p_spl_0,
    n2718_o2_p_spl_
  );


  buf

  (
    g1690_n_spl_,
    g1690_n
  );


  buf

  (
    n5663_o2_n_spl_,
    n5663_o2_n
  );


  buf

  (
    n5663_o2_n_spl_0,
    n5663_o2_n_spl_
  );


  buf

  (
    n5663_o2_n_spl_00,
    n5663_o2_n_spl_0
  );


  buf

  (
    n5663_o2_n_spl_1,
    n5663_o2_n_spl_
  );


  buf

  (
    n2753_o2_n_spl_,
    n2753_o2_n
  );


  buf

  (
    n2628_lo_p_spl_,
    n2628_lo_p
  );


  buf

  (
    n2628_lo_p_spl_0,
    n2628_lo_p_spl_
  );


  buf

  (
    n2628_lo_p_spl_1,
    n2628_lo_p_spl_
  );


  buf

  (
    n5802_o2_p_spl_,
    n5802_o2_p
  );


  buf

  (
    g1695_n_spl_,
    g1695_n
  );


  buf

  (
    n2715_o2_n_spl_,
    n2715_o2_n
  );


  buf

  (
    n2715_o2_p_spl_,
    n2715_o2_p
  );


  buf

  (
    n2715_o2_p_spl_0,
    n2715_o2_p_spl_
  );


  buf

  (
    n3010_o2_n_spl_,
    n3010_o2_n
  );


  buf

  (
    n3010_o2_p_spl_,
    n3010_o2_p
  );


  buf

  (
    n2653_o2_p_spl_,
    n2653_o2_p
  );


  buf

  (
    n2740_o2_p_spl_,
    n2740_o2_p
  );


  buf

  (
    n2740_o2_p_spl_0,
    n2740_o2_p_spl_
  );


  buf

  (
    n2736_o2_p_spl_,
    n2736_o2_p
  );


  buf

  (
    n2740_o2_n_spl_,
    n2740_o2_n
  );


  buf

  (
    n2614_inv_p_spl_,
    n2614_inv_p
  );


  buf

  (
    n2614_inv_p_spl_0,
    n2614_inv_p_spl_
  );


  buf

  (
    g1703_p_spl_,
    g1703_p
  );


  buf

  (
    g1703_p_spl_0,
    g1703_p_spl_
  );


  buf

  (
    n2614_inv_n_spl_,
    n2614_inv_n
  );


  buf

  (
    g1703_n_spl_,
    g1703_n
  );


  buf

  (
    n4632_lo_n_spl_,
    n4632_lo_n
  );


  buf

  (
    n4632_lo_n_spl_0,
    n4632_lo_n_spl_
  );


  buf

  (
    n4632_lo_n_spl_00,
    n4632_lo_n_spl_0
  );


  buf

  (
    n4632_lo_n_spl_000,
    n4632_lo_n_spl_00
  );


  buf

  (
    n4632_lo_n_spl_001,
    n4632_lo_n_spl_00
  );


  buf

  (
    n4632_lo_n_spl_01,
    n4632_lo_n_spl_0
  );


  buf

  (
    n4632_lo_n_spl_010,
    n4632_lo_n_spl_01
  );


  buf

  (
    n4632_lo_n_spl_011,
    n4632_lo_n_spl_01
  );


  buf

  (
    n4632_lo_n_spl_1,
    n4632_lo_n_spl_
  );


  buf

  (
    n4632_lo_n_spl_10,
    n4632_lo_n_spl_1
  );


  buf

  (
    n4632_lo_n_spl_11,
    n4632_lo_n_spl_1
  );


  buf

  (
    n4596_lo_p_spl_,
    n4596_lo_p
  );


  buf

  (
    n4596_lo_p_spl_0,
    n4596_lo_p_spl_
  );


  buf

  (
    n4596_lo_p_spl_00,
    n4596_lo_p_spl_0
  );


  buf

  (
    n4596_lo_p_spl_000,
    n4596_lo_p_spl_00
  );


  buf

  (
    n4596_lo_p_spl_001,
    n4596_lo_p_spl_00
  );


  buf

  (
    n4596_lo_p_spl_01,
    n4596_lo_p_spl_0
  );


  buf

  (
    n4596_lo_p_spl_010,
    n4596_lo_p_spl_01
  );


  buf

  (
    n4596_lo_p_spl_011,
    n4596_lo_p_spl_01
  );


  buf

  (
    n4596_lo_p_spl_1,
    n4596_lo_p_spl_
  );


  buf

  (
    n4596_lo_p_spl_10,
    n4596_lo_p_spl_1
  );


  buf

  (
    n4596_lo_p_spl_11,
    n4596_lo_p_spl_1
  );


  buf

  (
    n5914_o2_p_spl_,
    n5914_o2_p
  );


  buf

  (
    n5914_o2_p_spl_0,
    n5914_o2_p_spl_
  );


  buf

  (
    lo382_buf_o2_p_spl_,
    lo382_buf_o2_p
  );


  buf

  (
    lo382_buf_o2_p_spl_0,
    lo382_buf_o2_p_spl_
  );


  buf

  (
    lo382_buf_o2_p_spl_00,
    lo382_buf_o2_p_spl_0
  );


  buf

  (
    lo382_buf_o2_p_spl_01,
    lo382_buf_o2_p_spl_0
  );


  buf

  (
    lo382_buf_o2_p_spl_1,
    lo382_buf_o2_p_spl_
  );


  buf

  (
    n5914_o2_n_spl_,
    n5914_o2_n
  );


  buf

  (
    lo382_buf_o2_n_spl_,
    lo382_buf_o2_n
  );


  buf

  (
    lo382_buf_o2_n_spl_0,
    lo382_buf_o2_n_spl_
  );


  buf

  (
    lo382_buf_o2_n_spl_00,
    lo382_buf_o2_n_spl_0
  );


  buf

  (
    lo382_buf_o2_n_spl_1,
    lo382_buf_o2_n_spl_
  );


  buf

  (
    n2629_inv_p_spl_,
    n2629_inv_p
  );


  buf

  (
    n2353_inv_p_spl_,
    n2353_inv_p
  );


  buf

  (
    g1698_n_spl_,
    g1698_n
  );


  buf

  (
    g1698_n_spl_0,
    g1698_n_spl_
  );


  buf

  (
    g1698_n_spl_1,
    g1698_n_spl_
  );


  buf

  (
    g1698_p_spl_,
    g1698_p
  );


  buf

  (
    g1698_p_spl_0,
    g1698_p_spl_
  );


  buf

  (
    n2734_o2_n_spl_,
    n2734_o2_n
  );


  buf

  (
    n2734_o2_p_spl_,
    n2734_o2_p
  );


  buf

  (
    n2689_inv_p_spl_,
    n2689_inv_p
  );


  buf

  (
    n2689_inv_p_spl_0,
    n2689_inv_p_spl_
  );


  buf

  (
    n2689_inv_p_spl_1,
    n2689_inv_p_spl_
  );


  buf

  (
    n2711_o2_n_spl_,
    n2711_o2_n
  );


  buf

  (
    n2689_inv_n_spl_,
    n2689_inv_n
  );


  buf

  (
    n2689_inv_n_spl_0,
    n2689_inv_n_spl_
  );


  buf

  (
    n2711_o2_p_spl_,
    n2711_o2_p
  );


  buf

  (
    lo585_buf_o2_p_spl_,
    lo585_buf_o2_p
  );


  buf

  (
    lo585_buf_o2_p_spl_0,
    lo585_buf_o2_p_spl_
  );


  buf

  (
    lo585_buf_o2_p_spl_00,
    lo585_buf_o2_p_spl_0
  );


  buf

  (
    lo585_buf_o2_p_spl_1,
    lo585_buf_o2_p_spl_
  );


  buf

  (
    g1700_n_spl_,
    g1700_n
  );


  buf

  (
    g1700_n_spl_0,
    g1700_n_spl_
  );


  buf

  (
    lo585_buf_o2_n_spl_,
    lo585_buf_o2_n
  );


  buf

  (
    lo585_buf_o2_n_spl_0,
    lo585_buf_o2_n_spl_
  );


  buf

  (
    lo585_buf_o2_n_spl_1,
    lo585_buf_o2_n_spl_
  );


  buf

  (
    g1700_p_spl_,
    g1700_p
  );


  buf

  (
    g1717_n_spl_,
    g1717_n
  );


  buf

  (
    g1717_p_spl_,
    g1717_p
  );


  buf

  (
    g1696_p_spl_,
    g1696_p
  );


  buf

  (
    n5919_o2_p_spl_,
    n5919_o2_p
  );


  buf

  (
    g1723_n_spl_,
    g1723_n
  );


  buf

  (
    n2611_inv_p_spl_,
    n2611_inv_p
  );


  buf

  (
    n2611_inv_p_spl_0,
    n2611_inv_p_spl_
  );


  buf

  (
    n2611_inv_p_spl_1,
    n2611_inv_p_spl_
  );


  buf

  (
    n2682_o2_p_spl_,
    n2682_o2_p
  );


  buf

  (
    n2682_o2_p_spl_0,
    n2682_o2_p_spl_
  );


  buf

  (
    n2682_o2_p_spl_1,
    n2682_o2_p_spl_
  );


  buf

  (
    n2611_inv_n_spl_,
    n2611_inv_n
  );


  buf

  (
    n2682_o2_n_spl_,
    n2682_o2_n
  );


  buf

  (
    n5849_o2_p_spl_,
    n5849_o2_p
  );


  buf

  (
    n5849_o2_p_spl_0,
    n5849_o2_p_spl_
  );


  buf

  (
    n5598_o2_n_spl_,
    n5598_o2_n
  );


  buf

  (
    n5598_o2_n_spl_0,
    n5598_o2_n_spl_
  );


  buf

  (
    n5598_o2_n_spl_1,
    n5598_o2_n_spl_
  );


  buf

  (
    n4620_lo_n_spl_,
    n4620_lo_n
  );


  buf

  (
    n4620_lo_n_spl_0,
    n4620_lo_n_spl_
  );


  buf

  (
    n4620_lo_n_spl_00,
    n4620_lo_n_spl_0
  );


  buf

  (
    n4620_lo_n_spl_000,
    n4620_lo_n_spl_00
  );


  buf

  (
    n4620_lo_n_spl_001,
    n4620_lo_n_spl_00
  );


  buf

  (
    n4620_lo_n_spl_01,
    n4620_lo_n_spl_0
  );


  buf

  (
    n4620_lo_n_spl_010,
    n4620_lo_n_spl_01
  );


  buf

  (
    n4620_lo_n_spl_1,
    n4620_lo_n_spl_
  );


  buf

  (
    n4620_lo_n_spl_10,
    n4620_lo_n_spl_1
  );


  buf

  (
    n4620_lo_n_spl_11,
    n4620_lo_n_spl_1
  );


  buf

  (
    n5598_o2_p_spl_,
    n5598_o2_p
  );


  buf

  (
    n5598_o2_p_spl_0,
    n5598_o2_p_spl_
  );


  buf

  (
    n5598_o2_p_spl_1,
    n5598_o2_p_spl_
  );


  buf

  (
    n4608_lo_p_spl_,
    n4608_lo_p
  );


  buf

  (
    n4608_lo_p_spl_0,
    n4608_lo_p_spl_
  );


  buf

  (
    n4608_lo_p_spl_00,
    n4608_lo_p_spl_0
  );


  buf

  (
    n4608_lo_p_spl_000,
    n4608_lo_p_spl_00
  );


  buf

  (
    n4608_lo_p_spl_001,
    n4608_lo_p_spl_00
  );


  buf

  (
    n4608_lo_p_spl_01,
    n4608_lo_p_spl_0
  );


  buf

  (
    n4608_lo_p_spl_010,
    n4608_lo_p_spl_01
  );


  buf

  (
    n4608_lo_p_spl_1,
    n4608_lo_p_spl_
  );


  buf

  (
    n4608_lo_p_spl_10,
    n4608_lo_p_spl_1
  );


  buf

  (
    n4608_lo_p_spl_11,
    n4608_lo_p_spl_1
  );


  buf

  (
    n5325_o2_n_spl_,
    n5325_o2_n
  );


  buf

  (
    n5325_o2_n_spl_0,
    n5325_o2_n_spl_
  );


  buf

  (
    n5325_o2_p_spl_,
    n5325_o2_p
  );


  buf

  (
    n5325_o2_p_spl_0,
    n5325_o2_p_spl_
  );


  buf

  (
    n5833_o2_n_spl_,
    n5833_o2_n
  );


  buf

  (
    n5833_o2_n_spl_0,
    n5833_o2_n_spl_
  );


  buf

  (
    n5833_o2_p_spl_,
    n5833_o2_p
  );


  buf

  (
    n5833_o2_p_spl_0,
    n5833_o2_p_spl_
  );


  buf

  (
    n4293_lo_p_spl_,
    n4293_lo_p
  );


  buf

  (
    n4293_lo_p_spl_0,
    n4293_lo_p_spl_
  );


  buf

  (
    n4293_lo_p_spl_00,
    n4293_lo_p_spl_0
  );


  buf

  (
    n4293_lo_p_spl_1,
    n4293_lo_p_spl_
  );


  buf

  (
    g1711_n_spl_,
    g1711_n
  );


  buf

  (
    g1711_n_spl_0,
    g1711_n_spl_
  );


  buf

  (
    n4293_lo_n_spl_,
    n4293_lo_n
  );


  buf

  (
    n4293_lo_n_spl_0,
    n4293_lo_n_spl_
  );


  buf

  (
    n4293_lo_n_spl_1,
    n4293_lo_n_spl_
  );


  buf

  (
    g1711_p_spl_,
    g1711_p
  );


  buf

  (
    g1756_p_spl_,
    g1756_p
  );


  buf

  (
    lo494_buf_o2_p_spl_,
    lo494_buf_o2_p
  );


  buf

  (
    lo494_buf_o2_p_spl_0,
    lo494_buf_o2_p_spl_
  );


  buf

  (
    lo494_buf_o2_p_spl_00,
    lo494_buf_o2_p_spl_0
  );


  buf

  (
    lo494_buf_o2_p_spl_000,
    lo494_buf_o2_p_spl_00
  );


  buf

  (
    lo494_buf_o2_p_spl_001,
    lo494_buf_o2_p_spl_00
  );


  buf

  (
    lo494_buf_o2_p_spl_01,
    lo494_buf_o2_p_spl_0
  );


  buf

  (
    lo494_buf_o2_p_spl_1,
    lo494_buf_o2_p_spl_
  );


  buf

  (
    lo494_buf_o2_p_spl_10,
    lo494_buf_o2_p_spl_1
  );


  buf

  (
    lo494_buf_o2_p_spl_11,
    lo494_buf_o2_p_spl_1
  );


  buf

  (
    lo434_buf_o2_p_spl_,
    lo434_buf_o2_p
  );


  buf

  (
    lo494_buf_o2_n_spl_,
    lo494_buf_o2_n
  );


  buf

  (
    lo494_buf_o2_n_spl_0,
    lo494_buf_o2_n_spl_
  );


  buf

  (
    lo494_buf_o2_n_spl_00,
    lo494_buf_o2_n_spl_0
  );


  buf

  (
    lo494_buf_o2_n_spl_000,
    lo494_buf_o2_n_spl_00
  );


  buf

  (
    lo494_buf_o2_n_spl_01,
    lo494_buf_o2_n_spl_0
  );


  buf

  (
    lo494_buf_o2_n_spl_1,
    lo494_buf_o2_n_spl_
  );


  buf

  (
    lo494_buf_o2_n_spl_10,
    lo494_buf_o2_n_spl_1
  );


  buf

  (
    lo494_buf_o2_n_spl_11,
    lo494_buf_o2_n_spl_1
  );


  buf

  (
    lo557_buf_o2_p_spl_,
    lo557_buf_o2_p
  );


  buf

  (
    lo557_buf_o2_p_spl_0,
    lo557_buf_o2_p_spl_
  );


  buf

  (
    g1721_n_spl_,
    g1721_n
  );


  buf

  (
    g1721_n_spl_0,
    g1721_n_spl_
  );


  buf

  (
    lo573_buf_o2_p_spl_,
    lo573_buf_o2_p
  );


  buf

  (
    lo573_buf_o2_p_spl_0,
    lo573_buf_o2_p_spl_
  );


  buf

  (
    g1720_n_spl_,
    g1720_n
  );


  buf

  (
    g1720_n_spl_0,
    g1720_n_spl_
  );


  buf

  (
    lo466_buf_o2_p_spl_,
    lo466_buf_o2_p
  );


  buf

  (
    lo490_buf_o2_p_spl_,
    lo490_buf_o2_p
  );


  buf

  (
    lo490_buf_o2_p_spl_0,
    lo490_buf_o2_p_spl_
  );


  buf

  (
    lo490_buf_o2_p_spl_00,
    lo490_buf_o2_p_spl_0
  );


  buf

  (
    lo490_buf_o2_p_spl_000,
    lo490_buf_o2_p_spl_00
  );


  buf

  (
    lo490_buf_o2_p_spl_001,
    lo490_buf_o2_p_spl_00
  );


  buf

  (
    lo490_buf_o2_p_spl_01,
    lo490_buf_o2_p_spl_0
  );


  buf

  (
    lo490_buf_o2_p_spl_010,
    lo490_buf_o2_p_spl_01
  );


  buf

  (
    lo490_buf_o2_p_spl_011,
    lo490_buf_o2_p_spl_01
  );


  buf

  (
    lo490_buf_o2_p_spl_1,
    lo490_buf_o2_p_spl_
  );


  buf

  (
    lo490_buf_o2_p_spl_10,
    lo490_buf_o2_p_spl_1
  );


  buf

  (
    lo490_buf_o2_p_spl_11,
    lo490_buf_o2_p_spl_1
  );


  buf

  (
    lo490_buf_o2_n_spl_,
    lo490_buf_o2_n
  );


  buf

  (
    lo490_buf_o2_n_spl_0,
    lo490_buf_o2_n_spl_
  );


  buf

  (
    lo490_buf_o2_n_spl_00,
    lo490_buf_o2_n_spl_0
  );


  buf

  (
    lo490_buf_o2_n_spl_000,
    lo490_buf_o2_n_spl_00
  );


  buf

  (
    lo490_buf_o2_n_spl_001,
    lo490_buf_o2_n_spl_00
  );


  buf

  (
    lo490_buf_o2_n_spl_01,
    lo490_buf_o2_n_spl_0
  );


  buf

  (
    lo490_buf_o2_n_spl_010,
    lo490_buf_o2_n_spl_01
  );


  buf

  (
    lo490_buf_o2_n_spl_1,
    lo490_buf_o2_n_spl_
  );


  buf

  (
    lo490_buf_o2_n_spl_10,
    lo490_buf_o2_n_spl_1
  );


  buf

  (
    lo490_buf_o2_n_spl_11,
    lo490_buf_o2_n_spl_1
  );


  buf

  (
    g1704_p_spl_,
    g1704_p
  );


  buf

  (
    g1719_p_spl_,
    g1719_p
  );


  buf

  (
    g1719_p_spl_0,
    g1719_p_spl_
  );


  buf

  (
    g1772_n_spl_,
    g1772_n
  );


  buf

  (
    g1719_n_spl_,
    g1719_n
  );


  buf

  (
    g1772_p_spl_,
    g1772_p
  );


  buf

  (
    g1773_n_spl_,
    g1773_n
  );


  buf

  (
    g1773_p_spl_,
    g1773_p
  );


  buf

  (
    lo357_buf_o2_p_spl_,
    lo357_buf_o2_p
  );


  buf

  (
    lo417_buf_o2_p_spl_,
    lo417_buf_o2_p
  );


  buf

  (
    g1699_p_spl_,
    g1699_p
  );


  buf

  (
    g1699_p_spl_0,
    g1699_p_spl_
  );


  buf

  (
    g1781_p_spl_,
    g1781_p
  );


  buf

  (
    g1699_n_spl_,
    g1699_n
  );


  buf

  (
    g1699_n_spl_0,
    g1699_n_spl_
  );


  buf

  (
    g1699_n_spl_1,
    g1699_n_spl_
  );


  buf

  (
    g1781_n_spl_,
    g1781_n
  );


  buf

  (
    g1712_p_spl_,
    g1712_p
  );


  buf

  (
    g1712_p_spl_0,
    g1712_p_spl_
  );


  buf

  (
    g1785_p_spl_,
    g1785_p
  );


  buf

  (
    lo473_buf_o2_p_spl_,
    lo473_buf_o2_p
  );


  buf

  (
    lo536_buf_o2_p_spl_,
    lo536_buf_o2_p
  );


  buf

  (
    lo536_buf_o2_p_spl_0,
    lo536_buf_o2_p_spl_
  );


  buf

  (
    g1761_n_spl_,
    g1761_n
  );


  buf

  (
    g1761_n_spl_0,
    g1761_n_spl_
  );


  buf

  (
    lo553_buf_o2_p_spl_,
    lo553_buf_o2_p
  );


  buf

  (
    lo553_buf_o2_p_spl_0,
    lo553_buf_o2_p_spl_
  );


  buf

  (
    g1722_n_spl_,
    g1722_n
  );


  buf

  (
    g1722_n_spl_0,
    g1722_n_spl_
  );


  buf

  (
    g1763_n_spl_,
    g1763_n
  );


  buf

  (
    g1763_n_spl_0,
    g1763_n_spl_
  );


  buf

  (
    g1763_n_spl_1,
    g1763_n_spl_
  );


  buf

  (
    lo508_buf_o2_p_spl_,
    lo508_buf_o2_p
  );


  buf

  (
    lo512_buf_o2_p_spl_,
    lo512_buf_o2_p
  );


  buf

  (
    n4254_lo_p_spl_,
    n4254_lo_p
  );


  buf

  (
    n4254_lo_p_spl_0,
    n4254_lo_p_spl_
  );


  buf

  (
    g1780_n_spl_,
    g1780_n
  );


  buf

  (
    g1780_n_spl_0,
    g1780_n_spl_
  );


  buf

  (
    n4314_lo_p_spl_,
    n4314_lo_p
  );


  buf

  (
    n4314_lo_p_spl_0,
    n4314_lo_p_spl_
  );


  buf

  (
    g1777_n_spl_,
    g1777_n
  );


  buf

  (
    g1777_n_spl_0,
    g1777_n_spl_
  );


  buf

  (
    n4350_lo_p_spl_,
    n4350_lo_p
  );


  buf

  (
    n4350_lo_p_spl_0,
    n4350_lo_p_spl_
  );


  buf

  (
    g1790_n_spl_,
    g1790_n
  );


  buf

  (
    g1790_n_spl_0,
    g1790_n_spl_
  );


  buf

  (
    lo576_buf_o2_p_spl_,
    lo576_buf_o2_p
  );


  buf

  (
    lo576_buf_o2_p_spl_0,
    lo576_buf_o2_p_spl_
  );


  buf

  (
    g1767_n_spl_,
    g1767_n
  );


  buf

  (
    g1767_n_spl_0,
    g1767_n_spl_
  );


  buf

  (
    g1807_n_spl_,
    g1807_n
  );


  buf

  (
    g1797_p_spl_,
    g1797_p
  );


  buf

  (
    g1799_p_spl_,
    g1799_p
  );


  buf

  (
    g1799_p_spl_0,
    g1799_p_spl_
  );


  buf

  (
    n4728_lo_n_spl_,
    n4728_lo_n
  );


  buf

  (
    n4728_lo_n_spl_0,
    n4728_lo_n_spl_
  );


  buf

  (
    n4728_lo_n_spl_00,
    n4728_lo_n_spl_0
  );


  buf

  (
    n4728_lo_n_spl_000,
    n4728_lo_n_spl_00
  );


  buf

  (
    n4728_lo_n_spl_001,
    n4728_lo_n_spl_00
  );


  buf

  (
    n4728_lo_n_spl_01,
    n4728_lo_n_spl_0
  );


  buf

  (
    n4728_lo_n_spl_010,
    n4728_lo_n_spl_01
  );


  buf

  (
    n4728_lo_n_spl_1,
    n4728_lo_n_spl_
  );


  buf

  (
    n4728_lo_n_spl_10,
    n4728_lo_n_spl_1
  );


  buf

  (
    n4728_lo_n_spl_11,
    n4728_lo_n_spl_1
  );


  buf

  (
    n4728_lo_p_spl_,
    n4728_lo_p
  );


  buf

  (
    n4728_lo_p_spl_0,
    n4728_lo_p_spl_
  );


  buf

  (
    n4728_lo_p_spl_00,
    n4728_lo_p_spl_0
  );


  buf

  (
    n4728_lo_p_spl_000,
    n4728_lo_p_spl_00
  );


  buf

  (
    n4728_lo_p_spl_001,
    n4728_lo_p_spl_00
  );


  buf

  (
    n4728_lo_p_spl_01,
    n4728_lo_p_spl_0
  );


  buf

  (
    n4728_lo_p_spl_010,
    n4728_lo_p_spl_01
  );


  buf

  (
    n4728_lo_p_spl_011,
    n4728_lo_p_spl_01
  );


  buf

  (
    n4728_lo_p_spl_1,
    n4728_lo_p_spl_
  );


  buf

  (
    n4728_lo_p_spl_10,
    n4728_lo_p_spl_1
  );


  buf

  (
    n4728_lo_p_spl_100,
    n4728_lo_p_spl_10
  );


  buf

  (
    n4728_lo_p_spl_101,
    n4728_lo_p_spl_10
  );


  buf

  (
    n4728_lo_p_spl_11,
    n4728_lo_p_spl_1
  );


  buf

  (
    n5327_o2_n_spl_,
    n5327_o2_n
  );


  buf

  (
    n5327_o2_n_spl_0,
    n5327_o2_n_spl_
  );


  buf

  (
    n5327_o2_p_spl_,
    n5327_o2_p
  );


  buf

  (
    n5327_o2_p_spl_0,
    n5327_o2_p_spl_
  );


  buf

  (
    n4716_lo_n_spl_,
    n4716_lo_n
  );


  buf

  (
    n4716_lo_n_spl_0,
    n4716_lo_n_spl_
  );


  buf

  (
    n3252_lo_p_spl_,
    n3252_lo_p
  );


  buf

  (
    n4716_lo_p_spl_,
    n4716_lo_p
  );


  buf

  (
    n4716_lo_p_spl_0,
    n4716_lo_p_spl_
  );


  buf

  (
    n5918_o2_n_spl_,
    n5918_o2_n
  );


  buf

  (
    n5918_o2_p_spl_,
    n5918_o2_p
  );


  buf

  (
    n5920_o2_p_spl_,
    n5920_o2_p
  );


  buf

  (
    n5920_o2_p_spl_0,
    n5920_o2_p_spl_
  );


  buf

  (
    n2149_inv_p_spl_,
    n2149_inv_p
  );


  buf

  (
    n3478_o2_p_spl_,
    n3478_o2_p
  );


  buf

  (
    n3484_o2_p_spl_,
    n3484_o2_p
  );


  buf

  (
    n3478_o2_n_spl_,
    n3478_o2_n
  );


  buf

  (
    n3484_o2_n_spl_,
    n3484_o2_n
  );


  buf

  (
    g1831_p_spl_,
    g1831_p
  );


  buf

  (
    g1834_n_spl_,
    g1834_n
  );


  buf

  (
    g1831_n_spl_,
    g1831_n
  );


  buf

  (
    g1834_p_spl_,
    g1834_p
  );


  buf

  (
    n5663_o2_p_spl_,
    n5663_o2_p
  );


  buf

  (
    g1692_p_spl_,
    g1692_p
  );


  buf

  (
    g1692_p_spl_0,
    g1692_p_spl_
  );


  buf

  (
    g1840_n_spl_,
    g1840_n
  );


  buf

  (
    g1692_n_spl_,
    g1692_n
  );


  buf

  (
    g1692_n_spl_0,
    g1692_n_spl_
  );


  buf

  (
    g1840_p_spl_,
    g1840_p
  );


  buf

  (
    g1755_n_spl_,
    g1755_n
  );


  buf

  (
    g1737_n_spl_,
    g1737_n
  );


  buf

  (
    g1746_n_spl_,
    g1746_n
  );


  buf

  (
    g1854_p_spl_,
    g1854_p
  );


  buf

  (
    g1855_n_spl_,
    g1855_n
  );


  buf

  (
    g1854_n_spl_,
    g1854_n
  );


  buf

  (
    g1855_p_spl_,
    g1855_p
  );


  buf

  (
    n2502_o2_p_spl_,
    n2502_o2_p
  );


  buf

  (
    n2704_inv_p_spl_,
    n2704_inv_p
  );


  buf

  (
    g1859_p_spl_,
    g1859_p
  );


  buf

  (
    g1860_p_spl_,
    g1860_p
  );


  buf

  (
    g1859_n_spl_,
    g1859_n
  );


  buf

  (
    g1860_n_spl_,
    g1860_n
  );


  buf

  (
    n2620_inv_p_spl_,
    n2620_inv_p
  );


  buf

  (
    n2620_inv_p_spl_0,
    n2620_inv_p_spl_
  );


  buf

  (
    n2620_inv_p_spl_1,
    n2620_inv_p_spl_
  );


  buf

  (
    n2628_lo_n_spl_,
    n2628_lo_n
  );


  buf

  (
    n2620_inv_n_spl_,
    n2620_inv_n
  );


  buf

  (
    n2620_inv_n_spl_0,
    n2620_inv_n_spl_
  );


  buf

  (
    n2617_inv_n_spl_,
    n2617_inv_n
  );


  buf

  (
    n2617_inv_n_spl_0,
    n2617_inv_n_spl_
  );


  buf

  (
    n2617_inv_n_spl_1,
    n2617_inv_n_spl_
  );


  buf

  (
    n2617_inv_p_spl_,
    n2617_inv_p
  );


  buf

  (
    n2617_inv_p_spl_0,
    n2617_inv_p_spl_
  );


  buf

  (
    n2617_inv_p_spl_00,
    n2617_inv_p_spl_0
  );


  buf

  (
    n2617_inv_p_spl_1,
    n2617_inv_p_spl_
  );


  buf

  (
    g1872_n_spl_,
    g1872_n
  );


  buf

  (
    g1872_n_spl_0,
    g1872_n_spl_
  );


  buf

  (
    g1872_n_spl_00,
    g1872_n_spl_0
  );


  buf

  (
    g1872_n_spl_1,
    g1872_n_spl_
  );


  buf

  (
    g1872_p_spl_,
    g1872_p
  );


  buf

  (
    g1872_p_spl_0,
    g1872_p_spl_
  );


  buf

  (
    g1872_p_spl_00,
    g1872_p_spl_0
  );


  buf

  (
    g1872_p_spl_1,
    g1872_p_spl_
  );


  buf

  (
    n3048_o2_p_spl_,
    n3048_o2_p
  );


  buf

  (
    n3048_o2_n_spl_,
    n3048_o2_n
  );


  buf

  (
    n3048_o2_n_spl_0,
    n3048_o2_n_spl_
  );


  buf

  (
    g1877_n_spl_,
    g1877_n
  );


  buf

  (
    g1724_p_spl_,
    g1724_p
  );


  buf

  (
    n4188_lo_p_spl_,
    n4188_lo_p
  );


  buf

  (
    n4188_lo_p_spl_0,
    n4188_lo_p_spl_
  );


  buf

  (
    g1884_n_spl_,
    g1884_n
  );


  buf

  (
    n2863_o2_p_spl_,
    n2863_o2_p
  );


  buf

  (
    g1693_n_spl_,
    g1693_n
  );


  buf

  (
    g1891_p_spl_,
    g1891_p
  );


  buf

  (
    g1728_n_spl_,
    g1728_n
  );


  buf

  (
    n5823_o2_p_spl_,
    n5823_o2_p
  );


  buf

  (
    g1895_n_spl_,
    g1895_n
  );


  buf

  (
    n4098_lo_p_spl_,
    n4098_lo_p
  );


  buf

  (
    n2591_o2_n_spl_,
    n2591_o2_n
  );


  buf

  (
    n2591_o2_n_spl_0,
    n2591_o2_n_spl_
  );


  buf

  (
    g1708_n_spl_,
    g1708_n
  );


  buf

  (
    n5400_o2_p_spl_,
    n5400_o2_p
  );


  buf

  (
    n5400_o2_p_spl_0,
    n5400_o2_p_spl_
  );


  buf

  (
    n5400_o2_n_spl_,
    n5400_o2_n
  );


  buf

  (
    n5400_o2_n_spl_0,
    n5400_o2_n_spl_
  );


  buf

  (
    n5323_o2_p_spl_,
    n5323_o2_p
  );


  buf

  (
    n5323_o2_p_spl_0,
    n5323_o2_p_spl_
  );


  buf

  (
    n5323_o2_n_spl_,
    n5323_o2_n
  );


  buf

  (
    n5323_o2_n_spl_0,
    n5323_o2_n_spl_
  );


  buf

  (
    n5402_o2_p_spl_,
    n5402_o2_p
  );


  buf

  (
    n5402_o2_p_spl_0,
    n5402_o2_p_spl_
  );


  buf

  (
    n5402_o2_n_spl_,
    n5402_o2_n
  );


  buf

  (
    n5402_o2_n_spl_0,
    n5402_o2_n_spl_
  );


  buf

  (
    n5369_o2_n_spl_,
    n5369_o2_n
  );


  buf

  (
    n5369_o2_n_spl_0,
    n5369_o2_n_spl_
  );


  buf

  (
    n5369_o2_n_spl_1,
    n5369_o2_n_spl_
  );


  buf

  (
    n5369_o2_p_spl_,
    n5369_o2_p
  );


  buf

  (
    n5369_o2_p_spl_0,
    n5369_o2_p_spl_
  );


  buf

  (
    n5369_o2_p_spl_1,
    n5369_o2_p_spl_
  );


  buf

  (
    n5896_o2_n_spl_,
    n5896_o2_n
  );


  buf

  (
    n5896_o2_n_spl_0,
    n5896_o2_n_spl_
  );


  buf

  (
    n5896_o2_n_spl_1,
    n5896_o2_n_spl_
  );


  buf

  (
    n5896_o2_p_spl_,
    n5896_o2_p
  );


  buf

  (
    n5896_o2_p_spl_0,
    n5896_o2_p_spl_
  );


  buf

  (
    n5896_o2_p_spl_1,
    n5896_o2_p_spl_
  );


  buf

  (
    n5600_o2_n_spl_,
    n5600_o2_n
  );


  buf

  (
    n5600_o2_n_spl_0,
    n5600_o2_n_spl_
  );


  buf

  (
    n5600_o2_p_spl_,
    n5600_o2_p
  );


  buf

  (
    n5600_o2_p_spl_0,
    n5600_o2_p_spl_
  );


  buf

  (
    n5557_o2_n_spl_,
    n5557_o2_n
  );


  buf

  (
    n5557_o2_n_spl_0,
    n5557_o2_n_spl_
  );


  buf

  (
    n5557_o2_p_spl_,
    n5557_o2_p
  );


  buf

  (
    n5557_o2_p_spl_0,
    n5557_o2_p_spl_
  );


  buf

  (
    n3671_o2_n_spl_,
    n3671_o2_n
  );


  buf

  (
    n3680_o2_p_spl_,
    n3680_o2_p
  );


  buf

  (
    n3671_o2_p_spl_,
    n3671_o2_p
  );


  buf

  (
    n3680_o2_n_spl_,
    n3680_o2_n
  );


  buf

  (
    n3692_o2_n_spl_,
    n3692_o2_n
  );


  buf

  (
    n3692_o2_p_spl_,
    n3692_o2_p
  );


  buf

  (
    n2591_o2_p_spl_,
    n2591_o2_p
  );


  buf

  (
    n2591_o2_p_spl_0,
    n2591_o2_p_spl_
  );


  buf

  (
    g1982_n_spl_,
    g1982_n
  );


  buf

  (
    g1985_p_spl_,
    g1985_p
  );


  buf

  (
    g1982_p_spl_,
    g1982_p
  );


  buf

  (
    g1985_n_spl_,
    g1985_n
  );


  buf

  (
    n3707_o2_n_spl_,
    n3707_o2_n
  );


  buf

  (
    n3716_o2_p_spl_,
    n3716_o2_p
  );


  buf

  (
    n3707_o2_p_spl_,
    n3707_o2_p
  );


  buf

  (
    n3716_o2_n_spl_,
    n3716_o2_n
  );


  buf

  (
    n3749_o2_n_spl_,
    n3749_o2_n
  );


  buf

  (
    n3740_o2_n_spl_,
    n3740_o2_n
  );


  buf

  (
    n3749_o2_p_spl_,
    n3749_o2_p
  );


  buf

  (
    n3740_o2_p_spl_,
    n3740_o2_p
  );


  buf

  (
    g1991_p_spl_,
    g1991_p
  );


  buf

  (
    g1994_n_spl_,
    g1994_n
  );


  buf

  (
    g1991_n_spl_,
    g1991_n
  );


  buf

  (
    g1994_p_spl_,
    g1994_p
  );


  buf

  (
    n3936_lo_p_spl_,
    n3936_lo_p
  );


  buf

  (
    n3936_lo_p_spl_0,
    n3936_lo_p_spl_
  );


  buf

  (
    n5329_o2_p_spl_,
    n5329_o2_p
  );


  buf

  (
    n3936_lo_n_spl_,
    n3936_lo_n
  );


  buf

  (
    n3936_lo_n_spl_0,
    n3936_lo_n_spl_
  );


  buf

  (
    n5329_o2_n_spl_,
    n5329_o2_n
  );


  buf

  (
    n2818_o2_p_spl_,
    n2818_o2_p
  );


  buf

  (
    n2655_o2_p_spl_,
    n2655_o2_p
  );


  buf

  (
    lo450_buf_o2_p_spl_,
    lo450_buf_o2_p
  );


  buf

  (
    g2035_n_spl_,
    g2035_n
  );


  buf

  (
    g2038_p_spl_,
    g2038_p
  );


  buf

  (
    n4188_lo_n_spl_,
    n4188_lo_n
  );


  buf

  (
    n5653_o2_p_spl_,
    n5653_o2_p
  );


  buf

  (
    n5653_o2_n_spl_,
    n5653_o2_n
  );


  buf

  (
    g2046_n_spl_,
    g2046_n
  );


  buf

  (
    g2049_p_spl_,
    g2049_p
  );


  buf

  (
    g2054_n_spl_,
    g2054_n
  );


  buf

  (
    g2057_n_spl_,
    g2057_n
  );


  buf

  (
    g2069_p_spl_,
    g2069_p
  );


  buf

  (
    g2070_n_spl_,
    g2070_n
  );


  buf

  (
    g2069_n_spl_,
    g2069_n
  );


  buf

  (
    g2070_p_spl_,
    g2070_p
  );


  buf

  (
    n4488_lo_n_spl_,
    n4488_lo_n
  );


  buf

  (
    n4488_lo_n_spl_0,
    n4488_lo_n_spl_
  );


  buf

  (
    n4488_lo_n_spl_1,
    n4488_lo_n_spl_
  );


  buf

  (
    n4488_lo_p_spl_,
    n4488_lo_p
  );


  buf

  (
    n4488_lo_p_spl_0,
    n4488_lo_p_spl_
  );


  buf

  (
    n4488_lo_p_spl_1,
    n4488_lo_p_spl_
  );


  buf

  (
    g2075_p_spl_,
    g2075_p
  );


  buf

  (
    g2076_p_spl_,
    g2076_p
  );


  buf

  (
    g2075_n_spl_,
    g2075_n
  );


  buf

  (
    g2076_n_spl_,
    g2076_n
  );


  buf

  (
    g2082_n_spl_,
    g2082_n
  );


  buf

  (
    g2082_p_spl_,
    g2082_p
  );


  buf

  (
    g2085_p_spl_,
    g2085_p
  );


  buf

  (
    g2085_n_spl_,
    g2085_n
  );


  buf

  (
    g1793_p_spl_,
    g1793_p
  );


  buf

  (
    g1796_p_spl_,
    g1796_p
  );


  buf

  (
    g1796_p_spl_0,
    g1796_p_spl_
  );


  buf

  (
    g1762_p_spl_,
    g1762_p
  );


  buf

  (
    n5936_o2_n_spl_,
    n5936_o2_n
  );


  buf

  (
    lo398_buf_o2_n_spl_,
    lo398_buf_o2_n
  );


  buf

  (
    lo398_buf_o2_n_spl_0,
    lo398_buf_o2_n_spl_
  );


  buf

  (
    lo398_buf_o2_n_spl_00,
    lo398_buf_o2_n_spl_0
  );


  buf

  (
    lo398_buf_o2_n_spl_000,
    lo398_buf_o2_n_spl_00
  );


  buf

  (
    lo398_buf_o2_n_spl_001,
    lo398_buf_o2_n_spl_00
  );


  buf

  (
    lo398_buf_o2_n_spl_01,
    lo398_buf_o2_n_spl_0
  );


  buf

  (
    lo398_buf_o2_n_spl_010,
    lo398_buf_o2_n_spl_01
  );


  buf

  (
    lo398_buf_o2_n_spl_011,
    lo398_buf_o2_n_spl_01
  );


  buf

  (
    lo398_buf_o2_n_spl_1,
    lo398_buf_o2_n_spl_
  );


  buf

  (
    lo398_buf_o2_n_spl_10,
    lo398_buf_o2_n_spl_1
  );


  buf

  (
    lo398_buf_o2_n_spl_100,
    lo398_buf_o2_n_spl_10
  );


  buf

  (
    lo398_buf_o2_n_spl_101,
    lo398_buf_o2_n_spl_10
  );


  buf

  (
    lo398_buf_o2_n_spl_11,
    lo398_buf_o2_n_spl_1
  );


  buf

  (
    lo398_buf_o2_n_spl_110,
    lo398_buf_o2_n_spl_11
  );


  buf

  (
    lo398_buf_o2_n_spl_111,
    lo398_buf_o2_n_spl_11
  );


  buf

  (
    n5936_o2_p_spl_,
    n5936_o2_p
  );


  buf

  (
    n5936_o2_p_spl_0,
    n5936_o2_p_spl_
  );


  buf

  (
    lo402_buf_o2_n_spl_,
    lo402_buf_o2_n
  );


  buf

  (
    lo402_buf_o2_n_spl_0,
    lo402_buf_o2_n_spl_
  );


  buf

  (
    lo402_buf_o2_n_spl_00,
    lo402_buf_o2_n_spl_0
  );


  buf

  (
    lo402_buf_o2_n_spl_000,
    lo402_buf_o2_n_spl_00
  );


  buf

  (
    lo402_buf_o2_n_spl_001,
    lo402_buf_o2_n_spl_00
  );


  buf

  (
    lo402_buf_o2_n_spl_01,
    lo402_buf_o2_n_spl_0
  );


  buf

  (
    lo402_buf_o2_n_spl_010,
    lo402_buf_o2_n_spl_01
  );


  buf

  (
    lo402_buf_o2_n_spl_011,
    lo402_buf_o2_n_spl_01
  );


  buf

  (
    lo402_buf_o2_n_spl_1,
    lo402_buf_o2_n_spl_
  );


  buf

  (
    lo402_buf_o2_n_spl_10,
    lo402_buf_o2_n_spl_1
  );


  buf

  (
    lo402_buf_o2_n_spl_100,
    lo402_buf_o2_n_spl_10
  );


  buf

  (
    lo402_buf_o2_n_spl_101,
    lo402_buf_o2_n_spl_10
  );


  buf

  (
    lo402_buf_o2_n_spl_11,
    lo402_buf_o2_n_spl_1
  );


  buf

  (
    lo402_buf_o2_n_spl_110,
    lo402_buf_o2_n_spl_11
  );


  buf

  (
    lo406_buf_o2_p_spl_,
    lo406_buf_o2_p
  );


  buf

  (
    lo406_buf_o2_p_spl_0,
    lo406_buf_o2_p_spl_
  );


  buf

  (
    lo406_buf_o2_p_spl_00,
    lo406_buf_o2_p_spl_0
  );


  buf

  (
    lo406_buf_o2_p_spl_000,
    lo406_buf_o2_p_spl_00
  );


  buf

  (
    lo406_buf_o2_p_spl_001,
    lo406_buf_o2_p_spl_00
  );


  buf

  (
    lo406_buf_o2_p_spl_01,
    lo406_buf_o2_p_spl_0
  );


  buf

  (
    lo406_buf_o2_p_spl_010,
    lo406_buf_o2_p_spl_01
  );


  buf

  (
    lo406_buf_o2_p_spl_011,
    lo406_buf_o2_p_spl_01
  );


  buf

  (
    lo406_buf_o2_p_spl_1,
    lo406_buf_o2_p_spl_
  );


  buf

  (
    lo406_buf_o2_p_spl_10,
    lo406_buf_o2_p_spl_1
  );


  buf

  (
    lo406_buf_o2_p_spl_100,
    lo406_buf_o2_p_spl_10
  );


  buf

  (
    lo406_buf_o2_p_spl_101,
    lo406_buf_o2_p_spl_10
  );


  buf

  (
    lo406_buf_o2_p_spl_11,
    lo406_buf_o2_p_spl_1
  );


  buf

  (
    lo390_buf_o2_p_spl_,
    lo390_buf_o2_p
  );


  buf

  (
    lo390_buf_o2_p_spl_0,
    lo390_buf_o2_p_spl_
  );


  buf

  (
    lo390_buf_o2_p_spl_00,
    lo390_buf_o2_p_spl_0
  );


  buf

  (
    lo390_buf_o2_p_spl_000,
    lo390_buf_o2_p_spl_00
  );


  buf

  (
    lo390_buf_o2_p_spl_001,
    lo390_buf_o2_p_spl_00
  );


  buf

  (
    lo390_buf_o2_p_spl_01,
    lo390_buf_o2_p_spl_0
  );


  buf

  (
    lo390_buf_o2_p_spl_010,
    lo390_buf_o2_p_spl_01
  );


  buf

  (
    lo390_buf_o2_p_spl_011,
    lo390_buf_o2_p_spl_01
  );


  buf

  (
    lo390_buf_o2_p_spl_1,
    lo390_buf_o2_p_spl_
  );


  buf

  (
    lo390_buf_o2_p_spl_10,
    lo390_buf_o2_p_spl_1
  );


  buf

  (
    lo390_buf_o2_p_spl_100,
    lo390_buf_o2_p_spl_10
  );


  buf

  (
    lo390_buf_o2_p_spl_101,
    lo390_buf_o2_p_spl_10
  );


  buf

  (
    lo390_buf_o2_p_spl_11,
    lo390_buf_o2_p_spl_1
  );


  buf

  (
    lo390_buf_o2_p_spl_110,
    lo390_buf_o2_p_spl_11
  );


  buf

  (
    lo474_buf_o2_n_spl_,
    lo474_buf_o2_n
  );


  buf

  (
    lo474_buf_o2_p_spl_,
    lo474_buf_o2_p
  );


  buf

  (
    lo474_buf_o2_p_spl_0,
    lo474_buf_o2_p_spl_
  );


  buf

  (
    lo518_buf_o2_p_spl_,
    lo518_buf_o2_p
  );


  buf

  (
    lo458_buf_o2_p_spl_,
    lo458_buf_o2_p
  );


  buf

  (
    n3957_lo_p_spl_,
    n3957_lo_p
  );


  buf

  (
    n3957_lo_p_spl_0,
    n3957_lo_p_spl_
  );


  buf

  (
    n3834_lo_p_spl_,
    n3834_lo_p
  );


  buf

  (
    n4110_lo_p_spl_,
    n4110_lo_p
  );


  buf

  (
    n4122_lo_p_spl_,
    n4122_lo_p
  );


  buf

  (
    n2811_o2_p_spl_,
    n2811_o2_p
  );


  buf

  (
    n2811_o2_p_spl_0,
    n2811_o2_p_spl_
  );


  buf

  (
    n2811_o2_p_spl_1,
    n2811_o2_p_spl_
  );


  buf

  (
    n2811_o2_n_spl_,
    n2811_o2_n
  );


  buf

  (
    n2811_o2_n_spl_0,
    n2811_o2_n_spl_
  );


  buf

  (
    n2811_o2_n_spl_1,
    n2811_o2_n_spl_
  );


  buf

  (
    n2740_inv_p_spl_,
    n2740_inv_p
  );


  buf

  (
    g1758_p_spl_,
    g1758_p
  );


  buf

  (
    g1758_p_spl_0,
    g1758_p_spl_
  );


  buf

  (
    g2139_n_spl_,
    g2139_n
  );


  buf

  (
    g2139_n_spl_0,
    g2139_n_spl_
  );


  buf

  (
    n2779_inv_n_spl_,
    n2779_inv_n
  );


  buf

  (
    n2779_inv_n_spl_0,
    n2779_inv_n_spl_
  );


  buf

  (
    n2779_inv_n_spl_1,
    n2779_inv_n_spl_
  );


  buf

  (
    g1725_n_spl_,
    g1725_n
  );


  buf

  (
    g1758_n_spl_,
    g1758_n
  );


  buf

  (
    g1758_n_spl_0,
    g1758_n_spl_
  );


  buf

  (
    g1758_n_spl_1,
    g1758_n_spl_
  );


  buf

  (
    g2142_n_spl_,
    g2142_n
  );


  buf

  (
    n2317_inv_n_spl_,
    n2317_inv_n
  );


  buf

  (
    n2317_inv_p_spl_,
    n2317_inv_p
  );


  buf

  (
    n2317_inv_p_spl_0,
    n2317_inv_p_spl_
  );


  buf

  (
    n2572_inv_n_spl_,
    n2572_inv_n
  );


  buf

  (
    n2572_inv_n_spl_0,
    n2572_inv_n_spl_
  );


  buf

  (
    g2146_p_spl_,
    g2146_p
  );


  buf

  (
    n2572_inv_p_spl_,
    n2572_inv_p
  );


  buf

  (
    n2572_inv_p_spl_0,
    n2572_inv_p_spl_
  );


  buf

  (
    n2572_inv_p_spl_1,
    n2572_inv_p_spl_
  );


  buf

  (
    g2146_n_spl_,
    g2146_n
  );


  buf

  (
    n2689_o2_p_spl_,
    n2689_o2_p
  );


  buf

  (
    n2638_inv_p_spl_,
    n2638_inv_p
  );


  buf

  (
    n2779_inv_p_spl_,
    n2779_inv_p
  );


  buf

  (
    n2779_inv_p_spl_0,
    n2779_inv_p_spl_
  );


  buf

  (
    n2779_inv_p_spl_1,
    n2779_inv_p_spl_
  );


  buf

  (
    g2139_p_spl_,
    g2139_p
  );


  buf

  (
    g2139_p_spl_0,
    g2139_p_spl_
  );


  buf

  (
    g2151_n_spl_,
    g2151_n
  );


  buf

  (
    g2151_n_spl_0,
    g2151_n_spl_
  );


  buf

  (
    g2151_p_spl_,
    g2151_p
  );


  buf

  (
    g2151_p_spl_0,
    g2151_p_spl_
  );


  buf

  (
    g2157_n_spl_,
    g2157_n
  );


  buf

  (
    g1702_n_spl_,
    g1702_n
  );


  buf

  (
    g1702_n_spl_0,
    g1702_n_spl_
  );


  buf

  (
    g2161_p_spl_,
    g2161_p
  );


  buf

  (
    g1702_p_spl_,
    g1702_p
  );


  buf

  (
    g2161_n_spl_,
    g2161_n
  );


  buf

  (
    n2323_inv_n_spl_,
    n2323_inv_n
  );


  buf

  (
    n2323_inv_p_spl_,
    n2323_inv_p
  );


  buf

  (
    n2323_inv_p_spl_0,
    n2323_inv_p_spl_
  );


  buf

  (
    n2323_inv_p_spl_1,
    n2323_inv_p_spl_
  );


  buf

  (
    g2164_n_spl_,
    g2164_n
  );


  buf

  (
    g2165_p_spl_,
    g2165_p
  );


  buf

  (
    g1705_p_spl_,
    g1705_p
  );


  buf

  (
    n2662_o2_p_spl_,
    n2662_o2_p
  );


  buf

  (
    n2662_o2_p_spl_0,
    n2662_o2_p_spl_
  );


  buf

  (
    g2169_n_spl_,
    g2169_n
  );


  buf

  (
    n2662_o2_n_spl_,
    n2662_o2_n
  );


  buf

  (
    g2169_p_spl_,
    g2169_p
  );


  buf

  (
    g2167_n_spl_,
    g2167_n
  );


  buf

  (
    g2172_n_spl_,
    g2172_n
  );


  buf

  (
    g2172_n_spl_0,
    g2172_n_spl_
  );


  buf

  (
    g2096_n_spl_,
    g2096_n
  );


  buf

  (
    g1805_p_spl_,
    g1805_p
  );


  buf

  (
    g1808_p_spl_,
    g1808_p
  );


  buf

  (
    n5938_o2_p_spl_,
    n5938_o2_p
  );


  buf

  (
    n3969_lo_p_spl_,
    n3969_lo_p
  );


  buf

  (
    n5912_o2_n_spl_,
    n5912_o2_n
  );


  buf

  (
    n5912_o2_p_spl_,
    n5912_o2_p
  );


  buf

  (
    n5912_o2_p_spl_0,
    n5912_o2_p_spl_
  );


  buf

  (
    lo554_buf_o2_p_spl_,
    lo554_buf_o2_p
  );


  buf

  (
    n5910_o2_n_spl_,
    n5910_o2_n
  );


  buf

  (
    n5910_o2_p_spl_,
    n5910_o2_p
  );


  buf

  (
    n5910_o2_p_spl_0,
    n5910_o2_p_spl_
  );


  buf

  (
    lo558_buf_o2_p_spl_,
    lo558_buf_o2_p
  );


  buf

  (
    n5908_o2_n_spl_,
    n5908_o2_n
  );


  buf

  (
    n5908_o2_p_spl_,
    n5908_o2_p
  );


  buf

  (
    n5908_o2_p_spl_0,
    n5908_o2_p_spl_
  );


  buf

  (
    lo574_buf_o2_p_spl_,
    lo574_buf_o2_p
  );


  buf

  (
    n5934_o2_n_spl_,
    n5934_o2_n
  );


  buf

  (
    n5934_o2_p_spl_,
    n5934_o2_p
  );


  buf

  (
    n5934_o2_p_spl_0,
    n5934_o2_p_spl_
  );


  buf

  (
    lo538_buf_o2_p_spl_,
    lo538_buf_o2_p
  );


  buf

  (
    lo418_buf_o2_n_spl_,
    lo418_buf_o2_n
  );


  buf

  (
    lo418_buf_o2_p_spl_,
    lo418_buf_o2_p
  );


  buf

  (
    lo418_buf_o2_p_spl_0,
    lo418_buf_o2_p_spl_
  );


  buf

  (
    lo550_buf_o2_p_spl_,
    lo550_buf_o2_p
  );


  buf

  (
    lo358_buf_o2_n_spl_,
    lo358_buf_o2_n
  );


  buf

  (
    lo358_buf_o2_p_spl_,
    lo358_buf_o2_p
  );


  buf

  (
    lo358_buf_o2_p_spl_0,
    lo358_buf_o2_p_spl_
  );


  buf

  (
    lo570_buf_o2_p_spl_,
    lo570_buf_o2_p
  );


  buf

  (
    lo350_buf_o2_n_spl_,
    lo350_buf_o2_n
  );


  buf

  (
    lo350_buf_o2_p_spl_,
    lo350_buf_o2_p
  );


  buf

  (
    lo350_buf_o2_p_spl_0,
    lo350_buf_o2_p_spl_
  );


  buf

  (
    g1714_n_spl_,
    g1714_n
  );


  buf

  (
    g1714_n_spl_0,
    g1714_n_spl_
  );


  buf

  (
    g1714_p_spl_,
    g1714_p
  );


  buf

  (
    n2694_o2_p_spl_,
    n2694_o2_p
  );


  buf

  (
    g2253_n_spl_,
    g2253_n
  );


  buf

  (
    n2694_o2_n_spl_,
    n2694_o2_n
  );


  buf

  (
    g2253_p_spl_,
    g2253_p
  );


  buf

  (
    g2250_p_spl_,
    g2250_p
  );


  buf

  (
    g2259_n_spl_,
    g2259_n
  );


  buf

  (
    n3654_lo_p_spl_,
    n3654_lo_p
  );


  buf

  (
    g1768_n_spl_,
    g1768_n
  );


  buf

  (
    g2269_p_spl_,
    g2269_p
  );


  buf

  (
    g2272_p_spl_,
    g2272_p
  );


  buf

  (
    g1764_p_spl_,
    g1764_p
  );


  buf

  (
    g1764_p_spl_0,
    g1764_p_spl_
  );


  buf

  (
    g1809_p_spl_,
    g1809_p
  );


  buf

  (
    g2099_p_spl_,
    g2099_p
  );


  buf

  (
    g2099_p_spl_0,
    g2099_p_spl_
  );


  buf

  (
    g2275_n_spl_,
    g2275_n
  );


  buf

  (
    g2108_n_spl_,
    g2108_n
  );


  buf

  (
    g2108_n_spl_0,
    g2108_n_spl_
  );


  buf

  (
    g2123_n_spl_,
    g2123_n
  );


  buf

  (
    g2123_n_spl_0,
    g2123_n_spl_
  );


  buf

  (
    g2117_n_spl_,
    g2117_n
  );


  buf

  (
    g2117_n_spl_0,
    g2117_n_spl_
  );


  buf

  (
    g2126_p_spl_,
    g2126_p
  );


  buf

  (
    g2126_p_spl_0,
    g2126_p_spl_
  );


  buf

  (
    lo590_buf_o2_p_spl_,
    lo590_buf_o2_p
  );


  buf

  (
    lo590_buf_o2_p_spl_0,
    lo590_buf_o2_p_spl_
  );


  buf

  (
    lo590_buf_o2_n_spl_,
    lo590_buf_o2_n
  );


  buf

  (
    lo398_buf_o2_p_spl_,
    lo398_buf_o2_p
  );


  buf

  (
    lo398_buf_o2_p_spl_0,
    lo398_buf_o2_p_spl_
  );


  buf

  (
    lo398_buf_o2_p_spl_00,
    lo398_buf_o2_p_spl_0
  );


  buf

  (
    lo398_buf_o2_p_spl_1,
    lo398_buf_o2_p_spl_
  );


  buf

  (
    lo390_buf_o2_n_spl_,
    lo390_buf_o2_n
  );


  buf

  (
    lo390_buf_o2_n_spl_0,
    lo390_buf_o2_n_spl_
  );


  buf

  (
    lo390_buf_o2_n_spl_00,
    lo390_buf_o2_n_spl_0
  );


  buf

  (
    lo390_buf_o2_n_spl_1,
    lo390_buf_o2_n_spl_
  );


  buf

  (
    lo482_buf_o2_n_spl_,
    lo482_buf_o2_n
  );


  buf

  (
    lo482_buf_o2_n_spl_0,
    lo482_buf_o2_n_spl_
  );


  buf

  (
    lo482_buf_o2_n_spl_1,
    lo482_buf_o2_n_spl_
  );


  buf

  (
    lo482_buf_o2_p_spl_,
    lo482_buf_o2_p
  );


  buf

  (
    lo482_buf_o2_p_spl_0,
    lo482_buf_o2_p_spl_
  );


  buf

  (
    lo482_buf_o2_p_spl_00,
    lo482_buf_o2_p_spl_0
  );


  buf

  (
    lo482_buf_o2_p_spl_1,
    lo482_buf_o2_p_spl_
  );


  buf

  (
    lo402_buf_o2_p_spl_,
    lo402_buf_o2_p
  );


  buf

  (
    lo402_buf_o2_p_spl_0,
    lo402_buf_o2_p_spl_
  );


  buf

  (
    lo402_buf_o2_p_spl_1,
    lo402_buf_o2_p_spl_
  );


  buf

  (
    lo406_buf_o2_n_spl_,
    lo406_buf_o2_n
  );


  buf

  (
    lo406_buf_o2_n_spl_0,
    lo406_buf_o2_n_spl_
  );


  buf

  (
    lo406_buf_o2_n_spl_1,
    lo406_buf_o2_n_spl_
  );


  buf

  (
    g2120_n_spl_,
    g2120_n
  );


  buf

  (
    g2120_n_spl_0,
    g2120_n_spl_
  );


  buf

  (
    g2295_n_spl_,
    g2295_n
  );


  buf

  (
    lo510_buf_o2_n_spl_,
    lo510_buf_o2_n
  );


  buf

  (
    lo510_buf_o2_p_spl_,
    lo510_buf_o2_p
  );


  buf

  (
    lo510_buf_o2_p_spl_0,
    lo510_buf_o2_p_spl_
  );


  buf

  (
    lo598_buf_o2_p_spl_,
    lo598_buf_o2_p
  );


  buf

  (
    lo502_buf_o2_p_spl_,
    lo502_buf_o2_p
  );


  buf

  (
    lo502_buf_o2_p_spl_0,
    lo502_buf_o2_p_spl_
  );


  buf

  (
    lo502_buf_o2_n_spl_,
    lo502_buf_o2_n
  );


  buf

  (
    lo594_buf_o2_p_spl_,
    lo594_buf_o2_p
  );


  buf

  (
    g2306_n_spl_,
    g2306_n
  );


  buf

  (
    g2315_p_spl_,
    g2315_p
  );


  buf

  (
    n2641_inv_p_spl_,
    n2641_inv_p
  );


  buf

  (
    g1774_n_spl_,
    g1774_n
  );


  buf

  (
    g1787_n_spl_,
    g1787_n
  );


  buf

  (
    g1697_n_spl_,
    g1697_n
  );


  buf

  (
    g1697_n_spl_0,
    g1697_n_spl_
  );


  buf

  (
    g1701_p_spl_,
    g1701_p
  );


  buf

  (
    g1697_p_spl_,
    g1697_p
  );


  buf

  (
    g1701_n_spl_,
    g1701_n
  );


  buf

  (
    g1701_n_spl_0,
    g1701_n_spl_
  );


  buf

  (
    lo410_buf_o2_n_spl_,
    lo410_buf_o2_n
  );


  buf

  (
    lo410_buf_o2_n_spl_0,
    lo410_buf_o2_n_spl_
  );


  buf

  (
    lo410_buf_o2_n_spl_1,
    lo410_buf_o2_n_spl_
  );


  buf

  (
    lo410_buf_o2_p_spl_,
    lo410_buf_o2_p
  );


  buf

  (
    lo410_buf_o2_p_spl_0,
    lo410_buf_o2_p_spl_
  );


  buf

  (
    lo410_buf_o2_p_spl_00,
    lo410_buf_o2_p_spl_0
  );


  buf

  (
    lo410_buf_o2_p_spl_1,
    lo410_buf_o2_p_spl_
  );


  buf

  (
    lo546_buf_o2_p_spl_,
    lo546_buf_o2_p
  );


  buf

  (
    lo546_buf_o2_p_spl_0,
    lo546_buf_o2_p_spl_
  );


  buf

  (
    lo546_buf_o2_n_spl_,
    lo546_buf_o2_n
  );


  buf

  (
    n4545_lo_n_spl_,
    n4545_lo_n
  );


  buf

  (
    n4545_lo_p_spl_,
    n4545_lo_p
  );


  buf

  (
    g1716_n_spl_,
    g1716_n
  );


  buf

  (
    g1792_p_spl_,
    g1792_p
  );


  buf

  (
    n4386_lo_p_spl_,
    n4386_lo_p
  );


  buf

  (
    g2132_n_spl_,
    g2132_n
  );


  buf

  (
    n4398_lo_p_spl_,
    n4398_lo_p
  );


  buf

  (
    g1802_n_spl_,
    g1802_n
  );


  buf

  (
    g2133_n_spl_,
    g2133_n
  );


  buf

  (
    n3978_lo_p_spl_,
    n3978_lo_p
  );


  buf

  (
    n4050_lo_p_spl_,
    n4050_lo_p
  );


  buf

  (
    g2276_n_spl_,
    g2276_n
  );


  buf

  (
    g2276_n_spl_0,
    g2276_n_spl_
  );


  buf

  (
    g2137_p_spl_,
    g2137_p
  );


  buf

  (
    g2137_p_spl_0,
    g2137_p_spl_
  );


  buf

  (
    g2137_p_spl_1,
    g2137_p_spl_
  );


  buf

  (
    g2160_n_spl_,
    g2160_n
  );


  buf

  (
    g2160_n_spl_0,
    g2160_n_spl_
  );


  buf

  (
    g2175_p_spl_,
    g2175_p
  );


  buf

  (
    g2098_n_spl_,
    g2098_n
  );


  buf

  (
    g2135_p_spl_,
    g2135_p
  );


  buf

  (
    g1803_p_spl_,
    g1803_p
  );


  buf

  (
    g1804_p_spl_,
    g1804_p
  );


  buf

  (
    g2177_n_spl_,
    g2177_n
  );


  buf

  (
    n4302_lo_p_spl_,
    n4302_lo_p
  );


  buf

  (
    n4302_lo_p_spl_0,
    n4302_lo_p_spl_
  );


  buf

  (
    g2264_n_spl_,
    g2264_n
  );


  buf

  (
    g2264_n_spl_0,
    g2264_n_spl_
  );


  buf

  (
    g2267_p_spl_,
    g2267_p
  );


  buf

  (
    g2365_p_spl_,
    g2365_p
  );


  buf

  (
    n4374_lo_p_spl_,
    n4374_lo_p
  );


  buf

  (
    g1898_n_spl_,
    g1898_n
  );


  buf

  (
    g2268_n_spl_,
    g2268_n
  );


  buf

  (
    n4242_lo_p_spl_,
    n4242_lo_p
  );


  buf

  (
    g2129_n_spl_,
    g2129_n
  );


  buf

  (
    g2361_n_spl_,
    g2361_n
  );


  buf

  (
    g2362_n_spl_,
    g2362_n
  );


  buf

  (
    g2363_n_spl_,
    g2363_n
  );


  buf

  (
    G92_p_spl_,
    G92_p
  );


  buf

  (
    G124_p_spl_,
    G124_p
  );


  buf

  (
    G124_p_spl_0,
    G124_p_spl_
  );


  buf

  (
    G124_p_spl_1,
    G124_p_spl_
  );


  buf

  (
    G124_n_spl_,
    G124_n
  );


  buf

  (
    G124_n_spl_0,
    G124_n_spl_
  );


  buf

  (
    G94_p_spl_,
    G94_p
  );


  buf

  (
    G107_p_spl_,
    G107_p
  );


  buf

  (
    n4419_lo_n_spl_,
    n4419_lo_n
  );


  buf

  (
    n4419_lo_n_spl_0,
    n4419_lo_n_spl_
  );


  buf

  (
    n4431_lo_p_spl_,
    n4431_lo_p
  );


  buf

  (
    n2619_lo_n_spl_,
    n2619_lo_n
  );


  buf

  (
    n2619_lo_n_spl_0,
    n2619_lo_n_spl_
  );


  buf

  (
    n2619_lo_n_spl_1,
    n2619_lo_n_spl_
  );


  buf

  (
    n3975_lo_n_spl_,
    n3975_lo_n
  );


  buf

  (
    g1064_n_spl_,
    g1064_n
  );


  buf

  (
    g1102_n_spl_,
    g1102_n
  );


  buf

  (
    g1106_p_spl_,
    g1106_p
  );


  buf

  (
    g1126_p_spl_,
    g1126_p
  );


  buf

  (
    g1127_n_spl_,
    g1127_n
  );


endmodule
