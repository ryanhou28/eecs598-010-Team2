
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G1884,
  G1885,
  G1886,
  G1887,
  G1888,
  G1889,
  G1890,
  G1891,
  G1892,
  G1893,
  G1894,
  G1895,
  G1896,
  G1897,
  G1898,
  G1899,
  G1900,
  G1901,
  G1902,
  G1903,
  G1904,
  G1905,
  G1906,
  G1907,
  G1908
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;
  output G1884;output G1885;output G1886;output G1887;output G1888;output G1889;output G1890;output G1891;output G1892;output G1893;output G1894;output G1895;output G1896;output G1897;output G1898;output G1899;output G1900;output G1901;output G1902;output G1903;output G1904;output G1905;output G1906;output G1907;output G1908;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire g34_p;
  wire g34_n;
  wire g35_p;
  wire g35_n;
  wire g36_p;
  wire g36_n;
  wire g37_p;
  wire g37_n;
  wire g38_p;
  wire g38_n;
  wire g39_p;
  wire g39_n;
  wire g40_p;
  wire g40_n;
  wire g41_p;
  wire g41_n;
  wire g42_p;
  wire g42_n;
  wire g43_p;
  wire g43_n;
  wire g44_p;
  wire g44_n;
  wire g45_p;
  wire g45_n;
  wire g46_p;
  wire g46_n;
  wire g47_p;
  wire g47_n;
  wire g48_p;
  wire g48_n;
  wire g49_p;
  wire g49_n;
  wire g50_p;
  wire g50_n;
  wire g51_p;
  wire g51_n;
  wire g52_p;
  wire g52_n;
  wire g53_p;
  wire g53_n;
  wire g54_p;
  wire g54_n;
  wire g55_p;
  wire g55_n;
  wire g56_p;
  wire g56_n;
  wire g57_p;
  wire g57_n;
  wire g58_p;
  wire g58_n;
  wire g59_p;
  wire g59_n;
  wire g60_p;
  wire g60_n;
  wire g61_p;
  wire g61_n;
  wire g62_p;
  wire g62_n;
  wire g63_p;
  wire g63_n;
  wire g64_p;
  wire g64_n;
  wire g65_p;
  wire g65_n;
  wire g66_p;
  wire g66_n;
  wire g67_p;
  wire g67_n;
  wire g68_p;
  wire g68_n;
  wire g69_p;
  wire g69_n;
  wire g70_p;
  wire g70_n;
  wire g71_p;
  wire g71_n;
  wire g72_p;
  wire g72_n;
  wire g73_p;
  wire g73_n;
  wire g74_p;
  wire g74_n;
  wire g75_p;
  wire g75_n;
  wire g76_p;
  wire g76_n;
  wire g77_p;
  wire g77_n;
  wire g78_p;
  wire g78_n;
  wire g79_p;
  wire g79_n;
  wire g80_p;
  wire g80_n;
  wire g81_p;
  wire g81_n;
  wire g82_p;
  wire g82_n;
  wire g83_p;
  wire g83_n;
  wire g84_p;
  wire g84_n;
  wire g85_p;
  wire g85_n;
  wire g86_p;
  wire g86_n;
  wire g87_p;
  wire g87_n;
  wire g88_p;
  wire g88_n;
  wire g89_p;
  wire g89_n;
  wire g90_p;
  wire g90_n;
  wire g91_p;
  wire g91_n;
  wire g92_p;
  wire g92_n;
  wire g93_p;
  wire g93_n;
  wire g94_p;
  wire g94_n;
  wire g95_p;
  wire g95_n;
  wire g96_p;
  wire g96_n;
  wire g97_p;
  wire g97_n;
  wire g98_p;
  wire g98_n;
  wire g99_p;
  wire g99_n;
  wire g100_p;
  wire g100_n;
  wire g101_p;
  wire g101_n;
  wire g102_p;
  wire g102_n;
  wire g103_p;
  wire g103_n;
  wire g104_p;
  wire g104_n;
  wire g105_p;
  wire g105_n;
  wire g106_p;
  wire g106_n;
  wire g107_p;
  wire g107_n;
  wire g108_p;
  wire g108_n;
  wire g109_p;
  wire g109_n;
  wire g110_p;
  wire g110_n;
  wire g111_p;
  wire g111_n;
  wire g112_p;
  wire g112_n;
  wire g113_p;
  wire g113_n;
  wire g114_p;
  wire g114_n;
  wire g115_p;
  wire g115_n;
  wire g116_p;
  wire g116_n;
  wire g117_p;
  wire g117_n;
  wire g118_p;
  wire g118_n;
  wire g119_p;
  wire g119_n;
  wire g120_p;
  wire g120_n;
  wire g121_p;
  wire g121_n;
  wire g122_p;
  wire g122_n;
  wire g123_p;
  wire g123_n;
  wire g124_p;
  wire g124_n;
  wire g125_p;
  wire g125_n;
  wire g126_p;
  wire g126_n;
  wire g127_p;
  wire g127_n;
  wire g128_p;
  wire g128_n;
  wire g129_p;
  wire g129_n;
  wire g130_p;
  wire g130_n;
  wire g131_p;
  wire g131_n;
  wire g132_p;
  wire g132_n;
  wire g133_p;
  wire g133_n;
  wire g134_p;
  wire g134_n;
  wire g135_p;
  wire g135_n;
  wire g136_p;
  wire g136_n;
  wire g137_p;
  wire g137_n;
  wire g138_p;
  wire g138_n;
  wire g139_p;
  wire g139_n;
  wire g140_p;
  wire g140_n;
  wire g141_p;
  wire g141_n;
  wire g142_p;
  wire g142_n;
  wire g143_p;
  wire g143_n;
  wire g144_p;
  wire g144_n;
  wire g145_p;
  wire g145_n;
  wire g146_p;
  wire g146_n;
  wire g147_p;
  wire g147_n;
  wire g148_p;
  wire g148_n;
  wire g149_p;
  wire g149_n;
  wire g150_p;
  wire g150_n;
  wire g151_p;
  wire g151_n;
  wire g152_p;
  wire g152_n;
  wire g153_p;
  wire g153_n;
  wire g154_p;
  wire g154_n;
  wire g155_p;
  wire g155_n;
  wire g156_p;
  wire g156_n;
  wire g157_p;
  wire g157_n;
  wire g158_p;
  wire g158_n;
  wire g159_p;
  wire g159_n;
  wire g160_p;
  wire g160_n;
  wire g161_p;
  wire g161_n;
  wire g162_p;
  wire g162_n;
  wire g163_p;
  wire g163_n;
  wire g164_p;
  wire g164_n;
  wire g165_p;
  wire g165_n;
  wire g166_p;
  wire g166_n;
  wire g167_p;
  wire g167_n;
  wire g168_p;
  wire g168_n;
  wire g169_p;
  wire g169_n;
  wire g170_p;
  wire g170_n;
  wire g171_p;
  wire g171_n;
  wire g172_p;
  wire g172_n;
  wire g173_p;
  wire g173_n;
  wire g174_p;
  wire g174_n;
  wire g175_p;
  wire g175_n;
  wire g176_p;
  wire g176_n;
  wire g177_p;
  wire g177_n;
  wire g178_p;
  wire g178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire G29_n_spl_;
  wire G33_n_spl_;
  wire G33_n_spl_0;
  wire G33_n_spl_00;
  wire G33_n_spl_000;
  wire G33_n_spl_001;
  wire G33_n_spl_01;
  wire G33_n_spl_010;
  wire G33_n_spl_011;
  wire G33_n_spl_1;
  wire G33_n_spl_10;
  wire G33_n_spl_11;
  wire G29_p_spl_;
  wire G33_p_spl_;
  wire G33_p_spl_0;
  wire G33_p_spl_00;
  wire G33_p_spl_000;
  wire G33_p_spl_001;
  wire G33_p_spl_01;
  wire G33_p_spl_010;
  wire G33_p_spl_1;
  wire G33_p_spl_10;
  wire G33_p_spl_11;
  wire G23_n_spl_;
  wire G23_n_spl_0;
  wire G23_n_spl_1;
  wire G24_p_spl_;
  wire G24_p_spl_0;
  wire G24_p_spl_1;
  wire G23_p_spl_;
  wire G23_p_spl_0;
  wire G23_p_spl_1;
  wire G24_n_spl_;
  wire G24_n_spl_0;
  wire G24_n_spl_1;
  wire G31_n_spl_;
  wire G31_n_spl_0;
  wire G31_n_spl_00;
  wire G31_n_spl_000;
  wire G31_n_spl_001;
  wire G31_n_spl_01;
  wire G31_n_spl_010;
  wire G31_n_spl_011;
  wire G31_n_spl_1;
  wire G31_n_spl_10;
  wire G31_n_spl_11;
  wire g35_n_spl_;
  wire G31_p_spl_;
  wire G31_p_spl_0;
  wire G31_p_spl_00;
  wire G31_p_spl_000;
  wire G31_p_spl_001;
  wire G31_p_spl_01;
  wire G31_p_spl_010;
  wire G31_p_spl_011;
  wire G31_p_spl_1;
  wire G31_p_spl_10;
  wire G31_p_spl_100;
  wire G31_p_spl_101;
  wire G31_p_spl_11;
  wire G31_p_spl_110;
  wire g35_p_spl_;
  wire g34_p_spl_;
  wire g36_p_spl_;
  wire g34_n_spl_;
  wire g36_n_spl_;
  wire G32_n_spl_;
  wire g38_p_spl_;
  wire g38_p_spl_0;
  wire g38_p_spl_00;
  wire g38_p_spl_01;
  wire g38_p_spl_1;
  wire g38_p_spl_10;
  wire g39_n_spl_;
  wire g39_p_spl_;
  wire G20_p_spl_;
  wire g41_n_spl_;
  wire G20_n_spl_;
  wire g41_p_spl_;
  wire G22_p_spl_;
  wire G22_n_spl_;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_00;
  wire G4_p_spl_01;
  wire G4_p_spl_1;
  wire G4_p_spl_10;
  wire G14_n_spl_;
  wire G14_n_spl_0;
  wire G14_n_spl_00;
  wire G14_n_spl_1;
  wire G4_n_spl_;
  wire G4_n_spl_0;
  wire G4_n_spl_00;
  wire G4_n_spl_01;
  wire G4_n_spl_1;
  wire G4_n_spl_10;
  wire G14_p_spl_;
  wire G14_p_spl_0;
  wire G14_p_spl_00;
  wire G14_p_spl_1;
  wire g43_p_spl_;
  wire g46_p_spl_;
  wire g43_n_spl_;
  wire g46_n_spl_;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire G12_p_spl_00;
  wire G12_p_spl_1;
  wire G13_n_spl_;
  wire G13_n_spl_0;
  wire G13_n_spl_00;
  wire G13_n_spl_1;
  wire G12_n_spl_;
  wire G12_n_spl_0;
  wire G12_n_spl_00;
  wire G12_n_spl_1;
  wire G13_p_spl_;
  wire G13_p_spl_0;
  wire G13_p_spl_00;
  wire G13_p_spl_1;
  wire G11_p_spl_;
  wire G11_p_spl_0;
  wire G11_p_spl_00;
  wire G11_p_spl_1;
  wire g52_p_spl_;
  wire G11_n_spl_;
  wire G11_n_spl_0;
  wire G11_n_spl_00;
  wire G11_n_spl_1;
  wire g52_n_spl_;
  wire G10_n_spl_;
  wire G10_n_spl_0;
  wire G10_n_spl_00;
  wire G10_n_spl_1;
  wire G15_n_spl_;
  wire G15_n_spl_0;
  wire G15_n_spl_00;
  wire G15_n_spl_1;
  wire G10_p_spl_;
  wire G10_p_spl_0;
  wire G10_p_spl_00;
  wire G10_p_spl_1;
  wire G15_p_spl_;
  wire G15_p_spl_0;
  wire G15_p_spl_00;
  wire G15_p_spl_1;
  wire G16_p_spl_;
  wire G16_p_spl_0;
  wire G16_p_spl_00;
  wire G16_p_spl_1;
  wire g58_n_spl_;
  wire g58_n_spl_0;
  wire g58_n_spl_1;
  wire G16_n_spl_;
  wire G16_n_spl_0;
  wire G16_n_spl_00;
  wire G16_n_spl_1;
  wire g58_p_spl_;
  wire g58_p_spl_0;
  wire g58_p_spl_1;
  wire g55_n_spl_;
  wire g61_p_spl_;
  wire g61_p_spl_0;
  wire g61_p_spl_1;
  wire g55_p_spl_;
  wire g61_n_spl_;
  wire g61_n_spl_0;
  wire g61_n_spl_1;
  wire G2_p_spl_;
  wire G2_p_spl_0;
  wire G2_p_spl_00;
  wire G2_p_spl_1;
  wire G3_n_spl_;
  wire G3_n_spl_0;
  wire G3_n_spl_00;
  wire G3_n_spl_1;
  wire G2_n_spl_;
  wire G2_n_spl_0;
  wire G2_n_spl_00;
  wire G2_n_spl_1;
  wire G3_p_spl_;
  wire G3_p_spl_0;
  wire G3_p_spl_00;
  wire G3_p_spl_1;
  wire G1_p_spl_;
  wire G1_p_spl_0;
  wire G1_p_spl_00;
  wire G1_p_spl_1;
  wire g67_p_spl_;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire G1_n_spl_00;
  wire G1_n_spl_1;
  wire g67_n_spl_;
  wire g64_n_spl_;
  wire g64_n_spl_0;
  wire g64_n_spl_00;
  wire g64_n_spl_01;
  wire g64_n_spl_1;
  wire g70_n_spl_;
  wire g70_n_spl_0;
  wire g70_n_spl_1;
  wire g64_p_spl_;
  wire g64_p_spl_0;
  wire g64_p_spl_00;
  wire g64_p_spl_01;
  wire g64_p_spl_1;
  wire g70_p_spl_;
  wire g70_p_spl_0;
  wire g70_p_spl_1;
  wire g49_n_spl_;
  wire g73_n_spl_;
  wire g49_p_spl_;
  wire g73_p_spl_;
  wire g76_n_spl_;
  wire g76_p_spl_;
  wire G25_n_spl_;
  wire G25_n_spl_0;
  wire g77_p_spl_;
  wire G25_p_spl_;
  wire G25_p_spl_0;
  wire g77_n_spl_;
  wire g42_p_spl_;
  wire g42_p_spl_0;
  wire g80_n_spl_;
  wire g80_n_spl_0;
  wire g42_n_spl_;
  wire g80_p_spl_;
  wire G18_p_spl_;
  wire G18_n_spl_;
  wire g83_n_spl_;
  wire g83_p_spl_;
  wire g86_n_spl_;
  wire g86_p_spl_;
  wire G9_p_spl_;
  wire G9_p_spl_0;
  wire G9_p_spl_00;
  wire G9_p_spl_1;
  wire G9_n_spl_;
  wire G9_n_spl_0;
  wire G9_n_spl_00;
  wire G9_n_spl_1;
  wire g92_n_spl_;
  wire g92_n_spl_0;
  wire g92_n_spl_1;
  wire g92_p_spl_;
  wire g92_p_spl_0;
  wire g92_p_spl_1;
  wire g89_p_spl_;
  wire g95_p_spl_;
  wire g95_p_spl_0;
  wire g95_p_spl_1;
  wire g89_n_spl_;
  wire g95_n_spl_;
  wire g95_n_spl_0;
  wire g95_n_spl_1;
  wire G5_n_spl_;
  wire G5_n_spl_0;
  wire G5_n_spl_00;
  wire G5_n_spl_1;
  wire G8_n_spl_;
  wire G8_n_spl_0;
  wire G8_n_spl_00;
  wire G8_n_spl_01;
  wire G8_n_spl_1;
  wire G8_n_spl_10;
  wire G5_p_spl_;
  wire G5_p_spl_0;
  wire G5_p_spl_00;
  wire G5_p_spl_1;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire G8_p_spl_00;
  wire G8_p_spl_01;
  wire G8_p_spl_1;
  wire G8_p_spl_10;
  wire g101_p_spl_;
  wire g101_n_spl_;
  wire g98_n_spl_;
  wire g104_p_spl_;
  wire g98_p_spl_;
  wire g104_n_spl_;
  wire g107_n_spl_;
  wire G27_n_spl_;
  wire G27_n_spl_0;
  wire g108_p_spl_;
  wire G27_p_spl_;
  wire g108_n_spl_;
  wire G6_n_spl_;
  wire G6_n_spl_0;
  wire G6_n_spl_00;
  wire G6_n_spl_1;
  wire G6_p_spl_;
  wire G6_p_spl_0;
  wire G6_p_spl_00;
  wire G6_p_spl_1;
  wire g112_p_spl_;
  wire g112_n_spl_;
  wire g115_n_spl_;
  wire g118_n_spl_;
  wire g115_p_spl_;
  wire g118_p_spl_;
  wire G19_p_spl_;
  wire G19_n_spl_;
  wire g121_n_spl_;
  wire g123_n_spl_;
  wire g121_p_spl_;
  wire g123_p_spl_;
  wire g126_n_spl_;
  wire G28_n_spl_;
  wire G28_n_spl_0;
  wire g127_p_spl_;
  wire G28_p_spl_;
  wire g127_n_spl_;
  wire G7_n_spl_;
  wire G7_n_spl_0;
  wire G7_n_spl_00;
  wire G7_n_spl_1;
  wire G7_p_spl_;
  wire G7_p_spl_0;
  wire G7_p_spl_00;
  wire G7_p_spl_1;
  wire g133_p_spl_;
  wire g133_n_spl_;
  wire g136_n_spl_;
  wire g136_p_spl_;
  wire g141_p_spl_;
  wire g141_n_spl_;
  wire g139_n_spl_;
  wire g144_n_spl_;
  wire g139_p_spl_;
  wire g144_p_spl_;
  wire g147_n_spl_;
  wire g148_p_spl_;
  wire g149_n_spl_;
  wire g149_n_spl_0;
  wire g148_n_spl_;
  wire g149_p_spl_;
  wire G17_p_spl_;
  wire G17_n_spl_;
  wire g156_p_spl_;
  wire g156_n_spl_;
  wire g162_p_spl_;
  wire g162_n_spl_;
  wire g165_n_spl_;
  wire g165_n_spl_0;
  wire g165_n_spl_1;
  wire g165_p_spl_;
  wire g165_p_spl_0;
  wire g165_p_spl_1;
  wire g159_p_spl_;
  wire g168_p_spl_;
  wire g159_n_spl_;
  wire g168_n_spl_;
  wire g171_n_spl_;
  wire g171_p_spl_;
  wire G26_p_spl_;
  wire G26_p_spl_0;
  wire g172_n_spl_;
  wire G26_n_spl_;
  wire G26_n_spl_0;
  wire g172_p_spl_;
  wire g179_n_spl_;
  wire g179_p_spl_;
  wire G21_p_spl_;
  wire G21_n_spl_;
  wire g181_p_spl_;
  wire g184_p_spl_;
  wire g181_n_spl_;
  wire g184_n_spl_;
  wire g190_p_spl_;
  wire g193_n_spl_;
  wire g190_n_spl_;
  wire g193_p_spl_;
  wire g187_p_spl_;
  wire g196_n_spl_;
  wire g196_n_spl_0;
  wire g187_n_spl_;
  wire g196_p_spl_;
  wire g196_p_spl_0;
  wire g199_p_spl_;
  wire g199_n_spl_;
  wire g200_p_spl_;
  wire g201_n_spl_;
  wire g201_n_spl_0;
  wire g200_n_spl_;
  wire g201_p_spl_;
  wire g201_p_spl_0;
  wire g180_p_spl_;
  wire g180_p_spl_0;
  wire g204_n_spl_;
  wire g204_n_spl_0;
  wire g180_n_spl_;
  wire g204_p_spl_;
  wire g178_p_spl_;
  wire g178_n_spl_;
  wire g178_n_spl_0;
  wire g81_n_spl_;
  wire g206_p_spl_;
  wire g81_p_spl_;
  wire g206_n_spl_;
  wire g40_n_spl_;
  wire g207_p_spl_;
  wire g40_p_spl_;
  wire g207_n_spl_;
  wire g208_n_spl_;
  wire g208_n_spl_0;
  wire g208_n_spl_00;
  wire g208_n_spl_01;
  wire g208_n_spl_1;
  wire g208_n_spl_10;
  wire g208_p_spl_;
  wire g208_p_spl_0;
  wire g208_p_spl_00;
  wire g208_p_spl_01;
  wire g208_p_spl_1;
  wire g208_p_spl_10;
  wire G30_n_spl_;
  wire G30_p_spl_;
  wire g221_p_spl_;
  wire g221_n_spl_;
  wire g223_n_spl_;
  wire g223_n_spl_0;
  wire g223_p_spl_;
  wire g223_p_spl_0;
  wire g224_n_spl_;
  wire g224_n_spl_0;
  wire g224_n_spl_00;
  wire g224_n_spl_01;
  wire g224_n_spl_1;
  wire g224_p_spl_;
  wire g224_p_spl_0;
  wire g224_p_spl_00;
  wire g224_p_spl_01;
  wire g224_p_spl_1;
  wire g235_p_spl_;
  wire g235_n_spl_;
  wire g236_n_spl_;
  wire g236_n_spl_0;
  wire g236_n_spl_1;
  wire g236_p_spl_;
  wire g236_p_spl_0;
  wire g236_p_spl_1;
  wire g256_n_spl_;
  wire g256_n_spl_0;
  wire g256_n_spl_1;
  wire g256_p_spl_;
  wire g256_p_spl_0;
  wire g256_p_spl_1;
  wire g269_p_spl_;
  wire g269_p_spl_0;
  wire g269_p_spl_00;
  wire g269_p_spl_01;
  wire g269_p_spl_1;
  wire g269_p_spl_10;
  wire g269_n_spl_;
  wire g269_n_spl_0;
  wire g303_n_spl_;
  wire g303_p_spl_;
  wire g315_n_spl_;
  wire g315_p_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  and

  (
    g34_p,
    G29_n_spl_,
    G33_n_spl_000
  );


  or

  (
    g34_n,
    G29_p_spl_,
    G33_p_spl_000
  );


  and

  (
    g35_p,
    G23_n_spl_0,
    G24_p_spl_0
  );


  or

  (
    g35_n,
    G23_p_spl_0,
    G24_n_spl_0
  );


  and

  (
    g36_p,
    G31_n_spl_000,
    g35_n_spl_
  );


  or

  (
    g36_n,
    G31_p_spl_000,
    g35_p_spl_
  );


  and

  (
    g37_p,
    g34_p_spl_,
    g36_p_spl_
  );


  or

  (
    g37_n,
    g34_n_spl_,
    g36_n_spl_
  );


  and

  (
    g38_p,
    G32_n_spl_,
    G33_n_spl_000
  );


  or

  (
    g38_n,
    G32_p,
    G33_p_spl_000
  );


  and

  (
    g39_p,
    g35_n_spl_,
    g38_p_spl_00
  );


  or

  (
    g39_n,
    g35_p_spl_,
    g38_n
  );


  and

  (
    g40_p,
    g37_n,
    g39_n_spl_
  );


  or

  (
    g40_n,
    g37_p,
    g39_p_spl_
  );


  and

  (
    g41_p,
    G23_n_spl_0,
    G31_n_spl_000
  );


  or

  (
    g41_n,
    G23_p_spl_0,
    G31_p_spl_000
  );


  and

  (
    g42_p,
    G20_p_spl_,
    g41_n_spl_
  );


  or

  (
    g42_n,
    G20_n_spl_,
    g41_p_spl_
  );


  and

  (
    g43_p,
    G22_p_spl_,
    G33_n_spl_001
  );


  or

  (
    g43_n,
    G22_n_spl_,
    G33_p_spl_001
  );


  and

  (
    g44_p,
    G4_p_spl_00,
    G14_n_spl_00
  );


  or

  (
    g44_n,
    G4_n_spl_00,
    G14_p_spl_00
  );


  and

  (
    g45_p,
    G4_n_spl_00,
    G14_p_spl_00
  );


  or

  (
    g45_n,
    G4_p_spl_00,
    G14_n_spl_00
  );


  and

  (
    g46_p,
    g44_n,
    g45_n
  );


  or

  (
    g46_n,
    g44_p,
    g45_p
  );


  and

  (
    g47_p,
    g43_p_spl_,
    g46_p_spl_
  );


  or

  (
    g47_n,
    g43_n_spl_,
    g46_n_spl_
  );


  and

  (
    g48_p,
    g43_n_spl_,
    g46_n_spl_
  );


  or

  (
    g48_n,
    g43_p_spl_,
    g46_p_spl_
  );


  and

  (
    g49_p,
    g47_n,
    g48_n
  );


  or

  (
    g49_n,
    g47_p,
    g48_p
  );


  and

  (
    g50_p,
    G12_p_spl_00,
    G13_n_spl_00
  );


  or

  (
    g50_n,
    G12_n_spl_00,
    G13_p_spl_00
  );


  and

  (
    g51_p,
    G12_n_spl_00,
    G13_p_spl_00
  );


  or

  (
    g51_n,
    G12_p_spl_00,
    G13_n_spl_00
  );


  and

  (
    g52_p,
    g50_n,
    g51_n
  );


  or

  (
    g52_n,
    g50_p,
    g51_p
  );


  and

  (
    g53_p,
    G11_p_spl_00,
    g52_p_spl_
  );


  or

  (
    g53_n,
    G11_n_spl_00,
    g52_n_spl_
  );


  and

  (
    g54_p,
    G11_n_spl_00,
    g52_n_spl_
  );


  or

  (
    g54_n,
    G11_p_spl_00,
    g52_p_spl_
  );


  and

  (
    g55_p,
    g53_n,
    g54_n
  );


  or

  (
    g55_n,
    g53_p,
    g54_p
  );


  and

  (
    g56_p,
    G10_n_spl_00,
    G15_n_spl_00
  );


  or

  (
    g56_n,
    G10_p_spl_00,
    G15_p_spl_00
  );


  and

  (
    g57_p,
    G10_p_spl_00,
    G15_p_spl_00
  );


  or

  (
    g57_n,
    G10_n_spl_00,
    G15_n_spl_00
  );


  and

  (
    g58_p,
    g56_n,
    g57_n
  );


  or

  (
    g58_n,
    g56_p,
    g57_p
  );


  and

  (
    g59_p,
    G16_p_spl_00,
    g58_n_spl_0
  );


  or

  (
    g59_n,
    G16_n_spl_00,
    g58_p_spl_0
  );


  and

  (
    g60_p,
    G16_n_spl_00,
    g58_p_spl_0
  );


  or

  (
    g60_n,
    G16_p_spl_00,
    g58_n_spl_0
  );


  and

  (
    g61_p,
    g59_n,
    g60_n
  );


  or

  (
    g61_n,
    g59_p,
    g60_p
  );


  and

  (
    g62_p,
    g55_n_spl_,
    g61_p_spl_0
  );


  or

  (
    g62_n,
    g55_p_spl_,
    g61_n_spl_0
  );


  and

  (
    g63_p,
    g55_p_spl_,
    g61_n_spl_0
  );


  or

  (
    g63_n,
    g55_n_spl_,
    g61_p_spl_0
  );


  and

  (
    g64_p,
    g62_n,
    g63_n
  );


  or

  (
    g64_n,
    g62_p,
    g63_p
  );


  and

  (
    g65_p,
    G2_p_spl_00,
    G3_n_spl_00
  );


  or

  (
    g65_n,
    G2_n_spl_00,
    G3_p_spl_00
  );


  and

  (
    g66_p,
    G2_n_spl_00,
    G3_p_spl_00
  );


  or

  (
    g66_n,
    G2_p_spl_00,
    G3_n_spl_00
  );


  and

  (
    g67_p,
    g65_n,
    g66_n
  );


  or

  (
    g67_n,
    g65_p,
    g66_p
  );


  and

  (
    g68_p,
    G1_p_spl_00,
    g67_p_spl_
  );


  or

  (
    g68_n,
    G1_n_spl_00,
    g67_n_spl_
  );


  and

  (
    g69_p,
    G1_n_spl_00,
    g67_n_spl_
  );


  or

  (
    g69_n,
    G1_p_spl_00,
    g67_p_spl_
  );


  and

  (
    g70_p,
    g68_n,
    g69_n
  );


  or

  (
    g70_n,
    g68_p,
    g69_p
  );


  and

  (
    g71_p,
    g64_n_spl_00,
    g70_n_spl_0
  );


  or

  (
    g71_n,
    g64_p_spl_00,
    g70_p_spl_0
  );


  and

  (
    g72_p,
    g64_p_spl_00,
    g70_p_spl_0
  );


  or

  (
    g72_n,
    g64_n_spl_00,
    g70_n_spl_0
  );


  and

  (
    g73_p,
    g71_n,
    g72_n
  );


  or

  (
    g73_n,
    g71_p,
    g72_p
  );


  and

  (
    g74_p,
    g49_n_spl_,
    g73_n_spl_
  );


  or

  (
    g74_n,
    g49_p_spl_,
    g73_p_spl_
  );


  and

  (
    g75_p,
    g49_p_spl_,
    g73_p_spl_
  );


  or

  (
    g75_n,
    g49_n_spl_,
    g73_n_spl_
  );


  and

  (
    g76_p,
    g74_n,
    g75_n
  );


  or

  (
    g76_n,
    g74_p,
    g75_p
  );


  and

  (
    g77_p,
    G31_n_spl_001,
    g76_n_spl_
  );


  or

  (
    g77_n,
    G31_p_spl_001,
    g76_p_spl_
  );


  and

  (
    g78_p,
    G25_n_spl_0,
    g77_p_spl_
  );


  or

  (
    g78_n,
    G25_p_spl_0,
    g77_n_spl_
  );


  and

  (
    g79_p,
    G25_p_spl_0,
    g77_n_spl_
  );


  or

  (
    g79_n,
    G25_n_spl_0,
    g77_p_spl_
  );


  and

  (
    g80_p,
    g78_n,
    g79_n
  );


  or

  (
    g80_n,
    g78_p,
    g79_p
  );


  and

  (
    g81_p,
    g42_p_spl_0,
    g80_n_spl_0
  );


  or

  (
    g81_n,
    g42_n_spl_,
    g80_p_spl_
  );


  and

  (
    g82_p,
    G18_p_spl_,
    G33_n_spl_001
  );


  or

  (
    g82_n,
    G18_n_spl_,
    G33_p_spl_001
  );


  and

  (
    g83_p,
    G24_n_spl_0,
    g82_p
  );


  or

  (
    g83_n,
    G24_p_spl_0,
    g82_n
  );


  and

  (
    g84_p,
    G15_p_spl_0,
    g83_n_spl_
  );


  or

  (
    g84_n,
    G15_n_spl_0,
    g83_p_spl_
  );


  and

  (
    g85_p,
    G15_n_spl_1,
    g83_p_spl_
  );


  or

  (
    g85_n,
    G15_p_spl_1,
    g83_n_spl_
  );


  and

  (
    g86_p,
    g84_n,
    g85_n
  );


  or

  (
    g86_n,
    g84_p,
    g85_p
  );


  and

  (
    g87_p,
    G11_n_spl_0,
    g86_n_spl_
  );


  or

  (
    g87_n,
    G11_p_spl_0,
    g86_p_spl_
  );


  and

  (
    g88_p,
    G11_p_spl_1,
    g86_p_spl_
  );


  or

  (
    g88_n,
    G11_n_spl_1,
    g86_n_spl_
  );


  and

  (
    g89_p,
    g87_n,
    g88_n
  );


  or

  (
    g89_n,
    g87_p,
    g88_p
  );


  and

  (
    g90_p,
    G9_p_spl_00,
    G14_n_spl_0
  );


  or

  (
    g90_n,
    G9_n_spl_00,
    G14_p_spl_0
  );


  and

  (
    g91_p,
    G9_n_spl_00,
    G14_p_spl_1
  );


  or

  (
    g91_n,
    G9_p_spl_00,
    G14_n_spl_1
  );


  and

  (
    g92_p,
    g90_n,
    g91_n
  );


  or

  (
    g92_n,
    g90_p,
    g91_p
  );


  and

  (
    g93_p,
    G16_p_spl_0,
    g92_n_spl_0
  );


  or

  (
    g93_n,
    G16_n_spl_0,
    g92_p_spl_0
  );


  and

  (
    g94_p,
    G16_n_spl_1,
    g92_p_spl_0
  );


  or

  (
    g94_n,
    G16_p_spl_1,
    g92_n_spl_0
  );


  and

  (
    g95_p,
    g93_n,
    g94_n
  );


  or

  (
    g95_n,
    g93_p,
    g94_p
  );


  and

  (
    g96_p,
    g89_p_spl_,
    g95_p_spl_0
  );


  or

  (
    g96_n,
    g89_n_spl_,
    g95_n_spl_0
  );


  and

  (
    g97_p,
    g89_n_spl_,
    g95_n_spl_0
  );


  or

  (
    g97_n,
    g89_p_spl_,
    g95_p_spl_0
  );


  and

  (
    g98_p,
    g96_n,
    g97_n
  );


  or

  (
    g98_n,
    g96_p,
    g97_p
  );


  and

  (
    g99_p,
    G5_n_spl_00,
    G8_n_spl_00
  );


  or

  (
    g99_n,
    G5_p_spl_00,
    G8_p_spl_00
  );


  and

  (
    g100_p,
    G5_p_spl_00,
    G8_p_spl_00
  );


  or

  (
    g100_n,
    G5_n_spl_00,
    G8_n_spl_00
  );


  and

  (
    g101_p,
    g99_n,
    g100_n
  );


  or

  (
    g101_n,
    g99_p,
    g100_p
  );


  and

  (
    g102_p,
    G2_n_spl_0,
    g101_p_spl_
  );


  or

  (
    g102_n,
    G2_p_spl_0,
    g101_n_spl_
  );


  and

  (
    g103_p,
    G2_p_spl_1,
    g101_n_spl_
  );


  or

  (
    g103_n,
    G2_n_spl_1,
    g101_p_spl_
  );


  and

  (
    g104_p,
    g102_n,
    g103_n
  );


  or

  (
    g104_n,
    g102_p,
    g103_p
  );


  and

  (
    g105_p,
    g98_n_spl_,
    g104_p_spl_
  );


  or

  (
    g105_n,
    g98_p_spl_,
    g104_n_spl_
  );


  and

  (
    g106_p,
    g98_p_spl_,
    g104_n_spl_
  );


  or

  (
    g106_n,
    g98_n_spl_,
    g104_p_spl_
  );


  and

  (
    g107_p,
    g105_n,
    g106_n
  );


  or

  (
    g107_n,
    g105_p,
    g106_p
  );


  and

  (
    g108_p,
    G31_n_spl_001,
    g107_n_spl_
  );


  or

  (
    g108_n,
    G31_p_spl_001,
    g107_p
  );


  and

  (
    g109_p,
    G27_n_spl_0,
    g108_p_spl_
  );


  or

  (
    g109_n,
    G27_p_spl_,
    g108_n_spl_
  );


  and

  (
    g110_p,
    G6_n_spl_00,
    G8_n_spl_01
  );


  or

  (
    g110_n,
    G6_p_spl_00,
    G8_p_spl_01
  );


  and

  (
    g111_p,
    G6_p_spl_00,
    G8_p_spl_01
  );


  or

  (
    g111_n,
    G6_n_spl_00,
    G8_n_spl_01
  );


  and

  (
    g112_p,
    g110_n,
    g111_n
  );


  or

  (
    g112_n,
    g110_p,
    g111_p
  );


  and

  (
    g113_p,
    G3_n_spl_0,
    g112_p_spl_
  );


  or

  (
    g113_n,
    G3_p_spl_0,
    g112_n_spl_
  );


  and

  (
    g114_p,
    G3_p_spl_1,
    g112_n_spl_
  );


  or

  (
    g114_n,
    G3_n_spl_1,
    g112_p_spl_
  );


  and

  (
    g115_p,
    g113_n,
    g114_n
  );


  or

  (
    g115_n,
    g113_p,
    g114_p
  );


  and

  (
    g116_p,
    G12_n_spl_0,
    g58_n_spl_1
  );


  or

  (
    g116_n,
    G12_p_spl_0,
    g58_p_spl_1
  );


  and

  (
    g117_p,
    G12_p_spl_1,
    g58_p_spl_1
  );


  or

  (
    g117_n,
    G12_n_spl_1,
    g58_n_spl_1
  );


  and

  (
    g118_p,
    g116_n,
    g117_n
  );


  or

  (
    g118_n,
    g116_p,
    g117_p
  );


  and

  (
    g119_p,
    g115_n_spl_,
    g118_n_spl_
  );


  or

  (
    g119_n,
    g115_p_spl_,
    g118_p_spl_
  );


  and

  (
    g120_p,
    g115_p_spl_,
    g118_p_spl_
  );


  or

  (
    g120_n,
    g115_n_spl_,
    g118_n_spl_
  );


  and

  (
    g121_p,
    g119_n,
    g120_n
  );


  or

  (
    g121_n,
    g119_p,
    g120_p
  );


  and

  (
    g122_p,
    G19_p_spl_,
    G33_n_spl_010
  );


  or

  (
    g122_n,
    G19_n_spl_,
    G33_p_spl_010
  );


  and

  (
    g123_p,
    G23_n_spl_1,
    g122_p
  );


  or

  (
    g123_n,
    G23_p_spl_1,
    g122_n
  );


  and

  (
    g124_p,
    g121_n_spl_,
    g123_n_spl_
  );


  or

  (
    g124_n,
    g121_p_spl_,
    g123_p_spl_
  );


  and

  (
    g125_p,
    g121_p_spl_,
    g123_p_spl_
  );


  or

  (
    g125_n,
    g121_n_spl_,
    g123_n_spl_
  );


  and

  (
    g126_p,
    g124_n,
    g125_n
  );


  or

  (
    g126_n,
    g124_p,
    g125_p
  );


  and

  (
    g127_p,
    G31_n_spl_010,
    g126_n_spl_
  );


  or

  (
    g127_n,
    G31_p_spl_010,
    g126_p
  );


  and

  (
    g128_p,
    G28_n_spl_0,
    g127_p_spl_
  );


  or

  (
    g128_n,
    G28_p_spl_,
    g127_n_spl_
  );


  and

  (
    g129_p,
    G28_p_spl_,
    g127_n_spl_
  );


  or

  (
    g129_n,
    G28_n_spl_0,
    g127_p_spl_
  );


  and

  (
    g130_p,
    g128_n,
    g129_n
  );


  or

  (
    g130_n,
    g128_p,
    g129_p
  );


  and

  (
    g131_p,
    G7_n_spl_00,
    G10_n_spl_0
  );


  or

  (
    g131_n,
    G7_p_spl_00,
    G10_p_spl_0
  );


  and

  (
    g132_p,
    G7_p_spl_00,
    G10_p_spl_1
  );


  or

  (
    g132_n,
    G7_n_spl_00,
    G10_n_spl_1
  );


  and

  (
    g133_p,
    g131_n,
    g132_n
  );


  or

  (
    g133_n,
    g131_p,
    g132_p
  );


  and

  (
    g134_p,
    G4_n_spl_01,
    g133_p_spl_
  );


  or

  (
    g134_n,
    G4_p_spl_01,
    g133_n_spl_
  );


  and

  (
    g135_p,
    G4_p_spl_01,
    g133_n_spl_
  );


  or

  (
    g135_n,
    G4_n_spl_01,
    g133_p_spl_
  );


  and

  (
    g136_p,
    g134_n,
    g135_n
  );


  or

  (
    g136_n,
    g134_p,
    g135_p
  );


  and

  (
    g137_p,
    g95_n_spl_1,
    g136_n_spl_
  );


  or

  (
    g137_n,
    g95_p_spl_1,
    g136_p_spl_
  );


  and

  (
    g138_p,
    g95_p_spl_1,
    g136_p_spl_
  );


  or

  (
    g138_n,
    g95_n_spl_1,
    g136_n_spl_
  );


  and

  (
    g139_p,
    g137_n,
    g138_n
  );


  or

  (
    g139_n,
    g137_p,
    g138_p
  );


  and

  (
    g140_p,
    G20_p_spl_,
    G33_n_spl_010
  );


  or

  (
    g140_n,
    G20_n_spl_,
    G33_p_spl_010
  );


  and

  (
    g141_p,
    G23_n_spl_1,
    g140_p
  );


  or

  (
    g141_n,
    G23_p_spl_1,
    g140_n
  );


  and

  (
    g142_p,
    G13_n_spl_0,
    g141_p_spl_
  );


  or

  (
    g142_n,
    G13_p_spl_0,
    g141_n_spl_
  );


  and

  (
    g143_p,
    G13_p_spl_1,
    g141_n_spl_
  );


  or

  (
    g143_n,
    G13_n_spl_1,
    g141_p_spl_
  );


  and

  (
    g144_p,
    g142_n,
    g143_n
  );


  or

  (
    g144_n,
    g142_p,
    g143_p
  );


  and

  (
    g145_p,
    g139_n_spl_,
    g144_n_spl_
  );


  or

  (
    g145_n,
    g139_p_spl_,
    g144_p_spl_
  );


  and

  (
    g146_p,
    g139_p_spl_,
    g144_p_spl_
  );


  or

  (
    g146_n,
    g139_n_spl_,
    g144_n_spl_
  );


  and

  (
    g147_p,
    g145_n,
    g146_n
  );


  or

  (
    g147_n,
    g145_p,
    g146_p
  );


  and

  (
    g148_p,
    G31_n_spl_010,
    g147_n_spl_
  );


  or

  (
    g148_n,
    G31_p_spl_010,
    g147_p
  );


  and

  (
    g149_p,
    G19_p_spl_,
    g41_n_spl_
  );


  or

  (
    g149_n,
    G19_n_spl_,
    g41_p_spl_
  );


  and

  (
    g150_p,
    g148_p_spl_,
    g149_n_spl_0
  );


  or

  (
    g150_n,
    g148_n_spl_,
    g149_p_spl_
  );


  and

  (
    g151_p,
    g148_n_spl_,
    g149_p_spl_
  );


  or

  (
    g151_n,
    g148_p_spl_,
    g149_n_spl_0
  );


  and

  (
    g152_p,
    g150_n,
    g151_n
  );


  or

  (
    g152_n,
    g150_p,
    g151_p
  );


  and

  (
    g153_p,
    g130_p,
    g152_p
  );


  or

  (
    g153_n,
    g130_n,
    g152_n
  );


  and

  (
    g154_p,
    g109_n,
    g153_p
  );


  or

  (
    g154_n,
    g109_p,
    g153_n
  );


  and

  (
    g155_p,
    G17_p_spl_,
    G33_n_spl_011
  );


  or

  (
    g155_n,
    G17_n_spl_,
    G33_p_spl_01
  );


  and

  (
    g156_p,
    G24_n_spl_1,
    g155_p
  );


  or

  (
    g156_n,
    G24_p_spl_1,
    g155_n
  );


  and

  (
    g157_p,
    G1_p_spl_0,
    g156_p_spl_
  );


  or

  (
    g157_n,
    G1_n_spl_0,
    g156_n_spl_
  );


  and

  (
    g158_p,
    G1_n_spl_1,
    g156_n_spl_
  );


  or

  (
    g158_n,
    G1_p_spl_1,
    g156_p_spl_
  );


  and

  (
    g159_p,
    g157_n,
    g158_n
  );


  or

  (
    g159_n,
    g157_p,
    g158_p
  );


  and

  (
    g160_p,
    G6_p_spl_0,
    G7_n_spl_0
  );


  or

  (
    g160_n,
    G6_n_spl_0,
    G7_p_spl_0
  );


  and

  (
    g161_p,
    G6_n_spl_1,
    G7_p_spl_1
  );


  or

  (
    g161_n,
    G6_p_spl_1,
    G7_n_spl_1
  );


  and

  (
    g162_p,
    g160_n,
    g161_n
  );


  or

  (
    g162_n,
    g160_p,
    g161_p
  );


  and

  (
    g163_p,
    G5_p_spl_0,
    g162_p_spl_
  );


  or

  (
    g163_n,
    G5_n_spl_0,
    g162_n_spl_
  );


  and

  (
    g164_p,
    G5_n_spl_1,
    g162_n_spl_
  );


  or

  (
    g164_n,
    G5_p_spl_1,
    g162_p_spl_
  );


  and

  (
    g165_p,
    g163_n,
    g164_n
  );


  or

  (
    g165_n,
    g163_p,
    g164_p
  );


  and

  (
    g166_p,
    g64_n_spl_01,
    g165_n_spl_0
  );


  or

  (
    g166_n,
    g64_p_spl_01,
    g165_p_spl_0
  );


  and

  (
    g167_p,
    g64_p_spl_01,
    g165_p_spl_0
  );


  or

  (
    g167_n,
    g64_n_spl_01,
    g165_n_spl_0
  );


  and

  (
    g168_p,
    g166_n,
    g167_n
  );


  or

  (
    g168_n,
    g166_p,
    g167_p
  );


  and

  (
    g169_p,
    g159_p_spl_,
    g168_p_spl_
  );


  or

  (
    g169_n,
    g159_n_spl_,
    g168_n_spl_
  );


  and

  (
    g170_p,
    g159_n_spl_,
    g168_n_spl_
  );


  or

  (
    g170_n,
    g159_p_spl_,
    g168_p_spl_
  );


  and

  (
    g171_p,
    g169_n,
    g170_n
  );


  or

  (
    g171_n,
    g169_p,
    g170_p
  );


  and

  (
    g172_p,
    G31_n_spl_011,
    g171_n_spl_
  );


  or

  (
    g172_n,
    G31_p_spl_011,
    g171_p_spl_
  );


  and

  (
    g173_p,
    G26_p_spl_0,
    g172_n_spl_
  );


  or

  (
    g173_n,
    G26_n_spl_0,
    g172_p_spl_
  );


  and

  (
    g174_p,
    G27_p_spl_,
    g108_n_spl_
  );


  or

  (
    g174_n,
    G27_n_spl_0,
    g108_p_spl_
  );


  and

  (
    g175_p,
    G26_n_spl_0,
    g172_p_spl_
  );


  or

  (
    g175_n,
    G26_p_spl_0,
    g172_n_spl_
  );


  and

  (
    g176_p,
    g174_n,
    g175_n
  );


  or

  (
    g176_n,
    g174_p,
    g175_p
  );


  and

  (
    g177_p,
    g173_n,
    g176_p
  );


  or

  (
    g177_n,
    g173_p,
    g176_n
  );


  and

  (
    g178_p,
    g154_p,
    g177_p
  );


  or

  (
    g178_n,
    g154_n,
    g177_n
  );


  and

  (
    g179_p,
    G24_n_spl_1,
    G31_n_spl_011
  );


  or

  (
    g179_n,
    G24_p_spl_1,
    G31_p_spl_011
  );


  and

  (
    g180_p,
    G18_p_spl_,
    g179_n_spl_
  );


  or

  (
    g180_n,
    G18_n_spl_,
    g179_p_spl_
  );


  and

  (
    g181_p,
    G21_p_spl_,
    G33_n_spl_011
  );


  or

  (
    g181_n,
    G21_n_spl_,
    G33_p_spl_10
  );


  and

  (
    g182_p,
    G9_p_spl_0,
    g61_n_spl_1
  );


  or

  (
    g182_n,
    G9_n_spl_0,
    g61_p_spl_1
  );


  and

  (
    g183_p,
    G9_n_spl_1,
    g61_p_spl_1
  );


  or

  (
    g183_n,
    G9_p_spl_1,
    g61_n_spl_1
  );


  and

  (
    g184_p,
    g182_n,
    g183_n
  );


  or

  (
    g184_n,
    g182_p,
    g183_p
  );


  and

  (
    g185_p,
    g181_p_spl_,
    g184_p_spl_
  );


  or

  (
    g185_n,
    g181_n_spl_,
    g184_n_spl_
  );


  and

  (
    g186_p,
    g181_n_spl_,
    g184_n_spl_
  );


  or

  (
    g186_n,
    g181_p_spl_,
    g184_p_spl_
  );


  and

  (
    g187_p,
    g185_n,
    g186_n
  );


  or

  (
    g187_n,
    g185_p,
    g186_p
  );


  and

  (
    g188_p,
    g70_n_spl_1,
    g165_p_spl_1
  );


  or

  (
    g188_n,
    g70_p_spl_1,
    g165_n_spl_1
  );


  and

  (
    g189_p,
    g70_p_spl_1,
    g165_n_spl_1
  );


  or

  (
    g189_n,
    g70_n_spl_1,
    g165_p_spl_1
  );


  and

  (
    g190_p,
    g188_n,
    g189_n
  );


  or

  (
    g190_n,
    g188_p,
    g189_p
  );


  and

  (
    g191_p,
    G4_n_spl_10,
    G8_n_spl_10
  );


  or

  (
    g191_n,
    G4_p_spl_10,
    G8_p_spl_10
  );


  and

  (
    g192_p,
    G4_p_spl_10,
    G8_p_spl_10
  );


  or

  (
    g192_n,
    G4_n_spl_10,
    G8_n_spl_10
  );


  and

  (
    g193_p,
    g191_n,
    g192_n
  );


  or

  (
    g193_n,
    g191_p,
    g192_p
  );


  and

  (
    g194_p,
    g190_p_spl_,
    g193_n_spl_
  );


  or

  (
    g194_n,
    g190_n_spl_,
    g193_p_spl_
  );


  and

  (
    g195_p,
    g190_n_spl_,
    g193_p_spl_
  );


  or

  (
    g195_n,
    g190_p_spl_,
    g193_n_spl_
  );


  and

  (
    g196_p,
    g194_n,
    g195_n
  );


  or

  (
    g196_n,
    g194_p,
    g195_p
  );


  and

  (
    g197_p,
    g187_p_spl_,
    g196_n_spl_0
  );


  or

  (
    g197_n,
    g187_n_spl_,
    g196_p_spl_0
  );


  and

  (
    g198_p,
    g187_n_spl_,
    g196_p_spl_0
  );


  or

  (
    g198_n,
    g187_p_spl_,
    g196_n_spl_0
  );


  and

  (
    g199_p,
    g197_n,
    g198_n
  );


  or

  (
    g199_n,
    g197_p,
    g198_p
  );


  and

  (
    g200_p,
    G31_n_spl_10,
    g199_p_spl_
  );


  or

  (
    g200_n,
    G31_p_spl_100,
    g199_n_spl_
  );


  and

  (
    g201_p,
    G17_p_spl_,
    g179_n_spl_
  );


  or

  (
    g201_n,
    G17_n_spl_,
    g179_p_spl_
  );


  and

  (
    g202_p,
    g200_p_spl_,
    g201_n_spl_0
  );


  or

  (
    g202_n,
    g200_n_spl_,
    g201_p_spl_0
  );


  and

  (
    g203_p,
    g200_n_spl_,
    g201_p_spl_0
  );


  or

  (
    g203_n,
    g200_p_spl_,
    g201_n_spl_0
  );


  and

  (
    g204_p,
    g202_n,
    g203_n
  );


  or

  (
    g204_n,
    g202_p,
    g203_p
  );


  and

  (
    g205_p,
    g180_p_spl_0,
    g204_n_spl_0
  );


  or

  (
    g205_n,
    g180_n_spl_,
    g204_p_spl_
  );


  and

  (
    g206_p,
    g178_p_spl_,
    g205_n
  );


  or

  (
    g206_n,
    g178_n_spl_0,
    g205_p
  );


  and

  (
    g207_p,
    g81_n_spl_,
    g206_p_spl_
  );


  or

  (
    g207_n,
    g81_p_spl_,
    g206_n_spl_
  );


  and

  (
    g208_p,
    g40_n_spl_,
    g207_p_spl_
  );


  or

  (
    g208_n,
    g40_p_spl_,
    g207_n_spl_
  );


  and

  (
    g209_p,
    G1_p_spl_1,
    g208_n_spl_00
  );


  and

  (
    g210_p,
    G1_n_spl_1,
    g208_p_spl_00
  );


  or

  (
    g211_n,
    g209_p,
    g210_p
  );


  and

  (
    g212_p,
    G2_p_spl_1,
    g208_n_spl_00
  );


  and

  (
    g213_p,
    G2_n_spl_1,
    g208_p_spl_00
  );


  or

  (
    g214_n,
    g212_p,
    g213_p
  );


  and

  (
    g215_p,
    G3_p_spl_1,
    g208_n_spl_01
  );


  and

  (
    g216_p,
    G3_n_spl_1,
    g208_p_spl_01
  );


  or

  (
    g217_n,
    g215_p,
    g216_p
  );


  and

  (
    g218_p,
    G4_p_spl_1,
    g208_n_spl_01
  );


  and

  (
    g219_p,
    G4_n_spl_1,
    g208_p_spl_01
  );


  or

  (
    g220_n,
    g218_p,
    g219_p
  );


  and

  (
    g221_p,
    G30_n_spl_,
    G33_n_spl_10
  );


  or

  (
    g221_n,
    G30_p_spl_,
    G33_p_spl_10
  );


  and

  (
    g222_p,
    g36_p_spl_,
    g221_p_spl_
  );


  or

  (
    g222_n,
    g36_n_spl_,
    g221_n_spl_
  );


  and

  (
    g223_p,
    g39_n_spl_,
    g222_n
  );


  or

  (
    g223_n,
    g39_p_spl_,
    g222_p
  );


  and

  (
    g224_p,
    g207_p_spl_,
    g223_n_spl_0
  );


  or

  (
    g224_n,
    g207_n_spl_,
    g223_p_spl_0
  );


  and

  (
    g225_p,
    G10_p_spl_1,
    g224_n_spl_00
  );


  and

  (
    g226_p,
    G10_n_spl_1,
    g224_p_spl_00
  );


  or

  (
    g227_n,
    g225_p,
    g226_p
  );


  and

  (
    g228_p,
    G15_p_spl_1,
    g224_n_spl_00
  );


  and

  (
    g229_p,
    G15_n_spl_1,
    g224_p_spl_00
  );


  or

  (
    g230_n,
    g228_p,
    g229_p
  );


  and

  (
    g231_p,
    G16_p_spl_1,
    g224_n_spl_01
  );


  and

  (
    g232_p,
    G16_n_spl_1,
    g224_p_spl_01
  );


  or

  (
    g233_n,
    g231_p,
    g232_p
  );


  and

  (
    g234_p,
    g42_p_spl_0,
    g80_p_spl_
  );


  or

  (
    g234_n,
    g42_n_spl_,
    g80_n_spl_0
  );


  and

  (
    g235_p,
    g206_p_spl_,
    g234_p
  );


  or

  (
    g235_n,
    g206_n_spl_,
    g234_n
  );


  and

  (
    g236_p,
    g40_n_spl_,
    g235_p_spl_
  );


  or

  (
    g236_n,
    g40_p_spl_,
    g235_n_spl_
  );


  and

  (
    g237_p,
    G5_p_spl_1,
    g236_n_spl_0
  );


  and

  (
    g238_p,
    G5_n_spl_1,
    g236_p_spl_0
  );


  or

  (
    g239_n,
    g237_p,
    g238_p
  );


  and

  (
    g240_p,
    G6_p_spl_1,
    g236_n_spl_0
  );


  and

  (
    g241_p,
    G6_n_spl_1,
    g236_p_spl_0
  );


  or

  (
    g242_n,
    g240_p,
    g241_p
  );


  and

  (
    g243_p,
    G7_p_spl_1,
    g236_n_spl_1
  );


  and

  (
    g244_p,
    G7_n_spl_1,
    g236_p_spl_1
  );


  or

  (
    g245_n,
    g243_p,
    g244_p
  );


  and

  (
    g246_p,
    G8_p_spl_1,
    g236_n_spl_1
  );


  and

  (
    g247_p,
    G8_n_spl_1,
    g236_p_spl_1
  );


  or

  (
    g248_n,
    g246_p,
    g247_p
  );


  and

  (
    g249_p,
    g223_n_spl_0,
    g235_p_spl_
  );


  or

  (
    g249_n,
    g223_p_spl_0,
    g235_n_spl_
  );


  or

  (
    g250_n,
    G9_n_spl_1,
    g249_n
  );


  or

  (
    g251_n,
    G9_p_spl_1,
    g249_p
  );


  and

  (
    g252_p,
    g250_n,
    g251_n
  );


  and

  (
    g253_p,
    g178_p_spl_,
    g180_p_spl_0
  );


  or

  (
    g253_n,
    g178_n_spl_0,
    g180_n_spl_
  );


  and

  (
    g254_p,
    g81_n_spl_,
    g223_n_spl_
  );


  or

  (
    g254_n,
    g81_p_spl_,
    g223_p_spl_
  );


  and

  (
    g255_p,
    g204_p_spl_,
    g254_p
  );


  or

  (
    g255_n,
    g204_n_spl_0,
    g254_n
  );


  and

  (
    g256_p,
    g253_p,
    g255_p
  );


  or

  (
    g256_n,
    g253_n,
    g255_n
  );


  and

  (
    g257_p,
    G11_p_spl_1,
    g256_n_spl_0
  );


  and

  (
    g258_p,
    G11_n_spl_1,
    g256_p_spl_0
  );


  or

  (
    g259_n,
    g257_p,
    g258_p
  );


  and

  (
    g260_p,
    G12_p_spl_1,
    g256_n_spl_0
  );


  and

  (
    g261_p,
    G12_n_spl_1,
    g256_p_spl_0
  );


  or

  (
    g262_n,
    g260_p,
    g261_p
  );


  and

  (
    g263_p,
    G13_p_spl_1,
    g256_n_spl_1
  );


  and

  (
    g264_p,
    G13_n_spl_1,
    g256_p_spl_1
  );


  or

  (
    g265_n,
    g263_p,
    g264_p
  );


  and

  (
    g266_p,
    G14_p_spl_1,
    g256_n_spl_1
  );


  and

  (
    g267_p,
    G14_n_spl_1,
    g256_p_spl_1
  );


  or

  (
    g268_n,
    g266_p,
    g267_p
  );


  and

  (
    g269_p,
    g208_n_spl_10,
    g224_n_spl_01
  );


  or

  (
    g269_n,
    g208_p_spl_10,
    g224_p_spl_01
  );


  or

  (
    g270_n,
    G32_n_spl_,
    g269_p_spl_00
  );


  or

  (
    g271_n,
    g80_n_spl_,
    g204_n_spl_
  );


  or

  (
    g272_n,
    g42_p_spl_,
    g180_p_spl_
  );


  or

  (
    g273_n,
    g178_n_spl_,
    g272_n
  );


  or

  (
    g274_n,
    g271_n,
    g273_n
  );


  and

  (
    g275_p,
    g270_n,
    g274_n
  );


  and

  (
    g276_p,
    G33_n_spl_10,
    g275_p
  );


  and

  (
    g277_p,
    G31_n_spl_10,
    g201_p_spl_
  );


  or

  (
    g277_n,
    G31_p_spl_100,
    g201_n_spl_
  );


  and

  (
    g278_p,
    g269_n_spl_0,
    g277_p
  );


  or

  (
    g278_n,
    g269_p_spl_00,
    g277_n
  );


  or

  (
    g279_n,
    g199_n_spl_,
    g278_p
  );


  or

  (
    g280_n,
    g199_p_spl_,
    g278_n
  );


  and

  (
    g281_p,
    g279_n,
    g280_n
  );


  or

  (
    g282_n,
    g38_p_spl_00,
    g281_p
  );


  and

  (
    g283_p,
    G25_p_spl_,
    G31_n_spl_11
  );


  or

  (
    g283_n,
    G25_n_spl_,
    G31_p_spl_101
  );


  and

  (
    g284_p,
    g269_n_spl_0,
    g283_p
  );


  or

  (
    g284_n,
    g269_p_spl_01,
    g283_n
  );


  or

  (
    g285_n,
    g76_p_spl_,
    g284_p
  );


  or

  (
    g286_n,
    g76_n_spl_,
    g284_n
  );


  and

  (
    g287_p,
    g285_n,
    g286_n
  );


  or

  (
    g288_n,
    g38_p_spl_01,
    g287_p
  );


  or

  (
    g289_n,
    G27_n_spl_,
    G31_p_spl_101
  );


  or

  (
    g290_n,
    g269_p_spl_01,
    g289_n
  );


  and

  (
    g291_p,
    g107_n_spl_,
    g290_n
  );


  or

  (
    g292_n,
    g38_p_spl_01,
    g291_p
  );


  or

  (
    g293_n,
    G28_n_spl_,
    G31_p_spl_110
  );


  or

  (
    g294_n,
    g269_p_spl_10,
    g293_n
  );


  and

  (
    g295_p,
    g126_n_spl_,
    g294_n
  );


  or

  (
    g296_n,
    g38_p_spl_10,
    g295_p
  );


  or

  (
    g297_n,
    G31_p_spl_110,
    g149_n_spl_
  );


  or

  (
    g298_n,
    g269_p_spl_10,
    g297_n
  );


  and

  (
    g299_p,
    g147_n_spl_,
    g298_n
  );


  or

  (
    g300_n,
    g38_p_spl_10,
    g299_p
  );


  and

  (
    g301_p,
    G21_p_spl_,
    G29_p_spl_
  );


  or

  (
    g301_n,
    G21_n_spl_,
    G29_n_spl_
  );


  and

  (
    g302_p,
    G33_n_spl_11,
    g301_n
  );


  or

  (
    g302_n,
    G33_p_spl_11,
    g301_p
  );


  and

  (
    g303_p,
    g34_n_spl_,
    g196_p_spl_
  );


  or

  (
    g303_n,
    g34_p_spl_,
    g196_n_spl_
  );


  and

  (
    g304_p,
    g208_n_spl_10,
    g303_n_spl_
  );


  or

  (
    g304_n,
    g208_p_spl_10,
    g303_p_spl_
  );


  and

  (
    g305_p,
    g208_p_spl_1,
    g303_p_spl_
  );


  or

  (
    g305_n,
    g208_n_spl_1,
    g303_n_spl_
  );


  and

  (
    g306_p,
    g304_n,
    g305_n
  );


  or

  (
    g306_n,
    g304_p,
    g305_p
  );


  or

  (
    g307_n,
    g302_p,
    g306_n
  );


  or

  (
    g308_n,
    g302_n,
    g306_p
  );


  and

  (
    g309_p,
    g307_n,
    g308_n
  );


  and

  (
    g310_p,
    G22_p_spl_,
    G30_p_spl_
  );


  or

  (
    g310_n,
    G22_n_spl_,
    G30_n_spl_
  );


  and

  (
    g311_p,
    G33_n_spl_11,
    g310_n
  );


  or

  (
    g311_n,
    G33_p_spl_11,
    g310_p
  );


  and

  (
    g312_p,
    g64_p_spl_1,
    g92_n_spl_1
  );


  or

  (
    g312_n,
    g64_n_spl_1,
    g92_p_spl_1
  );


  and

  (
    g313_p,
    g64_n_spl_1,
    g92_p_spl_1
  );


  or

  (
    g313_n,
    g64_p_spl_1,
    g92_n_spl_1
  );


  and

  (
    g314_p,
    g312_n,
    g313_n
  );


  or

  (
    g314_n,
    g312_p,
    g313_p
  );


  and

  (
    g315_p,
    g221_n_spl_,
    g314_n
  );


  or

  (
    g315_n,
    g221_p_spl_,
    g314_p
  );


  and

  (
    g316_p,
    g224_n_spl_1,
    g315_n_spl_
  );


  or

  (
    g316_n,
    g224_p_spl_1,
    g315_p_spl_
  );


  and

  (
    g317_p,
    g224_p_spl_1,
    g315_p_spl_
  );


  or

  (
    g317_n,
    g224_n_spl_1,
    g315_n_spl_
  );


  and

  (
    g318_p,
    g316_n,
    g317_n
  );


  or

  (
    g318_n,
    g316_p,
    g317_p
  );


  or

  (
    g319_n,
    g311_p,
    g318_n
  );


  or

  (
    g320_n,
    g311_n,
    g318_p
  );


  and

  (
    g321_p,
    g319_n,
    g320_n
  );


  and

  (
    g322_p,
    G26_p_spl_,
    G31_n_spl_11
  );


  or

  (
    g322_n,
    G26_n_spl_,
    G31_p_spl_11
  );


  and

  (
    g323_p,
    g269_n_spl_,
    g322_p
  );


  or

  (
    g323_n,
    g269_p_spl_1,
    g322_n
  );


  or

  (
    g324_n,
    g171_p_spl_,
    g323_p
  );


  or

  (
    g325_n,
    g171_n_spl_,
    g323_n
  );


  and

  (
    g326_p,
    g324_n,
    g325_n
  );


  or

  (
    g327_n,
    g38_p_spl_1,
    g326_p
  );


  not

  (
    G1884,
    g211_n
  );


  not

  (
    G1885,
    g214_n
  );


  not

  (
    G1886,
    g217_n
  );


  not

  (
    G1887,
    g220_n
  );


  not

  (
    G1888,
    g227_n
  );


  not

  (
    G1889,
    g230_n
  );


  not

  (
    G1890,
    g233_n
  );


  not

  (
    G1891,
    g239_n
  );


  not

  (
    G1892,
    g242_n
  );


  not

  (
    G1893,
    g245_n
  );


  not

  (
    G1894,
    g248_n
  );


  not

  (
    G1895,
    g252_p
  );


  not

  (
    G1896,
    g259_n
  );


  not

  (
    G1897,
    g262_n
  );


  not

  (
    G1898,
    g265_n
  );


  not

  (
    G1899,
    g268_n
  );


  not

  (
    G1900,
    g276_p
  );


  not

  (
    G1901,
    g282_n
  );


  not

  (
    G1902,
    g288_n
  );


  not

  (
    G1903,
    g292_n
  );


  not

  (
    G1904,
    g296_n
  );


  not

  (
    G1905,
    g300_n
  );


  not

  (
    G1906,
    g309_p
  );


  not

  (
    G1907,
    g321_p
  );


  not

  (
    G1908,
    g327_n
  );


  buf

  (
    G29_n_spl_,
    G29_n
  );


  buf

  (
    G33_n_spl_,
    G33_n
  );


  buf

  (
    G33_n_spl_0,
    G33_n_spl_
  );


  buf

  (
    G33_n_spl_00,
    G33_n_spl_0
  );


  buf

  (
    G33_n_spl_000,
    G33_n_spl_00
  );


  buf

  (
    G33_n_spl_001,
    G33_n_spl_00
  );


  buf

  (
    G33_n_spl_01,
    G33_n_spl_0
  );


  buf

  (
    G33_n_spl_010,
    G33_n_spl_01
  );


  buf

  (
    G33_n_spl_011,
    G33_n_spl_01
  );


  buf

  (
    G33_n_spl_1,
    G33_n_spl_
  );


  buf

  (
    G33_n_spl_10,
    G33_n_spl_1
  );


  buf

  (
    G33_n_spl_11,
    G33_n_spl_1
  );


  buf

  (
    G29_p_spl_,
    G29_p
  );


  buf

  (
    G33_p_spl_,
    G33_p
  );


  buf

  (
    G33_p_spl_0,
    G33_p_spl_
  );


  buf

  (
    G33_p_spl_00,
    G33_p_spl_0
  );


  buf

  (
    G33_p_spl_000,
    G33_p_spl_00
  );


  buf

  (
    G33_p_spl_001,
    G33_p_spl_00
  );


  buf

  (
    G33_p_spl_01,
    G33_p_spl_0
  );


  buf

  (
    G33_p_spl_010,
    G33_p_spl_01
  );


  buf

  (
    G33_p_spl_1,
    G33_p_spl_
  );


  buf

  (
    G33_p_spl_10,
    G33_p_spl_1
  );


  buf

  (
    G33_p_spl_11,
    G33_p_spl_1
  );


  buf

  (
    G23_n_spl_,
    G23_n
  );


  buf

  (
    G23_n_spl_0,
    G23_n_spl_
  );


  buf

  (
    G23_n_spl_1,
    G23_n_spl_
  );


  buf

  (
    G24_p_spl_,
    G24_p
  );


  buf

  (
    G24_p_spl_0,
    G24_p_spl_
  );


  buf

  (
    G24_p_spl_1,
    G24_p_spl_
  );


  buf

  (
    G23_p_spl_,
    G23_p
  );


  buf

  (
    G23_p_spl_0,
    G23_p_spl_
  );


  buf

  (
    G23_p_spl_1,
    G23_p_spl_
  );


  buf

  (
    G24_n_spl_,
    G24_n
  );


  buf

  (
    G24_n_spl_0,
    G24_n_spl_
  );


  buf

  (
    G24_n_spl_1,
    G24_n_spl_
  );


  buf

  (
    G31_n_spl_,
    G31_n
  );


  buf

  (
    G31_n_spl_0,
    G31_n_spl_
  );


  buf

  (
    G31_n_spl_00,
    G31_n_spl_0
  );


  buf

  (
    G31_n_spl_000,
    G31_n_spl_00
  );


  buf

  (
    G31_n_spl_001,
    G31_n_spl_00
  );


  buf

  (
    G31_n_spl_01,
    G31_n_spl_0
  );


  buf

  (
    G31_n_spl_010,
    G31_n_spl_01
  );


  buf

  (
    G31_n_spl_011,
    G31_n_spl_01
  );


  buf

  (
    G31_n_spl_1,
    G31_n_spl_
  );


  buf

  (
    G31_n_spl_10,
    G31_n_spl_1
  );


  buf

  (
    G31_n_spl_11,
    G31_n_spl_1
  );


  buf

  (
    g35_n_spl_,
    g35_n
  );


  buf

  (
    G31_p_spl_,
    G31_p
  );


  buf

  (
    G31_p_spl_0,
    G31_p_spl_
  );


  buf

  (
    G31_p_spl_00,
    G31_p_spl_0
  );


  buf

  (
    G31_p_spl_000,
    G31_p_spl_00
  );


  buf

  (
    G31_p_spl_001,
    G31_p_spl_00
  );


  buf

  (
    G31_p_spl_01,
    G31_p_spl_0
  );


  buf

  (
    G31_p_spl_010,
    G31_p_spl_01
  );


  buf

  (
    G31_p_spl_011,
    G31_p_spl_01
  );


  buf

  (
    G31_p_spl_1,
    G31_p_spl_
  );


  buf

  (
    G31_p_spl_10,
    G31_p_spl_1
  );


  buf

  (
    G31_p_spl_100,
    G31_p_spl_10
  );


  buf

  (
    G31_p_spl_101,
    G31_p_spl_10
  );


  buf

  (
    G31_p_spl_11,
    G31_p_spl_1
  );


  buf

  (
    G31_p_spl_110,
    G31_p_spl_11
  );


  buf

  (
    g35_p_spl_,
    g35_p
  );


  buf

  (
    g34_p_spl_,
    g34_p
  );


  buf

  (
    g36_p_spl_,
    g36_p
  );


  buf

  (
    g34_n_spl_,
    g34_n
  );


  buf

  (
    g36_n_spl_,
    g36_n
  );


  buf

  (
    G32_n_spl_,
    G32_n
  );


  buf

  (
    g38_p_spl_,
    g38_p
  );


  buf

  (
    g38_p_spl_0,
    g38_p_spl_
  );


  buf

  (
    g38_p_spl_00,
    g38_p_spl_0
  );


  buf

  (
    g38_p_spl_01,
    g38_p_spl_0
  );


  buf

  (
    g38_p_spl_1,
    g38_p_spl_
  );


  buf

  (
    g38_p_spl_10,
    g38_p_spl_1
  );


  buf

  (
    g39_n_spl_,
    g39_n
  );


  buf

  (
    g39_p_spl_,
    g39_p
  );


  buf

  (
    G20_p_spl_,
    G20_p
  );


  buf

  (
    g41_n_spl_,
    g41_n
  );


  buf

  (
    G20_n_spl_,
    G20_n
  );


  buf

  (
    g41_p_spl_,
    g41_p
  );


  buf

  (
    G22_p_spl_,
    G22_p
  );


  buf

  (
    G22_n_spl_,
    G22_n
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_00,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_01,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_10,
    G4_p_spl_1
  );


  buf

  (
    G14_n_spl_,
    G14_n
  );


  buf

  (
    G14_n_spl_0,
    G14_n_spl_
  );


  buf

  (
    G14_n_spl_00,
    G14_n_spl_0
  );


  buf

  (
    G14_n_spl_1,
    G14_n_spl_
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    G4_n_spl_0,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_00,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_01,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_1,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_10,
    G4_n_spl_1
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G14_p_spl_0,
    G14_p_spl_
  );


  buf

  (
    G14_p_spl_00,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_1,
    G14_p_spl_
  );


  buf

  (
    g43_p_spl_,
    g43_p
  );


  buf

  (
    g46_p_spl_,
    g46_p
  );


  buf

  (
    g43_n_spl_,
    g43_n
  );


  buf

  (
    g46_n_spl_,
    g46_n
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_00,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_1,
    G12_p_spl_
  );


  buf

  (
    G13_n_spl_,
    G13_n
  );


  buf

  (
    G13_n_spl_0,
    G13_n_spl_
  );


  buf

  (
    G13_n_spl_00,
    G13_n_spl_0
  );


  buf

  (
    G13_n_spl_1,
    G13_n_spl_
  );


  buf

  (
    G12_n_spl_,
    G12_n
  );


  buf

  (
    G12_n_spl_0,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_00,
    G12_n_spl_0
  );


  buf

  (
    G12_n_spl_1,
    G12_n_spl_
  );


  buf

  (
    G13_p_spl_,
    G13_p
  );


  buf

  (
    G13_p_spl_0,
    G13_p_spl_
  );


  buf

  (
    G13_p_spl_00,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_1,
    G13_p_spl_
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    G11_p_spl_0,
    G11_p_spl_
  );


  buf

  (
    G11_p_spl_00,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_1,
    G11_p_spl_
  );


  buf

  (
    g52_p_spl_,
    g52_p
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    G11_n_spl_0,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_00,
    G11_n_spl_0
  );


  buf

  (
    G11_n_spl_1,
    G11_n_spl_
  );


  buf

  (
    g52_n_spl_,
    g52_n
  );


  buf

  (
    G10_n_spl_,
    G10_n
  );


  buf

  (
    G10_n_spl_0,
    G10_n_spl_
  );


  buf

  (
    G10_n_spl_00,
    G10_n_spl_0
  );


  buf

  (
    G10_n_spl_1,
    G10_n_spl_
  );


  buf

  (
    G15_n_spl_,
    G15_n
  );


  buf

  (
    G15_n_spl_0,
    G15_n_spl_
  );


  buf

  (
    G15_n_spl_00,
    G15_n_spl_0
  );


  buf

  (
    G15_n_spl_1,
    G15_n_spl_
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


  buf

  (
    G10_p_spl_0,
    G10_p_spl_
  );


  buf

  (
    G10_p_spl_00,
    G10_p_spl_0
  );


  buf

  (
    G10_p_spl_1,
    G10_p_spl_
  );


  buf

  (
    G15_p_spl_,
    G15_p
  );


  buf

  (
    G15_p_spl_0,
    G15_p_spl_
  );


  buf

  (
    G15_p_spl_00,
    G15_p_spl_0
  );


  buf

  (
    G15_p_spl_1,
    G15_p_spl_
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    G16_p_spl_0,
    G16_p_spl_
  );


  buf

  (
    G16_p_spl_00,
    G16_p_spl_0
  );


  buf

  (
    G16_p_spl_1,
    G16_p_spl_
  );


  buf

  (
    g58_n_spl_,
    g58_n
  );


  buf

  (
    g58_n_spl_0,
    g58_n_spl_
  );


  buf

  (
    g58_n_spl_1,
    g58_n_spl_
  );


  buf

  (
    G16_n_spl_,
    G16_n
  );


  buf

  (
    G16_n_spl_0,
    G16_n_spl_
  );


  buf

  (
    G16_n_spl_00,
    G16_n_spl_0
  );


  buf

  (
    G16_n_spl_1,
    G16_n_spl_
  );


  buf

  (
    g58_p_spl_,
    g58_p
  );


  buf

  (
    g58_p_spl_0,
    g58_p_spl_
  );


  buf

  (
    g58_p_spl_1,
    g58_p_spl_
  );


  buf

  (
    g55_n_spl_,
    g55_n
  );


  buf

  (
    g61_p_spl_,
    g61_p
  );


  buf

  (
    g61_p_spl_0,
    g61_p_spl_
  );


  buf

  (
    g61_p_spl_1,
    g61_p_spl_
  );


  buf

  (
    g55_p_spl_,
    g55_p
  );


  buf

  (
    g61_n_spl_,
    g61_n
  );


  buf

  (
    g61_n_spl_0,
    g61_n_spl_
  );


  buf

  (
    g61_n_spl_1,
    g61_n_spl_
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G2_p_spl_0,
    G2_p_spl_
  );


  buf

  (
    G2_p_spl_00,
    G2_p_spl_0
  );


  buf

  (
    G2_p_spl_1,
    G2_p_spl_
  );


  buf

  (
    G3_n_spl_,
    G3_n
  );


  buf

  (
    G3_n_spl_0,
    G3_n_spl_
  );


  buf

  (
    G3_n_spl_00,
    G3_n_spl_0
  );


  buf

  (
    G3_n_spl_1,
    G3_n_spl_
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G2_n_spl_0,
    G2_n_spl_
  );


  buf

  (
    G2_n_spl_00,
    G2_n_spl_0
  );


  buf

  (
    G2_n_spl_1,
    G2_n_spl_
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G3_p_spl_0,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_00,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_1,
    G3_p_spl_
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G1_p_spl_0,
    G1_p_spl_
  );


  buf

  (
    G1_p_spl_00,
    G1_p_spl_0
  );


  buf

  (
    G1_p_spl_1,
    G1_p_spl_
  );


  buf

  (
    g67_p_spl_,
    g67_p
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    G1_n_spl_00,
    G1_n_spl_0
  );


  buf

  (
    G1_n_spl_1,
    G1_n_spl_
  );


  buf

  (
    g67_n_spl_,
    g67_n
  );


  buf

  (
    g64_n_spl_,
    g64_n
  );


  buf

  (
    g64_n_spl_0,
    g64_n_spl_
  );


  buf

  (
    g64_n_spl_00,
    g64_n_spl_0
  );


  buf

  (
    g64_n_spl_01,
    g64_n_spl_0
  );


  buf

  (
    g64_n_spl_1,
    g64_n_spl_
  );


  buf

  (
    g70_n_spl_,
    g70_n
  );


  buf

  (
    g70_n_spl_0,
    g70_n_spl_
  );


  buf

  (
    g70_n_spl_1,
    g70_n_spl_
  );


  buf

  (
    g64_p_spl_,
    g64_p
  );


  buf

  (
    g64_p_spl_0,
    g64_p_spl_
  );


  buf

  (
    g64_p_spl_00,
    g64_p_spl_0
  );


  buf

  (
    g64_p_spl_01,
    g64_p_spl_0
  );


  buf

  (
    g64_p_spl_1,
    g64_p_spl_
  );


  buf

  (
    g70_p_spl_,
    g70_p
  );


  buf

  (
    g70_p_spl_0,
    g70_p_spl_
  );


  buf

  (
    g70_p_spl_1,
    g70_p_spl_
  );


  buf

  (
    g49_n_spl_,
    g49_n
  );


  buf

  (
    g73_n_spl_,
    g73_n
  );


  buf

  (
    g49_p_spl_,
    g49_p
  );


  buf

  (
    g73_p_spl_,
    g73_p
  );


  buf

  (
    g76_n_spl_,
    g76_n
  );


  buf

  (
    g76_p_spl_,
    g76_p
  );


  buf

  (
    G25_n_spl_,
    G25_n
  );


  buf

  (
    G25_n_spl_0,
    G25_n_spl_
  );


  buf

  (
    g77_p_spl_,
    g77_p
  );


  buf

  (
    G25_p_spl_,
    G25_p
  );


  buf

  (
    G25_p_spl_0,
    G25_p_spl_
  );


  buf

  (
    g77_n_spl_,
    g77_n
  );


  buf

  (
    g42_p_spl_,
    g42_p
  );


  buf

  (
    g42_p_spl_0,
    g42_p_spl_
  );


  buf

  (
    g80_n_spl_,
    g80_n
  );


  buf

  (
    g80_n_spl_0,
    g80_n_spl_
  );


  buf

  (
    g42_n_spl_,
    g42_n
  );


  buf

  (
    g80_p_spl_,
    g80_p
  );


  buf

  (
    G18_p_spl_,
    G18_p
  );


  buf

  (
    G18_n_spl_,
    G18_n
  );


  buf

  (
    g83_n_spl_,
    g83_n
  );


  buf

  (
    g83_p_spl_,
    g83_p
  );


  buf

  (
    g86_n_spl_,
    g86_n
  );


  buf

  (
    g86_p_spl_,
    g86_p
  );


  buf

  (
    G9_p_spl_,
    G9_p
  );


  buf

  (
    G9_p_spl_0,
    G9_p_spl_
  );


  buf

  (
    G9_p_spl_00,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_1,
    G9_p_spl_
  );


  buf

  (
    G9_n_spl_,
    G9_n
  );


  buf

  (
    G9_n_spl_0,
    G9_n_spl_
  );


  buf

  (
    G9_n_spl_00,
    G9_n_spl_0
  );


  buf

  (
    G9_n_spl_1,
    G9_n_spl_
  );


  buf

  (
    g92_n_spl_,
    g92_n
  );


  buf

  (
    g92_n_spl_0,
    g92_n_spl_
  );


  buf

  (
    g92_n_spl_1,
    g92_n_spl_
  );


  buf

  (
    g92_p_spl_,
    g92_p
  );


  buf

  (
    g92_p_spl_0,
    g92_p_spl_
  );


  buf

  (
    g92_p_spl_1,
    g92_p_spl_
  );


  buf

  (
    g89_p_spl_,
    g89_p
  );


  buf

  (
    g95_p_spl_,
    g95_p
  );


  buf

  (
    g95_p_spl_0,
    g95_p_spl_
  );


  buf

  (
    g95_p_spl_1,
    g95_p_spl_
  );


  buf

  (
    g89_n_spl_,
    g89_n
  );


  buf

  (
    g95_n_spl_,
    g95_n
  );


  buf

  (
    g95_n_spl_0,
    g95_n_spl_
  );


  buf

  (
    g95_n_spl_1,
    g95_n_spl_
  );


  buf

  (
    G5_n_spl_,
    G5_n
  );


  buf

  (
    G5_n_spl_0,
    G5_n_spl_
  );


  buf

  (
    G5_n_spl_00,
    G5_n_spl_0
  );


  buf

  (
    G5_n_spl_1,
    G5_n_spl_
  );


  buf

  (
    G8_n_spl_,
    G8_n
  );


  buf

  (
    G8_n_spl_0,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_00,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_01,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_1,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_10,
    G8_n_spl_1
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G5_p_spl_0,
    G5_p_spl_
  );


  buf

  (
    G5_p_spl_00,
    G5_p_spl_0
  );


  buf

  (
    G5_p_spl_1,
    G5_p_spl_
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_00,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_01,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_1,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_10,
    G8_p_spl_1
  );


  buf

  (
    g101_p_spl_,
    g101_p
  );


  buf

  (
    g101_n_spl_,
    g101_n
  );


  buf

  (
    g98_n_spl_,
    g98_n
  );


  buf

  (
    g104_p_spl_,
    g104_p
  );


  buf

  (
    g98_p_spl_,
    g98_p
  );


  buf

  (
    g104_n_spl_,
    g104_n
  );


  buf

  (
    g107_n_spl_,
    g107_n
  );


  buf

  (
    G27_n_spl_,
    G27_n
  );


  buf

  (
    G27_n_spl_0,
    G27_n_spl_
  );


  buf

  (
    g108_p_spl_,
    g108_p
  );


  buf

  (
    G27_p_spl_,
    G27_p
  );


  buf

  (
    g108_n_spl_,
    g108_n
  );


  buf

  (
    G6_n_spl_,
    G6_n
  );


  buf

  (
    G6_n_spl_0,
    G6_n_spl_
  );


  buf

  (
    G6_n_spl_00,
    G6_n_spl_0
  );


  buf

  (
    G6_n_spl_1,
    G6_n_spl_
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G6_p_spl_0,
    G6_p_spl_
  );


  buf

  (
    G6_p_spl_00,
    G6_p_spl_0
  );


  buf

  (
    G6_p_spl_1,
    G6_p_spl_
  );


  buf

  (
    g112_p_spl_,
    g112_p
  );


  buf

  (
    g112_n_spl_,
    g112_n
  );


  buf

  (
    g115_n_spl_,
    g115_n
  );


  buf

  (
    g118_n_spl_,
    g118_n
  );


  buf

  (
    g115_p_spl_,
    g115_p
  );


  buf

  (
    g118_p_spl_,
    g118_p
  );


  buf

  (
    G19_p_spl_,
    G19_p
  );


  buf

  (
    G19_n_spl_,
    G19_n
  );


  buf

  (
    g121_n_spl_,
    g121_n
  );


  buf

  (
    g123_n_spl_,
    g123_n
  );


  buf

  (
    g121_p_spl_,
    g121_p
  );


  buf

  (
    g123_p_spl_,
    g123_p
  );


  buf

  (
    g126_n_spl_,
    g126_n
  );


  buf

  (
    G28_n_spl_,
    G28_n
  );


  buf

  (
    G28_n_spl_0,
    G28_n_spl_
  );


  buf

  (
    g127_p_spl_,
    g127_p
  );


  buf

  (
    G28_p_spl_,
    G28_p
  );


  buf

  (
    g127_n_spl_,
    g127_n
  );


  buf

  (
    G7_n_spl_,
    G7_n
  );


  buf

  (
    G7_n_spl_0,
    G7_n_spl_
  );


  buf

  (
    G7_n_spl_00,
    G7_n_spl_0
  );


  buf

  (
    G7_n_spl_1,
    G7_n_spl_
  );


  buf

  (
    G7_p_spl_,
    G7_p
  );


  buf

  (
    G7_p_spl_0,
    G7_p_spl_
  );


  buf

  (
    G7_p_spl_00,
    G7_p_spl_0
  );


  buf

  (
    G7_p_spl_1,
    G7_p_spl_
  );


  buf

  (
    g133_p_spl_,
    g133_p
  );


  buf

  (
    g133_n_spl_,
    g133_n
  );


  buf

  (
    g136_n_spl_,
    g136_n
  );


  buf

  (
    g136_p_spl_,
    g136_p
  );


  buf

  (
    g141_p_spl_,
    g141_p
  );


  buf

  (
    g141_n_spl_,
    g141_n
  );


  buf

  (
    g139_n_spl_,
    g139_n
  );


  buf

  (
    g144_n_spl_,
    g144_n
  );


  buf

  (
    g139_p_spl_,
    g139_p
  );


  buf

  (
    g144_p_spl_,
    g144_p
  );


  buf

  (
    g147_n_spl_,
    g147_n
  );


  buf

  (
    g148_p_spl_,
    g148_p
  );


  buf

  (
    g149_n_spl_,
    g149_n
  );


  buf

  (
    g149_n_spl_0,
    g149_n_spl_
  );


  buf

  (
    g148_n_spl_,
    g148_n
  );


  buf

  (
    g149_p_spl_,
    g149_p
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    G17_n_spl_,
    G17_n
  );


  buf

  (
    g156_p_spl_,
    g156_p
  );


  buf

  (
    g156_n_spl_,
    g156_n
  );


  buf

  (
    g162_p_spl_,
    g162_p
  );


  buf

  (
    g162_n_spl_,
    g162_n
  );


  buf

  (
    g165_n_spl_,
    g165_n
  );


  buf

  (
    g165_n_spl_0,
    g165_n_spl_
  );


  buf

  (
    g165_n_spl_1,
    g165_n_spl_
  );


  buf

  (
    g165_p_spl_,
    g165_p
  );


  buf

  (
    g165_p_spl_0,
    g165_p_spl_
  );


  buf

  (
    g165_p_spl_1,
    g165_p_spl_
  );


  buf

  (
    g159_p_spl_,
    g159_p
  );


  buf

  (
    g168_p_spl_,
    g168_p
  );


  buf

  (
    g159_n_spl_,
    g159_n
  );


  buf

  (
    g168_n_spl_,
    g168_n
  );


  buf

  (
    g171_n_spl_,
    g171_n
  );


  buf

  (
    g171_p_spl_,
    g171_p
  );


  buf

  (
    G26_p_spl_,
    G26_p
  );


  buf

  (
    G26_p_spl_0,
    G26_p_spl_
  );


  buf

  (
    g172_n_spl_,
    g172_n
  );


  buf

  (
    G26_n_spl_,
    G26_n
  );


  buf

  (
    G26_n_spl_0,
    G26_n_spl_
  );


  buf

  (
    g172_p_spl_,
    g172_p
  );


  buf

  (
    g179_n_spl_,
    g179_n
  );


  buf

  (
    g179_p_spl_,
    g179_p
  );


  buf

  (
    G21_p_spl_,
    G21_p
  );


  buf

  (
    G21_n_spl_,
    G21_n
  );


  buf

  (
    g181_p_spl_,
    g181_p
  );


  buf

  (
    g184_p_spl_,
    g184_p
  );


  buf

  (
    g181_n_spl_,
    g181_n
  );


  buf

  (
    g184_n_spl_,
    g184_n
  );


  buf

  (
    g190_p_spl_,
    g190_p
  );


  buf

  (
    g193_n_spl_,
    g193_n
  );


  buf

  (
    g190_n_spl_,
    g190_n
  );


  buf

  (
    g193_p_spl_,
    g193_p
  );


  buf

  (
    g187_p_spl_,
    g187_p
  );


  buf

  (
    g196_n_spl_,
    g196_n
  );


  buf

  (
    g196_n_spl_0,
    g196_n_spl_
  );


  buf

  (
    g187_n_spl_,
    g187_n
  );


  buf

  (
    g196_p_spl_,
    g196_p
  );


  buf

  (
    g196_p_spl_0,
    g196_p_spl_
  );


  buf

  (
    g199_p_spl_,
    g199_p
  );


  buf

  (
    g199_n_spl_,
    g199_n
  );


  buf

  (
    g200_p_spl_,
    g200_p
  );


  buf

  (
    g201_n_spl_,
    g201_n
  );


  buf

  (
    g201_n_spl_0,
    g201_n_spl_
  );


  buf

  (
    g200_n_spl_,
    g200_n
  );


  buf

  (
    g201_p_spl_,
    g201_p
  );


  buf

  (
    g201_p_spl_0,
    g201_p_spl_
  );


  buf

  (
    g180_p_spl_,
    g180_p
  );


  buf

  (
    g180_p_spl_0,
    g180_p_spl_
  );


  buf

  (
    g204_n_spl_,
    g204_n
  );


  buf

  (
    g204_n_spl_0,
    g204_n_spl_
  );


  buf

  (
    g180_n_spl_,
    g180_n
  );


  buf

  (
    g204_p_spl_,
    g204_p
  );


  buf

  (
    g178_p_spl_,
    g178_p
  );


  buf

  (
    g178_n_spl_,
    g178_n
  );


  buf

  (
    g178_n_spl_0,
    g178_n_spl_
  );


  buf

  (
    g81_n_spl_,
    g81_n
  );


  buf

  (
    g206_p_spl_,
    g206_p
  );


  buf

  (
    g81_p_spl_,
    g81_p
  );


  buf

  (
    g206_n_spl_,
    g206_n
  );


  buf

  (
    g40_n_spl_,
    g40_n
  );


  buf

  (
    g207_p_spl_,
    g207_p
  );


  buf

  (
    g40_p_spl_,
    g40_p
  );


  buf

  (
    g207_n_spl_,
    g207_n
  );


  buf

  (
    g208_n_spl_,
    g208_n
  );


  buf

  (
    g208_n_spl_0,
    g208_n_spl_
  );


  buf

  (
    g208_n_spl_00,
    g208_n_spl_0
  );


  buf

  (
    g208_n_spl_01,
    g208_n_spl_0
  );


  buf

  (
    g208_n_spl_1,
    g208_n_spl_
  );


  buf

  (
    g208_n_spl_10,
    g208_n_spl_1
  );


  buf

  (
    g208_p_spl_,
    g208_p
  );


  buf

  (
    g208_p_spl_0,
    g208_p_spl_
  );


  buf

  (
    g208_p_spl_00,
    g208_p_spl_0
  );


  buf

  (
    g208_p_spl_01,
    g208_p_spl_0
  );


  buf

  (
    g208_p_spl_1,
    g208_p_spl_
  );


  buf

  (
    g208_p_spl_10,
    g208_p_spl_1
  );


  buf

  (
    G30_n_spl_,
    G30_n
  );


  buf

  (
    G30_p_spl_,
    G30_p
  );


  buf

  (
    g221_p_spl_,
    g221_p
  );


  buf

  (
    g221_n_spl_,
    g221_n
  );


  buf

  (
    g223_n_spl_,
    g223_n
  );


  buf

  (
    g223_n_spl_0,
    g223_n_spl_
  );


  buf

  (
    g223_p_spl_,
    g223_p
  );


  buf

  (
    g223_p_spl_0,
    g223_p_spl_
  );


  buf

  (
    g224_n_spl_,
    g224_n
  );


  buf

  (
    g224_n_spl_0,
    g224_n_spl_
  );


  buf

  (
    g224_n_spl_00,
    g224_n_spl_0
  );


  buf

  (
    g224_n_spl_01,
    g224_n_spl_0
  );


  buf

  (
    g224_n_spl_1,
    g224_n_spl_
  );


  buf

  (
    g224_p_spl_,
    g224_p
  );


  buf

  (
    g224_p_spl_0,
    g224_p_spl_
  );


  buf

  (
    g224_p_spl_00,
    g224_p_spl_0
  );


  buf

  (
    g224_p_spl_01,
    g224_p_spl_0
  );


  buf

  (
    g224_p_spl_1,
    g224_p_spl_
  );


  buf

  (
    g235_p_spl_,
    g235_p
  );


  buf

  (
    g235_n_spl_,
    g235_n
  );


  buf

  (
    g236_n_spl_,
    g236_n
  );


  buf

  (
    g236_n_spl_0,
    g236_n_spl_
  );


  buf

  (
    g236_n_spl_1,
    g236_n_spl_
  );


  buf

  (
    g236_p_spl_,
    g236_p
  );


  buf

  (
    g236_p_spl_0,
    g236_p_spl_
  );


  buf

  (
    g236_p_spl_1,
    g236_p_spl_
  );


  buf

  (
    g256_n_spl_,
    g256_n
  );


  buf

  (
    g256_n_spl_0,
    g256_n_spl_
  );


  buf

  (
    g256_n_spl_1,
    g256_n_spl_
  );


  buf

  (
    g256_p_spl_,
    g256_p
  );


  buf

  (
    g256_p_spl_0,
    g256_p_spl_
  );


  buf

  (
    g256_p_spl_1,
    g256_p_spl_
  );


  buf

  (
    g269_p_spl_,
    g269_p
  );


  buf

  (
    g269_p_spl_0,
    g269_p_spl_
  );


  buf

  (
    g269_p_spl_00,
    g269_p_spl_0
  );


  buf

  (
    g269_p_spl_01,
    g269_p_spl_0
  );


  buf

  (
    g269_p_spl_1,
    g269_p_spl_
  );


  buf

  (
    g269_p_spl_10,
    g269_p_spl_1
  );


  buf

  (
    g269_n_spl_,
    g269_n
  );


  buf

  (
    g269_n_spl_0,
    g269_n_spl_
  );


  buf

  (
    g303_n_spl_,
    g303_n
  );


  buf

  (
    g303_p_spl_,
    g303_p
  );


  buf

  (
    g315_n_spl_,
    g315_n
  );


  buf

  (
    g315_p_spl_,
    g315_p
  );


endmodule
