// Benchmark "mymod" written by ABC on Sun Oct 29 23:44:43 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33,
    G1884, G1885, G1886, G1887, G1888, G1889, G1890, G1891, G1892, G1893,
    G1894, G1895, G1896, G1897, G1898, G1899, G1900, G1901, G1902, G1903,
    G1904, G1905, G1906, G1907, G1908  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33;
  output G1884, G1885, G1886, G1887, G1888, G1889, G1890, G1891, G1892, G1893,
    G1894, G1895, G1896, G1897, G1898, G1899, G1900, G1901, G1902, G1903,
    G1904, G1905, G1906, G1907, G1908;
  reg n940_lo, n949_lo, n961_lo, n973_lo, n976_lo, n985_lo, n988_lo,
    n997_lo, n1009_lo, n1021_lo, n1033_lo, n1045_lo, n1057_lo, n1060_lo,
    n1069_lo, n1081_lo, n1093_lo, n1105_lo, n1117_lo, n1120_lo, n1129_lo,
    n1132_lo, n1156_lo, n1168_lo, n1180_lo, n1189_lo, n1192_lo, n1195_lo,
    n1201_lo, n1204_lo, n1228_lo, n1231_lo, n1234_lo, n1237_lo, n1240_lo,
    n1243_lo, n1249_lo, n1252_lo, n1255_lo, n1261_lo, n1264_lo, n1267_lo,
    n1273_lo, n1276_lo, n1279_lo, n1282_lo, n1285_lo, n1288_lo, n1291_lo,
    n1294_lo, n1297_lo, n1300_lo, n1303_lo, n1309_lo, n1312_lo, n1315_lo,
    n1318_lo, n1321_lo, n1333_lo, n1225_o2, n1229_o2, n1228_o2, n1259_o2,
    n1272_o2, n1269_o2, n1307_o2, n1201_o2, n1202_o2, n1203_o2, n1204_o2,
    n622_o2, n1205_o2, n1206_o2, n497_o2, n1212_o2, n1213_o2, n1214_o2,
    n1215_o2, n1216_o2, n1217_o2, n1218_o2, n1219_o2, n1242_o2, n1243_o2,
    n1273_o2, n1274_o2, n1275_o2, n1276_o2, n1277_o2, n1286_o2, n1299_o2,
    n601_o2, n625_o2, n463_o2, lo082_buf_o2, n455_o2, n642_o2, n459_o2,
    n501_o2, n599_o2, n485_o2, lo086_buf_o2, lo122_buf_o2, n502_o2,
    n627_o2, lo038_buf_o2, lo046_buf_o2, lo050_buf_o2, lo058_buf_o2,
    lo070_buf_o2, lo094_buf_o2, n462_o2, lo006_buf_o2, lo010_buf_o2,
    lo022_buf_o2, lo026_buf_o2, lo030_buf_o2, lo034_buf_o2, lo054_buf_o2,
    lo130_buf_o2, n547_o2, n424_inv, n617_o2, lo042_buf_o2, lo062_buf_o2,
    lo110_buf_o2, n733_o2, n734_o2, n570_o2, n461_o2, n644_o2, n628_o2,
    n528_o2, n460_inv, lo002_buf_o2, lo014_buf_o2, lo018_buf_o2,
    lo078_buf_o2, lo090_buf_o2, n513_o2, lo102_buf_o2, lo106_buf_o2,
    n600_o2, n529_o2, n593_o2, lo066_buf_o2, n549_o2, n550_o2, n571_o2,
    n572_o2, n495_o2, n496_o2, n620_o2, n482_o2, lo081_buf_o2, n576_o2,
    n520_o2, n521_o2, n562_o2, n508_o2, n509_o2, lo074_buf_o2, n539_o2,
    n536_o2, n516_o2, n491_o2, n557_o2, n586_o2, n483_o2, n484_o2,
    lo004_buf_o2, lo008_buf_o2, lo020_buf_o2, lo024_buf_o2, lo028_buf_o2,
    lo032_buf_o2, lo052_buf_o2, lo128_buf_o2, lo037_buf_o2, lo045_buf_o2,
    lo049_buf_o2, lo057_buf_o2, lo069_buf_o2, lo093_buf_o2;
  wire new_n427_, new_n429_, new_n431_, new_n433_, new_n435_, new_n437_,
    new_n439_, new_n441_, new_n443_, new_n445_, new_n447_, new_n449_,
    new_n451_, new_n453_, new_n455_, new_n457_, new_n459_, new_n461_,
    new_n463_, new_n465_, new_n467_, new_n469_, new_n471_, new_n473_,
    new_n475_, new_n477_, new_n479_, new_n481_, new_n483_, new_n485_,
    new_n487_, new_n489_, new_n491_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n537_, new_n539_,
    new_n541_, new_n543_, new_n544_, new_n545_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n555_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n563_,
    new_n566_, new_n567_, new_n569_, new_n571_, new_n573_, new_n575_,
    new_n576_, new_n577_, new_n579_, new_n581_, new_n583_, new_n585_,
    new_n586_, new_n587_, new_n589_, new_n591_, new_n593_, new_n594_,
    new_n595_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n603_, new_n605_, new_n607_, new_n609_, new_n610_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n617_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n629_, new_n631_,
    new_n633_, new_n634_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n645_, new_n647_, new_n649_, new_n651_,
    new_n653_, new_n655_, new_n657_, new_n659_, new_n661_, new_n663_,
    new_n665_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n713_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n737_, new_n739_, new_n741_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n786_, new_n788_, new_n789_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_,
    new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_,
    new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_,
    new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_,
    new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_,
    new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_,
    new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_,
    new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_,
    new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_,
    new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_,
    new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_,
    new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_,
    new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_,
    new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_,
    new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_,
    new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_,
    new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_,
    new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, n2248_li000_li000, n2257_li003_li003, n2269_li007_li007,
    n2281_li011_li011, n2284_li012_li012, n2293_li015_li015,
    n2296_li016_li016, n2305_li019_li019, n2317_li023_li023,
    n2329_li027_li027, n2341_li031_li031, n2353_li035_li035,
    n2365_li039_li039, n2368_li040_li040, n2377_li043_li043,
    n2389_li047_li047, n2401_li051_li051, n2413_li055_li055,
    n2425_li059_li059, n2428_li060_li060, n2437_li063_li063,
    n2440_li064_li064, n2464_li072_li072, n2476_li076_li076,
    n2488_li080_li080, n2497_li083_li083, n2500_li084_li084,
    n2503_li085_li085, n2509_li087_li087, n2512_li088_li088,
    n2536_li096_li096, n2539_li097_li097, n2542_li098_li098,
    n2545_li099_li099, n2548_li100_li100, n2551_li101_li101,
    n2557_li103_li103, n2560_li104_li104, n2563_li105_li105,
    n2569_li107_li107, n2572_li108_li108, n2575_li109_li109,
    n2581_li111_li111, n2584_li112_li112, n2587_li113_li113,
    n2590_li114_li114, n2593_li115_li115, n2596_li116_li116,
    n2599_li117_li117, n2602_li118_li118, n2605_li119_li119,
    n2608_li120_li120, n2611_li121_li121, n2617_li123_li123,
    n2620_li124_li124, n2623_li125_li125, n2626_li126_li126,
    n2629_li127_li127, n2641_li131_li131, n1225_i2, n1229_i2, n1228_i2,
    n1259_i2, n1272_i2, n1269_i2, n1307_i2, n1201_i2, n1202_i2, n1203_i2,
    n1204_i2, n622_i2, n1205_i2, n1206_i2, n497_i2, n1212_i2, n1213_i2,
    n1214_i2, n1215_i2, n1216_i2, n1217_i2, n1218_i2, n1219_i2, n1242_i2,
    n1243_i2, n1273_i2, n1274_i2, n1275_i2, n1276_i2, n1277_i2, n1286_i2,
    n1299_i2, n601_i2, n625_i2, n463_i2, lo082_buf_i2, n455_i2, n642_i2,
    n459_i2, n501_i2, n599_i2, n485_i2, lo086_buf_i2, lo122_buf_i2,
    n502_i2, n627_i2, lo038_buf_i2, lo046_buf_i2, lo050_buf_i2,
    lo058_buf_i2, lo070_buf_i2, lo094_buf_i2, n462_i2, lo006_buf_i2,
    lo010_buf_i2, lo022_buf_i2, lo026_buf_i2, lo030_buf_i2, lo034_buf_i2,
    lo054_buf_i2, lo130_buf_i2, n547_i2, n568_i2, n617_i2, lo042_buf_i2,
    lo062_buf_i2, lo110_buf_i2, n733_i2, n734_i2, n570_i2, n461_i2,
    n644_i2, n628_i2, n528_i2, n592_i2, lo002_buf_i2, lo014_buf_i2,
    lo018_buf_i2, lo078_buf_i2, lo090_buf_i2, n513_i2, lo102_buf_i2,
    lo106_buf_i2, n600_i2, n529_i2, n593_i2, lo066_buf_i2, n549_i2,
    n550_i2, n571_i2, n572_i2, n495_i2, n496_i2, n620_i2, n482_i2,
    lo081_buf_i2, n576_i2, n520_i2, n521_i2, n562_i2, n508_i2, n509_i2,
    lo074_buf_i2, n539_i2, n536_i2, n516_i2, n491_i2, n557_i2, n586_i2,
    n483_i2, n484_i2, lo004_buf_i2, lo008_buf_i2, lo020_buf_i2,
    lo024_buf_i2, lo028_buf_i2, lo032_buf_i2, lo052_buf_i2, lo128_buf_i2,
    lo037_buf_i2, lo045_buf_i2, lo049_buf_i2, lo057_buf_i2, lo069_buf_i2,
    lo093_buf_i2;
  assign new_n427_ = G1;
  assign new_n429_ = G2;
  assign new_n431_ = G3;
  assign new_n433_ = G4;
  assign new_n435_ = G5;
  assign new_n437_ = G6;
  assign new_n439_ = G7;
  assign new_n441_ = G8;
  assign new_n443_ = G9;
  assign new_n445_ = G10;
  assign new_n447_ = G11;
  assign new_n449_ = G12;
  assign new_n451_ = G13;
  assign new_n453_ = G14;
  assign new_n455_ = G15;
  assign new_n457_ = G16;
  assign new_n459_ = G17;
  assign new_n461_ = G18;
  assign new_n463_ = G19;
  assign new_n465_ = G20;
  assign new_n467_ = G21;
  assign new_n469_ = G22;
  assign new_n471_ = G23;
  assign new_n473_ = G24;
  assign new_n475_ = G25;
  assign new_n477_ = G26;
  assign new_n479_ = G27;
  assign new_n481_ = G28;
  assign new_n483_ = G29;
  assign new_n485_ = G30;
  assign new_n487_ = G31;
  assign new_n489_ = G32;
  assign new_n491_ = G33;
  assign new_n493_ = n940_lo;
  assign new_n494_ = ~n940_lo;
  assign new_n495_ = n949_lo;
  assign new_n496_ = ~n949_lo;
  assign new_n497_ = n961_lo;
  assign new_n498_ = ~n961_lo;
  assign new_n499_ = n973_lo;
  assign new_n500_ = ~n973_lo;
  assign new_n501_ = n976_lo;
  assign new_n502_ = ~n976_lo;
  assign new_n503_ = n985_lo;
  assign new_n504_ = ~n985_lo;
  assign new_n505_ = n988_lo;
  assign new_n506_ = ~n988_lo;
  assign new_n507_ = n997_lo;
  assign new_n508_ = ~n997_lo;
  assign new_n509_ = n1009_lo;
  assign new_n510_ = ~n1009_lo;
  assign new_n511_ = n1021_lo;
  assign new_n512_ = ~n1021_lo;
  assign new_n513_ = n1033_lo;
  assign new_n514_ = ~n1033_lo;
  assign new_n515_ = n1045_lo;
  assign new_n516_ = ~n1045_lo;
  assign new_n517_ = n1057_lo;
  assign new_n518_ = ~n1057_lo;
  assign new_n519_ = n1060_lo;
  assign new_n520_ = ~n1060_lo;
  assign new_n521_ = n1069_lo;
  assign new_n522_ = ~n1069_lo;
  assign new_n523_ = n1081_lo;
  assign new_n524_ = ~n1081_lo;
  assign new_n525_ = n1093_lo;
  assign new_n526_ = ~n1093_lo;
  assign new_n527_ = n1105_lo;
  assign new_n528_ = ~n1105_lo;
  assign new_n529_ = n1117_lo;
  assign new_n530_ = ~n1117_lo;
  assign new_n531_ = n1120_lo;
  assign new_n532_ = ~n1120_lo;
  assign new_n533_ = n1129_lo;
  assign new_n534_ = ~n1129_lo;
  assign new_n535_ = n1132_lo;
  assign new_n537_ = n1156_lo;
  assign new_n539_ = n1168_lo;
  assign new_n541_ = n1180_lo;
  assign new_n543_ = n1189_lo;
  assign new_n544_ = ~n1189_lo;
  assign new_n545_ = n1192_lo;
  assign new_n547_ = n1195_lo;
  assign new_n548_ = ~n1195_lo;
  assign new_n549_ = n1201_lo;
  assign new_n550_ = ~n1201_lo;
  assign new_n551_ = n1204_lo;
  assign new_n552_ = ~n1204_lo;
  assign new_n553_ = n1228_lo;
  assign new_n555_ = n1231_lo;
  assign new_n557_ = n1234_lo;
  assign new_n558_ = ~n1234_lo;
  assign new_n559_ = n1237_lo;
  assign new_n560_ = ~n1237_lo;
  assign new_n561_ = n1240_lo;
  assign new_n563_ = n1243_lo;
  assign new_n566_ = ~n1249_lo;
  assign new_n567_ = n1252_lo;
  assign new_n569_ = n1255_lo;
  assign new_n571_ = n1261_lo;
  assign new_n573_ = n1264_lo;
  assign new_n575_ = n1267_lo;
  assign new_n576_ = ~n1267_lo;
  assign new_n577_ = n1273_lo;
  assign new_n579_ = n1276_lo;
  assign new_n581_ = n1279_lo;
  assign new_n583_ = n1282_lo;
  assign new_n585_ = n1285_lo;
  assign new_n586_ = ~n1285_lo;
  assign new_n587_ = n1288_lo;
  assign new_n589_ = n1291_lo;
  assign new_n591_ = n1294_lo;
  assign new_n593_ = n1297_lo;
  assign new_n594_ = ~n1297_lo;
  assign new_n595_ = n1300_lo;
  assign new_n597_ = n1303_lo;
  assign new_n598_ = ~n1303_lo;
  assign new_n599_ = n1309_lo;
  assign new_n600_ = ~n1309_lo;
  assign new_n601_ = n1312_lo;
  assign new_n603_ = n1315_lo;
  assign new_n605_ = n1318_lo;
  assign new_n607_ = n1321_lo;
  assign new_n609_ = n1333_lo;
  assign new_n610_ = ~n1333_lo;
  assign new_n612_ = ~n1225_o2;
  assign new_n613_ = n1229_o2;
  assign new_n614_ = ~n1229_o2;
  assign new_n615_ = n1228_o2;
  assign new_n617_ = n1259_o2;
  assign new_n620_ = ~n1272_o2;
  assign new_n622_ = ~n1269_o2;
  assign new_n623_ = n1307_o2;
  assign new_n624_ = ~n1307_o2;
  assign new_n625_ = n1201_o2;
  assign new_n627_ = n1202_o2;
  assign new_n629_ = n1203_o2;
  assign new_n631_ = n1204_o2;
  assign new_n633_ = n622_o2;
  assign new_n634_ = ~n622_o2;
  assign new_n636_ = ~n1205_o2;
  assign new_n637_ = n1206_o2;
  assign new_n639_ = n497_o2;
  assign new_n640_ = ~n497_o2;
  assign new_n641_ = n1212_o2;
  assign new_n643_ = n1213_o2;
  assign new_n645_ = n1214_o2;
  assign new_n647_ = n1215_o2;
  assign new_n649_ = n1216_o2;
  assign new_n651_ = n1217_o2;
  assign new_n653_ = n1218_o2;
  assign new_n655_ = n1219_o2;
  assign new_n657_ = n1242_o2;
  assign new_n659_ = n1243_o2;
  assign new_n661_ = n1273_o2;
  assign new_n663_ = n1274_o2;
  assign new_n665_ = n1275_o2;
  assign new_n668_ = ~n1276_o2;
  assign new_n670_ = ~n1277_o2;
  assign new_n671_ = n1286_o2;
  assign new_n672_ = ~n1286_o2;
  assign new_n673_ = n1299_o2;
  assign new_n674_ = ~n1299_o2;
  assign new_n675_ = n601_o2;
  assign new_n676_ = ~n601_o2;
  assign new_n677_ = n625_o2;
  assign new_n678_ = ~n625_o2;
  assign new_n679_ = n463_o2;
  assign new_n680_ = ~n463_o2;
  assign new_n681_ = lo082_buf_o2;
  assign new_n683_ = n455_o2;
  assign new_n684_ = ~n455_o2;
  assign new_n685_ = n642_o2;
  assign new_n686_ = ~n642_o2;
  assign new_n687_ = n459_o2;
  assign new_n689_ = n501_o2;
  assign new_n690_ = ~n501_o2;
  assign new_n691_ = n599_o2;
  assign new_n692_ = ~n599_o2;
  assign new_n693_ = n485_o2;
  assign new_n694_ = ~n485_o2;
  assign new_n695_ = lo086_buf_o2;
  assign new_n697_ = lo122_buf_o2;
  assign new_n698_ = ~lo122_buf_o2;
  assign new_n699_ = n502_o2;
  assign new_n700_ = ~n502_o2;
  assign new_n701_ = n627_o2;
  assign new_n702_ = ~n627_o2;
  assign new_n703_ = lo038_buf_o2;
  assign new_n705_ = lo046_buf_o2;
  assign new_n707_ = lo050_buf_o2;
  assign new_n708_ = ~lo050_buf_o2;
  assign new_n709_ = lo058_buf_o2;
  assign new_n711_ = lo070_buf_o2;
  assign new_n713_ = lo094_buf_o2;
  assign new_n716_ = ~n462_o2;
  assign new_n717_ = lo006_buf_o2;
  assign new_n718_ = ~lo006_buf_o2;
  assign new_n719_ = lo010_buf_o2;
  assign new_n721_ = lo022_buf_o2;
  assign new_n723_ = lo026_buf_o2;
  assign new_n725_ = lo030_buf_o2;
  assign new_n726_ = ~lo030_buf_o2;
  assign new_n727_ = lo034_buf_o2;
  assign new_n728_ = ~lo034_buf_o2;
  assign new_n729_ = lo054_buf_o2;
  assign new_n730_ = ~lo054_buf_o2;
  assign new_n731_ = lo130_buf_o2;
  assign new_n732_ = ~lo130_buf_o2;
  assign new_n733_ = n547_o2;
  assign new_n735_ = n424_inv;
  assign new_n737_ = n617_o2;
  assign new_n739_ = lo042_buf_o2;
  assign new_n741_ = lo062_buf_o2;
  assign new_n743_ = lo110_buf_o2;
  assign new_n745_ = n733_o2;
  assign new_n746_ = ~n733_o2;
  assign new_n747_ = n734_o2;
  assign new_n748_ = ~n734_o2;
  assign new_n749_ = n570_o2;
  assign new_n751_ = n461_o2;
  assign new_n752_ = ~n461_o2;
  assign new_n753_ = n644_o2;
  assign new_n754_ = ~n644_o2;
  assign new_n755_ = n628_o2;
  assign new_n756_ = ~n628_o2;
  assign new_n757_ = n528_o2;
  assign new_n759_ = n460_inv;
  assign new_n761_ = lo002_buf_o2;
  assign new_n762_ = ~lo002_buf_o2;
  assign new_n763_ = lo014_buf_o2;
  assign new_n764_ = ~lo014_buf_o2;
  assign new_n765_ = lo018_buf_o2;
  assign new_n767_ = lo078_buf_o2;
  assign new_n769_ = lo090_buf_o2;
  assign new_n770_ = ~lo090_buf_o2;
  assign new_n771_ = n513_o2;
  assign new_n773_ = lo102_buf_o2;
  assign new_n774_ = ~lo102_buf_o2;
  assign new_n775_ = lo106_buf_o2;
  assign new_n776_ = ~lo106_buf_o2;
  assign new_n777_ = n600_o2;
  assign new_n778_ = ~n600_o2;
  assign new_n779_ = n529_o2;
  assign new_n780_ = ~n529_o2;
  assign new_n781_ = n593_o2;
  assign new_n782_ = ~n593_o2;
  assign new_n783_ = lo066_buf_o2;
  assign new_n786_ = ~n549_o2;
  assign new_n788_ = ~n550_o2;
  assign new_n789_ = n571_o2;
  assign new_n792_ = ~n572_o2;
  assign new_n793_ = n495_o2;
  assign new_n794_ = ~n495_o2;
  assign new_n795_ = n496_o2;
  assign new_n796_ = ~n496_o2;
  assign new_n797_ = n620_o2;
  assign new_n798_ = ~n620_o2;
  assign new_n799_ = n482_o2;
  assign new_n800_ = ~n482_o2;
  assign new_n801_ = lo081_buf_o2;
  assign new_n802_ = ~lo081_buf_o2;
  assign new_n803_ = n576_o2;
  assign new_n804_ = ~n576_o2;
  assign new_n805_ = n520_o2;
  assign new_n806_ = ~n520_o2;
  assign new_n807_ = n521_o2;
  assign new_n808_ = ~n521_o2;
  assign new_n809_ = n562_o2;
  assign new_n810_ = ~n562_o2;
  assign new_n811_ = n508_o2;
  assign new_n812_ = ~n508_o2;
  assign new_n813_ = n509_o2;
  assign new_n814_ = ~n509_o2;
  assign new_n815_ = lo074_buf_o2;
  assign new_n816_ = ~lo074_buf_o2;
  assign new_n817_ = n539_o2;
  assign new_n818_ = ~n539_o2;
  assign new_n819_ = n536_o2;
  assign new_n820_ = ~n536_o2;
  assign new_n821_ = n516_o2;
  assign new_n822_ = ~n516_o2;
  assign new_n823_ = n491_o2;
  assign new_n824_ = ~n491_o2;
  assign new_n825_ = n557_o2;
  assign new_n826_ = ~n557_o2;
  assign new_n827_ = n586_o2;
  assign new_n828_ = ~n586_o2;
  assign new_n829_ = n483_o2;
  assign new_n830_ = ~n483_o2;
  assign new_n831_ = n484_o2;
  assign new_n832_ = ~n484_o2;
  assign new_n833_ = lo004_buf_o2;
  assign new_n834_ = ~lo004_buf_o2;
  assign new_n835_ = lo008_buf_o2;
  assign new_n836_ = ~lo008_buf_o2;
  assign new_n837_ = lo020_buf_o2;
  assign new_n838_ = ~lo020_buf_o2;
  assign new_n839_ = lo024_buf_o2;
  assign new_n840_ = ~lo024_buf_o2;
  assign new_n841_ = lo028_buf_o2;
  assign new_n842_ = ~lo028_buf_o2;
  assign new_n843_ = lo032_buf_o2;
  assign new_n844_ = ~lo032_buf_o2;
  assign new_n845_ = lo052_buf_o2;
  assign new_n846_ = ~lo052_buf_o2;
  assign new_n847_ = lo128_buf_o2;
  assign new_n848_ = ~lo128_buf_o2;
  assign new_n849_ = lo037_buf_o2;
  assign new_n850_ = ~lo037_buf_o2;
  assign new_n851_ = lo045_buf_o2;
  assign new_n852_ = ~lo045_buf_o2;
  assign new_n853_ = lo049_buf_o2;
  assign new_n854_ = ~lo049_buf_o2;
  assign new_n855_ = lo057_buf_o2;
  assign new_n856_ = ~lo057_buf_o2;
  assign new_n857_ = lo069_buf_o2;
  assign new_n858_ = ~lo069_buf_o2;
  assign new_n859_ = lo093_buf_o2;
  assign new_n860_ = ~lo093_buf_o2;
  assign new_n861_ = new_n1464_ & new_n1465_;
  assign new_n862_ = new_n1466_ | new_n1467_;
  assign new_n863_ = new_n1470_ & new_n496_;
  assign new_n864_ = new_n1476_ & new_n495_;
  assign new_n865_ = new_n864_ | new_n863_;
  assign new_n866_ = new_n1470_ & new_n498_;
  assign new_n867_ = new_n1476_ & new_n497_;
  assign new_n868_ = new_n867_ | new_n866_;
  assign new_n869_ = new_n1471_ & new_n500_;
  assign new_n870_ = new_n1477_ & new_n499_;
  assign new_n871_ = new_n870_ | new_n869_;
  assign new_n872_ = new_n1471_ & new_n504_;
  assign new_n873_ = new_n1477_ & new_n503_;
  assign new_n874_ = new_n873_ | new_n872_;
  assign new_n875_ = new_n1464_ & new_n1481_;
  assign new_n876_ = new_n1466_ | new_n1483_;
  assign new_n877_ = new_n1486_ & new_n518_;
  assign new_n878_ = new_n1491_ & new_n517_;
  assign new_n879_ = new_n878_ | new_n877_;
  assign new_n880_ = new_n1486_ & new_n530_;
  assign new_n881_ = new_n1491_ & new_n529_;
  assign new_n882_ = new_n881_ | new_n880_;
  assign new_n883_ = new_n1487_ & new_n534_;
  assign new_n884_ = new_n1492_ & new_n533_;
  assign new_n885_ = new_n884_ | new_n883_;
  assign new_n886_ = new_n1494_ & new_n679_;
  assign new_n887_ = new_n689_ | new_n1495_;
  assign new_n888_ = new_n886_ & new_n701_;
  assign new_n889_ = new_n887_ | new_n702_;
  assign new_n890_ = new_n1496_ & new_n1465_;
  assign new_n891_ = new_n1497_ | new_n1467_;
  assign new_n892_ = new_n1499_ & new_n508_;
  assign new_n893_ = new_n1502_ & new_n507_;
  assign new_n894_ = new_n893_ | new_n892_;
  assign new_n895_ = new_n1499_ & new_n510_;
  assign new_n896_ = new_n1502_ & new_n509_;
  assign new_n897_ = new_n896_ | new_n895_;
  assign new_n898_ = new_n1500_ & new_n512_;
  assign new_n899_ = new_n1503_ & new_n511_;
  assign new_n900_ = new_n899_ | new_n898_;
  assign new_n901_ = new_n1500_ & new_n514_;
  assign new_n902_ = new_n1503_ & new_n513_;
  assign new_n903_ = new_n902_ | new_n901_;
  assign new_n904_ = new_n1496_ & new_n1481_;
  assign new_n905_ = new_n1497_ | new_n1483_;
  assign new_n906_ = new_n904_ & new_n515_;
  assign new_n907_ = new_n905_ & new_n516_;
  assign new_n908_ = new_n907_ | new_n906_;
  assign new_n909_ = new_n1480_ & new_n675_;
  assign new_n910_ = new_n1482_ | new_n1504_;
  assign new_n911_ = new_n909_ & new_n1505_;
  assign new_n912_ = new_n910_ | new_n678_;
  assign new_n913_ = new_n911_ & new_n700_;
  assign new_n914_ = new_n912_ | new_n699_;
  assign new_n915_ = new_n913_ & new_n1506_;
  assign new_n916_ = new_n914_ | new_n692_;
  assign new_n917_ = new_n1508_ & new_n522_;
  assign new_n918_ = new_n1511_ & new_n521_;
  assign new_n919_ = new_n918_ | new_n917_;
  assign new_n920_ = new_n1508_ & new_n524_;
  assign new_n921_ = new_n1511_ & new_n523_;
  assign new_n922_ = new_n921_ | new_n920_;
  assign new_n923_ = new_n1509_ & new_n526_;
  assign new_n924_ = new_n1512_ & new_n525_;
  assign new_n925_ = new_n924_ | new_n923_;
  assign new_n926_ = new_n1509_ & new_n528_;
  assign new_n927_ = new_n1512_ & new_n527_;
  assign new_n928_ = new_n927_ | new_n926_;
  assign new_n929_ = new_n1487_ & new_n1473_;
  assign new_n930_ = new_n1492_ | new_n1479_;
  assign new_n931_ = new_n1515_ & new_n607_;
  assign new_n932_ = new_n1495_ & new_n1504_;
  assign new_n933_ = new_n932_ & new_n1494_;
  assign new_n934_ = new_n933_ & new_n1505_;
  assign new_n935_ = new_n934_ & new_n1506_;
  assign new_n936_ = new_n935_ | new_n1519_;
  assign new_n937_ = new_n936_ | new_n931_;
  assign new_n938_ = new_n633_ & new_n1522_;
  assign new_n939_ = new_n634_ | new_n1525_;
  assign new_n940_ = new_n938_ & new_n1515_;
  assign new_n941_ = new_n939_ | new_n1527_;
  assign new_n942_ = new_n941_ & new_n624_;
  assign new_n943_ = new_n940_ & new_n623_;
  assign new_n944_ = new_n943_ | new_n942_;
  assign new_n945_ = new_n944_ & new_n1530_;
  assign new_n946_ = new_n1522_ & new_n559_;
  assign new_n947_ = new_n1525_ | new_n560_;
  assign new_n948_ = new_n946_ & new_n1516_;
  assign new_n949_ = new_n947_ | new_n1527_;
  assign new_n950_ = new_n949_ & new_n639_;
  assign new_n951_ = new_n948_ & new_n640_;
  assign new_n952_ = new_n951_ | new_n950_;
  assign new_n953_ = new_n952_ & new_n1530_;
  assign new_n954_ = new_n1521_ & new_n571_;
  assign new_n955_ = new_n954_ & new_n1516_;
  assign new_n956_ = new_n955_ | new_n622_;
  assign new_n957_ = new_n956_ & new_n1531_;
  assign new_n958_ = new_n1523_ & new_n577_;
  assign new_n959_ = new_n958_ & new_n1517_;
  assign new_n960_ = new_n959_ | new_n612_;
  assign new_n961_ = new_n960_ & new_n1531_;
  assign new_n962_ = new_n617_ & new_n1523_;
  assign new_n963_ = new_n962_ & new_n1517_;
  assign new_n964_ = new_n963_ | new_n615_;
  assign new_n965_ = new_n964_ & new_n1532_;
  assign new_n966_ = new_n585_ & new_n543_;
  assign new_n967_ = new_n586_ | new_n544_;
  assign new_n968_ = new_n967_ & new_n1533_;
  assign new_n969_ = new_n966_ | new_n1519_;
  assign new_n970_ = new_n683_ & new_n613_;
  assign new_n971_ = new_n684_ | new_n614_;
  assign new_n972_ = new_n1534_ & new_n1479_;
  assign new_n973_ = new_n1535_ | new_n1473_;
  assign new_n974_ = new_n1535_ & new_n1472_;
  assign new_n975_ = new_n1534_ | new_n1478_;
  assign new_n976_ = new_n975_ & new_n973_;
  assign new_n977_ = new_n974_ | new_n972_;
  assign new_n978_ = new_n977_ & new_n969_;
  assign new_n979_ = new_n976_ & new_n968_;
  assign new_n980_ = new_n979_ | new_n978_;
  assign new_n981_ = new_n593_ & new_n549_;
  assign new_n982_ = new_n594_ | new_n550_;
  assign new_n983_ = new_n982_ & new_n1533_;
  assign new_n984_ = new_n981_ | new_n1518_;
  assign new_n985_ = new_n748_ & new_n746_;
  assign new_n986_ = new_n747_ | new_n745_;
  assign new_n987_ = new_n986_ & new_n685_;
  assign new_n988_ = new_n985_ | new_n686_;
  assign new_n989_ = new_n1536_ & new_n1493_;
  assign new_n990_ = new_n1537_ | new_n1488_;
  assign new_n991_ = new_n1537_ & new_n1488_;
  assign new_n992_ = new_n1536_ | new_n1493_;
  assign new_n993_ = new_n992_ & new_n990_;
  assign new_n994_ = new_n991_ | new_n989_;
  assign new_n995_ = new_n994_ & new_n984_;
  assign new_n996_ = new_n993_ & new_n983_;
  assign new_n997_ = new_n996_ | new_n995_;
  assign new_n998_ = new_n1524_ | new_n566_;
  assign new_n999_ = new_n998_ | new_n1526_;
  assign new_n1000_ = new_n999_ & new_n620_;
  assign new_n1001_ = new_n1000_ & new_n1532_;
  assign new_n1002_ = new_n777_ & new_n673_;
  assign new_n1003_ = new_n1538_ | new_n674_;
  assign new_n1004_ = new_n796_ & new_n794_;
  assign new_n1005_ = new_n795_ | new_n793_;
  assign new_n1006_ = new_n1538_ | new_n636_;
  assign new_n1007_ = new_n798_ & new_n1539_;
  assign new_n1008_ = new_n1540_ | new_n1542_;
  assign new_n1009_ = new_n1008_ | new_n1544_;
  assign new_n1010_ = new_n1007_ | new_n1003_;
  assign new_n1011_ = new_n1010_ & new_n1009_;
  assign new_n1012_ = new_n716_ | new_n668_;
  assign new_n1013_ = new_n1546_ | new_n1548_;
  assign new_n1014_ = new_n1546_ | new_n1549_;
  assign new_n1015_ = new_n1547_ | new_n1550_;
  assign new_n1016_ = new_n1551_ & new_n1539_;
  assign new_n1017_ = new_n1004_ | new_n1542_;
  assign new_n1018_ = new_n1017_ | new_n1552_;
  assign new_n1019_ = new_n1016_ | new_n558_;
  assign new_n1020_ = new_n1019_ & new_n1018_;
  assign new_n1021_ = new_n780_ | new_n1553_;
  assign new_n1022_ = new_n788_ & new_n786_;
  assign new_n1023_ = new_n792_ & new_n789_;
  assign new_n1024_ = new_n1023_ & new_n1022_;
  assign new_n1025_ = new_n1024_ & new_n1021_;
  assign new_n1026_ = new_n782_ | new_n774_;
  assign new_n1027_ = new_n781_ | new_n1554_;
  assign new_n1028_ = new_n779_ | new_n776_;
  assign new_n1029_ = new_n1028_ & new_n1027_;
  assign new_n1030_ = new_n1029_ & new_n1026_;
  assign new_n1031_ = new_n1030_ & new_n1025_;
  assign new_n1032_ = new_n832_ & new_n830_;
  assign new_n1033_ = new_n831_ | new_n829_;
  assign new_n1034_ = new_n1555_ | new_n1556_;
  assign new_n1035_ = new_n1557_ | new_n1558_;
  assign new_n1036_ = new_n1035_ & new_n1559_;
  assign new_n1037_ = new_n1561_ | new_n1563_;
  assign new_n1038_ = new_n1565_ & new_n1566_;
  assign new_n1039_ = new_n1567_ | new_n1568_;
  assign new_n1040_ = new_n1567_ & new_n1568_;
  assign new_n1041_ = new_n1565_ | new_n1566_;
  assign new_n1042_ = new_n1041_ & new_n1039_;
  assign new_n1043_ = new_n1040_ | new_n1038_;
  assign new_n1044_ = new_n1569_ & new_n770_;
  assign new_n1045_ = new_n816_ | new_n1561_;
  assign new_n1046_ = new_n1044_ & new_n1571_;
  assign new_n1047_ = new_n1045_ | new_n1575_;
  assign new_n1048_ = new_n1047_ & new_n1043_;
  assign new_n1049_ = new_n1046_ & new_n1042_;
  assign new_n1050_ = new_n1049_ | new_n1048_;
  assign new_n1051_ = new_n1577_ & new_n1579_;
  assign new_n1052_ = new_n1581_ | new_n1583_;
  assign new_n1053_ = new_n1581_ & new_n1583_;
  assign new_n1054_ = new_n1577_ | new_n1579_;
  assign new_n1055_ = new_n1054_ & new_n1052_;
  assign new_n1056_ = new_n1053_ | new_n1051_;
  assign new_n1057_ = new_n1585_ & new_n1586_;
  assign new_n1058_ = new_n1587_ | new_n1589_;
  assign new_n1059_ = new_n1587_ & new_n1589_;
  assign new_n1060_ = new_n1585_ | new_n1586_;
  assign new_n1061_ = new_n1060_ & new_n1058_;
  assign new_n1062_ = new_n1059_ | new_n1057_;
  assign new_n1063_ = new_n1061_ | new_n1055_;
  assign new_n1064_ = new_n1062_ | new_n1056_;
  assign new_n1065_ = new_n1064_ & new_n1063_;
  assign new_n1066_ = new_n1591_ & new_n1594_;
  assign new_n1067_ = new_n1596_ | new_n1599_;
  assign new_n1068_ = new_n1596_ & new_n1599_;
  assign new_n1069_ = new_n1591_ | new_n1594_;
  assign new_n1070_ = new_n1069_ & new_n1067_;
  assign new_n1071_ = new_n1068_ | new_n1066_;
  assign new_n1072_ = new_n1602_ & new_n1604_;
  assign new_n1073_ = new_n1606_ | new_n1609_;
  assign new_n1074_ = new_n1606_ & new_n1609_;
  assign new_n1075_ = new_n1602_ | new_n1604_;
  assign new_n1076_ = new_n1075_ & new_n1073_;
  assign new_n1077_ = new_n1074_ | new_n1072_;
  assign new_n1078_ = new_n1610_ & new_n1611_;
  assign new_n1079_ = new_n1612_ | new_n1613_;
  assign new_n1080_ = new_n1612_ & new_n1613_;
  assign new_n1081_ = new_n1610_ | new_n1611_;
  assign new_n1082_ = new_n1081_ & new_n1079_;
  assign new_n1083_ = new_n1080_ | new_n1078_;
  assign new_n1084_ = new_n693_ & new_n672_;
  assign new_n1085_ = new_n694_ & new_n671_;
  assign new_n1086_ = new_n1614_ & new_n1569_;
  assign new_n1087_ = new_n670_ & new_n637_;
  assign new_n1088_ = new_n1615_ | new_n1543_;
  assign new_n1089_ = new_n1616_ | new_n1617_;
  assign new_n1090_ = new_n1615_ | new_n1618_;
  assign new_n1091_ = new_n1619_ & new_n1089_;
  assign new_n1092_ = new_n1616_ | new_n1620_;
  assign new_n1093_ = new_n1092_ & new_n1619_;
  assign new_n1094_ = new_n1621_ & new_n1622_;
  assign new_n1095_ = new_n814_ & new_n812_;
  assign new_n1096_ = new_n813_ | new_n811_;
  assign new_n1097_ = new_n1623_ & new_n1584_;
  assign new_n1098_ = new_n1624_ | new_n1580_;
  assign new_n1099_ = new_n1624_ & new_n1580_;
  assign new_n1100_ = new_n1623_ | new_n1584_;
  assign new_n1101_ = new_n1100_ & new_n1098_;
  assign new_n1102_ = new_n1099_ | new_n1097_;
  assign new_n1103_ = new_n808_ & new_n806_;
  assign new_n1104_ = new_n807_ | new_n805_;
  assign new_n1105_ = new_n1625_ & new_n1626_;
  assign new_n1106_ = new_n1627_ | new_n1629_;
  assign new_n1107_ = new_n1627_ & new_n1629_;
  assign new_n1108_ = new_n1625_ | new_n1626_;
  assign new_n1109_ = new_n1108_ & new_n1106_;
  assign new_n1110_ = new_n1107_ | new_n1105_;
  assign new_n1111_ = new_n1109_ & new_n1102_;
  assign new_n1112_ = new_n1110_ & new_n1101_;
  assign new_n1113_ = new_n1112_ | new_n1111_;
  assign new_n1114_ = new_n803_ & new_n1571_;
  assign new_n1115_ = new_n804_ | new_n1575_;
  assign new_n1116_ = new_n1630_ & new_n1632_;
  assign new_n1117_ = new_n1633_ | new_n1634_;
  assign new_n1118_ = new_n1633_ & new_n1634_;
  assign new_n1119_ = new_n1630_ | new_n1632_;
  assign new_n1120_ = new_n1119_ & new_n1117_;
  assign new_n1121_ = new_n1118_ | new_n1116_;
  assign new_n1122_ = new_n1636_ & new_n1592_;
  assign new_n1123_ = new_n1638_ | new_n1597_;
  assign new_n1124_ = new_n1638_ & new_n1597_;
  assign new_n1125_ = new_n1636_ | new_n1592_;
  assign new_n1126_ = new_n1125_ & new_n1123_;
  assign new_n1127_ = new_n1124_ | new_n1122_;
  assign new_n1128_ = new_n1127_ & new_n1120_;
  assign new_n1129_ = new_n1126_ & new_n1121_;
  assign new_n1130_ = new_n1129_ | new_n1128_;
  assign new_n1131_ = new_n1640_ & new_n1641_;
  assign new_n1132_ = new_n1643_ | new_n1645_;
  assign new_n1133_ = new_n1643_ & new_n1645_;
  assign new_n1134_ = new_n1640_ | new_n1641_;
  assign new_n1135_ = new_n1134_ & new_n1132_;
  assign new_n1136_ = new_n1133_ | new_n1131_;
  assign new_n1137_ = new_n1646_ | new_n1563_;
  assign new_n1138_ = new_n1647_ & new_n1649_;
  assign new_n1139_ = new_n1650_ & new_n1649_;
  assign new_n1140_ = new_n1651_ & new_n1648_;
  assign new_n1141_ = new_n1652_ & new_n1653_;
  assign new_n1142_ = new_n1652_ | new_n1653_;
  assign new_n1143_ = new_n1654_ | new_n1564_;
  assign new_n1144_ = new_n1655_ | new_n1657_;
  assign new_n1145_ = new_n1655_ & new_n1657_;
  assign new_n1146_ = new_n1572_ & new_n1658_;
  assign new_n1147_ = new_n1574_ | new_n548_;
  assign new_n1148_ = new_n1607_ & new_n1659_;
  assign new_n1149_ = new_n1601_ | new_n1661_;
  assign new_n1150_ = new_n1603_ & new_n1661_;
  assign new_n1151_ = new_n1607_ | new_n1659_;
  assign new_n1152_ = new_n1151_ & new_n1149_;
  assign new_n1153_ = new_n1150_ | new_n1148_;
  assign new_n1154_ = new_n1153_ & new_n1146_;
  assign new_n1155_ = new_n1152_ & new_n1147_;
  assign new_n1156_ = new_n1155_ | new_n1154_;
  assign new_n1157_ = new_n1639_ | new_n1598_;
  assign new_n1158_ = new_n1635_ | new_n1593_;
  assign new_n1159_ = new_n1158_ & new_n1157_;
  assign new_n1160_ = new_n1662_ & new_n1663_;
  assign new_n1161_ = new_n1662_ | new_n1663_;
  assign new_n1162_ = new_n1664_ & new_n1572_;
  assign new_n1163_ = new_n802_ | new_n1576_;
  assign new_n1164_ = new_n1665_ & new_n1667_;
  assign new_n1165_ = new_n1668_ | new_n1669_;
  assign new_n1166_ = new_n1668_ & new_n1669_;
  assign new_n1167_ = new_n1665_ | new_n1667_;
  assign new_n1168_ = new_n1167_ & new_n1165_;
  assign new_n1169_ = new_n1166_ | new_n1164_;
  assign new_n1170_ = new_n1670_ & new_n1671_;
  assign new_n1171_ = new_n1672_ | new_n1673_;
  assign new_n1172_ = new_n1672_ & new_n1673_;
  assign new_n1173_ = new_n1670_ | new_n1671_;
  assign new_n1174_ = new_n1173_ & new_n1171_;
  assign new_n1175_ = new_n1172_ | new_n1170_;
  assign new_n1176_ = new_n1174_ & new_n1083_;
  assign new_n1177_ = new_n1175_ & new_n1674_;
  assign new_n1178_ = new_n1177_ | new_n1176_;
  assign new_n1179_ = new_n1676_ & new_n1679_;
  assign new_n1180_ = new_n1682_ | new_n1685_;
  assign new_n1181_ = new_n1682_ & new_n1685_;
  assign new_n1182_ = new_n1676_ | new_n1679_;
  assign new_n1183_ = new_n1182_ & new_n1180_;
  assign new_n1184_ = new_n1181_ | new_n1179_;
  assign new_n1185_ = new_n1687_ & new_n1689_;
  assign new_n1186_ = new_n1690_ & new_n1691_;
  assign new_n1187_ = new_n1186_ | new_n1185_;
  assign new_n1188_ = new_n1692_ & new_n1693_;
  assign new_n1189_ = new_n1695_ & new_n1697_;
  assign new_n1190_ = new_n1699_ & new_n1701_;
  assign new_n1191_ = new_n552_ & new_n1702_;
  assign new_n1192_ = new_n1191_ & new_n1703_;
  assign new_n1193_ = new_n1692_ & new_n1704_;
  assign new_n1194_ = new_n1705_ | new_n858_;
  assign new_n1195_ = new_n1193_ & new_n1703_;
  assign new_n1196_ = new_n1194_ | new_n1706_;
  assign new_n1197_ = new_n1196_ & new_n1683_;
  assign new_n1198_ = new_n1195_ & new_n1675_;
  assign new_n1199_ = new_n1198_ | new_n1197_;
  assign new_n1200_ = new_n1707_ & new_n1709_;
  assign new_n1201_ = new_n1707_ | new_n1709_;
  assign new_n1202_ = new_n1687_ & new_n1711_;
  assign new_n1203_ = new_n1690_ & new_n1713_;
  assign new_n1204_ = new_n1203_ | new_n1202_;
  assign new_n1205_ = new_n1695_ & new_n1717_;
  assign new_n1206_ = new_n1699_ | new_n1720_;
  assign new_n1207_ = new_n1700_ & new_n1720_;
  assign new_n1208_ = new_n1694_ | new_n1717_;
  assign new_n1209_ = new_n1208_ & new_n1206_;
  assign new_n1210_ = new_n1207_ | new_n1205_;
  assign new_n1211_ = new_n1210_ & new_n1723_;
  assign new_n1212_ = new_n1209_ & new_n1725_;
  assign new_n1213_ = new_n1212_ | new_n1211_;
  assign new_n1214_ = new_n1136_ & new_n1689_;
  assign new_n1215_ = new_n1727_ & new_n1691_;
  assign new_n1216_ = new_n1215_ | new_n1214_;
  assign new_n1217_ = new_n1723_ & new_n1728_;
  assign new_n1218_ = new_n1725_ | new_n1730_;
  assign new_n1219_ = new_n1726_ & new_n1730_;
  assign new_n1220_ = new_n1722_ | new_n1728_;
  assign new_n1221_ = new_n1220_ & new_n1218_;
  assign new_n1222_ = new_n1219_ | new_n1217_;
  assign new_n1223_ = new_n1222_ & new_n1731_;
  assign new_n1224_ = new_n1221_ & new_n494_;
  assign new_n1225_ = new_n1224_ | new_n1223_;
  assign new_n1226_ = new_n1686_ & new_n1734_;
  assign new_n1227_ = new_n1678_ | new_n1737_;
  assign new_n1228_ = new_n1680_ & new_n1737_;
  assign new_n1229_ = new_n1686_ | new_n1734_;
  assign new_n1230_ = new_n1229_ & new_n1227_;
  assign new_n1231_ = new_n1228_ | new_n1226_;
  assign new_n1232_ = new_n1231_ & new_n502_;
  assign new_n1233_ = new_n1230_ & new_n1739_;
  assign new_n1234_ = new_n1233_ | new_n1232_;
  assign new_n1235_ = new_n1738_ & new_n1721_;
  assign new_n1236_ = new_n1733_ | new_n1716_;
  assign new_n1237_ = new_n1735_ & new_n1718_;
  assign new_n1238_ = new_n1738_ | new_n1721_;
  assign new_n1239_ = new_n1238_ & new_n1236_;
  assign new_n1240_ = new_n1237_ | new_n1235_;
  assign new_n1241_ = new_n1240_ & new_n1697_;
  assign new_n1242_ = new_n1239_ & new_n1701_;
  assign new_n1243_ = new_n1242_ | new_n1241_;
  assign new_n1244_ = new_n1740_ & new_n1711_;
  assign new_n1245_ = new_n1742_ | new_n1713_;
  assign new_n1246_ = new_n1742_ & new_n1714_;
  assign new_n1247_ = new_n1740_ | new_n1710_;
  assign new_n1248_ = new_n1247_ & new_n1245_;
  assign new_n1249_ = new_n1246_ | new_n1244_;
  assign new_n1250_ = new_n1249_ & new_n1743_;
  assign new_n1251_ = new_n1248_ & new_n1708_;
  assign new_n1252_ = new_n1251_ | new_n1250_;
  assign new_n1253_ = new_n1744_ & new_n1746_;
  assign new_n1254_ = new_n1744_ | new_n1746_;
  assign G1884 = new_n865_;
  assign G1885 = new_n868_;
  assign G1886 = new_n871_;
  assign G1887 = new_n874_;
  assign G1888 = new_n879_;
  assign G1889 = new_n882_;
  assign G1890 = new_n885_;
  assign G1891 = new_n894_;
  assign G1892 = new_n897_;
  assign G1893 = new_n900_;
  assign G1894 = new_n903_;
  assign G1895 = new_n908_;
  assign G1896 = new_n919_;
  assign G1897 = new_n922_;
  assign G1898 = new_n925_;
  assign G1899 = new_n928_;
  assign G1900 = new_n937_;
  assign G1901 = new_n945_;
  assign G1902 = new_n953_;
  assign G1903 = new_n957_;
  assign G1904 = new_n961_;
  assign G1905 = new_n965_;
  assign G1906 = new_n980_;
  assign G1907 = new_n997_;
  assign G1908 = new_n1001_;
  assign n2248_li000_li000 = new_n427_;
  assign n2257_li003_li003 = new_n661_;
  assign n2269_li007_li007 = new_n641_;
  assign n2281_li011_li011 = new_n643_;
  assign n2284_li012_li012 = new_n433_;
  assign n2293_li015_li015 = new_n663_;
  assign n2296_li016_li016 = new_n435_;
  assign n2305_li019_li019 = new_n665_;
  assign n2317_li023_li023 = new_n645_;
  assign n2329_li027_li027 = new_n647_;
  assign n2341_li031_li031 = new_n649_;
  assign n2353_li035_li035 = new_n651_;
  assign n2365_li039_li039 = new_n625_;
  assign n2368_li040_li040 = new_n447_;
  assign n2377_li043_li043 = new_n657_;
  assign n2389_li047_li047 = new_n627_;
  assign n2401_li051_li051 = new_n629_;
  assign n2413_li055_li055 = new_n653_;
  assign n2425_li059_li059 = new_n631_;
  assign n2428_li060_li060 = new_n457_;
  assign n2437_li063_li063 = new_n659_;
  assign n2440_li064_li064 = new_n459_;
  assign n2464_li072_li072 = new_n463_;
  assign n2476_li076_li076 = new_n465_;
  assign n2488_li080_li080 = new_n467_;
  assign n2497_li083_li083 = new_n681_;
  assign n2500_li084_li084 = new_n469_;
  assign n2503_li085_li085 = new_n545_;
  assign n2509_li087_li087 = new_n695_;
  assign n2512_li088_li088 = new_n471_;
  assign n2536_li096_li096 = new_n475_;
  assign n2539_li097_li097 = new_n553_;
  assign n2542_li098_li098 = new_n555_;
  assign n2545_li099_li099 = new_n1552_;
  assign n2548_li100_li100 = new_n477_;
  assign n2551_li101_li101 = new_n561_;
  assign n2557_li103_li103 = new_n1554_;
  assign n2560_li104_li104 = new_n479_;
  assign n2563_li105_li105 = new_n567_;
  assign n2569_li107_li107 = new_n1553_;
  assign n2572_li108_li108 = new_n481_;
  assign n2575_li109_li109 = new_n573_;
  assign n2581_li111_li111 = new_n743_;
  assign n2584_li112_li112 = new_n483_;
  assign n2587_li113_li113 = new_n579_;
  assign n2590_li114_li114 = new_n581_;
  assign n2593_li115_li115 = new_n1548_;
  assign n2596_li116_li116 = new_n485_;
  assign n2599_li117_li117 = new_n587_;
  assign n2602_li118_li118 = new_n589_;
  assign n2605_li119_li119 = new_n1549_;
  assign n2608_li120_li120 = new_n487_;
  assign n2611_li121_li121 = new_n595_;
  assign n2617_li123_li123 = new_n1543_;
  assign n2620_li124_li124 = new_n489_;
  assign n2623_li125_li125 = new_n601_;
  assign n2626_li126_li126 = new_n603_;
  assign n2629_li127_li127 = new_n1550_;
  assign n2641_li131_li131 = new_n1547_;
  assign n1225_i2 = new_n733_;
  assign n1229_i2 = new_n737_;
  assign n1228_i2 = new_n735_;
  assign n1259_i2 = new_n749_;
  assign n1272_i2 = new_n759_;
  assign n1269_i2 = new_n757_;
  assign n1307_i2 = new_n1540_;
  assign n1201_i2 = new_n703_;
  assign n1202_i2 = new_n705_;
  assign n1203_i2 = new_n1588_;
  assign n1204_i2 = new_n709_;
  assign n622_i2 = new_n1544_;
  assign n1205_i2 = new_n711_;
  assign n1206_i2 = new_n1646_;
  assign n497_i2 = new_n1551_;
  assign n1212_i2 = new_n1628_;
  assign n1213_i2 = new_n719_;
  assign n1214_i2 = new_n721_;
  assign n1215_i2 = new_n723_;
  assign n1216_i2 = new_n1608_;
  assign n1217_i2 = new_n1666_;
  assign n1218_i2 = new_n1660_;
  assign n1219_i2 = new_n1576_;
  assign n1242_i2 = new_n739_;
  assign n1243_i2 = new_n741_;
  assign n1273_i2 = new_n1631_;
  assign n1274_i2 = new_n1603_;
  assign n1275_i2 = new_n765_;
  assign n1276_i2 = new_n767_;
  assign n1277_i2 = new_n1560_;
  assign n1286_i2 = new_n771_;
  assign n1299_i2 = new_n783_;
  assign n601_i2 = ~new_n1558_;
  assign n625_i2 = new_n1557_;
  assign n463_i2 = ~new_n1556_;
  assign lo082_buf_i2 = new_n1664_;
  assign n455_i2 = new_n1617_;
  assign n642_i2 = new_n1620_;
  assign n459_i2 = new_n1618_;
  assign n501_i2 = ~new_n1555_;
  assign n599_i2 = new_n1559_;
  assign n485_i2 = new_n1639_;
  assign lo086_buf_i2 = new_n1658_;
  assign lo122_buf_i2 = new_n1564_;
  assign n502_i2 = ~new_n1622_;
  assign n627_i2 = new_n1621_;
  assign lo038_buf_i2 = new_n1680_;
  assign lo046_buf_i2 = new_n1714_;
  assign lo050_buf_i2 = new_n1741_;
  assign lo058_buf_i2 = new_n1683_;
  assign lo070_buf_i2 = new_n1704_;
  assign lo094_buf_i2 = new_n1705_;
  assign n462_i2 = new_n1614_;
  assign lo006_buf_i2 = new_n1729_;
  assign lo010_buf_i2 = new_n1726_;
  assign lo022_buf_i2 = new_n1718_;
  assign lo026_buf_i2 = new_n1735_;
  assign lo030_buf_i2 = new_n1700_;
  assign lo034_buf_i2 = new_n1644_;
  assign lo054_buf_i2 = new_n1642_;
  assign lo130_buf_i2 = new_n1706_;
  assign n547_i2 = new_n1651_;
  assign n568_i2 = new_n1654_;
  assign n617_i2 = new_n1674_;
  assign lo042_buf_i2 = new_n1743_;
  assign lo062_buf_i2 = new_n1688_;
  assign lo110_buf_i2 = new_n575_;
  assign n733_i2 = new_n1084_;
  assign n734_i2 = new_n1085_;
  assign n570_i2 = new_n1656_;
  assign n461_i2 = new_n1091_;
  assign n644_i2 = new_n1093_;
  assign n628_i2 = new_n1094_;
  assign n528_i2 = new_n1647_;
  assign n592_i2 = ~new_n1650_;
  assign lo002_buf_i2 = new_n1731_;
  assign lo014_buf_i2 = new_n1739_;
  assign lo018_buf_i2 = new_n1696_;
  assign lo078_buf_i2 = new_n1702_;
  assign lo090_buf_i2 = new_n551_;
  assign n513_i2 = new_n1727_;
  assign lo102_buf_i2 = new_n563_;
  assign lo106_buf_i2 = new_n569_;
  assign n600_i2 = new_n1137_;
  assign n529_i2 = new_n1138_;
  assign n593_i2 = ~new_n1139_;
  assign lo066_buf_i2 = new_n1693_;
  assign n549_i2 = new_n1141_;
  assign n550_i2 = ~new_n1142_;
  assign n571_i2 = new_n1144_;
  assign n572_i2 = new_n1145_;
  assign n495_i2 = new_n1160_;
  assign n496_i2 = ~new_n1161_;
  assign n620_i2 = new_n1178_;
  assign n482_i2 = ~new_n1745_;
  assign lo081_buf_i2 = new_n541_;
  assign n576_i2 = new_n1188_;
  assign n520_i2 = new_n1189_;
  assign n521_i2 = new_n1190_;
  assign n562_i2 = new_n1192_;
  assign n508_i2 = new_n1200_;
  assign n509_i2 = ~new_n1201_;
  assign lo074_buf_i2 = new_n537_;
  assign n539_i2 = new_n1204_;
  assign n536_i2 = new_n1213_;
  assign n516_i2 = new_n1216_;
  assign n491_i2 = new_n1225_;
  assign n557_i2 = new_n1234_;
  assign n586_i2 = new_n1243_;
  assign n483_i2 = new_n1253_;
  assign n484_i2 = ~new_n1254_;
  assign lo004_buf_i2 = new_n429_;
  assign lo008_buf_i2 = new_n431_;
  assign lo020_buf_i2 = new_n437_;
  assign lo024_buf_i2 = new_n439_;
  assign lo028_buf_i2 = new_n441_;
  assign lo032_buf_i2 = new_n443_;
  assign lo052_buf_i2 = new_n453_;
  assign lo128_buf_i2 = new_n491_;
  assign lo037_buf_i2 = new_n445_;
  assign lo045_buf_i2 = new_n449_;
  assign lo049_buf_i2 = new_n451_;
  assign lo057_buf_i2 = new_n455_;
  assign lo069_buf_i2 = new_n461_;
  assign lo093_buf_i2 = new_n473_;
  assign new_n1464_ = new_n755_;
  assign new_n1465_ = new_n752_;
  assign new_n1466_ = new_n756_;
  assign new_n1467_ = new_n751_;
  assign new_n1468_ = new_n862_;
  assign new_n1469_ = new_n1468_;
  assign new_n1470_ = new_n1469_;
  assign new_n1471_ = new_n1469_;
  assign new_n1472_ = new_n1468_;
  assign new_n1473_ = new_n1472_;
  assign new_n1474_ = new_n861_;
  assign new_n1475_ = new_n1474_;
  assign new_n1476_ = new_n1475_;
  assign new_n1477_ = new_n1475_;
  assign new_n1478_ = new_n1474_;
  assign new_n1479_ = new_n1478_;
  assign new_n1480_ = new_n754_;
  assign new_n1481_ = new_n1480_;
  assign new_n1482_ = new_n753_;
  assign new_n1483_ = new_n1482_;
  assign new_n1484_ = new_n876_;
  assign new_n1485_ = new_n1484_;
  assign new_n1486_ = new_n1485_;
  assign new_n1487_ = new_n1485_;
  assign new_n1488_ = new_n1484_;
  assign new_n1489_ = new_n875_;
  assign new_n1490_ = new_n1489_;
  assign new_n1491_ = new_n1490_;
  assign new_n1492_ = new_n1490_;
  assign new_n1493_ = new_n1489_;
  assign new_n1494_ = new_n690_;
  assign new_n1495_ = new_n680_;
  assign new_n1496_ = new_n888_;
  assign new_n1497_ = new_n889_;
  assign new_n1498_ = new_n891_;
  assign new_n1499_ = new_n1498_;
  assign new_n1500_ = new_n1498_;
  assign new_n1501_ = new_n890_;
  assign new_n1502_ = new_n1501_;
  assign new_n1503_ = new_n1501_;
  assign new_n1504_ = new_n676_;
  assign new_n1505_ = new_n677_;
  assign new_n1506_ = new_n691_;
  assign new_n1507_ = new_n916_;
  assign new_n1508_ = new_n1507_;
  assign new_n1509_ = new_n1507_;
  assign new_n1510_ = new_n915_;
  assign new_n1511_ = new_n1510_;
  assign new_n1512_ = new_n1510_;
  assign new_n1513_ = new_n930_;
  assign new_n1514_ = new_n1513_;
  assign new_n1515_ = new_n1514_;
  assign new_n1516_ = new_n1514_;
  assign new_n1517_ = new_n1513_;
  assign new_n1518_ = new_n609_;
  assign new_n1519_ = new_n1518_;
  assign new_n1520_ = new_n600_;
  assign new_n1521_ = new_n1520_;
  assign new_n1522_ = new_n1521_;
  assign new_n1523_ = new_n1520_;
  assign new_n1524_ = new_n599_;
  assign new_n1525_ = new_n1524_;
  assign new_n1526_ = new_n929_;
  assign new_n1527_ = new_n1526_;
  assign new_n1528_ = new_n687_;
  assign new_n1529_ = new_n1528_;
  assign new_n1530_ = new_n1529_;
  assign new_n1531_ = new_n1529_;
  assign new_n1532_ = new_n1528_;
  assign new_n1533_ = new_n610_;
  assign new_n1534_ = new_n971_;
  assign new_n1535_ = new_n970_;
  assign new_n1536_ = new_n988_;
  assign new_n1537_ = new_n987_;
  assign new_n1538_ = new_n778_;
  assign new_n1539_ = new_n698_;
  assign new_n1540_ = new_n797_;
  assign new_n1541_ = new_n697_;
  assign new_n1542_ = new_n1541_;
  assign new_n1543_ = new_n1541_;
  assign new_n1544_ = new_n1002_;
  assign new_n1545_ = new_n655_;
  assign new_n1546_ = new_n1545_;
  assign new_n1547_ = new_n1545_;
  assign new_n1548_ = new_n583_;
  assign new_n1549_ = new_n591_;
  assign new_n1550_ = new_n605_;
  assign new_n1551_ = new_n1005_;
  assign new_n1552_ = new_n557_;
  assign new_n1553_ = new_n775_;
  assign new_n1554_ = new_n773_;
  assign new_n1555_ = new_n1020_;
  assign new_n1556_ = new_n1012_;
  assign new_n1557_ = new_n1011_;
  assign new_n1558_ = new_n1006_;
  assign new_n1559_ = new_n1031_;
  assign new_n1560_ = new_n769_;
  assign new_n1561_ = new_n1560_;
  assign new_n1562_ = new_n597_;
  assign new_n1563_ = new_n1562_;
  assign new_n1564_ = new_n1562_;
  assign new_n1565_ = new_n819_;
  assign new_n1566_ = new_n818_;
  assign new_n1567_ = new_n820_;
  assign new_n1568_ = new_n817_;
  assign new_n1569_ = new_n815_;
  assign new_n1570_ = new_n732_;
  assign new_n1571_ = new_n1570_;
  assign new_n1572_ = new_n1570_;
  assign new_n1573_ = new_n731_;
  assign new_n1574_ = new_n1573_;
  assign new_n1575_ = new_n1574_;
  assign new_n1576_ = new_n1573_;
  assign new_n1577_ = new_n825_;
  assign new_n1578_ = new_n822_;
  assign new_n1579_ = new_n1578_;
  assign new_n1580_ = new_n1578_;
  assign new_n1581_ = new_n826_;
  assign new_n1582_ = new_n821_;
  assign new_n1583_ = new_n1582_;
  assign new_n1584_ = new_n1582_;
  assign new_n1585_ = new_n809_;
  assign new_n1586_ = new_n708_;
  assign new_n1587_ = new_n810_;
  assign new_n1588_ = new_n707_;
  assign new_n1589_ = new_n1588_;
  assign new_n1590_ = new_n827_;
  assign new_n1591_ = new_n1590_;
  assign new_n1592_ = new_n1590_;
  assign new_n1593_ = new_n823_;
  assign new_n1594_ = new_n1593_;
  assign new_n1595_ = new_n828_;
  assign new_n1596_ = new_n1595_;
  assign new_n1597_ = new_n1595_;
  assign new_n1598_ = new_n824_;
  assign new_n1599_ = new_n1598_;
  assign new_n1600_ = new_n763_;
  assign new_n1601_ = new_n1600_;
  assign new_n1602_ = new_n1601_;
  assign new_n1603_ = new_n1600_;
  assign new_n1604_ = new_n726_;
  assign new_n1605_ = new_n764_;
  assign new_n1606_ = new_n1605_;
  assign new_n1607_ = new_n1605_;
  assign new_n1608_ = new_n725_;
  assign new_n1609_ = new_n1608_;
  assign new_n1610_ = new_n1076_;
  assign new_n1611_ = new_n1071_;
  assign new_n1612_ = new_n1077_;
  assign new_n1613_ = new_n1070_;
  assign new_n1614_ = new_n1037_;
  assign new_n1615_ = new_n1087_;
  assign new_n1616_ = new_n1088_;
  assign new_n1617_ = new_n1013_;
  assign new_n1618_ = new_n1015_;
  assign new_n1619_ = new_n1090_;
  assign new_n1620_ = new_n1014_;
  assign new_n1621_ = new_n1036_;
  assign new_n1622_ = new_n1034_;
  assign new_n1623_ = new_n1095_;
  assign new_n1624_ = new_n1096_;
  assign new_n1625_ = new_n1104_;
  assign new_n1626_ = new_n718_;
  assign new_n1627_ = new_n1103_;
  assign new_n1628_ = new_n717_;
  assign new_n1629_ = new_n1628_;
  assign new_n1630_ = new_n1114_;
  assign new_n1631_ = new_n761_;
  assign new_n1632_ = new_n1631_;
  assign new_n1633_ = new_n1115_;
  assign new_n1634_ = new_n762_;
  assign new_n1635_ = new_n1032_;
  assign new_n1636_ = new_n1635_;
  assign new_n1637_ = new_n1033_;
  assign new_n1638_ = new_n1637_;
  assign new_n1639_ = new_n1637_;
  assign new_n1640_ = new_n846_;
  assign new_n1641_ = new_n844_;
  assign new_n1642_ = new_n845_;
  assign new_n1643_ = new_n1642_;
  assign new_n1644_ = new_n843_;
  assign new_n1645_ = new_n1644_;
  assign new_n1646_ = new_n713_;
  assign new_n1647_ = new_n1113_;
  assign new_n1648_ = new_n598_;
  assign new_n1649_ = new_n1648_;
  assign new_n1650_ = new_n1130_;
  assign new_n1651_ = new_n1050_;
  assign new_n1652_ = new_n1140_;
  assign new_n1653_ = new_n576_;
  assign new_n1654_ = new_n1065_;
  assign new_n1655_ = new_n1143_;
  assign new_n1656_ = new_n1086_;
  assign new_n1657_ = new_n1656_;
  assign new_n1658_ = new_n547_;
  assign new_n1659_ = new_n730_;
  assign new_n1660_ = new_n729_;
  assign new_n1661_ = new_n1660_;
  assign new_n1662_ = new_n1159_;
  assign new_n1663_ = new_n1156_;
  assign new_n1664_ = new_n801_;
  assign new_n1665_ = new_n800_;
  assign new_n1666_ = new_n727_;
  assign new_n1667_ = new_n1666_;
  assign new_n1668_ = new_n799_;
  assign new_n1669_ = new_n728_;
  assign new_n1670_ = new_n1169_;
  assign new_n1671_ = new_n1162_;
  assign new_n1672_ = new_n1168_;
  assign new_n1673_ = new_n1163_;
  assign new_n1674_ = new_n1082_;
  assign new_n1675_ = new_n856_;
  assign new_n1676_ = new_n1675_;
  assign new_n1677_ = new_n849_;
  assign new_n1678_ = new_n1677_;
  assign new_n1679_ = new_n1678_;
  assign new_n1680_ = new_n1677_;
  assign new_n1681_ = new_n855_;
  assign new_n1682_ = new_n1681_;
  assign new_n1683_ = new_n1681_;
  assign new_n1684_ = new_n850_;
  assign new_n1685_ = new_n1684_;
  assign new_n1686_ = new_n1684_;
  assign new_n1687_ = new_n1184_;
  assign new_n1688_ = new_n531_;
  assign new_n1689_ = new_n1688_;
  assign new_n1690_ = new_n1183_;
  assign new_n1691_ = new_n532_;
  assign new_n1692_ = new_n860_;
  assign new_n1693_ = new_n535_;
  assign new_n1694_ = new_n842_;
  assign new_n1695_ = new_n1694_;
  assign new_n1696_ = new_n505_;
  assign new_n1697_ = new_n1696_;
  assign new_n1698_ = new_n841_;
  assign new_n1699_ = new_n1698_;
  assign new_n1700_ = new_n1698_;
  assign new_n1701_ = new_n506_;
  assign new_n1702_ = new_n539_;
  assign new_n1703_ = new_n848_;
  assign new_n1704_ = new_n857_;
  assign new_n1705_ = new_n859_;
  assign new_n1706_ = new_n847_;
  assign new_n1707_ = new_n1199_;
  assign new_n1708_ = new_n520_;
  assign new_n1709_ = new_n1708_;
  assign new_n1710_ = new_n852_;
  assign new_n1711_ = new_n1710_;
  assign new_n1712_ = new_n851_;
  assign new_n1713_ = new_n1712_;
  assign new_n1714_ = new_n1712_;
  assign new_n1715_ = new_n837_;
  assign new_n1716_ = new_n1715_;
  assign new_n1717_ = new_n1716_;
  assign new_n1718_ = new_n1715_;
  assign new_n1719_ = new_n838_;
  assign new_n1720_ = new_n1719_;
  assign new_n1721_ = new_n1719_;
  assign new_n1722_ = new_n836_;
  assign new_n1723_ = new_n1722_;
  assign new_n1724_ = new_n835_;
  assign new_n1725_ = new_n1724_;
  assign new_n1726_ = new_n1724_;
  assign new_n1727_ = new_n1135_;
  assign new_n1728_ = new_n834_;
  assign new_n1729_ = new_n833_;
  assign new_n1730_ = new_n1729_;
  assign new_n1731_ = new_n493_;
  assign new_n1732_ = new_n839_;
  assign new_n1733_ = new_n1732_;
  assign new_n1734_ = new_n1733_;
  assign new_n1735_ = new_n1732_;
  assign new_n1736_ = new_n840_;
  assign new_n1737_ = new_n1736_;
  assign new_n1738_ = new_n1736_;
  assign new_n1739_ = new_n501_;
  assign new_n1740_ = new_n854_;
  assign new_n1741_ = new_n853_;
  assign new_n1742_ = new_n1741_;
  assign new_n1743_ = new_n519_;
  assign new_n1744_ = new_n1252_;
  assign new_n1745_ = new_n1187_;
  assign new_n1746_ = new_n1745_;
  always @ (posedge clock) begin
    n940_lo <= n2248_li000_li000;
    n949_lo <= n2257_li003_li003;
    n961_lo <= n2269_li007_li007;
    n973_lo <= n2281_li011_li011;
    n976_lo <= n2284_li012_li012;
    n985_lo <= n2293_li015_li015;
    n988_lo <= n2296_li016_li016;
    n997_lo <= n2305_li019_li019;
    n1009_lo <= n2317_li023_li023;
    n1021_lo <= n2329_li027_li027;
    n1033_lo <= n2341_li031_li031;
    n1045_lo <= n2353_li035_li035;
    n1057_lo <= n2365_li039_li039;
    n1060_lo <= n2368_li040_li040;
    n1069_lo <= n2377_li043_li043;
    n1081_lo <= n2389_li047_li047;
    n1093_lo <= n2401_li051_li051;
    n1105_lo <= n2413_li055_li055;
    n1117_lo <= n2425_li059_li059;
    n1120_lo <= n2428_li060_li060;
    n1129_lo <= n2437_li063_li063;
    n1132_lo <= n2440_li064_li064;
    n1156_lo <= n2464_li072_li072;
    n1168_lo <= n2476_li076_li076;
    n1180_lo <= n2488_li080_li080;
    n1189_lo <= n2497_li083_li083;
    n1192_lo <= n2500_li084_li084;
    n1195_lo <= n2503_li085_li085;
    n1201_lo <= n2509_li087_li087;
    n1204_lo <= n2512_li088_li088;
    n1228_lo <= n2536_li096_li096;
    n1231_lo <= n2539_li097_li097;
    n1234_lo <= n2542_li098_li098;
    n1237_lo <= n2545_li099_li099;
    n1240_lo <= n2548_li100_li100;
    n1243_lo <= n2551_li101_li101;
    n1249_lo <= n2557_li103_li103;
    n1252_lo <= n2560_li104_li104;
    n1255_lo <= n2563_li105_li105;
    n1261_lo <= n2569_li107_li107;
    n1264_lo <= n2572_li108_li108;
    n1267_lo <= n2575_li109_li109;
    n1273_lo <= n2581_li111_li111;
    n1276_lo <= n2584_li112_li112;
    n1279_lo <= n2587_li113_li113;
    n1282_lo <= n2590_li114_li114;
    n1285_lo <= n2593_li115_li115;
    n1288_lo <= n2596_li116_li116;
    n1291_lo <= n2599_li117_li117;
    n1294_lo <= n2602_li118_li118;
    n1297_lo <= n2605_li119_li119;
    n1300_lo <= n2608_li120_li120;
    n1303_lo <= n2611_li121_li121;
    n1309_lo <= n2617_li123_li123;
    n1312_lo <= n2620_li124_li124;
    n1315_lo <= n2623_li125_li125;
    n1318_lo <= n2626_li126_li126;
    n1321_lo <= n2629_li127_li127;
    n1333_lo <= n2641_li131_li131;
    n1225_o2 <= n1225_i2;
    n1229_o2 <= n1229_i2;
    n1228_o2 <= n1228_i2;
    n1259_o2 <= n1259_i2;
    n1272_o2 <= n1272_i2;
    n1269_o2 <= n1269_i2;
    n1307_o2 <= n1307_i2;
    n1201_o2 <= n1201_i2;
    n1202_o2 <= n1202_i2;
    n1203_o2 <= n1203_i2;
    n1204_o2 <= n1204_i2;
    n622_o2 <= n622_i2;
    n1205_o2 <= n1205_i2;
    n1206_o2 <= n1206_i2;
    n497_o2 <= n497_i2;
    n1212_o2 <= n1212_i2;
    n1213_o2 <= n1213_i2;
    n1214_o2 <= n1214_i2;
    n1215_o2 <= n1215_i2;
    n1216_o2 <= n1216_i2;
    n1217_o2 <= n1217_i2;
    n1218_o2 <= n1218_i2;
    n1219_o2 <= n1219_i2;
    n1242_o2 <= n1242_i2;
    n1243_o2 <= n1243_i2;
    n1273_o2 <= n1273_i2;
    n1274_o2 <= n1274_i2;
    n1275_o2 <= n1275_i2;
    n1276_o2 <= n1276_i2;
    n1277_o2 <= n1277_i2;
    n1286_o2 <= n1286_i2;
    n1299_o2 <= n1299_i2;
    n601_o2 <= n601_i2;
    n625_o2 <= n625_i2;
    n463_o2 <= n463_i2;
    lo082_buf_o2 <= lo082_buf_i2;
    n455_o2 <= n455_i2;
    n642_o2 <= n642_i2;
    n459_o2 <= n459_i2;
    n501_o2 <= n501_i2;
    n599_o2 <= n599_i2;
    n485_o2 <= n485_i2;
    lo086_buf_o2 <= lo086_buf_i2;
    lo122_buf_o2 <= lo122_buf_i2;
    n502_o2 <= n502_i2;
    n627_o2 <= n627_i2;
    lo038_buf_o2 <= lo038_buf_i2;
    lo046_buf_o2 <= lo046_buf_i2;
    lo050_buf_o2 <= lo050_buf_i2;
    lo058_buf_o2 <= lo058_buf_i2;
    lo070_buf_o2 <= lo070_buf_i2;
    lo094_buf_o2 <= lo094_buf_i2;
    n462_o2 <= n462_i2;
    lo006_buf_o2 <= lo006_buf_i2;
    lo010_buf_o2 <= lo010_buf_i2;
    lo022_buf_o2 <= lo022_buf_i2;
    lo026_buf_o2 <= lo026_buf_i2;
    lo030_buf_o2 <= lo030_buf_i2;
    lo034_buf_o2 <= lo034_buf_i2;
    lo054_buf_o2 <= lo054_buf_i2;
    lo130_buf_o2 <= lo130_buf_i2;
    n547_o2 <= n547_i2;
    n424_inv <= n568_i2;
    n617_o2 <= n617_i2;
    lo042_buf_o2 <= lo042_buf_i2;
    lo062_buf_o2 <= lo062_buf_i2;
    lo110_buf_o2 <= lo110_buf_i2;
    n733_o2 <= n733_i2;
    n734_o2 <= n734_i2;
    n570_o2 <= n570_i2;
    n461_o2 <= n461_i2;
    n644_o2 <= n644_i2;
    n628_o2 <= n628_i2;
    n528_o2 <= n528_i2;
    n460_inv <= n592_i2;
    lo002_buf_o2 <= lo002_buf_i2;
    lo014_buf_o2 <= lo014_buf_i2;
    lo018_buf_o2 <= lo018_buf_i2;
    lo078_buf_o2 <= lo078_buf_i2;
    lo090_buf_o2 <= lo090_buf_i2;
    n513_o2 <= n513_i2;
    lo102_buf_o2 <= lo102_buf_i2;
    lo106_buf_o2 <= lo106_buf_i2;
    n600_o2 <= n600_i2;
    n529_o2 <= n529_i2;
    n593_o2 <= n593_i2;
    lo066_buf_o2 <= lo066_buf_i2;
    n549_o2 <= n549_i2;
    n550_o2 <= n550_i2;
    n571_o2 <= n571_i2;
    n572_o2 <= n572_i2;
    n495_o2 <= n495_i2;
    n496_o2 <= n496_i2;
    n620_o2 <= n620_i2;
    n482_o2 <= n482_i2;
    lo081_buf_o2 <= lo081_buf_i2;
    n576_o2 <= n576_i2;
    n520_o2 <= n520_i2;
    n521_o2 <= n521_i2;
    n562_o2 <= n562_i2;
    n508_o2 <= n508_i2;
    n509_o2 <= n509_i2;
    lo074_buf_o2 <= lo074_buf_i2;
    n539_o2 <= n539_i2;
    n536_o2 <= n536_i2;
    n516_o2 <= n516_i2;
    n491_o2 <= n491_i2;
    n557_o2 <= n557_i2;
    n586_o2 <= n586_i2;
    n483_o2 <= n483_i2;
    n484_o2 <= n484_i2;
    lo004_buf_o2 <= lo004_buf_i2;
    lo008_buf_o2 <= lo008_buf_i2;
    lo020_buf_o2 <= lo020_buf_i2;
    lo024_buf_o2 <= lo024_buf_i2;
    lo028_buf_o2 <= lo028_buf_i2;
    lo032_buf_o2 <= lo032_buf_i2;
    lo052_buf_o2 <= lo052_buf_i2;
    lo128_buf_o2 <= lo128_buf_i2;
    lo037_buf_o2 <= lo037_buf_i2;
    lo045_buf_o2 <= lo045_buf_i2;
    lo049_buf_o2 <= lo049_buf_i2;
    lo057_buf_o2 <= lo057_buf_i2;
    lo069_buf_o2 <= lo069_buf_i2;
    lo093_buf_o2 <= lo093_buf_i2;
  end
  initial begin
    n940_lo <= 1'b0;
    n949_lo <= 1'b0;
    n961_lo <= 1'b0;
    n973_lo <= 1'b0;
    n976_lo <= 1'b0;
    n985_lo <= 1'b0;
    n988_lo <= 1'b0;
    n997_lo <= 1'b0;
    n1009_lo <= 1'b0;
    n1021_lo <= 1'b0;
    n1033_lo <= 1'b0;
    n1045_lo <= 1'b0;
    n1057_lo <= 1'b0;
    n1060_lo <= 1'b0;
    n1069_lo <= 1'b0;
    n1081_lo <= 1'b0;
    n1093_lo <= 1'b0;
    n1105_lo <= 1'b0;
    n1117_lo <= 1'b0;
    n1120_lo <= 1'b0;
    n1129_lo <= 1'b0;
    n1132_lo <= 1'b0;
    n1156_lo <= 1'b0;
    n1168_lo <= 1'b0;
    n1180_lo <= 1'b0;
    n1189_lo <= 1'b0;
    n1192_lo <= 1'b0;
    n1195_lo <= 1'b0;
    n1201_lo <= 1'b0;
    n1204_lo <= 1'b0;
    n1228_lo <= 1'b0;
    n1231_lo <= 1'b0;
    n1234_lo <= 1'b0;
    n1237_lo <= 1'b0;
    n1240_lo <= 1'b0;
    n1243_lo <= 1'b0;
    n1249_lo <= 1'b0;
    n1252_lo <= 1'b0;
    n1255_lo <= 1'b0;
    n1261_lo <= 1'b0;
    n1264_lo <= 1'b0;
    n1267_lo <= 1'b0;
    n1273_lo <= 1'b0;
    n1276_lo <= 1'b0;
    n1279_lo <= 1'b0;
    n1282_lo <= 1'b0;
    n1285_lo <= 1'b0;
    n1288_lo <= 1'b0;
    n1291_lo <= 1'b0;
    n1294_lo <= 1'b0;
    n1297_lo <= 1'b0;
    n1300_lo <= 1'b0;
    n1303_lo <= 1'b0;
    n1309_lo <= 1'b0;
    n1312_lo <= 1'b0;
    n1315_lo <= 1'b0;
    n1318_lo <= 1'b0;
    n1321_lo <= 1'b0;
    n1333_lo <= 1'b0;
    n1225_o2 <= 1'b0;
    n1229_o2 <= 1'b0;
    n1228_o2 <= 1'b0;
    n1259_o2 <= 1'b0;
    n1272_o2 <= 1'b0;
    n1269_o2 <= 1'b0;
    n1307_o2 <= 1'b0;
    n1201_o2 <= 1'b0;
    n1202_o2 <= 1'b0;
    n1203_o2 <= 1'b0;
    n1204_o2 <= 1'b0;
    n622_o2 <= 1'b0;
    n1205_o2 <= 1'b0;
    n1206_o2 <= 1'b0;
    n497_o2 <= 1'b0;
    n1212_o2 <= 1'b0;
    n1213_o2 <= 1'b0;
    n1214_o2 <= 1'b0;
    n1215_o2 <= 1'b0;
    n1216_o2 <= 1'b0;
    n1217_o2 <= 1'b0;
    n1218_o2 <= 1'b0;
    n1219_o2 <= 1'b0;
    n1242_o2 <= 1'b0;
    n1243_o2 <= 1'b0;
    n1273_o2 <= 1'b0;
    n1274_o2 <= 1'b0;
    n1275_o2 <= 1'b0;
    n1276_o2 <= 1'b0;
    n1277_o2 <= 1'b0;
    n1286_o2 <= 1'b0;
    n1299_o2 <= 1'b0;
    n601_o2 <= 1'b0;
    n625_o2 <= 1'b0;
    n463_o2 <= 1'b0;
    lo082_buf_o2 <= 1'b0;
    n455_o2 <= 1'b0;
    n642_o2 <= 1'b0;
    n459_o2 <= 1'b0;
    n501_o2 <= 1'b0;
    n599_o2 <= 1'b0;
    n485_o2 <= 1'b0;
    lo086_buf_o2 <= 1'b0;
    lo122_buf_o2 <= 1'b0;
    n502_o2 <= 1'b0;
    n627_o2 <= 1'b0;
    lo038_buf_o2 <= 1'b0;
    lo046_buf_o2 <= 1'b0;
    lo050_buf_o2 <= 1'b0;
    lo058_buf_o2 <= 1'b0;
    lo070_buf_o2 <= 1'b0;
    lo094_buf_o2 <= 1'b0;
    n462_o2 <= 1'b0;
    lo006_buf_o2 <= 1'b0;
    lo010_buf_o2 <= 1'b0;
    lo022_buf_o2 <= 1'b0;
    lo026_buf_o2 <= 1'b0;
    lo030_buf_o2 <= 1'b0;
    lo034_buf_o2 <= 1'b0;
    lo054_buf_o2 <= 1'b0;
    lo130_buf_o2 <= 1'b0;
    n547_o2 <= 1'b0;
    n424_inv <= 1'b0;
    n617_o2 <= 1'b0;
    lo042_buf_o2 <= 1'b0;
    lo062_buf_o2 <= 1'b0;
    lo110_buf_o2 <= 1'b0;
    n733_o2 <= 1'b0;
    n734_o2 <= 1'b0;
    n570_o2 <= 1'b0;
    n461_o2 <= 1'b0;
    n644_o2 <= 1'b0;
    n628_o2 <= 1'b0;
    n528_o2 <= 1'b0;
    n460_inv <= 1'b0;
    lo002_buf_o2 <= 1'b0;
    lo014_buf_o2 <= 1'b0;
    lo018_buf_o2 <= 1'b0;
    lo078_buf_o2 <= 1'b0;
    lo090_buf_o2 <= 1'b0;
    n513_o2 <= 1'b0;
    lo102_buf_o2 <= 1'b0;
    lo106_buf_o2 <= 1'b0;
    n600_o2 <= 1'b0;
    n529_o2 <= 1'b0;
    n593_o2 <= 1'b0;
    lo066_buf_o2 <= 1'b0;
    n549_o2 <= 1'b0;
    n550_o2 <= 1'b0;
    n571_o2 <= 1'b0;
    n572_o2 <= 1'b0;
    n495_o2 <= 1'b0;
    n496_o2 <= 1'b0;
    n620_o2 <= 1'b0;
    n482_o2 <= 1'b0;
    lo081_buf_o2 <= 1'b0;
    n576_o2 <= 1'b0;
    n520_o2 <= 1'b0;
    n521_o2 <= 1'b0;
    n562_o2 <= 1'b0;
    n508_o2 <= 1'b0;
    n509_o2 <= 1'b0;
    lo074_buf_o2 <= 1'b0;
    n539_o2 <= 1'b0;
    n536_o2 <= 1'b0;
    n516_o2 <= 1'b0;
    n491_o2 <= 1'b0;
    n557_o2 <= 1'b0;
    n586_o2 <= 1'b0;
    n483_o2 <= 1'b0;
    n484_o2 <= 1'b0;
    lo004_buf_o2 <= 1'b0;
    lo008_buf_o2 <= 1'b0;
    lo020_buf_o2 <= 1'b0;
    lo024_buf_o2 <= 1'b0;
    lo028_buf_o2 <= 1'b0;
    lo032_buf_o2 <= 1'b0;
    lo052_buf_o2 <= 1'b0;
    lo128_buf_o2 <= 1'b0;
    lo037_buf_o2 <= 1'b0;
    lo045_buf_o2 <= 1'b0;
    lo049_buf_o2 <= 1'b0;
    lo057_buf_o2 <= 1'b0;
    lo069_buf_o2 <= 1'b0;
    lo093_buf_o2 <= 1'b0;
  end
endmodule


