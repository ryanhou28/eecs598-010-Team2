
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  G42,
  G43,
  G44,
  G45,
  G46,
  G47,
  G48,
  G49,
  G50,
  G51,
  G52,
  G53,
  G54,
  G55,
  G56,
  G57,
  G58,
  G59,
  G60,
  n480_lo,
  n492_lo,
  n495_lo,
  n498_lo,
  n501_lo,
  n504_lo,
  n516_lo,
  n528_lo,
  n531_lo,
  n540_lo,
  n543_lo,
  n546_lo,
  n549_lo,
  n552_lo,
  n564_lo,
  n579_lo,
  n600_lo,
  n603_lo,
  n606_lo,
  n609_lo,
  n612_lo,
  n615_lo,
  n618_lo,
  n621_lo,
  n627_lo,
  n630_lo,
  n633_lo,
  n639_lo,
  n642_lo,
  n645_lo,
  n648_lo,
  n660_lo,
  n663_lo,
  n672_lo,
  n675_lo,
  n678_lo,
  n681_lo,
  n684_lo,
  n687_lo,
  n690_lo,
  n693_lo,
  n696_lo,
  n699_lo,
  n702_lo,
  n705_lo,
  n708_lo,
  n711_lo,
  n714_lo,
  n717_lo,
  n720_lo,
  n723_lo,
  n726_lo,
  n729_lo,
  n732_lo,
  n735_lo,
  n738_lo,
  n741_lo,
  n744_lo,
  n747_lo,
  n750_lo,
  n756_lo,
  n759_lo,
  n762_lo,
  n768_lo,
  n771_lo,
  n774_lo,
  n780_lo,
  n783_lo,
  n786_lo,
  n792_lo,
  n795_lo,
  n804_lo,
  n807_lo,
  n816_lo,
  n819_lo,
  n828_lo,
  n831_lo,
  n843_lo,
  n846_lo,
  n849_lo,
  n852_lo,
  n855_lo,
  n858_lo,
  n861_lo,
  n864_lo,
  n867_lo,
  n870_lo,
  n879_lo,
  n891_lo,
  n903_lo,
  n915_lo,
  n918_lo,
  n927_lo,
  n951_lo,
  n954_lo,
  n957_lo,
  n960_lo,
  n963_lo,
  n966_lo,
  n972_lo,
  n975_lo,
  n978_lo,
  n984_lo,
  n987_lo,
  n990_lo,
  n996_lo,
  n999_lo,
  n1002_lo,
  n1008_lo,
  n1011_lo,
  n1014_lo,
  n1020_lo,
  n1023_lo,
  n1026_lo,
  n1032_lo,
  n1035_lo,
  n1038_lo,
  n1044_lo,
  n1047_lo,
  n1050_lo,
  n1053_lo,
  n1056_lo,
  n1059_lo,
  n1062_lo,
  n1065_lo,
  n1068_lo,
  n1071_lo,
  n1074_lo,
  n1077_lo,
  n1080_lo,
  n1083_lo,
  n1086_lo,
  n1089_lo,
  n1092_lo,
  n1095_lo,
  n1098_lo,
  n1101_lo,
  n1104_lo,
  n1107_lo,
  n1110_lo,
  n1113_lo,
  n1116_lo,
  n1119_lo,
  n1122_lo,
  n1125_lo,
  n1128_lo,
  n1131_lo,
  n1134_lo,
  n1137_lo,
  n1140_lo,
  n1143_lo,
  n1146_lo,
  n1149_lo,
  n1152_lo,
  n1155_lo,
  n1158_lo,
  n1167_lo,
  n1170_lo,
  n1173_lo,
  n1176_lo,
  n1179_lo,
  n1529_o2,
  n1616_o2,
  n1655_o2,
  n1656_o2,
  n1657_o2,
  n1730_o2,
  n1731_o2,
  n1732_o2,
  n1729_o2,
  n1805_o2,
  n1808_o2,
  n1807_o2,
  n1809_o2,
  n1663_o2,
  n1664_o2,
  n1704_o2,
  n1705_o2,
  n1706_o2,
  n1707_o2,
  n1708_o2,
  n1709_o2,
  G280_o2,
  G655_o2,
  G663_o2,
  G672_o2,
  G538_o2,
  n1780_o2,
  n1781_o2,
  n1797_o2,
  n1798_o2,
  n1799_o2,
  n1800_o2,
  G578_o2,
  n1828_o2,
  n801_lo_buf_o2,
  G693_o2,
  G702_o2,
  G712_o2,
  G685_o2,
  G658_o2,
  G667_o2,
  G677_o2,
  G650_o2,
  G798_o2,
  n1017_lo_buf_o2,
  n1029_lo_buf_o2,
  n1041_lo_buf_o2,
  G558_o2,
  G562_o2,
  G566_o2,
  n1835_o2,
  n1836_o2,
  n1837_o2,
  n765_lo_buf_o2,
  n777_lo_buf_o2,
  n789_lo_buf_o2,
  G617_o2,
  G626_o2,
  G636_o2,
  n489_lo_buf_o2,
  n513_lo_buf_o2,
  n561_lo_buf_o2,
  n597_lo_buf_o2,
  n657_lo_buf_o2,
  G276_o2,
  n1005_lo_buf_o2,
  n1161_lo_buf_o2,
  G620_o2,
  G629_o2,
  G639_o2,
  G554_o2,
  G690_o2,
  G698_o2,
  G707_o2,
  G319_o2,
  G389_o2,
  n753_lo_buf_o2,
  G647_o2,
  G769_o2,
  G785_o2,
  G808_o2,
  G445_o2,
  G448_o2,
  G477_o2,
  G480_o2,
  G436_o2,
  G786_o2,
  G787_o2,
  G826_o2,
  G827_o2,
  G825_o2,
  G610_o2,
  n537_lo_buf_o2,
  n669_lo_buf_o2,
  n969_lo_buf_o2,
  n981_lo_buf_o2,
  n993_lo_buf_o2,
  G309_o2,
  G461_o2,
  G487_o2,
  G460_o2,
  G468_o2,
  G287_o2,
  G613_o2,
  n585_lo_buf_o2,
  n813_lo_buf_o2,
  n825_lo_buf_o2,
  n837_lo_buf_o2,
  n897_lo_buf_o2,
  n909_lo_buf_o2,
  n933_lo_buf_o2,
  G451_o2,
  G682_o2,
  G756_o2,
  G542_o2,
  G546_o2,
  G550_o2,
  G310_o2,
  n798_lo_buf_o2,
  n882_lo_buf_o2,
  G427_o2,
  G497_o2,
  G499_o2,
  G501_o2,
  G498_o2,
  G500_o2,
  G502_o2,
  G369_o2,
  n939_lo_buf_o2,
  n486_lo_buf_o2,
  n510_lo_buf_o2,
  n558_lo_buf_o2,
  n594_lo_buf_o2,
  n654_lo_buf_o2,
  n477_lo_buf_o2,
  n525_lo_buf_o2,
  n573_lo_buf_o2,
  G855,
  G856,
  G857,
  G858,
  G859,
  G860,
  G861,
  G862,
  G863,
  G864,
  G865,
  G866,
  G867,
  G868,
  G869,
  G870,
  G871,
  G872,
  G873,
  G874,
  G875,
  G876,
  G877,
  G878,
  G879,
  G880,
  n480_li,
  n492_li,
  n495_li,
  n498_li,
  n501_li,
  n504_li,
  n516_li,
  n528_li,
  n531_li,
  n540_li,
  n543_li,
  n546_li,
  n549_li,
  n552_li,
  n564_li,
  n579_li,
  n600_li,
  n603_li,
  n606_li,
  n609_li,
  n612_li,
  n615_li,
  n618_li,
  n621_li,
  n627_li,
  n630_li,
  n633_li,
  n639_li,
  n642_li,
  n645_li,
  n648_li,
  n660_li,
  n663_li,
  n672_li,
  n675_li,
  n678_li,
  n681_li,
  n684_li,
  n687_li,
  n690_li,
  n693_li,
  n696_li,
  n699_li,
  n702_li,
  n705_li,
  n708_li,
  n711_li,
  n714_li,
  n717_li,
  n720_li,
  n723_li,
  n726_li,
  n729_li,
  n732_li,
  n735_li,
  n738_li,
  n741_li,
  n744_li,
  n747_li,
  n750_li,
  n756_li,
  n759_li,
  n762_li,
  n768_li,
  n771_li,
  n774_li,
  n780_li,
  n783_li,
  n786_li,
  n792_li,
  n795_li,
  n804_li,
  n807_li,
  n816_li,
  n819_li,
  n828_li,
  n831_li,
  n843_li,
  n846_li,
  n849_li,
  n852_li,
  n855_li,
  n858_li,
  n861_li,
  n864_li,
  n867_li,
  n870_li,
  n879_li,
  n891_li,
  n903_li,
  n915_li,
  n918_li,
  n927_li,
  n951_li,
  n954_li,
  n957_li,
  n960_li,
  n963_li,
  n966_li,
  n972_li,
  n975_li,
  n978_li,
  n984_li,
  n987_li,
  n990_li,
  n996_li,
  n999_li,
  n1002_li,
  n1008_li,
  n1011_li,
  n1014_li,
  n1020_li,
  n1023_li,
  n1026_li,
  n1032_li,
  n1035_li,
  n1038_li,
  n1044_li,
  n1047_li,
  n1050_li,
  n1053_li,
  n1056_li,
  n1059_li,
  n1062_li,
  n1065_li,
  n1068_li,
  n1071_li,
  n1074_li,
  n1077_li,
  n1080_li,
  n1083_li,
  n1086_li,
  n1089_li,
  n1092_li,
  n1095_li,
  n1098_li,
  n1101_li,
  n1104_li,
  n1107_li,
  n1110_li,
  n1113_li,
  n1116_li,
  n1119_li,
  n1122_li,
  n1125_li,
  n1128_li,
  n1131_li,
  n1134_li,
  n1137_li,
  n1140_li,
  n1143_li,
  n1146_li,
  n1149_li,
  n1152_li,
  n1155_li,
  n1158_li,
  n1167_li,
  n1170_li,
  n1173_li,
  n1176_li,
  n1179_li,
  n1529_i2,
  n1616_i2,
  n1655_i2,
  n1656_i2,
  n1657_i2,
  n1730_i2,
  n1731_i2,
  n1732_i2,
  n1729_i2,
  n1805_i2,
  n1808_i2,
  n1807_i2,
  n1809_i2,
  n1663_i2,
  n1664_i2,
  n1704_i2,
  n1705_i2,
  n1706_i2,
  n1707_i2,
  n1708_i2,
  n1709_i2,
  G280_i2,
  G655_i2,
  G663_i2,
  G672_i2,
  G538_i2,
  n1780_i2,
  n1781_i2,
  n1797_i2,
  n1798_i2,
  n1799_i2,
  n1800_i2,
  G578_i2,
  n1828_i2,
  n801_lo_buf_i2,
  G693_i2,
  G702_i2,
  G712_i2,
  G685_i2,
  G658_i2,
  G667_i2,
  G677_i2,
  G650_i2,
  G798_i2,
  n1017_lo_buf_i2,
  n1029_lo_buf_i2,
  n1041_lo_buf_i2,
  G558_i2,
  G562_i2,
  G566_i2,
  n1835_i2,
  n1836_i2,
  n1837_i2,
  n765_lo_buf_i2,
  n777_lo_buf_i2,
  n789_lo_buf_i2,
  G617_i2,
  G626_i2,
  G636_i2,
  n489_lo_buf_i2,
  n513_lo_buf_i2,
  n561_lo_buf_i2,
  n597_lo_buf_i2,
  n657_lo_buf_i2,
  G276_i2,
  n1005_lo_buf_i2,
  n1161_lo_buf_i2,
  G620_i2,
  G629_i2,
  G639_i2,
  G554_i2,
  G690_i2,
  G698_i2,
  G707_i2,
  G319_i2,
  G389_i2,
  n753_lo_buf_i2,
  G647_i2,
  G769_i2,
  G785_i2,
  G808_i2,
  G445_i2,
  G448_i2,
  G477_i2,
  G480_i2,
  G436_i2,
  G786_i2,
  G787_i2,
  G826_i2,
  G827_i2,
  G825_i2,
  G610_i2,
  n537_lo_buf_i2,
  n669_lo_buf_i2,
  n969_lo_buf_i2,
  n981_lo_buf_i2,
  n993_lo_buf_i2,
  G309_i2,
  G461_i2,
  G487_i2,
  G460_i2,
  G468_i2,
  G287_i2,
  G613_i2,
  n585_lo_buf_i2,
  n813_lo_buf_i2,
  n825_lo_buf_i2,
  n837_lo_buf_i2,
  n897_lo_buf_i2,
  n909_lo_buf_i2,
  n933_lo_buf_i2,
  G451_i2,
  G682_i2,
  G756_i2,
  G542_i2,
  G546_i2,
  G550_i2,
  G310_i2,
  n798_lo_buf_i2,
  n882_lo_buf_i2,
  G427_i2,
  G497_i2,
  G499_i2,
  G501_i2,
  G498_i2,
  G500_i2,
  G502_i2,
  G369_i2,
  n939_lo_buf_i2,
  n486_lo_buf_i2,
  n510_lo_buf_i2,
  n558_lo_buf_i2,
  n594_lo_buf_i2,
  n654_lo_buf_i2,
  n477_lo_buf_i2,
  n525_lo_buf_i2,
  n573_lo_buf_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input G42;input G43;input G44;input G45;input G46;input G47;input G48;input G49;input G50;input G51;input G52;input G53;input G54;input G55;input G56;input G57;input G58;input G59;input G60;input n480_lo;input n492_lo;input n495_lo;input n498_lo;input n501_lo;input n504_lo;input n516_lo;input n528_lo;input n531_lo;input n540_lo;input n543_lo;input n546_lo;input n549_lo;input n552_lo;input n564_lo;input n579_lo;input n600_lo;input n603_lo;input n606_lo;input n609_lo;input n612_lo;input n615_lo;input n618_lo;input n621_lo;input n627_lo;input n630_lo;input n633_lo;input n639_lo;input n642_lo;input n645_lo;input n648_lo;input n660_lo;input n663_lo;input n672_lo;input n675_lo;input n678_lo;input n681_lo;input n684_lo;input n687_lo;input n690_lo;input n693_lo;input n696_lo;input n699_lo;input n702_lo;input n705_lo;input n708_lo;input n711_lo;input n714_lo;input n717_lo;input n720_lo;input n723_lo;input n726_lo;input n729_lo;input n732_lo;input n735_lo;input n738_lo;input n741_lo;input n744_lo;input n747_lo;input n750_lo;input n756_lo;input n759_lo;input n762_lo;input n768_lo;input n771_lo;input n774_lo;input n780_lo;input n783_lo;input n786_lo;input n792_lo;input n795_lo;input n804_lo;input n807_lo;input n816_lo;input n819_lo;input n828_lo;input n831_lo;input n843_lo;input n846_lo;input n849_lo;input n852_lo;input n855_lo;input n858_lo;input n861_lo;input n864_lo;input n867_lo;input n870_lo;input n879_lo;input n891_lo;input n903_lo;input n915_lo;input n918_lo;input n927_lo;input n951_lo;input n954_lo;input n957_lo;input n960_lo;input n963_lo;input n966_lo;input n972_lo;input n975_lo;input n978_lo;input n984_lo;input n987_lo;input n990_lo;input n996_lo;input n999_lo;input n1002_lo;input n1008_lo;input n1011_lo;input n1014_lo;input n1020_lo;input n1023_lo;input n1026_lo;input n1032_lo;input n1035_lo;input n1038_lo;input n1044_lo;input n1047_lo;input n1050_lo;input n1053_lo;input n1056_lo;input n1059_lo;input n1062_lo;input n1065_lo;input n1068_lo;input n1071_lo;input n1074_lo;input n1077_lo;input n1080_lo;input n1083_lo;input n1086_lo;input n1089_lo;input n1092_lo;input n1095_lo;input n1098_lo;input n1101_lo;input n1104_lo;input n1107_lo;input n1110_lo;input n1113_lo;input n1116_lo;input n1119_lo;input n1122_lo;input n1125_lo;input n1128_lo;input n1131_lo;input n1134_lo;input n1137_lo;input n1140_lo;input n1143_lo;input n1146_lo;input n1149_lo;input n1152_lo;input n1155_lo;input n1158_lo;input n1167_lo;input n1170_lo;input n1173_lo;input n1176_lo;input n1179_lo;input n1529_o2;input n1616_o2;input n1655_o2;input n1656_o2;input n1657_o2;input n1730_o2;input n1731_o2;input n1732_o2;input n1729_o2;input n1805_o2;input n1808_o2;input n1807_o2;input n1809_o2;input n1663_o2;input n1664_o2;input n1704_o2;input n1705_o2;input n1706_o2;input n1707_o2;input n1708_o2;input n1709_o2;input G280_o2;input G655_o2;input G663_o2;input G672_o2;input G538_o2;input n1780_o2;input n1781_o2;input n1797_o2;input n1798_o2;input n1799_o2;input n1800_o2;input G578_o2;input n1828_o2;input n801_lo_buf_o2;input G693_o2;input G702_o2;input G712_o2;input G685_o2;input G658_o2;input G667_o2;input G677_o2;input G650_o2;input G798_o2;input n1017_lo_buf_o2;input n1029_lo_buf_o2;input n1041_lo_buf_o2;input G558_o2;input G562_o2;input G566_o2;input n1835_o2;input n1836_o2;input n1837_o2;input n765_lo_buf_o2;input n777_lo_buf_o2;input n789_lo_buf_o2;input G617_o2;input G626_o2;input G636_o2;input n489_lo_buf_o2;input n513_lo_buf_o2;input n561_lo_buf_o2;input n597_lo_buf_o2;input n657_lo_buf_o2;input G276_o2;input n1005_lo_buf_o2;input n1161_lo_buf_o2;input G620_o2;input G629_o2;input G639_o2;input G554_o2;input G690_o2;input G698_o2;input G707_o2;input G319_o2;input G389_o2;input n753_lo_buf_o2;input G647_o2;input G769_o2;input G785_o2;input G808_o2;input G445_o2;input G448_o2;input G477_o2;input G480_o2;input G436_o2;input G786_o2;input G787_o2;input G826_o2;input G827_o2;input G825_o2;input G610_o2;input n537_lo_buf_o2;input n669_lo_buf_o2;input n969_lo_buf_o2;input n981_lo_buf_o2;input n993_lo_buf_o2;input G309_o2;input G461_o2;input G487_o2;input G460_o2;input G468_o2;input G287_o2;input G613_o2;input n585_lo_buf_o2;input n813_lo_buf_o2;input n825_lo_buf_o2;input n837_lo_buf_o2;input n897_lo_buf_o2;input n909_lo_buf_o2;input n933_lo_buf_o2;input G451_o2;input G682_o2;input G756_o2;input G542_o2;input G546_o2;input G550_o2;input G310_o2;input n798_lo_buf_o2;input n882_lo_buf_o2;input G427_o2;input G497_o2;input G499_o2;input G501_o2;input G498_o2;input G500_o2;input G502_o2;input G369_o2;input n939_lo_buf_o2;input n486_lo_buf_o2;input n510_lo_buf_o2;input n558_lo_buf_o2;input n594_lo_buf_o2;input n654_lo_buf_o2;input n477_lo_buf_o2;input n525_lo_buf_o2;input n573_lo_buf_o2;
  output G855;output G856;output G857;output G858;output G859;output G860;output G861;output G862;output G863;output G864;output G865;output G866;output G867;output G868;output G869;output G870;output G871;output G872;output G873;output G874;output G875;output G876;output G877;output G878;output G879;output G880;output n480_li;output n492_li;output n495_li;output n498_li;output n501_li;output n504_li;output n516_li;output n528_li;output n531_li;output n540_li;output n543_li;output n546_li;output n549_li;output n552_li;output n564_li;output n579_li;output n600_li;output n603_li;output n606_li;output n609_li;output n612_li;output n615_li;output n618_li;output n621_li;output n627_li;output n630_li;output n633_li;output n639_li;output n642_li;output n645_li;output n648_li;output n660_li;output n663_li;output n672_li;output n675_li;output n678_li;output n681_li;output n684_li;output n687_li;output n690_li;output n693_li;output n696_li;output n699_li;output n702_li;output n705_li;output n708_li;output n711_li;output n714_li;output n717_li;output n720_li;output n723_li;output n726_li;output n729_li;output n732_li;output n735_li;output n738_li;output n741_li;output n744_li;output n747_li;output n750_li;output n756_li;output n759_li;output n762_li;output n768_li;output n771_li;output n774_li;output n780_li;output n783_li;output n786_li;output n792_li;output n795_li;output n804_li;output n807_li;output n816_li;output n819_li;output n828_li;output n831_li;output n843_li;output n846_li;output n849_li;output n852_li;output n855_li;output n858_li;output n861_li;output n864_li;output n867_li;output n870_li;output n879_li;output n891_li;output n903_li;output n915_li;output n918_li;output n927_li;output n951_li;output n954_li;output n957_li;output n960_li;output n963_li;output n966_li;output n972_li;output n975_li;output n978_li;output n984_li;output n987_li;output n990_li;output n996_li;output n999_li;output n1002_li;output n1008_li;output n1011_li;output n1014_li;output n1020_li;output n1023_li;output n1026_li;output n1032_li;output n1035_li;output n1038_li;output n1044_li;output n1047_li;output n1050_li;output n1053_li;output n1056_li;output n1059_li;output n1062_li;output n1065_li;output n1068_li;output n1071_li;output n1074_li;output n1077_li;output n1080_li;output n1083_li;output n1086_li;output n1089_li;output n1092_li;output n1095_li;output n1098_li;output n1101_li;output n1104_li;output n1107_li;output n1110_li;output n1113_li;output n1116_li;output n1119_li;output n1122_li;output n1125_li;output n1128_li;output n1131_li;output n1134_li;output n1137_li;output n1140_li;output n1143_li;output n1146_li;output n1149_li;output n1152_li;output n1155_li;output n1158_li;output n1167_li;output n1170_li;output n1173_li;output n1176_li;output n1179_li;output n1529_i2;output n1616_i2;output n1655_i2;output n1656_i2;output n1657_i2;output n1730_i2;output n1731_i2;output n1732_i2;output n1729_i2;output n1805_i2;output n1808_i2;output n1807_i2;output n1809_i2;output n1663_i2;output n1664_i2;output n1704_i2;output n1705_i2;output n1706_i2;output n1707_i2;output n1708_i2;output n1709_i2;output G280_i2;output G655_i2;output G663_i2;output G672_i2;output G538_i2;output n1780_i2;output n1781_i2;output n1797_i2;output n1798_i2;output n1799_i2;output n1800_i2;output G578_i2;output n1828_i2;output n801_lo_buf_i2;output G693_i2;output G702_i2;output G712_i2;output G685_i2;output G658_i2;output G667_i2;output G677_i2;output G650_i2;output G798_i2;output n1017_lo_buf_i2;output n1029_lo_buf_i2;output n1041_lo_buf_i2;output G558_i2;output G562_i2;output G566_i2;output n1835_i2;output n1836_i2;output n1837_i2;output n765_lo_buf_i2;output n777_lo_buf_i2;output n789_lo_buf_i2;output G617_i2;output G626_i2;output G636_i2;output n489_lo_buf_i2;output n513_lo_buf_i2;output n561_lo_buf_i2;output n597_lo_buf_i2;output n657_lo_buf_i2;output G276_i2;output n1005_lo_buf_i2;output n1161_lo_buf_i2;output G620_i2;output G629_i2;output G639_i2;output G554_i2;output G690_i2;output G698_i2;output G707_i2;output G319_i2;output G389_i2;output n753_lo_buf_i2;output G647_i2;output G769_i2;output G785_i2;output G808_i2;output G445_i2;output G448_i2;output G477_i2;output G480_i2;output G436_i2;output G786_i2;output G787_i2;output G826_i2;output G827_i2;output G825_i2;output G610_i2;output n537_lo_buf_i2;output n669_lo_buf_i2;output n969_lo_buf_i2;output n981_lo_buf_i2;output n993_lo_buf_i2;output G309_i2;output G461_i2;output G487_i2;output G460_i2;output G468_i2;output G287_i2;output G613_i2;output n585_lo_buf_i2;output n813_lo_buf_i2;output n825_lo_buf_i2;output n837_lo_buf_i2;output n897_lo_buf_i2;output n909_lo_buf_i2;output n933_lo_buf_i2;output G451_i2;output G682_i2;output G756_i2;output G542_i2;output G546_i2;output G550_i2;output G310_i2;output n798_lo_buf_i2;output n882_lo_buf_i2;output G427_i2;output G497_i2;output G499_i2;output G501_i2;output G498_i2;output G500_i2;output G502_i2;output G369_i2;output n939_lo_buf_i2;output n486_lo_buf_i2;output n510_lo_buf_i2;output n558_lo_buf_i2;output n594_lo_buf_i2;output n654_lo_buf_i2;output n477_lo_buf_i2;output n525_lo_buf_i2;output n573_lo_buf_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire G51_p;
  wire G51_n;
  wire G52_p;
  wire G52_n;
  wire G53_p;
  wire G53_n;
  wire G54_p;
  wire G54_n;
  wire G55_p;
  wire G55_n;
  wire G56_p;
  wire G56_n;
  wire G57_p;
  wire G57_n;
  wire G58_p;
  wire G58_n;
  wire G59_p;
  wire G59_n;
  wire G60_p;
  wire G60_n;
  wire n480_lo_p;
  wire n480_lo_n;
  wire n492_lo_p;
  wire n492_lo_n;
  wire n495_lo_p;
  wire n495_lo_n;
  wire n498_lo_p;
  wire n498_lo_n;
  wire n501_lo_p;
  wire n501_lo_n;
  wire n504_lo_p;
  wire n504_lo_n;
  wire n516_lo_p;
  wire n516_lo_n;
  wire n528_lo_p;
  wire n528_lo_n;
  wire n531_lo_p;
  wire n531_lo_n;
  wire n540_lo_p;
  wire n540_lo_n;
  wire n543_lo_p;
  wire n543_lo_n;
  wire n546_lo_p;
  wire n546_lo_n;
  wire n549_lo_p;
  wire n549_lo_n;
  wire n552_lo_p;
  wire n552_lo_n;
  wire n564_lo_p;
  wire n564_lo_n;
  wire n579_lo_p;
  wire n579_lo_n;
  wire n600_lo_p;
  wire n600_lo_n;
  wire n603_lo_p;
  wire n603_lo_n;
  wire n606_lo_p;
  wire n606_lo_n;
  wire n609_lo_p;
  wire n609_lo_n;
  wire n612_lo_p;
  wire n612_lo_n;
  wire n615_lo_p;
  wire n615_lo_n;
  wire n618_lo_p;
  wire n618_lo_n;
  wire n621_lo_p;
  wire n621_lo_n;
  wire n627_lo_p;
  wire n627_lo_n;
  wire n630_lo_p;
  wire n630_lo_n;
  wire n633_lo_p;
  wire n633_lo_n;
  wire n639_lo_p;
  wire n639_lo_n;
  wire n642_lo_p;
  wire n642_lo_n;
  wire n645_lo_p;
  wire n645_lo_n;
  wire n648_lo_p;
  wire n648_lo_n;
  wire n660_lo_p;
  wire n660_lo_n;
  wire n663_lo_p;
  wire n663_lo_n;
  wire n672_lo_p;
  wire n672_lo_n;
  wire n675_lo_p;
  wire n675_lo_n;
  wire n678_lo_p;
  wire n678_lo_n;
  wire n681_lo_p;
  wire n681_lo_n;
  wire n684_lo_p;
  wire n684_lo_n;
  wire n687_lo_p;
  wire n687_lo_n;
  wire n690_lo_p;
  wire n690_lo_n;
  wire n693_lo_p;
  wire n693_lo_n;
  wire n696_lo_p;
  wire n696_lo_n;
  wire n699_lo_p;
  wire n699_lo_n;
  wire n702_lo_p;
  wire n702_lo_n;
  wire n705_lo_p;
  wire n705_lo_n;
  wire n708_lo_p;
  wire n708_lo_n;
  wire n711_lo_p;
  wire n711_lo_n;
  wire n714_lo_p;
  wire n714_lo_n;
  wire n717_lo_p;
  wire n717_lo_n;
  wire n720_lo_p;
  wire n720_lo_n;
  wire n723_lo_p;
  wire n723_lo_n;
  wire n726_lo_p;
  wire n726_lo_n;
  wire n729_lo_p;
  wire n729_lo_n;
  wire n732_lo_p;
  wire n732_lo_n;
  wire n735_lo_p;
  wire n735_lo_n;
  wire n738_lo_p;
  wire n738_lo_n;
  wire n741_lo_p;
  wire n741_lo_n;
  wire n744_lo_p;
  wire n744_lo_n;
  wire n747_lo_p;
  wire n747_lo_n;
  wire n750_lo_p;
  wire n750_lo_n;
  wire n756_lo_p;
  wire n756_lo_n;
  wire n759_lo_p;
  wire n759_lo_n;
  wire n762_lo_p;
  wire n762_lo_n;
  wire n768_lo_p;
  wire n768_lo_n;
  wire n771_lo_p;
  wire n771_lo_n;
  wire n774_lo_p;
  wire n774_lo_n;
  wire n780_lo_p;
  wire n780_lo_n;
  wire n783_lo_p;
  wire n783_lo_n;
  wire n786_lo_p;
  wire n786_lo_n;
  wire n792_lo_p;
  wire n792_lo_n;
  wire n795_lo_p;
  wire n795_lo_n;
  wire n804_lo_p;
  wire n804_lo_n;
  wire n807_lo_p;
  wire n807_lo_n;
  wire n816_lo_p;
  wire n816_lo_n;
  wire n819_lo_p;
  wire n819_lo_n;
  wire n828_lo_p;
  wire n828_lo_n;
  wire n831_lo_p;
  wire n831_lo_n;
  wire n843_lo_p;
  wire n843_lo_n;
  wire n846_lo_p;
  wire n846_lo_n;
  wire n849_lo_p;
  wire n849_lo_n;
  wire n852_lo_p;
  wire n852_lo_n;
  wire n855_lo_p;
  wire n855_lo_n;
  wire n858_lo_p;
  wire n858_lo_n;
  wire n861_lo_p;
  wire n861_lo_n;
  wire n864_lo_p;
  wire n864_lo_n;
  wire n867_lo_p;
  wire n867_lo_n;
  wire n870_lo_p;
  wire n870_lo_n;
  wire n879_lo_p;
  wire n879_lo_n;
  wire n891_lo_p;
  wire n891_lo_n;
  wire n903_lo_p;
  wire n903_lo_n;
  wire n915_lo_p;
  wire n915_lo_n;
  wire n918_lo_p;
  wire n918_lo_n;
  wire n927_lo_p;
  wire n927_lo_n;
  wire n951_lo_p;
  wire n951_lo_n;
  wire n954_lo_p;
  wire n954_lo_n;
  wire n957_lo_p;
  wire n957_lo_n;
  wire n960_lo_p;
  wire n960_lo_n;
  wire n963_lo_p;
  wire n963_lo_n;
  wire n966_lo_p;
  wire n966_lo_n;
  wire n972_lo_p;
  wire n972_lo_n;
  wire n975_lo_p;
  wire n975_lo_n;
  wire n978_lo_p;
  wire n978_lo_n;
  wire n984_lo_p;
  wire n984_lo_n;
  wire n987_lo_p;
  wire n987_lo_n;
  wire n990_lo_p;
  wire n990_lo_n;
  wire n996_lo_p;
  wire n996_lo_n;
  wire n999_lo_p;
  wire n999_lo_n;
  wire n1002_lo_p;
  wire n1002_lo_n;
  wire n1008_lo_p;
  wire n1008_lo_n;
  wire n1011_lo_p;
  wire n1011_lo_n;
  wire n1014_lo_p;
  wire n1014_lo_n;
  wire n1020_lo_p;
  wire n1020_lo_n;
  wire n1023_lo_p;
  wire n1023_lo_n;
  wire n1026_lo_p;
  wire n1026_lo_n;
  wire n1032_lo_p;
  wire n1032_lo_n;
  wire n1035_lo_p;
  wire n1035_lo_n;
  wire n1038_lo_p;
  wire n1038_lo_n;
  wire n1044_lo_p;
  wire n1044_lo_n;
  wire n1047_lo_p;
  wire n1047_lo_n;
  wire n1050_lo_p;
  wire n1050_lo_n;
  wire n1053_lo_p;
  wire n1053_lo_n;
  wire n1056_lo_p;
  wire n1056_lo_n;
  wire n1059_lo_p;
  wire n1059_lo_n;
  wire n1062_lo_p;
  wire n1062_lo_n;
  wire n1065_lo_p;
  wire n1065_lo_n;
  wire n1068_lo_p;
  wire n1068_lo_n;
  wire n1071_lo_p;
  wire n1071_lo_n;
  wire n1074_lo_p;
  wire n1074_lo_n;
  wire n1077_lo_p;
  wire n1077_lo_n;
  wire n1080_lo_p;
  wire n1080_lo_n;
  wire n1083_lo_p;
  wire n1083_lo_n;
  wire n1086_lo_p;
  wire n1086_lo_n;
  wire n1089_lo_p;
  wire n1089_lo_n;
  wire n1092_lo_p;
  wire n1092_lo_n;
  wire n1095_lo_p;
  wire n1095_lo_n;
  wire n1098_lo_p;
  wire n1098_lo_n;
  wire n1101_lo_p;
  wire n1101_lo_n;
  wire n1104_lo_p;
  wire n1104_lo_n;
  wire n1107_lo_p;
  wire n1107_lo_n;
  wire n1110_lo_p;
  wire n1110_lo_n;
  wire n1113_lo_p;
  wire n1113_lo_n;
  wire n1116_lo_p;
  wire n1116_lo_n;
  wire n1119_lo_p;
  wire n1119_lo_n;
  wire n1122_lo_p;
  wire n1122_lo_n;
  wire n1125_lo_p;
  wire n1125_lo_n;
  wire n1128_lo_p;
  wire n1128_lo_n;
  wire n1131_lo_p;
  wire n1131_lo_n;
  wire n1134_lo_p;
  wire n1134_lo_n;
  wire n1137_lo_p;
  wire n1137_lo_n;
  wire n1140_lo_p;
  wire n1140_lo_n;
  wire n1143_lo_p;
  wire n1143_lo_n;
  wire n1146_lo_p;
  wire n1146_lo_n;
  wire n1149_lo_p;
  wire n1149_lo_n;
  wire n1152_lo_p;
  wire n1152_lo_n;
  wire n1155_lo_p;
  wire n1155_lo_n;
  wire n1158_lo_p;
  wire n1158_lo_n;
  wire n1167_lo_p;
  wire n1167_lo_n;
  wire n1170_lo_p;
  wire n1170_lo_n;
  wire n1173_lo_p;
  wire n1173_lo_n;
  wire n1176_lo_p;
  wire n1176_lo_n;
  wire n1179_lo_p;
  wire n1179_lo_n;
  wire n1529_o2_p;
  wire n1529_o2_n;
  wire n1616_o2_p;
  wire n1616_o2_n;
  wire n1655_o2_p;
  wire n1655_o2_n;
  wire n1656_o2_p;
  wire n1656_o2_n;
  wire n1657_o2_p;
  wire n1657_o2_n;
  wire n1730_o2_p;
  wire n1730_o2_n;
  wire n1731_o2_p;
  wire n1731_o2_n;
  wire n1732_o2_p;
  wire n1732_o2_n;
  wire n1729_o2_p;
  wire n1729_o2_n;
  wire n1805_o2_p;
  wire n1805_o2_n;
  wire n1808_o2_p;
  wire n1808_o2_n;
  wire n1807_o2_p;
  wire n1807_o2_n;
  wire n1809_o2_p;
  wire n1809_o2_n;
  wire n1663_o2_p;
  wire n1663_o2_n;
  wire n1664_o2_p;
  wire n1664_o2_n;
  wire n1704_o2_p;
  wire n1704_o2_n;
  wire n1705_o2_p;
  wire n1705_o2_n;
  wire n1706_o2_p;
  wire n1706_o2_n;
  wire n1707_o2_p;
  wire n1707_o2_n;
  wire n1708_o2_p;
  wire n1708_o2_n;
  wire n1709_o2_p;
  wire n1709_o2_n;
  wire G280_o2_p;
  wire G280_o2_n;
  wire G655_o2_p;
  wire G655_o2_n;
  wire G663_o2_p;
  wire G663_o2_n;
  wire G672_o2_p;
  wire G672_o2_n;
  wire G538_o2_p;
  wire G538_o2_n;
  wire n1780_o2_p;
  wire n1780_o2_n;
  wire n1781_o2_p;
  wire n1781_o2_n;
  wire n1797_o2_p;
  wire n1797_o2_n;
  wire n1798_o2_p;
  wire n1798_o2_n;
  wire n1799_o2_p;
  wire n1799_o2_n;
  wire n1800_o2_p;
  wire n1800_o2_n;
  wire G578_o2_p;
  wire G578_o2_n;
  wire n1828_o2_p;
  wire n1828_o2_n;
  wire n801_lo_buf_o2_p;
  wire n801_lo_buf_o2_n;
  wire G693_o2_p;
  wire G693_o2_n;
  wire G702_o2_p;
  wire G702_o2_n;
  wire G712_o2_p;
  wire G712_o2_n;
  wire G685_o2_p;
  wire G685_o2_n;
  wire G658_o2_p;
  wire G658_o2_n;
  wire G667_o2_p;
  wire G667_o2_n;
  wire G677_o2_p;
  wire G677_o2_n;
  wire G650_o2_p;
  wire G650_o2_n;
  wire G798_o2_p;
  wire G798_o2_n;
  wire n1017_lo_buf_o2_p;
  wire n1017_lo_buf_o2_n;
  wire n1029_lo_buf_o2_p;
  wire n1029_lo_buf_o2_n;
  wire n1041_lo_buf_o2_p;
  wire n1041_lo_buf_o2_n;
  wire G558_o2_p;
  wire G558_o2_n;
  wire G562_o2_p;
  wire G562_o2_n;
  wire G566_o2_p;
  wire G566_o2_n;
  wire n1835_o2_p;
  wire n1835_o2_n;
  wire n1836_o2_p;
  wire n1836_o2_n;
  wire n1837_o2_p;
  wire n1837_o2_n;
  wire n765_lo_buf_o2_p;
  wire n765_lo_buf_o2_n;
  wire n777_lo_buf_o2_p;
  wire n777_lo_buf_o2_n;
  wire n789_lo_buf_o2_p;
  wire n789_lo_buf_o2_n;
  wire G617_o2_p;
  wire G617_o2_n;
  wire G626_o2_p;
  wire G626_o2_n;
  wire G636_o2_p;
  wire G636_o2_n;
  wire n489_lo_buf_o2_p;
  wire n489_lo_buf_o2_n;
  wire n513_lo_buf_o2_p;
  wire n513_lo_buf_o2_n;
  wire n561_lo_buf_o2_p;
  wire n561_lo_buf_o2_n;
  wire n597_lo_buf_o2_p;
  wire n597_lo_buf_o2_n;
  wire n657_lo_buf_o2_p;
  wire n657_lo_buf_o2_n;
  wire G276_o2_p;
  wire G276_o2_n;
  wire n1005_lo_buf_o2_p;
  wire n1005_lo_buf_o2_n;
  wire n1161_lo_buf_o2_p;
  wire n1161_lo_buf_o2_n;
  wire G620_o2_p;
  wire G620_o2_n;
  wire G629_o2_p;
  wire G629_o2_n;
  wire G639_o2_p;
  wire G639_o2_n;
  wire G554_o2_p;
  wire G554_o2_n;
  wire G690_o2_p;
  wire G690_o2_n;
  wire G698_o2_p;
  wire G698_o2_n;
  wire G707_o2_p;
  wire G707_o2_n;
  wire G319_o2_p;
  wire G319_o2_n;
  wire G389_o2_p;
  wire G389_o2_n;
  wire n753_lo_buf_o2_p;
  wire n753_lo_buf_o2_n;
  wire G647_o2_p;
  wire G647_o2_n;
  wire G769_o2_p;
  wire G769_o2_n;
  wire G785_o2_p;
  wire G785_o2_n;
  wire G808_o2_p;
  wire G808_o2_n;
  wire G445_o2_p;
  wire G445_o2_n;
  wire G448_o2_p;
  wire G448_o2_n;
  wire G477_o2_p;
  wire G477_o2_n;
  wire G480_o2_p;
  wire G480_o2_n;
  wire G436_o2_p;
  wire G436_o2_n;
  wire G786_o2_p;
  wire G786_o2_n;
  wire G787_o2_p;
  wire G787_o2_n;
  wire G826_o2_p;
  wire G826_o2_n;
  wire G827_o2_p;
  wire G827_o2_n;
  wire G825_o2_p;
  wire G825_o2_n;
  wire G610_o2_p;
  wire G610_o2_n;
  wire n537_lo_buf_o2_p;
  wire n537_lo_buf_o2_n;
  wire n669_lo_buf_o2_p;
  wire n669_lo_buf_o2_n;
  wire n969_lo_buf_o2_p;
  wire n969_lo_buf_o2_n;
  wire n981_lo_buf_o2_p;
  wire n981_lo_buf_o2_n;
  wire n993_lo_buf_o2_p;
  wire n993_lo_buf_o2_n;
  wire G309_o2_p;
  wire G309_o2_n;
  wire G461_o2_p;
  wire G461_o2_n;
  wire G487_o2_p;
  wire G487_o2_n;
  wire G460_o2_p;
  wire G460_o2_n;
  wire G468_o2_p;
  wire G468_o2_n;
  wire G287_o2_p;
  wire G287_o2_n;
  wire G613_o2_p;
  wire G613_o2_n;
  wire n585_lo_buf_o2_p;
  wire n585_lo_buf_o2_n;
  wire n813_lo_buf_o2_p;
  wire n813_lo_buf_o2_n;
  wire n825_lo_buf_o2_p;
  wire n825_lo_buf_o2_n;
  wire n837_lo_buf_o2_p;
  wire n837_lo_buf_o2_n;
  wire n897_lo_buf_o2_p;
  wire n897_lo_buf_o2_n;
  wire n909_lo_buf_o2_p;
  wire n909_lo_buf_o2_n;
  wire n933_lo_buf_o2_p;
  wire n933_lo_buf_o2_n;
  wire G451_o2_p;
  wire G451_o2_n;
  wire G682_o2_p;
  wire G682_o2_n;
  wire G756_o2_p;
  wire G756_o2_n;
  wire G542_o2_p;
  wire G542_o2_n;
  wire G546_o2_p;
  wire G546_o2_n;
  wire G550_o2_p;
  wire G550_o2_n;
  wire G310_o2_p;
  wire G310_o2_n;
  wire n798_lo_buf_o2_p;
  wire n798_lo_buf_o2_n;
  wire n882_lo_buf_o2_p;
  wire n882_lo_buf_o2_n;
  wire G427_o2_p;
  wire G427_o2_n;
  wire G497_o2_p;
  wire G497_o2_n;
  wire G499_o2_p;
  wire G499_o2_n;
  wire G501_o2_p;
  wire G501_o2_n;
  wire G498_o2_p;
  wire G498_o2_n;
  wire G500_o2_p;
  wire G500_o2_n;
  wire G502_o2_p;
  wire G502_o2_n;
  wire G369_o2_p;
  wire G369_o2_n;
  wire n939_lo_buf_o2_p;
  wire n939_lo_buf_o2_n;
  wire n486_lo_buf_o2_p;
  wire n486_lo_buf_o2_n;
  wire n510_lo_buf_o2_p;
  wire n510_lo_buf_o2_n;
  wire n558_lo_buf_o2_p;
  wire n558_lo_buf_o2_n;
  wire n594_lo_buf_o2_p;
  wire n594_lo_buf_o2_n;
  wire n654_lo_buf_o2_p;
  wire n654_lo_buf_o2_n;
  wire n477_lo_buf_o2_p;
  wire n477_lo_buf_o2_n;
  wire n525_lo_buf_o2_p;
  wire n525_lo_buf_o2_n;
  wire n573_lo_buf_o2_p;
  wire n573_lo_buf_o2_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire n540_lo_n_spl_;
  wire n540_lo_n_spl_0;
  wire n564_lo_n_spl_;
  wire n564_lo_n_spl_0;
  wire n552_lo_n_spl_;
  wire g361_n_spl_;
  wire n672_lo_n_spl_;
  wire n480_lo_n_spl_;
  wire n504_lo_n_spl_;
  wire n516_lo_n_spl_;
  wire g363_n_spl_;
  wire g363_n_spl_0;
  wire n600_lo_n_spl_;
  wire g374_n_spl_;
  wire g377_n_spl_;
  wire n612_lo_n_spl_;
  wire G280_o2_n_spl_;
  wire G445_o2_p_spl_;
  wire n852_lo_p_spl_;
  wire n852_lo_p_spl_0;
  wire n852_lo_p_spl_1;
  wire G445_o2_n_spl_;
  wire n852_lo_n_spl_;
  wire n852_lo_n_spl_0;
  wire n852_lo_n_spl_1;
  wire G448_o2_p_spl_;
  wire n864_lo_p_spl_;
  wire G448_o2_n_spl_;
  wire n864_lo_n_spl_;
  wire G477_o2_p_spl_;
  wire G477_o2_n_spl_;
  wire G480_o2_p_spl_;
  wire n1056_lo_p_spl_;
  wire G480_o2_n_spl_;
  wire n1056_lo_n_spl_;
  wire n1068_lo_n_spl_;
  wire n1068_lo_n_spl_0;
  wire n1068_lo_n_spl_00;
  wire n1068_lo_n_spl_01;
  wire n1068_lo_n_spl_1;
  wire n1068_lo_n_spl_10;
  wire n1068_lo_n_spl_11;
  wire n1080_lo_n_spl_;
  wire n1080_lo_n_spl_0;
  wire n1080_lo_n_spl_00;
  wire n1080_lo_n_spl_01;
  wire n1080_lo_n_spl_1;
  wire n1080_lo_n_spl_10;
  wire n1080_lo_n_spl_11;
  wire n1092_lo_n_spl_;
  wire n1092_lo_n_spl_0;
  wire n1092_lo_n_spl_00;
  wire n1092_lo_n_spl_01;
  wire n1092_lo_n_spl_1;
  wire n1092_lo_n_spl_10;
  wire n1092_lo_n_spl_11;
  wire n1104_lo_n_spl_;
  wire n1104_lo_n_spl_0;
  wire n1104_lo_n_spl_00;
  wire n1104_lo_n_spl_01;
  wire n1104_lo_n_spl_1;
  wire n1104_lo_n_spl_10;
  wire n1104_lo_n_spl_11;
  wire n1128_lo_n_spl_;
  wire n1128_lo_n_spl_0;
  wire n1116_lo_n_spl_;
  wire n1116_lo_n_spl_0;
  wire n1116_lo_n_spl_00;
  wire n1116_lo_n_spl_01;
  wire n1116_lo_n_spl_1;
  wire n1116_lo_n_spl_10;
  wire n1116_lo_n_spl_11;
  wire G436_o2_n_spl_;
  wire G436_o2_n_spl_0;
  wire G436_o2_n_spl_00;
  wire G436_o2_n_spl_01;
  wire G436_o2_n_spl_1;
  wire G436_o2_n_spl_10;
  wire G436_o2_n_spl_11;
  wire G647_o2_n_spl_;
  wire G542_o2_p_spl_;
  wire G542_o2_p_spl_0;
  wire n969_lo_buf_o2_p_spl_;
  wire n969_lo_buf_o2_p_spl_0;
  wire n969_lo_buf_o2_p_spl_00;
  wire n969_lo_buf_o2_p_spl_1;
  wire G542_o2_n_spl_;
  wire n969_lo_buf_o2_n_spl_;
  wire n969_lo_buf_o2_n_spl_0;
  wire n969_lo_buf_o2_n_spl_1;
  wire G546_o2_p_spl_;
  wire G546_o2_p_spl_0;
  wire n981_lo_buf_o2_p_spl_;
  wire n981_lo_buf_o2_p_spl_0;
  wire n981_lo_buf_o2_p_spl_00;
  wire n981_lo_buf_o2_p_spl_1;
  wire G546_o2_n_spl_;
  wire n981_lo_buf_o2_n_spl_;
  wire n981_lo_buf_o2_n_spl_0;
  wire n981_lo_buf_o2_n_spl_1;
  wire G550_o2_p_spl_;
  wire G550_o2_p_spl_0;
  wire n993_lo_buf_o2_p_spl_;
  wire n993_lo_buf_o2_p_spl_0;
  wire n993_lo_buf_o2_p_spl_00;
  wire n993_lo_buf_o2_p_spl_1;
  wire G550_o2_n_spl_;
  wire n993_lo_buf_o2_n_spl_;
  wire n993_lo_buf_o2_n_spl_0;
  wire n993_lo_buf_o2_n_spl_1;
  wire g508_p_spl_;
  wire n957_lo_n_spl_;
  wire n957_lo_n_spl_0;
  wire n957_lo_n_spl_1;
  wire g508_n_spl_;
  wire g508_n_spl_0;
  wire n957_lo_p_spl_;
  wire n957_lo_p_spl_0;
  wire n957_lo_p_spl_00;
  wire n957_lo_p_spl_1;
  wire G629_o2_p_spl_;
  wire G629_o2_p_spl_0;
  wire G629_o2_n_spl_;
  wire G629_o2_n_spl_0;
  wire G639_o2_p_spl_;
  wire G639_o2_p_spl_0;
  wire G639_o2_n_spl_;
  wire G639_o2_n_spl_0;
  wire G613_o2_p_spl_;
  wire G613_o2_n_spl_;
  wire g514_n_spl_;
  wire g514_n_spl_0;
  wire g503_n_spl_;
  wire g514_p_spl_;
  wire g514_p_spl_0;
  wire g503_p_spl_;
  wire g503_p_spl_0;
  wire g516_n_spl_;
  wire g516_n_spl_0;
  wire g516_n_spl_1;
  wire g504_n_spl_;
  wire g504_n_spl_0;
  wire g516_p_spl_;
  wire g516_p_spl_0;
  wire g516_p_spl_1;
  wire g504_p_spl_;
  wire g504_p_spl_0;
  wire g504_p_spl_1;
  wire g518_n_spl_;
  wire g518_n_spl_0;
  wire g518_n_spl_1;
  wire g505_n_spl_;
  wire g505_n_spl_0;
  wire g505_n_spl_1;
  wire g518_p_spl_;
  wire g518_p_spl_0;
  wire g518_p_spl_1;
  wire g505_p_spl_;
  wire g505_p_spl_0;
  wire g505_p_spl_00;
  wire g505_p_spl_1;
  wire g509_n_spl_;
  wire g520_p_spl_;
  wire g523_p_spl_;
  wire g523_n_spl_;
  wire G756_o2_p_spl_;
  wire G756_o2_n_spl_;
  wire G682_o2_p_spl_;
  wire g526_n_spl_;
  wire g526_n_spl_0;
  wire g526_n_spl_1;
  wire g526_p_spl_;
  wire g526_p_spl_0;
  wire g526_p_spl_1;
  wire G369_o2_p_spl_;
  wire g532_n_spl_;
  wire g532_n_spl_0;
  wire g532_n_spl_1;
  wire g534_p_spl_;
  wire g534_p_spl_0;
  wire n1014_lo_n_spl_;
  wire g536_p_spl_;
  wire g536_p_spl_0;
  wire n1026_lo_n_spl_;
  wire g538_p_spl_;
  wire g538_p_spl_0;
  wire n1038_lo_n_spl_;
  wire n525_lo_buf_o2_p_spl_;
  wire n477_lo_buf_o2_p_spl_;
  wire n477_lo_buf_o2_p_spl_0;
  wire n477_lo_buf_o2_n_spl_;
  wire n573_lo_buf_o2_p_spl_;
  wire n573_lo_buf_o2_p_spl_0;
  wire n882_lo_buf_o2_n_spl_;
  wire G451_o2_n_spl_;
  wire G451_o2_n_spl_0;
  wire G451_o2_n_spl_1;
  wire n594_lo_buf_o2_n_spl_;
  wire g512_p_spl_;
  wire n1161_lo_buf_o2_p_spl_;
  wire n1161_lo_buf_o2_p_spl_0;
  wire n1161_lo_buf_o2_n_spl_;
  wire n1161_lo_buf_o2_n_spl_0;
  wire g513_p_spl_;
  wire g519_p_spl_;
  wire n753_lo_buf_o2_p_spl_;
  wire n753_lo_buf_o2_p_spl_0;
  wire n765_lo_buf_o2_p_spl_;
  wire n765_lo_buf_o2_p_spl_0;
  wire n753_lo_buf_o2_n_spl_;
  wire n765_lo_buf_o2_n_spl_;
  wire n789_lo_buf_o2_p_spl_;
  wire n789_lo_buf_o2_p_spl_0;
  wire n777_lo_buf_o2_p_spl_;
  wire n777_lo_buf_o2_p_spl_0;
  wire n789_lo_buf_o2_n_spl_;
  wire n777_lo_buf_o2_n_spl_;
  wire n801_lo_buf_o2_p_spl_;
  wire n801_lo_buf_o2_p_spl_0;
  wire n1798_o2_p_spl_;
  wire n1798_o2_p_spl_0;
  wire n801_lo_buf_o2_n_spl_;
  wire n1798_o2_n_spl_;
  wire n1800_o2_p_spl_;
  wire n1799_o2_p_spl_;
  wire n1799_o2_p_spl_0;
  wire n1800_o2_n_spl_;
  wire n1799_o2_n_spl_;
  wire n1005_lo_buf_o2_p_spl_;
  wire n1005_lo_buf_o2_p_spl_0;
  wire n1017_lo_buf_o2_p_spl_;
  wire n1017_lo_buf_o2_p_spl_0;
  wire n1005_lo_buf_o2_n_spl_;
  wire n1017_lo_buf_o2_n_spl_;
  wire n1041_lo_buf_o2_p_spl_;
  wire n1041_lo_buf_o2_p_spl_0;
  wire n1029_lo_buf_o2_p_spl_;
  wire n1029_lo_buf_o2_p_spl_0;
  wire n1041_lo_buf_o2_n_spl_;
  wire n1029_lo_buf_o2_n_spl_;
  wire g502_n_spl_;
  wire G707_o2_p_spl_;
  wire G707_o2_p_spl_0;
  wire G707_o2_n_spl_;
  wire G698_o2_p_spl_;
  wire g510_p_spl_;
  wire g511_p_spl_;
  wire g515_p_spl_;
  wire g517_p_spl_;
  wire g531_n_spl_;
  wire g521_p_spl_;
  wire g550_p_spl_;
  wire g550_p_spl_0;
  wire n1002_lo_n_spl_;
  wire n489_lo_buf_o2_p_spl_;
  wire G389_o2_n_spl_;
  wire n513_lo_buf_o2_n_spl_;
  wire n750_lo_p_spl_;
  wire g638_n_spl_;
  wire g638_n_spl_0;
  wire g638_n_spl_1;
  wire g551_n_spl_;
  wire g543_p_spl_;
  wire g543_p_spl_0;
  wire g543_p_spl_1;
  wire n510_lo_buf_o2_p_spl_;
  wire n510_lo_buf_o2_p_spl_0;
  wire n510_lo_buf_o2_p_spl_1;
  wire n654_lo_buf_o2_n_spl_;
  wire n558_lo_buf_o2_p_spl_;
  wire n558_lo_buf_o2_n_spl_;
  wire n594_lo_buf_o2_p_spl_;
  wire n486_lo_buf_o2_p_spl_;
  wire g544_p_spl_;
  wire g544_p_spl_0;
  wire g540_n_spl_;
  wire g540_n_spl_0;
  wire g545_p_spl_;
  wire g660_n_spl_;
  wire g541_n_spl_;
  wire g541_n_spl_0;
  wire g546_p_spl_;
  wire g539_n_spl_;
  wire g539_n_spl_0;
  wire n870_lo_n_spl_;
  wire n870_lo_n_spl_0;
  wire g635_n_spl_;
  wire g635_n_spl_0;
  wire g635_n_spl_1;
  wire g644_n_spl_;
  wire g642_n_spl_;
  wire g642_n_spl_0;
  wire g642_n_spl_1;
  wire n891_lo_p_spl_;
  wire n903_lo_p_spl_;
  wire n927_lo_p_spl_;
  wire g658_n_spl_;
  wire g658_n_spl_0;
  wire g658_n_spl_1;
  wire n807_lo_p_spl_;
  wire n819_lo_p_spl_;
  wire n831_lo_p_spl_;
  wire g631_n_spl_;
  wire n1179_lo_p_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  buf

  (
    G42_p,
    G42
  );


  not

  (
    G42_n,
    G42
  );


  buf

  (
    G43_p,
    G43
  );


  not

  (
    G43_n,
    G43
  );


  buf

  (
    G44_p,
    G44
  );


  not

  (
    G44_n,
    G44
  );


  buf

  (
    G45_p,
    G45
  );


  not

  (
    G45_n,
    G45
  );


  buf

  (
    G46_p,
    G46
  );


  not

  (
    G46_n,
    G46
  );


  buf

  (
    G47_p,
    G47
  );


  not

  (
    G47_n,
    G47
  );


  buf

  (
    G48_p,
    G48
  );


  not

  (
    G48_n,
    G48
  );


  buf

  (
    G49_p,
    G49
  );


  not

  (
    G49_n,
    G49
  );


  buf

  (
    G50_p,
    G50
  );


  not

  (
    G50_n,
    G50
  );


  buf

  (
    G51_p,
    G51
  );


  not

  (
    G51_n,
    G51
  );


  buf

  (
    G52_p,
    G52
  );


  not

  (
    G52_n,
    G52
  );


  buf

  (
    G53_p,
    G53
  );


  not

  (
    G53_n,
    G53
  );


  buf

  (
    G54_p,
    G54
  );


  not

  (
    G54_n,
    G54
  );


  buf

  (
    G55_p,
    G55
  );


  not

  (
    G55_n,
    G55
  );


  buf

  (
    G56_p,
    G56
  );


  not

  (
    G56_n,
    G56
  );


  buf

  (
    G57_p,
    G57
  );


  not

  (
    G57_n,
    G57
  );


  buf

  (
    G58_p,
    G58
  );


  not

  (
    G58_n,
    G58
  );


  buf

  (
    G59_p,
    G59
  );


  not

  (
    G59_n,
    G59
  );


  buf

  (
    G60_p,
    G60
  );


  not

  (
    G60_n,
    G60
  );


  buf

  (
    n480_lo_p,
    n480_lo
  );


  not

  (
    n480_lo_n,
    n480_lo
  );


  buf

  (
    n492_lo_p,
    n492_lo
  );


  not

  (
    n492_lo_n,
    n492_lo
  );


  buf

  (
    n495_lo_p,
    n495_lo
  );


  not

  (
    n495_lo_n,
    n495_lo
  );


  buf

  (
    n498_lo_p,
    n498_lo
  );


  not

  (
    n498_lo_n,
    n498_lo
  );


  buf

  (
    n501_lo_p,
    n501_lo
  );


  not

  (
    n501_lo_n,
    n501_lo
  );


  buf

  (
    n504_lo_p,
    n504_lo
  );


  not

  (
    n504_lo_n,
    n504_lo
  );


  buf

  (
    n516_lo_p,
    n516_lo
  );


  not

  (
    n516_lo_n,
    n516_lo
  );


  buf

  (
    n528_lo_p,
    n528_lo
  );


  not

  (
    n528_lo_n,
    n528_lo
  );


  buf

  (
    n531_lo_p,
    n531_lo
  );


  not

  (
    n531_lo_n,
    n531_lo
  );


  buf

  (
    n540_lo_p,
    n540_lo
  );


  not

  (
    n540_lo_n,
    n540_lo
  );


  buf

  (
    n543_lo_p,
    n543_lo
  );


  not

  (
    n543_lo_n,
    n543_lo
  );


  buf

  (
    n546_lo_p,
    n546_lo
  );


  not

  (
    n546_lo_n,
    n546_lo
  );


  buf

  (
    n549_lo_p,
    n549_lo
  );


  not

  (
    n549_lo_n,
    n549_lo
  );


  buf

  (
    n552_lo_p,
    n552_lo
  );


  not

  (
    n552_lo_n,
    n552_lo
  );


  buf

  (
    n564_lo_p,
    n564_lo
  );


  not

  (
    n564_lo_n,
    n564_lo
  );


  buf

  (
    n579_lo_p,
    n579_lo
  );


  not

  (
    n579_lo_n,
    n579_lo
  );


  buf

  (
    n600_lo_p,
    n600_lo
  );


  not

  (
    n600_lo_n,
    n600_lo
  );


  buf

  (
    n603_lo_p,
    n603_lo
  );


  not

  (
    n603_lo_n,
    n603_lo
  );


  buf

  (
    n606_lo_p,
    n606_lo
  );


  not

  (
    n606_lo_n,
    n606_lo
  );


  buf

  (
    n609_lo_p,
    n609_lo
  );


  not

  (
    n609_lo_n,
    n609_lo
  );


  buf

  (
    n612_lo_p,
    n612_lo
  );


  not

  (
    n612_lo_n,
    n612_lo
  );


  buf

  (
    n615_lo_p,
    n615_lo
  );


  not

  (
    n615_lo_n,
    n615_lo
  );


  buf

  (
    n618_lo_p,
    n618_lo
  );


  not

  (
    n618_lo_n,
    n618_lo
  );


  buf

  (
    n621_lo_p,
    n621_lo
  );


  not

  (
    n621_lo_n,
    n621_lo
  );


  buf

  (
    n627_lo_p,
    n627_lo
  );


  not

  (
    n627_lo_n,
    n627_lo
  );


  buf

  (
    n630_lo_p,
    n630_lo
  );


  not

  (
    n630_lo_n,
    n630_lo
  );


  buf

  (
    n633_lo_p,
    n633_lo
  );


  not

  (
    n633_lo_n,
    n633_lo
  );


  buf

  (
    n639_lo_p,
    n639_lo
  );


  not

  (
    n639_lo_n,
    n639_lo
  );


  buf

  (
    n642_lo_p,
    n642_lo
  );


  not

  (
    n642_lo_n,
    n642_lo
  );


  buf

  (
    n645_lo_p,
    n645_lo
  );


  not

  (
    n645_lo_n,
    n645_lo
  );


  buf

  (
    n648_lo_p,
    n648_lo
  );


  not

  (
    n648_lo_n,
    n648_lo
  );


  buf

  (
    n660_lo_p,
    n660_lo
  );


  not

  (
    n660_lo_n,
    n660_lo
  );


  buf

  (
    n663_lo_p,
    n663_lo
  );


  not

  (
    n663_lo_n,
    n663_lo
  );


  buf

  (
    n672_lo_p,
    n672_lo
  );


  not

  (
    n672_lo_n,
    n672_lo
  );


  buf

  (
    n675_lo_p,
    n675_lo
  );


  not

  (
    n675_lo_n,
    n675_lo
  );


  buf

  (
    n678_lo_p,
    n678_lo
  );


  not

  (
    n678_lo_n,
    n678_lo
  );


  buf

  (
    n681_lo_p,
    n681_lo
  );


  not

  (
    n681_lo_n,
    n681_lo
  );


  buf

  (
    n684_lo_p,
    n684_lo
  );


  not

  (
    n684_lo_n,
    n684_lo
  );


  buf

  (
    n687_lo_p,
    n687_lo
  );


  not

  (
    n687_lo_n,
    n687_lo
  );


  buf

  (
    n690_lo_p,
    n690_lo
  );


  not

  (
    n690_lo_n,
    n690_lo
  );


  buf

  (
    n693_lo_p,
    n693_lo
  );


  not

  (
    n693_lo_n,
    n693_lo
  );


  buf

  (
    n696_lo_p,
    n696_lo
  );


  not

  (
    n696_lo_n,
    n696_lo
  );


  buf

  (
    n699_lo_p,
    n699_lo
  );


  not

  (
    n699_lo_n,
    n699_lo
  );


  buf

  (
    n702_lo_p,
    n702_lo
  );


  not

  (
    n702_lo_n,
    n702_lo
  );


  buf

  (
    n705_lo_p,
    n705_lo
  );


  not

  (
    n705_lo_n,
    n705_lo
  );


  buf

  (
    n708_lo_p,
    n708_lo
  );


  not

  (
    n708_lo_n,
    n708_lo
  );


  buf

  (
    n711_lo_p,
    n711_lo
  );


  not

  (
    n711_lo_n,
    n711_lo
  );


  buf

  (
    n714_lo_p,
    n714_lo
  );


  not

  (
    n714_lo_n,
    n714_lo
  );


  buf

  (
    n717_lo_p,
    n717_lo
  );


  not

  (
    n717_lo_n,
    n717_lo
  );


  buf

  (
    n720_lo_p,
    n720_lo
  );


  not

  (
    n720_lo_n,
    n720_lo
  );


  buf

  (
    n723_lo_p,
    n723_lo
  );


  not

  (
    n723_lo_n,
    n723_lo
  );


  buf

  (
    n726_lo_p,
    n726_lo
  );


  not

  (
    n726_lo_n,
    n726_lo
  );


  buf

  (
    n729_lo_p,
    n729_lo
  );


  not

  (
    n729_lo_n,
    n729_lo
  );


  buf

  (
    n732_lo_p,
    n732_lo
  );


  not

  (
    n732_lo_n,
    n732_lo
  );


  buf

  (
    n735_lo_p,
    n735_lo
  );


  not

  (
    n735_lo_n,
    n735_lo
  );


  buf

  (
    n738_lo_p,
    n738_lo
  );


  not

  (
    n738_lo_n,
    n738_lo
  );


  buf

  (
    n741_lo_p,
    n741_lo
  );


  not

  (
    n741_lo_n,
    n741_lo
  );


  buf

  (
    n744_lo_p,
    n744_lo
  );


  not

  (
    n744_lo_n,
    n744_lo
  );


  buf

  (
    n747_lo_p,
    n747_lo
  );


  not

  (
    n747_lo_n,
    n747_lo
  );


  buf

  (
    n750_lo_p,
    n750_lo
  );


  not

  (
    n750_lo_n,
    n750_lo
  );


  buf

  (
    n756_lo_p,
    n756_lo
  );


  not

  (
    n756_lo_n,
    n756_lo
  );


  buf

  (
    n759_lo_p,
    n759_lo
  );


  not

  (
    n759_lo_n,
    n759_lo
  );


  buf

  (
    n762_lo_p,
    n762_lo
  );


  not

  (
    n762_lo_n,
    n762_lo
  );


  buf

  (
    n768_lo_p,
    n768_lo
  );


  not

  (
    n768_lo_n,
    n768_lo
  );


  buf

  (
    n771_lo_p,
    n771_lo
  );


  not

  (
    n771_lo_n,
    n771_lo
  );


  buf

  (
    n774_lo_p,
    n774_lo
  );


  not

  (
    n774_lo_n,
    n774_lo
  );


  buf

  (
    n780_lo_p,
    n780_lo
  );


  not

  (
    n780_lo_n,
    n780_lo
  );


  buf

  (
    n783_lo_p,
    n783_lo
  );


  not

  (
    n783_lo_n,
    n783_lo
  );


  buf

  (
    n786_lo_p,
    n786_lo
  );


  not

  (
    n786_lo_n,
    n786_lo
  );


  buf

  (
    n792_lo_p,
    n792_lo
  );


  not

  (
    n792_lo_n,
    n792_lo
  );


  buf

  (
    n795_lo_p,
    n795_lo
  );


  not

  (
    n795_lo_n,
    n795_lo
  );


  buf

  (
    n804_lo_p,
    n804_lo
  );


  not

  (
    n804_lo_n,
    n804_lo
  );


  buf

  (
    n807_lo_p,
    n807_lo
  );


  not

  (
    n807_lo_n,
    n807_lo
  );


  buf

  (
    n816_lo_p,
    n816_lo
  );


  not

  (
    n816_lo_n,
    n816_lo
  );


  buf

  (
    n819_lo_p,
    n819_lo
  );


  not

  (
    n819_lo_n,
    n819_lo
  );


  buf

  (
    n828_lo_p,
    n828_lo
  );


  not

  (
    n828_lo_n,
    n828_lo
  );


  buf

  (
    n831_lo_p,
    n831_lo
  );


  not

  (
    n831_lo_n,
    n831_lo
  );


  buf

  (
    n843_lo_p,
    n843_lo
  );


  not

  (
    n843_lo_n,
    n843_lo
  );


  buf

  (
    n846_lo_p,
    n846_lo
  );


  not

  (
    n846_lo_n,
    n846_lo
  );


  buf

  (
    n849_lo_p,
    n849_lo
  );


  not

  (
    n849_lo_n,
    n849_lo
  );


  buf

  (
    n852_lo_p,
    n852_lo
  );


  not

  (
    n852_lo_n,
    n852_lo
  );


  buf

  (
    n855_lo_p,
    n855_lo
  );


  not

  (
    n855_lo_n,
    n855_lo
  );


  buf

  (
    n858_lo_p,
    n858_lo
  );


  not

  (
    n858_lo_n,
    n858_lo
  );


  buf

  (
    n861_lo_p,
    n861_lo
  );


  not

  (
    n861_lo_n,
    n861_lo
  );


  buf

  (
    n864_lo_p,
    n864_lo
  );


  not

  (
    n864_lo_n,
    n864_lo
  );


  buf

  (
    n867_lo_p,
    n867_lo
  );


  not

  (
    n867_lo_n,
    n867_lo
  );


  buf

  (
    n870_lo_p,
    n870_lo
  );


  not

  (
    n870_lo_n,
    n870_lo
  );


  buf

  (
    n879_lo_p,
    n879_lo
  );


  not

  (
    n879_lo_n,
    n879_lo
  );


  buf

  (
    n891_lo_p,
    n891_lo
  );


  not

  (
    n891_lo_n,
    n891_lo
  );


  buf

  (
    n903_lo_p,
    n903_lo
  );


  not

  (
    n903_lo_n,
    n903_lo
  );


  buf

  (
    n915_lo_p,
    n915_lo
  );


  not

  (
    n915_lo_n,
    n915_lo
  );


  buf

  (
    n918_lo_p,
    n918_lo
  );


  not

  (
    n918_lo_n,
    n918_lo
  );


  buf

  (
    n927_lo_p,
    n927_lo
  );


  not

  (
    n927_lo_n,
    n927_lo
  );


  buf

  (
    n951_lo_p,
    n951_lo
  );


  not

  (
    n951_lo_n,
    n951_lo
  );


  buf

  (
    n954_lo_p,
    n954_lo
  );


  not

  (
    n954_lo_n,
    n954_lo
  );


  buf

  (
    n957_lo_p,
    n957_lo
  );


  not

  (
    n957_lo_n,
    n957_lo
  );


  buf

  (
    n960_lo_p,
    n960_lo
  );


  not

  (
    n960_lo_n,
    n960_lo
  );


  buf

  (
    n963_lo_p,
    n963_lo
  );


  not

  (
    n963_lo_n,
    n963_lo
  );


  buf

  (
    n966_lo_p,
    n966_lo
  );


  not

  (
    n966_lo_n,
    n966_lo
  );


  buf

  (
    n972_lo_p,
    n972_lo
  );


  not

  (
    n972_lo_n,
    n972_lo
  );


  buf

  (
    n975_lo_p,
    n975_lo
  );


  not

  (
    n975_lo_n,
    n975_lo
  );


  buf

  (
    n978_lo_p,
    n978_lo
  );


  not

  (
    n978_lo_n,
    n978_lo
  );


  buf

  (
    n984_lo_p,
    n984_lo
  );


  not

  (
    n984_lo_n,
    n984_lo
  );


  buf

  (
    n987_lo_p,
    n987_lo
  );


  not

  (
    n987_lo_n,
    n987_lo
  );


  buf

  (
    n990_lo_p,
    n990_lo
  );


  not

  (
    n990_lo_n,
    n990_lo
  );


  buf

  (
    n996_lo_p,
    n996_lo
  );


  not

  (
    n996_lo_n,
    n996_lo
  );


  buf

  (
    n999_lo_p,
    n999_lo
  );


  not

  (
    n999_lo_n,
    n999_lo
  );


  buf

  (
    n1002_lo_p,
    n1002_lo
  );


  not

  (
    n1002_lo_n,
    n1002_lo
  );


  buf

  (
    n1008_lo_p,
    n1008_lo
  );


  not

  (
    n1008_lo_n,
    n1008_lo
  );


  buf

  (
    n1011_lo_p,
    n1011_lo
  );


  not

  (
    n1011_lo_n,
    n1011_lo
  );


  buf

  (
    n1014_lo_p,
    n1014_lo
  );


  not

  (
    n1014_lo_n,
    n1014_lo
  );


  buf

  (
    n1020_lo_p,
    n1020_lo
  );


  not

  (
    n1020_lo_n,
    n1020_lo
  );


  buf

  (
    n1023_lo_p,
    n1023_lo
  );


  not

  (
    n1023_lo_n,
    n1023_lo
  );


  buf

  (
    n1026_lo_p,
    n1026_lo
  );


  not

  (
    n1026_lo_n,
    n1026_lo
  );


  buf

  (
    n1032_lo_p,
    n1032_lo
  );


  not

  (
    n1032_lo_n,
    n1032_lo
  );


  buf

  (
    n1035_lo_p,
    n1035_lo
  );


  not

  (
    n1035_lo_n,
    n1035_lo
  );


  buf

  (
    n1038_lo_p,
    n1038_lo
  );


  not

  (
    n1038_lo_n,
    n1038_lo
  );


  buf

  (
    n1044_lo_p,
    n1044_lo
  );


  not

  (
    n1044_lo_n,
    n1044_lo
  );


  buf

  (
    n1047_lo_p,
    n1047_lo
  );


  not

  (
    n1047_lo_n,
    n1047_lo
  );


  buf

  (
    n1050_lo_p,
    n1050_lo
  );


  not

  (
    n1050_lo_n,
    n1050_lo
  );


  buf

  (
    n1053_lo_p,
    n1053_lo
  );


  not

  (
    n1053_lo_n,
    n1053_lo
  );


  buf

  (
    n1056_lo_p,
    n1056_lo
  );


  not

  (
    n1056_lo_n,
    n1056_lo
  );


  buf

  (
    n1059_lo_p,
    n1059_lo
  );


  not

  (
    n1059_lo_n,
    n1059_lo
  );


  buf

  (
    n1062_lo_p,
    n1062_lo
  );


  not

  (
    n1062_lo_n,
    n1062_lo
  );


  buf

  (
    n1065_lo_p,
    n1065_lo
  );


  not

  (
    n1065_lo_n,
    n1065_lo
  );


  buf

  (
    n1068_lo_p,
    n1068_lo
  );


  not

  (
    n1068_lo_n,
    n1068_lo
  );


  buf

  (
    n1071_lo_p,
    n1071_lo
  );


  not

  (
    n1071_lo_n,
    n1071_lo
  );


  buf

  (
    n1074_lo_p,
    n1074_lo
  );


  not

  (
    n1074_lo_n,
    n1074_lo
  );


  buf

  (
    n1077_lo_p,
    n1077_lo
  );


  not

  (
    n1077_lo_n,
    n1077_lo
  );


  buf

  (
    n1080_lo_p,
    n1080_lo
  );


  not

  (
    n1080_lo_n,
    n1080_lo
  );


  buf

  (
    n1083_lo_p,
    n1083_lo
  );


  not

  (
    n1083_lo_n,
    n1083_lo
  );


  buf

  (
    n1086_lo_p,
    n1086_lo
  );


  not

  (
    n1086_lo_n,
    n1086_lo
  );


  buf

  (
    n1089_lo_p,
    n1089_lo
  );


  not

  (
    n1089_lo_n,
    n1089_lo
  );


  buf

  (
    n1092_lo_p,
    n1092_lo
  );


  not

  (
    n1092_lo_n,
    n1092_lo
  );


  buf

  (
    n1095_lo_p,
    n1095_lo
  );


  not

  (
    n1095_lo_n,
    n1095_lo
  );


  buf

  (
    n1098_lo_p,
    n1098_lo
  );


  not

  (
    n1098_lo_n,
    n1098_lo
  );


  buf

  (
    n1101_lo_p,
    n1101_lo
  );


  not

  (
    n1101_lo_n,
    n1101_lo
  );


  buf

  (
    n1104_lo_p,
    n1104_lo
  );


  not

  (
    n1104_lo_n,
    n1104_lo
  );


  buf

  (
    n1107_lo_p,
    n1107_lo
  );


  not

  (
    n1107_lo_n,
    n1107_lo
  );


  buf

  (
    n1110_lo_p,
    n1110_lo
  );


  not

  (
    n1110_lo_n,
    n1110_lo
  );


  buf

  (
    n1113_lo_p,
    n1113_lo
  );


  not

  (
    n1113_lo_n,
    n1113_lo
  );


  buf

  (
    n1116_lo_p,
    n1116_lo
  );


  not

  (
    n1116_lo_n,
    n1116_lo
  );


  buf

  (
    n1119_lo_p,
    n1119_lo
  );


  not

  (
    n1119_lo_n,
    n1119_lo
  );


  buf

  (
    n1122_lo_p,
    n1122_lo
  );


  not

  (
    n1122_lo_n,
    n1122_lo
  );


  buf

  (
    n1125_lo_p,
    n1125_lo
  );


  not

  (
    n1125_lo_n,
    n1125_lo
  );


  buf

  (
    n1128_lo_p,
    n1128_lo
  );


  not

  (
    n1128_lo_n,
    n1128_lo
  );


  buf

  (
    n1131_lo_p,
    n1131_lo
  );


  not

  (
    n1131_lo_n,
    n1131_lo
  );


  buf

  (
    n1134_lo_p,
    n1134_lo
  );


  not

  (
    n1134_lo_n,
    n1134_lo
  );


  buf

  (
    n1137_lo_p,
    n1137_lo
  );


  not

  (
    n1137_lo_n,
    n1137_lo
  );


  buf

  (
    n1140_lo_p,
    n1140_lo
  );


  not

  (
    n1140_lo_n,
    n1140_lo
  );


  buf

  (
    n1143_lo_p,
    n1143_lo
  );


  not

  (
    n1143_lo_n,
    n1143_lo
  );


  buf

  (
    n1146_lo_p,
    n1146_lo
  );


  not

  (
    n1146_lo_n,
    n1146_lo
  );


  buf

  (
    n1149_lo_p,
    n1149_lo
  );


  not

  (
    n1149_lo_n,
    n1149_lo
  );


  buf

  (
    n1152_lo_p,
    n1152_lo
  );


  not

  (
    n1152_lo_n,
    n1152_lo
  );


  buf

  (
    n1155_lo_p,
    n1155_lo
  );


  not

  (
    n1155_lo_n,
    n1155_lo
  );


  buf

  (
    n1158_lo_p,
    n1158_lo
  );


  not

  (
    n1158_lo_n,
    n1158_lo
  );


  buf

  (
    n1167_lo_p,
    n1167_lo
  );


  not

  (
    n1167_lo_n,
    n1167_lo
  );


  buf

  (
    n1170_lo_p,
    n1170_lo
  );


  not

  (
    n1170_lo_n,
    n1170_lo
  );


  buf

  (
    n1173_lo_p,
    n1173_lo
  );


  not

  (
    n1173_lo_n,
    n1173_lo
  );


  buf

  (
    n1176_lo_p,
    n1176_lo
  );


  not

  (
    n1176_lo_n,
    n1176_lo
  );


  buf

  (
    n1179_lo_p,
    n1179_lo
  );


  not

  (
    n1179_lo_n,
    n1179_lo
  );


  buf

  (
    n1529_o2_p,
    n1529_o2
  );


  not

  (
    n1529_o2_n,
    n1529_o2
  );


  buf

  (
    n1616_o2_p,
    n1616_o2
  );


  not

  (
    n1616_o2_n,
    n1616_o2
  );


  buf

  (
    n1655_o2_p,
    n1655_o2
  );


  not

  (
    n1655_o2_n,
    n1655_o2
  );


  buf

  (
    n1656_o2_p,
    n1656_o2
  );


  not

  (
    n1656_o2_n,
    n1656_o2
  );


  buf

  (
    n1657_o2_p,
    n1657_o2
  );


  not

  (
    n1657_o2_n,
    n1657_o2
  );


  buf

  (
    n1730_o2_p,
    n1730_o2
  );


  not

  (
    n1730_o2_n,
    n1730_o2
  );


  buf

  (
    n1731_o2_p,
    n1731_o2
  );


  not

  (
    n1731_o2_n,
    n1731_o2
  );


  buf

  (
    n1732_o2_p,
    n1732_o2
  );


  not

  (
    n1732_o2_n,
    n1732_o2
  );


  buf

  (
    n1729_o2_p,
    n1729_o2
  );


  not

  (
    n1729_o2_n,
    n1729_o2
  );


  buf

  (
    n1805_o2_p,
    n1805_o2
  );


  not

  (
    n1805_o2_n,
    n1805_o2
  );


  buf

  (
    n1808_o2_p,
    n1808_o2
  );


  not

  (
    n1808_o2_n,
    n1808_o2
  );


  buf

  (
    n1807_o2_p,
    n1807_o2
  );


  not

  (
    n1807_o2_n,
    n1807_o2
  );


  buf

  (
    n1809_o2_p,
    n1809_o2
  );


  not

  (
    n1809_o2_n,
    n1809_o2
  );


  buf

  (
    n1663_o2_p,
    n1663_o2
  );


  not

  (
    n1663_o2_n,
    n1663_o2
  );


  buf

  (
    n1664_o2_p,
    n1664_o2
  );


  not

  (
    n1664_o2_n,
    n1664_o2
  );


  buf

  (
    n1704_o2_p,
    n1704_o2
  );


  not

  (
    n1704_o2_n,
    n1704_o2
  );


  buf

  (
    n1705_o2_p,
    n1705_o2
  );


  not

  (
    n1705_o2_n,
    n1705_o2
  );


  buf

  (
    n1706_o2_p,
    n1706_o2
  );


  not

  (
    n1706_o2_n,
    n1706_o2
  );


  buf

  (
    n1707_o2_p,
    n1707_o2
  );


  not

  (
    n1707_o2_n,
    n1707_o2
  );


  buf

  (
    n1708_o2_p,
    n1708_o2
  );


  not

  (
    n1708_o2_n,
    n1708_o2
  );


  buf

  (
    n1709_o2_p,
    n1709_o2
  );


  not

  (
    n1709_o2_n,
    n1709_o2
  );


  buf

  (
    G280_o2_p,
    G280_o2
  );


  not

  (
    G280_o2_n,
    G280_o2
  );


  buf

  (
    G655_o2_p,
    G655_o2
  );


  not

  (
    G655_o2_n,
    G655_o2
  );


  buf

  (
    G663_o2_p,
    G663_o2
  );


  not

  (
    G663_o2_n,
    G663_o2
  );


  buf

  (
    G672_o2_p,
    G672_o2
  );


  not

  (
    G672_o2_n,
    G672_o2
  );


  buf

  (
    G538_o2_p,
    G538_o2
  );


  not

  (
    G538_o2_n,
    G538_o2
  );


  buf

  (
    n1780_o2_p,
    n1780_o2
  );


  not

  (
    n1780_o2_n,
    n1780_o2
  );


  buf

  (
    n1781_o2_p,
    n1781_o2
  );


  not

  (
    n1781_o2_n,
    n1781_o2
  );


  buf

  (
    n1797_o2_p,
    n1797_o2
  );


  not

  (
    n1797_o2_n,
    n1797_o2
  );


  buf

  (
    n1798_o2_p,
    n1798_o2
  );


  not

  (
    n1798_o2_n,
    n1798_o2
  );


  buf

  (
    n1799_o2_p,
    n1799_o2
  );


  not

  (
    n1799_o2_n,
    n1799_o2
  );


  buf

  (
    n1800_o2_p,
    n1800_o2
  );


  not

  (
    n1800_o2_n,
    n1800_o2
  );


  buf

  (
    G578_o2_p,
    G578_o2
  );


  not

  (
    G578_o2_n,
    G578_o2
  );


  buf

  (
    n1828_o2_p,
    n1828_o2
  );


  not

  (
    n1828_o2_n,
    n1828_o2
  );


  buf

  (
    n801_lo_buf_o2_p,
    n801_lo_buf_o2
  );


  not

  (
    n801_lo_buf_o2_n,
    n801_lo_buf_o2
  );


  buf

  (
    G693_o2_p,
    G693_o2
  );


  not

  (
    G693_o2_n,
    G693_o2
  );


  buf

  (
    G702_o2_p,
    G702_o2
  );


  not

  (
    G702_o2_n,
    G702_o2
  );


  buf

  (
    G712_o2_p,
    G712_o2
  );


  not

  (
    G712_o2_n,
    G712_o2
  );


  buf

  (
    G685_o2_p,
    G685_o2
  );


  not

  (
    G685_o2_n,
    G685_o2
  );


  buf

  (
    G658_o2_p,
    G658_o2
  );


  not

  (
    G658_o2_n,
    G658_o2
  );


  buf

  (
    G667_o2_p,
    G667_o2
  );


  not

  (
    G667_o2_n,
    G667_o2
  );


  buf

  (
    G677_o2_p,
    G677_o2
  );


  not

  (
    G677_o2_n,
    G677_o2
  );


  buf

  (
    G650_o2_p,
    G650_o2
  );


  not

  (
    G650_o2_n,
    G650_o2
  );


  buf

  (
    G798_o2_p,
    G798_o2
  );


  not

  (
    G798_o2_n,
    G798_o2
  );


  buf

  (
    n1017_lo_buf_o2_p,
    n1017_lo_buf_o2
  );


  not

  (
    n1017_lo_buf_o2_n,
    n1017_lo_buf_o2
  );


  buf

  (
    n1029_lo_buf_o2_p,
    n1029_lo_buf_o2
  );


  not

  (
    n1029_lo_buf_o2_n,
    n1029_lo_buf_o2
  );


  buf

  (
    n1041_lo_buf_o2_p,
    n1041_lo_buf_o2
  );


  not

  (
    n1041_lo_buf_o2_n,
    n1041_lo_buf_o2
  );


  buf

  (
    G558_o2_p,
    G558_o2
  );


  not

  (
    G558_o2_n,
    G558_o2
  );


  buf

  (
    G562_o2_p,
    G562_o2
  );


  not

  (
    G562_o2_n,
    G562_o2
  );


  buf

  (
    G566_o2_p,
    G566_o2
  );


  not

  (
    G566_o2_n,
    G566_o2
  );


  buf

  (
    n1835_o2_p,
    n1835_o2
  );


  not

  (
    n1835_o2_n,
    n1835_o2
  );


  buf

  (
    n1836_o2_p,
    n1836_o2
  );


  not

  (
    n1836_o2_n,
    n1836_o2
  );


  buf

  (
    n1837_o2_p,
    n1837_o2
  );


  not

  (
    n1837_o2_n,
    n1837_o2
  );


  buf

  (
    n765_lo_buf_o2_p,
    n765_lo_buf_o2
  );


  not

  (
    n765_lo_buf_o2_n,
    n765_lo_buf_o2
  );


  buf

  (
    n777_lo_buf_o2_p,
    n777_lo_buf_o2
  );


  not

  (
    n777_lo_buf_o2_n,
    n777_lo_buf_o2
  );


  buf

  (
    n789_lo_buf_o2_p,
    n789_lo_buf_o2
  );


  not

  (
    n789_lo_buf_o2_n,
    n789_lo_buf_o2
  );


  buf

  (
    G617_o2_p,
    G617_o2
  );


  not

  (
    G617_o2_n,
    G617_o2
  );


  buf

  (
    G626_o2_p,
    G626_o2
  );


  not

  (
    G626_o2_n,
    G626_o2
  );


  buf

  (
    G636_o2_p,
    G636_o2
  );


  not

  (
    G636_o2_n,
    G636_o2
  );


  buf

  (
    n489_lo_buf_o2_p,
    n489_lo_buf_o2
  );


  not

  (
    n489_lo_buf_o2_n,
    n489_lo_buf_o2
  );


  buf

  (
    n513_lo_buf_o2_p,
    n513_lo_buf_o2
  );


  not

  (
    n513_lo_buf_o2_n,
    n513_lo_buf_o2
  );


  buf

  (
    n561_lo_buf_o2_p,
    n561_lo_buf_o2
  );


  not

  (
    n561_lo_buf_o2_n,
    n561_lo_buf_o2
  );


  buf

  (
    n597_lo_buf_o2_p,
    n597_lo_buf_o2
  );


  not

  (
    n597_lo_buf_o2_n,
    n597_lo_buf_o2
  );


  buf

  (
    n657_lo_buf_o2_p,
    n657_lo_buf_o2
  );


  not

  (
    n657_lo_buf_o2_n,
    n657_lo_buf_o2
  );


  buf

  (
    G276_o2_p,
    G276_o2
  );


  not

  (
    G276_o2_n,
    G276_o2
  );


  buf

  (
    n1005_lo_buf_o2_p,
    n1005_lo_buf_o2
  );


  not

  (
    n1005_lo_buf_o2_n,
    n1005_lo_buf_o2
  );


  buf

  (
    n1161_lo_buf_o2_p,
    n1161_lo_buf_o2
  );


  not

  (
    n1161_lo_buf_o2_n,
    n1161_lo_buf_o2
  );


  buf

  (
    G620_o2_p,
    G620_o2
  );


  not

  (
    G620_o2_n,
    G620_o2
  );


  buf

  (
    G629_o2_p,
    G629_o2
  );


  not

  (
    G629_o2_n,
    G629_o2
  );


  buf

  (
    G639_o2_p,
    G639_o2
  );


  not

  (
    G639_o2_n,
    G639_o2
  );


  buf

  (
    G554_o2_p,
    G554_o2
  );


  not

  (
    G554_o2_n,
    G554_o2
  );


  buf

  (
    G690_o2_p,
    G690_o2
  );


  not

  (
    G690_o2_n,
    G690_o2
  );


  buf

  (
    G698_o2_p,
    G698_o2
  );


  not

  (
    G698_o2_n,
    G698_o2
  );


  buf

  (
    G707_o2_p,
    G707_o2
  );


  not

  (
    G707_o2_n,
    G707_o2
  );


  buf

  (
    G319_o2_p,
    G319_o2
  );


  not

  (
    G319_o2_n,
    G319_o2
  );


  buf

  (
    G389_o2_p,
    G389_o2
  );


  not

  (
    G389_o2_n,
    G389_o2
  );


  buf

  (
    n753_lo_buf_o2_p,
    n753_lo_buf_o2
  );


  not

  (
    n753_lo_buf_o2_n,
    n753_lo_buf_o2
  );


  buf

  (
    G647_o2_p,
    G647_o2
  );


  not

  (
    G647_o2_n,
    G647_o2
  );


  buf

  (
    G769_o2_p,
    G769_o2
  );


  not

  (
    G769_o2_n,
    G769_o2
  );


  buf

  (
    G785_o2_p,
    G785_o2
  );


  not

  (
    G785_o2_n,
    G785_o2
  );


  buf

  (
    G808_o2_p,
    G808_o2
  );


  not

  (
    G808_o2_n,
    G808_o2
  );


  buf

  (
    G445_o2_p,
    G445_o2
  );


  not

  (
    G445_o2_n,
    G445_o2
  );


  buf

  (
    G448_o2_p,
    G448_o2
  );


  not

  (
    G448_o2_n,
    G448_o2
  );


  buf

  (
    G477_o2_p,
    G477_o2
  );


  not

  (
    G477_o2_n,
    G477_o2
  );


  buf

  (
    G480_o2_p,
    G480_o2
  );


  not

  (
    G480_o2_n,
    G480_o2
  );


  buf

  (
    G436_o2_p,
    G436_o2
  );


  not

  (
    G436_o2_n,
    G436_o2
  );


  buf

  (
    G786_o2_p,
    G786_o2
  );


  not

  (
    G786_o2_n,
    G786_o2
  );


  buf

  (
    G787_o2_p,
    G787_o2
  );


  not

  (
    G787_o2_n,
    G787_o2
  );


  buf

  (
    G826_o2_p,
    G826_o2
  );


  not

  (
    G826_o2_n,
    G826_o2
  );


  buf

  (
    G827_o2_p,
    G827_o2
  );


  not

  (
    G827_o2_n,
    G827_o2
  );


  buf

  (
    G825_o2_p,
    G825_o2
  );


  not

  (
    G825_o2_n,
    G825_o2
  );


  buf

  (
    G610_o2_p,
    G610_o2
  );


  not

  (
    G610_o2_n,
    G610_o2
  );


  buf

  (
    n537_lo_buf_o2_p,
    n537_lo_buf_o2
  );


  not

  (
    n537_lo_buf_o2_n,
    n537_lo_buf_o2
  );


  buf

  (
    n669_lo_buf_o2_p,
    n669_lo_buf_o2
  );


  not

  (
    n669_lo_buf_o2_n,
    n669_lo_buf_o2
  );


  buf

  (
    n969_lo_buf_o2_p,
    n969_lo_buf_o2
  );


  not

  (
    n969_lo_buf_o2_n,
    n969_lo_buf_o2
  );


  buf

  (
    n981_lo_buf_o2_p,
    n981_lo_buf_o2
  );


  not

  (
    n981_lo_buf_o2_n,
    n981_lo_buf_o2
  );


  buf

  (
    n993_lo_buf_o2_p,
    n993_lo_buf_o2
  );


  not

  (
    n993_lo_buf_o2_n,
    n993_lo_buf_o2
  );


  buf

  (
    G309_o2_p,
    G309_o2
  );


  not

  (
    G309_o2_n,
    G309_o2
  );


  buf

  (
    G461_o2_p,
    G461_o2
  );


  not

  (
    G461_o2_n,
    G461_o2
  );


  buf

  (
    G487_o2_p,
    G487_o2
  );


  not

  (
    G487_o2_n,
    G487_o2
  );


  buf

  (
    G460_o2_p,
    G460_o2
  );


  not

  (
    G460_o2_n,
    G460_o2
  );


  buf

  (
    G468_o2_p,
    G468_o2
  );


  not

  (
    G468_o2_n,
    G468_o2
  );


  buf

  (
    G287_o2_p,
    G287_o2
  );


  not

  (
    G287_o2_n,
    G287_o2
  );


  buf

  (
    G613_o2_p,
    G613_o2
  );


  not

  (
    G613_o2_n,
    G613_o2
  );


  buf

  (
    n585_lo_buf_o2_p,
    n585_lo_buf_o2
  );


  not

  (
    n585_lo_buf_o2_n,
    n585_lo_buf_o2
  );


  buf

  (
    n813_lo_buf_o2_p,
    n813_lo_buf_o2
  );


  not

  (
    n813_lo_buf_o2_n,
    n813_lo_buf_o2
  );


  buf

  (
    n825_lo_buf_o2_p,
    n825_lo_buf_o2
  );


  not

  (
    n825_lo_buf_o2_n,
    n825_lo_buf_o2
  );


  buf

  (
    n837_lo_buf_o2_p,
    n837_lo_buf_o2
  );


  not

  (
    n837_lo_buf_o2_n,
    n837_lo_buf_o2
  );


  buf

  (
    n897_lo_buf_o2_p,
    n897_lo_buf_o2
  );


  not

  (
    n897_lo_buf_o2_n,
    n897_lo_buf_o2
  );


  buf

  (
    n909_lo_buf_o2_p,
    n909_lo_buf_o2
  );


  not

  (
    n909_lo_buf_o2_n,
    n909_lo_buf_o2
  );


  buf

  (
    n933_lo_buf_o2_p,
    n933_lo_buf_o2
  );


  not

  (
    n933_lo_buf_o2_n,
    n933_lo_buf_o2
  );


  buf

  (
    G451_o2_p,
    G451_o2
  );


  not

  (
    G451_o2_n,
    G451_o2
  );


  buf

  (
    G682_o2_p,
    G682_o2
  );


  not

  (
    G682_o2_n,
    G682_o2
  );


  buf

  (
    G756_o2_p,
    G756_o2
  );


  not

  (
    G756_o2_n,
    G756_o2
  );


  buf

  (
    G542_o2_p,
    G542_o2
  );


  not

  (
    G542_o2_n,
    G542_o2
  );


  buf

  (
    G546_o2_p,
    G546_o2
  );


  not

  (
    G546_o2_n,
    G546_o2
  );


  buf

  (
    G550_o2_p,
    G550_o2
  );


  not

  (
    G550_o2_n,
    G550_o2
  );


  buf

  (
    G310_o2_p,
    G310_o2
  );


  not

  (
    G310_o2_n,
    G310_o2
  );


  buf

  (
    n798_lo_buf_o2_p,
    n798_lo_buf_o2
  );


  not

  (
    n798_lo_buf_o2_n,
    n798_lo_buf_o2
  );


  buf

  (
    n882_lo_buf_o2_p,
    n882_lo_buf_o2
  );


  not

  (
    n882_lo_buf_o2_n,
    n882_lo_buf_o2
  );


  buf

  (
    G427_o2_p,
    G427_o2
  );


  not

  (
    G427_o2_n,
    G427_o2
  );


  buf

  (
    G497_o2_p,
    G497_o2
  );


  not

  (
    G497_o2_n,
    G497_o2
  );


  buf

  (
    G499_o2_p,
    G499_o2
  );


  not

  (
    G499_o2_n,
    G499_o2
  );


  buf

  (
    G501_o2_p,
    G501_o2
  );


  not

  (
    G501_o2_n,
    G501_o2
  );


  buf

  (
    G498_o2_p,
    G498_o2
  );


  not

  (
    G498_o2_n,
    G498_o2
  );


  buf

  (
    G500_o2_p,
    G500_o2
  );


  not

  (
    G500_o2_n,
    G500_o2
  );


  buf

  (
    G502_o2_p,
    G502_o2
  );


  not

  (
    G502_o2_n,
    G502_o2
  );


  buf

  (
    G369_o2_p,
    G369_o2
  );


  not

  (
    G369_o2_n,
    G369_o2
  );


  buf

  (
    n939_lo_buf_o2_p,
    n939_lo_buf_o2
  );


  not

  (
    n939_lo_buf_o2_n,
    n939_lo_buf_o2
  );


  buf

  (
    n486_lo_buf_o2_p,
    n486_lo_buf_o2
  );


  not

  (
    n486_lo_buf_o2_n,
    n486_lo_buf_o2
  );


  buf

  (
    n510_lo_buf_o2_p,
    n510_lo_buf_o2
  );


  not

  (
    n510_lo_buf_o2_n,
    n510_lo_buf_o2
  );


  buf

  (
    n558_lo_buf_o2_p,
    n558_lo_buf_o2
  );


  not

  (
    n558_lo_buf_o2_n,
    n558_lo_buf_o2
  );


  buf

  (
    n594_lo_buf_o2_p,
    n594_lo_buf_o2
  );


  not

  (
    n594_lo_buf_o2_n,
    n594_lo_buf_o2
  );


  buf

  (
    n654_lo_buf_o2_p,
    n654_lo_buf_o2
  );


  not

  (
    n654_lo_buf_o2_n,
    n654_lo_buf_o2
  );


  buf

  (
    n477_lo_buf_o2_p,
    n477_lo_buf_o2
  );


  not

  (
    n477_lo_buf_o2_n,
    n477_lo_buf_o2
  );


  buf

  (
    n525_lo_buf_o2_p,
    n525_lo_buf_o2
  );


  not

  (
    n525_lo_buf_o2_n,
    n525_lo_buf_o2
  );


  buf

  (
    n573_lo_buf_o2_p,
    n573_lo_buf_o2
  );


  not

  (
    n573_lo_buf_o2_n,
    n573_lo_buf_o2
  );


  or

  (
    g359_n,
    n660_lo_n,
    n540_lo_n_spl_0
  );


  or

  (
    g360_n,
    g359_n,
    n564_lo_n_spl_0
  );


  or

  (
    g361_n,
    n552_lo_n_spl_,
    n540_lo_n_spl_0
  );


  or

  (
    g362_n,
    g361_n_spl_,
    n672_lo_n_spl_
  );


  or

  (
    g363_n,
    g361_n_spl_,
    n564_lo_n_spl_0
  );


  or

  (
    g364_n,
    n696_lo_n,
    n684_lo_n
  );


  or

  (
    g365_n,
    n492_lo_n,
    n480_lo_n_spl_
  );


  or

  (
    g366_n,
    g365_n,
    n504_lo_n_spl_
  );


  or

  (
    g367_n,
    g366_n,
    n516_lo_n_spl_
  );


  and

  (
    g368_p,
    n528_lo_p,
    n480_lo_p
  );


  or

  (
    g368_n,
    n528_lo_n,
    n480_lo_n_spl_
  );


  and

  (
    g369_p,
    g368_p,
    n504_lo_p
  );


  or

  (
    g369_n,
    g368_n,
    n504_lo_n_spl_
  );


  and

  (
    g370_p,
    g369_p,
    n516_lo_p
  );


  or

  (
    g370_n,
    g369_n,
    n516_lo_n_spl_
  );


  and

  (
    g371_p,
    g370_p,
    g363_n_spl_0
  );


  and

  (
    g372_p,
    n660_lo_p,
    n600_lo_p
  );


  and

  (
    g373_p,
    g372_p,
    n672_lo_p
  );


  or

  (
    g374_n,
    n600_lo_n_spl_,
    n552_lo_n_spl_
  );


  or

  (
    g375_n,
    g374_n_spl_,
    n672_lo_n_spl_
  );


  or

  (
    g376_n,
    g374_n_spl_,
    n564_lo_n_spl_
  );


  or

  (
    g377_n,
    n720_lo_p,
    n708_lo_p
  );


  and

  (
    g378_p,
    g377_n_spl_,
    n744_lo_p
  );


  or

  (
    g379_n,
    g370_n,
    g363_n_spl_0
  );


  or

  (
    g380_n,
    n612_lo_n_spl_,
    n540_lo_n_spl_
  );


  or

  (
    g381_n,
    g380_n,
    G280_o2_n_spl_
  );


  or

  (
    g382_n,
    n612_lo_n_spl_,
    n600_lo_n_spl_
  );


  or

  (
    g383_n,
    g382_n,
    n648_lo_n
  );


  or

  (
    g384_n,
    g383_n,
    G280_o2_n_spl_
  );


  and

  (
    g385_p,
    g377_n_spl_,
    n732_lo_p
  );


  and

  (
    g386_p,
    G445_o2_p_spl_,
    n852_lo_p_spl_0
  );


  or

  (
    g386_n,
    G445_o2_n_spl_,
    n852_lo_n_spl_0
  );


  and

  (
    g387_p,
    G445_o2_n_spl_,
    n852_lo_n_spl_0
  );


  or

  (
    g387_n,
    G445_o2_p_spl_,
    n852_lo_p_spl_0
  );


  and

  (
    g388_p,
    g387_n,
    g386_n
  );


  or

  (
    g388_n,
    g387_p,
    g386_p
  );


  and

  (
    g389_p,
    G448_o2_p_spl_,
    n864_lo_p_spl_
  );


  or

  (
    g389_n,
    G448_o2_n_spl_,
    n864_lo_n_spl_
  );


  and

  (
    g390_p,
    G448_o2_n_spl_,
    n864_lo_n_spl_
  );


  or

  (
    g390_n,
    G448_o2_p_spl_,
    n864_lo_p_spl_
  );


  and

  (
    g391_p,
    g390_n,
    g389_n
  );


  or

  (
    g391_n,
    g390_p,
    g389_p
  );


  and

  (
    g392_p,
    g391_n,
    g388_n
  );


  and

  (
    g393_p,
    g391_p,
    g388_p
  );


  or

  (
    g394_n,
    g393_p,
    g392_p
  );


  and

  (
    g395_p,
    G477_o2_p_spl_,
    n852_lo_p_spl_1
  );


  or

  (
    g395_n,
    G477_o2_n_spl_,
    n852_lo_n_spl_1
  );


  and

  (
    g396_p,
    G477_o2_n_spl_,
    n852_lo_n_spl_1
  );


  or

  (
    g396_n,
    G477_o2_p_spl_,
    n852_lo_p_spl_1
  );


  and

  (
    g397_p,
    g396_n,
    g395_n
  );


  or

  (
    g397_n,
    g396_p,
    g395_p
  );


  and

  (
    g398_p,
    G480_o2_p_spl_,
    n1056_lo_p_spl_
  );


  or

  (
    g398_n,
    G480_o2_n_spl_,
    n1056_lo_n_spl_
  );


  and

  (
    g399_p,
    G480_o2_n_spl_,
    n1056_lo_n_spl_
  );


  or

  (
    g399_n,
    G480_o2_p_spl_,
    n1056_lo_p_spl_
  );


  and

  (
    g400_p,
    g399_n,
    g398_n
  );


  or

  (
    g400_n,
    g399_p,
    g398_p
  );


  and

  (
    g401_p,
    g400_n,
    g397_n
  );


  and

  (
    g402_p,
    g400_p,
    g397_p
  );


  or

  (
    g403_n,
    g402_p,
    g401_p
  );


  or

  (
    g404_n,
    n1068_lo_n_spl_00,
    n828_lo_n
  );


  or

  (
    g405_n,
    G769_o2_n,
    n1080_lo_n_spl_00
  );


  and

  (
    g406_p,
    g405_n,
    g404_n
  );


  or

  (
    g407_n,
    G712_o2_n,
    n1092_lo_n_spl_00
  );


  or

  (
    g408_n,
    n1732_o2_n,
    n1104_lo_n_spl_00
  );


  and

  (
    g409_p,
    g408_n,
    g407_n
  );


  or

  (
    g410_n,
    n1176_lo_n,
    n1128_lo_n_spl_0
  );


  or

  (
    g411_n,
    n1657_o2_n,
    n1116_lo_n_spl_00
  );


  and

  (
    g412_p,
    g411_n,
    g410_n
  );


  or

  (
    g413_n,
    G436_o2_n_spl_00,
    n1044_lo_n
  );


  and

  (
    g414_p,
    g409_p,
    g406_p
  );


  and

  (
    g415_p,
    g414_p,
    g412_p
  );


  and

  (
    g416_p,
    g415_p,
    g413_n
  );


  or

  (
    g417_n,
    n1068_lo_n_spl_00,
    n792_lo_n
  );


  or

  (
    g418_n,
    G785_o2_n,
    n1080_lo_n_spl_00
  );


  and

  (
    g419_p,
    g418_n,
    g417_n
  );


  or

  (
    g420_n,
    G685_o2_n,
    n1092_lo_n_spl_00
  );


  or

  (
    g421_n,
    n1805_o2_n,
    n1104_lo_n_spl_00
  );


  and

  (
    g422_p,
    g421_n,
    g420_n
  );


  or

  (
    g423_n,
    n1729_o2_n,
    n1116_lo_n_spl_00
  );


  or

  (
    g424_n,
    G436_o2_n_spl_00,
    n1008_lo_n
  );


  and

  (
    g425_p,
    g424_n,
    g423_n
  );


  and

  (
    g426_p,
    g422_p,
    g419_p
  );


  and

  (
    g427_p,
    g426_p,
    g425_p
  );


  or

  (
    g428_n,
    n1068_lo_n_spl_01,
    n804_lo_n
  );


  or

  (
    g429_n,
    G786_o2_n,
    n1080_lo_n_spl_01
  );


  and

  (
    g430_p,
    g429_n,
    g428_n
  );


  or

  (
    g431_n,
    G693_o2_n,
    n1092_lo_n_spl_01
  );


  or

  (
    g432_n,
    n1730_o2_n,
    n1104_lo_n_spl_01
  );


  and

  (
    g433_p,
    g432_n,
    g431_n
  );


  or

  (
    g434_n,
    n1140_lo_n,
    n1128_lo_n_spl_0
  );


  or

  (
    g435_n,
    n1655_o2_n,
    n1116_lo_n_spl_01
  );


  and

  (
    g436_p,
    g435_n,
    g434_n
  );


  or

  (
    g437_n,
    G436_o2_n_spl_01,
    n1020_lo_n
  );


  and

  (
    g438_p,
    g433_p,
    g430_p
  );


  and

  (
    g439_p,
    g438_p,
    g436_p
  );


  and

  (
    g440_p,
    g439_p,
    g437_n
  );


  or

  (
    g441_n,
    n1068_lo_n_spl_01,
    n816_lo_n
  );


  or

  (
    g442_n,
    G787_o2_n,
    n1080_lo_n_spl_01
  );


  and

  (
    g443_p,
    g442_n,
    g441_n
  );


  or

  (
    g444_n,
    G702_o2_n,
    n1092_lo_n_spl_01
  );


  or

  (
    g445_n,
    n1731_o2_n,
    n1104_lo_n_spl_01
  );


  and

  (
    g446_p,
    g445_n,
    g444_n
  );


  or

  (
    g447_n,
    n1152_lo_n,
    n1128_lo_n_spl_
  );


  or

  (
    g448_n,
    n1656_o2_n,
    n1116_lo_n_spl_01
  );


  and

  (
    g449_p,
    g448_n,
    g447_n
  );


  or

  (
    g450_n,
    G436_o2_n_spl_01,
    n1032_lo_n
  );


  and

  (
    g451_p,
    g446_p,
    g443_p
  );


  and

  (
    g452_p,
    g451_p,
    g449_p
  );


  and

  (
    g453_p,
    g452_p,
    g450_n
  );


  or

  (
    g454_n,
    G798_o2_n,
    G578_o2_n
  );


  and

  (
    g455_p,
    g454_n,
    G647_o2_n_spl_
  );


  or

  (
    g456_n,
    n1068_lo_n_spl_10,
    n780_lo_n
  );


  or

  (
    g457_n,
    G808_o2_n,
    n1080_lo_n_spl_10
  );


  and

  (
    g458_p,
    g457_n,
    g456_n
  );


  or

  (
    g459_n,
    G677_o2_n,
    n1092_lo_n_spl_10
  );


  or

  (
    g460_n,
    G672_o2_n,
    n1104_lo_n_spl_10
  );


  and

  (
    g461_p,
    g460_n,
    g459_n
  );


  or

  (
    g462_n,
    n1809_o2_n,
    n1116_lo_n_spl_10
  );


  or

  (
    g463_n,
    G436_o2_n_spl_10,
    n996_lo_n
  );


  and

  (
    g464_p,
    g463_n,
    g462_n
  );


  and

  (
    g465_p,
    g461_p,
    g458_p
  );


  and

  (
    g466_p,
    g465_p,
    g464_p
  );


  or

  (
    g467_n,
    n1616_o2_n,
    n1068_lo_n_spl_10
  );


  or

  (
    g468_n,
    G825_o2_n,
    n1080_lo_n_spl_10
  );


  and

  (
    g469_p,
    g468_n,
    g467_n
  );


  or

  (
    g470_n,
    G650_o2_n,
    n1092_lo_n_spl_10
  );


  or

  (
    g471_n,
    G647_o2_n_spl_,
    n1104_lo_n_spl_10
  );


  and

  (
    g472_p,
    g471_n,
    g470_n
  );


  or

  (
    g473_n,
    G538_o2_n,
    n1116_lo_n_spl_10
  );


  or

  (
    g474_n,
    G436_o2_n_spl_10,
    n960_lo_n
  );


  and

  (
    g475_p,
    g474_n,
    g473_n
  );


  and

  (
    g476_p,
    g472_p,
    g469_p
  );


  and

  (
    g477_p,
    g476_p,
    g475_p
  );


  or

  (
    g478_n,
    n1068_lo_n_spl_11,
    n756_lo_n
  );


  or

  (
    g479_n,
    G826_o2_n,
    n1080_lo_n_spl_11
  );


  and

  (
    g480_p,
    g479_n,
    g478_n
  );


  or

  (
    g481_n,
    G658_o2_n,
    n1092_lo_n_spl_11
  );


  or

  (
    g482_n,
    G655_o2_n,
    n1104_lo_n_spl_11
  );


  and

  (
    g483_p,
    g482_n,
    g481_n
  );


  or

  (
    g484_n,
    n1807_o2_n,
    n1116_lo_n_spl_11
  );


  or

  (
    g485_n,
    G436_o2_n_spl_11,
    n972_lo_n
  );


  and

  (
    g486_p,
    g485_n,
    g484_n
  );


  and

  (
    g487_p,
    g483_p,
    g480_p
  );


  and

  (
    g488_p,
    g487_p,
    g486_p
  );


  or

  (
    g489_n,
    n1068_lo_n_spl_11,
    n768_lo_n
  );


  or

  (
    g490_n,
    G827_o2_n,
    n1080_lo_n_spl_11
  );


  and

  (
    g491_p,
    g490_n,
    g489_n
  );


  or

  (
    g492_n,
    G667_o2_n,
    n1092_lo_n_spl_11
  );


  or

  (
    g493_n,
    G663_o2_n,
    n1104_lo_n_spl_11
  );


  and

  (
    g494_p,
    g493_n,
    g492_n
  );


  or

  (
    g495_n,
    n1808_o2_n,
    n1116_lo_n_spl_11
  );


  or

  (
    g496_n,
    G436_o2_n_spl_11,
    n984_lo_n
  );


  and

  (
    g497_p,
    g496_n,
    g495_n
  );


  and

  (
    g498_p,
    g494_p,
    g491_p
  );


  and

  (
    g499_p,
    g498_p,
    g497_p
  );


  or

  (
    g500_n,
    n1704_o2_n,
    n1663_o2_n
  );


  or

  (
    g501_n,
    g500_n,
    n501_lo_n
  );


  or

  (
    g502_n,
    g501_n,
    n1797_o2_n
  );


  and

  (
    g503_p,
    G542_o2_p_spl_0,
    n969_lo_buf_o2_p_spl_00
  );


  or

  (
    g503_n,
    G542_o2_n_spl_,
    n969_lo_buf_o2_n_spl_0
  );


  and

  (
    g504_p,
    G546_o2_p_spl_0,
    n981_lo_buf_o2_p_spl_00
  );


  or

  (
    g504_n,
    G546_o2_n_spl_,
    n981_lo_buf_o2_n_spl_0
  );


  and

  (
    g505_p,
    G550_o2_p_spl_0,
    n993_lo_buf_o2_p_spl_00
  );


  or

  (
    g505_n,
    G550_o2_n_spl_,
    n993_lo_buf_o2_n_spl_0
  );


  and

  (
    g506_p,
    G487_o2_n,
    G309_o2_n
  );


  or

  (
    g506_n,
    G487_o2_p,
    G309_o2_p
  );


  and

  (
    g507_p,
    G460_o2_n,
    G461_o2_n
  );


  or

  (
    g507_n,
    G460_o2_p,
    G461_o2_p
  );


  and

  (
    g508_p,
    g507_p,
    g506_p
  );


  or

  (
    g508_n,
    g507_n,
    g506_n
  );


  and

  (
    g509_p,
    g508_p_spl_,
    n957_lo_n_spl_0
  );


  or

  (
    g509_n,
    g508_n_spl_0,
    n957_lo_p_spl_00
  );


  and

  (
    g510_p,
    G620_o2_p,
    G617_o2_n
  );


  or

  (
    g510_n,
    G620_o2_n,
    G617_o2_p
  );


  and

  (
    g511_p,
    G629_o2_p_spl_0,
    G626_o2_n
  );


  or

  (
    g511_n,
    G629_o2_n_spl_0,
    G626_o2_p
  );


  and

  (
    g512_p,
    G639_o2_p_spl_0,
    G636_o2_n
  );


  or

  (
    g512_n,
    G639_o2_n_spl_0,
    G636_o2_p
  );


  and

  (
    g513_p,
    G613_o2_p_spl_,
    G610_o2_n
  );


  or

  (
    g513_n,
    G613_o2_n_spl_,
    G610_o2_p
  );


  and

  (
    g514_p,
    G542_o2_n_spl_,
    n969_lo_buf_o2_n_spl_0
  );


  or

  (
    g514_n,
    G542_o2_p_spl_0,
    n969_lo_buf_o2_p_spl_00
  );


  and

  (
    g515_p,
    g514_n_spl_0,
    g503_n_spl_
  );


  or

  (
    g515_n,
    g514_p_spl_0,
    g503_p_spl_0
  );


  and

  (
    g516_p,
    G546_o2_n_spl_,
    n981_lo_buf_o2_n_spl_0
  );


  or

  (
    g516_n,
    G546_o2_p_spl_0,
    n981_lo_buf_o2_p_spl_00
  );


  and

  (
    g517_p,
    g516_n_spl_0,
    g504_n_spl_0
  );


  or

  (
    g517_n,
    g516_p_spl_0,
    g504_p_spl_0
  );


  and

  (
    g518_p,
    G550_o2_n_spl_,
    n993_lo_buf_o2_n_spl_0
  );


  or

  (
    g518_n,
    G550_o2_p_spl_0,
    n993_lo_buf_o2_p_spl_00
  );


  and

  (
    g519_p,
    g518_n_spl_0,
    g505_n_spl_0
  );


  or

  (
    g519_n,
    g518_p_spl_0,
    g505_p_spl_00
  );


  and

  (
    g520_p,
    g508_n_spl_0,
    n957_lo_p_spl_00
  );


  or

  (
    g520_n,
    g508_p_spl_,
    n957_lo_n_spl_0
  );


  and

  (
    g521_p,
    g520_n,
    g509_n_spl_
  );


  or

  (
    g521_n,
    g520_p_spl_,
    g509_p
  );


  and

  (
    g522_p,
    g514_n_spl_0,
    g504_p_spl_0
  );


  or

  (
    g522_n,
    g514_p_spl_0,
    g504_n_spl_0
  );


  and

  (
    g523_p,
    g516_n_spl_0,
    g514_n_spl_
  );


  or

  (
    g523_n,
    g516_p_spl_0,
    g514_p_spl_
  );


  and

  (
    g524_p,
    g523_p_spl_,
    g505_p_spl_00
  );


  or

  (
    g524_n,
    g523_n_spl_,
    g505_n_spl_0
  );


  and

  (
    g525_p,
    G756_o2_p_spl_,
    G613_o2_p_spl_
  );


  or

  (
    g525_n,
    G756_o2_n_spl_,
    G613_o2_n_spl_
  );


  and

  (
    g526_p,
    g525_n,
    G682_o2_n
  );


  or

  (
    g526_n,
    g525_p,
    G682_o2_p_spl_
  );


  and

  (
    g527_p,
    g523_p_spl_,
    g518_n_spl_0
  );


  or

  (
    g527_n,
    g523_n_spl_,
    g518_p_spl_0
  );


  and

  (
    g528_p,
    g527_p,
    g526_n_spl_0
  );


  or

  (
    g528_n,
    g527_n,
    g526_p_spl_0
  );


  and

  (
    g529_p,
    g522_n,
    g503_n_spl_
  );


  or

  (
    g529_n,
    g522_p,
    g503_p_spl_0
  );


  and

  (
    g530_p,
    g529_p,
    g524_n
  );


  or

  (
    g530_n,
    g529_n,
    g524_p
  );


  and

  (
    g531_p,
    g530_p,
    g528_n
  );


  or

  (
    g531_n,
    g530_n,
    g528_p
  );


  or

  (
    g532_n,
    G369_o2_p_spl_,
    G427_o2_n
  );


  and

  (
    g533_p,
    G498_o2_n,
    G497_o2_n
  );


  and

  (
    g534_p,
    g533_p,
    g532_n_spl_0
  );


  and

  (
    g535_p,
    G500_o2_n,
    G499_o2_n
  );


  and

  (
    g536_p,
    g535_p,
    g532_n_spl_0
  );


  and

  (
    g537_p,
    G502_o2_n,
    G501_o2_n
  );


  and

  (
    g538_p,
    g537_p,
    g532_n_spl_1
  );


  or

  (
    g539_n,
    g534_p_spl_0,
    n1014_lo_n_spl_
  );


  or

  (
    g540_n,
    g536_p_spl_0,
    n1026_lo_n_spl_
  );


  or

  (
    g541_n,
    g538_p_spl_0,
    n1038_lo_n_spl_
  );


  and

  (
    g542_p,
    n525_lo_buf_o2_p_spl_,
    n477_lo_buf_o2_p_spl_0
  );


  or

  (
    g542_n,
    n525_lo_buf_o2_n,
    n477_lo_buf_o2_n_spl_
  );


  and

  (
    g543_p,
    g542_p,
    n573_lo_buf_o2_p_spl_0
  );


  or

  (
    g543_n,
    g542_n,
    n573_lo_buf_o2_n
  );


  and

  (
    g544_p,
    g534_p_spl_0,
    n1014_lo_n_spl_
  );


  and

  (
    g545_p,
    g536_p_spl_0,
    n1026_lo_n_spl_
  );


  and

  (
    g546_p,
    g538_p_spl_0,
    n1038_lo_n_spl_
  );


  or

  (
    g547_n,
    n882_lo_buf_o2_n_spl_,
    G468_o2_p
  );


  or

  (
    g548_n,
    n798_lo_buf_o2_n,
    G451_o2_n_spl_0
  );


  and

  (
    g549_p,
    g548_n,
    g547_n
  );


  and

  (
    g550_p,
    g549_p,
    g532_n_spl_1
  );


  or

  (
    g551_n,
    n594_lo_buf_o2_n_spl_,
    n939_lo_buf_o2_n
  );


  or

  (
    g552_n,
    g512_p_spl_,
    n1161_lo_buf_o2_p_spl_0
  );


  or

  (
    g553_n,
    g512_n,
    n1161_lo_buf_o2_n_spl_0
  );


  and

  (
    g554_p,
    g553_n,
    g552_n
  );


  or

  (
    g555_n,
    g513_p_spl_,
    G756_o2_p_spl_
  );


  or

  (
    g556_n,
    g513_n,
    G756_o2_n_spl_
  );


  and

  (
    g557_p,
    g556_n,
    g555_n
  );


  or

  (
    g558_n,
    g526_n_spl_0,
    g519_p_spl_
  );


  or

  (
    g559_n,
    g526_p_spl_0,
    g519_n
  );


  and

  (
    g560_p,
    g559_n,
    g558_n
  );


  and

  (
    g561_p,
    n753_lo_buf_o2_p_spl_0,
    n765_lo_buf_o2_p_spl_0
  );


  or

  (
    g561_n,
    n753_lo_buf_o2_n_spl_,
    n765_lo_buf_o2_n_spl_
  );


  and

  (
    g562_p,
    n753_lo_buf_o2_n_spl_,
    n765_lo_buf_o2_n_spl_
  );


  or

  (
    g562_n,
    n753_lo_buf_o2_p_spl_0,
    n765_lo_buf_o2_p_spl_0
  );


  and

  (
    g563_p,
    g562_n,
    g561_n
  );


  or

  (
    g563_n,
    g562_p,
    g561_p
  );


  and

  (
    g564_p,
    n789_lo_buf_o2_p_spl_0,
    n777_lo_buf_o2_p_spl_0
  );


  or

  (
    g564_n,
    n789_lo_buf_o2_n_spl_,
    n777_lo_buf_o2_n_spl_
  );


  and

  (
    g565_p,
    n789_lo_buf_o2_n_spl_,
    n777_lo_buf_o2_n_spl_
  );


  or

  (
    g565_n,
    n789_lo_buf_o2_p_spl_0,
    n777_lo_buf_o2_p_spl_0
  );


  and

  (
    g566_p,
    g565_n,
    g564_n
  );


  or

  (
    g566_n,
    g565_p,
    g564_p
  );


  or

  (
    g567_n,
    g566_p,
    g563_p
  );


  or

  (
    g568_n,
    g566_n,
    g563_n
  );


  and

  (
    g569_p,
    g568_n,
    g567_n
  );


  and

  (
    g570_p,
    n801_lo_buf_o2_p_spl_0,
    n1798_o2_p_spl_0
  );


  or

  (
    g570_n,
    n801_lo_buf_o2_n_spl_,
    n1798_o2_n_spl_
  );


  and

  (
    g571_p,
    n801_lo_buf_o2_n_spl_,
    n1798_o2_n_spl_
  );


  or

  (
    g571_n,
    n801_lo_buf_o2_p_spl_0,
    n1798_o2_p_spl_0
  );


  and

  (
    g572_p,
    g571_n,
    g570_n
  );


  or

  (
    g572_n,
    g571_p,
    g570_p
  );


  and

  (
    g573_p,
    n1800_o2_p_spl_,
    n1799_o2_p_spl_0
  );


  or

  (
    g573_n,
    n1800_o2_n_spl_,
    n1799_o2_n_spl_
  );


  and

  (
    g574_p,
    n1800_o2_n_spl_,
    n1799_o2_n_spl_
  );


  or

  (
    g574_n,
    n1800_o2_p_spl_,
    n1799_o2_p_spl_0
  );


  and

  (
    g575_p,
    g574_n,
    g573_n
  );


  or

  (
    g575_n,
    g574_p,
    g573_p
  );


  or

  (
    g576_n,
    g575_p,
    g572_p
  );


  or

  (
    g577_n,
    g575_n,
    g572_n
  );


  and

  (
    g578_p,
    g577_n,
    g576_n
  );


  and

  (
    g579_p,
    n969_lo_buf_o2_p_spl_0,
    n957_lo_p_spl_0
  );


  or

  (
    g579_n,
    n969_lo_buf_o2_n_spl_1,
    n957_lo_n_spl_1
  );


  and

  (
    g580_p,
    n969_lo_buf_o2_n_spl_1,
    n957_lo_n_spl_1
  );


  or

  (
    g580_n,
    n969_lo_buf_o2_p_spl_1,
    n957_lo_p_spl_1
  );


  and

  (
    g581_p,
    g580_n,
    g579_n
  );


  or

  (
    g581_n,
    g580_p,
    g579_p
  );


  and

  (
    g582_p,
    n993_lo_buf_o2_p_spl_0,
    n981_lo_buf_o2_p_spl_0
  );


  or

  (
    g582_n,
    n993_lo_buf_o2_n_spl_1,
    n981_lo_buf_o2_n_spl_1
  );


  and

  (
    g583_p,
    n993_lo_buf_o2_n_spl_1,
    n981_lo_buf_o2_n_spl_1
  );


  or

  (
    g583_n,
    n993_lo_buf_o2_p_spl_1,
    n981_lo_buf_o2_p_spl_1
  );


  and

  (
    g584_p,
    g583_n,
    g582_n
  );


  or

  (
    g584_n,
    g583_p,
    g582_p
  );


  or

  (
    g585_n,
    g584_p,
    g581_p
  );


  or

  (
    g586_n,
    g584_n,
    g581_n
  );


  and

  (
    g587_p,
    g586_n,
    g585_n
  );


  and

  (
    g588_p,
    n1005_lo_buf_o2_p_spl_0,
    n1017_lo_buf_o2_p_spl_0
  );


  or

  (
    g588_n,
    n1005_lo_buf_o2_n_spl_,
    n1017_lo_buf_o2_n_spl_
  );


  and

  (
    g589_p,
    n1005_lo_buf_o2_n_spl_,
    n1017_lo_buf_o2_n_spl_
  );


  or

  (
    g589_n,
    n1005_lo_buf_o2_p_spl_0,
    n1017_lo_buf_o2_p_spl_0
  );


  and

  (
    g590_p,
    g589_n,
    g588_n
  );


  or

  (
    g590_n,
    g589_p,
    g588_p
  );


  and

  (
    g591_p,
    n1041_lo_buf_o2_p_spl_0,
    n1029_lo_buf_o2_p_spl_0
  );


  or

  (
    g591_n,
    n1041_lo_buf_o2_n_spl_,
    n1029_lo_buf_o2_n_spl_
  );


  and

  (
    g592_p,
    n1041_lo_buf_o2_n_spl_,
    n1029_lo_buf_o2_n_spl_
  );


  or

  (
    g592_n,
    n1041_lo_buf_o2_p_spl_0,
    n1029_lo_buf_o2_p_spl_0
  );


  and

  (
    g593_p,
    g592_n,
    g591_n
  );


  or

  (
    g593_n,
    g592_p,
    g591_p
  );


  or

  (
    g594_n,
    g593_p,
    g590_p
  );


  or

  (
    g595_n,
    g593_n,
    g590_n
  );


  and

  (
    g596_p,
    g595_n,
    g594_n
  );


  or

  (
    g597_n,
    n1707_o2_n,
    n1706_o2_n
  );


  or

  (
    g598_n,
    g597_n,
    n609_lo_n
  );


  or

  (
    g599_n,
    g598_n,
    n621_lo_n
  );


  or

  (
    g600_n,
    g599_n,
    g502_n_spl_
  );


  or

  (
    g601_n,
    g600_n,
    n633_lo_n
  );


  and

  (
    g602_p,
    G707_o2_p_spl_0,
    G629_o2_p_spl_0
  );


  or

  (
    g602_n,
    G707_o2_n_spl_,
    G629_o2_n_spl_0
  );


  and

  (
    g603_p,
    G639_o2_p_spl_0,
    G629_o2_p_spl_
  );


  or

  (
    g603_n,
    G639_o2_n_spl_0,
    G629_o2_n_spl_
  );


  and

  (
    g604_p,
    g603_p,
    n1161_lo_buf_o2_p_spl_0
  );


  or

  (
    g604_n,
    g603_n,
    n1161_lo_buf_o2_n_spl_0
  );


  and

  (
    g605_p,
    g602_n,
    G698_o2_n
  );


  or

  (
    g605_n,
    g602_p,
    G698_o2_p_spl_
  );


  and

  (
    g606_p,
    g605_p,
    g604_n
  );


  or

  (
    g606_n,
    g605_n,
    g604_p
  );


  or

  (
    g607_n,
    g606_n,
    g510_p_spl_
  );


  or

  (
    g608_n,
    g606_p,
    g510_n
  );


  and

  (
    g609_p,
    g608_n,
    g607_n
  );


  and

  (
    g610_p,
    G639_o2_p_spl_,
    n1161_lo_buf_o2_p_spl_
  );


  or

  (
    g610_n,
    G639_o2_n_spl_,
    n1161_lo_buf_o2_n_spl_
  );


  and

  (
    g611_p,
    g610_n,
    G707_o2_n_spl_
  );


  or

  (
    g611_n,
    g610_p,
    G707_o2_p_spl_0
  );


  or

  (
    g612_n,
    g611_n,
    g511_p_spl_
  );


  or

  (
    g613_n,
    g611_p,
    g511_n
  );


  and

  (
    g614_p,
    g613_n,
    g612_n
  );


  and

  (
    g615_p,
    g516_n_spl_1,
    g505_p_spl_0
  );


  or

  (
    g615_n,
    g516_p_spl_1,
    g505_n_spl_1
  );


  and

  (
    g616_p,
    g518_n_spl_1,
    g516_n_spl_1
  );


  or

  (
    g616_n,
    g518_p_spl_1,
    g516_p_spl_1
  );


  and

  (
    g617_p,
    g616_p,
    g526_n_spl_1
  );


  or

  (
    g617_n,
    g616_n,
    g526_p_spl_1
  );


  and

  (
    g618_p,
    g615_n,
    g504_n_spl_
  );


  or

  (
    g618_n,
    g615_p,
    g504_p_spl_1
  );


  and

  (
    g619_p,
    g618_p,
    g617_n
  );


  or

  (
    g619_n,
    g618_n,
    g617_p
  );


  or

  (
    g620_n,
    g619_n,
    g515_p_spl_
  );


  or

  (
    g621_n,
    g619_p,
    g515_n
  );


  and

  (
    g622_p,
    g621_n,
    g620_n
  );


  and

  (
    g623_p,
    g526_n_spl_1,
    g518_n_spl_1
  );


  or

  (
    g623_n,
    g526_p_spl_1,
    g518_p_spl_1
  );


  and

  (
    g624_p,
    g623_n,
    g505_n_spl_1
  );


  or

  (
    g624_n,
    g623_p,
    g505_p_spl_1
  );


  or

  (
    g625_n,
    g624_n,
    g517_p_spl_
  );


  or

  (
    g626_n,
    g624_p,
    g517_n
  );


  and

  (
    g627_p,
    g626_n,
    g625_n
  );


  or

  (
    g628_n,
    g531_n_spl_,
    g521_p_spl_
  );


  or

  (
    g629_n,
    g531_p,
    g521_n
  );


  and

  (
    g630_p,
    g629_n,
    g628_n
  );


  or

  (
    g631_n,
    g550_p_spl_0,
    n1002_lo_n_spl_
  );


  and

  (
    g632_p,
    n489_lo_buf_o2_p_spl_,
    n870_lo_p
  );


  or

  (
    g633_n,
    G389_o2_n_spl_,
    n513_lo_buf_o2_n_spl_
  );


  or

  (
    g634_n,
    g633_n,
    G287_o2_n
  );


  or

  (
    g635_n,
    g634_n,
    G310_o2_p
  );


  and

  (
    g636_p,
    G451_o2_p,
    n750_lo_p_spl_
  );


  or

  (
    g637_n,
    G389_o2_n_spl_,
    G319_o2_p
  );


  or

  (
    g638_n,
    g637_n,
    n585_lo_buf_o2_n
  );


  or

  (
    g639_n,
    g638_n_spl_0,
    n882_lo_buf_o2_n_spl_
  );


  and

  (
    g640_p,
    g551_n_spl_,
    g543_p_spl_0
  );


  and

  (
    g641_p,
    g640_p,
    n510_lo_buf_o2_p_spl_0
  );


  or

  (
    g642_n,
    g641_p,
    n477_lo_buf_o2_n_spl_
  );


  or

  (
    g643_n,
    n654_lo_buf_o2_n_spl_,
    n531_lo_n
  );


  or

  (
    g644_n,
    g643_n,
    n663_lo_n
  );


  and

  (
    g645_p,
    g550_p_spl_0,
    n1002_lo_n_spl_
  );


  or

  (
    g646_n,
    n558_lo_buf_o2_p_spl_,
    n510_lo_buf_o2_p_spl_0
  );


  or

  (
    g647_n,
    n558_lo_buf_o2_n_spl_,
    n510_lo_buf_o2_n
  );


  and

  (
    g648_p,
    g647_n,
    g646_n
  );


  and

  (
    g649_p,
    g648_p,
    n594_lo_buf_o2_p_spl_
  );


  and

  (
    g650_p,
    g649_p,
    n939_lo_buf_o2_p
  );


  and

  (
    g651_p,
    g650_p,
    g543_p_spl_0
  );


  and

  (
    g652_p,
    n477_lo_buf_o2_p_spl_0,
    n486_lo_buf_o2_p_spl_
  );


  and

  (
    g653_p,
    g652_p,
    n573_lo_buf_o2_p_spl_0
  );


  and

  (
    g654_p,
    g653_p,
    n510_lo_buf_o2_p_spl_1
  );


  or

  (
    g655_n,
    n654_lo_buf_o2_n_spl_,
    n594_lo_buf_o2_n_spl_
  );


  or

  (
    g656_n,
    g655_n,
    n558_lo_buf_o2_n_spl_
  );


  and

  (
    g657_p,
    g656_n,
    g654_p
  );


  or

  (
    g658_n,
    g657_p,
    g651_p
  );


  or

  (
    g659_n,
    g544_p_spl_0,
    g540_n_spl_0
  );


  or

  (
    g660_n,
    g545_p_spl_,
    g544_p_spl_0
  );


  or

  (
    g661_n,
    g660_n_spl_,
    g541_n_spl_0
  );


  or

  (
    g662_n,
    g660_n_spl_,
    g546_p_spl_
  );


  or

  (
    g663_n,
    g662_n,
    n1158_lo_n
  );


  and

  (
    g664_p,
    g659_n,
    g539_n_spl_0
  );


  and

  (
    g665_p,
    g664_p,
    g661_n
  );


  and

  (
    g666_p,
    g665_p,
    g663_n
  );


  or

  (
    g667_n,
    n1837_o2_n,
    n870_lo_n_spl_0
  );


  or

  (
    g668_n,
    G451_o2_n_spl_0,
    n762_lo_n
  );


  and

  (
    g669_p,
    g668_n,
    g667_n
  );


  or

  (
    g670_n,
    g638_n_spl_0,
    n897_lo_buf_o2_n
  );


  and

  (
    g671_p,
    g670_n,
    g635_n_spl_0
  );


  and

  (
    g672_p,
    g671_p,
    g669_p
  );


  or

  (
    g673_n,
    n513_lo_buf_o2_n_spl_,
    n870_lo_n_spl_0
  );


  or

  (
    g674_n,
    G451_o2_n_spl_1,
    n774_lo_n
  );


  and

  (
    g675_p,
    g674_n,
    g673_n
  );


  or

  (
    g676_n,
    g638_n_spl_1,
    n909_lo_buf_o2_n
  );


  and

  (
    g677_p,
    g676_n,
    g635_n_spl_0
  );


  and

  (
    g678_p,
    g677_p,
    g675_p
  );


  or

  (
    g679_n,
    n918_lo_n,
    n870_lo_n_spl_
  );


  or

  (
    g680_n,
    G451_o2_n_spl_1,
    n786_lo_n
  );


  and

  (
    g681_p,
    g680_n,
    g679_n
  );


  or

  (
    g682_n,
    g638_n_spl_1,
    n933_lo_buf_o2_n
  );


  and

  (
    g683_p,
    g682_n,
    g635_n_spl_1
  );


  and

  (
    g684_p,
    g683_p,
    g681_p
  );


  or

  (
    g685_n,
    g644_n_spl_,
    g543_n
  );


  or

  (
    g686_n,
    g685_n,
    n579_lo_n
  );


  and

  (
    g687_p,
    g642_n_spl_0,
    n891_lo_p_spl_
  );


  and

  (
    g688_p,
    g642_n_spl_0,
    n903_lo_p_spl_
  );


  and

  (
    g689_p,
    g642_n_spl_1,
    n927_lo_p_spl_
  );


  and

  (
    g690_p,
    g658_n_spl_0,
    n807_lo_p_spl_
  );


  and

  (
    g691_p,
    g658_n_spl_0,
    n819_lo_p_spl_
  );


  and

  (
    g692_p,
    g658_n_spl_1,
    n831_lo_p_spl_
  );


  buf

  (
    G855,
    g360_n
  );


  buf

  (
    G856,
    g362_n
  );


  buf

  (
    G857,
    g363_n_spl_
  );


  buf

  (
    G858,
    g364_n
  );


  buf

  (
    G859,
    g367_n
  );


  buf

  (
    G860,
    g371_p
  );


  buf

  (
    G861,
    g373_p
  );


  not

  (
    G862,
    g375_n
  );


  not

  (
    G863,
    g376_n
  );


  not

  (
    G864,
    g378_p
  );


  not

  (
    G865,
    g379_n
  );


  buf

  (
    G866,
    n1529_o2_n
  );


  buf

  (
    G867,
    g381_n
  );


  buf

  (
    G868,
    g384_n
  );


  not

  (
    G869,
    g385_p
  );


  buf

  (
    G870,
    g394_n
  );


  buf

  (
    G871,
    g403_n
  );


  buf

  (
    G872,
    g416_p
  );


  buf

  (
    G873,
    g427_p
  );


  buf

  (
    G874,
    g440_p
  );


  buf

  (
    G875,
    g453_p
  );


  buf

  (
    G876,
    g455_p
  );


  buf

  (
    G877,
    g466_p
  );


  buf

  (
    G878,
    g477_p
  );


  buf

  (
    G879,
    g488_p
  );


  buf

  (
    G880,
    g499_p
  );


  buf

  (
    n480_li,
    n1663_o2_p
  );


  buf

  (
    n492_li,
    n1704_o2_p
  );


  buf

  (
    n495_li,
    G3_p
  );


  buf

  (
    n498_li,
    n495_lo_p
  );


  buf

  (
    n501_li,
    n498_lo_p
  );


  buf

  (
    n504_li,
    n501_lo_p
  );


  buf

  (
    n516_li,
    n1705_o2_p
  );


  buf

  (
    n528_li,
    n1664_o2_p
  );


  buf

  (
    n531_li,
    G6_p
  );


  buf

  (
    n540_li,
    n1780_o2_p
  );


  buf

  (
    n543_li,
    G7_p
  );


  buf

  (
    n546_li,
    n543_lo_p
  );


  buf

  (
    n549_li,
    n546_lo_p
  );


  buf

  (
    n552_li,
    n549_lo_p
  );


  buf

  (
    n564_li,
    n1706_o2_p
  );


  buf

  (
    n579_li,
    G10_p
  );


  buf

  (
    n600_li,
    n1707_o2_p
  );


  buf

  (
    n603_li,
    G12_p
  );


  buf

  (
    n606_li,
    n603_lo_p
  );


  buf

  (
    n609_li,
    n606_lo_p
  );


  buf

  (
    n612_li,
    n609_lo_p
  );


  buf

  (
    n615_li,
    G13_p
  );


  buf

  (
    n618_li,
    n615_lo_p
  );


  buf

  (
    n621_li,
    n618_lo_p
  );


  buf

  (
    n627_li,
    G14_p
  );


  buf

  (
    n630_li,
    n627_lo_p
  );


  buf

  (
    n633_li,
    n630_lo_p
  );


  buf

  (
    n639_li,
    G15_p
  );


  buf

  (
    n642_li,
    n639_lo_p
  );


  buf

  (
    n645_li,
    n642_lo_p
  );


  buf

  (
    n648_li,
    n645_lo_p
  );


  buf

  (
    n660_li,
    n1708_o2_p
  );


  buf

  (
    n663_li,
    G17_p
  );


  buf

  (
    n672_li,
    n1781_o2_p
  );


  buf

  (
    n675_li,
    G18_p
  );


  buf

  (
    n678_li,
    n675_lo_p
  );


  buf

  (
    n681_li,
    n678_lo_p
  );


  buf

  (
    n684_li,
    n681_lo_p
  );


  buf

  (
    n687_li,
    G19_p
  );


  buf

  (
    n690_li,
    n687_lo_p
  );


  buf

  (
    n693_li,
    n690_lo_p
  );


  buf

  (
    n696_li,
    n693_lo_p
  );


  buf

  (
    n699_li,
    G20_p
  );


  buf

  (
    n702_li,
    n699_lo_p
  );


  buf

  (
    n705_li,
    n702_lo_p
  );


  buf

  (
    n708_li,
    n705_lo_p
  );


  buf

  (
    n711_li,
    G21_p
  );


  buf

  (
    n714_li,
    n711_lo_p
  );


  buf

  (
    n717_li,
    n714_lo_p
  );


  buf

  (
    n720_li,
    n717_lo_p
  );


  buf

  (
    n723_li,
    G22_p
  );


  buf

  (
    n726_li,
    n723_lo_p
  );


  buf

  (
    n729_li,
    n726_lo_p
  );


  buf

  (
    n732_li,
    n729_lo_p
  );


  buf

  (
    n735_li,
    G23_p
  );


  buf

  (
    n738_li,
    n735_lo_p
  );


  buf

  (
    n741_li,
    n738_lo_p
  );


  buf

  (
    n744_li,
    n741_lo_p
  );


  buf

  (
    n747_li,
    G24_p
  );


  buf

  (
    n750_li,
    n747_lo_p
  );


  buf

  (
    n756_li,
    n753_lo_buf_o2_p_spl_
  );


  buf

  (
    n759_li,
    G25_p
  );


  buf

  (
    n762_li,
    n759_lo_p
  );


  buf

  (
    n768_li,
    n765_lo_buf_o2_p_spl_
  );


  buf

  (
    n771_li,
    G26_p
  );


  buf

  (
    n774_li,
    n771_lo_p
  );


  buf

  (
    n780_li,
    n777_lo_buf_o2_p_spl_
  );


  buf

  (
    n783_li,
    G27_p
  );


  buf

  (
    n786_li,
    n783_lo_p
  );


  buf

  (
    n792_li,
    n789_lo_buf_o2_p_spl_
  );


  buf

  (
    n795_li,
    G28_p
  );


  buf

  (
    n804_li,
    n801_lo_buf_o2_p_spl_
  );


  buf

  (
    n807_li,
    G29_p
  );


  buf

  (
    n816_li,
    n1798_o2_p_spl_
  );


  buf

  (
    n819_li,
    G30_p
  );


  buf

  (
    n828_li,
    n1799_o2_p_spl_
  );


  buf

  (
    n831_li,
    G31_p
  );


  buf

  (
    n843_li,
    G32_p
  );


  buf

  (
    n846_li,
    n843_lo_p
  );


  buf

  (
    n849_li,
    n846_lo_p
  );


  buf

  (
    n852_li,
    n849_lo_p
  );


  buf

  (
    n855_li,
    G33_p
  );


  buf

  (
    n858_li,
    n855_lo_p
  );


  buf

  (
    n861_li,
    n858_lo_p
  );


  buf

  (
    n864_li,
    n861_lo_p
  );


  buf

  (
    n867_li,
    G34_p
  );


  buf

  (
    n870_li,
    n867_lo_p
  );


  buf

  (
    n879_li,
    G35_p
  );


  buf

  (
    n891_li,
    G36_p
  );


  buf

  (
    n903_li,
    G37_p
  );


  buf

  (
    n915_li,
    G38_p
  );


  buf

  (
    n918_li,
    n915_lo_p
  );


  buf

  (
    n927_li,
    G39_p
  );


  buf

  (
    n951_li,
    G41_p
  );


  buf

  (
    n954_li,
    n951_lo_p
  );


  buf

  (
    n957_li,
    n954_lo_p
  );


  buf

  (
    n960_li,
    n957_lo_p_spl_1
  );


  buf

  (
    n963_li,
    G42_p
  );


  buf

  (
    n966_li,
    n963_lo_p
  );


  buf

  (
    n972_li,
    n969_lo_buf_o2_p_spl_1
  );


  buf

  (
    n975_li,
    G43_p
  );


  buf

  (
    n978_li,
    n975_lo_p
  );


  buf

  (
    n984_li,
    n981_lo_buf_o2_p_spl_1
  );


  buf

  (
    n987_li,
    G44_p
  );


  buf

  (
    n990_li,
    n987_lo_p
  );


  buf

  (
    n996_li,
    n993_lo_buf_o2_p_spl_1
  );


  buf

  (
    n999_li,
    G45_p
  );


  buf

  (
    n1002_li,
    n999_lo_p
  );


  buf

  (
    n1008_li,
    n1005_lo_buf_o2_p_spl_
  );


  buf

  (
    n1011_li,
    G46_p
  );


  buf

  (
    n1014_li,
    n1011_lo_p
  );


  buf

  (
    n1020_li,
    n1017_lo_buf_o2_p_spl_
  );


  buf

  (
    n1023_li,
    G47_p
  );


  buf

  (
    n1026_li,
    n1023_lo_p
  );


  buf

  (
    n1032_li,
    n1029_lo_buf_o2_p_spl_
  );


  buf

  (
    n1035_li,
    G48_p
  );


  buf

  (
    n1038_li,
    n1035_lo_p
  );


  buf

  (
    n1044_li,
    n1041_lo_buf_o2_p_spl_
  );


  buf

  (
    n1047_li,
    G49_p
  );


  buf

  (
    n1050_li,
    n1047_lo_p
  );


  buf

  (
    n1053_li,
    n1050_lo_p
  );


  buf

  (
    n1056_li,
    n1053_lo_p
  );


  buf

  (
    n1059_li,
    G50_p
  );


  buf

  (
    n1062_li,
    n1059_lo_p
  );


  buf

  (
    n1065_li,
    n1062_lo_p
  );


  buf

  (
    n1068_li,
    n1065_lo_p
  );


  buf

  (
    n1071_li,
    G51_p
  );


  buf

  (
    n1074_li,
    n1071_lo_p
  );


  buf

  (
    n1077_li,
    n1074_lo_p
  );


  buf

  (
    n1080_li,
    n1077_lo_p
  );


  buf

  (
    n1083_li,
    G52_p
  );


  buf

  (
    n1086_li,
    n1083_lo_p
  );


  buf

  (
    n1089_li,
    n1086_lo_p
  );


  buf

  (
    n1092_li,
    n1089_lo_p
  );


  buf

  (
    n1095_li,
    G53_p
  );


  buf

  (
    n1098_li,
    n1095_lo_p
  );


  buf

  (
    n1101_li,
    n1098_lo_p
  );


  buf

  (
    n1104_li,
    n1101_lo_p
  );


  buf

  (
    n1107_li,
    G54_p
  );


  buf

  (
    n1110_li,
    n1107_lo_p
  );


  buf

  (
    n1113_li,
    n1110_lo_p
  );


  buf

  (
    n1116_li,
    n1113_lo_p
  );


  buf

  (
    n1119_li,
    G55_p
  );


  buf

  (
    n1122_li,
    n1119_lo_p
  );


  buf

  (
    n1125_li,
    n1122_lo_p
  );


  buf

  (
    n1128_li,
    n1125_lo_p
  );


  buf

  (
    n1131_li,
    G56_p
  );


  buf

  (
    n1134_li,
    n1131_lo_p
  );


  buf

  (
    n1137_li,
    n1134_lo_p
  );


  buf

  (
    n1140_li,
    n1137_lo_p
  );


  buf

  (
    n1143_li,
    G57_p
  );


  buf

  (
    n1146_li,
    n1143_lo_p
  );


  buf

  (
    n1149_li,
    n1146_lo_p
  );


  buf

  (
    n1152_li,
    n1149_lo_p
  );


  buf

  (
    n1155_li,
    G58_p
  );


  buf

  (
    n1158_li,
    n1155_lo_p
  );


  buf

  (
    n1167_li,
    G59_p
  );


  buf

  (
    n1170_li,
    n1167_lo_p
  );


  buf

  (
    n1173_li,
    n1170_lo_p
  );


  buf

  (
    n1176_li,
    n1173_lo_p
  );


  buf

  (
    n1179_li,
    G60_p
  );


  buf

  (
    n1529_i2,
    n1709_o2_p
  );


  buf

  (
    n1616_i2,
    n1828_o2_p
  );


  buf

  (
    n1655_i2,
    G558_o2_p
  );


  buf

  (
    n1656_i2,
    G562_o2_p
  );


  buf

  (
    n1657_i2,
    G566_o2_p
  );


  buf

  (
    n1730_i2,
    G690_o2_p
  );


  buf

  (
    n1731_i2,
    G698_o2_p_spl_
  );


  buf

  (
    n1732_i2,
    G707_o2_p_spl_
  );


  buf

  (
    n1729_i2,
    G554_o2_p
  );


  buf

  (
    n1805_i2,
    G682_o2_p_spl_
  );


  buf

  (
    n1808_i2,
    G546_o2_p_spl_
  );


  buf

  (
    n1807_i2,
    G542_o2_p_spl_
  );


  buf

  (
    n1809_i2,
    G550_o2_p_spl_
  );


  buf

  (
    n1663_i2,
    n1835_o2_p
  );


  buf

  (
    n1664_i2,
    n1836_o2_p
  );


  buf

  (
    n1704_i2,
    n489_lo_buf_o2_p_spl_
  );


  buf

  (
    n1705_i2,
    n513_lo_buf_o2_p
  );


  buf

  (
    n1706_i2,
    n561_lo_buf_o2_p
  );


  buf

  (
    n1707_i2,
    n597_lo_buf_o2_p
  );


  buf

  (
    n1708_i2,
    n657_lo_buf_o2_p
  );


  buf

  (
    n1709_i2,
    G276_o2_p
  );


  not

  (
    G280_i2,
    g502_n_spl_
  );


  buf

  (
    G655_i2,
    g503_p_spl_
  );


  buf

  (
    G663_i2,
    g504_p_spl_1
  );


  buf

  (
    G672_i2,
    g505_p_spl_1
  );


  buf

  (
    G538_i2,
    g508_n_spl_
  );


  buf

  (
    n1780_i2,
    n537_lo_buf_o2_p
  );


  buf

  (
    n1781_i2,
    n669_lo_buf_o2_p
  );


  buf

  (
    n1797_i2,
    n585_lo_buf_o2_p
  );


  buf

  (
    n1798_i2,
    n813_lo_buf_o2_p
  );


  buf

  (
    n1799_i2,
    n825_lo_buf_o2_p
  );


  buf

  (
    n1800_i2,
    n837_lo_buf_o2_p
  );


  buf

  (
    G578_i2,
    g509_n_spl_
  );


  buf

  (
    n1828_i2,
    G369_o2_p_spl_
  );


  buf

  (
    n801_lo_buf_i2,
    n798_lo_buf_o2_p
  );


  buf

  (
    G693_i2,
    g510_p_spl_
  );


  buf

  (
    G702_i2,
    g511_p_spl_
  );


  buf

  (
    G712_i2,
    g512_p_spl_
  );


  buf

  (
    G685_i2,
    g513_p_spl_
  );


  buf

  (
    G658_i2,
    g515_p_spl_
  );


  buf

  (
    G667_i2,
    g517_p_spl_
  );


  buf

  (
    G677_i2,
    g519_p_spl_
  );


  buf

  (
    G650_i2,
    g521_p_spl_
  );


  buf

  (
    G798_i2,
    g531_n_spl_
  );


  buf

  (
    n1017_lo_buf_i2,
    n1014_lo_p
  );


  buf

  (
    n1029_lo_buf_i2,
    n1026_lo_p
  );


  buf

  (
    n1041_lo_buf_i2,
    n1038_lo_p
  );


  not

  (
    G558_i2,
    g534_p_spl_
  );


  not

  (
    G562_i2,
    g536_p_spl_
  );


  not

  (
    G566_i2,
    g538_p_spl_
  );


  buf

  (
    n1835_i2,
    n477_lo_buf_o2_p_spl_
  );


  buf

  (
    n1836_i2,
    n525_lo_buf_o2_p_spl_
  );


  buf

  (
    n1837_i2,
    n573_lo_buf_o2_p_spl_
  );


  buf

  (
    n765_lo_buf_i2,
    n762_lo_p
  );


  buf

  (
    n777_lo_buf_i2,
    n774_lo_p
  );


  buf

  (
    n789_lo_buf_i2,
    n786_lo_p
  );


  not

  (
    G617_i2,
    g539_n_spl_0
  );


  not

  (
    G626_i2,
    g540_n_spl_0
  );


  not

  (
    G636_i2,
    g541_n_spl_0
  );


  buf

  (
    n489_lo_buf_i2,
    n486_lo_buf_o2_p_spl_
  );


  buf

  (
    n513_lo_buf_i2,
    n510_lo_buf_o2_p_spl_1
  );


  buf

  (
    n561_lo_buf_i2,
    n558_lo_buf_o2_p_spl_
  );


  buf

  (
    n597_lo_buf_i2,
    n594_lo_buf_o2_p_spl_
  );


  buf

  (
    n657_lo_buf_i2,
    n654_lo_buf_o2_p
  );


  buf

  (
    G276_i2,
    g543_p_spl_1
  );


  buf

  (
    n1005_lo_buf_i2,
    n1002_lo_p
  );


  buf

  (
    n1161_lo_buf_i2,
    n1158_lo_p
  );


  not

  (
    G620_i2,
    g544_p_spl_
  );


  not

  (
    G629_i2,
    g545_p_spl_
  );


  not

  (
    G639_i2,
    g546_p_spl_
  );


  not

  (
    G554_i2,
    g550_p_spl_
  );


  not

  (
    G690_i2,
    g539_n_spl_
  );


  not

  (
    G698_i2,
    g540_n_spl_
  );


  not

  (
    G707_i2,
    g541_n_spl_
  );


  not

  (
    G319_i2,
    g551_n_spl_
  );


  buf

  (
    G389_i2,
    g543_p_spl_1
  );


  buf

  (
    n753_lo_buf_i2,
    n750_lo_p_spl_
  );


  buf

  (
    G647_i2,
    g520_p_spl_
  );


  buf

  (
    G769_i2,
    g554_p
  );


  buf

  (
    G785_i2,
    g557_p
  );


  buf

  (
    G808_i2,
    g560_p
  );


  buf

  (
    G445_i2,
    g569_p
  );


  buf

  (
    G448_i2,
    g578_p
  );


  buf

  (
    G477_i2,
    g587_p
  );


  buf

  (
    G480_i2,
    g596_p
  );


  not

  (
    G436_i2,
    g601_n
  );


  buf

  (
    G786_i2,
    g609_p
  );


  buf

  (
    G787_i2,
    g614_p
  );


  buf

  (
    G826_i2,
    g622_p
  );


  buf

  (
    G827_i2,
    g627_p
  );


  buf

  (
    G825_i2,
    g630_p
  );


  not

  (
    G610_i2,
    g631_n_spl_
  );


  buf

  (
    n537_lo_buf_i2,
    n531_lo_p
  );


  buf

  (
    n669_lo_buf_i2,
    n663_lo_p
  );


  buf

  (
    n969_lo_buf_i2,
    n966_lo_p
  );


  buf

  (
    n981_lo_buf_i2,
    n978_lo_p
  );


  buf

  (
    n993_lo_buf_i2,
    n990_lo_p
  );


  buf

  (
    G309_i2,
    g632_p
  );


  not

  (
    G461_i2,
    g635_n_spl_1
  );


  buf

  (
    G487_i2,
    g636_p
  );


  not

  (
    G460_i2,
    g639_n
  );


  not

  (
    G468_i2,
    g642_n_spl_1
  );


  not

  (
    G287_i2,
    g644_n_spl_
  );


  not

  (
    G613_i2,
    g645_p
  );


  buf

  (
    n585_lo_buf_i2,
    n579_lo_p
  );


  buf

  (
    n813_lo_buf_i2,
    n807_lo_p_spl_
  );


  buf

  (
    n825_lo_buf_i2,
    n819_lo_p_spl_
  );


  buf

  (
    n837_lo_buf_i2,
    n831_lo_p_spl_
  );


  buf

  (
    n897_lo_buf_i2,
    n891_lo_p_spl_
  );


  buf

  (
    n909_lo_buf_i2,
    n903_lo_p_spl_
  );


  buf

  (
    n933_lo_buf_i2,
    n927_lo_p_spl_
  );


  buf

  (
    G451_i2,
    g658_n_spl_1
  );


  not

  (
    G682_i2,
    g631_n_spl_
  );


  not

  (
    G756_i2,
    g666_p
  );


  not

  (
    G542_i2,
    g672_p
  );


  not

  (
    G546_i2,
    g678_p
  );


  not

  (
    G550_i2,
    g684_p
  );


  buf

  (
    G310_i2,
    n1179_lo_p_spl_
  );


  buf

  (
    n798_lo_buf_i2,
    n795_lo_p
  );


  buf

  (
    n882_lo_buf_i2,
    n879_lo_p
  );


  not

  (
    G427_i2,
    g686_n
  );


  buf

  (
    G497_i2,
    g687_p
  );


  buf

  (
    G499_i2,
    g688_p
  );


  buf

  (
    G501_i2,
    g689_p
  );


  buf

  (
    G498_i2,
    g690_p
  );


  buf

  (
    G500_i2,
    g691_p
  );


  buf

  (
    G502_i2,
    g692_p
  );


  buf

  (
    G369_i2,
    n1179_lo_p_spl_
  );


  buf

  (
    n939_lo_buf_i2,
    G40_p
  );


  buf

  (
    n486_lo_buf_i2,
    G2_p
  );


  buf

  (
    n510_lo_buf_i2,
    G4_p
  );


  buf

  (
    n558_lo_buf_i2,
    G8_p
  );


  buf

  (
    n594_lo_buf_i2,
    G11_p
  );


  buf

  (
    n654_lo_buf_i2,
    G16_p
  );


  buf

  (
    n477_lo_buf_i2,
    G1_p
  );


  buf

  (
    n525_lo_buf_i2,
    G5_p
  );


  buf

  (
    n573_lo_buf_i2,
    G9_p
  );


  buf

  (
    n540_lo_n_spl_,
    n540_lo_n
  );


  buf

  (
    n540_lo_n_spl_0,
    n540_lo_n_spl_
  );


  buf

  (
    n564_lo_n_spl_,
    n564_lo_n
  );


  buf

  (
    n564_lo_n_spl_0,
    n564_lo_n_spl_
  );


  buf

  (
    n552_lo_n_spl_,
    n552_lo_n
  );


  buf

  (
    g361_n_spl_,
    g361_n
  );


  buf

  (
    n672_lo_n_spl_,
    n672_lo_n
  );


  buf

  (
    n480_lo_n_spl_,
    n480_lo_n
  );


  buf

  (
    n504_lo_n_spl_,
    n504_lo_n
  );


  buf

  (
    n516_lo_n_spl_,
    n516_lo_n
  );


  buf

  (
    g363_n_spl_,
    g363_n
  );


  buf

  (
    g363_n_spl_0,
    g363_n_spl_
  );


  buf

  (
    n600_lo_n_spl_,
    n600_lo_n
  );


  buf

  (
    g374_n_spl_,
    g374_n
  );


  buf

  (
    g377_n_spl_,
    g377_n
  );


  buf

  (
    n612_lo_n_spl_,
    n612_lo_n
  );


  buf

  (
    G280_o2_n_spl_,
    G280_o2_n
  );


  buf

  (
    G445_o2_p_spl_,
    G445_o2_p
  );


  buf

  (
    n852_lo_p_spl_,
    n852_lo_p
  );


  buf

  (
    n852_lo_p_spl_0,
    n852_lo_p_spl_
  );


  buf

  (
    n852_lo_p_spl_1,
    n852_lo_p_spl_
  );


  buf

  (
    G445_o2_n_spl_,
    G445_o2_n
  );


  buf

  (
    n852_lo_n_spl_,
    n852_lo_n
  );


  buf

  (
    n852_lo_n_spl_0,
    n852_lo_n_spl_
  );


  buf

  (
    n852_lo_n_spl_1,
    n852_lo_n_spl_
  );


  buf

  (
    G448_o2_p_spl_,
    G448_o2_p
  );


  buf

  (
    n864_lo_p_spl_,
    n864_lo_p
  );


  buf

  (
    G448_o2_n_spl_,
    G448_o2_n
  );


  buf

  (
    n864_lo_n_spl_,
    n864_lo_n
  );


  buf

  (
    G477_o2_p_spl_,
    G477_o2_p
  );


  buf

  (
    G477_o2_n_spl_,
    G477_o2_n
  );


  buf

  (
    G480_o2_p_spl_,
    G480_o2_p
  );


  buf

  (
    n1056_lo_p_spl_,
    n1056_lo_p
  );


  buf

  (
    G480_o2_n_spl_,
    G480_o2_n
  );


  buf

  (
    n1056_lo_n_spl_,
    n1056_lo_n
  );


  buf

  (
    n1068_lo_n_spl_,
    n1068_lo_n
  );


  buf

  (
    n1068_lo_n_spl_0,
    n1068_lo_n_spl_
  );


  buf

  (
    n1068_lo_n_spl_00,
    n1068_lo_n_spl_0
  );


  buf

  (
    n1068_lo_n_spl_01,
    n1068_lo_n_spl_0
  );


  buf

  (
    n1068_lo_n_spl_1,
    n1068_lo_n_spl_
  );


  buf

  (
    n1068_lo_n_spl_10,
    n1068_lo_n_spl_1
  );


  buf

  (
    n1068_lo_n_spl_11,
    n1068_lo_n_spl_1
  );


  buf

  (
    n1080_lo_n_spl_,
    n1080_lo_n
  );


  buf

  (
    n1080_lo_n_spl_0,
    n1080_lo_n_spl_
  );


  buf

  (
    n1080_lo_n_spl_00,
    n1080_lo_n_spl_0
  );


  buf

  (
    n1080_lo_n_spl_01,
    n1080_lo_n_spl_0
  );


  buf

  (
    n1080_lo_n_spl_1,
    n1080_lo_n_spl_
  );


  buf

  (
    n1080_lo_n_spl_10,
    n1080_lo_n_spl_1
  );


  buf

  (
    n1080_lo_n_spl_11,
    n1080_lo_n_spl_1
  );


  buf

  (
    n1092_lo_n_spl_,
    n1092_lo_n
  );


  buf

  (
    n1092_lo_n_spl_0,
    n1092_lo_n_spl_
  );


  buf

  (
    n1092_lo_n_spl_00,
    n1092_lo_n_spl_0
  );


  buf

  (
    n1092_lo_n_spl_01,
    n1092_lo_n_spl_0
  );


  buf

  (
    n1092_lo_n_spl_1,
    n1092_lo_n_spl_
  );


  buf

  (
    n1092_lo_n_spl_10,
    n1092_lo_n_spl_1
  );


  buf

  (
    n1092_lo_n_spl_11,
    n1092_lo_n_spl_1
  );


  buf

  (
    n1104_lo_n_spl_,
    n1104_lo_n
  );


  buf

  (
    n1104_lo_n_spl_0,
    n1104_lo_n_spl_
  );


  buf

  (
    n1104_lo_n_spl_00,
    n1104_lo_n_spl_0
  );


  buf

  (
    n1104_lo_n_spl_01,
    n1104_lo_n_spl_0
  );


  buf

  (
    n1104_lo_n_spl_1,
    n1104_lo_n_spl_
  );


  buf

  (
    n1104_lo_n_spl_10,
    n1104_lo_n_spl_1
  );


  buf

  (
    n1104_lo_n_spl_11,
    n1104_lo_n_spl_1
  );


  buf

  (
    n1128_lo_n_spl_,
    n1128_lo_n
  );


  buf

  (
    n1128_lo_n_spl_0,
    n1128_lo_n_spl_
  );


  buf

  (
    n1116_lo_n_spl_,
    n1116_lo_n
  );


  buf

  (
    n1116_lo_n_spl_0,
    n1116_lo_n_spl_
  );


  buf

  (
    n1116_lo_n_spl_00,
    n1116_lo_n_spl_0
  );


  buf

  (
    n1116_lo_n_spl_01,
    n1116_lo_n_spl_0
  );


  buf

  (
    n1116_lo_n_spl_1,
    n1116_lo_n_spl_
  );


  buf

  (
    n1116_lo_n_spl_10,
    n1116_lo_n_spl_1
  );


  buf

  (
    n1116_lo_n_spl_11,
    n1116_lo_n_spl_1
  );


  buf

  (
    G436_o2_n_spl_,
    G436_o2_n
  );


  buf

  (
    G436_o2_n_spl_0,
    G436_o2_n_spl_
  );


  buf

  (
    G436_o2_n_spl_00,
    G436_o2_n_spl_0
  );


  buf

  (
    G436_o2_n_spl_01,
    G436_o2_n_spl_0
  );


  buf

  (
    G436_o2_n_spl_1,
    G436_o2_n_spl_
  );


  buf

  (
    G436_o2_n_spl_10,
    G436_o2_n_spl_1
  );


  buf

  (
    G436_o2_n_spl_11,
    G436_o2_n_spl_1
  );


  buf

  (
    G647_o2_n_spl_,
    G647_o2_n
  );


  buf

  (
    G542_o2_p_spl_,
    G542_o2_p
  );


  buf

  (
    G542_o2_p_spl_0,
    G542_o2_p_spl_
  );


  buf

  (
    n969_lo_buf_o2_p_spl_,
    n969_lo_buf_o2_p
  );


  buf

  (
    n969_lo_buf_o2_p_spl_0,
    n969_lo_buf_o2_p_spl_
  );


  buf

  (
    n969_lo_buf_o2_p_spl_00,
    n969_lo_buf_o2_p_spl_0
  );


  buf

  (
    n969_lo_buf_o2_p_spl_1,
    n969_lo_buf_o2_p_spl_
  );


  buf

  (
    G542_o2_n_spl_,
    G542_o2_n
  );


  buf

  (
    n969_lo_buf_o2_n_spl_,
    n969_lo_buf_o2_n
  );


  buf

  (
    n969_lo_buf_o2_n_spl_0,
    n969_lo_buf_o2_n_spl_
  );


  buf

  (
    n969_lo_buf_o2_n_spl_1,
    n969_lo_buf_o2_n_spl_
  );


  buf

  (
    G546_o2_p_spl_,
    G546_o2_p
  );


  buf

  (
    G546_o2_p_spl_0,
    G546_o2_p_spl_
  );


  buf

  (
    n981_lo_buf_o2_p_spl_,
    n981_lo_buf_o2_p
  );


  buf

  (
    n981_lo_buf_o2_p_spl_0,
    n981_lo_buf_o2_p_spl_
  );


  buf

  (
    n981_lo_buf_o2_p_spl_00,
    n981_lo_buf_o2_p_spl_0
  );


  buf

  (
    n981_lo_buf_o2_p_spl_1,
    n981_lo_buf_o2_p_spl_
  );


  buf

  (
    G546_o2_n_spl_,
    G546_o2_n
  );


  buf

  (
    n981_lo_buf_o2_n_spl_,
    n981_lo_buf_o2_n
  );


  buf

  (
    n981_lo_buf_o2_n_spl_0,
    n981_lo_buf_o2_n_spl_
  );


  buf

  (
    n981_lo_buf_o2_n_spl_1,
    n981_lo_buf_o2_n_spl_
  );


  buf

  (
    G550_o2_p_spl_,
    G550_o2_p
  );


  buf

  (
    G550_o2_p_spl_0,
    G550_o2_p_spl_
  );


  buf

  (
    n993_lo_buf_o2_p_spl_,
    n993_lo_buf_o2_p
  );


  buf

  (
    n993_lo_buf_o2_p_spl_0,
    n993_lo_buf_o2_p_spl_
  );


  buf

  (
    n993_lo_buf_o2_p_spl_00,
    n993_lo_buf_o2_p_spl_0
  );


  buf

  (
    n993_lo_buf_o2_p_spl_1,
    n993_lo_buf_o2_p_spl_
  );


  buf

  (
    G550_o2_n_spl_,
    G550_o2_n
  );


  buf

  (
    n993_lo_buf_o2_n_spl_,
    n993_lo_buf_o2_n
  );


  buf

  (
    n993_lo_buf_o2_n_spl_0,
    n993_lo_buf_o2_n_spl_
  );


  buf

  (
    n993_lo_buf_o2_n_spl_1,
    n993_lo_buf_o2_n_spl_
  );


  buf

  (
    g508_p_spl_,
    g508_p
  );


  buf

  (
    n957_lo_n_spl_,
    n957_lo_n
  );


  buf

  (
    n957_lo_n_spl_0,
    n957_lo_n_spl_
  );


  buf

  (
    n957_lo_n_spl_1,
    n957_lo_n_spl_
  );


  buf

  (
    g508_n_spl_,
    g508_n
  );


  buf

  (
    g508_n_spl_0,
    g508_n_spl_
  );


  buf

  (
    n957_lo_p_spl_,
    n957_lo_p
  );


  buf

  (
    n957_lo_p_spl_0,
    n957_lo_p_spl_
  );


  buf

  (
    n957_lo_p_spl_00,
    n957_lo_p_spl_0
  );


  buf

  (
    n957_lo_p_spl_1,
    n957_lo_p_spl_
  );


  buf

  (
    G629_o2_p_spl_,
    G629_o2_p
  );


  buf

  (
    G629_o2_p_spl_0,
    G629_o2_p_spl_
  );


  buf

  (
    G629_o2_n_spl_,
    G629_o2_n
  );


  buf

  (
    G629_o2_n_spl_0,
    G629_o2_n_spl_
  );


  buf

  (
    G639_o2_p_spl_,
    G639_o2_p
  );


  buf

  (
    G639_o2_p_spl_0,
    G639_o2_p_spl_
  );


  buf

  (
    G639_o2_n_spl_,
    G639_o2_n
  );


  buf

  (
    G639_o2_n_spl_0,
    G639_o2_n_spl_
  );


  buf

  (
    G613_o2_p_spl_,
    G613_o2_p
  );


  buf

  (
    G613_o2_n_spl_,
    G613_o2_n
  );


  buf

  (
    g514_n_spl_,
    g514_n
  );


  buf

  (
    g514_n_spl_0,
    g514_n_spl_
  );


  buf

  (
    g503_n_spl_,
    g503_n
  );


  buf

  (
    g514_p_spl_,
    g514_p
  );


  buf

  (
    g514_p_spl_0,
    g514_p_spl_
  );


  buf

  (
    g503_p_spl_,
    g503_p
  );


  buf

  (
    g503_p_spl_0,
    g503_p_spl_
  );


  buf

  (
    g516_n_spl_,
    g516_n
  );


  buf

  (
    g516_n_spl_0,
    g516_n_spl_
  );


  buf

  (
    g516_n_spl_1,
    g516_n_spl_
  );


  buf

  (
    g504_n_spl_,
    g504_n
  );


  buf

  (
    g504_n_spl_0,
    g504_n_spl_
  );


  buf

  (
    g516_p_spl_,
    g516_p
  );


  buf

  (
    g516_p_spl_0,
    g516_p_spl_
  );


  buf

  (
    g516_p_spl_1,
    g516_p_spl_
  );


  buf

  (
    g504_p_spl_,
    g504_p
  );


  buf

  (
    g504_p_spl_0,
    g504_p_spl_
  );


  buf

  (
    g504_p_spl_1,
    g504_p_spl_
  );


  buf

  (
    g518_n_spl_,
    g518_n
  );


  buf

  (
    g518_n_spl_0,
    g518_n_spl_
  );


  buf

  (
    g518_n_spl_1,
    g518_n_spl_
  );


  buf

  (
    g505_n_spl_,
    g505_n
  );


  buf

  (
    g505_n_spl_0,
    g505_n_spl_
  );


  buf

  (
    g505_n_spl_1,
    g505_n_spl_
  );


  buf

  (
    g518_p_spl_,
    g518_p
  );


  buf

  (
    g518_p_spl_0,
    g518_p_spl_
  );


  buf

  (
    g518_p_spl_1,
    g518_p_spl_
  );


  buf

  (
    g505_p_spl_,
    g505_p
  );


  buf

  (
    g505_p_spl_0,
    g505_p_spl_
  );


  buf

  (
    g505_p_spl_00,
    g505_p_spl_0
  );


  buf

  (
    g505_p_spl_1,
    g505_p_spl_
  );


  buf

  (
    g509_n_spl_,
    g509_n
  );


  buf

  (
    g520_p_spl_,
    g520_p
  );


  buf

  (
    g523_p_spl_,
    g523_p
  );


  buf

  (
    g523_n_spl_,
    g523_n
  );


  buf

  (
    G756_o2_p_spl_,
    G756_o2_p
  );


  buf

  (
    G756_o2_n_spl_,
    G756_o2_n
  );


  buf

  (
    G682_o2_p_spl_,
    G682_o2_p
  );


  buf

  (
    g526_n_spl_,
    g526_n
  );


  buf

  (
    g526_n_spl_0,
    g526_n_spl_
  );


  buf

  (
    g526_n_spl_1,
    g526_n_spl_
  );


  buf

  (
    g526_p_spl_,
    g526_p
  );


  buf

  (
    g526_p_spl_0,
    g526_p_spl_
  );


  buf

  (
    g526_p_spl_1,
    g526_p_spl_
  );


  buf

  (
    G369_o2_p_spl_,
    G369_o2_p
  );


  buf

  (
    g532_n_spl_,
    g532_n
  );


  buf

  (
    g532_n_spl_0,
    g532_n_spl_
  );


  buf

  (
    g532_n_spl_1,
    g532_n_spl_
  );


  buf

  (
    g534_p_spl_,
    g534_p
  );


  buf

  (
    g534_p_spl_0,
    g534_p_spl_
  );


  buf

  (
    n1014_lo_n_spl_,
    n1014_lo_n
  );


  buf

  (
    g536_p_spl_,
    g536_p
  );


  buf

  (
    g536_p_spl_0,
    g536_p_spl_
  );


  buf

  (
    n1026_lo_n_spl_,
    n1026_lo_n
  );


  buf

  (
    g538_p_spl_,
    g538_p
  );


  buf

  (
    g538_p_spl_0,
    g538_p_spl_
  );


  buf

  (
    n1038_lo_n_spl_,
    n1038_lo_n
  );


  buf

  (
    n525_lo_buf_o2_p_spl_,
    n525_lo_buf_o2_p
  );


  buf

  (
    n477_lo_buf_o2_p_spl_,
    n477_lo_buf_o2_p
  );


  buf

  (
    n477_lo_buf_o2_p_spl_0,
    n477_lo_buf_o2_p_spl_
  );


  buf

  (
    n477_lo_buf_o2_n_spl_,
    n477_lo_buf_o2_n
  );


  buf

  (
    n573_lo_buf_o2_p_spl_,
    n573_lo_buf_o2_p
  );


  buf

  (
    n573_lo_buf_o2_p_spl_0,
    n573_lo_buf_o2_p_spl_
  );


  buf

  (
    n882_lo_buf_o2_n_spl_,
    n882_lo_buf_o2_n
  );


  buf

  (
    G451_o2_n_spl_,
    G451_o2_n
  );


  buf

  (
    G451_o2_n_spl_0,
    G451_o2_n_spl_
  );


  buf

  (
    G451_o2_n_spl_1,
    G451_o2_n_spl_
  );


  buf

  (
    n594_lo_buf_o2_n_spl_,
    n594_lo_buf_o2_n
  );


  buf

  (
    g512_p_spl_,
    g512_p
  );


  buf

  (
    n1161_lo_buf_o2_p_spl_,
    n1161_lo_buf_o2_p
  );


  buf

  (
    n1161_lo_buf_o2_p_spl_0,
    n1161_lo_buf_o2_p_spl_
  );


  buf

  (
    n1161_lo_buf_o2_n_spl_,
    n1161_lo_buf_o2_n
  );


  buf

  (
    n1161_lo_buf_o2_n_spl_0,
    n1161_lo_buf_o2_n_spl_
  );


  buf

  (
    g513_p_spl_,
    g513_p
  );


  buf

  (
    g519_p_spl_,
    g519_p
  );


  buf

  (
    n753_lo_buf_o2_p_spl_,
    n753_lo_buf_o2_p
  );


  buf

  (
    n753_lo_buf_o2_p_spl_0,
    n753_lo_buf_o2_p_spl_
  );


  buf

  (
    n765_lo_buf_o2_p_spl_,
    n765_lo_buf_o2_p
  );


  buf

  (
    n765_lo_buf_o2_p_spl_0,
    n765_lo_buf_o2_p_spl_
  );


  buf

  (
    n753_lo_buf_o2_n_spl_,
    n753_lo_buf_o2_n
  );


  buf

  (
    n765_lo_buf_o2_n_spl_,
    n765_lo_buf_o2_n
  );


  buf

  (
    n789_lo_buf_o2_p_spl_,
    n789_lo_buf_o2_p
  );


  buf

  (
    n789_lo_buf_o2_p_spl_0,
    n789_lo_buf_o2_p_spl_
  );


  buf

  (
    n777_lo_buf_o2_p_spl_,
    n777_lo_buf_o2_p
  );


  buf

  (
    n777_lo_buf_o2_p_spl_0,
    n777_lo_buf_o2_p_spl_
  );


  buf

  (
    n789_lo_buf_o2_n_spl_,
    n789_lo_buf_o2_n
  );


  buf

  (
    n777_lo_buf_o2_n_spl_,
    n777_lo_buf_o2_n
  );


  buf

  (
    n801_lo_buf_o2_p_spl_,
    n801_lo_buf_o2_p
  );


  buf

  (
    n801_lo_buf_o2_p_spl_0,
    n801_lo_buf_o2_p_spl_
  );


  buf

  (
    n1798_o2_p_spl_,
    n1798_o2_p
  );


  buf

  (
    n1798_o2_p_spl_0,
    n1798_o2_p_spl_
  );


  buf

  (
    n801_lo_buf_o2_n_spl_,
    n801_lo_buf_o2_n
  );


  buf

  (
    n1798_o2_n_spl_,
    n1798_o2_n
  );


  buf

  (
    n1800_o2_p_spl_,
    n1800_o2_p
  );


  buf

  (
    n1799_o2_p_spl_,
    n1799_o2_p
  );


  buf

  (
    n1799_o2_p_spl_0,
    n1799_o2_p_spl_
  );


  buf

  (
    n1800_o2_n_spl_,
    n1800_o2_n
  );


  buf

  (
    n1799_o2_n_spl_,
    n1799_o2_n
  );


  buf

  (
    n1005_lo_buf_o2_p_spl_,
    n1005_lo_buf_o2_p
  );


  buf

  (
    n1005_lo_buf_o2_p_spl_0,
    n1005_lo_buf_o2_p_spl_
  );


  buf

  (
    n1017_lo_buf_o2_p_spl_,
    n1017_lo_buf_o2_p
  );


  buf

  (
    n1017_lo_buf_o2_p_spl_0,
    n1017_lo_buf_o2_p_spl_
  );


  buf

  (
    n1005_lo_buf_o2_n_spl_,
    n1005_lo_buf_o2_n
  );


  buf

  (
    n1017_lo_buf_o2_n_spl_,
    n1017_lo_buf_o2_n
  );


  buf

  (
    n1041_lo_buf_o2_p_spl_,
    n1041_lo_buf_o2_p
  );


  buf

  (
    n1041_lo_buf_o2_p_spl_0,
    n1041_lo_buf_o2_p_spl_
  );


  buf

  (
    n1029_lo_buf_o2_p_spl_,
    n1029_lo_buf_o2_p
  );


  buf

  (
    n1029_lo_buf_o2_p_spl_0,
    n1029_lo_buf_o2_p_spl_
  );


  buf

  (
    n1041_lo_buf_o2_n_spl_,
    n1041_lo_buf_o2_n
  );


  buf

  (
    n1029_lo_buf_o2_n_spl_,
    n1029_lo_buf_o2_n
  );


  buf

  (
    g502_n_spl_,
    g502_n
  );


  buf

  (
    G707_o2_p_spl_,
    G707_o2_p
  );


  buf

  (
    G707_o2_p_spl_0,
    G707_o2_p_spl_
  );


  buf

  (
    G707_o2_n_spl_,
    G707_o2_n
  );


  buf

  (
    G698_o2_p_spl_,
    G698_o2_p
  );


  buf

  (
    g510_p_spl_,
    g510_p
  );


  buf

  (
    g511_p_spl_,
    g511_p
  );


  buf

  (
    g515_p_spl_,
    g515_p
  );


  buf

  (
    g517_p_spl_,
    g517_p
  );


  buf

  (
    g531_n_spl_,
    g531_n
  );


  buf

  (
    g521_p_spl_,
    g521_p
  );


  buf

  (
    g550_p_spl_,
    g550_p
  );


  buf

  (
    g550_p_spl_0,
    g550_p_spl_
  );


  buf

  (
    n1002_lo_n_spl_,
    n1002_lo_n
  );


  buf

  (
    n489_lo_buf_o2_p_spl_,
    n489_lo_buf_o2_p
  );


  buf

  (
    G389_o2_n_spl_,
    G389_o2_n
  );


  buf

  (
    n513_lo_buf_o2_n_spl_,
    n513_lo_buf_o2_n
  );


  buf

  (
    n750_lo_p_spl_,
    n750_lo_p
  );


  buf

  (
    g638_n_spl_,
    g638_n
  );


  buf

  (
    g638_n_spl_0,
    g638_n_spl_
  );


  buf

  (
    g638_n_spl_1,
    g638_n_spl_
  );


  buf

  (
    g551_n_spl_,
    g551_n
  );


  buf

  (
    g543_p_spl_,
    g543_p
  );


  buf

  (
    g543_p_spl_0,
    g543_p_spl_
  );


  buf

  (
    g543_p_spl_1,
    g543_p_spl_
  );


  buf

  (
    n510_lo_buf_o2_p_spl_,
    n510_lo_buf_o2_p
  );


  buf

  (
    n510_lo_buf_o2_p_spl_0,
    n510_lo_buf_o2_p_spl_
  );


  buf

  (
    n510_lo_buf_o2_p_spl_1,
    n510_lo_buf_o2_p_spl_
  );


  buf

  (
    n654_lo_buf_o2_n_spl_,
    n654_lo_buf_o2_n
  );


  buf

  (
    n558_lo_buf_o2_p_spl_,
    n558_lo_buf_o2_p
  );


  buf

  (
    n558_lo_buf_o2_n_spl_,
    n558_lo_buf_o2_n
  );


  buf

  (
    n594_lo_buf_o2_p_spl_,
    n594_lo_buf_o2_p
  );


  buf

  (
    n486_lo_buf_o2_p_spl_,
    n486_lo_buf_o2_p
  );


  buf

  (
    g544_p_spl_,
    g544_p
  );


  buf

  (
    g544_p_spl_0,
    g544_p_spl_
  );


  buf

  (
    g540_n_spl_,
    g540_n
  );


  buf

  (
    g540_n_spl_0,
    g540_n_spl_
  );


  buf

  (
    g545_p_spl_,
    g545_p
  );


  buf

  (
    g660_n_spl_,
    g660_n
  );


  buf

  (
    g541_n_spl_,
    g541_n
  );


  buf

  (
    g541_n_spl_0,
    g541_n_spl_
  );


  buf

  (
    g546_p_spl_,
    g546_p
  );


  buf

  (
    g539_n_spl_,
    g539_n
  );


  buf

  (
    g539_n_spl_0,
    g539_n_spl_
  );


  buf

  (
    n870_lo_n_spl_,
    n870_lo_n
  );


  buf

  (
    n870_lo_n_spl_0,
    n870_lo_n_spl_
  );


  buf

  (
    g635_n_spl_,
    g635_n
  );


  buf

  (
    g635_n_spl_0,
    g635_n_spl_
  );


  buf

  (
    g635_n_spl_1,
    g635_n_spl_
  );


  buf

  (
    g644_n_spl_,
    g644_n
  );


  buf

  (
    g642_n_spl_,
    g642_n
  );


  buf

  (
    g642_n_spl_0,
    g642_n_spl_
  );


  buf

  (
    g642_n_spl_1,
    g642_n_spl_
  );


  buf

  (
    n891_lo_p_spl_,
    n891_lo_p
  );


  buf

  (
    n903_lo_p_spl_,
    n903_lo_p
  );


  buf

  (
    n927_lo_p_spl_,
    n927_lo_p
  );


  buf

  (
    g658_n_spl_,
    g658_n
  );


  buf

  (
    g658_n_spl_0,
    g658_n_spl_
  );


  buf

  (
    g658_n_spl_1,
    g658_n_spl_
  );


  buf

  (
    n807_lo_p_spl_,
    n807_lo_p
  );


  buf

  (
    n819_lo_p_spl_,
    n819_lo_p
  );


  buf

  (
    n831_lo_p_spl_,
    n831_lo_p
  );


  buf

  (
    g631_n_spl_,
    g631_n
  );


  buf

  (
    n1179_lo_p_spl_,
    n1179_lo_p
  );


endmodule
