
module mymod
(
  G1_p,
  G1_n,
  G2_p,
  G2_n,
  G3_p,
  G3_n,
  G4_p,
  G4_n,
  G5_p,
  G5_n,
  G6_p,
  G6_n,
  G7_p,
  G7_n,
  G8_p,
  G8_n,
  G9_p,
  G9_n,
  G10_p,
  G10_n,
  G11_p,
  G11_n,
  G12_p,
  G12_n,
  G13_p,
  G13_n,
  G14_p,
  G14_n,
  G15_p,
  G15_n,
  G16_p,
  G16_n,
  G17_p,
  G17_n,
  G18_p,
  G18_n,
  G19_p,
  G19_n,
  G20_p,
  G20_n,
  G21_p,
  G21_n,
  G22_p,
  G22_n,
  G23_p,
  G23_n,
  G24_p,
  G24_n,
  G25_p,
  G25_n,
  G26_p,
  G26_n,
  G27_p,
  G27_n,
  G28_p,
  G28_n,
  G29_p,
  G29_n,
  G30_p,
  G30_n,
  G31_p,
  G31_n,
  G32_p,
  G32_n,
  G33_p,
  G33_n,
  G34_p,
  G34_n,
  G35_p,
  G35_n,
  G36_p,
  G36_n,
  G37_p,
  G37_n,
  G38_p,
  G38_n,
  G39_p,
  G39_n,
  G40_p,
  G40_n,
  G41_p,
  G41_n,
  G42_p,
  G42_n,
  G43_p,
  G43_n,
  G44_p,
  G44_n,
  G45_p,
  G45_n,
  G46_p,
  G46_n,
  G47_p,
  G47_n,
  G48_p,
  G48_n,
  G49_p,
  G49_n,
  G50_p,
  G50_n,
  G3519_p,
  G3520_p,
  G3521_p,
  G3522_p,
  G3523_p,
  G3524_p,
  G3525_p,
  G3526_p,
  G3527_p,
  G3528_p,
  G3529_p,
  G3530_p,
  G3531_p,
  G3532_p,
  G3533_p,
  G3534_p,
  G3535_p,
  G3536_p,
  G3537_p,
  G3538_n,
  G3539_p,
  G3540_p
);

  input G1_p;input G1_n;input G2_p;input G2_n;input G3_p;input G3_n;input G4_p;input G4_n;input G5_p;input G5_n;input G6_p;input G6_n;input G7_p;input G7_n;input G8_p;input G8_n;input G9_p;input G9_n;input G10_p;input G10_n;input G11_p;input G11_n;input G12_p;input G12_n;input G13_p;input G13_n;input G14_p;input G14_n;input G15_p;input G15_n;input G16_p;input G16_n;input G17_p;input G17_n;input G18_p;input G18_n;input G19_p;input G19_n;input G20_p;input G20_n;input G21_p;input G21_n;input G22_p;input G22_n;input G23_p;input G23_n;input G24_p;input G24_n;input G25_p;input G25_n;input G26_p;input G26_n;input G27_p;input G27_n;input G28_p;input G28_n;input G29_p;input G29_n;input G30_p;input G30_n;input G31_p;input G31_n;input G32_p;input G32_n;input G33_p;input G33_n;input G34_p;input G34_n;input G35_p;input G35_n;input G36_p;input G36_n;input G37_p;input G37_n;input G38_p;input G38_n;input G39_p;input G39_n;input G40_p;input G40_n;input G41_p;input G41_n;input G42_p;input G42_n;input G43_p;input G43_n;input G44_p;input G44_n;input G45_p;input G45_n;input G46_p;input G46_n;input G47_p;input G47_n;input G48_p;input G48_n;input G49_p;input G49_n;input G50_p;input G50_n;
  output G3519_p;output G3520_p;output G3521_p;output G3522_p;output G3523_p;output G3524_p;output G3525_p;output G3526_p;output G3527_p;output G3528_p;output G3529_p;output G3530_p;output G3531_p;output G3532_p;output G3533_p;output G3534_p;output G3535_p;output G3536_p;output G3537_p;output G3538_n;output G3539_p;output G3540_p;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire ffc_0_p;
  wire ffc_0_n;
  wire ffc_1_p;
  wire ffc_1_n;
  wire ffc_2_p;
  wire ffc_2_n;
  wire ffc_3_p;
  wire ffc_3_n;
  wire ffc_4_p;
  wire ffc_4_n;
  wire ffc_5_p;
  wire ffc_5_n;
  wire ffc_6_p;
  wire ffc_6_n;
  wire ffc_7_p;
  wire ffc_7_n;
  wire ffc_8_p;
  wire ffc_8_n;
  wire ffc_9_p;
  wire ffc_9_n;
  wire ffc_10_p;
  wire ffc_10_n;
  wire ffc_11_p;
  wire ffc_11_n;
  wire ffc_12_p;
  wire ffc_12_n;
  wire ffc_13_p;
  wire ffc_13_n;
  wire ffc_14_p;
  wire ffc_14_n;
  wire ffc_15_p;
  wire ffc_15_n;
  wire ffc_16_p;
  wire ffc_16_n;
  wire ffc_17_p;
  wire ffc_17_n;
  wire ffc_18_p;
  wire ffc_18_n;
  wire ffc_19_p;
  wire ffc_19_n;
  wire ffc_20_p;
  wire ffc_20_n;
  wire ffc_21_p;
  wire ffc_21_n;
  wire ffc_22_p;
  wire ffc_22_n;
  wire ffc_23_p;
  wire ffc_23_n;
  wire ffc_24_p;
  wire ffc_24_n;
  wire ffc_25_p;
  wire ffc_25_n;
  wire ffc_26_p;
  wire ffc_26_n;
  wire ffc_27_p;
  wire ffc_27_n;
  wire ffc_28_p;
  wire ffc_28_n;
  wire ffc_29_p;
  wire ffc_29_n;
  wire ffc_30_p;
  wire ffc_30_n;
  wire ffc_31_p;
  wire ffc_31_n;
  wire ffc_32_p;
  wire ffc_32_n;
  wire ffc_33_p;
  wire ffc_33_n;
  wire ffc_34_p;
  wire ffc_34_n;
  wire ffc_35_p;
  wire ffc_35_n;
  wire ffc_36_p;
  wire ffc_36_n;
  wire ffc_37_p;
  wire ffc_37_n;
  wire ffc_38_p;
  wire ffc_38_n;
  wire ffc_39_p;
  wire ffc_39_n;
  wire ffc_40_p;
  wire ffc_40_n;
  wire ffc_41_p;
  wire ffc_41_n;
  wire ffc_42_p;
  wire ffc_42_n;
  wire ffc_43_p;
  wire ffc_43_n;
  wire ffc_44_p;
  wire ffc_44_n;
  wire ffc_45_p;
  wire ffc_45_n;
  wire ffc_46_p;
  wire ffc_46_n;
  wire ffc_47_p;
  wire ffc_47_n;
  wire ffc_48_p;
  wire ffc_48_n;
  wire ffc_49_p;
  wire ffc_49_n;
  wire ffc_50_p;
  wire ffc_50_n;
  wire ffc_51_p;
  wire ffc_51_n;
  wire ffc_52_p;
  wire ffc_52_n;
  wire ffc_53_p;
  wire ffc_53_n;
  wire ffc_54_p;
  wire ffc_54_n;
  wire ffc_55_p;
  wire ffc_55_n;
  wire ffc_56_p;
  wire ffc_56_n;
  wire ffc_57_p;
  wire ffc_57_n;
  wire ffc_58_p;
  wire ffc_58_n;
  wire ffc_59_p;
  wire ffc_59_n;
  wire ffc_60_p;
  wire ffc_60_n;
  wire ffc_61_p;
  wire ffc_61_n;
  wire ffc_62_p;
  wire ffc_62_n;
  wire ffc_63_p;
  wire ffc_63_n;
  wire ffc_64_p;
  wire ffc_64_n;
  wire ffc_65_p;
  wire ffc_65_n;
  wire ffc_66_p;
  wire ffc_66_n;
  wire ffc_67_p;
  wire ffc_67_n;
  wire ffc_68_p;
  wire ffc_68_n;
  wire ffc_69_p;
  wire ffc_69_n;
  wire ffc_70_p;
  wire ffc_70_n;
  wire ffc_71_p;
  wire ffc_71_n;
  wire ffc_72_p;
  wire ffc_72_n;
  wire ffc_73_p;
  wire ffc_73_n;
  wire ffc_74_p;
  wire ffc_74_n;
  wire ffc_75_p;
  wire ffc_75_n;
  wire ffc_76_p;
  wire ffc_76_n;
  wire ffc_77_p;
  wire ffc_77_n;
  wire ffc_78_p;
  wire ffc_78_n;
  wire ffc_79_p;
  wire ffc_79_n;
  wire ffc_80_p;
  wire ffc_80_n;
  wire ffc_81_p;
  wire ffc_81_n;
  wire ffc_82_p;
  wire ffc_82_n;
  wire ffc_83_p;
  wire ffc_83_n;
  wire ffc_84_p;
  wire ffc_84_n;
  wire ffc_85_p;
  wire ffc_85_n;
  wire ffc_86_p;
  wire ffc_86_n;
  wire ffc_87_p;
  wire ffc_87_n;
  wire ffc_88_p;
  wire ffc_88_n;
  wire ffc_89_p;
  wire ffc_89_n;
  wire ffc_90_p;
  wire ffc_90_n;
  wire ffc_91_p;
  wire ffc_91_n;
  wire ffc_92_p;
  wire ffc_92_n;
  wire ffc_93_p;
  wire ffc_93_n;
  wire ffc_94_p;
  wire ffc_94_n;
  wire ffc_95_p;
  wire ffc_95_n;
  wire ffc_96_p;
  wire ffc_96_n;
  wire ffc_97_p;
  wire ffc_97_n;
  wire ffc_98_p;
  wire ffc_98_n;
  wire ffc_99_p;
  wire ffc_99_n;
  wire ffc_100_p;
  wire ffc_100_n;
  wire ffc_101_p;
  wire ffc_101_n;
  wire ffc_102_p;
  wire ffc_102_n;
  wire ffc_103_p;
  wire ffc_103_n;
  wire ffc_104_p;
  wire ffc_104_n;
  wire ffc_105_p;
  wire ffc_105_n;
  wire ffc_106_p;
  wire ffc_106_n;
  wire ffc_107_p;
  wire ffc_107_n;
  wire ffc_108_p;
  wire ffc_108_n;
  wire ffc_109_p;
  wire ffc_109_n;
  wire ffc_110_p;
  wire ffc_110_n;
  wire ffc_111_p;
  wire ffc_111_n;
  wire ffc_112_p;
  wire ffc_112_n;
  wire ffc_113_p;
  wire ffc_113_n;
  wire ffc_114_p;
  wire ffc_114_n;
  wire ffc_115_p;
  wire ffc_115_n;
  wire ffc_116_p;
  wire ffc_116_n;
  wire ffc_117_p;
  wire ffc_117_n;
  wire ffc_118_p;
  wire ffc_118_n;
  wire ffc_119_p;
  wire ffc_119_n;
  wire ffc_120_p;
  wire ffc_120_n;
  wire ffc_121_p;
  wire ffc_121_n;
  wire ffc_122_p;
  wire ffc_122_n;
  wire ffc_123_p;
  wire ffc_123_n;
  wire ffc_124_p;
  wire ffc_124_n;
  wire ffc_125_p;
  wire ffc_125_n;
  wire ffc_126_p;
  wire ffc_126_n;
  wire ffc_127_p;
  wire ffc_127_n;
  wire ffc_128_p;
  wire ffc_128_n;
  wire ffc_129_p;
  wire ffc_129_n;
  wire ffc_130_p;
  wire ffc_130_n;
  wire ffc_131_p;
  wire ffc_131_n;
  wire ffc_132_p;
  wire ffc_132_n;
  wire ffc_133_p;
  wire ffc_133_n;
  wire ffc_134_p;
  wire ffc_134_n;
  wire ffc_135_p;
  wire ffc_135_n;
  wire ffc_136_p;
  wire ffc_136_n;
  wire ffc_137_p;
  wire ffc_137_n;
  wire ffc_138_p;
  wire ffc_138_n;
  wire ffc_139_p;
  wire ffc_139_n;
  wire ffc_140_p;
  wire ffc_140_n;
  wire ffc_141_p;
  wire ffc_141_n;
  wire ffc_142_p;
  wire ffc_142_n;
  wire ffc_143_p;
  wire ffc_143_n;
  wire ffc_144_p;
  wire ffc_144_n;
  wire ffc_145_p;
  wire ffc_145_n;
  wire ffc_146_p;
  wire ffc_146_n;
  wire ffc_147_p;
  wire ffc_147_n;
  wire ffc_148_p;
  wire ffc_148_n;
  wire ffc_149_p;
  wire ffc_149_n;
  wire ffc_150_p;
  wire ffc_150_n;
  wire ffc_151_p;
  wire ffc_151_n;
  wire ffc_152_p;
  wire ffc_152_n;
  wire ffc_153_p;
  wire ffc_153_n;
  wire ffc_154_p;
  wire ffc_154_n;
  wire ffc_155_p;
  wire ffc_155_n;
  wire ffc_156_p;
  wire ffc_156_n;
  wire ffc_157_p;
  wire ffc_157_n;
  wire ffc_158_p;
  wire ffc_158_n;
  wire ffc_159_p;
  wire ffc_159_n;
  wire ffc_160_p;
  wire ffc_160_n;
  wire ffc_161_p;
  wire ffc_161_n;
  wire ffc_162_p;
  wire ffc_162_n;
  wire ffc_163_p;
  wire ffc_163_n;
  wire ffc_164_p;
  wire ffc_164_n;
  wire ffc_165_p;
  wire ffc_165_n;
  wire ffc_166_p;
  wire ffc_166_n;
  wire ffc_167_p;
  wire ffc_167_n;
  wire ffc_168_p;
  wire ffc_168_n;
  wire ffc_169_p;
  wire ffc_169_n;
  wire ffc_170_p;
  wire ffc_170_n;
  wire ffc_171_p;
  wire ffc_171_n;
  wire ffc_172_p;
  wire ffc_172_n;
  wire ffc_173_p;
  wire ffc_173_n;
  wire ffc_174_p;
  wire ffc_174_n;
  wire ffc_175_p;
  wire ffc_175_n;
  wire ffc_176_p;
  wire ffc_176_n;
  wire ffc_177_p;
  wire ffc_177_n;
  wire ffc_178_p;
  wire ffc_178_n;
  wire ffc_179_p;
  wire ffc_179_n;
  wire ffc_180_p;
  wire ffc_180_n;
  wire ffc_181_p;
  wire ffc_181_n;
  wire ffc_182_p;
  wire ffc_182_n;
  wire ffc_183_p;
  wire ffc_183_n;
  wire ffc_184_p;
  wire ffc_184_n;
  wire ffc_185_p;
  wire ffc_185_n;
  wire ffc_186_p;
  wire ffc_186_n;
  wire ffc_187_p;
  wire ffc_187_n;
  wire ffc_188_p;
  wire ffc_188_n;
  wire ffc_189_p;
  wire ffc_189_n;
  wire ffc_190_p;
  wire ffc_190_n;
  wire ffc_191_p;
  wire ffc_191_n;
  wire ffc_192_p;
  wire ffc_192_n;
  wire ffc_193_p;
  wire ffc_193_n;
  wire ffc_194_p;
  wire ffc_194_n;
  wire ffc_195_p;
  wire ffc_195_n;
  wire ffc_196_p;
  wire ffc_196_n;
  wire ffc_197_p;
  wire ffc_197_n;
  wire ffc_198_p;
  wire ffc_198_n;
  wire ffc_199_p;
  wire ffc_199_n;
  wire ffc_200_p;
  wire ffc_200_n;
  wire ffc_201_p;
  wire ffc_201_n;
  wire ffc_202_p;
  wire ffc_202_n;
  wire ffc_203_p;
  wire ffc_203_n;
  wire ffc_204_p;
  wire ffc_204_n;
  wire ffc_205_p;
  wire ffc_205_n;
  wire ffc_206_p;
  wire ffc_206_n;
  wire ffc_207_p;
  wire ffc_207_n;
  wire ffc_208_p;
  wire ffc_208_n;
  wire ffc_209_p;
  wire ffc_209_n;
  wire ffc_210_p;
  wire ffc_210_n;
  wire ffc_211_p;
  wire ffc_211_n;
  wire ffc_212_p;
  wire ffc_212_n;
  wire ffc_213_p;
  wire ffc_213_n;
  wire ffc_214_p;
  wire ffc_214_n;
  wire ffc_215_p;
  wire ffc_215_n;
  wire ffc_216_p;
  wire ffc_216_n;
  wire ffc_217_p;
  wire ffc_217_n;
  wire ffc_218_p;
  wire ffc_218_n;
  wire ffc_219_p;
  wire ffc_219_n;
  wire ffc_220_p;
  wire ffc_220_n;
  wire ffc_221_p;
  wire ffc_221_n;
  wire ffc_222_p;
  wire ffc_222_n;
  wire ffc_223_p;
  wire ffc_223_n;
  wire ffc_224_p;
  wire ffc_224_n;
  wire ffc_225_p;
  wire ffc_225_n;
  wire ffc_226_p;
  wire ffc_226_n;
  wire ffc_227_p;
  wire ffc_227_n;
  wire ffc_228_p;
  wire ffc_228_n;
  wire ffc_229_p;
  wire ffc_229_n;
  wire ffc_230_p;
  wire ffc_230_n;
  wire ffc_231_p;
  wire ffc_231_n;
  wire ffc_232_p;
  wire ffc_232_n;
  wire ffc_233_p;
  wire ffc_233_n;
  wire ffc_234_p;
  wire ffc_234_n;
  wire ffc_235_p;
  wire ffc_235_n;
  wire ffc_236_p;
  wire ffc_236_n;
  wire ffc_237_p;
  wire ffc_237_n;
  wire ffc_238_p;
  wire ffc_238_n;
  wire ffc_239_p;
  wire ffc_239_n;
  wire ffc_240_p;
  wire ffc_240_n;
  wire ffc_241_p;
  wire ffc_241_n;
  wire ffc_242_p;
  wire ffc_242_n;
  wire ffc_243_p;
  wire ffc_243_n;
  wire ffc_244_p;
  wire ffc_244_n;
  wire ffc_245_p;
  wire ffc_245_n;
  wire ffc_246_p;
  wire ffc_246_n;
  wire ffc_247_p;
  wire ffc_247_n;
  wire ffc_248_p;
  wire ffc_248_n;
  wire ffc_249_p;
  wire ffc_249_n;
  wire ffc_250_p;
  wire ffc_250_n;
  wire ffc_251_p;
  wire ffc_251_n;
  wire ffc_252_p;
  wire ffc_252_n;
  wire ffc_253_p;
  wire ffc_253_n;
  wire ffc_254_p;
  wire ffc_254_n;
  wire ffc_255_p;
  wire ffc_255_n;
  wire ffc_256_p;
  wire ffc_256_n;
  wire ffc_257_p;
  wire ffc_257_n;
  wire ffc_258_p;
  wire ffc_258_n;
  wire ffc_259_p;
  wire ffc_259_n;
  wire ffc_260_p;
  wire ffc_260_n;
  wire ffc_261_p;
  wire ffc_261_n;
  wire ffc_262_p;
  wire ffc_262_n;
  wire ffc_263_p;
  wire ffc_263_n;
  wire ffc_264_p;
  wire ffc_264_n;
  wire ffc_265_p;
  wire ffc_265_n;
  wire ffc_266_p;
  wire ffc_266_n;
  wire ffc_267_p;
  wire ffc_267_n;
  wire ffc_268_p;
  wire ffc_268_n;
  wire ffc_269_p;
  wire ffc_269_n;
  wire ffc_270_p;
  wire ffc_270_n;
  wire ffc_271_p;
  wire ffc_271_n;
  wire ffc_272_p;
  wire ffc_272_n;
  wire ffc_273_p;
  wire ffc_273_n;
  wire ffc_274_p;
  wire ffc_274_n;
  wire ffc_275_p;
  wire ffc_275_n;
  wire ffc_276_p;
  wire ffc_276_n;
  wire ffc_277_p;
  wire ffc_277_n;
  wire ffc_278_p;
  wire ffc_278_n;
  wire ffc_279_p;
  wire ffc_279_n;
  wire ffc_280_p;
  wire ffc_280_n;
  wire ffc_281_p;
  wire ffc_281_n;
  wire ffc_282_p;
  wire ffc_282_n;
  wire ffc_283_p;
  wire ffc_283_n;
  wire ffc_284_p;
  wire ffc_284_n;
  wire ffc_285_p;
  wire ffc_285_n;
  wire ffc_286_p;
  wire ffc_286_n;
  wire ffc_287_p;
  wire ffc_287_n;
  wire ffc_288_p;
  wire ffc_288_n;
  wire ffc_289_p;
  wire ffc_289_n;
  wire ffc_290_p;
  wire ffc_290_n;
  wire ffc_291_p;
  wire ffc_291_n;
  wire ffc_292_p;
  wire ffc_292_n;
  wire ffc_293_p;
  wire ffc_293_n;
  wire ffc_294_p;
  wire ffc_294_n;
  wire ffc_295_p;
  wire ffc_295_n;
  wire ffc_296_p;
  wire ffc_296_n;
  wire ffc_297_p;
  wire ffc_297_n;
  wire ffc_298_p;
  wire ffc_298_n;
  wire ffc_299_p;
  wire ffc_299_n;
  wire ffc_300_p;
  wire ffc_300_n;
  wire ffc_301_p;
  wire ffc_301_n;
  wire ffc_302_p;
  wire ffc_302_n;
  wire ffc_303_p;
  wire ffc_303_n;
  wire ffc_304_p;
  wire ffc_304_n;
  wire ffc_305_p;
  wire ffc_305_n;
  wire ffc_306_p;
  wire ffc_306_n;
  wire ffc_307_p;
  wire ffc_307_n;
  wire ffc_308_p;
  wire ffc_308_n;
  wire ffc_309_p;
  wire ffc_309_n;
  wire ffc_310_p;
  wire ffc_310_n;
  wire ffc_311_p;
  wire ffc_311_n;
  wire ffc_312_p;
  wire ffc_312_n;
  wire ffc_313_p;
  wire ffc_313_n;
  wire ffc_314_p;
  wire ffc_314_n;
  wire ffc_315_p;
  wire ffc_315_n;
  wire ffc_316_p;
  wire ffc_316_n;
  wire ffc_317_p;
  wire ffc_317_n;
  wire ffc_318_p;
  wire ffc_318_n;
  wire ffc_319_p;
  wire ffc_319_n;
  wire ffc_320_p;
  wire ffc_320_n;
  wire ffc_321_p;
  wire ffc_321_n;
  wire ffc_322_p;
  wire ffc_322_n;
  wire ffc_323_p;
  wire ffc_323_n;
  wire ffc_324_p;
  wire ffc_324_n;
  wire ffc_325_p;
  wire ffc_325_n;
  wire ffc_326_p;
  wire ffc_326_n;
  wire ffc_327_p;
  wire ffc_327_n;
  wire ffc_328_p;
  wire ffc_328_n;
  wire ffc_329_p;
  wire ffc_329_n;
  wire ffc_330_p;
  wire ffc_330_n;
  wire ffc_331_p;
  wire ffc_331_n;
  wire ffc_332_p;
  wire ffc_332_n;
  wire ffc_333_p;
  wire ffc_333_n;
  wire ffc_334_p;
  wire ffc_334_n;
  wire ffc_335_p;
  wire ffc_335_n;
  wire ffc_336_p;
  wire ffc_336_n;
  wire ffc_337_p;
  wire ffc_337_n;
  wire ffc_338_p;
  wire ffc_338_n;
  wire ffc_339_p;
  wire ffc_339_n;
  wire ffc_340_p;
  wire ffc_340_n;
  wire ffc_341_p;
  wire ffc_341_n;
  wire ffc_342_p;
  wire ffc_342_n;
  wire ffc_343_p;
  wire ffc_343_n;
  wire ffc_344_p;
  wire ffc_344_n;
  wire ffc_345_p;
  wire ffc_345_n;
  wire ffc_346_p;
  wire ffc_346_n;
  wire ffc_347_p;
  wire ffc_347_n;
  wire ffc_348_p;
  wire ffc_348_n;
  wire ffc_349_p;
  wire ffc_349_n;
  wire ffc_350_p;
  wire ffc_350_n;
  wire ffc_351_p;
  wire ffc_351_n;
  wire ffc_352_p;
  wire ffc_352_n;
  wire ffc_353_p;
  wire ffc_353_n;
  wire ffc_354_p;
  wire ffc_354_n;
  wire ffc_355_p;
  wire ffc_355_n;
  wire ffc_356_p;
  wire ffc_356_n;
  wire ffc_357_p;
  wire ffc_357_n;
  wire ffc_358_p;
  wire ffc_358_n;
  wire ffc_359_p;
  wire ffc_359_n;
  wire ffc_360_p;
  wire ffc_360_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire g693_p;
  wire g693_n;
  wire g694_p;
  wire g694_n;
  wire g695_p;
  wire g695_n;
  wire g696_p;
  wire g696_n;
  wire g697_p;
  wire g697_n;
  wire g698_p;
  wire g698_n;
  wire g699_p;
  wire g699_n;
  wire g700_p;
  wire g700_n;
  wire g701_p;
  wire g701_n;
  wire g702_p;
  wire g702_n;
  wire g703_p;
  wire g703_n;
  wire g704_p;
  wire g704_n;
  wire g705_p;
  wire g705_n;
  wire g706_p;
  wire g706_n;
  wire g707_p;
  wire g707_n;
  wire g708_p;
  wire g708_n;
  wire g709_p;
  wire g709_n;
  wire g710_p;
  wire g710_n;
  wire g711_p;
  wire g711_n;
  wire g712_p;
  wire g712_n;
  wire g713_p;
  wire g713_n;
  wire g714_p;
  wire g714_n;
  wire g715_p;
  wire g715_n;
  wire g716_p;
  wire g716_n;
  wire g717_p;
  wire g717_n;
  wire g718_p;
  wire g718_n;
  wire g719_p;
  wire g719_n;
  wire g720_p;
  wire g720_n;
  wire g721_p;
  wire g721_n;
  wire g722_p;
  wire g722_n;
  wire g723_p;
  wire g723_n;
  wire g724_p;
  wire g724_n;
  wire g725_p;
  wire g725_n;
  wire g726_p;
  wire g726_n;
  wire g727_p;
  wire g727_n;
  wire g728_p;
  wire g728_n;
  wire g729_p;
  wire g729_n;
  wire g730_p;
  wire g730_n;
  wire g731_p;
  wire g731_n;
  wire g732_p;
  wire g732_n;
  wire g733_p;
  wire g733_n;
  wire g734_p;
  wire g734_n;
  wire g735_p;
  wire g735_n;
  wire g736_p;
  wire g736_n;
  wire g737_p;
  wire g737_n;
  wire g738_p;
  wire g738_n;
  wire g739_p;
  wire g739_n;
  wire g740_p;
  wire g740_n;
  wire g741_p;
  wire g741_n;
  wire g742_p;
  wire g742_n;
  wire g743_p;
  wire g743_n;
  wire g744_p;
  wire g744_n;
  wire g745_p;
  wire g745_n;
  wire g746_p;
  wire g746_n;
  wire g747_p;
  wire g747_n;
  wire g748_p;
  wire g748_n;
  wire g749_p;
  wire g749_n;
  wire g750_p;
  wire g750_n;
  wire g751_p;
  wire g751_n;
  wire g752_p;
  wire g752_n;
  wire g753_p;
  wire g753_n;
  wire g754_p;
  wire g754_n;
  wire g755_p;
  wire g755_n;
  wire g756_p;
  wire g756_n;
  wire g757_p;
  wire g757_n;
  wire g758_p;
  wire g758_n;
  wire g759_p;
  wire g759_n;
  wire g760_p;
  wire g760_n;
  wire g761_p;
  wire g761_n;
  wire g762_p;
  wire g762_n;
  wire g763_p;
  wire g763_n;
  wire g764_p;
  wire g764_n;
  wire g765_p;
  wire g765_n;
  wire g766_p;
  wire g766_n;
  wire g767_p;
  wire g767_n;
  wire g768_p;
  wire g768_n;
  wire g769_p;
  wire g769_n;
  wire g770_p;
  wire g770_n;
  wire g771_p;
  wire g771_n;
  wire g772_p;
  wire g772_n;
  wire g773_p;
  wire g773_n;
  wire g774_p;
  wire g774_n;
  wire g775_p;
  wire g775_n;
  wire g776_p;
  wire g776_n;
  wire g777_p;
  wire g777_n;
  wire g778_p;
  wire g778_n;
  wire g779_p;
  wire g779_n;
  wire g780_p;
  wire g780_n;
  wire g781_p;
  wire g781_n;
  wire g782_p;
  wire g782_n;
  wire g783_p;
  wire g783_n;
  wire g784_p;
  wire g784_n;
  wire g785_p;
  wire g785_n;
  wire g786_p;
  wire g786_n;
  wire g787_p;
  wire g787_n;
  wire g788_p;
  wire g788_n;
  wire g789_p;
  wire g789_n;
  wire g790_p;
  wire g790_n;
  wire g791_p;
  wire g791_n;
  wire g792_p;
  wire g792_n;
  wire g793_p;
  wire g793_n;
  wire g794_p;
  wire g794_n;
  wire g795_p;
  wire g795_n;
  wire g796_p;
  wire g796_n;
  wire g797_p;
  wire g797_n;
  wire g798_p;
  wire g798_n;
  wire g799_p;
  wire g799_n;
  wire g800_p;
  wire g800_n;
  wire g801_p;
  wire g801_n;
  wire g802_p;
  wire g802_n;
  wire g803_p;
  wire g803_n;
  wire g804_p;
  wire g804_n;
  wire g805_p;
  wire g805_n;
  wire g806_p;
  wire g806_n;
  wire g807_p;
  wire g807_n;
  wire g808_p;
  wire g808_n;
  wire g809_p;
  wire g809_n;
  wire g810_p;
  wire g810_n;
  wire g811_p;
  wire g811_n;
  wire g812_p;
  wire g812_n;
  wire g813_p;
  wire g813_n;
  wire g814_p;
  wire g814_n;
  wire g815_p;
  wire g815_n;
  wire g816_p;
  wire g816_n;
  wire g817_p;
  wire g817_n;
  wire g818_p;
  wire g818_n;
  wire g819_p;
  wire g819_n;
  wire g820_p;
  wire g820_n;
  wire g821_p;
  wire g821_n;
  wire g822_p;
  wire g822_n;
  wire g823_p;
  wire g823_n;
  wire g824_p;
  wire g824_n;
  wire g825_p;
  wire g825_n;
  wire g826_p;
  wire g826_n;
  wire g827_p;
  wire g827_n;
  wire g828_p;
  wire g828_n;
  wire g829_p;
  wire g829_n;
  wire g830_p;
  wire g830_n;
  wire g831_p;
  wire g831_n;
  wire g832_p;
  wire g832_n;
  wire g833_p;
  wire g833_n;
  wire g834_p;
  wire g834_n;
  wire g835_p;
  wire g835_n;
  wire g836_p;
  wire g836_n;
  wire g837_p;
  wire g837_n;
  wire g838_p;
  wire g838_n;
  wire g839_p;
  wire g839_n;
  wire g840_p;
  wire g840_n;
  wire g841_p;
  wire g841_n;
  wire g842_p;
  wire g842_n;
  wire g843_p;
  wire g843_n;
  wire g844_p;
  wire g844_n;
  wire g845_p;
  wire g845_n;
  wire g846_p;
  wire g846_n;
  wire g847_p;
  wire g847_n;
  wire g848_p;
  wire g848_n;
  wire g849_p;
  wire g849_n;
  wire g850_p;
  wire g850_n;
  wire g851_p;
  wire g851_n;
  wire g852_p;
  wire g852_n;
  wire g853_p;
  wire g853_n;
  wire g854_p;
  wire g854_n;
  wire g855_p;
  wire g855_n;
  wire g856_p;
  wire g856_n;
  wire g857_p;
  wire g857_n;
  wire g858_p;
  wire g858_n;
  wire g859_p;
  wire g859_n;
  wire g860_p;
  wire g860_n;
  wire g861_p;
  wire g861_n;
  wire g862_p;
  wire g862_n;
  wire g863_p;
  wire g863_n;
  wire g864_p;
  wire g864_n;
  wire g865_p;
  wire g865_n;
  wire g866_p;
  wire g866_n;
  wire g867_p;
  wire g867_n;
  wire g868_p;
  wire g868_n;
  wire g869_p;
  wire g869_n;
  wire g870_p;
  wire g870_n;
  wire g871_p;
  wire g871_n;
  wire g872_p;
  wire g872_n;
  wire g873_p;
  wire g873_n;
  wire g874_p;
  wire g874_n;
  wire g875_p;
  wire g875_n;
  wire g876_p;
  wire g876_n;
  wire g877_p;
  wire g877_n;
  wire g878_p;
  wire g878_n;
  wire g879_p;
  wire g879_n;
  wire g880_p;
  wire g880_n;
  wire g881_p;
  wire g881_n;
  wire g882_p;
  wire g882_n;
  wire g883_p;
  wire g883_n;
  wire g884_p;
  wire g884_n;
  wire g885_p;
  wire g885_n;
  wire g886_p;
  wire g886_n;
  wire g887_p;
  wire g887_n;
  wire g888_p;
  wire g888_n;
  wire g889_p;
  wire g889_n;
  wire g890_p;
  wire g890_n;
  wire g891_p;
  wire g891_n;
  wire g892_p;
  wire g892_n;
  wire g893_p;
  wire g893_n;
  wire g894_p;
  wire g894_n;
  wire g895_p;
  wire g895_n;
  wire g896_p;
  wire g896_n;
  wire g897_p;
  wire g897_n;
  wire g898_p;
  wire g898_n;
  wire g899_p;
  wire g899_n;
  wire g900_p;
  wire g900_n;
  wire g901_p;
  wire g901_n;
  wire g902_p;
  wire g902_n;
  wire g903_p;
  wire g903_n;
  wire g904_p;
  wire g904_n;
  wire g905_p;
  wire g905_n;
  wire g906_p;
  wire g906_n;
  wire g907_p;
  wire g907_n;
  wire g908_p;
  wire g908_n;
  wire g909_p;
  wire g909_n;
  wire g910_p;
  wire g910_n;
  wire g911_p;
  wire g911_n;
  wire g912_p;
  wire g912_n;
  wire g913_p;
  wire g913_n;
  wire g914_p;
  wire g914_n;
  wire g915_p;
  wire g915_n;
  wire g916_p;
  wire g916_n;
  wire g917_p;
  wire g917_n;
  wire g918_p;
  wire g918_n;
  wire g919_p;
  wire g919_n;
  wire g920_p;
  wire g920_n;
  wire g921_p;
  wire g921_n;
  wire g922_p;
  wire g922_n;
  wire g923_p;
  wire g923_n;
  wire g924_p;
  wire g924_n;
  wire g925_p;
  wire g925_n;
  wire g926_p;
  wire g926_n;
  wire g927_p;
  wire g927_n;
  wire g928_p;
  wire g928_n;
  wire g929_p;
  wire g929_n;
  wire g930_p;
  wire g930_n;
  wire g931_p;
  wire g931_n;
  wire g932_p;
  wire g932_n;
  wire g933_p;
  wire g933_n;
  wire g934_p;
  wire g934_n;
  wire g935_p;
  wire g935_n;
  wire g936_p;
  wire g936_n;
  wire g937_p;
  wire g937_n;
  wire g938_p;
  wire g938_n;
  wire g939_p;
  wire g939_n;
  wire g940_p;
  wire g940_n;
  wire g941_p;
  wire g941_n;
  wire g942_p;
  wire g942_n;
  wire g943_p;
  wire g943_n;
  wire g944_p;
  wire g944_n;
  wire g945_p;
  wire g945_n;
  wire g946_p;
  wire g946_n;
  wire g947_p;
  wire g947_n;
  wire g948_p;
  wire g948_n;
  wire g949_p;
  wire g949_n;
  wire g950_p;
  wire g950_n;
  wire g951_p;
  wire g951_n;
  wire g952_p;
  wire g952_n;
  wire g953_p;
  wire g953_n;
  wire g954_p;
  wire g954_n;
  wire g955_p;
  wire g955_n;
  wire g956_p;
  wire g956_n;
  wire g957_p;
  wire g957_n;
  wire g958_p;
  wire g958_n;
  wire g959_p;
  wire g959_n;
  wire g960_p;
  wire g960_n;
  wire g961_p;
  wire g961_n;
  wire g962_p;
  wire g962_n;
  wire g963_p;
  wire g963_n;
  wire g964_p;
  wire g964_n;
  wire g965_p;
  wire g965_n;
  wire g966_p;
  wire g966_n;
  wire g967_p;
  wire g967_n;
  wire g968_p;
  wire g968_n;
  wire g969_p;
  wire g969_n;
  wire g970_p;
  wire g970_n;
  wire g971_p;
  wire g971_n;
  wire g972_p;
  wire g972_n;
  wire g973_p;
  wire g973_n;
  wire g974_p;
  wire g974_n;
  wire g975_p;
  wire g975_n;
  wire g976_p;
  wire g976_n;
  wire g977_p;
  wire g977_n;
  wire g978_p;
  wire g978_n;
  wire g979_p;
  wire g979_n;
  wire g980_p;
  wire g980_n;
  wire g981_p;
  wire g981_n;
  wire g982_p;
  wire g982_n;
  wire g983_p;
  wire g983_n;
  wire g984_p;
  wire g984_n;
  wire g985_p;
  wire g985_n;
  wire g986_p;
  wire g986_n;
  wire g987_p;
  wire g987_n;
  wire g988_p;
  wire g988_n;
  wire g989_p;
  wire g989_n;
  wire g990_p;
  wire g990_n;
  wire g991_p;
  wire g991_n;
  wire g992_p;
  wire g992_n;
  wire g993_p;
  wire g993_n;
  wire g994_p;
  wire g994_n;
  wire g995_p;
  wire g995_n;
  wire g996_p;
  wire g996_n;
  wire g997_p;
  wire g997_n;
  wire g998_p;
  wire g998_n;
  wire g999_p;
  wire g999_n;
  wire g1000_p;
  wire g1000_n;
  wire g1001_p;
  wire g1001_n;
  wire g1002_p;
  wire g1002_n;
  wire g1003_p;
  wire g1003_n;
  wire g1004_p;
  wire g1004_n;
  wire g1005_p;
  wire g1005_n;
  wire g1006_p;
  wire g1006_n;
  wire g1007_p;
  wire g1007_n;
  wire g1008_p;
  wire g1008_n;
  wire g1009_p;
  wire g1009_n;
  wire g1010_p;
  wire g1010_n;
  wire g1011_p;
  wire g1011_n;
  wire g1012_p;
  wire g1012_n;
  wire g1013_p;
  wire g1013_n;
  wire g1014_p;
  wire g1014_n;
  wire g1015_p;
  wire g1015_n;
  wire g1016_p;
  wire g1016_n;
  wire g1017_p;
  wire g1017_n;
  wire g1018_p;
  wire g1018_n;
  wire g1019_p;
  wire g1019_n;
  wire g1020_p;
  wire g1020_n;
  wire g1021_p;
  wire g1021_n;
  wire g1022_p;
  wire g1022_n;
  wire g1023_p;
  wire g1023_n;
  wire g1024_p;
  wire g1024_n;
  wire g1025_p;
  wire g1025_n;
  wire g1026_p;
  wire g1026_n;
  wire g1027_p;
  wire g1027_n;
  wire g1028_p;
  wire g1028_n;
  wire g1029_p;
  wire g1029_n;
  wire g1030_p;
  wire g1030_n;
  wire g1031_p;
  wire g1031_n;
  wire g1032_p;
  wire g1032_n;
  wire g1033_p;
  wire g1033_n;
  wire g1034_p;
  wire g1034_n;
  wire g1035_p;
  wire g1035_n;
  wire g1036_p;
  wire g1036_n;
  wire g1037_p;
  wire g1037_n;
  wire g1038_p;
  wire g1038_n;
  wire g1039_p;
  wire g1039_n;
  wire g1040_p;
  wire g1040_n;
  wire g1041_p;
  wire g1041_n;
  wire g1042_p;
  wire g1042_n;
  wire g1043_p;
  wire g1043_n;
  wire g1044_p;
  wire g1044_n;
  wire g1045_p;
  wire g1045_n;
  wire g1046_p;
  wire g1046_n;
  wire g1047_p;
  wire g1047_n;
  wire g1048_p;
  wire g1048_n;
  wire g1049_p;
  wire g1049_n;
  wire g1050_p;
  wire g1050_n;
  wire g1051_p;
  wire g1051_n;
  wire g1052_p;
  wire g1052_n;
  wire g1053_p;
  wire g1053_n;
  wire g1054_p;
  wire g1054_n;
  wire g1055_p;
  wire g1055_n;
  wire g1056_p;
  wire g1056_n;
  wire g1057_p;
  wire g1057_n;
  wire g1058_p;
  wire g1058_n;
  wire g1059_p;
  wire g1059_n;
  wire g1060_p;
  wire g1060_n;
  wire g1061_p;
  wire g1061_n;
  wire g1062_p;
  wire g1062_n;
  wire g1063_p;
  wire g1063_n;
  wire g1064_p;
  wire g1064_n;
  wire g1065_p;
  wire g1065_n;
  wire g1066_p;
  wire g1066_n;
  wire g1067_p;
  wire g1067_n;
  wire g1068_p;
  wire g1068_n;
  wire g1069_p;
  wire g1069_n;
  wire g1070_p;
  wire g1070_n;
  wire g1071_p;
  wire g1071_n;
  wire g1072_p;
  wire g1072_n;
  wire g1073_p;
  wire g1073_n;
  wire g1074_p;
  wire g1074_n;
  wire g1075_p;
  wire g1075_n;
  wire g1076_p;
  wire g1076_n;
  wire g1077_p;
  wire g1077_n;
  wire g1078_p;
  wire g1078_n;
  wire g1079_p;
  wire g1079_n;
  wire g1080_p;
  wire g1080_n;
  wire g1081_p;
  wire g1081_n;
  wire g1082_p;
  wire g1082_n;
  wire g1083_p;
  wire g1083_n;
  wire g1084_p;
  wire g1084_n;
  wire g1085_p;
  wire g1085_n;
  wire g1086_p;
  wire g1086_n;
  wire g1087_p;
  wire g1087_n;
  wire g1088_p;
  wire g1088_n;
  wire g1089_p;
  wire g1089_n;
  wire g1090_p;
  wire g1090_n;
  wire g1091_p;
  wire g1091_n;
  wire g1092_p;
  wire g1092_n;
  wire g1093_p;
  wire g1093_n;
  wire g1094_p;
  wire g1094_n;
  wire g1095_p;
  wire g1095_n;
  wire g1096_p;
  wire g1096_n;
  wire g1097_p;
  wire g1097_n;
  wire g1098_p;
  wire g1098_n;
  wire g1099_p;
  wire g1099_n;
  wire g1100_p;
  wire g1100_n;
  wire g1101_p;
  wire g1101_n;
  wire g1102_p;
  wire g1102_n;
  wire g1103_p;
  wire g1103_n;
  wire g1104_p;
  wire g1104_n;
  wire g1105_p;
  wire g1105_n;
  wire g1106_p;
  wire g1106_n;
  wire g1107_p;
  wire g1107_n;
  wire g1108_p;
  wire g1108_n;
  wire g1109_p;
  wire g1109_n;
  wire g1110_p;
  wire g1110_n;
  wire g1111_p;
  wire g1111_n;
  wire g1112_p;
  wire g1112_n;
  wire g1113_p;
  wire g1113_n;
  wire g1114_p;
  wire g1114_n;
  wire g1115_p;
  wire g1115_n;
  wire g1116_p;
  wire g1116_n;
  wire g1117_p;
  wire g1117_n;
  wire g1118_p;
  wire g1118_n;
  wire g1119_p;
  wire g1119_n;
  wire g1120_p;
  wire g1120_n;
  wire g1121_p;
  wire g1121_n;
  wire g1122_p;
  wire g1122_n;
  wire g1123_p;
  wire g1123_n;
  wire g1124_p;
  wire g1124_n;
  wire g1125_p;
  wire g1125_n;
  wire g1126_p;
  wire g1126_n;
  wire g1127_p;
  wire g1127_n;
  wire g1128_p;
  wire g1128_n;
  wire g1129_p;
  wire g1129_n;
  wire g1130_p;
  wire g1130_n;
  wire g1131_p;
  wire g1131_n;
  wire g1132_p;
  wire g1132_n;
  wire g1133_p;
  wire g1133_n;
  wire g1134_p;
  wire g1134_n;
  wire g1135_p;
  wire g1135_n;
  wire g1136_p;
  wire g1136_n;
  wire g1137_p;
  wire g1137_n;
  wire g1138_p;
  wire g1138_n;
  wire g1139_p;
  wire g1139_n;
  wire g1140_p;
  wire g1140_n;
  wire g1141_p;
  wire g1141_n;
  wire g1142_p;
  wire g1142_n;
  wire g1143_p;
  wire g1143_n;
  wire g1144_p;
  wire g1144_n;
  wire g1145_p;
  wire g1145_n;
  wire g1146_p;
  wire g1146_n;
  wire g1147_p;
  wire g1147_n;
  wire g1148_p;
  wire g1148_n;
  wire g1149_p;
  wire g1149_n;
  wire g1150_p;
  wire g1150_n;
  wire g1151_p;
  wire g1151_n;
  wire g1152_p;
  wire g1152_n;
  wire g1153_p;
  wire g1153_n;
  wire g1154_p;
  wire g1154_n;
  wire g1155_p;
  wire g1155_n;
  wire g1156_p;
  wire g1156_n;
  wire g1157_p;
  wire g1157_n;
  wire g1158_p;
  wire g1158_n;
  wire g1159_p;
  wire g1159_n;
  wire g1160_p;
  wire g1160_n;
  wire g1161_p;
  wire g1161_n;
  wire g1162_p;
  wire g1162_n;
  wire g1163_p;
  wire g1163_n;
  wire g1164_p;
  wire g1164_n;
  wire g1165_p;
  wire g1165_n;
  wire g1166_p;
  wire g1166_n;
  wire g1167_p;
  wire g1167_n;
  wire g1168_p;
  wire g1168_n;
  wire g1169_p;
  wire g1169_n;
  wire g1170_p;
  wire g1170_n;
  wire g1171_p;
  wire g1171_n;
  wire g1172_p;
  wire g1172_n;
  wire g1173_p;
  wire g1173_n;
  wire g1174_p;
  wire g1174_n;
  wire g1175_p;
  wire g1175_n;
  wire g1176_p;
  wire g1176_n;
  wire g1177_p;
  wire g1177_n;
  wire g1178_p;
  wire g1178_n;
  wire g1179_p;
  wire g1179_n;
  wire g1180_p;
  wire g1180_n;
  wire g1181_p;
  wire g1181_n;
  wire g1182_p;
  wire g1182_n;
  wire g1183_p;
  wire g1183_n;
  wire g1184_p;
  wire g1184_n;
  wire g1185_p;
  wire g1185_n;
  wire g1186_p;
  wire g1186_n;
  wire g1187_p;
  wire g1187_n;
  wire g1188_p;
  wire g1188_n;
  wire g1189_p;
  wire g1189_n;
  wire g1190_p;
  wire g1190_n;
  wire g1191_p;
  wire g1191_n;
  wire g1192_p;
  wire g1192_n;
  wire g1193_p;
  wire g1193_n;
  wire g1194_p;
  wire g1194_n;
  wire g1195_p;
  wire g1195_n;
  wire g1196_p;
  wire g1196_n;
  wire g1197_p;
  wire g1197_n;
  wire g1198_p;
  wire g1198_n;
  wire g1199_p;
  wire g1199_n;
  wire g1200_p;
  wire g1200_n;
  wire g1201_p;
  wire g1201_n;
  wire g1202_p;
  wire g1202_n;
  wire g1203_p;
  wire g1203_n;
  wire g1204_p;
  wire g1204_n;
  wire g1205_p;
  wire g1205_n;
  wire g1206_p;
  wire g1206_n;
  wire g1207_p;
  wire g1207_n;
  wire g1208_p;
  wire g1208_n;
  wire g1209_p;
  wire g1209_n;
  wire g1210_p;
  wire g1210_n;
  wire g1211_p;
  wire g1211_n;
  wire g1212_p;
  wire g1212_n;
  wire g1213_p;
  wire g1213_n;
  wire g1214_p;
  wire g1214_n;
  wire g1215_p;
  wire g1215_n;
  wire g1216_p;
  wire g1216_n;
  wire g1217_p;
  wire g1217_n;
  wire g1218_p;
  wire g1218_n;
  wire g1219_p;
  wire g1219_n;
  wire g1220_p;
  wire g1220_n;
  wire g1221_p;
  wire g1221_n;
  wire g1222_p;
  wire g1222_n;
  wire g1223_p;
  wire g1223_n;
  wire g1224_p;
  wire g1224_n;
  wire g1225_p;
  wire g1225_n;
  wire g1226_p;
  wire g1226_n;
  wire g1227_p;
  wire g1227_n;
  wire g1228_p;
  wire g1228_n;
  wire g1229_p;
  wire g1229_n;
  wire g1230_p;
  wire g1230_n;
  wire g1231_p;
  wire g1231_n;
  wire g1232_p;
  wire g1232_n;
  wire g1233_p;
  wire g1233_n;
  wire g1234_p;
  wire g1234_n;
  wire g1235_p;
  wire g1235_n;
  wire ffc_5_n_spl_;
  wire ffc_0_n_spl_;
  wire ffc_1_n_spl_;
  wire ffc_6_p_spl_;
  wire ffc_32_n_spl_;
  wire ffc_32_n_spl_0;
  wire ffc_32_n_spl_1;
  wire ffc_30_n_spl_;
  wire ffc_30_n_spl_0;
  wire ffc_2_p_spl_;
  wire ffc_28_n_spl_;
  wire ffc_28_n_spl_0;
  wire ffc_31_n_spl_;
  wire ffc_31_n_spl_0;
  wire ffc_9_p_spl_;
  wire ffc_9_p_spl_0;
  wire ffc_35_n_spl_;
  wire ffc_35_n_spl_0;
  wire ffc_29_n_spl_;
  wire ffc_29_n_spl_0;
  wire ffc_7_p_spl_;
  wire ffc_33_n_spl_;
  wire ffc_33_n_spl_0;
  wire ffc_33_n_spl_1;
  wire ffc_8_p_spl_;
  wire ffc_8_p_spl_0;
  wire ffc_34_n_spl_;
  wire ffc_34_n_spl_0;
  wire ffc_34_n_spl_1;
  wire g430_n_spl_;
  wire ffc_34_p_spl_;
  wire ffc_35_p_spl_;
  wire ffc_32_p_spl_;
  wire ffc_33_p_spl_;
  wire g439_n_spl_;
  wire g442_p_spl_;
  wire g439_p_spl_;
  wire g442_n_spl_;
  wire ffc_30_p_spl_;
  wire ffc_31_p_spl_;
  wire ffc_28_p_spl_;
  wire ffc_29_p_spl_;
  wire g448_p_spl_;
  wire g451_n_spl_;
  wire g448_n_spl_;
  wire g451_p_spl_;
  wire ffc_9_n_spl_;
  wire ffc_9_n_spl_0;
  wire ffc_8_n_spl_;
  wire g459_p_spl_;
  wire g462_p_spl_;
  wire g459_n_spl_;
  wire g462_n_spl_;
  wire ffc_79_p_spl_;
  wire ffc_106_n_spl_;
  wire ffc_106_n_spl_0;
  wire ffc_115_n_spl_;
  wire ffc_115_p_spl_;
  wire ffc_90_p_spl_;
  wire g481_n_spl_;
  wire ffc_90_n_spl_;
  wire g481_p_spl_;
  wire ffc_101_p_spl_;
  wire ffc_102_p_spl_;
  wire ffc_101_n_spl_;
  wire ffc_102_n_spl_;
  wire ffc_106_p_spl_;
  wire g480_p_spl_;
  wire g514_p_spl_;
  wire g480_n_spl_;
  wire g480_n_spl_0;
  wire g514_n_spl_;
  wire g514_n_spl_0;
  wire g505_p_spl_;
  wire g511_p_spl_;
  wire g505_n_spl_;
  wire g505_n_spl_0;
  wire g511_n_spl_;
  wire g511_n_spl_0;
  wire g477_p_spl_;
  wire g508_p_spl_;
  wire g477_n_spl_;
  wire g477_n_spl_0;
  wire g508_n_spl_;
  wire g508_n_spl_0;
  wire g516_n_spl_;
  wire g517_n_spl_;
  wire g515_n_spl_;
  wire ffc_233_p_spl_;
  wire ffc_233_p_spl_0;
  wire ffc_25_p_spl_;
  wire g521_n_spl_;
  wire g520_n_spl_;
  wire g526_p_spl_;
  wire g528_n_spl_;
  wire g526_n_spl_;
  wire g528_p_spl_;
  wire ffc_55_p_spl_;
  wire g534_n_spl_;
  wire g534_n_spl_0;
  wire g534_n_spl_1;
  wire ffc_55_n_spl_;
  wire g534_p_spl_;
  wire g534_p_spl_0;
  wire g534_p_spl_1;
  wire g533_p_spl_;
  wire g533_p_spl_0;
  wire g533_p_spl_1;
  wire g538_p_spl_;
  wire g533_n_spl_;
  wire g533_n_spl_0;
  wire g533_n_spl_1;
  wire g538_n_spl_;
  wire g531_n_spl_;
  wire g531_p_spl_;
  wire ffc_103_p_spl_;
  wire ffc_103_p_spl_0;
  wire ffc_103_p_spl_1;
  wire ffc_72_n_spl_;
  wire ffc_235_n_spl_;
  wire ffc_235_n_spl_0;
  wire ffc_235_p_spl_;
  wire ffc_290_p_spl_;
  wire ffc_118_n_spl_;
  wire ffc_118_p_spl_;
  wire ffc_118_p_spl_0;
  wire ffc_71_p_spl_;
  wire ffc_71_n_spl_;
  wire ffc_254_p_spl_;
  wire ffc_67_p_spl_;
  wire g556_p_spl_;
  wire g556_p_spl_0;
  wire g561_p_spl_;
  wire g556_n_spl_;
  wire g556_n_spl_0;
  wire g556_n_spl_1;
  wire g561_n_spl_;
  wire g561_n_spl_0;
  wire g561_n_spl_00;
  wire g561_n_spl_01;
  wire g561_n_spl_1;
  wire ffc_329_p_spl_;
  wire ffc_330_p_spl_;
  wire ffc_329_n_spl_;
  wire ffc_330_n_spl_;
  wire ffc_328_n_spl_;
  wire ffc_328_n_spl_0;
  wire ffc_328_n_spl_00;
  wire ffc_328_n_spl_000;
  wire ffc_328_n_spl_001;
  wire ffc_328_n_spl_01;
  wire ffc_328_n_spl_1;
  wire ffc_328_n_spl_10;
  wire ffc_328_n_spl_11;
  wire ffc_328_p_spl_;
  wire ffc_328_p_spl_0;
  wire ffc_328_p_spl_00;
  wire ffc_328_p_spl_000;
  wire ffc_328_p_spl_001;
  wire ffc_328_p_spl_01;
  wire ffc_328_p_spl_010;
  wire ffc_328_p_spl_011;
  wire ffc_328_p_spl_1;
  wire ffc_328_p_spl_10;
  wire ffc_328_p_spl_11;
  wire g563_p_spl_;
  wire ffc_319_n_spl_;
  wire ffc_319_n_spl_0;
  wire ffc_319_p_spl_;
  wire g568_n_spl_;
  wire g568_n_spl_0;
  wire g569_n_spl_;
  wire g568_p_spl_;
  wire g569_p_spl_;
  wire ffc_320_n_spl_;
  wire ffc_320_n_spl_0;
  wire ffc_320_p_spl_;
  wire g573_n_spl_;
  wire g573_n_spl_0;
  wire g574_n_spl_;
  wire g573_p_spl_;
  wire g574_p_spl_;
  wire ffc_124_p_spl_;
  wire ffc_124_p_spl_0;
  wire ffc_124_p_spl_00;
  wire ffc_124_p_spl_1;
  wire ffc_124_n_spl_;
  wire ffc_124_n_spl_0;
  wire ffc_167_n_spl_;
  wire g579_p_spl_;
  wire g579_p_spl_0;
  wire g579_p_spl_00;
  wire g579_p_spl_01;
  wire g579_p_spl_1;
  wire g578_p_spl_;
  wire g578_p_spl_0;
  wire g578_p_spl_1;
  wire ffc_167_p_spl_;
  wire ffc_297_n_spl_;
  wire ffc_239_p_spl_;
  wire ffc_200_p_spl_;
  wire ffc_240_p_spl_;
  wire g567_p_spl_;
  wire g567_p_spl_0;
  wire g572_p_spl_;
  wire g572_p_spl_0;
  wire ffc_19_p_spl_;
  wire ffc_19_p_spl_0;
  wire ffc_162_n_spl_;
  wire g589_n_spl_;
  wire g578_n_spl_;
  wire g593_n_spl_;
  wire g593_p_spl_;
  wire g579_n_spl_;
  wire g579_n_spl_0;
  wire g579_n_spl_1;
  wire g594_p_spl_;
  wire g594_n_spl_;
  wire g596_p_spl_;
  wire g596_n_spl_;
  wire ffc_275_n_spl_;
  wire ffc_275_p_spl_;
  wire ffc_155_p_spl_;
  wire ffc_155_p_spl_0;
  wire ffc_155_p_spl_1;
  wire ffc_267_p_spl_;
  wire ffc_155_n_spl_;
  wire ffc_155_n_spl_0;
  wire ffc_155_n_spl_1;
  wire g555_p_spl_;
  wire g601_n_spl_;
  wire g601_n_spl_0;
  wire g603_n_spl_;
  wire g601_p_spl_;
  wire g603_p_spl_;
  wire g604_n_spl_;
  wire g600_n_spl_;
  wire g600_n_spl_0;
  wire ffc_70_n_spl_;
  wire ffc_70_n_spl_0;
  wire ffc_70_n_spl_00;
  wire ffc_70_n_spl_01;
  wire ffc_70_n_spl_1;
  wire ffc_70_n_spl_10;
  wire g609_n_spl_;
  wire g609_n_spl_0;
  wire g609_n_spl_1;
  wire ffc_68_p_spl_;
  wire ffc_84_p_spl_;
  wire g612_p_spl_;
  wire g612_p_spl_0;
  wire g612_p_spl_00;
  wire g612_p_spl_01;
  wire g612_p_spl_1;
  wire g612_p_spl_10;
  wire g562_p_spl_;
  wire g562_p_spl_0;
  wire g562_p_spl_00;
  wire g562_p_spl_01;
  wire g562_p_spl_1;
  wire g562_p_spl_10;
  wire g622_n_spl_;
  wire g622_n_spl_0;
  wire g554_n_spl_;
  wire g554_n_spl_0;
  wire g554_p_spl_;
  wire g622_p_spl_;
  wire ffc_333_p_spl_;
  wire ffc_333_p_spl_0;
  wire ffc_333_p_spl_1;
  wire ffc_357_p_spl_;
  wire ffc_357_p_spl_0;
  wire ffc_357_p_spl_00;
  wire ffc_357_p_spl_1;
  wire ffc_312_n_spl_;
  wire ffc_182_n_spl_;
  wire ffc_312_p_spl_;
  wire g648_p_spl_;
  wire g648_p_spl_0;
  wire g648_n_spl_;
  wire g648_n_spl_0;
  wire ffc_181_p_spl_;
  wire ffc_181_n_spl_;
  wire g651_n_spl_;
  wire g651_p_spl_;
  wire ffc_291_n_spl_;
  wire ffc_291_n_spl_0;
  wire g652_n_spl_;
  wire g652_n_spl_0;
  wire g653_n_spl_;
  wire g652_p_spl_;
  wire g653_p_spl_;
  wire ffc_332_p_spl_;
  wire ffc_332_p_spl_0;
  wire ffc_332_p_spl_1;
  wire ffc_335_n_spl_;
  wire ffc_334_p_spl_;
  wire ffc_335_p_spl_;
  wire ffc_335_p_spl_0;
  wire ffc_336_p_spl_;
  wire ffc_337_p_spl_;
  wire ffc_129_n_spl_;
  wire g599_n_spl_;
  wire g599_n_spl_0;
  wire ffc_131_p_spl_;
  wire g597_p_spl_;
  wire g597_p_spl_0;
  wire g598_p_spl_;
  wire ffc_150_n_spl_;
  wire g597_n_spl_;
  wire g597_n_spl_0;
  wire g597_n_spl_1;
  wire ffc_151_p_spl_;
  wire ffc_151_p_spl_0;
  wire ffc_151_p_spl_00;
  wire ffc_151_p_spl_1;
  wire g595_p_spl_;
  wire ffc_17_p_spl_;
  wire ffc_17_p_spl_0;
  wire ffc_197_p_spl_;
  wire ffc_197_p_spl_0;
  wire g592_n_spl_;
  wire g657_n_spl_;
  wire ffc_353_n_spl_;
  wire ffc_245_p_spl_;
  wire ffc_245_p_spl_0;
  wire ffc_245_p_spl_00;
  wire ffc_245_p_spl_1;
  wire g668_n_spl_;
  wire g668_n_spl_0;
  wire g668_n_spl_1;
  wire ffc_245_n_spl_;
  wire ffc_245_n_spl_0;
  wire ffc_245_n_spl_1;
  wire g668_p_spl_;
  wire g668_p_spl_0;
  wire g668_p_spl_1;
  wire ffc_315_n_spl_;
  wire ffc_315_n_spl_0;
  wire ffc_315_n_spl_1;
  wire ffc_315_p_spl_;
  wire ffc_315_p_spl_0;
  wire ffc_315_p_spl_00;
  wire ffc_315_p_spl_01;
  wire ffc_315_p_spl_1;
  wire ffc_315_p_spl_10;
  wire ffc_339_n_spl_;
  wire ffc_339_n_spl_0;
  wire ffc_339_n_spl_1;
  wire ffc_357_n_spl_;
  wire ffc_357_n_spl_0;
  wire ffc_357_n_spl_1;
  wire ffc_339_p_spl_;
  wire ffc_339_p_spl_0;
  wire ffc_323_p_spl_;
  wire ffc_323_p_spl_0;
  wire ffc_323_p_spl_00;
  wire ffc_323_p_spl_000;
  wire ffc_323_p_spl_01;
  wire ffc_323_p_spl_1;
  wire ffc_323_p_spl_10;
  wire ffc_323_p_spl_11;
  wire ffc_323_n_spl_;
  wire ffc_323_n_spl_0;
  wire ffc_323_n_spl_00;
  wire ffc_323_n_spl_1;
  wire ffc_246_p_spl_;
  wire ffc_246_p_spl_0;
  wire ffc_246_p_spl_1;
  wire ffc_246_n_spl_;
  wire ffc_246_n_spl_0;
  wire ffc_246_n_spl_1;
  wire ffc_340_n_spl_;
  wire ffc_340_n_spl_0;
  wire ffc_340_n_spl_1;
  wire ffc_358_p_spl_;
  wire ffc_358_p_spl_0;
  wire ffc_358_p_spl_00;
  wire ffc_358_p_spl_1;
  wire ffc_358_n_spl_;
  wire ffc_333_n_spl_;
  wire ffc_333_n_spl_0;
  wire ffc_333_n_spl_1;
  wire g646_n_spl_;
  wire ffc_201_p_spl_;
  wire ffc_201_p_spl_0;
  wire ffc_201_p_spl_1;
  wire ffc_242_p_spl_;
  wire ffc_348_n_spl_;
  wire ffc_348_n_spl_0;
  wire ffc_348_n_spl_00;
  wire ffc_348_n_spl_01;
  wire ffc_348_n_spl_1;
  wire ffc_348_n_spl_10;
  wire ffc_348_p_spl_;
  wire ffc_348_p_spl_0;
  wire ffc_348_p_spl_00;
  wire ffc_348_p_spl_01;
  wire ffc_348_p_spl_1;
  wire ffc_348_p_spl_10;
  wire ffc_244_p_spl_;
  wire ffc_301_p_spl_;
  wire g688_p_spl_;
  wire g688_p_spl_0;
  wire g690_p_spl_;
  wire g690_p_spl_0;
  wire g688_n_spl_;
  wire g688_n_spl_0;
  wire g690_n_spl_;
  wire g690_n_spl_0;
  wire ffc_202_p_spl_;
  wire ffc_202_p_spl_0;
  wire ffc_202_p_spl_00;
  wire ffc_202_p_spl_1;
  wire ffc_202_n_spl_;
  wire g692_n_spl_;
  wire g692_p_spl_;
  wire g692_p_spl_0;
  wire ffc_247_n_spl_;
  wire ffc_247_n_spl_0;
  wire g693_n_spl_;
  wire ffc_247_p_spl_;
  wire ffc_247_p_spl_0;
  wire ffc_248_p_spl_;
  wire ffc_248_p_spl_0;
  wire ffc_248_p_spl_1;
  wire ffc_314_p_spl_;
  wire ffc_314_p_spl_0;
  wire ffc_248_n_spl_;
  wire ffc_248_n_spl_0;
  wire ffc_314_n_spl_;
  wire g658_p_spl_;
  wire g658_p_spl_0;
  wire g658_p_spl_1;
  wire g705_n_spl_;
  wire ffc_324_n_spl_;
  wire ffc_324_n_spl_0;
  wire ffc_324_p_spl_;
  wire ffc_324_p_spl_0;
  wire g708_n_spl_;
  wire g708_n_spl_0;
  wire g708_p_spl_;
  wire g708_p_spl_0;
  wire g711_n_spl_;
  wire ffc_148_n_spl_;
  wire ffc_127_p_spl_;
  wire ffc_127_p_spl_0;
  wire g661_n_spl_;
  wire ffc_236_n_spl_;
  wire g717_n_spl_;
  wire g717_n_spl_0;
  wire g717_n_spl_1;
  wire ffc_150_p_spl_;
  wire ffc_150_p_spl_0;
  wire ffc_150_p_spl_1;
  wire g599_p_spl_;
  wire ffc_236_p_spl_;
  wire ffc_289_p_spl_;
  wire ffc_289_n_spl_;
  wire g722_n_spl_;
  wire g724_n_spl_;
  wire g722_p_spl_;
  wire g722_p_spl_0;
  wire g724_p_spl_;
  wire ffc_120_n_spl_;
  wire ffc_264_n_spl_;
  wire ffc_120_p_spl_;
  wire ffc_264_p_spl_;
  wire g553_n_spl_;
  wire g731_n_spl_;
  wire g553_p_spl_;
  wire g553_p_spl_0;
  wire g731_p_spl_;
  wire g730_p_spl_;
  wire g730_p_spl_0;
  wire g730_p_spl_1;
  wire g732_p_spl_;
  wire g730_n_spl_;
  wire g730_n_spl_0;
  wire g730_n_spl_00;
  wire g730_n_spl_1;
  wire g732_n_spl_;
  wire g727_p_spl_;
  wire g735_p_spl_;
  wire ffc_171_p_spl_;
  wire ffc_171_p_spl_0;
  wire ffc_171_p_spl_1;
  wire g727_n_spl_;
  wire g727_n_spl_0;
  wire g735_n_spl_;
  wire ffc_70_p_spl_;
  wire ffc_70_p_spl_0;
  wire ffc_70_p_spl_00;
  wire ffc_70_p_spl_01;
  wire ffc_70_p_spl_1;
  wire ffc_70_p_spl_10;
  wire ffc_75_n_spl_;
  wire ffc_75_n_spl_0;
  wire ffc_75_n_spl_1;
  wire g559_n_spl_;
  wire g551_n_spl_;
  wire g552_n_spl_;
  wire g612_n_spl_;
  wire ffc_174_p_spl_;
  wire ffc_174_p_spl_0;
  wire ffc_174_p_spl_00;
  wire ffc_174_p_spl_1;
  wire ffc_159_n_spl_;
  wire ffc_159_n_spl_0;
  wire ffc_159_n_spl_1;
  wire ffc_173_p_spl_;
  wire ffc_173_p_spl_0;
  wire ffc_173_p_spl_1;
  wire ffc_89_n_spl_;
  wire ffc_175_p_spl_;
  wire ffc_175_p_spl_0;
  wire ffc_158_p_spl_;
  wire ffc_158_p_spl_0;
  wire ffc_158_p_spl_1;
  wire ffc_83_n_spl_;
  wire ffc_172_n_spl_;
  wire ffc_172_n_spl_0;
  wire g760_p_spl_;
  wire ffc_104_p_spl_;
  wire ffc_104_p_spl_0;
  wire ffc_73_p_spl_;
  wire g771_n_spl_;
  wire g562_n_spl_;
  wire ffc_75_p_spl_;
  wire ffc_72_p_spl_;
  wire ffc_74_p_spl_;
  wire ffc_74_n_spl_;
  wire ffc_172_p_spl_;
  wire ffc_172_p_spl_0;
  wire ffc_172_p_spl_00;
  wire ffc_172_p_spl_1;
  wire ffc_158_n_spl_;
  wire ffc_158_n_spl_0;
  wire ffc_158_n_spl_00;
  wire ffc_158_n_spl_01;
  wire ffc_158_n_spl_1;
  wire ffc_158_n_spl_10;
  wire ffc_78_p_spl_;
  wire ffc_78_p_spl_0;
  wire ffc_78_p_spl_1;
  wire ffc_204_p_spl_;
  wire ffc_174_n_spl_;
  wire ffc_174_n_spl_0;
  wire ffc_174_n_spl_00;
  wire ffc_174_n_spl_000;
  wire ffc_174_n_spl_01;
  wire ffc_174_n_spl_1;
  wire ffc_174_n_spl_10;
  wire ffc_174_n_spl_11;
  wire ffc_73_n_spl_;
  wire ffc_83_p_spl_;
  wire ffc_83_p_spl_0;
  wire ffc_173_n_spl_;
  wire ffc_173_n_spl_0;
  wire ffc_173_n_spl_00;
  wire ffc_173_n_spl_01;
  wire ffc_173_n_spl_1;
  wire ffc_175_n_spl_;
  wire ffc_175_n_spl_0;
  wire ffc_175_n_spl_00;
  wire ffc_175_n_spl_01;
  wire ffc_175_n_spl_1;
  wire ffc_175_n_spl_10;
  wire ffc_89_p_spl_;
  wire ffc_159_p_spl_;
  wire ffc_159_p_spl_0;
  wire ffc_159_p_spl_00;
  wire ffc_159_p_spl_01;
  wire ffc_159_p_spl_1;
  wire ffc_159_p_spl_10;
  wire ffc_112_p_spl_;
  wire ffc_112_p_spl_0;
  wire g849_p_spl_;
  wire g848_n_spl_;
  wire ffc_113_p_spl_;
  wire ffc_113_p_spl_0;
  wire ffc_262_n_spl_;
  wire ffc_103_n_spl_;
  wire ffc_122_p_spl_;
  wire ffc_122_n_spl_;
  wire ffc_119_n_spl_;
  wire g870_n_spl_;
  wire ffc_119_p_spl_;
  wire g870_p_spl_;
  wire g873_n_spl_;
  wire g873_n_spl_0;
  wire g687_n_spl_;
  wire g878_n_spl_;
  wire g877_p_spl_;
  wire g877_p_spl_0;
  wire g883_n_spl_;
  wire g883_n_spl_0;
  wire g883_n_spl_1;
  wire g884_n_spl_;
  wire g885_n_spl_;
  wire ffc_171_n_spl_;
  wire ffc_171_n_spl_0;
  wire g888_n_spl_;
  wire g577_n_spl_;
  wire g577_n_spl_0;
  wire g656_n_spl_;
  wire ffc_252_p_spl_;
  wire ffc_130_p_spl_;
  wire ffc_163_p_spl_;
  wire ffc_163_p_spl_0;
  wire g960_p_spl_;
  wire g873_p_spl_;
  wire g960_n_spl_;
  wire g621_n_spl_;
  wire g621_n_spl_0;
  wire g645_n_spl_;
  wire g645_n_spl_0;
  wire ffc_251_p_spl_;
  wire ffc_326_p_spl_;
  wire g990_n_spl_;
  wire g659_n_spl_;
  wire g659_n_spl_0;
  wire g659_n_spl_00;
  wire g659_n_spl_01;
  wire g659_n_spl_1;
  wire g659_n_spl_10;
  wire g705_p_spl_;
  wire g676_n_spl_;
  wire g707_n_spl_;
  wire g711_p_spl_;
  wire g684_n_spl_;
  wire g713_n_spl_;
  wire ffc_126_p_spl_;
  wire ffc_129_p_spl_;
  wire ffc_162_p_spl_;
  wire ffc_132_p_spl_;
  wire ffc_132_n_spl_;
  wire g581_n_spl_;
  wire g581_n_spl_0;
  wire g581_n_spl_00;
  wire g581_n_spl_01;
  wire g581_n_spl_1;
  wire ffc_145_p_spl_;
  wire ffc_15_p_spl_;
  wire ffc_15_p_spl_0;
  wire g583_n_spl_;
  wire g583_n_spl_0;
  wire g583_n_spl_00;
  wire g583_n_spl_01;
  wire g583_n_spl_1;
  wire g890_n_spl_;
  wire g1013_p_spl_;
  wire g1013_p_spl_0;
  wire g886_n_spl_;
  wire g886_n_spl_0;
  wire ffc_13_p_spl_;
  wire ffc_48_n_spl_;
  wire g976_n_spl_;
  wire ffc_39_p_spl_;
  wire ffc_37_p_spl_;
  wire g1020_n_spl_;
  wire ffc_48_p_spl_;
  wire g590_p_spl_;
  wire g577_p_spl_;
  wire g577_p_spl_0;
  wire g1026_p_spl_;
  wire g656_p_spl_;
  wire g656_p_spl_0;
  wire g1025_n_spl_;
  wire g1025_n_spl_0;
  wire g1031_n_spl_;
  wire G1_p_spl_;
  wire G1_p_spl_0;
  wire G2_n_spl_;
  wire G6_p_spl_;
  wire g662_n_spl_;
  wire g664_n_spl_;
  wire g716_p_spl_;
  wire ffc_196_p_spl_;
  wire ffc_196_p_spl_0;
  wire g591_n_spl_;
  wire ffc_21_p_spl_;
  wire ffc_21_p_spl_0;
  wire g598_n_spl_;
  wire g598_n_spl_0;
  wire g598_n_spl_1;
  wire ffc_137_p_spl_;
  wire g719_n_spl_;
  wire ffc_135_p_spl_;
  wire ffc_135_p_spl_0;
  wire g720_n_spl_;
  wire g950_n_spl_;
  wire g595_n_spl_;
  wire g595_n_spl_0;
  wire g875_n_spl_;
  wire g972_n_spl_;
  wire g876_n_spl_;
  wire ffc_313_p_spl_;
  wire ffc_313_p_spl_0;
  wire g1082_p_spl_;
  wire g1082_p_spl_0;
  wire g1082_p_spl_1;
  wire g666_p_spl_;
  wire g1086_n_spl_;
  wire g1088_p_spl_;
  wire g665_n_spl_;
  wire ffc_352_p_spl_;
  wire ffc_302_p_spl_;
  wire ffc_304_n_spl_;
  wire ffc_304_n_spl_0;
  wire ffc_304_p_spl_;
  wire ffc_304_p_spl_0;
  wire g1108_n_spl_;
  wire g663_p_spl_;
  wire g660_p_spl_;
  wire g990_p_spl_;
  wire g701_n_spl_;
  wire g992_n_spl_;
  wire g995_p_spl_;
  wire g998_p_spl_;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_00;
  wire G4_p_spl_000;
  wire G4_p_spl_001;
  wire G4_p_spl_01;
  wire G4_p_spl_1;
  wire G4_p_spl_10;
  wire G4_p_spl_11;
  wire G11_p_spl_;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire G12_p_spl_1;
  wire G13_p_spl_;
  wire G13_p_spl_0;
  wire ffc_22_p_spl_;
  wire g667_n_spl_;
  wire ffc_23_p_spl_;
  wire g686_p_spl_;
  wire ffc_351_p_spl_;
  wire ffc_351_p_spl_0;
  wire ffc_243_p_spl_;
  wire ffc_243_p_spl_0;
  wire ffc_243_p_spl_00;
  wire ffc_243_p_spl_1;
  wire ffc_27_p_spl_;
  wire ffc_243_n_spl_;
  wire ffc_243_n_spl_0;
  wire ffc_243_n_spl_1;
  wire g1108_p_spl_;
  wire ffc_359_p_spl_;
  wire g691_p_spl_;
  wire G3_p_spl_;
  wire G3_p_spl_0;
  wire G3_p_spl_00;
  wire G3_p_spl_1;
  wire G4_n_spl_;
  wire G4_n_spl_0;
  wire G4_n_spl_00;
  wire G4_n_spl_1;
  wire G3_n_spl_;
  wire g1034_n_spl_;
  wire G5_p_spl_;
  wire G5_p_spl_0;
  wire ffc_325_n_spl_;
  wire ffc_359_n_spl_;
  wire g691_n_spl_;
  wire g658_n_spl_;
  wire g658_n_spl_0;
  wire g1179_p_spl_;
  wire g1085_n_spl_;
  wire g1085_n_spl_0;
  wire g1190_p_spl_;
  wire g1098_n_spl_;
  wire g1098_n_spl_0;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire g1197_n_spl_;
  wire g1035_n_spl_;
  wire g1035_n_spl_0;
  wire g1074_n_spl_;
  wire g985_n_spl_;
  wire g1110_n_spl_;
  wire g1120_p_spl_;
  wire g1121_p_spl_;
  wire G13_n_spl_;
  wire g1124_n_spl_;
  wire g1123_n_spl_;
  wire g1208_p_spl_;
  wire G41_p_spl_;
  wire g1162_n_spl_;
  wire g1162_n_spl_0;
  wire g1162_n_spl_1;
  wire G34_n_spl_;
  wire g1122_n_spl_;
  wire g1122_n_spl_0;
  wire g1122_n_spl_1;
  wire g1164_p_spl_;
  wire G35_p_spl_;
  wire G35_p_spl_0;
  wire g1201_n_spl_;
  wire g1163_n_spl_;
  wire g1200_p_spl_;
  wire G40_p_spl_;
  wire G33_p_spl_;
  wire G14_p_spl_;
  wire G34_p_spl_;
  wire g1210_n_spl_;

  LA
  g_g412_p
  (
    .dout(g412_p),
    .din1(ffc_5_n_spl_),
    .din2(ffc_59_n)
  );


  LA
  g_g413_p
  (
    .dout(g413_p),
    .din1(ffc_0_n_spl_),
    .din2(ffc_1_n_spl_)
  );


  FA
  g_g414_n
  (
    .dout(g414_n),
    .din1(ffc_6_p_spl_),
    .din2(ffc_32_n_spl_0)
  );


  FA
  g_g415_n
  (
    .dout(g415_n),
    .din1(ffc_4_p),
    .din2(ffc_30_n_spl_0)
  );


  LA
  g_g416_p
  (
    .dout(g416_p),
    .din1(g414_n),
    .din2(g415_n)
  );


  FA
  g_g417_n
  (
    .dout(g417_n),
    .din1(ffc_2_p_spl_),
    .din2(ffc_28_n_spl_0)
  );


  FA
  g_g418_n
  (
    .dout(g418_n),
    .din1(ffc_5_p),
    .din2(ffc_31_n_spl_0)
  );


  LA
  g_g419_p
  (
    .dout(g419_p),
    .din1(g417_n),
    .din2(g418_n)
  );


  LA
  g_g420_p
  (
    .dout(g420_p),
    .din1(g416_p),
    .din2(g419_p)
  );


  FA
  g_g421_n
  (
    .dout(g421_n),
    .din1(ffc_9_p_spl_0),
    .din2(ffc_35_n_spl_0)
  );


  FA
  g_g422_n
  (
    .dout(g422_n),
    .din1(ffc_3_p),
    .din2(ffc_29_n_spl_0)
  );


  LA
  g_g423_p
  (
    .dout(g423_p),
    .din1(g421_n),
    .din2(g422_n)
  );


  FA
  g_g424_n
  (
    .dout(g424_n),
    .din1(ffc_7_p_spl_),
    .din2(ffc_33_n_spl_0)
  );


  FA
  g_g425_n
  (
    .dout(g425_n),
    .din1(ffc_8_p_spl_0),
    .din2(ffc_34_n_spl_0)
  );


  LA
  g_g426_p
  (
    .dout(g426_p),
    .din1(g424_n),
    .din2(g425_n)
  );


  LA
  g_g427_p
  (
    .dout(g427_p),
    .din1(g423_p),
    .din2(g426_p)
  );


  LA
  g_g428_p
  (
    .dout(g428_p),
    .din1(g420_p),
    .din2(g427_p)
  );


  FA
  g_g429_n
  (
    .dout(g429_n),
    .din1(g413_p),
    .din2(g428_p)
  );


  LA
  g_g430_p
  (
    .dout(g430_p),
    .din1(ffc_1_n_spl_),
    .din2(ffc_56_p)
  );


  FA
  g_g430_n
  (
    .dout(g430_n),
    .din1(ffc_1_p),
    .din2(ffc_56_n)
  );


  FA
  g_g431_n
  (
    .dout(g431_n),
    .din1(ffc_96_n),
    .din2(g430_n_spl_)
  );


  LA
  g_g432_p
  (
    .dout(g432_p),
    .din1(ffc_33_n_spl_0),
    .din2(ffc_34_n_spl_0)
  );


  FA
  g_g433_n
  (
    .dout(g433_n),
    .din1(ffc_32_n_spl_0),
    .din2(g432_p)
  );


  FA
  g_g434_n
  (
    .dout(g434_n),
    .din1(ffc_62_p),
    .din2(g433_n)
  );


  LA
  g_g435_p
  (
    .dout(g435_p),
    .din1(g431_n),
    .din2(g434_n)
  );


  LA
  g_g436_p
  (
    .dout(g436_p),
    .din1(g429_n),
    .din2(g435_p)
  );


  LA
  g_g437_p
  (
    .dout(g437_p),
    .din1(ffc_34_p_spl_),
    .din2(ffc_35_n_spl_0)
  );


  FA
  g_g437_n
  (
    .dout(g437_n),
    .din1(ffc_34_n_spl_1),
    .din2(ffc_35_p_spl_)
  );


  LA
  g_g438_p
  (
    .dout(g438_p),
    .din1(ffc_34_n_spl_1),
    .din2(ffc_35_p_spl_)
  );


  FA
  g_g438_n
  (
    .dout(g438_n),
    .din1(ffc_34_p_spl_),
    .din2(ffc_35_n_spl_)
  );


  LA
  g_g439_p
  (
    .dout(g439_p),
    .din1(g437_n),
    .din2(g438_n)
  );


  FA
  g_g439_n
  (
    .dout(g439_n),
    .din1(g437_p),
    .din2(g438_p)
  );


  LA
  g_g440_p
  (
    .dout(g440_p),
    .din1(ffc_32_p_spl_),
    .din2(ffc_33_n_spl_1)
  );


  FA
  g_g440_n
  (
    .dout(g440_n),
    .din1(ffc_32_n_spl_1),
    .din2(ffc_33_p_spl_)
  );


  LA
  g_g441_p
  (
    .dout(g441_p),
    .din1(ffc_32_n_spl_1),
    .din2(ffc_33_p_spl_)
  );


  FA
  g_g441_n
  (
    .dout(g441_n),
    .din1(ffc_32_p_spl_),
    .din2(ffc_33_n_spl_1)
  );


  LA
  g_g442_p
  (
    .dout(g442_p),
    .din1(g440_n),
    .din2(g441_n)
  );


  FA
  g_g442_n
  (
    .dout(g442_n),
    .din1(g440_p),
    .din2(g441_p)
  );


  LA
  g_g443_p
  (
    .dout(g443_p),
    .din1(g439_n_spl_),
    .din2(g442_p_spl_)
  );


  FA
  g_g443_n
  (
    .dout(g443_n),
    .din1(g439_p_spl_),
    .din2(g442_n_spl_)
  );


  LA
  g_g444_p
  (
    .dout(g444_p),
    .din1(g439_p_spl_),
    .din2(g442_n_spl_)
  );


  FA
  g_g444_n
  (
    .dout(g444_n),
    .din1(g439_n_spl_),
    .din2(g442_p_spl_)
  );


  LA
  g_g445_p
  (
    .dout(g445_p),
    .din1(g443_n),
    .din2(g444_n)
  );


  FA
  g_g445_n
  (
    .dout(g445_n),
    .din1(g443_p),
    .din2(g444_p)
  );


  LA
  g_g446_p
  (
    .dout(g446_p),
    .din1(ffc_30_p_spl_),
    .din2(ffc_31_n_spl_0)
  );


  FA
  g_g446_n
  (
    .dout(g446_n),
    .din1(ffc_30_n_spl_0),
    .din2(ffc_31_p_spl_)
  );


  LA
  g_g447_p
  (
    .dout(g447_p),
    .din1(ffc_30_n_spl_),
    .din2(ffc_31_p_spl_)
  );


  FA
  g_g447_n
  (
    .dout(g447_n),
    .din1(ffc_30_p_spl_),
    .din2(ffc_31_n_spl_)
  );


  LA
  g_g448_p
  (
    .dout(g448_p),
    .din1(g446_n),
    .din2(g447_n)
  );


  FA
  g_g448_n
  (
    .dout(g448_n),
    .din1(g446_p),
    .din2(g447_p)
  );


  LA
  g_g449_p
  (
    .dout(g449_p),
    .din1(ffc_28_p_spl_),
    .din2(ffc_29_n_spl_0)
  );


  FA
  g_g449_n
  (
    .dout(g449_n),
    .din1(ffc_28_n_spl_0),
    .din2(ffc_29_p_spl_)
  );


  LA
  g_g450_p
  (
    .dout(g450_p),
    .din1(ffc_28_n_spl_),
    .din2(ffc_29_p_spl_)
  );


  FA
  g_g450_n
  (
    .dout(g450_n),
    .din1(ffc_28_p_spl_),
    .din2(ffc_29_n_spl_)
  );


  LA
  g_g451_p
  (
    .dout(g451_p),
    .din1(g449_n),
    .din2(g450_n)
  );


  FA
  g_g451_n
  (
    .dout(g451_n),
    .din1(g449_p),
    .din2(g450_p)
  );


  LA
  g_g452_p
  (
    .dout(g452_p),
    .din1(g448_p_spl_),
    .din2(g451_n_spl_)
  );


  FA
  g_g452_n
  (
    .dout(g452_n),
    .din1(g448_n_spl_),
    .din2(g451_p_spl_)
  );


  LA
  g_g453_p
  (
    .dout(g453_p),
    .din1(g448_n_spl_),
    .din2(g451_p_spl_)
  );


  FA
  g_g453_n
  (
    .dout(g453_n),
    .din1(g448_p_spl_),
    .din2(g451_n_spl_)
  );


  LA
  g_g454_p
  (
    .dout(g454_p),
    .din1(g452_n),
    .din2(g453_n)
  );


  FA
  g_g454_n
  (
    .dout(g454_n),
    .din1(g452_p),
    .din2(g453_p)
  );


  FA
  g_g455_n
  (
    .dout(g455_n),
    .din1(g445_p),
    .din2(g454_p)
  );


  FA
  g_g456_n
  (
    .dout(g456_n),
    .din1(g445_n),
    .din2(g454_n)
  );


  LA
  g_g457_p
  (
    .dout(g457_p),
    .din1(g455_n),
    .din2(g456_n)
  );


  LA
  g_g458_p
  (
    .dout(g458_p),
    .din1(ffc_6_p_spl_),
    .din2(ffc_7_p_spl_)
  );


  FA
  g_g458_n
  (
    .dout(g458_n),
    .din1(ffc_6_n),
    .din2(ffc_7_n)
  );


  LA
  g_g459_p
  (
    .dout(g459_p),
    .din1(ffc_57_p),
    .din2(g458_n)
  );


  FA
  g_g459_n
  (
    .dout(g459_n),
    .din1(ffc_57_n),
    .din2(g458_p)
  );


  LA
  g_g460_p
  (
    .dout(g460_p),
    .din1(ffc_8_p_spl_0),
    .din2(ffc_9_n_spl_0)
  );


  FA
  g_g460_n
  (
    .dout(g460_n),
    .din1(ffc_8_n_spl_),
    .din2(ffc_9_p_spl_0)
  );


  LA
  g_g461_p
  (
    .dout(g461_p),
    .din1(ffc_8_n_spl_),
    .din2(ffc_9_p_spl_)
  );


  FA
  g_g461_n
  (
    .dout(g461_n),
    .din1(ffc_8_p_spl_),
    .din2(ffc_9_n_spl_0)
  );


  LA
  g_g462_p
  (
    .dout(g462_p),
    .din1(g460_n),
    .din2(g461_n)
  );


  FA
  g_g462_n
  (
    .dout(g462_n),
    .din1(g460_p),
    .din2(g461_p)
  );


  LA
  g_g463_p
  (
    .dout(g463_p),
    .din1(g459_p_spl_),
    .din2(g462_p_spl_)
  );


  FA
  g_g463_n
  (
    .dout(g463_n),
    .din1(g459_n_spl_),
    .din2(g462_n_spl_)
  );


  LA
  g_g464_p
  (
    .dout(g464_p),
    .din1(g459_n_spl_),
    .din2(g462_n_spl_)
  );


  FA
  g_g464_n
  (
    .dout(g464_n),
    .din1(g459_p_spl_),
    .din2(g462_p_spl_)
  );


  LA
  g_g465_p
  (
    .dout(g465_p),
    .din1(g463_n),
    .din2(g464_n)
  );


  FA
  g_g465_n
  (
    .dout(g465_n),
    .din1(g463_p),
    .din2(g464_p)
  );


  LA
  g_g466_p
  (
    .dout(g466_p),
    .din1(ffc_108_n),
    .din2(g465_n)
  );


  LA
  g_g467_p
  (
    .dout(g467_p),
    .din1(ffc_108_p),
    .din2(g465_p)
  );


  FA
  g_g468_n
  (
    .dout(g468_n),
    .din1(g466_p),
    .din2(g467_p)
  );


  LA
  g_g469_p
  (
    .dout(g469_p),
    .din1(ffc_63_p),
    .din2(ffc_79_p_spl_)
  );


  LA
  g_g470_p
  (
    .dout(g470_p),
    .din1(ffc_64_p),
    .din2(ffc_79_p_spl_)
  );


  FA
  g_g471_n
  (
    .dout(g471_n),
    .din1(ffc_91_p),
    .din2(g470_p)
  );


  LA
  g_g472_p
  (
    .dout(g472_p),
    .din1(ffc_96_p),
    .din2(ffc_106_n_spl_0)
  );


  LA
  g_g473_p
  (
    .dout(g473_p),
    .din1(ffc_0_n_spl_),
    .din2(ffc_66_p)
  );


  FA
  g_g474_n
  (
    .dout(g474_n),
    .din1(g472_p),
    .din2(g473_p)
  );


  LA
  g_g475_p
  (
    .dout(g475_p),
    .din1(ffc_115_n_spl_),
    .din2(ffc_215_n)
  );


  FA
  g_g475_n
  (
    .dout(g475_n),
    .din1(ffc_115_p_spl_),
    .din2(ffc_215_p)
  );


  LA
  g_g476_p
  (
    .dout(g476_p),
    .din1(ffc_208_n),
    .din2(ffc_216_p)
  );


  FA
  g_g476_n
  (
    .dout(g476_n),
    .din1(ffc_208_p),
    .din2(ffc_216_n)
  );


  LA
  g_g477_p
  (
    .dout(g477_p),
    .din1(g475_n),
    .din2(g476_n)
  );


  FA
  g_g477_n
  (
    .dout(g477_n),
    .din1(g475_p),
    .din2(g476_p)
  );


  LA
  g_g478_p
  (
    .dout(g478_p),
    .din1(ffc_206_n),
    .din2(ffc_217_p)
  );


  FA
  g_g478_n
  (
    .dout(g478_n),
    .din1(ffc_206_p),
    .din2(ffc_217_n)
  );


  LA
  g_g479_p
  (
    .dout(g479_p),
    .din1(ffc_115_n_spl_),
    .din2(ffc_231_p)
  );


  FA
  g_g479_n
  (
    .dout(g479_n),
    .din1(ffc_115_p_spl_),
    .din2(ffc_231_n)
  );


  LA
  g_g480_p
  (
    .dout(g480_p),
    .din1(g478_n),
    .din2(g479_n)
  );


  FA
  g_g480_n
  (
    .dout(g480_n),
    .din1(g478_p),
    .din2(g479_p)
  );


  LA
  g_g481_p
  (
    .dout(g481_p),
    .din1(ffc_65_p),
    .din2(ffc_80_p)
  );


  FA
  g_g481_n
  (
    .dout(g481_n),
    .din1(ffc_65_n),
    .din2(ffc_80_n)
  );


  LA
  g_g482_p
  (
    .dout(g482_p),
    .din1(ffc_90_p_spl_),
    .din2(g481_n_spl_)
  );


  FA
  g_g482_n
  (
    .dout(g482_n),
    .din1(ffc_90_n_spl_),
    .din2(g481_p_spl_)
  );


  LA
  g_g483_p
  (
    .dout(g483_p),
    .din1(ffc_90_n_spl_),
    .din2(g481_p_spl_)
  );


  FA
  g_g483_n
  (
    .dout(g483_n),
    .din1(ffc_90_p_spl_),
    .din2(g481_n_spl_)
  );


  LA
  g_g484_p
  (
    .dout(g484_p),
    .din1(g482_n),
    .din2(g483_n)
  );


  FA
  g_g484_n
  (
    .dout(g484_n),
    .din1(g482_p),
    .din2(g483_p)
  );


  LA
  g_g485_p
  (
    .dout(g485_p),
    .din1(ffc_49_p),
    .din2(g484_n)
  );


  FA
  g_g485_n
  (
    .dout(g485_n),
    .din1(ffc_49_n),
    .din2(g484_p)
  );


  LA
  g_g486_p
  (
    .dout(g486_p),
    .din1(ffc_101_p_spl_),
    .din2(ffc_102_p_spl_)
  );


  FA
  g_g486_n
  (
    .dout(g486_n),
    .din1(ffc_101_n_spl_),
    .din2(ffc_102_n_spl_)
  );


  LA
  g_g487_p
  (
    .dout(g487_p),
    .din1(ffc_101_n_spl_),
    .din2(ffc_102_n_spl_)
  );


  FA
  g_g487_n
  (
    .dout(g487_n),
    .din1(ffc_101_p_spl_),
    .din2(ffc_102_p_spl_)
  );


  LA
  g_g488_p
  (
    .dout(g488_p),
    .din1(g486_n),
    .din2(g487_n)
  );


  FA
  g_g488_n
  (
    .dout(g488_n),
    .din1(g486_p),
    .din2(g487_p)
  );


  LA
  g_g489_p
  (
    .dout(g489_p),
    .din1(g485_p),
    .din2(g488_p)
  );


  LA
  g_g490_p
  (
    .dout(g490_p),
    .din1(g485_n),
    .din2(g488_n)
  );


  FA
  g_g491_n
  (
    .dout(g491_n),
    .din1(g489_p),
    .din2(g490_p)
  );


  LA
  g_g492_p
  (
    .dout(g492_p),
    .din1(ffc_61_p),
    .din2(g430_n_spl_)
  );


  LA
  g_g493_p
  (
    .dout(g493_p),
    .din1(g491_n),
    .din2(g492_p)
  );


  LA
  g_g494_p
  (
    .dout(g494_p),
    .din1(ffc_9_n_spl_),
    .din2(g430_p)
  );


  LA
  g_g495_p
  (
    .dout(g495_p),
    .din1(ffc_58_n),
    .din2(g494_p)
  );


  LA
  g_g496_p
  (
    .dout(g496_p),
    .din1(ffc_5_n_spl_),
    .din2(ffc_60_n)
  );


  FA
  g_g497_n
  (
    .dout(g497_n),
    .din1(ffc_2_p_spl_),
    .din2(g496_p)
  );


  FA
  g_g498_n
  (
    .dout(g498_n),
    .din1(ffc_2_n),
    .din2(ffc_4_n)
  );


  LA
  g_g499_p
  (
    .dout(g499_p),
    .din1(ffc_61_n),
    .din2(g498_n)
  );


  LA
  g_g500_p
  (
    .dout(g500_p),
    .din1(g497_n),
    .din2(g499_p)
  );


  FA
  g_g501_n
  (
    .dout(g501_n),
    .din1(g495_p),
    .din2(g500_p)
  );


  FA
  g_g502_n
  (
    .dout(g502_n),
    .din1(g493_p),
    .din2(g501_n)
  );


  LA
  g_g503_p
  (
    .dout(g503_p),
    .din1(ffc_218_p),
    .din2(ffc_220_n)
  );


  FA
  g_g503_n
  (
    .dout(g503_n),
    .din1(ffc_218_n),
    .din2(ffc_220_p)
  );


  LA
  g_g504_p
  (
    .dout(g504_p),
    .din1(ffc_212_n),
    .din2(ffc_232_p)
  );


  FA
  g_g504_n
  (
    .dout(g504_n),
    .din1(ffc_212_p),
    .din2(ffc_232_n)
  );


  LA
  g_g505_p
  (
    .dout(g505_p),
    .din1(g503_n),
    .din2(g504_n)
  );


  FA
  g_g505_n
  (
    .dout(g505_n),
    .din1(g503_p),
    .din2(g504_p)
  );


  LA
  g_g506_p
  (
    .dout(g506_p),
    .din1(ffc_106_n_spl_0),
    .din2(ffc_224_p)
  );


  FA
  g_g506_n
  (
    .dout(g506_n),
    .din1(ffc_106_p_spl_),
    .din2(ffc_224_n)
  );


  LA
  g_g507_p
  (
    .dout(g507_p),
    .din1(ffc_213_n),
    .din2(ffc_226_n)
  );


  FA
  g_g507_n
  (
    .dout(g507_n),
    .din1(ffc_213_p),
    .din2(ffc_226_p)
  );


  LA
  g_g508_p
  (
    .dout(g508_p),
    .din1(g506_n),
    .din2(g507_p)
  );


  FA
  g_g508_n
  (
    .dout(g508_n),
    .din1(g506_p),
    .din2(g507_n)
  );


  LA
  g_g509_p
  (
    .dout(g509_p),
    .din1(ffc_106_n_spl_),
    .din2(ffc_229_p)
  );


  FA
  g_g509_n
  (
    .dout(g509_n),
    .din1(ffc_106_p_spl_),
    .din2(ffc_229_n)
  );


  LA
  g_g510_p
  (
    .dout(g510_p),
    .din1(ffc_214_n),
    .din2(ffc_228_n)
  );


  FA
  g_g510_n
  (
    .dout(g510_n),
    .din1(ffc_214_p),
    .din2(ffc_228_p)
  );


  LA
  g_g511_p
  (
    .dout(g511_p),
    .din1(g509_n),
    .din2(g510_p)
  );


  FA
  g_g511_n
  (
    .dout(g511_n),
    .din1(g509_p),
    .din2(g510_n)
  );


  LA
  g_g512_p
  (
    .dout(g512_p),
    .din1(ffc_205_n),
    .din2(ffc_219_p)
  );


  FA
  g_g512_n
  (
    .dout(g512_n),
    .din1(ffc_205_p),
    .din2(ffc_219_n)
  );


  LA
  g_g513_p
  (
    .dout(g513_p),
    .din1(ffc_211_n),
    .din2(ffc_227_p)
  );


  FA
  g_g513_n
  (
    .dout(g513_n),
    .din1(ffc_211_p),
    .din2(ffc_227_n)
  );


  LA
  g_g514_p
  (
    .dout(g514_p),
    .din1(g512_n),
    .din2(g513_n)
  );


  FA
  g_g514_n
  (
    .dout(g514_n),
    .din1(g512_p),
    .din2(g513_p)
  );


  LA
  g_g515_p
  (
    .dout(g515_p),
    .din1(g480_p_spl_),
    .din2(g514_p_spl_)
  );


  FA
  g_g515_n
  (
    .dout(g515_n),
    .din1(g480_n_spl_0),
    .din2(g514_n_spl_0)
  );


  LA
  g_g516_p
  (
    .dout(g516_p),
    .din1(g505_p_spl_),
    .din2(g511_p_spl_)
  );


  FA
  g_g516_n
  (
    .dout(g516_n),
    .din1(g505_n_spl_0),
    .din2(g511_n_spl_0)
  );


  LA
  g_g517_p
  (
    .dout(g517_p),
    .din1(g477_p_spl_),
    .din2(g508_p_spl_)
  );


  FA
  g_g517_n
  (
    .dout(g517_n),
    .din1(g477_n_spl_0),
    .din2(g508_n_spl_0)
  );


  FA
  g_g518_n
  (
    .dout(g518_n),
    .din1(g516_n_spl_),
    .din2(g517_n_spl_)
  );


  FA
  g_g519_n
  (
    .dout(g519_n),
    .din1(g515_n_spl_),
    .din2(g518_n)
  );


  FA
  g_g520_n
  (
    .dout(g520_n),
    .din1(ffc_233_p_spl_0),
    .din2(g519_n)
  );


  LA
  g_g521_p
  (
    .dout(g521_p),
    .din1(ffc_25_p_spl_),
    .din2(ffc_51_p)
  );


  FA
  g_g521_n
  (
    .dout(g521_n),
    .din1(ffc_25_n),
    .din2(ffc_51_n)
  );


  FA
  g_g522_n
  (
    .dout(g522_n),
    .din1(ffc_233_p_spl_0),
    .din2(g521_n_spl_)
  );


  LA
  g_g523_p
  (
    .dout(g523_p),
    .din1(ffc_25_p_spl_),
    .din2(g522_n)
  );


  LA
  g_g524_p
  (
    .dout(g524_p),
    .din1(g520_n_spl_),
    .din2(g523_p)
  );


  LA
  g_g525_p
  (
    .dout(g525_p),
    .din1(g477_n_spl_0),
    .din2(g508_n_spl_0)
  );


  FA
  g_g525_n
  (
    .dout(g525_n),
    .din1(g477_p_spl_),
    .din2(g508_p_spl_)
  );


  LA
  g_g526_p
  (
    .dout(g526_p),
    .din1(g517_n_spl_),
    .din2(g525_n)
  );


  FA
  g_g526_n
  (
    .dout(g526_n),
    .din1(g517_p),
    .din2(g525_p)
  );


  LA
  g_g527_p
  (
    .dout(g527_p),
    .din1(g505_n_spl_0),
    .din2(g511_n_spl_0)
  );


  FA
  g_g527_n
  (
    .dout(g527_n),
    .din1(g505_p_spl_),
    .din2(g511_p_spl_)
  );


  LA
  g_g528_p
  (
    .dout(g528_p),
    .din1(g516_n_spl_),
    .din2(g527_n)
  );


  FA
  g_g528_n
  (
    .dout(g528_n),
    .din1(g516_p),
    .din2(g527_p)
  );


  LA
  g_g529_p
  (
    .dout(g529_p),
    .din1(g526_p_spl_),
    .din2(g528_n_spl_)
  );


  FA
  g_g529_n
  (
    .dout(g529_n),
    .din1(g526_n_spl_),
    .din2(g528_p_spl_)
  );


  LA
  g_g530_p
  (
    .dout(g530_p),
    .din1(g526_n_spl_),
    .din2(g528_p_spl_)
  );


  FA
  g_g530_n
  (
    .dout(g530_n),
    .din1(g526_p_spl_),
    .din2(g528_n_spl_)
  );


  LA
  g_g531_p
  (
    .dout(g531_p),
    .din1(g529_n),
    .din2(g530_n)
  );


  FA
  g_g531_n
  (
    .dout(g531_n),
    .din1(g529_p),
    .din2(g530_p)
  );


  LA
  g_g532_p
  (
    .dout(g532_p),
    .din1(g480_n_spl_0),
    .din2(g514_n_spl_0)
  );


  FA
  g_g532_n
  (
    .dout(g532_n),
    .din1(g480_p_spl_),
    .din2(g514_p_spl_)
  );


  LA
  g_g533_p
  (
    .dout(g533_p),
    .din1(g515_n_spl_),
    .din2(g532_n)
  );


  FA
  g_g533_n
  (
    .dout(g533_n),
    .din1(g515_p),
    .din2(g532_p)
  );


  LA
  g_g534_p
  (
    .dout(g534_p),
    .din1(ffc_233_p_spl_),
    .din2(ffc_234_n)
  );


  FA
  g_g534_n
  (
    .dout(g534_n),
    .din1(ffc_233_n),
    .din2(ffc_234_p)
  );


  LA
  g_g535_p
  (
    .dout(g535_p),
    .din1(ffc_55_p_spl_),
    .din2(g534_n_spl_0)
  );


  FA
  g_g535_n
  (
    .dout(g535_n),
    .din1(ffc_55_n_spl_),
    .din2(g534_p_spl_0)
  );


  LA
  g_g536_p
  (
    .dout(g536_p),
    .din1(ffc_55_n_spl_),
    .din2(g534_p_spl_0)
  );


  FA
  g_g536_n
  (
    .dout(g536_n),
    .din1(ffc_55_p_spl_),
    .din2(g534_n_spl_0)
  );


  LA
  g_g537_p
  (
    .dout(g537_p),
    .din1(g535_n),
    .din2(g536_n)
  );


  FA
  g_g537_n
  (
    .dout(g537_n),
    .din1(g535_p),
    .din2(g536_p)
  );


  LA
  g_g538_p
  (
    .dout(g538_p),
    .din1(g521_n_spl_),
    .din2(g537_n)
  );


  FA
  g_g538_n
  (
    .dout(g538_n),
    .din1(g521_p),
    .din2(g537_p)
  );


  LA
  g_g539_p
  (
    .dout(g539_p),
    .din1(g533_p_spl_0),
    .din2(g538_p_spl_)
  );


  FA
  g_g539_n
  (
    .dout(g539_n),
    .din1(g533_n_spl_0),
    .din2(g538_n_spl_)
  );


  LA
  g_g540_p
  (
    .dout(g540_p),
    .din1(g533_n_spl_0),
    .din2(g538_n_spl_)
  );


  FA
  g_g540_n
  (
    .dout(g540_n),
    .din1(g533_p_spl_0),
    .din2(g538_p_spl_)
  );


  LA
  g_g541_p
  (
    .dout(g541_p),
    .din1(g539_n),
    .din2(g540_n)
  );


  FA
  g_g541_n
  (
    .dout(g541_n),
    .din1(g539_p),
    .din2(g540_p)
  );


  LA
  g_g542_p
  (
    .dout(g542_p),
    .din1(g531_n_spl_),
    .din2(g541_n)
  );


  LA
  g_g543_p
  (
    .dout(g543_p),
    .din1(g531_p_spl_),
    .din2(g541_p)
  );


  FA
  g_g544_n
  (
    .dout(g544_n),
    .din1(g542_p),
    .din2(g543_p)
  );


  LA
  g_g545_p
  (
    .dout(g545_p),
    .din1(g533_n_spl_1),
    .din2(g534_n_spl_1)
  );


  FA
  g_g545_n
  (
    .dout(g545_n),
    .din1(g533_p_spl_1),
    .din2(g534_p_spl_1)
  );


  LA
  g_g546_p
  (
    .dout(g546_p),
    .din1(g533_p_spl_1),
    .din2(g534_p_spl_1)
  );


  FA
  g_g546_n
  (
    .dout(g546_n),
    .din1(g533_n_spl_1),
    .din2(g534_n_spl_1)
  );


  LA
  g_g547_p
  (
    .dout(g547_p),
    .din1(g545_n),
    .din2(g546_n)
  );


  FA
  g_g547_n
  (
    .dout(g547_n),
    .din1(g545_p),
    .din2(g546_p)
  );


  FA
  g_g548_n
  (
    .dout(g548_n),
    .din1(g531_p_spl_),
    .din2(g547_p)
  );


  FA
  g_g549_n
  (
    .dout(g549_n),
    .din1(g531_n_spl_),
    .din2(g547_n)
  );


  LA
  g_g550_p
  (
    .dout(g550_p),
    .din1(g548_n),
    .din2(g549_n)
  );


  FA
  g_g551_n
  (
    .dout(g551_n),
    .din1(ffc_103_p_spl_0),
    .din2(ffc_107_n)
  );


  FA
  g_g552_n
  (
    .dout(g552_n),
    .din1(ffc_72_n_spl_),
    .din2(ffc_86_n)
  );


  LA
  g_g553_p
  (
    .dout(g553_p),
    .din1(ffc_235_n_spl_0),
    .din2(ffc_269_p)
  );


  FA
  g_g553_n
  (
    .dout(g553_n),
    .din1(ffc_235_p_spl_),
    .din2(ffc_269_n)
  );


  LA
  g_g554_p
  (
    .dout(g554_p),
    .din1(ffc_266_n),
    .din2(ffc_288_n)
  );


  FA
  g_g554_n
  (
    .dout(g554_n),
    .din1(ffc_266_p),
    .din2(ffc_288_p)
  );


  LA
  g_g555_p
  (
    .dout(g555_p),
    .din1(ffc_274_p),
    .din2(ffc_290_n)
  );


  FA
  g_g555_n
  (
    .dout(g555_n),
    .din1(ffc_274_n),
    .din2(ffc_290_p_spl_)
  );


  LA
  g_g556_p
  (
    .dout(g556_p),
    .din1(ffc_81_p),
    .din2(ffc_118_n_spl_)
  );


  FA
  g_g556_n
  (
    .dout(g556_n),
    .din1(ffc_81_n),
    .din2(ffc_118_p_spl_0)
  );


  LA
  g_g557_p
  (
    .dout(g557_p),
    .din1(ffc_263_p),
    .din2(ffc_284_n)
  );


  LA
  g_g558_p
  (
    .dout(g558_p),
    .din1(ffc_263_n),
    .din2(ffc_284_p)
  );


  FA
  g_g559_n
  (
    .dout(g559_n),
    .din1(g557_p),
    .din2(g558_p)
  );


  LA
  g_g560_p
  (
    .dout(g560_p),
    .din1(ffc_71_p_spl_),
    .din2(ffc_254_n)
  );


  FA
  g_g560_n
  (
    .dout(g560_n),
    .din1(ffc_71_n_spl_),
    .din2(ffc_254_p_spl_)
  );


  LA
  g_g561_p
  (
    .dout(g561_p),
    .din1(ffc_67_n),
    .din2(g560_n)
  );


  FA
  g_g561_n
  (
    .dout(g561_n),
    .din1(ffc_67_p_spl_),
    .din2(g560_p)
  );


  LA
  g_g562_p
  (
    .dout(g562_p),
    .din1(g556_p_spl_0),
    .din2(g561_p_spl_)
  );


  FA
  g_g562_n
  (
    .dout(g562_n),
    .din1(g556_n_spl_0),
    .din2(g561_n_spl_00)
  );


  LA
  g_g563_p
  (
    .dout(g563_p),
    .din1(ffc_329_p_spl_),
    .din2(ffc_330_p_spl_)
  );


  FA
  g_g563_n
  (
    .dout(g563_n),
    .din1(ffc_329_n_spl_),
    .din2(ffc_330_n_spl_)
  );


  LA
  g_g564_p
  (
    .dout(g564_p),
    .din1(ffc_310_n),
    .din2(ffc_311_n)
  );


  FA
  g_g564_n
  (
    .dout(g564_n),
    .din1(ffc_310_p),
    .din2(ffc_311_p)
  );


  LA
  g_g565_p
  (
    .dout(g565_p),
    .din1(ffc_328_n_spl_000),
    .din2(g564_p)
  );


  FA
  g_g565_n
  (
    .dout(g565_n),
    .din1(ffc_328_p_spl_000),
    .din2(g564_n)
  );


  LA
  g_g566_p
  (
    .dout(g566_p),
    .din1(ffc_328_p_spl_000),
    .din2(g563_p_spl_)
  );


  FA
  g_g566_n
  (
    .dout(g566_n),
    .din1(ffc_328_n_spl_000),
    .din2(g563_n)
  );


  LA
  g_g567_p
  (
    .dout(g567_p),
    .din1(g565_n),
    .din2(g566_n)
  );


  FA
  g_g567_n
  (
    .dout(g567_n),
    .din1(g565_p),
    .din2(g566_p)
  );


  LA
  g_g568_p
  (
    .dout(g568_p),
    .din1(ffc_319_n_spl_0),
    .din2(ffc_321_p)
  );


  FA
  g_g568_n
  (
    .dout(g568_n),
    .din1(ffc_319_p_spl_),
    .din2(ffc_321_n)
  );


  LA
  g_g569_p
  (
    .dout(g569_p),
    .din1(ffc_292_p),
    .din2(ffc_328_p_spl_001)
  );


  FA
  g_g569_n
  (
    .dout(g569_n),
    .din1(ffc_292_n),
    .din2(ffc_328_n_spl_001)
  );


  LA
  g_g570_p
  (
    .dout(g570_p),
    .din1(g568_n_spl_0),
    .din2(g569_n_spl_)
  );


  FA
  g_g570_n
  (
    .dout(g570_n),
    .din1(g568_p_spl_),
    .din2(g569_p_spl_)
  );


  LA
  g_g571_p
  (
    .dout(g571_p),
    .din1(g568_p_spl_),
    .din2(g569_p_spl_)
  );


  FA
  g_g571_n
  (
    .dout(g571_n),
    .din1(g568_n_spl_0),
    .din2(g569_n_spl_)
  );


  LA
  g_g572_p
  (
    .dout(g572_p),
    .din1(g570_n),
    .din2(g571_n)
  );


  FA
  g_g572_n
  (
    .dout(g572_n),
    .din1(g570_p),
    .din2(g571_p)
  );


  LA
  g_g573_p
  (
    .dout(g573_p),
    .din1(ffc_320_n_spl_0),
    .din2(ffc_322_p)
  );


  FA
  g_g573_n
  (
    .dout(g573_n),
    .din1(ffc_320_p_spl_),
    .din2(ffc_322_n)
  );


  LA
  g_g574_p
  (
    .dout(g574_p),
    .din1(ffc_295_p),
    .din2(ffc_328_p_spl_001)
  );


  FA
  g_g574_n
  (
    .dout(g574_n),
    .din1(ffc_295_n),
    .din2(ffc_328_n_spl_001)
  );


  LA
  g_g575_p
  (
    .dout(g575_p),
    .din1(g573_n_spl_0),
    .din2(g574_n_spl_)
  );


  FA
  g_g575_n
  (
    .dout(g575_n),
    .din1(g573_p_spl_),
    .din2(g574_p_spl_)
  );


  LA
  g_g576_p
  (
    .dout(g576_p),
    .din1(g573_p_spl_),
    .din2(g574_p_spl_)
  );


  FA
  g_g576_n
  (
    .dout(g576_n),
    .din1(g573_n_spl_0),
    .din2(g574_n_spl_)
  );


  LA
  g_g577_p
  (
    .dout(g577_p),
    .din1(g575_n),
    .din2(g576_n)
  );


  FA
  g_g577_n
  (
    .dout(g577_n),
    .din1(g575_p),
    .din2(g576_p)
  );


  LA
  g_g578_p
  (
    .dout(g578_p),
    .din1(ffc_124_p_spl_00),
    .din2(ffc_165_p)
  );


  FA
  g_g578_n
  (
    .dout(g578_n),
    .din1(ffc_124_n_spl_0),
    .din2(ffc_165_n)
  );


  LA
  g_g579_p
  (
    .dout(g579_p),
    .din1(ffc_124_p_spl_00),
    .din2(ffc_166_p)
  );


  FA
  g_g579_n
  (
    .dout(g579_n),
    .din1(ffc_124_n_spl_0),
    .din2(ffc_166_n)
  );


  FA
  g_g580_n
  (
    .dout(g580_n),
    .din1(ffc_167_n_spl_),
    .din2(g579_p_spl_00)
  );


  FA
  g_g581_n
  (
    .dout(g581_n),
    .din1(g578_p_spl_0),
    .din2(g580_n)
  );


  FA
  g_g582_n
  (
    .dout(g582_n),
    .din1(ffc_167_p_spl_),
    .din2(g579_p_spl_00)
  );


  FA
  g_g583_n
  (
    .dout(g583_n),
    .din1(g578_p_spl_0),
    .din2(g582_n)
  );


  LA
  g_g584_p
  (
    .dout(g584_p),
    .din1(ffc_297_p),
    .din2(ffc_330_p_spl_)
  );


  FA
  g_g584_n
  (
    .dout(g584_n),
    .din1(ffc_297_n_spl_),
    .din2(ffc_330_n_spl_)
  );


  LA
  g_g585_p
  (
    .dout(g585_p),
    .din1(ffc_239_p_spl_),
    .din2(ffc_300_p)
  );


  FA
  g_g585_n
  (
    .dout(g585_n),
    .din1(ffc_239_n),
    .din2(ffc_300_n)
  );


  LA
  g_g586_p
  (
    .dout(g586_p),
    .din1(ffc_200_p_spl_),
    .din2(ffc_240_p_spl_)
  );


  FA
  g_g586_n
  (
    .dout(g586_n),
    .din1(ffc_200_n),
    .din2(ffc_240_n)
  );


  LA
  g_g587_p
  (
    .dout(g587_p),
    .din1(ffc_199_n),
    .din2(g586_n)
  );


  FA
  g_g587_n
  (
    .dout(g587_n),
    .din1(ffc_199_p),
    .din2(g586_p)
  );


  LA
  g_g588_p
  (
    .dout(g588_p),
    .din1(g585_n),
    .din2(g587_p)
  );


  FA
  g_g588_n
  (
    .dout(g588_n),
    .din1(g585_p),
    .din2(g587_n)
  );


  LA
  g_g589_p
  (
    .dout(g589_p),
    .din1(g584_n),
    .din2(g588_p)
  );


  FA
  g_g589_n
  (
    .dout(g589_n),
    .din1(g584_p),
    .din2(g588_n)
  );


  LA
  g_g590_p
  (
    .dout(g590_p),
    .din1(g567_p_spl_0),
    .din2(g572_p_spl_0)
  );


  FA
  g_g590_n
  (
    .dout(g590_n),
    .din1(g567_n),
    .din2(g572_n)
  );


  FA
  g_g591_n
  (
    .dout(g591_n),
    .din1(ffc_19_p_spl_0),
    .din2(ffc_162_n_spl_)
  );


  LA
  g_g592_p
  (
    .dout(g592_p),
    .din1(ffc_328_n_spl_01),
    .din2(g589_n_spl_)
  );


  FA
  g_g592_n
  (
    .dout(g592_n),
    .din1(ffc_328_p_spl_010),
    .din2(g589_p)
  );


  LA
  g_g593_p
  (
    .dout(g593_p),
    .din1(ffc_124_p_spl_0),
    .din2(ffc_167_p_spl_)
  );


  FA
  g_g593_n
  (
    .dout(g593_n),
    .din1(ffc_124_n_spl_),
    .din2(ffc_167_n_spl_)
  );


  LA
  g_g594_p
  (
    .dout(g594_p),
    .din1(g578_n_spl_),
    .din2(g593_n_spl_)
  );


  FA
  g_g594_n
  (
    .dout(g594_n),
    .din1(g578_p_spl_1),
    .din2(g593_p_spl_)
  );


  LA
  g_g595_p
  (
    .dout(g595_p),
    .din1(g579_n_spl_0),
    .din2(g594_p_spl_)
  );


  FA
  g_g595_n
  (
    .dout(g595_n),
    .din1(g579_p_spl_01),
    .din2(g594_n_spl_)
  );


  LA
  g_g596_p
  (
    .dout(g596_p),
    .din1(g578_n_spl_),
    .din2(g593_p_spl_)
  );


  FA
  g_g596_n
  (
    .dout(g596_n),
    .din1(g578_p_spl_1),
    .din2(g593_n_spl_)
  );


  LA
  g_g597_p
  (
    .dout(g597_p),
    .din1(g579_p_spl_01),
    .din2(g596_p_spl_)
  );


  FA
  g_g597_n
  (
    .dout(g597_n),
    .din1(g579_n_spl_0),
    .din2(g596_n_spl_)
  );


  LA
  g_g598_p
  (
    .dout(g598_p),
    .din1(g579_p_spl_1),
    .din2(g594_p_spl_)
  );


  FA
  g_g598_n
  (
    .dout(g598_n),
    .din1(g579_n_spl_1),
    .din2(g594_n_spl_)
  );


  LA
  g_g599_p
  (
    .dout(g599_p),
    .din1(g579_n_spl_1),
    .din2(g596_p_spl_)
  );


  FA
  g_g599_n
  (
    .dout(g599_n),
    .din1(g579_p_spl_1),
    .din2(g596_n_spl_)
  );


  LA
  g_g600_p
  (
    .dout(g600_p),
    .din1(ffc_275_n_spl_),
    .din2(ffc_276_n)
  );


  FA
  g_g600_n
  (
    .dout(g600_n),
    .din1(ffc_275_p_spl_),
    .din2(ffc_276_p)
  );


  LA
  g_g601_p
  (
    .dout(g601_p),
    .din1(ffc_293_p),
    .din2(ffc_294_n)
  );


  FA
  g_g601_n
  (
    .dout(g601_n),
    .din1(ffc_293_n),
    .din2(ffc_294_p)
  );


  LA
  g_g602_p
  (
    .dout(g602_p),
    .din1(ffc_155_p_spl_0),
    .din2(ffc_267_p_spl_)
  );


  FA
  g_g602_n
  (
    .dout(g602_n),
    .din1(ffc_155_n_spl_0),
    .din2(ffc_267_n)
  );


  LA
  g_g603_p
  (
    .dout(g603_p),
    .din1(g555_n),
    .din2(g602_p)
  );


  FA
  g_g603_n
  (
    .dout(g603_n),
    .din1(g555_p_spl_),
    .din2(g602_n)
  );


  LA
  g_g604_p
  (
    .dout(g604_p),
    .din1(g601_n_spl_0),
    .din2(g603_n_spl_)
  );


  FA
  g_g604_n
  (
    .dout(g604_n),
    .din1(g601_p_spl_),
    .din2(g603_p_spl_)
  );


  LA
  g_g605_p
  (
    .dout(g605_p),
    .din1(g600_p),
    .din2(g604_n_spl_)
  );


  LA
  g_g606_p
  (
    .dout(g606_p),
    .din1(g600_n_spl_0),
    .din2(g604_p)
  );


  FA
  g_g607_n
  (
    .dout(g607_n),
    .din1(g605_p),
    .din2(g606_p)
  );


  LA
  g_g608_p
  (
    .dout(g608_p),
    .din1(g556_n_spl_0),
    .din2(g607_n)
  );


  FA
  g_g609_n
  (
    .dout(g609_n),
    .din1(ffc_69_p),
    .din2(ffc_70_n_spl_00)
  );


  FA
  g_g610_n
  (
    .dout(g610_n),
    .din1(ffc_179_n),
    .din2(g609_n_spl_0)
  );


  LA
  g_g611_p
  (
    .dout(g611_p),
    .din1(ffc_68_p_spl_),
    .din2(ffc_105_n)
  );


  FA
  g_g611_n
  (
    .dout(g611_n),
    .din1(ffc_68_n),
    .din2(ffc_105_p)
  );


  LA
  g_g612_p
  (
    .dout(g612_p),
    .din1(ffc_84_p_spl_),
    .din2(g611_n)
  );


  FA
  g_g612_n
  (
    .dout(g612_n),
    .din1(ffc_84_n),
    .din2(g611_p)
  );


  FA
  g_g613_n
  (
    .dout(g613_n),
    .din1(ffc_281_n),
    .din2(ffc_287_p)
  );


  FA
  g_g614_n
  (
    .dout(g614_n),
    .din1(ffc_280_n),
    .din2(ffc_298_n)
  );


  LA
  g_g615_p
  (
    .dout(g615_p),
    .din1(g613_n),
    .din2(g614_n)
  );


  FA
  g_g616_n
  (
    .dout(g616_n),
    .din1(g612_p_spl_00),
    .din2(g615_p)
  );


  LA
  g_g617_p
  (
    .dout(g617_p),
    .din1(g562_p_spl_00),
    .din2(g616_n)
  );


  LA
  g_g618_p
  (
    .dout(g618_p),
    .din1(g610_n),
    .din2(g617_p)
  );


  LA
  g_g619_p
  (
    .dout(g619_p),
    .din1(g561_n_spl_00),
    .din2(g600_n_spl_0)
  );


  FA
  g_g620_n
  (
    .dout(g620_n),
    .din1(g618_p),
    .din2(g619_p)
  );


  FA
  g_g621_n
  (
    .dout(g621_n),
    .din1(g608_p),
    .din2(g620_n)
  );


  LA
  g_g622_p
  (
    .dout(g622_p),
    .din1(ffc_272_p),
    .din2(ffc_273_n)
  );


  FA
  g_g622_n
  (
    .dout(g622_n),
    .din1(ffc_272_n),
    .din2(ffc_273_p)
  );


  FA
  g_g623_n
  (
    .dout(g623_n),
    .din1(g609_n_spl_0),
    .din2(g622_n_spl_0)
  );


  FA
  g_g624_n
  (
    .dout(g624_n),
    .din1(ffc_268_p),
    .din2(ffc_296_p)
  );


  FA
  g_g625_n
  (
    .dout(g625_n),
    .din1(ffc_259_n),
    .din2(ffc_286_p)
  );


  FA
  g_g626_n
  (
    .dout(g626_n),
    .din1(g624_n),
    .din2(g625_n)
  );


  FA
  g_g627_n
  (
    .dout(g627_n),
    .din1(ffc_257_n),
    .din2(ffc_283_n)
  );


  FA
  g_g628_n
  (
    .dout(g628_n),
    .din1(ffc_282_n),
    .din2(ffc_285_n)
  );


  FA
  g_g629_n
  (
    .dout(g629_n),
    .din1(g627_n),
    .din2(g628_n)
  );


  LA
  g_g630_p
  (
    .dout(g630_p),
    .din1(g626_n),
    .din2(g629_n)
  );


  FA
  g_g631_n
  (
    .dout(g631_n),
    .din1(g612_p_spl_00),
    .din2(g630_p)
  );


  LA
  g_g632_p
  (
    .dout(g632_p),
    .din1(g562_p_spl_00),
    .din2(g631_n)
  );


  LA
  g_g633_p
  (
    .dout(g633_p),
    .din1(g623_n),
    .din2(g632_p)
  );


  LA
  g_g634_p
  (
    .dout(g634_p),
    .din1(g554_n_spl_0),
    .din2(g622_n_spl_0)
  );


  FA
  g_g634_n
  (
    .dout(g634_n),
    .din1(g554_p_spl_),
    .din2(g622_p_spl_)
  );


  LA
  g_g635_p
  (
    .dout(g635_p),
    .din1(g554_p_spl_),
    .din2(g622_p_spl_)
  );


  FA
  g_g635_n
  (
    .dout(g635_n),
    .din1(g554_n_spl_0),
    .din2(g622_n_spl_)
  );


  LA
  g_g636_p
  (
    .dout(g636_p),
    .din1(g634_n),
    .din2(g635_n)
  );


  FA
  g_g636_n
  (
    .dout(g636_n),
    .din1(g634_p),
    .din2(g635_p)
  );


  LA
  g_g637_p
  (
    .dout(g637_p),
    .din1(ffc_275_n_spl_),
    .din2(g636_n)
  );


  LA
  g_g638_p
  (
    .dout(g638_p),
    .din1(ffc_275_p_spl_),
    .din2(g636_p)
  );


  FA
  g_g639_n
  (
    .dout(g639_n),
    .din1(g637_p),
    .din2(g638_p)
  );


  LA
  g_g640_p
  (
    .dout(g640_p),
    .din1(g600_n_spl_),
    .din2(g601_n_spl_0)
  );


  FA
  g_g641_n
  (
    .dout(g641_n),
    .din1(g603_n_spl_),
    .din2(g640_p)
  );


  LA
  g_g642_p
  (
    .dout(g642_p),
    .din1(g556_n_spl_1),
    .din2(g641_n)
  );


  FA
  g_g643_n
  (
    .dout(g643_n),
    .din1(g561_n_spl_01),
    .din2(g642_p)
  );


  LA
  g_g644_p
  (
    .dout(g644_p),
    .din1(g639_n),
    .din2(g643_n)
  );


  FA
  g_g645_n
  (
    .dout(g645_n),
    .din1(g633_p),
    .din2(g644_p)
  );


  FA
  g_g646_n
  (
    .dout(g646_n),
    .din1(ffc_333_p_spl_0),
    .din2(ffc_357_p_spl_00)
  );


  LA
  g_g647_p
  (
    .dout(g647_p),
    .din1(ffc_182_p),
    .din2(ffc_312_n_spl_)
  );


  FA
  g_g647_n
  (
    .dout(g647_n),
    .din1(ffc_182_n_spl_),
    .din2(ffc_312_p_spl_)
  );


  LA
  g_g648_p
  (
    .dout(g648_p),
    .din1(ffc_308_n),
    .din2(ffc_318_n)
  );


  FA
  g_g648_n
  (
    .dout(g648_n),
    .din1(ffc_308_p),
    .din2(ffc_318_p)
  );


  LA
  g_g649_p
  (
    .dout(g649_p),
    .din1(g647_n),
    .din2(g648_p_spl_0)
  );


  FA
  g_g649_n
  (
    .dout(g649_n),
    .din1(g647_p),
    .din2(g648_n_spl_0)
  );


  LA
  g_g650_p
  (
    .dout(g650_p),
    .din1(ffc_181_p_spl_),
    .din2(ffc_312_n_spl_)
  );


  FA
  g_g650_n
  (
    .dout(g650_n),
    .din1(ffc_181_n_spl_),
    .din2(ffc_312_p_spl_)
  );


  LA
  g_g651_p
  (
    .dout(g651_p),
    .din1(g648_n_spl_0),
    .din2(g650_p)
  );


  FA
  g_g651_n
  (
    .dout(g651_n),
    .din1(g648_p_spl_0),
    .din2(g650_n)
  );


  LA
  g_g652_p
  (
    .dout(g652_p),
    .din1(g649_n),
    .din2(g651_n_spl_)
  );


  FA
  g_g652_n
  (
    .dout(g652_n),
    .din1(g649_p),
    .din2(g651_p_spl_)
  );


  LA
  g_g653_p
  (
    .dout(g653_p),
    .din1(ffc_291_p),
    .din2(g648_n_spl_)
  );


  FA
  g_g653_n
  (
    .dout(g653_n),
    .din1(ffc_291_n_spl_0),
    .din2(g648_p_spl_)
  );


  LA
  g_g654_p
  (
    .dout(g654_p),
    .din1(g652_n_spl_0),
    .din2(g653_n_spl_)
  );


  FA
  g_g654_n
  (
    .dout(g654_n),
    .din1(g652_p_spl_),
    .din2(g653_p_spl_)
  );


  LA
  g_g655_p
  (
    .dout(g655_p),
    .din1(g652_p_spl_),
    .din2(g653_p_spl_)
  );


  FA
  g_g655_n
  (
    .dout(g655_n),
    .din1(g652_n_spl_0),
    .din2(g653_n_spl_)
  );


  LA
  g_g656_p
  (
    .dout(g656_p),
    .din1(g654_n),
    .din2(g655_n)
  );


  FA
  g_g656_n
  (
    .dout(g656_n),
    .din1(g654_p),
    .din2(g655_p)
  );


  FA
  g_g657_n
  (
    .dout(g657_n),
    .din1(ffc_332_p_spl_0),
    .din2(ffc_333_p_spl_0)
  );


  LA
  g_g658_p
  (
    .dout(g658_p),
    .din1(ffc_334_n),
    .din2(ffc_335_n_spl_)
  );


  FA
  g_g658_n
  (
    .dout(g658_n),
    .din1(ffc_334_p_spl_),
    .din2(ffc_335_p_spl_0)
  );


  FA
  g_g659_n
  (
    .dout(g659_n),
    .din1(ffc_336_p_spl_),
    .din2(ffc_337_p_spl_)
  );


  LA
  g_g660_p
  (
    .dout(g660_p),
    .din1(ffc_129_n_spl_),
    .din2(g599_n_spl_0)
  );


  FA
  g_g661_n
  (
    .dout(g661_n),
    .din1(ffc_131_p_spl_),
    .din2(g597_p_spl_0)
  );


  FA
  g_g662_n
  (
    .dout(g662_n),
    .din1(ffc_139_n),
    .din2(g598_p_spl_)
  );


  LA
  g_g663_p
  (
    .dout(g663_p),
    .din1(ffc_150_n_spl_),
    .din2(g597_n_spl_0)
  );


  FA
  g_g664_n
  (
    .dout(g664_n),
    .din1(ffc_151_p_spl_00),
    .din2(g595_p_spl_)
  );


  FA
  g_g665_n
  (
    .dout(g665_n),
    .din1(ffc_17_p_spl_0),
    .din2(ffc_197_p_spl_0)
  );


  LA
  g_g666_p
  (
    .dout(g666_p),
    .din1(g572_p_spl_0),
    .din2(g592_n_spl_)
  );


  FA
  g_g667_n
  (
    .dout(g667_n),
    .din1(ffc_357_p_spl_00),
    .din2(g657_n_spl_)
  );


  LA
  g_g668_p
  (
    .dout(g668_p),
    .din1(ffc_338_n),
    .din2(ffc_353_n_spl_)
  );


  FA
  g_g668_n
  (
    .dout(g668_n),
    .din1(ffc_338_p),
    .din2(ffc_353_p)
  );


  LA
  g_g669_p
  (
    .dout(g669_p),
    .din1(ffc_245_p_spl_00),
    .din2(g668_n_spl_0)
  );


  FA
  g_g669_n
  (
    .dout(g669_n),
    .din1(ffc_245_n_spl_0),
    .din2(g668_p_spl_0)
  );


  LA
  g_g670_p
  (
    .dout(g670_p),
    .din1(ffc_245_n_spl_0),
    .din2(ffc_315_n_spl_0)
  );


  FA
  g_g670_n
  (
    .dout(g670_n),
    .din1(ffc_245_p_spl_00),
    .din2(ffc_315_p_spl_00)
  );


  LA
  g_g671_p
  (
    .dout(g671_p),
    .din1(g669_n),
    .din2(g670_n)
  );


  FA
  g_g671_n
  (
    .dout(g671_n),
    .din1(g669_p),
    .din2(g670_p)
  );


  LA
  g_g672_p
  (
    .dout(g672_p),
    .din1(ffc_339_n_spl_0),
    .din2(ffc_357_n_spl_0)
  );


  FA
  g_g672_n
  (
    .dout(g672_n),
    .din1(ffc_339_p_spl_0),
    .din2(ffc_357_p_spl_0)
  );


  LA
  g_g673_p
  (
    .dout(g673_p),
    .din1(ffc_341_n),
    .din2(ffc_345_n)
  );


  FA
  g_g673_n
  (
    .dout(g673_n),
    .din1(ffc_341_p),
    .din2(ffc_345_p)
  );


  LA
  g_g674_p
  (
    .dout(g674_p),
    .din1(g672_n),
    .din2(g673_p)
  );


  FA
  g_g674_n
  (
    .dout(g674_n),
    .din1(g672_p),
    .din2(g673_n)
  );


  LA
  g_g675_p
  (
    .dout(g675_p),
    .din1(ffc_323_p_spl_000),
    .din2(g674_n)
  );


  FA
  g_g675_n
  (
    .dout(g675_n),
    .din1(ffc_323_n_spl_00),
    .din2(g674_p)
  );


  LA
  g_g676_p
  (
    .dout(g676_p),
    .din1(g671_n),
    .din2(g675_n)
  );


  FA
  g_g676_n
  (
    .dout(g676_n),
    .din1(g671_p),
    .din2(g675_p)
  );


  LA
  g_g677_p
  (
    .dout(g677_p),
    .din1(ffc_246_p_spl_0),
    .din2(g668_n_spl_0)
  );


  FA
  g_g677_n
  (
    .dout(g677_n),
    .din1(ffc_246_n_spl_0),
    .din2(g668_p_spl_0)
  );


  LA
  g_g678_p
  (
    .dout(g678_p),
    .din1(ffc_246_n_spl_0),
    .din2(ffc_315_n_spl_0)
  );


  FA
  g_g678_n
  (
    .dout(g678_n),
    .din1(ffc_246_p_spl_0),
    .din2(ffc_315_p_spl_00)
  );


  LA
  g_g679_p
  (
    .dout(g679_p),
    .din1(g677_n),
    .din2(g678_n)
  );


  FA
  g_g679_n
  (
    .dout(g679_n),
    .din1(g677_p),
    .din2(g678_p)
  );


  LA
  g_g680_p
  (
    .dout(g680_p),
    .din1(ffc_340_n_spl_0),
    .din2(ffc_358_p_spl_00)
  );


  FA
  g_g680_n
  (
    .dout(g680_n),
    .din1(ffc_340_p),
    .din2(ffc_358_n_spl_)
  );


  LA
  g_g681_p
  (
    .dout(g681_p),
    .din1(ffc_342_n),
    .din2(ffc_346_n)
  );


  FA
  g_g681_n
  (
    .dout(g681_n),
    .din1(ffc_342_p),
    .din2(ffc_346_p)
  );


  LA
  g_g682_p
  (
    .dout(g682_p),
    .din1(g680_n),
    .din2(g681_p)
  );


  FA
  g_g682_n
  (
    .dout(g682_n),
    .din1(g680_p),
    .din2(g681_n)
  );


  LA
  g_g683_p
  (
    .dout(g683_p),
    .din1(ffc_323_p_spl_000),
    .din2(g682_n)
  );


  FA
  g_g683_n
  (
    .dout(g683_n),
    .din1(ffc_323_n_spl_00),
    .din2(g682_p)
  );


  LA
  g_g684_p
  (
    .dout(g684_p),
    .din1(g679_n),
    .din2(g683_n)
  );


  FA
  g_g684_n
  (
    .dout(g684_n),
    .din1(g679_p),
    .din2(g683_p)
  );


  FA
  g_g685_n
  (
    .dout(g685_n),
    .din1(ffc_333_n_spl_0),
    .din2(ffc_357_n_spl_0)
  );


  LA
  g_g686_p
  (
    .dout(g686_p),
    .din1(g646_n_spl_),
    .din2(g685_n)
  );


  FA
  g_g687_n
  (
    .dout(g687_n),
    .din1(ffc_201_p_spl_0),
    .din2(ffc_242_p_spl_)
  );


  LA
  g_g688_p
  (
    .dout(g688_p),
    .din1(ffc_348_n_spl_00),
    .din2(ffc_360_p)
  );


  FA
  g_g688_n
  (
    .dout(g688_n),
    .din1(ffc_348_p_spl_00),
    .din2(ffc_360_n)
  );


  LA
  g_g689_p
  (
    .dout(g689_p),
    .din1(ffc_244_n),
    .din2(ffc_301_n)
  );


  FA
  g_g689_n
  (
    .dout(g689_n),
    .din1(ffc_244_p_spl_),
    .din2(ffc_301_p_spl_)
  );


  LA
  g_g690_p
  (
    .dout(g690_p),
    .din1(ffc_201_n),
    .din2(g689_n)
  );


  FA
  g_g690_n
  (
    .dout(g690_n),
    .din1(ffc_201_p_spl_0),
    .din2(g689_p)
  );


  LA
  g_g691_p
  (
    .dout(g691_p),
    .din1(g688_p_spl_0),
    .din2(g690_p_spl_0)
  );


  FA
  g_g691_n
  (
    .dout(g691_n),
    .din1(g688_n_spl_0),
    .din2(g690_n_spl_0)
  );


  LA
  g_g692_p
  (
    .dout(g692_p),
    .din1(ffc_202_p_spl_00),
    .din2(ffc_323_p_spl_00)
  );


  FA
  g_g692_n
  (
    .dout(g692_n),
    .din1(ffc_202_n_spl_),
    .din2(ffc_323_n_spl_0)
  );


  LA
  g_g693_p
  (
    .dout(g693_p),
    .din1(ffc_315_n_spl_1),
    .din2(g692_n_spl_)
  );


  FA
  g_g693_n
  (
    .dout(g693_n),
    .din1(ffc_315_p_spl_01),
    .din2(g692_p_spl_0)
  );


  LA
  g_g694_p
  (
    .dout(g694_p),
    .din1(ffc_247_n_spl_0),
    .din2(g693_n_spl_)
  );


  FA
  g_g694_n
  (
    .dout(g694_n),
    .din1(ffc_247_p_spl_0),
    .din2(g693_p)
  );


  LA
  g_g695_p
  (
    .dout(g695_p),
    .din1(ffc_245_n_spl_1),
    .din2(ffc_339_n_spl_0)
  );


  FA
  g_g695_n
  (
    .dout(g695_n),
    .din1(ffc_245_p_spl_0),
    .din2(ffc_339_p_spl_0)
  );


  LA
  g_g696_p
  (
    .dout(g696_p),
    .din1(ffc_248_p_spl_0),
    .din2(ffc_314_p_spl_0)
  );


  FA
  g_g696_n
  (
    .dout(g696_n),
    .din1(ffc_248_n_spl_0),
    .din2(ffc_314_n_spl_)
  );


  LA
  g_g697_p
  (
    .dout(g697_p),
    .din1(g695_n),
    .din2(g696_n)
  );


  FA
  g_g697_n
  (
    .dout(g697_n),
    .din1(g695_p),
    .din2(g696_p)
  );


  LA
  g_g698_p
  (
    .dout(g698_p),
    .din1(ffc_323_p_spl_01),
    .din2(g697_n)
  );


  FA
  g_g698_n
  (
    .dout(g698_n),
    .din1(ffc_323_n_spl_1),
    .din2(g697_p)
  );


  LA
  g_g699_p
  (
    .dout(g699_p),
    .din1(ffc_247_p_spl_0),
    .din2(g668_p_spl_1)
  );


  FA
  g_g699_n
  (
    .dout(g699_n),
    .din1(ffc_247_n_spl_0),
    .din2(g668_n_spl_1)
  );


  LA
  g_g700_p
  (
    .dout(g700_p),
    .din1(g698_n),
    .din2(g699_n)
  );


  FA
  g_g700_n
  (
    .dout(g700_n),
    .din1(g698_p),
    .din2(g699_p)
  );


  LA
  g_g701_p
  (
    .dout(g701_p),
    .din1(g694_n),
    .din2(g700_p)
  );


  FA
  g_g701_n
  (
    .dout(g701_n),
    .din1(g694_p),
    .din2(g700_n)
  );


  LA
  g_g702_p
  (
    .dout(g702_p),
    .din1(ffc_278_n),
    .din2(g688_p_spl_0)
  );


  FA
  g_g702_n
  (
    .dout(g702_n),
    .din1(ffc_278_p),
    .din2(g688_n_spl_0)
  );


  LA
  g_g703_p
  (
    .dout(g703_p),
    .din1(ffc_350_n),
    .din2(ffc_356_n)
  );


  FA
  g_g703_n
  (
    .dout(g703_n),
    .din1(ffc_350_p),
    .din2(ffc_356_p)
  );


  LA
  g_g704_p
  (
    .dout(g704_p),
    .din1(ffc_348_n_spl_00),
    .din2(g703_n)
  );


  FA
  g_g704_n
  (
    .dout(g704_n),
    .din1(ffc_348_p_spl_00),
    .din2(g703_p)
  );


  LA
  g_g705_p
  (
    .dout(g705_p),
    .din1(g702_n),
    .din2(g704_n)
  );


  FA
  g_g705_n
  (
    .dout(g705_n),
    .din1(g702_p),
    .din2(g704_p)
  );


  FA
  g_g706_n
  (
    .dout(g706_n),
    .din1(g658_p_spl_0),
    .din2(g705_n_spl_)
  );


  FA
  g_g707_n
  (
    .dout(g707_n),
    .din1(g676_p),
    .din2(g706_n)
  );


  LA
  g_g708_p
  (
    .dout(g708_p),
    .din1(ffc_324_n_spl_0),
    .din2(g688_p_spl_)
  );


  FA
  g_g708_n
  (
    .dout(g708_n),
    .din1(ffc_324_p_spl_0),
    .din2(g688_n_spl_)
  );


  LA
  g_g709_p
  (
    .dout(g709_p),
    .din1(ffc_349_n),
    .din2(ffc_355_n)
  );


  FA
  g_g709_n
  (
    .dout(g709_n),
    .din1(ffc_349_p),
    .din2(ffc_355_p)
  );


  LA
  g_g710_p
  (
    .dout(g710_p),
    .din1(ffc_348_n_spl_01),
    .din2(g709_n)
  );


  FA
  g_g710_n
  (
    .dout(g710_n),
    .din1(ffc_348_p_spl_01),
    .din2(g709_p)
  );


  LA
  g_g711_p
  (
    .dout(g711_p),
    .din1(g708_n_spl_0),
    .din2(g710_n)
  );


  FA
  g_g711_n
  (
    .dout(g711_n),
    .din1(g708_p_spl_0),
    .din2(g710_p)
  );


  FA
  g_g712_n
  (
    .dout(g712_n),
    .din1(g658_p_spl_0),
    .din2(g711_n_spl_)
  );


  FA
  g_g713_n
  (
    .dout(g713_n),
    .din1(g684_p),
    .din2(g712_n)
  );


  FA
  g_g714_n
  (
    .dout(g714_n),
    .din1(ffc_149_n),
    .din2(g609_n_spl_1)
  );


  FA
  g_g715_n
  (
    .dout(g715_n),
    .din1(ffc_148_n_spl_),
    .din2(g609_n_spl_1)
  );


  LA
  g_g716_p
  (
    .dout(g716_p),
    .din1(ffc_127_p_spl_0),
    .din2(g661_n_spl_)
  );


  FA
  g_g717_n
  (
    .dout(g717_n),
    .din1(ffc_70_n_spl_00),
    .din2(ffc_254_p_spl_)
  );


  FA
  g_g718_n
  (
    .dout(g718_n),
    .din1(ffc_236_n_spl_),
    .din2(g717_n_spl_0)
  );


  FA
  g_g719_n
  (
    .dout(g719_n),
    .din1(ffc_150_p_spl_0),
    .din2(g595_p_spl_)
  );


  FA
  g_g720_n
  (
    .dout(g720_n),
    .din1(ffc_151_p_spl_00),
    .din2(g599_p_spl_)
  );


  LA
  g_g721_p
  (
    .dout(g721_p),
    .din1(g601_p_spl_),
    .din2(g603_p_spl_)
  );


  LA
  g_g722_p
  (
    .dout(g722_p),
    .din1(ffc_155_p_spl_0),
    .din2(ffc_236_n_spl_)
  );


  FA
  g_g722_n
  (
    .dout(g722_n),
    .din1(ffc_155_n_spl_0),
    .din2(ffc_236_p_spl_)
  );


  LA
  g_g723_p
  (
    .dout(g723_p),
    .din1(ffc_221_p),
    .din2(ffc_235_p_spl_)
  );


  FA
  g_g723_n
  (
    .dout(g723_n),
    .din1(ffc_221_n),
    .din2(ffc_235_n_spl_0)
  );


  LA
  g_g724_p
  (
    .dout(g724_p),
    .din1(ffc_289_p_spl_),
    .din2(g723_n)
  );


  FA
  g_g724_n
  (
    .dout(g724_n),
    .din1(ffc_289_n_spl_),
    .din2(g723_p)
  );


  LA
  g_g725_p
  (
    .dout(g725_p),
    .din1(g722_n_spl_),
    .din2(g724_n_spl_)
  );


  FA
  g_g725_n
  (
    .dout(g725_n),
    .din1(g722_p_spl_0),
    .din2(g724_p_spl_)
  );


  LA
  g_g726_p
  (
    .dout(g726_p),
    .din1(g722_p_spl_0),
    .din2(g724_p_spl_)
  );


  FA
  g_g726_n
  (
    .dout(g726_n),
    .din1(g722_n_spl_),
    .din2(g724_n_spl_)
  );


  LA
  g_g727_p
  (
    .dout(g727_p),
    .din1(g725_n),
    .din2(g726_n)
  );


  FA
  g_g727_n
  (
    .dout(g727_n),
    .din1(g725_p),
    .din2(g726_p)
  );


  LA
  g_g728_p
  (
    .dout(g728_p),
    .din1(ffc_120_n_spl_),
    .din2(ffc_264_n_spl_)
  );


  FA
  g_g728_n
  (
    .dout(g728_n),
    .din1(ffc_120_p_spl_),
    .din2(ffc_264_p_spl_)
  );


  LA
  g_g729_p
  (
    .dout(g729_p),
    .din1(ffc_120_p_spl_),
    .din2(ffc_264_p_spl_)
  );


  FA
  g_g729_n
  (
    .dout(g729_n),
    .din1(ffc_120_n_spl_),
    .din2(ffc_264_n_spl_)
  );


  LA
  g_g730_p
  (
    .dout(g730_p),
    .din1(g728_n),
    .din2(g729_n)
  );


  FA
  g_g730_n
  (
    .dout(g730_n),
    .din1(g728_p),
    .din2(g729_p)
  );


  LA
  g_g731_p
  (
    .dout(g731_p),
    .din1(ffc_265_n),
    .din2(ffc_289_p_spl_)
  );


  FA
  g_g731_n
  (
    .dout(g731_n),
    .din1(ffc_265_p),
    .din2(ffc_289_n_spl_)
  );


  LA
  g_g732_p
  (
    .dout(g732_p),
    .din1(g553_n_spl_),
    .din2(g731_n_spl_)
  );


  FA
  g_g732_n
  (
    .dout(g732_n),
    .din1(g553_p_spl_0),
    .din2(g731_p_spl_)
  );


  LA
  g_g733_p
  (
    .dout(g733_p),
    .din1(g730_p_spl_0),
    .din2(g732_p_spl_)
  );


  FA
  g_g733_n
  (
    .dout(g733_n),
    .din1(g730_n_spl_00),
    .din2(g732_n_spl_)
  );


  LA
  g_g734_p
  (
    .dout(g734_p),
    .din1(g730_n_spl_00),
    .din2(g732_n_spl_)
  );


  FA
  g_g734_n
  (
    .dout(g734_n),
    .din1(g730_p_spl_0),
    .din2(g732_p_spl_)
  );


  LA
  g_g735_p
  (
    .dout(g735_p),
    .din1(g733_n),
    .din2(g734_n)
  );


  FA
  g_g735_n
  (
    .dout(g735_n),
    .din1(g733_p),
    .din2(g734_p)
  );


  FA
  g_g736_n
  (
    .dout(g736_n),
    .din1(g727_p_spl_),
    .din2(g735_p_spl_)
  );


  LA
  g_g737_p
  (
    .dout(g737_p),
    .din1(ffc_171_p_spl_0),
    .din2(g736_n)
  );


  FA
  g_g738_n
  (
    .dout(g738_n),
    .din1(g556_p_spl_0),
    .din2(g737_p)
  );


  LA
  g_g739_p
  (
    .dout(g739_p),
    .din1(g561_p_spl_),
    .din2(g738_n)
  );


  LA
  g_g740_p
  (
    .dout(g740_p),
    .din1(g561_n_spl_01),
    .din2(g727_n_spl_0)
  );


  LA
  g_g741_p
  (
    .dout(g741_p),
    .din1(g561_n_spl_1),
    .din2(g735_n_spl_)
  );


  LA
  g_g742_p
  (
    .dout(g742_p),
    .din1(ffc_155_n_spl_1),
    .din2(ffc_236_p_spl_)
  );


  FA
  g_g743_n
  (
    .dout(g743_n),
    .din1(g722_p_spl_),
    .din2(g742_p)
  );


  LA
  g_g744_p
  (
    .dout(g744_p),
    .din1(ffc_70_n_spl_01),
    .din2(ffc_118_n_spl_)
  );


  FA
  g_g744_n
  (
    .dout(g744_n),
    .din1(ffc_70_p_spl_00),
    .din2(ffc_118_p_spl_0)
  );


  FA
  g_g745_n
  (
    .dout(g745_n),
    .din1(ffc_75_n_spl_0),
    .din2(g744_p)
  );


  LA
  g_g746_p
  (
    .dout(g746_p),
    .din1(ffc_71_n_spl_),
    .din2(g559_n_spl_)
  );


  LA
  g_g747_p
  (
    .dout(g747_p),
    .din1(ffc_71_p_spl_),
    .din2(g551_n_spl_)
  );


  FA
  g_g748_n
  (
    .dout(g748_n),
    .din1(g552_n_spl_),
    .din2(g744_n)
  );


  FA
  g_g749_n
  (
    .dout(g749_n),
    .din1(g747_p),
    .din2(g748_n)
  );


  FA
  g_g750_n
  (
    .dout(g750_n),
    .din1(g746_p),
    .din2(g749_n)
  );


  LA
  g_g751_p
  (
    .dout(g751_p),
    .din1(g745_n),
    .din2(g750_n)
  );


  FA
  g_g752_n
  (
    .dout(g752_n),
    .din1(g612_n_spl_),
    .din2(g751_p)
  );


  FA
  g_g753_n
  (
    .dout(g753_n),
    .din1(ffc_46_n),
    .din2(ffc_174_p_spl_00)
  );


  FA
  g_g754_n
  (
    .dout(g754_n),
    .din1(ffc_159_n_spl_0),
    .din2(ffc_252_n)
  );


  FA
  g_g755_n
  (
    .dout(g755_n),
    .din1(ffc_173_p_spl_0),
    .din2(ffc_204_n)
  );


  LA
  g_g756_p
  (
    .dout(g756_p),
    .din1(g754_n),
    .din2(g755_n)
  );


  LA
  g_g757_p
  (
    .dout(g757_p),
    .din1(g753_n),
    .din2(g756_p)
  );


  FA
  g_g758_n
  (
    .dout(g758_n),
    .din1(ffc_78_n),
    .din2(ffc_173_p_spl_0)
  );


  FA
  g_g759_n
  (
    .dout(g759_n),
    .din1(ffc_174_p_spl_00),
    .din2(ffc_203_n)
  );


  LA
  g_g760_p
  (
    .dout(g760_p),
    .din1(g758_n),
    .din2(g759_n)
  );


  FA
  g_g761_n
  (
    .dout(g761_n),
    .din1(ffc_89_n_spl_),
    .din2(ffc_175_p_spl_0)
  );


  LA
  g_g762_p
  (
    .dout(g762_p),
    .din1(ffc_70_p_spl_00),
    .din2(g761_n)
  );


  FA
  g_g763_n
  (
    .dout(g763_n),
    .din1(ffc_158_p_spl_0),
    .din2(ffc_253_n)
  );


  FA
  g_g764_n
  (
    .dout(g764_n),
    .din1(ffc_83_n_spl_),
    .din2(ffc_172_n_spl_0)
  );


  LA
  g_g765_p
  (
    .dout(g765_p),
    .din1(g763_n),
    .din2(g764_n)
  );


  LA
  g_g766_p
  (
    .dout(g766_p),
    .din1(g762_p),
    .din2(g765_p)
  );


  LA
  g_g767_p
  (
    .dout(g767_p),
    .din1(g760_p_spl_),
    .din2(g766_p)
  );


  LA
  g_g768_p
  (
    .dout(g768_p),
    .din1(g757_p),
    .din2(g767_p)
  );


  FA
  g_g769_n
  (
    .dout(g769_n),
    .din1(ffc_104_p_spl_0),
    .din2(ffc_159_n_spl_0)
  );


  LA
  g_g770_p
  (
    .dout(g770_p),
    .din1(ffc_186_p),
    .din2(g769_n)
  );


  FA
  g_g771_n
  (
    .dout(g771_n),
    .din1(ffc_73_p_spl_),
    .din2(ffc_172_n_spl_0)
  );


  LA
  g_g772_p
  (
    .dout(g772_p),
    .din1(ffc_184_p),
    .din2(g771_n_spl_)
  );


  LA
  g_g773_p
  (
    .dout(g773_p),
    .din1(g770_p),
    .din2(g772_p)
  );


  FA
  g_g774_n
  (
    .dout(g774_n),
    .din1(ffc_174_p_spl_0),
    .din2(ffc_261_p)
  );


  LA
  g_g775_p
  (
    .dout(g775_p),
    .din1(ffc_70_n_spl_01),
    .din2(g774_n)
  );


  FA
  g_g776_n
  (
    .dout(g776_n),
    .din1(ffc_103_p_spl_0),
    .din2(ffc_158_p_spl_0)
  );


  LA
  g_g777_p
  (
    .dout(g777_p),
    .din1(ffc_183_p),
    .din2(g776_n)
  );


  LA
  g_g778_p
  (
    .dout(g778_p),
    .din1(g775_p),
    .din2(g777_p)
  );


  LA
  g_g779_p
  (
    .dout(g779_p),
    .din1(g773_p),
    .din2(g778_p)
  );


  FA
  g_g780_n
  (
    .dout(g780_n),
    .din1(g612_p_spl_01),
    .din2(g779_p)
  );


  FA
  g_g781_n
  (
    .dout(g781_n),
    .din1(g768_p),
    .din2(g780_n)
  );


  LA
  g_g782_p
  (
    .dout(g782_p),
    .din1(g752_n),
    .din2(g781_n)
  );


  FA
  g_g783_n
  (
    .dout(g783_n),
    .din1(g562_n_spl_),
    .din2(g782_p)
  );


  FA
  g_g784_n
  (
    .dout(g784_n),
    .din1(ffc_75_p_spl_),
    .din2(ffc_174_p_spl_1)
  );


  FA
  g_g785_n
  (
    .dout(g785_n),
    .din1(ffc_72_p_spl_),
    .din2(ffc_173_p_spl_1)
  );


  FA
  g_g786_n
  (
    .dout(g786_n),
    .din1(ffc_89_n_spl_),
    .din2(ffc_158_p_spl_1)
  );


  LA
  g_g787_p
  (
    .dout(g787_p),
    .din1(g785_n),
    .din2(g786_n)
  );


  LA
  g_g788_p
  (
    .dout(g788_p),
    .din1(g784_n),
    .din2(g787_p)
  );


  LA
  g_g789_p
  (
    .dout(g789_p),
    .din1(ffc_70_p_spl_01),
    .din2(g771_n_spl_)
  );


  FA
  g_g790_n
  (
    .dout(g790_n),
    .din1(ffc_74_p_spl_),
    .din2(ffc_175_p_spl_0)
  );


  FA
  g_g791_n
  (
    .dout(g791_n),
    .din1(ffc_83_n_spl_),
    .din2(ffc_159_n_spl_1)
  );


  LA
  g_g792_p
  (
    .dout(g792_p),
    .din1(g790_n),
    .din2(g791_n)
  );


  LA
  g_g793_p
  (
    .dout(g793_p),
    .din1(g789_p),
    .din2(g792_p)
  );


  LA
  g_g794_p
  (
    .dout(g794_p),
    .din1(g760_p_spl_),
    .din2(g793_p)
  );


  LA
  g_g795_p
  (
    .dout(g795_p),
    .din1(g788_p),
    .din2(g794_p)
  );


  FA
  g_g796_n
  (
    .dout(g796_n),
    .din1(ffc_104_p_spl_0),
    .din2(ffc_172_n_spl_)
  );


  FA
  g_g797_n
  (
    .dout(g797_n),
    .din1(ffc_153_n),
    .din2(ffc_158_p_spl_1)
  );


  FA
  g_g798_n
  (
    .dout(g798_n),
    .din1(ffc_154_n),
    .din2(ffc_159_n_spl_1)
  );


  LA
  g_g799_p
  (
    .dout(g799_p),
    .din1(g797_n),
    .din2(g798_n)
  );


  LA
  g_g800_p
  (
    .dout(g800_p),
    .din1(g796_n),
    .din2(g799_p)
  );


  FA
  g_g801_n
  (
    .dout(g801_n),
    .din1(ffc_174_p_spl_1),
    .din2(ffc_188_n)
  );


  LA
  g_g802_p
  (
    .dout(g802_p),
    .din1(ffc_70_n_spl_10),
    .din2(g801_n)
  );


  FA
  g_g803_n
  (
    .dout(g803_n),
    .din1(ffc_103_p_spl_1),
    .din2(ffc_175_p_spl_)
  );


  FA
  g_g804_n
  (
    .dout(g804_n),
    .din1(ffc_173_p_spl_1),
    .din2(ffc_260_p)
  );


  LA
  g_g805_p
  (
    .dout(g805_p),
    .din1(g803_n),
    .din2(g804_n)
  );


  LA
  g_g806_p
  (
    .dout(g806_p),
    .din1(g802_p),
    .din2(g805_p)
  );


  LA
  g_g807_p
  (
    .dout(g807_p),
    .din1(g800_p),
    .din2(g806_p)
  );


  FA
  g_g808_n
  (
    .dout(g808_n),
    .din1(g795_p),
    .din2(g807_p)
  );


  LA
  g_g809_p
  (
    .dout(g809_p),
    .din1(g612_n_spl_),
    .din2(g808_n)
  );


  FA
  g_g810_n
  (
    .dout(g810_n),
    .din1(g562_n_spl_),
    .din2(g809_p)
  );


  LA
  g_g811_p
  (
    .dout(g811_p),
    .din1(ffc_74_n_spl_),
    .din2(ffc_172_p_spl_00)
  );


  LA
  g_g812_p
  (
    .dout(g812_p),
    .din1(ffc_158_n_spl_00),
    .din2(ffc_203_p)
  );


  FA
  g_g813_n
  (
    .dout(g813_n),
    .din1(ffc_78_p_spl_0),
    .din2(ffc_204_p_spl_)
  );


  LA
  g_g814_p
  (
    .dout(g814_p),
    .din1(ffc_174_n_spl_000),
    .din2(g813_n)
  );


  FA
  g_g815_n
  (
    .dout(g815_n),
    .din1(g812_p),
    .din2(g814_p)
  );


  FA
  g_g816_n
  (
    .dout(g816_n),
    .din1(g811_p),
    .din2(g815_n)
  );


  FA
  g_g817_n
  (
    .dout(g817_n),
    .din1(ffc_73_n_spl_),
    .din2(ffc_83_p_spl_0)
  );


  LA
  g_g818_p
  (
    .dout(g818_p),
    .din1(ffc_173_n_spl_00),
    .din2(g817_n)
  );


  FA
  g_g819_n
  (
    .dout(g819_n),
    .din1(ffc_70_n_spl_10),
    .din2(g818_p)
  );


  LA
  g_g820_p
  (
    .dout(g820_p),
    .din1(ffc_75_n_spl_0),
    .din2(ffc_175_n_spl_00)
  );


  LA
  g_g821_p
  (
    .dout(g821_p),
    .din1(ffc_89_p_spl_),
    .din2(ffc_159_p_spl_00)
  );


  FA
  g_g822_n
  (
    .dout(g822_n),
    .din1(g820_p),
    .din2(g821_p)
  );


  FA
  g_g823_n
  (
    .dout(g823_n),
    .din1(g819_n),
    .din2(g822_n)
  );


  FA
  g_g824_n
  (
    .dout(g824_n),
    .din1(g816_n),
    .din2(g823_n)
  );


  LA
  g_g825_p
  (
    .dout(g825_p),
    .din1(ffc_112_p_spl_0),
    .din2(ffc_159_p_spl_00)
  );


  LA
  g_g826_p
  (
    .dout(g826_p),
    .din1(ffc_154_p),
    .din2(ffc_158_n_spl_00)
  );


  LA
  g_g827_p
  (
    .dout(g827_p),
    .din1(ffc_173_n_spl_00),
    .din2(ffc_261_n)
  );


  FA
  g_g828_n
  (
    .dout(g828_n),
    .din1(g826_p),
    .din2(g827_p)
  );


  FA
  g_g829_n
  (
    .dout(g829_n),
    .din1(g825_p),
    .din2(g828_n)
  );


  LA
  g_g830_p
  (
    .dout(g830_p),
    .din1(ffc_170_n),
    .din2(ffc_174_n_spl_000)
  );


  FA
  g_g831_n
  (
    .dout(g831_n),
    .din1(ffc_70_p_spl_01),
    .din2(g830_p)
  );


  LA
  g_g832_p
  (
    .dout(g832_p),
    .din1(ffc_104_n),
    .din2(ffc_175_n_spl_00)
  );


  FA
  g_g833_n
  (
    .dout(g833_n),
    .din1(ffc_209_p),
    .din2(g832_p)
  );


  FA
  g_g834_n
  (
    .dout(g834_n),
    .din1(g831_n),
    .din2(g833_n)
  );


  FA
  g_g835_n
  (
    .dout(g835_n),
    .din1(g829_n),
    .din2(g834_n)
  );


  LA
  g_g836_p
  (
    .dout(g836_p),
    .din1(g824_n),
    .din2(g835_n)
  );


  FA
  g_g837_n
  (
    .dout(g837_n),
    .din1(g612_p_spl_01),
    .din2(g836_p)
  );


  LA
  g_g838_p
  (
    .dout(g838_p),
    .din1(g562_p_spl_01),
    .din2(g837_n)
  );


  LA
  g_g839_p
  (
    .dout(g839_p),
    .din1(ffc_74_n_spl_),
    .din2(ffc_174_n_spl_00)
  );


  LA
  g_g840_p
  (
    .dout(g840_p),
    .din1(ffc_78_p_spl_0),
    .din2(ffc_159_p_spl_01)
  );


  FA
  g_g841_n
  (
    .dout(g841_n),
    .din1(g839_p),
    .din2(g840_p)
  );


  LA
  g_g842_p
  (
    .dout(g842_p),
    .din1(ffc_83_p_spl_0),
    .din2(ffc_158_n_spl_01)
  );


  FA
  g_g843_n
  (
    .dout(g843_n),
    .din1(ffc_75_n_spl_1),
    .din2(ffc_94_n)
  );


  LA
  g_g844_p
  (
    .dout(g844_p),
    .din1(ffc_173_n_spl_01),
    .din2(g843_n)
  );


  FA
  g_g845_n
  (
    .dout(g845_n),
    .din1(g842_p),
    .din2(g844_p)
  );


  FA
  g_g846_n
  (
    .dout(g846_n),
    .din1(g841_n),
    .din2(g845_n)
  );


  LA
  g_g847_p
  (
    .dout(g847_p),
    .din1(ffc_89_p_spl_),
    .din2(ffc_174_n_spl_01)
  );


  FA
  g_g848_n
  (
    .dout(g848_n),
    .din1(ffc_70_n_spl_1),
    .din2(g847_p)
  );


  LA
  g_g849_p
  (
    .dout(g849_p),
    .din1(ffc_72_n_spl_),
    .din2(ffc_172_p_spl_00)
  );


  LA
  g_g850_p
  (
    .dout(g850_p),
    .din1(ffc_73_n_spl_),
    .din2(ffc_175_n_spl_01)
  );


  FA
  g_g851_n
  (
    .dout(g851_n),
    .din1(g849_p_spl_),
    .din2(g850_p)
  );


  FA
  g_g852_n
  (
    .dout(g852_n),
    .din1(g848_n_spl_),
    .din2(g851_n)
  );


  FA
  g_g853_n
  (
    .dout(g853_n),
    .din1(g846_n),
    .din2(g852_n)
  );


  FA
  g_g854_n
  (
    .dout(g854_n),
    .din1(ffc_112_p_spl_0),
    .din2(ffc_168_p)
  );


  LA
  g_g855_p
  (
    .dout(g855_p),
    .din1(ffc_174_n_spl_01),
    .din2(g854_n)
  );


  LA
  g_g856_p
  (
    .dout(g856_p),
    .din1(ffc_113_p_spl_0),
    .din2(ffc_175_n_spl_01)
  );


  LA
  g_g857_p
  (
    .dout(g857_p),
    .din1(ffc_173_n_spl_01),
    .din2(ffc_262_n_spl_)
  );


  FA
  g_g858_n
  (
    .dout(g858_n),
    .din1(g856_p),
    .din2(g857_p)
  );


  FA
  g_g859_n
  (
    .dout(g859_n),
    .din1(g855_p),
    .din2(g858_n)
  );


  LA
  g_g860_p
  (
    .dout(g860_p),
    .din1(ffc_103_n_spl_),
    .din2(ffc_172_p_spl_0)
  );


  LA
  g_g861_p
  (
    .dout(g861_p),
    .din1(ffc_153_p),
    .din2(ffc_159_p_spl_01)
  );


  FA
  g_g862_n
  (
    .dout(g862_n),
    .din1(g860_p),
    .din2(g861_p)
  );


  LA
  g_g863_p
  (
    .dout(g863_p),
    .din1(ffc_158_n_spl_01),
    .din2(ffc_169_p)
  );


  FA
  g_g864_n
  (
    .dout(g864_n),
    .din1(ffc_70_p_spl_10),
    .din2(g863_p)
  );


  FA
  g_g865_n
  (
    .dout(g865_n),
    .din1(g862_n),
    .din2(g864_n)
  );


  FA
  g_g866_n
  (
    .dout(g866_n),
    .din1(g859_n),
    .din2(g865_n)
  );


  LA
  g_g867_p
  (
    .dout(g867_p),
    .din1(g853_n),
    .din2(g866_n)
  );


  FA
  g_g868_n
  (
    .dout(g868_n),
    .din1(g612_p_spl_10),
    .din2(g867_p)
  );


  LA
  g_g869_p
  (
    .dout(g869_p),
    .din1(g562_p_spl_01),
    .din2(g868_n)
  );


  LA
  g_g870_p
  (
    .dout(g870_p),
    .din1(ffc_110_p),
    .din2(ffc_122_p_spl_)
  );


  FA
  g_g870_n
  (
    .dout(g870_n),
    .din1(ffc_110_n),
    .din2(ffc_122_n_spl_)
  );


  LA
  g_g871_p
  (
    .dout(g871_p),
    .din1(ffc_119_n_spl_),
    .din2(g870_n_spl_)
  );


  FA
  g_g871_n
  (
    .dout(g871_n),
    .din1(ffc_119_p_spl_),
    .din2(g870_p_spl_)
  );


  LA
  g_g872_p
  (
    .dout(g872_p),
    .din1(ffc_119_p_spl_),
    .din2(g870_p_spl_)
  );


  FA
  g_g872_n
  (
    .dout(g872_n),
    .din1(ffc_119_n_spl_),
    .din2(g870_n_spl_)
  );


  LA
  g_g873_p
  (
    .dout(g873_p),
    .din1(g871_n),
    .din2(g872_n)
  );


  FA
  g_g873_n
  (
    .dout(g873_n),
    .din1(g871_p),
    .din2(g872_p)
  );


  FA
  g_g874_n
  (
    .dout(g874_n),
    .din1(g717_n_spl_0),
    .din2(g873_n_spl_0)
  );


  FA
  g_g875_n
  (
    .dout(g875_n),
    .din1(ffc_297_n_spl_),
    .din2(ffc_328_p_spl_010)
  );


  FA
  g_g876_n
  (
    .dout(g876_n),
    .din1(ffc_202_p_spl_00),
    .din2(g687_n_spl_)
  );


  LA
  g_g877_p
  (
    .dout(g877_p),
    .din1(ffc_307_n),
    .din2(ffc_317_n)
  );


  FA
  g_g877_n
  (
    .dout(g877_n),
    .din1(ffc_307_p),
    .din2(ffc_317_p)
  );


  LA
  g_g878_p
  (
    .dout(g878_p),
    .din1(ffc_195_n),
    .din2(ffc_309_n)
  );


  FA
  g_g878_n
  (
    .dout(g878_n),
    .din1(ffc_195_p),
    .din2(ffc_309_p)
  );


  FA
  g_g879_n
  (
    .dout(g879_n),
    .din1(ffc_182_n_spl_),
    .din2(g878_n_spl_)
  );


  LA
  g_g880_p
  (
    .dout(g880_p),
    .din1(g877_p_spl_0),
    .din2(g879_n)
  );


  LA
  g_g881_p
  (
    .dout(g881_p),
    .din1(ffc_181_p_spl_),
    .din2(g877_n)
  );


  FA
  g_g881_n
  (
    .dout(g881_n),
    .din1(ffc_181_n_spl_),
    .din2(g877_p_spl_0)
  );


  LA
  g_g882_p
  (
    .dout(g882_p),
    .din1(g878_p),
    .din2(g881_p)
  );


  FA
  g_g882_n
  (
    .dout(g882_n),
    .din1(g878_n_spl_),
    .din2(g881_n)
  );


  FA
  g_g883_n
  (
    .dout(g883_n),
    .din1(g880_p),
    .din2(g882_p)
  );


  FA
  g_g884_n
  (
    .dout(g884_n),
    .din1(g652_n_spl_),
    .din2(g883_n_spl_0)
  );


  FA
  g_g885_n
  (
    .dout(g885_n),
    .din1(g573_n_spl_),
    .din2(g884_n_spl_)
  );


  FA
  g_g886_n
  (
    .dout(g886_n),
    .din1(g568_n_spl_),
    .din2(g885_n_spl_)
  );


  FA
  g_g887_n
  (
    .dout(g887_n),
    .din1(ffc_171_n_spl_0),
    .din2(g727_n_spl_0)
  );


  LA
  g_g888_p
  (
    .dout(g888_p),
    .din1(ffc_171_n_spl_0),
    .din2(g727_n_spl_)
  );


  FA
  g_g888_n
  (
    .dout(g888_n),
    .din1(ffc_171_p_spl_0),
    .din2(g727_p_spl_)
  );


  LA
  g_g889_p
  (
    .dout(g889_p),
    .din1(g887_n),
    .din2(g888_n_spl_)
  );


  FA
  g_g890_n
  (
    .dout(g890_n),
    .din1(g577_n_spl_0),
    .din2(g656_n_spl_)
  );


  FA
  g_g891_n
  (
    .dout(g891_n),
    .din1(ffc_235_n_spl_),
    .din2(g717_n_spl_1)
  );


  LA
  g_g892_p
  (
    .dout(g892_p),
    .din1(ffc_158_n_spl_10),
    .din2(ffc_252_p_spl_)
  );


  LA
  g_g893_p
  (
    .dout(g893_p),
    .din1(ffc_78_p_spl_1),
    .din2(ffc_172_p_spl_1)
  );


  FA
  g_g894_n
  (
    .dout(g894_n),
    .din1(g892_p),
    .din2(g893_p)
  );


  LA
  g_g895_p
  (
    .dout(g895_p),
    .din1(ffc_173_n_spl_1),
    .din2(ffc_256_n)
  );


  LA
  g_g896_p
  (
    .dout(g896_p),
    .din1(ffc_159_p_spl_10),
    .din2(ffc_204_p_spl_)
  );


  FA
  g_g897_n
  (
    .dout(g897_n),
    .din1(g895_p),
    .din2(g896_p)
  );


  FA
  g_g898_n
  (
    .dout(g898_n),
    .din1(g894_n),
    .din2(g897_n)
  );


  LA
  g_g899_p
  (
    .dout(g899_p),
    .din1(ffc_83_p_spl_),
    .din2(ffc_175_n_spl_10)
  );


  LA
  g_g900_p
  (
    .dout(g900_p),
    .din1(ffc_174_n_spl_10),
    .din2(ffc_253_p)
  );


  FA
  g_g901_n
  (
    .dout(g901_n),
    .din1(g899_p),
    .din2(g900_p)
  );


  FA
  g_g902_n
  (
    .dout(g902_n),
    .din1(g848_n_spl_),
    .din2(g901_n)
  );


  FA
  g_g903_n
  (
    .dout(g903_n),
    .din1(g898_n),
    .din2(g902_n)
  );


  LA
  g_g904_p
  (
    .dout(g904_p),
    .din1(ffc_113_p_spl_0),
    .din2(ffc_158_n_spl_10)
  );


  LA
  g_g905_p
  (
    .dout(g905_p),
    .din1(ffc_174_n_spl_10),
    .din2(ffc_260_n)
  );


  FA
  g_g906_n
  (
    .dout(g906_n),
    .din1(g904_p),
    .din2(g905_p)
  );


  FA
  g_g907_n
  (
    .dout(g907_n),
    .din1(ffc_210_n),
    .din2(g906_n)
  );


  LA
  g_g908_p
  (
    .dout(g908_p),
    .din1(ffc_103_n_spl_),
    .din2(ffc_159_p_spl_10)
  );


  FA
  g_g909_n
  (
    .dout(g909_n),
    .din1(g849_p_spl_),
    .din2(g908_p)
  );


  FA
  g_g910_n
  (
    .dout(g910_n),
    .din1(ffc_70_p_spl_10),
    .din2(ffc_230_n)
  );


  FA
  g_g911_n
  (
    .dout(g911_n),
    .din1(g909_n),
    .din2(g910_n)
  );


  FA
  g_g912_n
  (
    .dout(g912_n),
    .din1(g907_n),
    .din2(g911_n)
  );


  LA
  g_g913_p
  (
    .dout(g913_p),
    .din1(g903_n),
    .din2(g912_n)
  );


  FA
  g_g914_n
  (
    .dout(g914_n),
    .din1(g612_p_spl_10),
    .din2(g913_p)
  );


  LA
  g_g915_p
  (
    .dout(g915_p),
    .din1(g562_p_spl_10),
    .din2(g914_n)
  );


  LA
  g_g916_p
  (
    .dout(g916_p),
    .din1(g891_n),
    .din2(g915_p)
  );


  LA
  g_g917_p
  (
    .dout(g917_p),
    .din1(g561_n_spl_1),
    .din2(g601_n_spl_)
  );


  LA
  g_g918_p
  (
    .dout(g918_p),
    .din1(g556_n_spl_1),
    .din2(g604_n_spl_)
  );


  FA
  g_g919_n
  (
    .dout(g919_n),
    .din1(g917_p),
    .din2(g918_p)
  );


  FA
  g_g920_n
  (
    .dout(g920_n),
    .din1(g717_n_spl_1),
    .din2(g730_n_spl_0)
  );


  LA
  g_g921_p
  (
    .dout(g921_p),
    .din1(ffc_93_n),
    .din2(ffc_175_n_spl_10)
  );


  LA
  g_g922_p
  (
    .dout(g922_p),
    .din1(ffc_112_p_spl_),
    .din2(ffc_158_n_spl_1)
  );


  LA
  g_g923_p
  (
    .dout(g923_p),
    .din1(ffc_113_p_spl_),
    .din2(ffc_159_p_spl_1)
  );


  FA
  g_g924_n
  (
    .dout(g924_n),
    .din1(g922_p),
    .din2(g923_p)
  );


  FA
  g_g925_n
  (
    .dout(g925_n),
    .din1(g921_p),
    .din2(g924_n)
  );


  LA
  g_g926_p
  (
    .dout(g926_p),
    .din1(ffc_174_n_spl_11),
    .din2(ffc_262_n_spl_)
  );


  FA
  g_g927_n
  (
    .dout(g927_n),
    .din1(ffc_70_p_spl_1),
    .din2(g926_p)
  );


  LA
  g_g928_p
  (
    .dout(g928_p),
    .din1(ffc_173_n_spl_1),
    .din2(ffc_255_n)
  );


  FA
  g_g929_n
  (
    .dout(g929_n),
    .din1(ffc_187_p),
    .din2(g928_p)
  );


  FA
  g_g930_n
  (
    .dout(g930_n),
    .din1(g927_n),
    .din2(g929_n)
  );


  FA
  g_g931_n
  (
    .dout(g931_n),
    .din1(g925_n),
    .din2(g930_n)
  );


  LA
  g_g932_p
  (
    .dout(g932_p),
    .din1(ffc_78_p_spl_1),
    .din2(ffc_175_n_spl_1)
  );


  LA
  g_g933_p
  (
    .dout(g933_p),
    .din1(ffc_174_n_spl_11),
    .din2(ffc_252_p_spl_)
  );


  LA
  g_g934_p
  (
    .dout(g934_p),
    .din1(ffc_75_n_spl_1),
    .din2(ffc_172_p_spl_1)
  );


  FA
  g_g935_n
  (
    .dout(g935_n),
    .din1(g933_p),
    .din2(g934_p)
  );


  FA
  g_g936_n
  (
    .dout(g936_n),
    .din1(g932_p),
    .din2(g935_n)
  );


  FA
  g_g937_n
  (
    .dout(g937_n),
    .din1(ffc_185_p),
    .din2(ffc_270_p)
  );


  FA
  g_g938_n
  (
    .dout(g938_n),
    .din1(ffc_258_p),
    .din2(ffc_271_p)
  );


  FA
  g_g939_n
  (
    .dout(g939_n),
    .din1(g937_n),
    .din2(g938_n)
  );


  FA
  g_g940_n
  (
    .dout(g940_n),
    .din1(ffc_207_n),
    .din2(g939_n)
  );


  FA
  g_g941_n
  (
    .dout(g941_n),
    .din1(g936_n),
    .din2(g940_n)
  );


  LA
  g_g942_p
  (
    .dout(g942_p),
    .din1(g931_n),
    .din2(g941_n)
  );


  FA
  g_g943_n
  (
    .dout(g943_n),
    .din1(g612_p_spl_1),
    .din2(g942_p)
  );


  LA
  g_g944_p
  (
    .dout(g944_p),
    .din1(g562_p_spl_10),
    .din2(g943_n)
  );


  LA
  g_g945_p
  (
    .dout(g945_p),
    .din1(g920_n),
    .din2(g944_p)
  );


  LA
  g_g946_p
  (
    .dout(g946_p),
    .din1(g735_p_spl_),
    .din2(g888_n_spl_)
  );


  LA
  g_g947_p
  (
    .dout(g947_p),
    .din1(g735_n_spl_),
    .din2(g888_p)
  );


  FA
  g_g948_n
  (
    .dout(g948_n),
    .din1(g946_p),
    .din2(g947_p)
  );


  LA
  g_g949_p
  (
    .dout(g949_p),
    .din1(ffc_130_p_spl_),
    .din2(ffc_163_p_spl_0)
  );


  FA
  g_g950_n
  (
    .dout(g950_n),
    .din1(g597_p_spl_0),
    .din2(g949_p)
  );


  LA
  g_g951_p
  (
    .dout(g951_p),
    .din1(ffc_147_n),
    .din2(ffc_155_p_spl_1)
  );


  FA
  g_g951_n
  (
    .dout(g951_n),
    .din1(ffc_147_p),
    .din2(ffc_155_n_spl_1)
  );


  LA
  g_g952_p
  (
    .dout(g952_p),
    .din1(ffc_148_n_spl_),
    .din2(ffc_171_p_spl_1)
  );


  FA
  g_g952_n
  (
    .dout(g952_n),
    .din1(ffc_148_p),
    .din2(ffc_171_n_spl_)
  );


  LA
  g_g953_p
  (
    .dout(g953_p),
    .din1(ffc_189_n),
    .din2(g952_n)
  );


  FA
  g_g953_n
  (
    .dout(g953_n),
    .din1(ffc_189_p),
    .din2(g952_p)
  );


  LA
  g_g954_p
  (
    .dout(g954_p),
    .din1(g951_p),
    .din2(g953_p)
  );


  LA
  g_g955_p
  (
    .dout(g955_p),
    .din1(g951_n),
    .din2(g953_n)
  );


  FA
  g_g956_n
  (
    .dout(g956_n),
    .din1(g954_p),
    .din2(g955_p)
  );


  LA
  g_g957_p
  (
    .dout(g957_p),
    .din1(g553_p_spl_0),
    .din2(g730_n_spl_1)
  );


  FA
  g_g957_n
  (
    .dout(g957_n),
    .din1(g553_n_spl_),
    .din2(g730_p_spl_1)
  );


  LA
  g_g958_p
  (
    .dout(g958_p),
    .din1(ffc_116_p),
    .din2(ffc_122_n_spl_)
  );


  FA
  g_g958_n
  (
    .dout(g958_n),
    .din1(ffc_116_n),
    .din2(ffc_122_p_spl_)
  );


  LA
  g_g959_p
  (
    .dout(g959_p),
    .din1(g730_n_spl_1),
    .din2(g731_n_spl_)
  );


  FA
  g_g959_n
  (
    .dout(g959_n),
    .din1(g730_p_spl_1),
    .din2(g731_p_spl_)
  );


  LA
  g_g960_p
  (
    .dout(g960_p),
    .din1(g958_n),
    .din2(g959_n)
  );


  FA
  g_g960_n
  (
    .dout(g960_n),
    .din1(g958_p),
    .din2(g959_p)
  );


  LA
  g_g961_p
  (
    .dout(g961_p),
    .din1(g873_n_spl_0),
    .din2(g960_p_spl_)
  );


  FA
  g_g961_n
  (
    .dout(g961_n),
    .din1(g873_p_spl_),
    .din2(g960_n_spl_)
  );


  LA
  g_g962_p
  (
    .dout(g962_p),
    .din1(g873_p_spl_),
    .din2(g960_n_spl_)
  );


  FA
  g_g962_n
  (
    .dout(g962_n),
    .din1(g873_n_spl_),
    .din2(g960_p_spl_)
  );


  LA
  g_g963_p
  (
    .dout(g963_p),
    .din1(g961_n),
    .din2(g962_n)
  );


  FA
  g_g963_n
  (
    .dout(g963_n),
    .din1(g961_p),
    .din2(g962_p)
  );


  LA
  g_g964_p
  (
    .dout(g964_p),
    .din1(g957_n),
    .din2(g963_n)
  );


  LA
  g_g965_p
  (
    .dout(g965_p),
    .din1(g957_p),
    .din2(g963_p)
  );


  FA
  g_g966_n
  (
    .dout(g966_n),
    .din1(g964_p),
    .din2(g965_p)
  );


  FA
  g_g967_n
  (
    .dout(g967_n),
    .din1(g621_n_spl_0),
    .din2(g645_n_spl_0)
  );


  LA
  g_g968_p
  (
    .dout(g968_p),
    .din1(g621_n_spl_0),
    .din2(g645_n_spl_0)
  );


  LA
  g_g969_p
  (
    .dout(g969_p),
    .din1(ffc_198_p),
    .din2(ffc_328_p_spl_011)
  );


  FA
  g_g969_n
  (
    .dout(g969_n),
    .din1(ffc_198_n),
    .din2(ffc_328_n_spl_01)
  );


  LA
  g_g970_p
  (
    .dout(g970_p),
    .din1(ffc_299_n),
    .din2(g969_n)
  );


  LA
  g_g971_p
  (
    .dout(g971_p),
    .din1(ffc_299_p),
    .din2(g969_p)
  );


  FA
  g_g972_n
  (
    .dout(g972_n),
    .din1(g970_p),
    .din2(g971_p)
  );


  LA
  g_g973_p
  (
    .dout(g973_p),
    .din1(ffc_238_p),
    .din2(ffc_328_p_spl_011)
  );


  FA
  g_g973_n
  (
    .dout(g973_n),
    .din1(ffc_238_n),
    .din2(ffc_328_n_spl_10)
  );


  LA
  g_g974_p
  (
    .dout(g974_p),
    .din1(ffc_329_n_spl_),
    .din2(g973_n)
  );


  LA
  g_g975_p
  (
    .dout(g975_p),
    .din1(ffc_329_p_spl_),
    .din2(g973_p)
  );


  FA
  g_g976_n
  (
    .dout(g976_n),
    .din1(g974_p),
    .din2(g975_p)
  );


  LA
  g_g977_p
  (
    .dout(g977_p),
    .din1(ffc_246_n_spl_1),
    .din2(ffc_339_n_spl_1)
  );


  FA
  g_g977_n
  (
    .dout(g977_n),
    .din1(ffc_246_p_spl_1),
    .din2(ffc_339_p_spl_)
  );


  LA
  g_g978_p
  (
    .dout(g978_p),
    .din1(ffc_251_p_spl_),
    .din2(ffc_314_p_spl_0)
  );


  FA
  g_g978_n
  (
    .dout(g978_n),
    .din1(ffc_251_n),
    .din2(ffc_314_n_spl_)
  );


  LA
  g_g979_p
  (
    .dout(g979_p),
    .din1(g977_n),
    .din2(g978_n)
  );


  FA
  g_g979_n
  (
    .dout(g979_n),
    .din1(g977_p),
    .din2(g978_p)
  );


  LA
  g_g980_p
  (
    .dout(g980_p),
    .din1(ffc_323_p_spl_01),
    .din2(g979_n)
  );


  FA
  g_g980_n
  (
    .dout(g980_n),
    .din1(ffc_323_n_spl_1),
    .din2(g979_p)
  );


  LA
  g_g981_p
  (
    .dout(g981_p),
    .din1(ffc_248_n_spl_0),
    .din2(ffc_315_n_spl_1)
  );


  FA
  g_g981_n
  (
    .dout(g981_n),
    .din1(ffc_248_p_spl_0),
    .din2(ffc_315_p_spl_01)
  );


  LA
  g_g982_p
  (
    .dout(g982_p),
    .din1(ffc_248_p_spl_1),
    .din2(g692_n_spl_)
  );


  FA
  g_g982_n
  (
    .dout(g982_n),
    .din1(ffc_248_n_spl_),
    .din2(g692_p_spl_0)
  );


  LA
  g_g983_p
  (
    .dout(g983_p),
    .din1(g668_n_spl_1),
    .din2(g982_p)
  );


  FA
  g_g983_n
  (
    .dout(g983_n),
    .din1(g668_p_spl_1),
    .din2(g982_n)
  );


  LA
  g_g984_p
  (
    .dout(g984_p),
    .din1(g981_n),
    .din2(g983_n)
  );


  FA
  g_g984_n
  (
    .dout(g984_n),
    .din1(g981_p),
    .din2(g983_p)
  );


  LA
  g_g985_p
  (
    .dout(g985_p),
    .din1(g980_n),
    .din2(g984_n)
  );


  FA
  g_g985_n
  (
    .dout(g985_n),
    .din1(g980_p),
    .din2(g984_p)
  );


  LA
  g_g986_p
  (
    .dout(g986_p),
    .din1(ffc_324_p_spl_0),
    .din2(ffc_326_p_spl_)
  );


  FA
  g_g986_n
  (
    .dout(g986_n),
    .din1(ffc_324_n_spl_0),
    .din2(ffc_326_n)
  );


  LA
  g_g987_p
  (
    .dout(g987_p),
    .din1(ffc_347_n),
    .din2(ffc_354_n)
  );


  FA
  g_g987_n
  (
    .dout(g987_n),
    .din1(ffc_347_p),
    .din2(ffc_354_p)
  );


  LA
  g_g988_p
  (
    .dout(g988_p),
    .din1(g986_n),
    .din2(g987_p)
  );


  FA
  g_g988_n
  (
    .dout(g988_n),
    .din1(g986_p),
    .din2(g987_n)
  );


  LA
  g_g989_p
  (
    .dout(g989_p),
    .din1(ffc_348_n_spl_01),
    .din2(g988_n)
  );


  FA
  g_g989_n
  (
    .dout(g989_n),
    .din1(ffc_348_p_spl_01),
    .din2(g988_p)
  );


  LA
  g_g990_p
  (
    .dout(g990_p),
    .din1(g708_n_spl_0),
    .din2(g989_n)
  );


  FA
  g_g990_n
  (
    .dout(g990_n),
    .din1(g708_p_spl_0),
    .din2(g989_p)
  );


  FA
  g_g991_n
  (
    .dout(g991_n),
    .din1(g658_p_spl_1),
    .din2(g990_n_spl_)
  );


  FA
  g_g992_n
  (
    .dout(g992_n),
    .din1(g701_p),
    .din2(g991_n)
  );


  LA
  g_g993_p
  (
    .dout(g993_p),
    .din1(g659_n_spl_00),
    .din2(g705_p_spl_)
  );


  FA
  g_g994_n
  (
    .dout(g994_n),
    .din1(g676_n_spl_),
    .din2(g993_p)
  );


  LA
  g_g995_p
  (
    .dout(g995_p),
    .din1(g707_n_spl_),
    .din2(g994_n)
  );


  LA
  g_g996_p
  (
    .dout(g996_p),
    .din1(g659_n_spl_00),
    .din2(g711_p_spl_)
  );


  FA
  g_g997_n
  (
    .dout(g997_n),
    .din1(g684_n_spl_),
    .din2(g996_p)
  );


  LA
  g_g998_p
  (
    .dout(g998_p),
    .din1(g713_n_spl_),
    .din2(g997_n)
  );


  FA
  g_g999_n
  (
    .dout(g999_n),
    .din1(ffc_124_p_spl_1),
    .din2(ffc_126_p_spl_)
  );


  LA
  g_g1000_p
  (
    .dout(g1000_p),
    .din1(ffc_129_p_spl_),
    .din2(ffc_162_p_spl_)
  );


  LA
  g_g1001_p
  (
    .dout(g1001_p),
    .din1(ffc_37_n),
    .din2(ffc_132_p_spl_)
  );


  LA
  g_g1002_p
  (
    .dout(g1002_p),
    .din1(ffc_132_n_spl_),
    .din2(g581_n_spl_00)
  );


  LA
  g_g1003_p
  (
    .dout(g1003_p),
    .din1(ffc_145_p_spl_),
    .din2(g597_n_spl_0)
  );


  LA
  g_g1004_p
  (
    .dout(g1004_p),
    .din1(ffc_15_p_spl_0),
    .din2(g583_n_spl_00)
  );


  FA
  g_g1005_n
  (
    .dout(g1005_n),
    .din1(ffc_142_n),
    .din2(g1004_p)
  );


  LA
  g_g1006_p
  (
    .dout(g1006_p),
    .din1(ffc_150_p_spl_0),
    .din2(ffc_196_n)
  );


  LA
  g_g1007_p
  (
    .dout(g1007_p),
    .din1(ffc_151_p_spl_0),
    .din2(ffc_197_n)
  );


  LA
  g_g1008_p
  (
    .dout(g1008_p),
    .din1(ffc_21_n),
    .din2(ffc_163_p_spl_0)
  );


  FA
  g_g1009_n
  (
    .dout(g1009_n),
    .din1(ffc_162_n_spl_),
    .din2(ffc_163_n)
  );


  LA
  g_g1010_p
  (
    .dout(g1010_p),
    .din1(ffc_180_p),
    .din2(g1009_n)
  );


  LA
  g_g1011_p
  (
    .dout(g1011_p),
    .din1(ffc_192_p),
    .din2(ffc_328_p_spl_10)
  );


  LA
  g_g1012_p
  (
    .dout(g1012_p),
    .din1(ffc_239_p_spl_),
    .din2(ffc_328_n_spl_10)
  );


  LA
  g_g1013_p
  (
    .dout(g1013_p),
    .din1(ffc_319_p_spl_),
    .din2(ffc_328_n_spl_11)
  );


  FA
  g_g1013_n
  (
    .dout(g1013_n),
    .din1(ffc_319_n_spl_0),
    .din2(ffc_328_p_spl_10)
  );


  FA
  g_g1014_n
  (
    .dout(g1014_n),
    .din1(g890_n_spl_),
    .din2(g1013_p_spl_0)
  );


  LA
  g_g1015_p
  (
    .dout(g1015_p),
    .din1(g567_p_spl_0),
    .din2(g886_n_spl_0)
  );


  LA
  g_g1016_p
  (
    .dout(g1016_p),
    .din1(ffc_13_p_spl_),
    .din2(g581_n_spl_00)
  );


  FA
  g_g1017_n
  (
    .dout(g1017_n),
    .din1(ffc_48_n_spl_),
    .din2(g976_n_spl_)
  );


  LA
  g_g1018_p
  (
    .dout(g1018_p),
    .din1(ffc_39_p_spl_),
    .din2(g581_n_spl_01)
  );


  LA
  g_g1019_p
  (
    .dout(g1019_p),
    .din1(ffc_37_p_spl_),
    .din2(g583_n_spl_00)
  );


  FA
  g_g1020_n
  (
    .dout(g1020_n),
    .din1(ffc_291_n_spl_0),
    .din2(g877_p_spl_)
  );


  LA
  g_g1021_p
  (
    .dout(g1021_p),
    .din1(g883_n_spl_0),
    .din2(g1020_n_spl_)
  );


  FA
  g_g1022_n
  (
    .dout(g1022_n),
    .din1(g883_n_spl_1),
    .din2(g1020_n_spl_)
  );


  LA
  g_g1023_p
  (
    .dout(g1023_p),
    .din1(g592_n_spl_),
    .din2(g886_n_spl_0)
  );


  LA
  g_g1024_p
  (
    .dout(g1024_p),
    .din1(ffc_48_p_spl_),
    .din2(g590_p_spl_)
  );


  FA
  g_g1024_n
  (
    .dout(g1024_n),
    .din1(ffc_48_n_spl_),
    .din2(g590_n)
  );


  FA
  g_g1025_n
  (
    .dout(g1025_n),
    .din1(g577_n_spl_0),
    .din2(g1024_n)
  );


  LA
  g_g1026_p
  (
    .dout(g1026_p),
    .din1(ffc_320_p_spl_),
    .din2(ffc_328_n_spl_11)
  );


  FA
  g_g1026_n
  (
    .dout(g1026_n),
    .din1(ffc_320_n_spl_0),
    .din2(ffc_328_p_spl_11)
  );


  LA
  g_g1027_p
  (
    .dout(g1027_p),
    .din1(g577_p_spl_0),
    .din2(g1013_n)
  );


  FA
  g_g1027_n
  (
    .dout(g1027_n),
    .din1(g577_n_spl_),
    .din2(g1013_p_spl_0)
  );


  LA
  g_g1028_p
  (
    .dout(g1028_p),
    .din1(g1026_n),
    .din2(g1027_n)
  );


  FA
  g_g1028_n
  (
    .dout(g1028_n),
    .din1(g1026_p_spl_),
    .din2(g1027_p)
  );


  LA
  g_g1029_p
  (
    .dout(g1029_p),
    .din1(g656_p_spl_0),
    .din2(g1028_p)
  );


  LA
  g_g1030_p
  (
    .dout(g1030_p),
    .din1(g656_n_spl_),
    .din2(g1028_n)
  );


  FA
  g_g1031_n
  (
    .dout(g1031_n),
    .din1(g1029_p),
    .din2(g1030_p)
  );


  FA
  g_g1032_n
  (
    .dout(g1032_n),
    .din1(g1025_n_spl_0),
    .din2(g1031_n_spl_)
  );


  LA
  g_g1033_p
  (
    .dout(g1033_p),
    .din1(g1025_n_spl_0),
    .din2(g1031_n_spl_)
  );


  FA
  g_g1034_n
  (
    .dout(g1034_n),
    .din1(G1_p_spl_0),
    .din2(G2_n_spl_)
  );


  FA
  g_g1035_n
  (
    .dout(g1035_n),
    .din1(G1_p_spl_0),
    .din2(G6_p_spl_)
  );


  LA
  g_g1036_p
  (
    .dout(g1036_p),
    .din1(g662_n_spl_),
    .din2(g664_n_spl_)
  );


  LA
  g_g1037_p
  (
    .dout(g1037_p),
    .din1(g716_p_spl_),
    .din2(g1036_p)
  );


  LA
  g_g1038_p
  (
    .dout(g1038_p),
    .din1(ffc_196_p_spl_0),
    .din2(g599_n_spl_0)
  );


  LA
  g_g1039_p
  (
    .dout(g1039_p),
    .din1(g591_n_spl_),
    .din2(g597_n_spl_1)
  );


  FA
  g_g1040_n
  (
    .dout(g1040_n),
    .din1(g1038_p),
    .din2(g1039_p)
  );


  FA
  g_g1041_n
  (
    .dout(g1041_n),
    .din1(ffc_13_p_spl_),
    .din2(ffc_21_p_spl_0)
  );


  LA
  g_g1042_p
  (
    .dout(g1042_p),
    .din1(g598_n_spl_0),
    .din2(g1041_n)
  );


  FA
  g_g1043_n
  (
    .dout(g1043_n),
    .din1(ffc_127_p_spl_0),
    .din2(g1042_p)
  );


  FA
  g_g1044_n
  (
    .dout(g1044_n),
    .din1(g1040_n),
    .din2(g1043_n)
  );


  LA
  g_g1045_p
  (
    .dout(g1045_p),
    .din1(ffc_127_n),
    .din2(ffc_137_p_spl_)
  );


  LA
  g_g1046_p
  (
    .dout(g1046_p),
    .din1(g719_n_spl_),
    .din2(g1045_p)
  );


  LA
  g_g1047_p
  (
    .dout(g1047_p),
    .din1(ffc_131_n),
    .din2(g583_n_spl_01)
  );


  FA
  g_g1048_n
  (
    .dout(g1048_n),
    .din1(ffc_129_n_spl_),
    .din2(ffc_135_p_spl_0)
  );


  LA
  g_g1049_p
  (
    .dout(g1049_p),
    .din1(g598_n_spl_0),
    .din2(g1048_n)
  );


  FA
  g_g1050_n
  (
    .dout(g1050_n),
    .din1(g1047_p),
    .din2(g1049_p)
  );


  FA
  g_g1051_n
  (
    .dout(g1051_n),
    .din1(ffc_150_p_spl_1),
    .din2(ffc_151_p_spl_1)
  );


  FA
  g_g1052_n
  (
    .dout(g1052_n),
    .din1(ffc_150_n_spl_),
    .din2(ffc_151_n)
  );


  LA
  g_g1053_p
  (
    .dout(g1053_p),
    .din1(g1051_n),
    .din2(g1052_n)
  );


  LA
  g_g1054_p
  (
    .dout(g1054_p),
    .din1(g720_n_spl_),
    .din2(g950_n_spl_)
  );


  FA
  g_g1055_n
  (
    .dout(g1055_n),
    .din1(ffc_11_p),
    .din2(ffc_19_p_spl_0)
  );


  LA
  g_g1056_p
  (
    .dout(g1056_p),
    .din1(g598_n_spl_1),
    .din2(g1055_n)
  );


  LA
  g_g1057_p
  (
    .dout(g1057_p),
    .din1(ffc_196_p_spl_0),
    .din2(g595_n_spl_0)
  );


  FA
  g_g1058_n
  (
    .dout(g1058_n),
    .din1(g1056_p),
    .din2(g1057_p)
  );


  LA
  g_g1059_p
  (
    .dout(g1059_p),
    .din1(ffc_197_p_spl_0),
    .din2(g595_n_spl_0)
  );


  LA
  g_g1060_p
  (
    .dout(g1060_p),
    .din1(ffc_15_p_spl_0),
    .din2(g581_n_spl_01)
  );


  LA
  g_g1061_p
  (
    .dout(g1061_p),
    .din1(ffc_17_p_spl_0),
    .din2(g583_n_spl_01)
  );


  FA
  g_g1062_n
  (
    .dout(g1062_n),
    .din1(g1060_p),
    .din2(g1061_p)
  );


  FA
  g_g1063_n
  (
    .dout(g1063_n),
    .din1(g1059_p),
    .din2(g1062_n)
  );


  LA
  g_g1064_p
  (
    .dout(g1064_p),
    .din1(g656_p_spl_0),
    .din2(g1026_p_spl_)
  );


  LA
  g_g1065_p
  (
    .dout(g1065_p),
    .din1(ffc_291_n_spl_),
    .din2(g651_p_spl_)
  );


  FA
  g_g1066_n
  (
    .dout(g1066_n),
    .din1(g1064_p),
    .din2(g1065_p)
  );


  LA
  g_g1067_p
  (
    .dout(g1067_p),
    .din1(g875_n_spl_),
    .din2(g972_n_spl_)
  );


  FA
  g_g1068_n
  (
    .dout(g1068_n),
    .din1(ffc_319_n_spl_),
    .din2(g885_n_spl_)
  );


  FA
  g_g1069_n
  (
    .dout(g1069_n),
    .din1(ffc_320_n_spl_),
    .din2(g884_n_spl_)
  );


  FA
  g_g1070_n
  (
    .dout(g1070_n),
    .din1(g651_n_spl_),
    .din2(g883_n_spl_1)
  );


  LA
  g_g1071_p
  (
    .dout(g1071_p),
    .din1(g882_n),
    .din2(g1070_n)
  );


  LA
  g_g1072_p
  (
    .dout(g1072_p),
    .din1(g1069_n),
    .din2(g1071_p)
  );


  LA
  g_g1073_p
  (
    .dout(g1073_p),
    .din1(g1068_n),
    .din2(g1072_p)
  );


  FA
  g_g1074_n
  (
    .dout(g1074_n),
    .din1(ffc_24_n),
    .din2(g876_n_spl_)
  );


  LA
  g_g1075_p
  (
    .dout(g1075_p),
    .din1(ffc_333_n_spl_0),
    .din2(ffc_339_n_spl_1)
  );


  LA
  g_g1076_p
  (
    .dout(g1076_p),
    .din1(ffc_245_n_spl_1),
    .din2(ffc_313_p_spl_0)
  );


  FA
  g_g1077_n
  (
    .dout(g1077_n),
    .din1(g1075_p),
    .din2(g1076_p)
  );


  LA
  g_g1078_p
  (
    .dout(g1078_p),
    .din1(ffc_323_p_spl_10),
    .din2(g1077_n)
  );


  FA
  g_g1079_n
  (
    .dout(g1079_n),
    .din1(ffc_315_p_spl_10),
    .din2(ffc_358_p_spl_00)
  );


  FA
  g_g1080_n
  (
    .dout(g1080_n),
    .din1(ffc_358_n_spl_),
    .din2(g692_p_spl_)
  );


  FA
  g_g1081_n
  (
    .dout(g1081_n),
    .din1(ffc_201_p_spl_1),
    .din2(ffc_202_n_spl_)
  );


  LA
  g_g1082_p
  (
    .dout(g1082_p),
    .din1(ffc_353_n_spl_),
    .din2(g1081_n)
  );


  FA
  g_g1083_n
  (
    .dout(g1083_n),
    .din1(g1080_n),
    .din2(g1082_p_spl_0)
  );


  LA
  g_g1084_p
  (
    .dout(g1084_p),
    .din1(g1079_n),
    .din2(g1083_n)
  );


  FA
  g_g1085_n
  (
    .dout(g1085_n),
    .din1(g1078_p),
    .din2(g1084_p)
  );


  FA
  g_g1086_n
  (
    .dout(g1086_n),
    .din1(g666_p_spl_),
    .din2(g1013_p_spl_)
  );


  FA
  g_g1087_n
  (
    .dout(g1087_n),
    .din1(g577_p_spl_0),
    .din2(g1024_p)
  );


  LA
  g_g1088_p
  (
    .dout(g1088_p),
    .din1(g1025_n_spl_),
    .din2(g1087_n)
  );


  FA
  g_g1089_n
  (
    .dout(g1089_n),
    .din1(g1086_n_spl_),
    .din2(g1088_p_spl_)
  );


  LA
  g_g1090_p
  (
    .dout(g1090_p),
    .din1(g1086_n_spl_),
    .din2(g1088_p_spl_)
  );


  LA
  g_g1091_p
  (
    .dout(g1091_p),
    .din1(ffc_357_n_spl_1),
    .din2(g693_n_spl_)
  );


  LA
  g_g1092_p
  (
    .dout(g1092_p),
    .din1(ffc_332_p_spl_0),
    .din2(ffc_340_n_spl_0)
  );


  LA
  g_g1093_p
  (
    .dout(g1093_p),
    .din1(ffc_314_p_spl_),
    .din2(ffc_358_p_spl_0)
  );


  FA
  g_g1094_n
  (
    .dout(g1094_n),
    .din1(g1092_p),
    .din2(g1093_p)
  );


  LA
  g_g1095_p
  (
    .dout(g1095_p),
    .din1(ffc_323_p_spl_10),
    .din2(g1094_n)
  );


  LA
  g_g1096_p
  (
    .dout(g1096_p),
    .din1(ffc_357_p_spl_1),
    .din2(g1082_p_spl_0)
  );


  FA
  g_g1097_n
  (
    .dout(g1097_n),
    .din1(g1095_p),
    .din2(g1096_p)
  );


  FA
  g_g1098_n
  (
    .dout(g1098_n),
    .din1(g1091_p),
    .din2(g1097_n)
  );


  LA
  g_g1099_p
  (
    .dout(g1099_p),
    .din1(ffc_21_p_spl_0),
    .din2(g599_n_spl_)
  );


  LA
  g_g1100_p
  (
    .dout(g1100_p),
    .din1(g597_n_spl_1),
    .din2(g665_n_spl_)
  );


  FA
  g_g1101_n
  (
    .dout(g1101_n),
    .din1(g1099_p),
    .din2(g1100_p)
  );


  LA
  g_g1102_p
  (
    .dout(g1102_p),
    .din1(ffc_324_p_spl_),
    .din2(ffc_352_p_spl_)
  );


  FA
  g_g1102_n
  (
    .dout(g1102_n),
    .din1(ffc_324_n_spl_),
    .din2(ffc_352_n)
  );


  LA
  g_g1103_p
  (
    .dout(g1103_p),
    .din1(ffc_343_p),
    .din2(ffc_344_n)
  );


  FA
  g_g1103_n
  (
    .dout(g1103_n),
    .din1(ffc_343_n),
    .din2(ffc_344_p)
  );


  LA
  g_g1104_p
  (
    .dout(g1104_p),
    .din1(ffc_302_p_spl_),
    .din2(ffc_304_n_spl_0)
  );


  FA
  g_g1104_n
  (
    .dout(g1104_n),
    .din1(ffc_302_n),
    .din2(ffc_304_p_spl_0)
  );


  LA
  g_g1105_p
  (
    .dout(g1105_p),
    .din1(g1103_n),
    .din2(g1104_n)
  );


  FA
  g_g1105_n
  (
    .dout(g1105_n),
    .din1(g1103_p),
    .din2(g1104_p)
  );


  LA
  g_g1106_p
  (
    .dout(g1106_p),
    .din1(g1102_n),
    .din2(g1105_p)
  );


  FA
  g_g1106_n
  (
    .dout(g1106_n),
    .din1(g1102_p),
    .din2(g1105_n)
  );


  LA
  g_g1107_p
  (
    .dout(g1107_p),
    .din1(ffc_348_n_spl_10),
    .din2(g1106_n)
  );


  FA
  g_g1107_n
  (
    .dout(g1107_n),
    .din1(ffc_348_p_spl_10),
    .din2(g1106_p)
  );


  LA
  g_g1108_p
  (
    .dout(g1108_p),
    .din1(g708_n_spl_),
    .din2(g1107_n)
  );


  FA
  g_g1108_n
  (
    .dout(g1108_n),
    .din1(g708_p_spl_),
    .din2(g1107_p)
  );


  FA
  g_g1109_n
  (
    .dout(g1109_n),
    .din1(g658_p_spl_1),
    .din2(g1108_n_spl_)
  );


  FA
  g_g1110_n
  (
    .dout(g1110_n),
    .din1(g985_p),
    .din2(g1109_n)
  );


  LA
  g_g1111_p
  (
    .dout(g1111_p),
    .din1(ffc_130_n),
    .din2(g598_n_spl_1)
  );


  FA
  g_g1112_n
  (
    .dout(g1112_n),
    .din1(g663_p_spl_),
    .din2(g1111_p)
  );


  LA
  g_g1113_p
  (
    .dout(g1113_p),
    .din1(ffc_135_p_spl_0),
    .din2(g581_n_spl_1)
  );


  LA
  g_g1114_p
  (
    .dout(g1114_p),
    .din1(ffc_132_n_spl_),
    .din2(g583_n_spl_1)
  );


  FA
  g_g1115_n
  (
    .dout(g1115_n),
    .din1(g1113_p),
    .din2(g1114_p)
  );


  FA
  g_g1116_n
  (
    .dout(g1116_n),
    .din1(g660_p_spl_),
    .din2(g1115_n)
  );


  FA
  g_g1117_n
  (
    .dout(g1117_n),
    .din1(g1112_n),
    .din2(g1116_n)
  );


  LA
  g_g1118_p
  (
    .dout(g1118_p),
    .din1(g659_n_spl_01),
    .din2(g990_p_spl_)
  );


  FA
  g_g1119_n
  (
    .dout(g1119_n),
    .din1(g701_n_spl_),
    .din2(g1118_p)
  );


  LA
  g_g1120_p
  (
    .dout(g1120_p),
    .din1(g992_n_spl_),
    .din2(g1119_n)
  );


  LA
  g_g1121_p
  (
    .dout(g1121_p),
    .din1(g995_p_spl_),
    .din2(g998_p_spl_)
  );


  FA
  g_g1122_n
  (
    .dout(g1122_n),
    .din1(G4_p_spl_000),
    .din2(G49_p)
  );


  FA
  g_g1123_n
  (
    .dout(g1123_n),
    .din1(G11_p_spl_),
    .din2(G12_p_spl_0)
  );


  FA
  g_g1124_n
  (
    .dout(g1124_n),
    .din1(G12_p_spl_0),
    .din2(G13_p_spl_0)
  );


  LA
  g_g1125_p
  (
    .dout(g1125_p),
    .din1(ffc_22_p_spl_),
    .din2(ffc_340_n_spl_1)
  );


  LA
  g_g1126_p
  (
    .dout(g1126_p),
    .din1(ffc_313_p_spl_0),
    .din2(ffc_333_n_spl_1)
  );


  LA
  g_g1127_p
  (
    .dout(g1127_p),
    .din1(ffc_202_p_spl_0),
    .din2(g667_n_spl_)
  );


  FA
  g_g1128_n
  (
    .dout(g1128_n),
    .din1(g1126_p),
    .din2(g1127_p)
  );


  FA
  g_g1129_n
  (
    .dout(g1129_n),
    .din1(g1125_p),
    .din2(g1128_n)
  );


  LA
  g_g1130_p
  (
    .dout(g1130_p),
    .din1(ffc_323_p_spl_11),
    .din2(g1129_n)
  );


  LA
  g_g1131_p
  (
    .dout(g1131_p),
    .din1(ffc_23_p_spl_),
    .din2(ffc_340_n_spl_1)
  );


  LA
  g_g1132_p
  (
    .dout(g1132_p),
    .din1(ffc_313_p_spl_),
    .din2(ffc_357_n_spl_1)
  );


  LA
  g_g1133_p
  (
    .dout(g1133_p),
    .din1(ffc_202_p_spl_1),
    .din2(g686_p_spl_)
  );


  FA
  g_g1134_n
  (
    .dout(g1134_n),
    .din1(g1132_p),
    .din2(g1133_p)
  );


  FA
  g_g1135_n
  (
    .dout(g1135_n),
    .din1(g1131_p),
    .din2(g1134_n)
  );


  LA
  g_g1136_p
  (
    .dout(g1136_p),
    .din1(ffc_323_p_spl_11),
    .din2(g1135_n)
  );


  LA
  g_g1137_p
  (
    .dout(g1137_p),
    .din1(ffc_351_p_spl_0),
    .din2(g690_n_spl_0)
  );


  FA
  g_g1138_n
  (
    .dout(g1138_n),
    .din1(ffc_243_p_spl_00),
    .din2(ffc_358_p_spl_1)
  );


  FA
  g_g1139_n
  (
    .dout(g1139_n),
    .din1(ffc_27_p_spl_),
    .din2(ffc_243_n_spl_0)
  );


  LA
  g_g1140_p
  (
    .dout(g1140_p),
    .din1(g1138_n),
    .din2(g1139_n)
  );


  LA
  g_g1141_p
  (
    .dout(g1141_p),
    .din1(ffc_26_p),
    .din2(ffc_304_n_spl_0)
  );


  FA
  g_g1142_n
  (
    .dout(g1142_n),
    .din1(g1140_p),
    .din2(g1141_p)
  );


  FA
  g_g1143_n
  (
    .dout(g1143_n),
    .din1(g1137_p),
    .din2(g1142_n)
  );


  LA
  g_g1144_p
  (
    .dout(g1144_p),
    .din1(ffc_348_n_spl_10),
    .din2(g1143_n)
  );


  FA
  g_g1145_n
  (
    .dout(g1145_n),
    .din1(g990_p_spl_),
    .din2(g1108_p_spl_)
  );


  FA
  g_g1146_n
  (
    .dout(g1146_n),
    .din1(g705_p_spl_),
    .din2(g711_p_spl_)
  );


  FA
  g_g1147_n
  (
    .dout(g1147_n),
    .din1(g1145_n),
    .din2(g1146_n)
  );


  LA
  g_g1148_p
  (
    .dout(g1148_p),
    .din1(ffc_335_p_spl_0),
    .din2(g1147_n)
  );


  FA
  g_g1149_n
  (
    .dout(g1149_n),
    .din1(g990_n_spl_),
    .din2(g1108_n_spl_)
  );


  FA
  g_g1150_n
  (
    .dout(g1150_n),
    .din1(g705_n_spl_),
    .din2(g711_n_spl_)
  );


  FA
  g_g1151_n
  (
    .dout(g1151_n),
    .din1(g1149_n),
    .din2(g1150_n)
  );


  LA
  g_g1152_p
  (
    .dout(g1152_p),
    .din1(ffc_335_n_spl_),
    .din2(g1151_n)
  );


  LA
  g_g1153_p
  (
    .dout(g1153_p),
    .din1(ffc_359_p_spl_),
    .din2(g690_n_spl_)
  );


  FA
  g_g1154_n
  (
    .dout(g1154_n),
    .din1(ffc_243_p_spl_00),
    .din2(ffc_245_p_spl_1)
  );


  FA
  g_g1155_n
  (
    .dout(g1155_n),
    .din1(ffc_243_n_spl_0),
    .din2(ffc_351_p_spl_0)
  );


  LA
  g_g1156_p
  (
    .dout(g1156_p),
    .din1(g1154_n),
    .din2(g1155_n)
  );


  LA
  g_g1157_p
  (
    .dout(g1157_p),
    .din1(ffc_27_p_spl_),
    .din2(ffc_304_n_spl_)
  );


  FA
  g_g1158_n
  (
    .dout(g1158_n),
    .din1(g1156_p),
    .din2(g1157_p)
  );


  FA
  g_g1159_n
  (
    .dout(g1159_n),
    .din1(g1153_p),
    .din2(g1158_n)
  );


  LA
  g_g1160_p
  (
    .dout(g1160_p),
    .din1(ffc_348_n_spl_1),
    .din2(g1159_n)
  );


  FA
  g_g1161_n
  (
    .dout(g1161_n),
    .din1(g691_p_spl_),
    .din2(g1160_p)
  );


  FA
  g_g1162_n
  (
    .dout(g1162_n),
    .din1(G3_p_spl_00),
    .din2(G4_n_spl_00)
  );


  FA
  g_g1163_n
  (
    .dout(g1163_n),
    .din1(G3_n_spl_),
    .din2(g1034_n_spl_)
  );


  LA
  g_g1164_p
  (
    .dout(g1164_p),
    .din1(G4_p_spl_000),
    .din2(G5_p_spl_0)
  );


  FA
  g_g1165_n
  (
    .dout(g1165_n),
    .din1(ffc_332_n),
    .din2(g1082_p_spl_1)
  );


  FA
  g_g1166_n
  (
    .dout(g1166_n),
    .din1(ffc_315_p_spl_10),
    .din2(ffc_332_p_spl_1)
  );


  LA
  g_g1167_p
  (
    .dout(g1167_p),
    .din1(g1165_n),
    .din2(g1166_n)
  );


  FA
  g_g1168_n
  (
    .dout(g1168_n),
    .din1(ffc_333_n_spl_1),
    .din2(g1082_p_spl_1)
  );


  FA
  g_g1169_n
  (
    .dout(g1169_n),
    .din1(ffc_315_p_spl_1),
    .din2(ffc_333_p_spl_1)
  );


  LA
  g_g1170_p
  (
    .dout(g1170_p),
    .din1(g1168_n),
    .din2(g1169_n)
  );


  FA
  g_g1171_n
  (
    .dout(g1171_n),
    .din1(ffc_249_n),
    .din2(g690_p_spl_0)
  );


  LA
  g_g1172_p
  (
    .dout(g1172_p),
    .din1(ffc_243_n_spl_1),
    .din2(ffc_247_n_spl_)
  );


  LA
  g_g1173_p
  (
    .dout(g1173_p),
    .din1(ffc_243_p_spl_0),
    .din2(ffc_325_n_spl_)
  );


  FA
  g_g1174_n
  (
    .dout(g1174_n),
    .din1(g1172_p),
    .din2(g1173_p)
  );


  FA
  g_g1175_n
  (
    .dout(g1175_n),
    .din1(ffc_304_p_spl_0),
    .din2(ffc_359_n_spl_)
  );


  LA
  g_g1176_p
  (
    .dout(g1176_p),
    .din1(g1174_n),
    .din2(g1175_n)
  );


  LA
  g_g1177_p
  (
    .dout(g1177_p),
    .din1(g1171_n),
    .din2(g1176_p)
  );


  FA
  g_g1178_n
  (
    .dout(g1178_n),
    .din1(ffc_348_p_spl_10),
    .din2(g1177_p)
  );


  LA
  g_g1179_p
  (
    .dout(g1179_p),
    .din1(g691_n_spl_),
    .din2(g1178_n)
  );


  LA
  g_g1180_p
  (
    .dout(g1180_p),
    .din1(g658_n_spl_0),
    .din2(g1179_p_spl_)
  );


  LA
  g_g1181_p
  (
    .dout(g1181_p),
    .din1(g1085_n_spl_0),
    .din2(g1180_p)
  );


  FA
  g_g1182_n
  (
    .dout(g1182_n),
    .din1(ffc_325_n_spl_),
    .din2(g690_p_spl_)
  );


  LA
  g_g1183_p
  (
    .dout(g1183_p),
    .din1(ffc_243_n_spl_1),
    .din2(ffc_246_n_spl_1)
  );


  LA
  g_g1184_p
  (
    .dout(g1184_p),
    .din1(ffc_243_p_spl_1),
    .din2(ffc_359_n_spl_)
  );


  FA
  g_g1185_n
  (
    .dout(g1185_n),
    .din1(g1183_p),
    .din2(g1184_p)
  );


  FA
  g_g1186_n
  (
    .dout(g1186_n),
    .din1(ffc_304_p_spl_),
    .din2(ffc_351_n)
  );


  LA
  g_g1187_p
  (
    .dout(g1187_p),
    .din1(g1185_n),
    .din2(g1186_n)
  );


  LA
  g_g1188_p
  (
    .dout(g1188_p),
    .din1(g1182_n),
    .din2(g1187_p)
  );


  FA
  g_g1189_n
  (
    .dout(g1189_n),
    .din1(ffc_348_p_spl_1),
    .din2(g1188_p)
  );


  LA
  g_g1190_p
  (
    .dout(g1190_p),
    .din1(g691_n_spl_),
    .din2(g1189_n)
  );


  LA
  g_g1191_p
  (
    .dout(g1191_p),
    .din1(g658_n_spl_0),
    .din2(g1190_p_spl_)
  );


  LA
  g_g1192_p
  (
    .dout(g1192_p),
    .din1(g1098_n_spl_0),
    .din2(g1191_p)
  );


  LA
  g_g1193_p
  (
    .dout(g1193_p),
    .din1(g659_n_spl_01),
    .din2(g1179_p_spl_)
  );


  FA
  g_g1194_n
  (
    .dout(g1194_n),
    .din1(g1085_n_spl_0),
    .din2(g1193_p)
  );


  LA
  g_g1195_p
  (
    .dout(g1195_p),
    .din1(g659_n_spl_10),
    .din2(g1190_p_spl_)
  );


  FA
  g_g1196_n
  (
    .dout(g1196_n),
    .din1(g1098_n_spl_0),
    .din2(g1195_p)
  );


  FA
  g_g1197_n
  (
    .dout(g1197_n),
    .din1(G1_n_spl_0),
    .din2(G2_n_spl_)
  );


  FA
  g_g1198_n
  (
    .dout(g1198_n),
    .din1(G1_n_spl_0),
    .din2(G3_n_spl_)
  );


  FA
  g_g1199_n
  (
    .dout(g1199_n),
    .din1(G4_n_spl_00),
    .din2(g1198_n)
  );


  LA
  g_g1200_p
  (
    .dout(g1200_p),
    .din1(g1197_n_spl_),
    .din2(g1199_n)
  );


  FA
  g_g1201_n
  (
    .dout(g1201_n),
    .din1(G5_p_spl_0),
    .din2(g1035_n_spl_0)
  );


  FA
  g_g1202_n
  (
    .dout(g1202_n),
    .din1(ffc_50_n),
    .din2(g1074_n_spl_)
  );


  LA
  g_g1203_p
  (
    .dout(g1203_p),
    .din1(g659_n_spl_10),
    .din2(g1108_p_spl_)
  );


  FA
  g_g1204_n
  (
    .dout(g1204_n),
    .din1(g985_n_spl_),
    .din2(g1203_p)
  );


  LA
  g_g1205_p
  (
    .dout(g1205_p),
    .din1(g1110_n_spl_),
    .din2(g1204_n)
  );


  LA
  g_g1206_p
  (
    .dout(g1206_p),
    .din1(g1120_p_spl_),
    .din2(g1121_p_spl_)
  );


  FA
  g_g1207_n
  (
    .dout(g1207_n),
    .din1(G12_n),
    .din2(G13_n_spl_)
  );


  LA
  g_g1208_p
  (
    .dout(g1208_p),
    .din1(g1124_n_spl_),
    .din2(g1207_n)
  );


  LA
  g_g1209_p
  (
    .dout(g1209_p),
    .din1(G1_n_spl_),
    .din2(G4_p_spl_001)
  );


  FA
  g_g1210_n
  (
    .dout(g1210_n),
    .din1(G3_p_spl_00),
    .din2(G4_p_spl_001)
  );


  FA
  g_g1211_n
  (
    .dout(g1211_n),
    .din1(G13_p_spl_0),
    .din2(g1123_n_spl_)
  );


  LA
  g_g1212_p
  (
    .dout(g1212_p),
    .din1(G3_p_spl_0),
    .din2(g1211_n)
  );


  LA
  g_g1213_p
  (
    .dout(g1213_p),
    .din1(G3_p_spl_1),
    .din2(g1208_p_spl_)
  );


  FA
  g_g1214_n
  (
    .dout(g1214_n),
    .din1(G4_p_spl_01),
    .din2(G41_p_spl_)
  );


  LA
  g_g1215_p
  (
    .dout(g1215_p),
    .din1(G4_p_spl_01),
    .din2(G36_n)
  );


  FA
  g_g1216_n
  (
    .dout(g1216_n),
    .din1(G12_p_spl_1),
    .din2(g1162_n_spl_0)
  );


  FA
  g_g1217_n
  (
    .dout(g1217_n),
    .din1(G13_n_spl_),
    .din2(g1162_n_spl_0)
  );


  FA
  g_g1218_n
  (
    .dout(g1218_n),
    .din1(G34_n_spl_),
    .din2(g1122_n_spl_0)
  );


  FA
  g_g1219_n
  (
    .dout(g1219_n),
    .din1(g1164_p_spl_),
    .din2(g1197_n_spl_)
  );


  LA
  g_g1220_p
  (
    .dout(g1220_p),
    .din1(G35_p_spl_0),
    .din2(g1201_n_spl_)
  );


  FA
  g_g1221_n
  (
    .dout(g1221_n),
    .din1(G32_n),
    .din2(g1122_n_spl_0)
  );


  LA
  g_g1222_p
  (
    .dout(g1222_p),
    .din1(g1163_n_spl_),
    .din2(g1200_p_spl_)
  );


  FA
  g_g1223_n
  (
    .dout(g1223_n),
    .din1(G4_p_spl_10),
    .din2(G40_p_spl_)
  );


  FA
  g_g1224_n
  (
    .dout(g1224_n),
    .din1(G4_n_spl_0),
    .din2(G35_p_spl_0)
  );


  LA
  g_g1225_p
  (
    .dout(g1225_p),
    .din1(g1223_n),
    .din2(g1224_n)
  );


  LA
  g_g1226_p
  (
    .dout(g1226_p),
    .din1(G4_n_spl_1),
    .din2(G39_n)
  );


  LA
  g_g1227_p
  (
    .dout(g1227_p),
    .din1(G4_p_spl_10),
    .din2(G34_n_spl_)
  );


  FA
  g_g1228_n
  (
    .dout(g1228_n),
    .din1(g1226_p),
    .din2(g1227_p)
  );


  FA
  g_g1229_n
  (
    .dout(g1229_n),
    .din1(G33_n),
    .din2(g1122_n_spl_1)
  );


  LA
  g_g1230_p
  (
    .dout(g1230_p),
    .din1(g1228_n),
    .din2(g1229_n)
  );


  LA
  g_g1231_p
  (
    .dout(g1231_p),
    .din1(G4_p_spl_11),
    .din2(G33_p_spl_)
  );


  LA
  g_g1232_p
  (
    .dout(g1232_p),
    .din1(G4_n_spl_1),
    .din2(G14_p_spl_)
  );


  FA
  g_g1233_n
  (
    .dout(g1233_n),
    .din1(g1231_p),
    .din2(g1232_p)
  );


  LA
  g_g1234_p
  (
    .dout(g1234_p),
    .din1(G34_p_spl_),
    .din2(g1035_n_spl_0)
  );


  FA
  g_g1235_n
  (
    .dout(g1235_n),
    .din1(g1233_n),
    .din2(g1234_p)
  );


  buf

  (
    G3519_p,
    g412_p
  );


  buf

  (
    G3520_p,
    ffc_97_n
  );


  buf

  (
    G3521_p,
    g436_p
  );


  buf

  (
    G3522_p,
    g457_p
  );


  buf

  (
    G3523_p,
    g468_n
  );


  buf

  (
    G3524_p,
    g469_p
  );


  buf

  (
    G3525_p,
    g471_n
  );


  buf

  (
    G3526_p,
    ffc_100_p
  );


  buf

  (
    G3527_p,
    g474_n
  );


  buf

  (
    G3528_p,
    g477_n_spl_
  );


  buf

  (
    G3529_p,
    g480_n_spl_
  );


  buf

  (
    G3530_p,
    g502_n
  );


  buf

  (
    G3531_p,
    g505_n_spl_
  );


  buf

  (
    G3532_p,
    g508_n_spl_
  );


  buf

  (
    G3533_p,
    g511_n_spl_
  );


  buf

  (
    G3534_p,
    ffc_176_p
  );


  buf

  (
    G3535_p,
    ffc_177_p
  );


  buf

  (
    G3536_p,
    g514_n_spl_
  );


  buf

  (
    G3537_p,
    g520_n_spl_
  );


  buf

  (
    G3538_n,
    g524_p
  );


  buf

  (
    G3539_p,
    g544_n
  );


  buf

  (
    G3540_p,
    g550_p
  );


  DROC
  ffc_0_3
  (
    .doutp(ffc_0_p),
    .doutn(ffc_0_n),
    .din(ffc_67_p_spl_)
  );


  DROC
  ffc_1_3
  (
    .doutp(ffc_1_p),
    .doutn(ffc_1_n),
    .din(ffc_68_p_spl_)
  );


  DROC
  ffc_2_3
  (
    .doutp(ffc_2_p),
    .doutn(ffc_2_n),
    .din(ffc_103_p_spl_1)
  );


  DROC
  ffc_3_3
  (
    .doutp(ffc_3_p),
    .doutn(ffc_3_n),
    .din(ffc_104_p_spl_)
  );


  DROC
  ffc_4_3
  (
    .doutp(ffc_4_p),
    .doutn(ffc_4_n),
    .din(ffc_93_p)
  );


  DROC
  ffc_5_3
  (
    .doutp(ffc_5_p),
    .doutn(ffc_5_n),
    .din(ffc_94_p)
  );


  DROC
  ffc_6_3
  (
    .doutp(ffc_6_p),
    .doutn(ffc_6_n),
    .din(ffc_72_p_spl_)
  );


  DROC
  ffc_7_3
  (
    .doutp(ffc_7_p),
    .doutn(ffc_7_n),
    .din(ffc_73_p_spl_)
  );


  DROC
  ffc_8_3
  (
    .doutp(ffc_8_p),
    .doutn(ffc_8_n),
    .din(ffc_74_p_spl_)
  );


  DROC
  ffc_9_3
  (
    .doutp(ffc_9_p),
    .doutn(ffc_9_n),
    .din(ffc_75_p_spl_)
  );


  DROC
  ffc_10_0
  (
    .doutp(ffc_10_p),
    .doutn(ffc_10_n),
    .din(G15_p)
  );


  DROC
  ffc_11_1
  (
    .doutp(ffc_11_p),
    .doutn(ffc_11_n),
    .din(ffc_10_p)
  );


  DROC
  ffc_12_0
  (
    .doutp(ffc_12_p),
    .doutn(ffc_12_n),
    .din(G16_p)
  );


  DROC
  ffc_13_1
  (
    .doutp(ffc_13_p),
    .doutn(ffc_13_n),
    .din(ffc_12_p)
  );


  DROC
  ffc_14_0
  (
    .doutp(ffc_14_p),
    .doutn(ffc_14_n),
    .din(G17_p)
  );


  DROC
  ffc_15_1
  (
    .doutp(ffc_15_p),
    .doutn(ffc_15_n),
    .din(ffc_14_p)
  );


  DROC
  ffc_16_0
  (
    .doutp(ffc_16_p),
    .doutn(ffc_16_n),
    .din(G18_p)
  );


  DROC
  ffc_17_1
  (
    .doutp(ffc_17_p),
    .doutn(ffc_17_n),
    .din(ffc_16_p)
  );


  DROC
  ffc_18_0
  (
    .doutp(ffc_18_p),
    .doutn(ffc_18_n),
    .din(G19_p)
  );


  DROC
  ffc_19_1
  (
    .doutp(ffc_19_p),
    .doutn(ffc_19_n),
    .din(ffc_18_p)
  );


  DROC
  ffc_20_0
  (
    .doutp(ffc_20_p),
    .doutn(ffc_20_n),
    .din(G20_p)
  );


  DROC
  ffc_21_1
  (
    .doutp(ffc_21_p),
    .doutn(ffc_21_n),
    .din(ffc_20_p)
  );


  DROC
  ffc_22_0
  (
    .doutp(ffc_22_p),
    .doutn(ffc_22_n),
    .din(G21_p)
  );


  DROC
  ffc_23_0
  (
    .doutp(ffc_23_p),
    .doutn(ffc_23_n),
    .din(G22_p)
  );


  DROC
  ffc_24_0
  (
    .doutp(ffc_24_p),
    .doutn(ffc_24_n),
    .din(G27_p)
  );


  DROC
  ffc_25_3
  (
    .doutp(ffc_25_p),
    .doutn(ffc_25_n),
    .din(ffc_117_p)
  );


  DROC
  ffc_26_0
  (
    .doutp(ffc_26_p),
    .doutn(ffc_26_n),
    .din(G28_p)
  );


  DROC
  ffc_27_0
  (
    .doutp(ffc_27_p),
    .doutn(ffc_27_n),
    .din(G29_p)
  );


  DROC
  ffc_28_3
  (
    .doutp(ffc_28_p),
    .doutn(ffc_28_n),
    .din(ffc_98_p)
  );


  DROC
  ffc_29_3
  (
    .doutp(ffc_29_p),
    .doutn(ffc_29_n),
    .din(ffc_95_p)
  );


  DROC
  ffc_30_3
  (
    .doutp(ffc_30_p),
    .doutn(ffc_30_n),
    .din(ffc_87_p)
  );


  DROC
  ffc_31_3
  (
    .doutp(ffc_31_p),
    .doutn(ffc_31_n),
    .din(ffc_76_p)
  );


  DROC
  ffc_32_3
  (
    .doutp(ffc_32_p),
    .doutn(ffc_32_n),
    .din(ffc_77_p)
  );


  DROC
  ffc_33_3
  (
    .doutp(ffc_33_p),
    .doutn(ffc_33_n),
    .din(ffc_82_p)
  );


  DROC
  ffc_34_3
  (
    .doutp(ffc_34_p),
    .doutn(ffc_34_n),
    .din(ffc_88_p)
  );


  DROC
  ffc_35_3
  (
    .doutp(ffc_35_p),
    .doutn(ffc_35_n),
    .din(ffc_99_p)
  );


  DROC
  ffc_36_0
  (
    .doutp(ffc_36_p),
    .doutn(ffc_36_n),
    .din(G42_p)
  );


  DROC
  ffc_37_1
  (
    .doutp(ffc_37_p),
    .doutn(ffc_37_n),
    .din(ffc_36_p)
  );


  DROC
  ffc_38_0
  (
    .doutp(ffc_38_p),
    .doutn(ffc_38_n),
    .din(G43_p)
  );


  DROC
  ffc_39_1
  (
    .doutp(ffc_39_p),
    .doutn(ffc_39_n),
    .din(ffc_38_p)
  );


  DROC
  ffc_40_0
  (
    .doutp(ffc_40_p),
    .doutn(ffc_40_n),
    .din(G44_p)
  );


  DROC
  ffc_41_1
  (
    .doutp(ffc_41_p),
    .doutn(ffc_41_n),
    .din(ffc_40_p)
  );


  DROC
  ffc_42_0
  (
    .doutp(ffc_42_p),
    .doutn(ffc_42_n),
    .din(G45_p)
  );


  DROC
  ffc_43_1
  (
    .doutp(ffc_43_p),
    .doutn(ffc_43_n),
    .din(ffc_42_p)
  );


  DROC
  ffc_44_0
  (
    .doutp(ffc_44_p),
    .doutn(ffc_44_n),
    .din(G46_p)
  );


  DROC
  ffc_45_1
  (
    .doutp(ffc_45_p),
    .doutn(ffc_45_n),
    .din(ffc_44_p)
  );


  DROC
  ffc_46_2
  (
    .doutp(ffc_46_p),
    .doutn(ffc_46_n),
    .din(ffc_45_p)
  );


  DROC
  ffc_47_0
  (
    .doutp(ffc_47_p),
    .doutn(ffc_47_n),
    .din(G47_p)
  );


  DROC
  ffc_48_1
  (
    .doutp(ffc_48_p),
    .doutn(ffc_48_n),
    .din(ffc_47_p)
  );


  DROC
  ffc_49_3
  (
    .doutp(ffc_49_p),
    .doutn(ffc_49_n),
    .din(ffc_155_p_spl_1)
  );


  DROC
  ffc_50_0
  (
    .doutp(ffc_50_p),
    .doutn(ffc_50_n),
    .din(G48_p)
  );


  DROC
  ffc_51_3
  (
    .doutp(ffc_51_p),
    .doutn(ffc_51_n),
    .din(ffc_121_p)
  );


  DROC
  ffc_52_0
  (
    .doutp(ffc_52_p),
    .doutn(ffc_52_n),
    .din(G50_p)
  );


  DROC
  ffc_53_1
  (
    .doutp(ffc_53_p),
    .doutn(ffc_53_n),
    .din(ffc_52_p)
  );


  DROC
  ffc_54_2
  (
    .doutp(ffc_54_p),
    .doutn(ffc_54_n),
    .din(ffc_53_p)
  );


  DROC
  ffc_55_3
  (
    .doutp(ffc_55_p),
    .doutn(ffc_55_n),
    .din(ffc_54_p)
  );


  DROC
  ffc_56_3
  (
    .doutp(ffc_56_p),
    .doutn(ffc_56_n),
    .din(ffc_84_p_spl_)
  );


  DROC
  ffc_57_3
  (
    .doutp(ffc_57_p),
    .doutn(ffc_57_n),
    .din(ffc_85_p)
  );


  DROC
  ffc_58_3
  (
    .doutp(ffc_58_p),
    .doutn(ffc_58_n),
    .din(ffc_92_p)
  );


  DROC
  ffc_59_3
  (
    .doutp(ffc_59_p),
    .doutn(ffc_59_n),
    .din(ffc_109_p)
  );


  DROC
  ffc_60_3
  (
    .doutp(ffc_60_p),
    .doutn(ffc_60_n),
    .din(ffc_111_p)
  );


  DROC
  ffc_61_3
  (
    .doutp(ffc_61_p),
    .doutn(ffc_61_n),
    .din(ffc_114_p)
  );


  DROC
  ffc_62_3
  (
    .doutp(ffc_62_p),
    .doutn(ffc_62_n),
    .din(ffc_118_p_spl_)
  );


  DROC
  ffc_63_3
  (
    .doutp(ffc_63_p),
    .doutn(ffc_63_n),
    .din(ffc_125_p)
  );


  DROC
  ffc_64_3
  (
    .doutp(ffc_64_p),
    .doutn(ffc_64_n),
    .din(ffc_160_p)
  );


  DROC
  ffc_65_3
  (
    .doutp(ffc_65_p),
    .doutn(ffc_65_n),
    .din(ffc_161_p)
  );


  DROC
  ffc_66_3
  (
    .doutp(ffc_66_p),
    .doutn(ffc_66_n),
    .din(ffc_171_p_spl_1)
  );


  DROC
  ffc_67_2
  (
    .doutp(ffc_67_p),
    .doutn(ffc_67_n),
    .din(ffc_123_p)
  );


  DROC
  ffc_68_2
  (
    .doutp(ffc_68_p),
    .doutn(ffc_68_n),
    .din(ffc_124_p_spl_1)
  );


  DROC
  ffc_69_2
  (
    .doutp(ffc_69_p),
    .doutn(ffc_69_n),
    .din(ffc_126_p_spl_)
  );


  DROC
  ffc_70_2
  (
    .doutp(ffc_70_p),
    .doutn(ffc_70_n),
    .din(ffc_127_p_spl_)
  );


  DROC
  ffc_71_2
  (
    .doutp(ffc_71_p),
    .doutn(ffc_71_n),
    .din(ffc_128_p)
  );


  DROC
  ffc_72_2
  (
    .doutp(ffc_72_p),
    .doutn(ffc_72_n),
    .din(ffc_129_p_spl_)
  );


  DROC
  ffc_73_2
  (
    .doutp(ffc_73_p),
    .doutn(ffc_73_n),
    .din(ffc_130_p_spl_)
  );


  DROC
  ffc_74_2
  (
    .doutp(ffc_74_p),
    .doutn(ffc_74_n),
    .din(ffc_131_p_spl_)
  );


  DROC
  ffc_75_2
  (
    .doutp(ffc_75_p),
    .doutn(ffc_75_n),
    .din(ffc_132_p_spl_)
  );


  DROC
  ffc_76_2
  (
    .doutp(ffc_76_p),
    .doutn(ffc_76_n),
    .din(ffc_133_p)
  );


  DROC
  ffc_77_2
  (
    .doutp(ffc_77_p),
    .doutn(ffc_77_n),
    .din(ffc_134_p)
  );


  DROC
  ffc_78_2
  (
    .doutp(ffc_78_p),
    .doutn(ffc_78_n),
    .din(ffc_135_p_spl_)
  );


  DROC
  ffc_79_3
  (
    .doutp(ffc_79_p),
    .doutn(ffc_79_n),
    .din(ffc_223_p)
  );


  DROC
  ffc_80_3
  (
    .doutp(ffc_80_p),
    .doutn(ffc_80_n),
    .din(ffc_225_p)
  );


  DROC
  ffc_81_2
  (
    .doutp(ffc_81_p),
    .doutn(ffc_81_n),
    .din(ffc_137_p_spl_)
  );


  DROC
  ffc_82_2
  (
    .doutp(ffc_82_p),
    .doutn(ffc_82_n),
    .din(ffc_138_p)
  );


  DROC
  ffc_83_2
  (
    .doutp(ffc_83_p),
    .doutn(ffc_83_n),
    .din(ffc_139_p)
  );


  DROC
  ffc_84_2
  (
    .doutp(ffc_84_p),
    .doutn(ffc_84_n),
    .din(ffc_136_p)
  );


  DROC
  ffc_85_2
  (
    .doutp(ffc_85_p),
    .doutn(ffc_85_n),
    .din(ffc_140_p)
  );


  DROC
  ffc_86_2
  (
    .doutp(ffc_86_p),
    .doutn(ffc_86_n),
    .din(ffc_141_p)
  );


  DROC
  ffc_87_2
  (
    .doutp(ffc_87_p),
    .doutn(ffc_87_n),
    .din(ffc_143_p)
  );


  DROC
  ffc_88_2
  (
    .doutp(ffc_88_p),
    .doutn(ffc_88_n),
    .din(ffc_144_p)
  );


  DROC
  ffc_89_2
  (
    .doutp(ffc_89_p),
    .doutn(ffc_89_n),
    .din(ffc_145_p_spl_)
  );


  DROC
  ffc_90_3
  (
    .doutp(ffc_90_p),
    .doutn(ffc_90_n),
    .din(ffc_267_p_spl_)
  );


  DROC
  ffc_91_3
  (
    .doutp(ffc_91_p),
    .doutn(ffc_91_n),
    .din(ffc_290_p_spl_)
  );


  DROC
  ffc_92_2
  (
    .doutp(ffc_92_p),
    .doutn(ffc_92_n),
    .din(ffc_146_p)
  );


  DROC
  ffc_93_2
  (
    .doutp(ffc_93_p),
    .doutn(ffc_93_n),
    .din(ffc_150_p_spl_1)
  );


  DROC
  ffc_94_2
  (
    .doutp(ffc_94_p),
    .doutn(ffc_94_n),
    .din(ffc_151_p_spl_1)
  );


  DROC
  ffc_95_2
  (
    .doutp(ffc_95_p),
    .doutn(ffc_95_n),
    .din(ffc_152_p)
  );


  DROC
  ffc_96_3
  (
    .doutp(ffc_96_n),
    .doutn(ffc_96_p),
    .din(g551_n_spl_)
  );


  DROC
  ffc_97_3
  (
    .doutp(ffc_97_n),
    .doutn(ffc_97_p),
    .din(g552_n_spl_)
  );


  DROC
  ffc_98_2
  (
    .doutp(ffc_98_p),
    .doutn(ffc_98_n),
    .din(ffc_156_p)
  );


  DROC
  ffc_99_2
  (
    .doutp(ffc_99_p),
    .doutn(ffc_99_n),
    .din(ffc_157_p)
  );


  DROC
  ffc_100_3
  (
    .doutp(ffc_100_p),
    .doutn(ffc_100_n),
    .din(g553_p_spl_)
  );


  DROC
  ffc_101_3
  (
    .doutp(ffc_101_p),
    .doutn(ffc_101_n),
    .din(g554_n_spl_)
  );


  DROC
  ffc_102_3
  (
    .doutp(ffc_102_p),
    .doutn(ffc_102_n),
    .din(g555_p_spl_)
  );


  DROC
  ffc_103_2
  (
    .doutp(ffc_103_p),
    .doutn(ffc_103_n),
    .din(ffc_162_p_spl_)
  );


  DROC
  ffc_104_2
  (
    .doutp(ffc_104_p),
    .doutn(ffc_104_n),
    .din(ffc_163_p_spl_)
  );


  DROC
  ffc_105_2
  (
    .doutp(ffc_105_p),
    .doutn(ffc_105_n),
    .din(ffc_164_p)
  );


  DROC
  ffc_106_3
  (
    .doutp(ffc_106_p),
    .doutn(ffc_106_n),
    .din(g556_p_spl_)
  );


  DROC
  ffc_107_2
  (
    .doutp(ffc_107_p),
    .doutn(ffc_107_n),
    .din(ffc_178_p)
  );


  DROC
  ffc_108_3
  (
    .doutp(ffc_108_p),
    .doutn(ffc_108_n),
    .din(g559_n_spl_)
  );


  DROC
  ffc_109_2
  (
    .doutp(ffc_109_p),
    .doutn(ffc_109_n),
    .din(ffc_190_p)
  );


  DROC
  ffc_110_2
  (
    .doutp(ffc_110_p),
    .doutn(ffc_110_n),
    .din(ffc_191_p)
  );


  DROC
  ffc_111_2
  (
    .doutp(ffc_111_p),
    .doutn(ffc_111_n),
    .din(ffc_193_p)
  );


  DROC
  ffc_112_2
  (
    .doutp(ffc_112_p),
    .doutn(ffc_112_n),
    .din(ffc_196_p_spl_)
  );


  DROC
  ffc_113_2
  (
    .doutp(ffc_113_p),
    .doutn(ffc_113_n),
    .din(ffc_197_p_spl_)
  );


  DROC
  ffc_114_2
  (
    .doutp(ffc_114_p),
    .doutn(ffc_114_n),
    .din(ffc_194_p)
  );


  DROC
  ffc_115_3
  (
    .doutp(ffc_115_p),
    .doutn(ffc_115_n),
    .din(g562_p_spl_1)
  );


  DROC
  ffc_116_2
  (
    .doutp(ffc_116_p),
    .doutn(ffc_116_n),
    .din(ffc_200_p_spl_)
  );


  DROC
  ffc_117_2
  (
    .doutp(ffc_117_p),
    .doutn(ffc_117_n),
    .din(ffc_237_p)
  );


  DROC
  ffc_118_2
  (
    .doutp(ffc_118_p),
    .doutn(ffc_118_n),
    .din(ffc_222_p)
  );


  DROC
  ffc_119_2
  (
    .doutp(ffc_119_p),
    .doutn(ffc_119_n),
    .din(ffc_240_p_spl_)
  );


  DROC
  ffc_120_2
  (
    .doutp(ffc_120_p),
    .doutn(ffc_120_n),
    .din(ffc_241_p)
  );


  DROC
  ffc_121_2
  (
    .doutp(ffc_121_p),
    .doutn(ffc_121_n),
    .din(ffc_279_p)
  );


  DROC
  ffc_122_2
  (
    .doutp(ffc_122_p),
    .doutn(ffc_122_n),
    .din(ffc_328_p_spl_11)
  );


  DROC
  ffc_123_1
  (
    .doutp(ffc_123_p),
    .doutn(ffc_123_n),
    .din(ffc_201_p_spl_1)
  );


  DROC
  ffc_124_1
  (
    .doutp(ffc_124_p),
    .doutn(ffc_124_n),
    .din(ffc_202_p_spl_1)
  );


  DROC
  ffc_125_2
  (
    .doutp(ffc_125_p),
    .doutn(ffc_125_n),
    .din(g563_p_spl_)
  );


  DROC
  ffc_126_1
  (
    .doutp(ffc_126_p),
    .doutn(ffc_126_n),
    .din(ffc_242_p_spl_)
  );


  DROC
  ffc_127_1
  (
    .doutp(ffc_127_p),
    .doutn(ffc_127_n),
    .din(ffc_243_p_spl_1)
  );


  DROC
  ffc_128_1
  (
    .doutp(ffc_128_p),
    .doutn(ffc_128_n),
    .din(ffc_244_p_spl_)
  );


  DROC
  ffc_129_1
  (
    .doutp(ffc_129_p),
    .doutn(ffc_129_n),
    .din(ffc_245_p_spl_1)
  );


  DROC
  ffc_130_1
  (
    .doutp(ffc_130_p),
    .doutn(ffc_130_n),
    .din(ffc_246_p_spl_1)
  );


  DROC
  ffc_131_1
  (
    .doutp(ffc_131_p),
    .doutn(ffc_131_n),
    .din(ffc_247_p_spl_)
  );


  DROC
  ffc_132_1
  (
    .doutp(ffc_132_p),
    .doutn(ffc_132_n),
    .din(ffc_248_p_spl_1)
  );


  DROC
  ffc_133_1
  (
    .doutp(ffc_133_p),
    .doutn(ffc_133_n),
    .din(ffc_249_p)
  );


  DROC
  ffc_134_1
  (
    .doutp(ffc_134_p),
    .doutn(ffc_134_n),
    .din(ffc_250_p)
  );


  DROC
  ffc_135_1
  (
    .doutp(ffc_135_p),
    .doutn(ffc_135_n),
    .din(ffc_251_p_spl_)
  );


  DROC
  ffc_136_1
  (
    .doutp(ffc_136_p),
    .doutn(ffc_136_n),
    .din(ffc_277_p)
  );


  DROC
  ffc_137_1
  (
    .doutp(ffc_137_p),
    .doutn(ffc_137_n),
    .din(ffc_301_p_spl_)
  );


  DROC
  ffc_138_1
  (
    .doutp(ffc_138_p),
    .doutn(ffc_138_n),
    .din(ffc_302_p_spl_)
  );


  DROC
  ffc_139_1
  (
    .doutp(ffc_139_p),
    .doutn(ffc_139_n),
    .din(ffc_303_p)
  );


  DROC
  ffc_140_1
  (
    .doutp(ffc_140_p),
    .doutn(ffc_140_n),
    .din(ffc_305_p)
  );


  DROC
  ffc_141_1
  (
    .doutp(ffc_141_p),
    .doutn(ffc_141_n),
    .din(ffc_306_p)
  );


  DROC
  ffc_142_1
  (
    .doutp(ffc_142_p),
    .doutn(ffc_142_n),
    .din(ffc_316_p)
  );


  DROC
  ffc_143_1
  (
    .doutp(ffc_143_p),
    .doutn(ffc_143_n),
    .din(ffc_325_p)
  );


  DROC
  ffc_144_1
  (
    .doutp(ffc_144_p),
    .doutn(ffc_144_n),
    .din(ffc_326_p_spl_)
  );


  DROC
  ffc_145_1
  (
    .doutp(ffc_145_p),
    .doutn(ffc_145_n),
    .din(ffc_327_p)
  );


  DROC
  ffc_146_1
  (
    .doutp(ffc_146_p),
    .doutn(ffc_146_n),
    .din(ffc_331_p)
  );


  DROC
  ffc_147_2
  (
    .doutp(ffc_147_p),
    .doutn(ffc_147_n),
    .din(g567_p_spl_)
  );


  DROC
  ffc_148_2
  (
    .doutp(ffc_148_p),
    .doutn(ffc_148_n),
    .din(g572_p_spl_)
  );


  DROC
  ffc_149_2
  (
    .doutp(ffc_149_p),
    .doutn(ffc_149_n),
    .din(g577_p_spl_)
  );


  DROC
  ffc_150_1
  (
    .doutp(ffc_150_p),
    .doutn(ffc_150_n),
    .din(ffc_357_p_spl_1)
  );


  DROC
  ffc_151_1
  (
    .doutp(ffc_151_p),
    .doutn(ffc_151_n),
    .din(ffc_358_p_spl_1)
  );


  DROC
  ffc_152_1
  (
    .doutp(ffc_152_p),
    .doutn(ffc_152_n),
    .din(ffc_359_p_spl_)
  );


  DROC
  ffc_153_2
  (
    .doutp(ffc_153_p),
    .doutn(ffc_153_n),
    .din(ffc_19_p_spl_)
  );


  DROC
  ffc_154_2
  (
    .doutp(ffc_154_p),
    .doutn(ffc_154_n),
    .din(ffc_21_p_spl_)
  );


  DROC
  ffc_155_2
  (
    .doutp(ffc_155_p),
    .doutn(ffc_155_n),
    .din(ffc_48_p_spl_)
  );


  DROC
  ffc_156_1
  (
    .doutp(ffc_156_p),
    .doutn(ffc_156_n),
    .din(ffc_351_p_spl_)
  );


  DROC
  ffc_157_1
  (
    .doutp(ffc_157_p),
    .doutn(ffc_157_n),
    .din(ffc_352_p_spl_)
  );


  DROC
  ffc_158_2
  (
    .doutp(ffc_158_n),
    .doutn(ffc_158_p),
    .din(g581_n_spl_1)
  );


  DROC
  ffc_159_2
  (
    .doutp(ffc_159_p),
    .doutn(ffc_159_n),
    .din(g583_n_spl_1)
  );


  DROC
  ffc_160_2
  (
    .doutp(ffc_160_p),
    .doutn(ffc_160_n),
    .din(g589_n_spl_)
  );


  DROC
  ffc_161_2
  (
    .doutp(ffc_161_p),
    .doutn(ffc_161_n),
    .din(g590_p_spl_)
  );


  DROC
  ffc_162_1
  (
    .doutp(ffc_162_p),
    .doutn(ffc_162_n),
    .din(ffc_332_p_spl_1)
  );


  DROC
  ffc_163_1
  (
    .doutp(ffc_163_p),
    .doutn(ffc_163_n),
    .din(ffc_333_p_spl_1)
  );


  DROC
  ffc_164_1
  (
    .doutp(ffc_164_p),
    .doutn(ffc_164_n),
    .din(ffc_334_p_spl_)
  );


  DROC
  ffc_165_1
  (
    .doutp(ffc_165_p),
    .doutn(ffc_165_n),
    .din(ffc_335_p_spl_)
  );


  DROC
  ffc_166_1
  (
    .doutp(ffc_166_p),
    .doutn(ffc_166_n),
    .din(ffc_336_p_spl_)
  );


  DROC
  ffc_167_1
  (
    .doutp(ffc_167_p),
    .doutn(ffc_167_n),
    .din(ffc_337_p_spl_)
  );


  DROC
  ffc_168_2
  (
    .doutp(ffc_168_p),
    .doutn(ffc_168_n),
    .din(ffc_15_p_spl_)
  );


  DROC
  ffc_169_2
  (
    .doutp(ffc_169_p),
    .doutn(ffc_169_n),
    .din(ffc_17_p_spl_)
  );


  DROC
  ffc_170_2
  (
    .doutp(ffc_170_n),
    .doutn(ffc_170_p),
    .din(g591_n_spl_)
  );


  DROC
  ffc_171_2
  (
    .doutp(ffc_171_p),
    .doutn(ffc_171_n),
    .din(g592_p)
  );


  DROC
  ffc_172_2
  (
    .doutp(ffc_172_p),
    .doutn(ffc_172_n),
    .din(g595_n_spl_)
  );


  DROC
  ffc_173_2
  (
    .doutp(ffc_173_p),
    .doutn(ffc_173_n),
    .din(g597_p_spl_)
  );


  DROC
  ffc_174_2
  (
    .doutp(ffc_174_p),
    .doutn(ffc_174_n),
    .din(g598_p_spl_)
  );


  DROC
  ffc_175_2
  (
    .doutp(ffc_175_p),
    .doutn(ffc_175_n),
    .din(g599_p_spl_)
  );


  DROC
  ffc_176_3
  (
    .doutp(ffc_176_p),
    .doutn(ffc_176_n),
    .din(g621_n_spl_)
  );


  DROC
  ffc_177_3
  (
    .doutp(ffc_177_p),
    .doutn(ffc_177_n),
    .din(g645_n_spl_)
  );


  DROC
  ffc_178_1
  (
    .doutp(ffc_178_p),
    .doutn(ffc_178_n),
    .din(g646_n_spl_)
  );


  DROC
  ffc_179_2
  (
    .doutp(ffc_179_p),
    .doutn(ffc_179_n),
    .din(g656_p_spl_)
  );


  DROC
  ffc_180_1
  (
    .doutp(ffc_180_p),
    .doutn(ffc_180_n),
    .din(g657_n_spl_)
  );


  DROC
  ffc_181_1
  (
    .doutp(ffc_181_p),
    .doutn(ffc_181_n),
    .din(g658_n_spl_)
  );


  DROC
  ffc_182_1
  (
    .doutp(ffc_182_p),
    .doutn(ffc_182_n),
    .din(g659_n_spl_1)
  );


  DROC
  ffc_183_2
  (
    .doutp(ffc_183_n),
    .doutn(ffc_183_p),
    .din(g660_p_spl_)
  );


  DROC
  ffc_184_2
  (
    .doutp(ffc_184_p),
    .doutn(ffc_184_n),
    .din(g661_n_spl_)
  );


  DROC
  ffc_185_2
  (
    .doutp(ffc_185_n),
    .doutn(ffc_185_p),
    .din(g662_n_spl_)
  );


  DROC
  ffc_186_2
  (
    .doutp(ffc_186_n),
    .doutn(ffc_186_p),
    .din(g663_p_spl_)
  );


  DROC
  ffc_187_2
  (
    .doutp(ffc_187_n),
    .doutn(ffc_187_p),
    .din(g664_n_spl_)
  );


  DROC
  ffc_188_2
  (
    .doutp(ffc_188_p),
    .doutn(ffc_188_n),
    .din(g665_n_spl_)
  );


  DROC
  ffc_189_2
  (
    .doutp(ffc_189_p),
    .doutn(ffc_189_n),
    .din(g666_p_spl_)
  );


  DROC
  ffc_190_1
  (
    .doutp(ffc_190_p),
    .doutn(ffc_190_n),
    .din(g667_n_spl_)
  );


  DROC
  ffc_191_1
  (
    .doutp(ffc_191_p),
    .doutn(ffc_191_n),
    .din(g676_n_spl_)
  );


  DROC
  ffc_192_1
  (
    .doutp(ffc_192_p),
    .doutn(ffc_192_n),
    .din(g684_n_spl_)
  );


  DROC
  ffc_193_1
  (
    .doutp(ffc_193_p),
    .doutn(ffc_193_n),
    .din(g686_p_spl_)
  );


  DROC
  ffc_194_1
  (
    .doutp(ffc_194_p),
    .doutn(ffc_194_n),
    .din(g687_n_spl_)
  );


  DROC
  ffc_195_1
  (
    .doutp(ffc_195_p),
    .doutn(ffc_195_n),
    .din(g691_p_spl_)
  );


  DROC
  ffc_196_1
  (
    .doutp(ffc_196_p),
    .doutn(ffc_196_n),
    .din(ffc_22_p_spl_)
  );


  DROC
  ffc_197_1
  (
    .doutp(ffc_197_p),
    .doutn(ffc_197_n),
    .din(ffc_23_p_spl_)
  );


  DROC
  ffc_198_1
  (
    .doutp(ffc_198_p),
    .doutn(ffc_198_n),
    .din(g701_n_spl_)
  );


  DROC
  ffc_199_1
  (
    .doutp(ffc_199_n),
    .doutn(ffc_199_p),
    .din(g707_n_spl_)
  );


  DROC
  ffc_200_1
  (
    .doutp(ffc_200_n),
    .doutn(ffc_200_p),
    .din(g713_n_spl_)
  );


  DROC
  ffc_201_0
  (
    .doutp(ffc_201_p),
    .doutn(ffc_201_n),
    .din(G1_p_spl_)
  );


  DROC
  ffc_202_0
  (
    .doutp(ffc_202_p),
    .doutn(ffc_202_n),
    .din(G3_p_spl_1)
  );


  DROC
  ffc_203_2
  (
    .doutp(ffc_203_p),
    .doutn(ffc_203_n),
    .din(ffc_37_p_spl_)
  );


  DROC
  ffc_204_2
  (
    .doutp(ffc_204_p),
    .doutn(ffc_204_n),
    .din(ffc_39_p_spl_)
  );


  DROC
  ffc_205_3
  (
    .doutp(ffc_205_n),
    .doutn(ffc_205_p),
    .din(g714_n)
  );


  DROC
  ffc_206_3
  (
    .doutp(ffc_206_n),
    .doutn(ffc_206_p),
    .din(g715_n)
  );


  DROC
  ffc_207_2
  (
    .doutp(ffc_207_p),
    .doutn(ffc_207_n),
    .din(g716_p_spl_)
  );


  DROC
  ffc_208_3
  (
    .doutp(ffc_208_n),
    .doutn(ffc_208_p),
    .din(g718_n)
  );


  DROC
  ffc_209_2
  (
    .doutp(ffc_209_n),
    .doutn(ffc_209_p),
    .din(g719_n_spl_)
  );


  DROC
  ffc_210_2
  (
    .doutp(ffc_210_p),
    .doutn(ffc_210_n),
    .din(g720_n_spl_)
  );


  DROC
  ffc_211_3
  (
    .doutp(ffc_211_p),
    .doutn(ffc_211_n),
    .din(g721_p)
  );


  DROC
  ffc_212_3
  (
    .doutp(ffc_212_p),
    .doutn(ffc_212_n),
    .din(g739_p)
  );


  DROC
  ffc_213_3
  (
    .doutp(ffc_213_p),
    .doutn(ffc_213_n),
    .din(g740_p)
  );


  DROC
  ffc_214_3
  (
    .doutp(ffc_214_p),
    .doutn(ffc_214_n),
    .din(g741_p)
  );


  DROC
  ffc_215_3
  (
    .doutp(ffc_215_p),
    .doutn(ffc_215_n),
    .din(g743_n)
  );


  DROC
  ffc_216_3
  (
    .doutp(ffc_216_n),
    .doutn(ffc_216_p),
    .din(g783_n)
  );


  DROC
  ffc_217_3
  (
    .doutp(ffc_217_n),
    .doutn(ffc_217_p),
    .din(g810_n)
  );


  DROC
  ffc_218_3
  (
    .doutp(ffc_218_p),
    .doutn(ffc_218_n),
    .din(g838_p)
  );


  DROC
  ffc_219_3
  (
    .doutp(ffc_219_p),
    .doutn(ffc_219_n),
    .din(g869_p)
  );


  DROC
  ffc_220_3
  (
    .doutp(ffc_220_n),
    .doutn(ffc_220_p),
    .din(g874_n)
  );


  DROC
  ffc_221_2
  (
    .doutp(ffc_221_n),
    .doutn(ffc_221_p),
    .din(g875_n_spl_)
  );


  DROC
  ffc_222_1
  (
    .doutp(ffc_222_p),
    .doutn(ffc_222_n),
    .din(g876_n_spl_)
  );


  DROC
  ffc_223_2
  (
    .doutp(ffc_223_n),
    .doutn(ffc_223_p),
    .din(g886_n_spl_)
  );


  DROC
  ffc_224_3
  (
    .doutp(ffc_224_p),
    .doutn(ffc_224_n),
    .din(g889_p)
  );


  DROC
  ffc_225_2
  (
    .doutp(ffc_225_n),
    .doutn(ffc_225_p),
    .din(g890_n_spl_)
  );


  DROC
  ffc_226_3
  (
    .doutp(ffc_226_p),
    .doutn(ffc_226_n),
    .din(g916_p)
  );


  DROC
  ffc_227_3
  (
    .doutp(ffc_227_p),
    .doutn(ffc_227_n),
    .din(g919_n)
  );


  DROC
  ffc_228_3
  (
    .doutp(ffc_228_p),
    .doutn(ffc_228_n),
    .din(g945_p)
  );


  DROC
  ffc_229_3
  (
    .doutp(ffc_229_p),
    .doutn(ffc_229_n),
    .din(g948_n)
  );


  DROC
  ffc_230_2
  (
    .doutp(ffc_230_p),
    .doutn(ffc_230_n),
    .din(g950_n_spl_)
  );


  DROC
  ffc_231_3
  (
    .doutp(ffc_231_p),
    .doutn(ffc_231_n),
    .din(g956_n)
  );


  DROC
  ffc_232_3
  (
    .doutp(ffc_232_p),
    .doutn(ffc_232_n),
    .din(g966_n)
  );


  DROC
  ffc_233_3
  (
    .doutp(ffc_233_p),
    .doutn(ffc_233_n),
    .din(g967_n)
  );


  DROC
  ffc_234_3
  (
    .doutp(ffc_234_p),
    .doutn(ffc_234_n),
    .din(g968_p)
  );


  DROC
  ffc_235_2
  (
    .doutp(ffc_235_n),
    .doutn(ffc_235_p),
    .din(g972_n_spl_)
  );


  DROC
  ffc_236_2
  (
    .doutp(ffc_236_n),
    .doutn(ffc_236_p),
    .din(g976_n_spl_)
  );


  DROC
  ffc_237_1
  (
    .doutp(ffc_237_p),
    .doutn(ffc_237_n),
    .din(ffc_24_p)
  );


  DROC
  ffc_238_1
  (
    .doutp(ffc_238_p),
    .doutn(ffc_238_n),
    .din(g985_n_spl_)
  );


  DROC
  ffc_239_1
  (
    .doutp(ffc_239_n),
    .doutn(ffc_239_p),
    .din(g992_n_spl_)
  );


  DROC
  ffc_240_1
  (
    .doutp(ffc_240_p),
    .doutn(ffc_240_n),
    .din(g995_p_spl_)
  );


  DROC
  ffc_241_1
  (
    .doutp(ffc_241_p),
    .doutn(ffc_241_n),
    .din(g998_p_spl_)
  );


  DROC
  ffc_242_0
  (
    .doutp(ffc_242_p),
    .doutn(ffc_242_n),
    .din(G2_p)
  );


  DROC
  ffc_243_0
  (
    .doutp(ffc_243_p),
    .doutn(ffc_243_n),
    .din(G4_p_spl_11)
  );


  DROC
  ffc_244_0
  (
    .doutp(ffc_244_p),
    .doutn(ffc_244_n),
    .din(G6_p_spl_)
  );


  DROC
  ffc_245_0
  (
    .doutp(ffc_245_p),
    .doutn(ffc_245_n),
    .din(G11_p_spl_)
  );


  DROC
  ffc_246_0
  (
    .doutp(ffc_246_p),
    .doutn(ffc_246_n),
    .din(G12_p_spl_1)
  );


  DROC
  ffc_247_0
  (
    .doutp(ffc_247_p),
    .doutn(ffc_247_n),
    .din(G13_p_spl_)
  );


  DROC
  ffc_248_0
  (
    .doutp(ffc_248_p),
    .doutn(ffc_248_n),
    .din(G14_p_spl_)
  );


  DROC
  ffc_249_0
  (
    .doutp(ffc_249_p),
    .doutn(ffc_249_n),
    .din(G33_p_spl_)
  );


  DROC
  ffc_250_0
  (
    .doutp(ffc_250_p),
    .doutn(ffc_250_n),
    .din(G34_p_spl_)
  );


  DROC
  ffc_251_0
  (
    .doutp(ffc_251_p),
    .doutn(ffc_251_n),
    .din(G39_p)
  );


  DROC
  ffc_252_2
  (
    .doutp(ffc_252_p),
    .doutn(ffc_252_n),
    .din(ffc_41_p)
  );


  DROC
  ffc_253_2
  (
    .doutp(ffc_253_p),
    .doutn(ffc_253_n),
    .din(ffc_43_p)
  );


  DROC
  ffc_254_2
  (
    .doutp(ffc_254_p),
    .doutn(ffc_254_n),
    .din(g999_n)
  );


  DROC
  ffc_255_2
  (
    .doutp(ffc_255_p),
    .doutn(ffc_255_n),
    .din(g1000_p)
  );


  DROC
  ffc_256_2
  (
    .doutp(ffc_256_p),
    .doutn(ffc_256_n),
    .din(g1001_p)
  );


  DROC
  ffc_257_2
  (
    .doutp(ffc_257_n),
    .doutn(ffc_257_p),
    .din(g1002_p)
  );


  DROC
  ffc_258_2
  (
    .doutp(ffc_258_p),
    .doutn(ffc_258_n),
    .din(g1003_p)
  );


  DROC
  ffc_259_2
  (
    .doutp(ffc_259_n),
    .doutn(ffc_259_p),
    .din(g1005_n)
  );


  DROC
  ffc_260_2
  (
    .doutp(ffc_260_p),
    .doutn(ffc_260_n),
    .din(g1006_p)
  );


  DROC
  ffc_261_2
  (
    .doutp(ffc_261_p),
    .doutn(ffc_261_n),
    .din(g1007_p)
  );


  DROC
  ffc_262_2
  (
    .doutp(ffc_262_p),
    .doutn(ffc_262_n),
    .din(g1008_p)
  );


  DROC
  ffc_263_2
  (
    .doutp(ffc_263_p),
    .doutn(ffc_263_n),
    .din(g1010_p)
  );


  DROC
  ffc_264_2
  (
    .doutp(ffc_264_p),
    .doutn(ffc_264_n),
    .din(g1011_p)
  );


  DROC
  ffc_265_2
  (
    .doutp(ffc_265_p),
    .doutn(ffc_265_n),
    .din(g1012_p)
  );


  DROC
  ffc_266_2
  (
    .doutp(ffc_266_n),
    .doutn(ffc_266_p),
    .din(g1014_n)
  );


  DROC
  ffc_267_2
  (
    .doutp(ffc_267_p),
    .doutn(ffc_267_n),
    .din(g1015_p)
  );


  DROC
  ffc_268_2
  (
    .doutp(ffc_268_p),
    .doutn(ffc_268_n),
    .din(g1016_p)
  );


  DROC
  ffc_269_2
  (
    .doutp(ffc_269_n),
    .doutn(ffc_269_p),
    .din(g1017_n)
  );


  DROC
  ffc_270_2
  (
    .doutp(ffc_270_p),
    .doutn(ffc_270_n),
    .din(g1018_p)
  );


  DROC
  ffc_271_2
  (
    .doutp(ffc_271_p),
    .doutn(ffc_271_n),
    .din(g1019_p)
  );


  DROC
  ffc_272_2
  (
    .doutp(ffc_272_n),
    .doutn(ffc_272_p),
    .din(g1021_p)
  );


  DROC
  ffc_273_2
  (
    .doutp(ffc_273_n),
    .doutn(ffc_273_p),
    .din(g1022_n)
  );


  DROC
  ffc_274_2
  (
    .doutp(ffc_274_n),
    .doutn(ffc_274_p),
    .din(g1023_p)
  );


  DROC
  ffc_275_2
  (
    .doutp(ffc_275_n),
    .doutn(ffc_275_p),
    .din(g1032_n)
  );


  DROC
  ffc_276_2
  (
    .doutp(ffc_276_p),
    .doutn(ffc_276_n),
    .din(g1033_p)
  );


  DROC
  ffc_277_0
  (
    .doutp(ffc_277_n),
    .doutn(ffc_277_p),
    .din(g1034_n_spl_)
  );


  DROC
  ffc_278_0
  (
    .doutp(ffc_278_p),
    .doutn(ffc_278_n),
    .din(g1035_n_spl_)
  );


  DROC
  ffc_279_1
  (
    .doutp(ffc_279_p),
    .doutn(ffc_279_n),
    .din(ffc_50_p)
  );


  DROC
  ffc_280_2
  (
    .doutp(ffc_280_p),
    .doutn(ffc_280_n),
    .din(g1037_p)
  );


  DROC
  ffc_281_2
  (
    .doutp(ffc_281_n),
    .doutn(ffc_281_p),
    .din(g1044_n)
  );


  DROC
  ffc_282_2
  (
    .doutp(ffc_282_p),
    .doutn(ffc_282_n),
    .din(g1046_p)
  );


  DROC
  ffc_283_2
  (
    .doutp(ffc_283_n),
    .doutn(ffc_283_p),
    .din(g1050_n)
  );


  DROC
  ffc_284_2
  (
    .doutp(ffc_284_p),
    .doutn(ffc_284_n),
    .din(g1053_p)
  );


  DROC
  ffc_285_2
  (
    .doutp(ffc_285_p),
    .doutn(ffc_285_n),
    .din(g1054_p)
  );


  DROC
  ffc_286_2
  (
    .doutp(ffc_286_p),
    .doutn(ffc_286_n),
    .din(g1058_n)
  );


  DROC
  ffc_287_2
  (
    .doutp(ffc_287_p),
    .doutn(ffc_287_n),
    .din(g1063_n)
  );


  DROC
  ffc_288_2
  (
    .doutp(ffc_288_p),
    .doutn(ffc_288_n),
    .din(g1066_n)
  );


  DROC
  ffc_289_2
  (
    .doutp(ffc_289_n),
    .doutn(ffc_289_p),
    .din(g1067_p)
  );


  DROC
  ffc_290_2
  (
    .doutp(ffc_290_n),
    .doutn(ffc_290_p),
    .din(g1073_p)
  );


  DROC
  ffc_291_1
  (
    .doutp(ffc_291_n),
    .doutn(ffc_291_p),
    .din(g1074_n_spl_)
  );


  DROC
  ffc_292_1
  (
    .doutp(ffc_292_p),
    .doutn(ffc_292_n),
    .din(g1085_n_spl_)
  );


  DROC
  ffc_293_2
  (
    .doutp(ffc_293_p),
    .doutn(ffc_293_n),
    .din(g1089_n)
  );


  DROC
  ffc_294_2
  (
    .doutp(ffc_294_p),
    .doutn(ffc_294_n),
    .din(g1090_p)
  );


  DROC
  ffc_295_1
  (
    .doutp(ffc_295_p),
    .doutn(ffc_295_n),
    .din(g1098_n_spl_)
  );


  DROC
  ffc_296_2
  (
    .doutp(ffc_296_p),
    .doutn(ffc_296_n),
    .din(g1101_n)
  );


  DROC
  ffc_297_1
  (
    .doutp(ffc_297_n),
    .doutn(ffc_297_p),
    .din(g1110_n_spl_)
  );


  DROC
  ffc_298_2
  (
    .doutp(ffc_298_n),
    .doutn(ffc_298_p),
    .din(g1117_n)
  );


  DROC
  ffc_299_1
  (
    .doutp(ffc_299_p),
    .doutn(ffc_299_n),
    .din(g1120_p_spl_)
  );


  DROC
  ffc_300_1
  (
    .doutp(ffc_300_p),
    .doutn(ffc_300_n),
    .din(g1121_p_spl_)
  );


  DROC
  ffc_301_0
  (
    .doutp(ffc_301_p),
    .doutn(ffc_301_n),
    .din(G5_p_spl_)
  );


  DROC
  ffc_302_0
  (
    .doutp(ffc_302_p),
    .doutn(ffc_302_n),
    .din(G35_p_spl_)
  );


  DROC
  ffc_303_0
  (
    .doutp(ffc_303_p),
    .doutn(ffc_303_n),
    .din(G40_p_spl_)
  );


  DROC
  ffc_304_0
  (
    .doutp(ffc_304_p),
    .doutn(ffc_304_n),
    .din(g1122_n_spl_1)
  );


  DROC
  ffc_305_0
  (
    .doutp(ffc_305_p),
    .doutn(ffc_305_n),
    .din(g1123_n_spl_)
  );


  DROC
  ffc_306_0
  (
    .doutp(ffc_306_p),
    .doutn(ffc_306_n),
    .din(g1124_n_spl_)
  );


  DROC
  ffc_307_1
  (
    .doutp(ffc_307_p),
    .doutn(ffc_307_n),
    .din(g1130_p)
  );


  DROC
  ffc_308_1
  (
    .doutp(ffc_308_p),
    .doutn(ffc_308_n),
    .din(g1136_p)
  );


  DROC
  ffc_309_1
  (
    .doutp(ffc_309_p),
    .doutn(ffc_309_n),
    .din(g1144_p)
  );


  DROC
  ffc_310_1
  (
    .doutp(ffc_310_p),
    .doutn(ffc_310_n),
    .din(g1148_p)
  );


  DROC
  ffc_311_1
  (
    .doutp(ffc_311_p),
    .doutn(ffc_311_n),
    .din(g1152_p)
  );


  DROC
  ffc_312_1
  (
    .doutp(ffc_312_p),
    .doutn(ffc_312_n),
    .din(g1161_n)
  );


  DROC
  ffc_313_0
  (
    .doutp(ffc_313_n),
    .doutn(ffc_313_p),
    .din(g1162_n_spl_1)
  );


  DROC
  ffc_314_0
  (
    .doutp(ffc_314_n),
    .doutn(ffc_314_p),
    .din(g1162_n_spl_1)
  );


  DROC
  ffc_315_0
  (
    .doutp(ffc_315_n),
    .doutn(ffc_315_p),
    .din(g1163_n_spl_)
  );


  DROC
  ffc_316_0
  (
    .doutp(ffc_316_p),
    .doutn(ffc_316_n),
    .din(g1164_p_spl_)
  );


  DROC
  ffc_317_1
  (
    .doutp(ffc_317_p),
    .doutn(ffc_317_n),
    .din(g1167_p)
  );


  DROC
  ffc_318_1
  (
    .doutp(ffc_318_p),
    .doutn(ffc_318_n),
    .din(g1170_p)
  );


  DROC
  ffc_319_1
  (
    .doutp(ffc_319_p),
    .doutn(ffc_319_n),
    .din(g1181_p)
  );


  DROC
  ffc_320_1
  (
    .doutp(ffc_320_p),
    .doutn(ffc_320_n),
    .din(g1192_p)
  );


  DROC
  ffc_321_1
  (
    .doutp(ffc_321_p),
    .doutn(ffc_321_n),
    .din(g1194_n)
  );


  DROC
  ffc_322_1
  (
    .doutp(ffc_322_p),
    .doutn(ffc_322_n),
    .din(g1196_n)
  );


  DROC
  ffc_323_0
  (
    .doutp(ffc_323_n),
    .doutn(ffc_323_p),
    .din(g1200_p_spl_)
  );


  DROC
  ffc_324_0
  (
    .doutp(ffc_324_p),
    .doutn(ffc_324_n),
    .din(g1201_n_spl_)
  );


  DROC
  ffc_325_0
  (
    .doutp(ffc_325_p),
    .doutn(ffc_325_n),
    .din(G32_p)
  );


  DROC
  ffc_326_0
  (
    .doutp(ffc_326_p),
    .doutn(ffc_326_n),
    .din(G36_p)
  );


  DROC
  ffc_327_0
  (
    .doutp(ffc_327_p),
    .doutn(ffc_327_n),
    .din(G41_p_spl_)
  );


  DROC
  ffc_328_1
  (
    .doutp(ffc_328_n),
    .doutn(ffc_328_p),
    .din(g1202_n)
  );


  DROC
  ffc_329_1
  (
    .doutp(ffc_329_p),
    .doutn(ffc_329_n),
    .din(g1205_p)
  );


  DROC
  ffc_330_1
  (
    .doutp(ffc_330_p),
    .doutn(ffc_330_n),
    .din(g1206_p)
  );


  DROC
  ffc_331_0
  (
    .doutp(ffc_331_p),
    .doutn(ffc_331_n),
    .din(g1208_p_spl_)
  );


  DROC
  ffc_332_0
  (
    .doutp(ffc_332_p),
    .doutn(ffc_332_n),
    .din(G7_p)
  );


  DROC
  ffc_333_0
  (
    .doutp(ffc_333_p),
    .doutn(ffc_333_n),
    .din(G8_p)
  );


  DROC
  ffc_334_0
  (
    .doutp(ffc_334_p),
    .doutn(ffc_334_n),
    .din(G23_p)
  );


  DROC
  ffc_335_0
  (
    .doutp(ffc_335_p),
    .doutn(ffc_335_n),
    .din(G24_p)
  );


  DROC
  ffc_336_0
  (
    .doutp(ffc_336_p),
    .doutn(ffc_336_n),
    .din(G25_p)
  );


  DROC
  ffc_337_0
  (
    .doutp(ffc_337_p),
    .doutn(ffc_337_n),
    .din(G26_p)
  );


  DROC
  ffc_338_0
  (
    .doutp(ffc_338_p),
    .doutn(ffc_338_n),
    .din(g1209_p)
  );


  DROC
  ffc_339_0
  (
    .doutp(ffc_339_p),
    .doutn(ffc_339_n),
    .din(g1210_n_spl_)
  );


  DROC
  ffc_340_0
  (
    .doutp(ffc_340_p),
    .doutn(ffc_340_n),
    .din(g1210_n_spl_)
  );


  DROC
  ffc_341_0
  (
    .doutp(ffc_341_p),
    .doutn(ffc_341_n),
    .din(g1212_p)
  );


  DROC
  ffc_342_0
  (
    .doutp(ffc_342_p),
    .doutn(ffc_342_n),
    .din(g1213_p)
  );


  DROC
  ffc_343_0
  (
    .doutp(ffc_343_p),
    .doutn(ffc_343_n),
    .din(g1214_n)
  );


  DROC
  ffc_344_0
  (
    .doutp(ffc_344_p),
    .doutn(ffc_344_n),
    .din(g1215_p)
  );


  DROC
  ffc_345_0
  (
    .doutp(ffc_345_n),
    .doutn(ffc_345_p),
    .din(g1216_n)
  );


  DROC
  ffc_346_0
  (
    .doutp(ffc_346_n),
    .doutn(ffc_346_p),
    .din(g1217_n)
  );


  DROC
  ffc_347_0
  (
    .doutp(ffc_347_n),
    .doutn(ffc_347_p),
    .din(g1218_n)
  );


  DROC
  ffc_348_0
  (
    .doutp(ffc_348_n),
    .doutn(ffc_348_p),
    .din(g1219_n)
  );


  DROC
  ffc_349_0
  (
    .doutp(ffc_349_p),
    .doutn(ffc_349_n),
    .din(g1220_p)
  );


  DROC
  ffc_350_0
  (
    .doutp(ffc_350_n),
    .doutn(ffc_350_p),
    .din(g1221_n)
  );


  DROC
  ffc_351_0
  (
    .doutp(ffc_351_p),
    .doutn(ffc_351_n),
    .din(G30_p)
  );


  DROC
  ffc_352_0
  (
    .doutp(ffc_352_p),
    .doutn(ffc_352_n),
    .din(G37_p)
  );


  DROC
  ffc_353_0
  (
    .doutp(ffc_353_n),
    .doutn(ffc_353_p),
    .din(g1222_p)
  );


  DROC
  ffc_354_0
  (
    .doutp(ffc_354_p),
    .doutn(ffc_354_n),
    .din(g1225_p)
  );


  DROC
  ffc_355_0
  (
    .doutp(ffc_355_n),
    .doutn(ffc_355_p),
    .din(g1230_p)
  );


  DROC
  ffc_356_0
  (
    .doutp(ffc_356_p),
    .doutn(ffc_356_n),
    .din(g1235_n)
  );


  DROC
  ffc_357_0
  (
    .doutp(ffc_357_p),
    .doutn(ffc_357_n),
    .din(G9_p)
  );


  DROC
  ffc_358_0
  (
    .doutp(ffc_358_p),
    .doutn(ffc_358_n),
    .din(G10_p)
  );


  DROC
  ffc_359_0
  (
    .doutp(ffc_359_p),
    .doutn(ffc_359_n),
    .din(G31_p)
  );


  DROC
  ffc_360_0
  (
    .doutp(ffc_360_p),
    .doutn(ffc_360_n),
    .din(G38_p)
  );


  buf

  (
    ffc_5_n_spl_,
    ffc_5_n
  );


  buf

  (
    ffc_0_n_spl_,
    ffc_0_n
  );


  buf

  (
    ffc_1_n_spl_,
    ffc_1_n
  );


  buf

  (
    ffc_6_p_spl_,
    ffc_6_p
  );


  buf

  (
    ffc_32_n_spl_,
    ffc_32_n
  );


  buf

  (
    ffc_32_n_spl_0,
    ffc_32_n_spl_
  );


  buf

  (
    ffc_32_n_spl_1,
    ffc_32_n_spl_
  );


  buf

  (
    ffc_30_n_spl_,
    ffc_30_n
  );


  buf

  (
    ffc_30_n_spl_0,
    ffc_30_n_spl_
  );


  buf

  (
    ffc_2_p_spl_,
    ffc_2_p
  );


  buf

  (
    ffc_28_n_spl_,
    ffc_28_n
  );


  buf

  (
    ffc_28_n_spl_0,
    ffc_28_n_spl_
  );


  buf

  (
    ffc_31_n_spl_,
    ffc_31_n
  );


  buf

  (
    ffc_31_n_spl_0,
    ffc_31_n_spl_
  );


  buf

  (
    ffc_9_p_spl_,
    ffc_9_p
  );


  buf

  (
    ffc_9_p_spl_0,
    ffc_9_p_spl_
  );


  buf

  (
    ffc_35_n_spl_,
    ffc_35_n
  );


  buf

  (
    ffc_35_n_spl_0,
    ffc_35_n_spl_
  );


  buf

  (
    ffc_29_n_spl_,
    ffc_29_n
  );


  buf

  (
    ffc_29_n_spl_0,
    ffc_29_n_spl_
  );


  buf

  (
    ffc_7_p_spl_,
    ffc_7_p
  );


  buf

  (
    ffc_33_n_spl_,
    ffc_33_n
  );


  buf

  (
    ffc_33_n_spl_0,
    ffc_33_n_spl_
  );


  buf

  (
    ffc_33_n_spl_1,
    ffc_33_n_spl_
  );


  buf

  (
    ffc_8_p_spl_,
    ffc_8_p
  );


  buf

  (
    ffc_8_p_spl_0,
    ffc_8_p_spl_
  );


  buf

  (
    ffc_34_n_spl_,
    ffc_34_n
  );


  buf

  (
    ffc_34_n_spl_0,
    ffc_34_n_spl_
  );


  buf

  (
    ffc_34_n_spl_1,
    ffc_34_n_spl_
  );


  buf

  (
    g430_n_spl_,
    g430_n
  );


  buf

  (
    ffc_34_p_spl_,
    ffc_34_p
  );


  buf

  (
    ffc_35_p_spl_,
    ffc_35_p
  );


  buf

  (
    ffc_32_p_spl_,
    ffc_32_p
  );


  buf

  (
    ffc_33_p_spl_,
    ffc_33_p
  );


  buf

  (
    g439_n_spl_,
    g439_n
  );


  buf

  (
    g442_p_spl_,
    g442_p
  );


  buf

  (
    g439_p_spl_,
    g439_p
  );


  buf

  (
    g442_n_spl_,
    g442_n
  );


  buf

  (
    ffc_30_p_spl_,
    ffc_30_p
  );


  buf

  (
    ffc_31_p_spl_,
    ffc_31_p
  );


  buf

  (
    ffc_28_p_spl_,
    ffc_28_p
  );


  buf

  (
    ffc_29_p_spl_,
    ffc_29_p
  );


  buf

  (
    g448_p_spl_,
    g448_p
  );


  buf

  (
    g451_n_spl_,
    g451_n
  );


  buf

  (
    g448_n_spl_,
    g448_n
  );


  buf

  (
    g451_p_spl_,
    g451_p
  );


  buf

  (
    ffc_9_n_spl_,
    ffc_9_n
  );


  buf

  (
    ffc_9_n_spl_0,
    ffc_9_n_spl_
  );


  buf

  (
    ffc_8_n_spl_,
    ffc_8_n
  );


  buf

  (
    g459_p_spl_,
    g459_p
  );


  buf

  (
    g462_p_spl_,
    g462_p
  );


  buf

  (
    g459_n_spl_,
    g459_n
  );


  buf

  (
    g462_n_spl_,
    g462_n
  );


  buf

  (
    ffc_79_p_spl_,
    ffc_79_p
  );


  buf

  (
    ffc_106_n_spl_,
    ffc_106_n
  );


  buf

  (
    ffc_106_n_spl_0,
    ffc_106_n_spl_
  );


  buf

  (
    ffc_115_n_spl_,
    ffc_115_n
  );


  buf

  (
    ffc_115_p_spl_,
    ffc_115_p
  );


  buf

  (
    ffc_90_p_spl_,
    ffc_90_p
  );


  buf

  (
    g481_n_spl_,
    g481_n
  );


  buf

  (
    ffc_90_n_spl_,
    ffc_90_n
  );


  buf

  (
    g481_p_spl_,
    g481_p
  );


  buf

  (
    ffc_101_p_spl_,
    ffc_101_p
  );


  buf

  (
    ffc_102_p_spl_,
    ffc_102_p
  );


  buf

  (
    ffc_101_n_spl_,
    ffc_101_n
  );


  buf

  (
    ffc_102_n_spl_,
    ffc_102_n
  );


  buf

  (
    ffc_106_p_spl_,
    ffc_106_p
  );


  buf

  (
    g480_p_spl_,
    g480_p
  );


  buf

  (
    g514_p_spl_,
    g514_p
  );


  buf

  (
    g480_n_spl_,
    g480_n
  );


  buf

  (
    g480_n_spl_0,
    g480_n_spl_
  );


  buf

  (
    g514_n_spl_,
    g514_n
  );


  buf

  (
    g514_n_spl_0,
    g514_n_spl_
  );


  buf

  (
    g505_p_spl_,
    g505_p
  );


  buf

  (
    g511_p_spl_,
    g511_p
  );


  buf

  (
    g505_n_spl_,
    g505_n
  );


  buf

  (
    g505_n_spl_0,
    g505_n_spl_
  );


  buf

  (
    g511_n_spl_,
    g511_n
  );


  buf

  (
    g511_n_spl_0,
    g511_n_spl_
  );


  buf

  (
    g477_p_spl_,
    g477_p
  );


  buf

  (
    g508_p_spl_,
    g508_p
  );


  buf

  (
    g477_n_spl_,
    g477_n
  );


  buf

  (
    g477_n_spl_0,
    g477_n_spl_
  );


  buf

  (
    g508_n_spl_,
    g508_n
  );


  buf

  (
    g508_n_spl_0,
    g508_n_spl_
  );


  buf

  (
    g516_n_spl_,
    g516_n
  );


  buf

  (
    g517_n_spl_,
    g517_n
  );


  buf

  (
    g515_n_spl_,
    g515_n
  );


  buf

  (
    ffc_233_p_spl_,
    ffc_233_p
  );


  buf

  (
    ffc_233_p_spl_0,
    ffc_233_p_spl_
  );


  buf

  (
    ffc_25_p_spl_,
    ffc_25_p
  );


  buf

  (
    g521_n_spl_,
    g521_n
  );


  buf

  (
    g520_n_spl_,
    g520_n
  );


  buf

  (
    g526_p_spl_,
    g526_p
  );


  buf

  (
    g528_n_spl_,
    g528_n
  );


  buf

  (
    g526_n_spl_,
    g526_n
  );


  buf

  (
    g528_p_spl_,
    g528_p
  );


  buf

  (
    ffc_55_p_spl_,
    ffc_55_p
  );


  buf

  (
    g534_n_spl_,
    g534_n
  );


  buf

  (
    g534_n_spl_0,
    g534_n_spl_
  );


  buf

  (
    g534_n_spl_1,
    g534_n_spl_
  );


  buf

  (
    ffc_55_n_spl_,
    ffc_55_n
  );


  buf

  (
    g534_p_spl_,
    g534_p
  );


  buf

  (
    g534_p_spl_0,
    g534_p_spl_
  );


  buf

  (
    g534_p_spl_1,
    g534_p_spl_
  );


  buf

  (
    g533_p_spl_,
    g533_p
  );


  buf

  (
    g533_p_spl_0,
    g533_p_spl_
  );


  buf

  (
    g533_p_spl_1,
    g533_p_spl_
  );


  buf

  (
    g538_p_spl_,
    g538_p
  );


  buf

  (
    g533_n_spl_,
    g533_n
  );


  buf

  (
    g533_n_spl_0,
    g533_n_spl_
  );


  buf

  (
    g533_n_spl_1,
    g533_n_spl_
  );


  buf

  (
    g538_n_spl_,
    g538_n
  );


  buf

  (
    g531_n_spl_,
    g531_n
  );


  buf

  (
    g531_p_spl_,
    g531_p
  );


  buf

  (
    ffc_103_p_spl_,
    ffc_103_p
  );


  buf

  (
    ffc_103_p_spl_0,
    ffc_103_p_spl_
  );


  buf

  (
    ffc_103_p_spl_1,
    ffc_103_p_spl_
  );


  buf

  (
    ffc_72_n_spl_,
    ffc_72_n
  );


  buf

  (
    ffc_235_n_spl_,
    ffc_235_n
  );


  buf

  (
    ffc_235_n_spl_0,
    ffc_235_n_spl_
  );


  buf

  (
    ffc_235_p_spl_,
    ffc_235_p
  );


  buf

  (
    ffc_290_p_spl_,
    ffc_290_p
  );


  buf

  (
    ffc_118_n_spl_,
    ffc_118_n
  );


  buf

  (
    ffc_118_p_spl_,
    ffc_118_p
  );


  buf

  (
    ffc_118_p_spl_0,
    ffc_118_p_spl_
  );


  buf

  (
    ffc_71_p_spl_,
    ffc_71_p
  );


  buf

  (
    ffc_71_n_spl_,
    ffc_71_n
  );


  buf

  (
    ffc_254_p_spl_,
    ffc_254_p
  );


  buf

  (
    ffc_67_p_spl_,
    ffc_67_p
  );


  buf

  (
    g556_p_spl_,
    g556_p
  );


  buf

  (
    g556_p_spl_0,
    g556_p_spl_
  );


  buf

  (
    g561_p_spl_,
    g561_p
  );


  buf

  (
    g556_n_spl_,
    g556_n
  );


  buf

  (
    g556_n_spl_0,
    g556_n_spl_
  );


  buf

  (
    g556_n_spl_1,
    g556_n_spl_
  );


  buf

  (
    g561_n_spl_,
    g561_n
  );


  buf

  (
    g561_n_spl_0,
    g561_n_spl_
  );


  buf

  (
    g561_n_spl_00,
    g561_n_spl_0
  );


  buf

  (
    g561_n_spl_01,
    g561_n_spl_0
  );


  buf

  (
    g561_n_spl_1,
    g561_n_spl_
  );


  buf

  (
    ffc_329_p_spl_,
    ffc_329_p
  );


  buf

  (
    ffc_330_p_spl_,
    ffc_330_p
  );


  buf

  (
    ffc_329_n_spl_,
    ffc_329_n
  );


  buf

  (
    ffc_330_n_spl_,
    ffc_330_n
  );


  buf

  (
    ffc_328_n_spl_,
    ffc_328_n
  );


  buf

  (
    ffc_328_n_spl_0,
    ffc_328_n_spl_
  );


  buf

  (
    ffc_328_n_spl_00,
    ffc_328_n_spl_0
  );


  buf

  (
    ffc_328_n_spl_000,
    ffc_328_n_spl_00
  );


  buf

  (
    ffc_328_n_spl_001,
    ffc_328_n_spl_00
  );


  buf

  (
    ffc_328_n_spl_01,
    ffc_328_n_spl_0
  );


  buf

  (
    ffc_328_n_spl_1,
    ffc_328_n_spl_
  );


  buf

  (
    ffc_328_n_spl_10,
    ffc_328_n_spl_1
  );


  buf

  (
    ffc_328_n_spl_11,
    ffc_328_n_spl_1
  );


  buf

  (
    ffc_328_p_spl_,
    ffc_328_p
  );


  buf

  (
    ffc_328_p_spl_0,
    ffc_328_p_spl_
  );


  buf

  (
    ffc_328_p_spl_00,
    ffc_328_p_spl_0
  );


  buf

  (
    ffc_328_p_spl_000,
    ffc_328_p_spl_00
  );


  buf

  (
    ffc_328_p_spl_001,
    ffc_328_p_spl_00
  );


  buf

  (
    ffc_328_p_spl_01,
    ffc_328_p_spl_0
  );


  buf

  (
    ffc_328_p_spl_010,
    ffc_328_p_spl_01
  );


  buf

  (
    ffc_328_p_spl_011,
    ffc_328_p_spl_01
  );


  buf

  (
    ffc_328_p_spl_1,
    ffc_328_p_spl_
  );


  buf

  (
    ffc_328_p_spl_10,
    ffc_328_p_spl_1
  );


  buf

  (
    ffc_328_p_spl_11,
    ffc_328_p_spl_1
  );


  buf

  (
    g563_p_spl_,
    g563_p
  );


  buf

  (
    ffc_319_n_spl_,
    ffc_319_n
  );


  buf

  (
    ffc_319_n_spl_0,
    ffc_319_n_spl_
  );


  buf

  (
    ffc_319_p_spl_,
    ffc_319_p
  );


  buf

  (
    g568_n_spl_,
    g568_n
  );


  buf

  (
    g568_n_spl_0,
    g568_n_spl_
  );


  buf

  (
    g569_n_spl_,
    g569_n
  );


  buf

  (
    g568_p_spl_,
    g568_p
  );


  buf

  (
    g569_p_spl_,
    g569_p
  );


  buf

  (
    ffc_320_n_spl_,
    ffc_320_n
  );


  buf

  (
    ffc_320_n_spl_0,
    ffc_320_n_spl_
  );


  buf

  (
    ffc_320_p_spl_,
    ffc_320_p
  );


  buf

  (
    g573_n_spl_,
    g573_n
  );


  buf

  (
    g573_n_spl_0,
    g573_n_spl_
  );


  buf

  (
    g574_n_spl_,
    g574_n
  );


  buf

  (
    g573_p_spl_,
    g573_p
  );


  buf

  (
    g574_p_spl_,
    g574_p
  );


  buf

  (
    ffc_124_p_spl_,
    ffc_124_p
  );


  buf

  (
    ffc_124_p_spl_0,
    ffc_124_p_spl_
  );


  buf

  (
    ffc_124_p_spl_00,
    ffc_124_p_spl_0
  );


  buf

  (
    ffc_124_p_spl_1,
    ffc_124_p_spl_
  );


  buf

  (
    ffc_124_n_spl_,
    ffc_124_n
  );


  buf

  (
    ffc_124_n_spl_0,
    ffc_124_n_spl_
  );


  buf

  (
    ffc_167_n_spl_,
    ffc_167_n
  );


  buf

  (
    g579_p_spl_,
    g579_p
  );


  buf

  (
    g579_p_spl_0,
    g579_p_spl_
  );


  buf

  (
    g579_p_spl_00,
    g579_p_spl_0
  );


  buf

  (
    g579_p_spl_01,
    g579_p_spl_0
  );


  buf

  (
    g579_p_spl_1,
    g579_p_spl_
  );


  buf

  (
    g578_p_spl_,
    g578_p
  );


  buf

  (
    g578_p_spl_0,
    g578_p_spl_
  );


  buf

  (
    g578_p_spl_1,
    g578_p_spl_
  );


  buf

  (
    ffc_167_p_spl_,
    ffc_167_p
  );


  buf

  (
    ffc_297_n_spl_,
    ffc_297_n
  );


  buf

  (
    ffc_239_p_spl_,
    ffc_239_p
  );


  buf

  (
    ffc_200_p_spl_,
    ffc_200_p
  );


  buf

  (
    ffc_240_p_spl_,
    ffc_240_p
  );


  buf

  (
    g567_p_spl_,
    g567_p
  );


  buf

  (
    g567_p_spl_0,
    g567_p_spl_
  );


  buf

  (
    g572_p_spl_,
    g572_p
  );


  buf

  (
    g572_p_spl_0,
    g572_p_spl_
  );


  buf

  (
    ffc_19_p_spl_,
    ffc_19_p
  );


  buf

  (
    ffc_19_p_spl_0,
    ffc_19_p_spl_
  );


  buf

  (
    ffc_162_n_spl_,
    ffc_162_n
  );


  buf

  (
    g589_n_spl_,
    g589_n
  );


  buf

  (
    g578_n_spl_,
    g578_n
  );


  buf

  (
    g593_n_spl_,
    g593_n
  );


  buf

  (
    g593_p_spl_,
    g593_p
  );


  buf

  (
    g579_n_spl_,
    g579_n
  );


  buf

  (
    g579_n_spl_0,
    g579_n_spl_
  );


  buf

  (
    g579_n_spl_1,
    g579_n_spl_
  );


  buf

  (
    g594_p_spl_,
    g594_p
  );


  buf

  (
    g594_n_spl_,
    g594_n
  );


  buf

  (
    g596_p_spl_,
    g596_p
  );


  buf

  (
    g596_n_spl_,
    g596_n
  );


  buf

  (
    ffc_275_n_spl_,
    ffc_275_n
  );


  buf

  (
    ffc_275_p_spl_,
    ffc_275_p
  );


  buf

  (
    ffc_155_p_spl_,
    ffc_155_p
  );


  buf

  (
    ffc_155_p_spl_0,
    ffc_155_p_spl_
  );


  buf

  (
    ffc_155_p_spl_1,
    ffc_155_p_spl_
  );


  buf

  (
    ffc_267_p_spl_,
    ffc_267_p
  );


  buf

  (
    ffc_155_n_spl_,
    ffc_155_n
  );


  buf

  (
    ffc_155_n_spl_0,
    ffc_155_n_spl_
  );


  buf

  (
    ffc_155_n_spl_1,
    ffc_155_n_spl_
  );


  buf

  (
    g555_p_spl_,
    g555_p
  );


  buf

  (
    g601_n_spl_,
    g601_n
  );


  buf

  (
    g601_n_spl_0,
    g601_n_spl_
  );


  buf

  (
    g603_n_spl_,
    g603_n
  );


  buf

  (
    g601_p_spl_,
    g601_p
  );


  buf

  (
    g603_p_spl_,
    g603_p
  );


  buf

  (
    g604_n_spl_,
    g604_n
  );


  buf

  (
    g600_n_spl_,
    g600_n
  );


  buf

  (
    g600_n_spl_0,
    g600_n_spl_
  );


  buf

  (
    ffc_70_n_spl_,
    ffc_70_n
  );


  buf

  (
    ffc_70_n_spl_0,
    ffc_70_n_spl_
  );


  buf

  (
    ffc_70_n_spl_00,
    ffc_70_n_spl_0
  );


  buf

  (
    ffc_70_n_spl_01,
    ffc_70_n_spl_0
  );


  buf

  (
    ffc_70_n_spl_1,
    ffc_70_n_spl_
  );


  buf

  (
    ffc_70_n_spl_10,
    ffc_70_n_spl_1
  );


  buf

  (
    g609_n_spl_,
    g609_n
  );


  buf

  (
    g609_n_spl_0,
    g609_n_spl_
  );


  buf

  (
    g609_n_spl_1,
    g609_n_spl_
  );


  buf

  (
    ffc_68_p_spl_,
    ffc_68_p
  );


  buf

  (
    ffc_84_p_spl_,
    ffc_84_p
  );


  buf

  (
    g612_p_spl_,
    g612_p
  );


  buf

  (
    g612_p_spl_0,
    g612_p_spl_
  );


  buf

  (
    g612_p_spl_00,
    g612_p_spl_0
  );


  buf

  (
    g612_p_spl_01,
    g612_p_spl_0
  );


  buf

  (
    g612_p_spl_1,
    g612_p_spl_
  );


  buf

  (
    g612_p_spl_10,
    g612_p_spl_1
  );


  buf

  (
    g562_p_spl_,
    g562_p
  );


  buf

  (
    g562_p_spl_0,
    g562_p_spl_
  );


  buf

  (
    g562_p_spl_00,
    g562_p_spl_0
  );


  buf

  (
    g562_p_spl_01,
    g562_p_spl_0
  );


  buf

  (
    g562_p_spl_1,
    g562_p_spl_
  );


  buf

  (
    g562_p_spl_10,
    g562_p_spl_1
  );


  buf

  (
    g622_n_spl_,
    g622_n
  );


  buf

  (
    g622_n_spl_0,
    g622_n_spl_
  );


  buf

  (
    g554_n_spl_,
    g554_n
  );


  buf

  (
    g554_n_spl_0,
    g554_n_spl_
  );


  buf

  (
    g554_p_spl_,
    g554_p
  );


  buf

  (
    g622_p_spl_,
    g622_p
  );


  buf

  (
    ffc_333_p_spl_,
    ffc_333_p
  );


  buf

  (
    ffc_333_p_spl_0,
    ffc_333_p_spl_
  );


  buf

  (
    ffc_333_p_spl_1,
    ffc_333_p_spl_
  );


  buf

  (
    ffc_357_p_spl_,
    ffc_357_p
  );


  buf

  (
    ffc_357_p_spl_0,
    ffc_357_p_spl_
  );


  buf

  (
    ffc_357_p_spl_00,
    ffc_357_p_spl_0
  );


  buf

  (
    ffc_357_p_spl_1,
    ffc_357_p_spl_
  );


  buf

  (
    ffc_312_n_spl_,
    ffc_312_n
  );


  buf

  (
    ffc_182_n_spl_,
    ffc_182_n
  );


  buf

  (
    ffc_312_p_spl_,
    ffc_312_p
  );


  buf

  (
    g648_p_spl_,
    g648_p
  );


  buf

  (
    g648_p_spl_0,
    g648_p_spl_
  );


  buf

  (
    g648_n_spl_,
    g648_n
  );


  buf

  (
    g648_n_spl_0,
    g648_n_spl_
  );


  buf

  (
    ffc_181_p_spl_,
    ffc_181_p
  );


  buf

  (
    ffc_181_n_spl_,
    ffc_181_n
  );


  buf

  (
    g651_n_spl_,
    g651_n
  );


  buf

  (
    g651_p_spl_,
    g651_p
  );


  buf

  (
    ffc_291_n_spl_,
    ffc_291_n
  );


  buf

  (
    ffc_291_n_spl_0,
    ffc_291_n_spl_
  );


  buf

  (
    g652_n_spl_,
    g652_n
  );


  buf

  (
    g652_n_spl_0,
    g652_n_spl_
  );


  buf

  (
    g653_n_spl_,
    g653_n
  );


  buf

  (
    g652_p_spl_,
    g652_p
  );


  buf

  (
    g653_p_spl_,
    g653_p
  );


  buf

  (
    ffc_332_p_spl_,
    ffc_332_p
  );


  buf

  (
    ffc_332_p_spl_0,
    ffc_332_p_spl_
  );


  buf

  (
    ffc_332_p_spl_1,
    ffc_332_p_spl_
  );


  buf

  (
    ffc_335_n_spl_,
    ffc_335_n
  );


  buf

  (
    ffc_334_p_spl_,
    ffc_334_p
  );


  buf

  (
    ffc_335_p_spl_,
    ffc_335_p
  );


  buf

  (
    ffc_335_p_spl_0,
    ffc_335_p_spl_
  );


  buf

  (
    ffc_336_p_spl_,
    ffc_336_p
  );


  buf

  (
    ffc_337_p_spl_,
    ffc_337_p
  );


  buf

  (
    ffc_129_n_spl_,
    ffc_129_n
  );


  buf

  (
    g599_n_spl_,
    g599_n
  );


  buf

  (
    g599_n_spl_0,
    g599_n_spl_
  );


  buf

  (
    ffc_131_p_spl_,
    ffc_131_p
  );


  buf

  (
    g597_p_spl_,
    g597_p
  );


  buf

  (
    g597_p_spl_0,
    g597_p_spl_
  );


  buf

  (
    g598_p_spl_,
    g598_p
  );


  buf

  (
    ffc_150_n_spl_,
    ffc_150_n
  );


  buf

  (
    g597_n_spl_,
    g597_n
  );


  buf

  (
    g597_n_spl_0,
    g597_n_spl_
  );


  buf

  (
    g597_n_spl_1,
    g597_n_spl_
  );


  buf

  (
    ffc_151_p_spl_,
    ffc_151_p
  );


  buf

  (
    ffc_151_p_spl_0,
    ffc_151_p_spl_
  );


  buf

  (
    ffc_151_p_spl_00,
    ffc_151_p_spl_0
  );


  buf

  (
    ffc_151_p_spl_1,
    ffc_151_p_spl_
  );


  buf

  (
    g595_p_spl_,
    g595_p
  );


  buf

  (
    ffc_17_p_spl_,
    ffc_17_p
  );


  buf

  (
    ffc_17_p_spl_0,
    ffc_17_p_spl_
  );


  buf

  (
    ffc_197_p_spl_,
    ffc_197_p
  );


  buf

  (
    ffc_197_p_spl_0,
    ffc_197_p_spl_
  );


  buf

  (
    g592_n_spl_,
    g592_n
  );


  buf

  (
    g657_n_spl_,
    g657_n
  );


  buf

  (
    ffc_353_n_spl_,
    ffc_353_n
  );


  buf

  (
    ffc_245_p_spl_,
    ffc_245_p
  );


  buf

  (
    ffc_245_p_spl_0,
    ffc_245_p_spl_
  );


  buf

  (
    ffc_245_p_spl_00,
    ffc_245_p_spl_0
  );


  buf

  (
    ffc_245_p_spl_1,
    ffc_245_p_spl_
  );


  buf

  (
    g668_n_spl_,
    g668_n
  );


  buf

  (
    g668_n_spl_0,
    g668_n_spl_
  );


  buf

  (
    g668_n_spl_1,
    g668_n_spl_
  );


  buf

  (
    ffc_245_n_spl_,
    ffc_245_n
  );


  buf

  (
    ffc_245_n_spl_0,
    ffc_245_n_spl_
  );


  buf

  (
    ffc_245_n_spl_1,
    ffc_245_n_spl_
  );


  buf

  (
    g668_p_spl_,
    g668_p
  );


  buf

  (
    g668_p_spl_0,
    g668_p_spl_
  );


  buf

  (
    g668_p_spl_1,
    g668_p_spl_
  );


  buf

  (
    ffc_315_n_spl_,
    ffc_315_n
  );


  buf

  (
    ffc_315_n_spl_0,
    ffc_315_n_spl_
  );


  buf

  (
    ffc_315_n_spl_1,
    ffc_315_n_spl_
  );


  buf

  (
    ffc_315_p_spl_,
    ffc_315_p
  );


  buf

  (
    ffc_315_p_spl_0,
    ffc_315_p_spl_
  );


  buf

  (
    ffc_315_p_spl_00,
    ffc_315_p_spl_0
  );


  buf

  (
    ffc_315_p_spl_01,
    ffc_315_p_spl_0
  );


  buf

  (
    ffc_315_p_spl_1,
    ffc_315_p_spl_
  );


  buf

  (
    ffc_315_p_spl_10,
    ffc_315_p_spl_1
  );


  buf

  (
    ffc_339_n_spl_,
    ffc_339_n
  );


  buf

  (
    ffc_339_n_spl_0,
    ffc_339_n_spl_
  );


  buf

  (
    ffc_339_n_spl_1,
    ffc_339_n_spl_
  );


  buf

  (
    ffc_357_n_spl_,
    ffc_357_n
  );


  buf

  (
    ffc_357_n_spl_0,
    ffc_357_n_spl_
  );


  buf

  (
    ffc_357_n_spl_1,
    ffc_357_n_spl_
  );


  buf

  (
    ffc_339_p_spl_,
    ffc_339_p
  );


  buf

  (
    ffc_339_p_spl_0,
    ffc_339_p_spl_
  );


  buf

  (
    ffc_323_p_spl_,
    ffc_323_p
  );


  buf

  (
    ffc_323_p_spl_0,
    ffc_323_p_spl_
  );


  buf

  (
    ffc_323_p_spl_00,
    ffc_323_p_spl_0
  );


  buf

  (
    ffc_323_p_spl_000,
    ffc_323_p_spl_00
  );


  buf

  (
    ffc_323_p_spl_01,
    ffc_323_p_spl_0
  );


  buf

  (
    ffc_323_p_spl_1,
    ffc_323_p_spl_
  );


  buf

  (
    ffc_323_p_spl_10,
    ffc_323_p_spl_1
  );


  buf

  (
    ffc_323_p_spl_11,
    ffc_323_p_spl_1
  );


  buf

  (
    ffc_323_n_spl_,
    ffc_323_n
  );


  buf

  (
    ffc_323_n_spl_0,
    ffc_323_n_spl_
  );


  buf

  (
    ffc_323_n_spl_00,
    ffc_323_n_spl_0
  );


  buf

  (
    ffc_323_n_spl_1,
    ffc_323_n_spl_
  );


  buf

  (
    ffc_246_p_spl_,
    ffc_246_p
  );


  buf

  (
    ffc_246_p_spl_0,
    ffc_246_p_spl_
  );


  buf

  (
    ffc_246_p_spl_1,
    ffc_246_p_spl_
  );


  buf

  (
    ffc_246_n_spl_,
    ffc_246_n
  );


  buf

  (
    ffc_246_n_spl_0,
    ffc_246_n_spl_
  );


  buf

  (
    ffc_246_n_spl_1,
    ffc_246_n_spl_
  );


  buf

  (
    ffc_340_n_spl_,
    ffc_340_n
  );


  buf

  (
    ffc_340_n_spl_0,
    ffc_340_n_spl_
  );


  buf

  (
    ffc_340_n_spl_1,
    ffc_340_n_spl_
  );


  buf

  (
    ffc_358_p_spl_,
    ffc_358_p
  );


  buf

  (
    ffc_358_p_spl_0,
    ffc_358_p_spl_
  );


  buf

  (
    ffc_358_p_spl_00,
    ffc_358_p_spl_0
  );


  buf

  (
    ffc_358_p_spl_1,
    ffc_358_p_spl_
  );


  buf

  (
    ffc_358_n_spl_,
    ffc_358_n
  );


  buf

  (
    ffc_333_n_spl_,
    ffc_333_n
  );


  buf

  (
    ffc_333_n_spl_0,
    ffc_333_n_spl_
  );


  buf

  (
    ffc_333_n_spl_1,
    ffc_333_n_spl_
  );


  buf

  (
    g646_n_spl_,
    g646_n
  );


  buf

  (
    ffc_201_p_spl_,
    ffc_201_p
  );


  buf

  (
    ffc_201_p_spl_0,
    ffc_201_p_spl_
  );


  buf

  (
    ffc_201_p_spl_1,
    ffc_201_p_spl_
  );


  buf

  (
    ffc_242_p_spl_,
    ffc_242_p
  );


  buf

  (
    ffc_348_n_spl_,
    ffc_348_n
  );


  buf

  (
    ffc_348_n_spl_0,
    ffc_348_n_spl_
  );


  buf

  (
    ffc_348_n_spl_00,
    ffc_348_n_spl_0
  );


  buf

  (
    ffc_348_n_spl_01,
    ffc_348_n_spl_0
  );


  buf

  (
    ffc_348_n_spl_1,
    ffc_348_n_spl_
  );


  buf

  (
    ffc_348_n_spl_10,
    ffc_348_n_spl_1
  );


  buf

  (
    ffc_348_p_spl_,
    ffc_348_p
  );


  buf

  (
    ffc_348_p_spl_0,
    ffc_348_p_spl_
  );


  buf

  (
    ffc_348_p_spl_00,
    ffc_348_p_spl_0
  );


  buf

  (
    ffc_348_p_spl_01,
    ffc_348_p_spl_0
  );


  buf

  (
    ffc_348_p_spl_1,
    ffc_348_p_spl_
  );


  buf

  (
    ffc_348_p_spl_10,
    ffc_348_p_spl_1
  );


  buf

  (
    ffc_244_p_spl_,
    ffc_244_p
  );


  buf

  (
    ffc_301_p_spl_,
    ffc_301_p
  );


  buf

  (
    g688_p_spl_,
    g688_p
  );


  buf

  (
    g688_p_spl_0,
    g688_p_spl_
  );


  buf

  (
    g690_p_spl_,
    g690_p
  );


  buf

  (
    g690_p_spl_0,
    g690_p_spl_
  );


  buf

  (
    g688_n_spl_,
    g688_n
  );


  buf

  (
    g688_n_spl_0,
    g688_n_spl_
  );


  buf

  (
    g690_n_spl_,
    g690_n
  );


  buf

  (
    g690_n_spl_0,
    g690_n_spl_
  );


  buf

  (
    ffc_202_p_spl_,
    ffc_202_p
  );


  buf

  (
    ffc_202_p_spl_0,
    ffc_202_p_spl_
  );


  buf

  (
    ffc_202_p_spl_00,
    ffc_202_p_spl_0
  );


  buf

  (
    ffc_202_p_spl_1,
    ffc_202_p_spl_
  );


  buf

  (
    ffc_202_n_spl_,
    ffc_202_n
  );


  buf

  (
    g692_n_spl_,
    g692_n
  );


  buf

  (
    g692_p_spl_,
    g692_p
  );


  buf

  (
    g692_p_spl_0,
    g692_p_spl_
  );


  buf

  (
    ffc_247_n_spl_,
    ffc_247_n
  );


  buf

  (
    ffc_247_n_spl_0,
    ffc_247_n_spl_
  );


  buf

  (
    g693_n_spl_,
    g693_n
  );


  buf

  (
    ffc_247_p_spl_,
    ffc_247_p
  );


  buf

  (
    ffc_247_p_spl_0,
    ffc_247_p_spl_
  );


  buf

  (
    ffc_248_p_spl_,
    ffc_248_p
  );


  buf

  (
    ffc_248_p_spl_0,
    ffc_248_p_spl_
  );


  buf

  (
    ffc_248_p_spl_1,
    ffc_248_p_spl_
  );


  buf

  (
    ffc_314_p_spl_,
    ffc_314_p
  );


  buf

  (
    ffc_314_p_spl_0,
    ffc_314_p_spl_
  );


  buf

  (
    ffc_248_n_spl_,
    ffc_248_n
  );


  buf

  (
    ffc_248_n_spl_0,
    ffc_248_n_spl_
  );


  buf

  (
    ffc_314_n_spl_,
    ffc_314_n
  );


  buf

  (
    g658_p_spl_,
    g658_p
  );


  buf

  (
    g658_p_spl_0,
    g658_p_spl_
  );


  buf

  (
    g658_p_spl_1,
    g658_p_spl_
  );


  buf

  (
    g705_n_spl_,
    g705_n
  );


  buf

  (
    ffc_324_n_spl_,
    ffc_324_n
  );


  buf

  (
    ffc_324_n_spl_0,
    ffc_324_n_spl_
  );


  buf

  (
    ffc_324_p_spl_,
    ffc_324_p
  );


  buf

  (
    ffc_324_p_spl_0,
    ffc_324_p_spl_
  );


  buf

  (
    g708_n_spl_,
    g708_n
  );


  buf

  (
    g708_n_spl_0,
    g708_n_spl_
  );


  buf

  (
    g708_p_spl_,
    g708_p
  );


  buf

  (
    g708_p_spl_0,
    g708_p_spl_
  );


  buf

  (
    g711_n_spl_,
    g711_n
  );


  buf

  (
    ffc_148_n_spl_,
    ffc_148_n
  );


  buf

  (
    ffc_127_p_spl_,
    ffc_127_p
  );


  buf

  (
    ffc_127_p_spl_0,
    ffc_127_p_spl_
  );


  buf

  (
    g661_n_spl_,
    g661_n
  );


  buf

  (
    ffc_236_n_spl_,
    ffc_236_n
  );


  buf

  (
    g717_n_spl_,
    g717_n
  );


  buf

  (
    g717_n_spl_0,
    g717_n_spl_
  );


  buf

  (
    g717_n_spl_1,
    g717_n_spl_
  );


  buf

  (
    ffc_150_p_spl_,
    ffc_150_p
  );


  buf

  (
    ffc_150_p_spl_0,
    ffc_150_p_spl_
  );


  buf

  (
    ffc_150_p_spl_1,
    ffc_150_p_spl_
  );


  buf

  (
    g599_p_spl_,
    g599_p
  );


  buf

  (
    ffc_236_p_spl_,
    ffc_236_p
  );


  buf

  (
    ffc_289_p_spl_,
    ffc_289_p
  );


  buf

  (
    ffc_289_n_spl_,
    ffc_289_n
  );


  buf

  (
    g722_n_spl_,
    g722_n
  );


  buf

  (
    g724_n_spl_,
    g724_n
  );


  buf

  (
    g722_p_spl_,
    g722_p
  );


  buf

  (
    g722_p_spl_0,
    g722_p_spl_
  );


  buf

  (
    g724_p_spl_,
    g724_p
  );


  buf

  (
    ffc_120_n_spl_,
    ffc_120_n
  );


  buf

  (
    ffc_264_n_spl_,
    ffc_264_n
  );


  buf

  (
    ffc_120_p_spl_,
    ffc_120_p
  );


  buf

  (
    ffc_264_p_spl_,
    ffc_264_p
  );


  buf

  (
    g553_n_spl_,
    g553_n
  );


  buf

  (
    g731_n_spl_,
    g731_n
  );


  buf

  (
    g553_p_spl_,
    g553_p
  );


  buf

  (
    g553_p_spl_0,
    g553_p_spl_
  );


  buf

  (
    g731_p_spl_,
    g731_p
  );


  buf

  (
    g730_p_spl_,
    g730_p
  );


  buf

  (
    g730_p_spl_0,
    g730_p_spl_
  );


  buf

  (
    g730_p_spl_1,
    g730_p_spl_
  );


  buf

  (
    g732_p_spl_,
    g732_p
  );


  buf

  (
    g730_n_spl_,
    g730_n
  );


  buf

  (
    g730_n_spl_0,
    g730_n_spl_
  );


  buf

  (
    g730_n_spl_00,
    g730_n_spl_0
  );


  buf

  (
    g730_n_spl_1,
    g730_n_spl_
  );


  buf

  (
    g732_n_spl_,
    g732_n
  );


  buf

  (
    g727_p_spl_,
    g727_p
  );


  buf

  (
    g735_p_spl_,
    g735_p
  );


  buf

  (
    ffc_171_p_spl_,
    ffc_171_p
  );


  buf

  (
    ffc_171_p_spl_0,
    ffc_171_p_spl_
  );


  buf

  (
    ffc_171_p_spl_1,
    ffc_171_p_spl_
  );


  buf

  (
    g727_n_spl_,
    g727_n
  );


  buf

  (
    g727_n_spl_0,
    g727_n_spl_
  );


  buf

  (
    g735_n_spl_,
    g735_n
  );


  buf

  (
    ffc_70_p_spl_,
    ffc_70_p
  );


  buf

  (
    ffc_70_p_spl_0,
    ffc_70_p_spl_
  );


  buf

  (
    ffc_70_p_spl_00,
    ffc_70_p_spl_0
  );


  buf

  (
    ffc_70_p_spl_01,
    ffc_70_p_spl_0
  );


  buf

  (
    ffc_70_p_spl_1,
    ffc_70_p_spl_
  );


  buf

  (
    ffc_70_p_spl_10,
    ffc_70_p_spl_1
  );


  buf

  (
    ffc_75_n_spl_,
    ffc_75_n
  );


  buf

  (
    ffc_75_n_spl_0,
    ffc_75_n_spl_
  );


  buf

  (
    ffc_75_n_spl_1,
    ffc_75_n_spl_
  );


  buf

  (
    g559_n_spl_,
    g559_n
  );


  buf

  (
    g551_n_spl_,
    g551_n
  );


  buf

  (
    g552_n_spl_,
    g552_n
  );


  buf

  (
    g612_n_spl_,
    g612_n
  );


  buf

  (
    ffc_174_p_spl_,
    ffc_174_p
  );


  buf

  (
    ffc_174_p_spl_0,
    ffc_174_p_spl_
  );


  buf

  (
    ffc_174_p_spl_00,
    ffc_174_p_spl_0
  );


  buf

  (
    ffc_174_p_spl_1,
    ffc_174_p_spl_
  );


  buf

  (
    ffc_159_n_spl_,
    ffc_159_n
  );


  buf

  (
    ffc_159_n_spl_0,
    ffc_159_n_spl_
  );


  buf

  (
    ffc_159_n_spl_1,
    ffc_159_n_spl_
  );


  buf

  (
    ffc_173_p_spl_,
    ffc_173_p
  );


  buf

  (
    ffc_173_p_spl_0,
    ffc_173_p_spl_
  );


  buf

  (
    ffc_173_p_spl_1,
    ffc_173_p_spl_
  );


  buf

  (
    ffc_89_n_spl_,
    ffc_89_n
  );


  buf

  (
    ffc_175_p_spl_,
    ffc_175_p
  );


  buf

  (
    ffc_175_p_spl_0,
    ffc_175_p_spl_
  );


  buf

  (
    ffc_158_p_spl_,
    ffc_158_p
  );


  buf

  (
    ffc_158_p_spl_0,
    ffc_158_p_spl_
  );


  buf

  (
    ffc_158_p_spl_1,
    ffc_158_p_spl_
  );


  buf

  (
    ffc_83_n_spl_,
    ffc_83_n
  );


  buf

  (
    ffc_172_n_spl_,
    ffc_172_n
  );


  buf

  (
    ffc_172_n_spl_0,
    ffc_172_n_spl_
  );


  buf

  (
    g760_p_spl_,
    g760_p
  );


  buf

  (
    ffc_104_p_spl_,
    ffc_104_p
  );


  buf

  (
    ffc_104_p_spl_0,
    ffc_104_p_spl_
  );


  buf

  (
    ffc_73_p_spl_,
    ffc_73_p
  );


  buf

  (
    g771_n_spl_,
    g771_n
  );


  buf

  (
    g562_n_spl_,
    g562_n
  );


  buf

  (
    ffc_75_p_spl_,
    ffc_75_p
  );


  buf

  (
    ffc_72_p_spl_,
    ffc_72_p
  );


  buf

  (
    ffc_74_p_spl_,
    ffc_74_p
  );


  buf

  (
    ffc_74_n_spl_,
    ffc_74_n
  );


  buf

  (
    ffc_172_p_spl_,
    ffc_172_p
  );


  buf

  (
    ffc_172_p_spl_0,
    ffc_172_p_spl_
  );


  buf

  (
    ffc_172_p_spl_00,
    ffc_172_p_spl_0
  );


  buf

  (
    ffc_172_p_spl_1,
    ffc_172_p_spl_
  );


  buf

  (
    ffc_158_n_spl_,
    ffc_158_n
  );


  buf

  (
    ffc_158_n_spl_0,
    ffc_158_n_spl_
  );


  buf

  (
    ffc_158_n_spl_00,
    ffc_158_n_spl_0
  );


  buf

  (
    ffc_158_n_spl_01,
    ffc_158_n_spl_0
  );


  buf

  (
    ffc_158_n_spl_1,
    ffc_158_n_spl_
  );


  buf

  (
    ffc_158_n_spl_10,
    ffc_158_n_spl_1
  );


  buf

  (
    ffc_78_p_spl_,
    ffc_78_p
  );


  buf

  (
    ffc_78_p_spl_0,
    ffc_78_p_spl_
  );


  buf

  (
    ffc_78_p_spl_1,
    ffc_78_p_spl_
  );


  buf

  (
    ffc_204_p_spl_,
    ffc_204_p
  );


  buf

  (
    ffc_174_n_spl_,
    ffc_174_n
  );


  buf

  (
    ffc_174_n_spl_0,
    ffc_174_n_spl_
  );


  buf

  (
    ffc_174_n_spl_00,
    ffc_174_n_spl_0
  );


  buf

  (
    ffc_174_n_spl_000,
    ffc_174_n_spl_00
  );


  buf

  (
    ffc_174_n_spl_01,
    ffc_174_n_spl_0
  );


  buf

  (
    ffc_174_n_spl_1,
    ffc_174_n_spl_
  );


  buf

  (
    ffc_174_n_spl_10,
    ffc_174_n_spl_1
  );


  buf

  (
    ffc_174_n_spl_11,
    ffc_174_n_spl_1
  );


  buf

  (
    ffc_73_n_spl_,
    ffc_73_n
  );


  buf

  (
    ffc_83_p_spl_,
    ffc_83_p
  );


  buf

  (
    ffc_83_p_spl_0,
    ffc_83_p_spl_
  );


  buf

  (
    ffc_173_n_spl_,
    ffc_173_n
  );


  buf

  (
    ffc_173_n_spl_0,
    ffc_173_n_spl_
  );


  buf

  (
    ffc_173_n_spl_00,
    ffc_173_n_spl_0
  );


  buf

  (
    ffc_173_n_spl_01,
    ffc_173_n_spl_0
  );


  buf

  (
    ffc_173_n_spl_1,
    ffc_173_n_spl_
  );


  buf

  (
    ffc_175_n_spl_,
    ffc_175_n
  );


  buf

  (
    ffc_175_n_spl_0,
    ffc_175_n_spl_
  );


  buf

  (
    ffc_175_n_spl_00,
    ffc_175_n_spl_0
  );


  buf

  (
    ffc_175_n_spl_01,
    ffc_175_n_spl_0
  );


  buf

  (
    ffc_175_n_spl_1,
    ffc_175_n_spl_
  );


  buf

  (
    ffc_175_n_spl_10,
    ffc_175_n_spl_1
  );


  buf

  (
    ffc_89_p_spl_,
    ffc_89_p
  );


  buf

  (
    ffc_159_p_spl_,
    ffc_159_p
  );


  buf

  (
    ffc_159_p_spl_0,
    ffc_159_p_spl_
  );


  buf

  (
    ffc_159_p_spl_00,
    ffc_159_p_spl_0
  );


  buf

  (
    ffc_159_p_spl_01,
    ffc_159_p_spl_0
  );


  buf

  (
    ffc_159_p_spl_1,
    ffc_159_p_spl_
  );


  buf

  (
    ffc_159_p_spl_10,
    ffc_159_p_spl_1
  );


  buf

  (
    ffc_112_p_spl_,
    ffc_112_p
  );


  buf

  (
    ffc_112_p_spl_0,
    ffc_112_p_spl_
  );


  buf

  (
    g849_p_spl_,
    g849_p
  );


  buf

  (
    g848_n_spl_,
    g848_n
  );


  buf

  (
    ffc_113_p_spl_,
    ffc_113_p
  );


  buf

  (
    ffc_113_p_spl_0,
    ffc_113_p_spl_
  );


  buf

  (
    ffc_262_n_spl_,
    ffc_262_n
  );


  buf

  (
    ffc_103_n_spl_,
    ffc_103_n
  );


  buf

  (
    ffc_122_p_spl_,
    ffc_122_p
  );


  buf

  (
    ffc_122_n_spl_,
    ffc_122_n
  );


  buf

  (
    ffc_119_n_spl_,
    ffc_119_n
  );


  buf

  (
    g870_n_spl_,
    g870_n
  );


  buf

  (
    ffc_119_p_spl_,
    ffc_119_p
  );


  buf

  (
    g870_p_spl_,
    g870_p
  );


  buf

  (
    g873_n_spl_,
    g873_n
  );


  buf

  (
    g873_n_spl_0,
    g873_n_spl_
  );


  buf

  (
    g687_n_spl_,
    g687_n
  );


  buf

  (
    g878_n_spl_,
    g878_n
  );


  buf

  (
    g877_p_spl_,
    g877_p
  );


  buf

  (
    g877_p_spl_0,
    g877_p_spl_
  );


  buf

  (
    g883_n_spl_,
    g883_n
  );


  buf

  (
    g883_n_spl_0,
    g883_n_spl_
  );


  buf

  (
    g883_n_spl_1,
    g883_n_spl_
  );


  buf

  (
    g884_n_spl_,
    g884_n
  );


  buf

  (
    g885_n_spl_,
    g885_n
  );


  buf

  (
    ffc_171_n_spl_,
    ffc_171_n
  );


  buf

  (
    ffc_171_n_spl_0,
    ffc_171_n_spl_
  );


  buf

  (
    g888_n_spl_,
    g888_n
  );


  buf

  (
    g577_n_spl_,
    g577_n
  );


  buf

  (
    g577_n_spl_0,
    g577_n_spl_
  );


  buf

  (
    g656_n_spl_,
    g656_n
  );


  buf

  (
    ffc_252_p_spl_,
    ffc_252_p
  );


  buf

  (
    ffc_130_p_spl_,
    ffc_130_p
  );


  buf

  (
    ffc_163_p_spl_,
    ffc_163_p
  );


  buf

  (
    ffc_163_p_spl_0,
    ffc_163_p_spl_
  );


  buf

  (
    g960_p_spl_,
    g960_p
  );


  buf

  (
    g873_p_spl_,
    g873_p
  );


  buf

  (
    g960_n_spl_,
    g960_n
  );


  buf

  (
    g621_n_spl_,
    g621_n
  );


  buf

  (
    g621_n_spl_0,
    g621_n_spl_
  );


  buf

  (
    g645_n_spl_,
    g645_n
  );


  buf

  (
    g645_n_spl_0,
    g645_n_spl_
  );


  buf

  (
    ffc_251_p_spl_,
    ffc_251_p
  );


  buf

  (
    ffc_326_p_spl_,
    ffc_326_p
  );


  buf

  (
    g990_n_spl_,
    g990_n
  );


  buf

  (
    g659_n_spl_,
    g659_n
  );


  buf

  (
    g659_n_spl_0,
    g659_n_spl_
  );


  buf

  (
    g659_n_spl_00,
    g659_n_spl_0
  );


  buf

  (
    g659_n_spl_01,
    g659_n_spl_0
  );


  buf

  (
    g659_n_spl_1,
    g659_n_spl_
  );


  buf

  (
    g659_n_spl_10,
    g659_n_spl_1
  );


  buf

  (
    g705_p_spl_,
    g705_p
  );


  buf

  (
    g676_n_spl_,
    g676_n
  );


  buf

  (
    g707_n_spl_,
    g707_n
  );


  buf

  (
    g711_p_spl_,
    g711_p
  );


  buf

  (
    g684_n_spl_,
    g684_n
  );


  buf

  (
    g713_n_spl_,
    g713_n
  );


  buf

  (
    ffc_126_p_spl_,
    ffc_126_p
  );


  buf

  (
    ffc_129_p_spl_,
    ffc_129_p
  );


  buf

  (
    ffc_162_p_spl_,
    ffc_162_p
  );


  buf

  (
    ffc_132_p_spl_,
    ffc_132_p
  );


  buf

  (
    ffc_132_n_spl_,
    ffc_132_n
  );


  buf

  (
    g581_n_spl_,
    g581_n
  );


  buf

  (
    g581_n_spl_0,
    g581_n_spl_
  );


  buf

  (
    g581_n_spl_00,
    g581_n_spl_0
  );


  buf

  (
    g581_n_spl_01,
    g581_n_spl_0
  );


  buf

  (
    g581_n_spl_1,
    g581_n_spl_
  );


  buf

  (
    ffc_145_p_spl_,
    ffc_145_p
  );


  buf

  (
    ffc_15_p_spl_,
    ffc_15_p
  );


  buf

  (
    ffc_15_p_spl_0,
    ffc_15_p_spl_
  );


  buf

  (
    g583_n_spl_,
    g583_n
  );


  buf

  (
    g583_n_spl_0,
    g583_n_spl_
  );


  buf

  (
    g583_n_spl_00,
    g583_n_spl_0
  );


  buf

  (
    g583_n_spl_01,
    g583_n_spl_0
  );


  buf

  (
    g583_n_spl_1,
    g583_n_spl_
  );


  buf

  (
    g890_n_spl_,
    g890_n
  );


  buf

  (
    g1013_p_spl_,
    g1013_p
  );


  buf

  (
    g1013_p_spl_0,
    g1013_p_spl_
  );


  buf

  (
    g886_n_spl_,
    g886_n
  );


  buf

  (
    g886_n_spl_0,
    g886_n_spl_
  );


  buf

  (
    ffc_13_p_spl_,
    ffc_13_p
  );


  buf

  (
    ffc_48_n_spl_,
    ffc_48_n
  );


  buf

  (
    g976_n_spl_,
    g976_n
  );


  buf

  (
    ffc_39_p_spl_,
    ffc_39_p
  );


  buf

  (
    ffc_37_p_spl_,
    ffc_37_p
  );


  buf

  (
    g1020_n_spl_,
    g1020_n
  );


  buf

  (
    ffc_48_p_spl_,
    ffc_48_p
  );


  buf

  (
    g590_p_spl_,
    g590_p
  );


  buf

  (
    g577_p_spl_,
    g577_p
  );


  buf

  (
    g577_p_spl_0,
    g577_p_spl_
  );


  buf

  (
    g1026_p_spl_,
    g1026_p
  );


  buf

  (
    g656_p_spl_,
    g656_p
  );


  buf

  (
    g656_p_spl_0,
    g656_p_spl_
  );


  buf

  (
    g1025_n_spl_,
    g1025_n
  );


  buf

  (
    g1025_n_spl_0,
    g1025_n_spl_
  );


  buf

  (
    g1031_n_spl_,
    g1031_n
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G1_p_spl_0,
    G1_p_spl_
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    g662_n_spl_,
    g662_n
  );


  buf

  (
    g664_n_spl_,
    g664_n
  );


  buf

  (
    g716_p_spl_,
    g716_p
  );


  buf

  (
    ffc_196_p_spl_,
    ffc_196_p
  );


  buf

  (
    ffc_196_p_spl_0,
    ffc_196_p_spl_
  );


  buf

  (
    g591_n_spl_,
    g591_n
  );


  buf

  (
    ffc_21_p_spl_,
    ffc_21_p
  );


  buf

  (
    ffc_21_p_spl_0,
    ffc_21_p_spl_
  );


  buf

  (
    g598_n_spl_,
    g598_n
  );


  buf

  (
    g598_n_spl_0,
    g598_n_spl_
  );


  buf

  (
    g598_n_spl_1,
    g598_n_spl_
  );


  buf

  (
    ffc_137_p_spl_,
    ffc_137_p
  );


  buf

  (
    g719_n_spl_,
    g719_n
  );


  buf

  (
    ffc_135_p_spl_,
    ffc_135_p
  );


  buf

  (
    ffc_135_p_spl_0,
    ffc_135_p_spl_
  );


  buf

  (
    g720_n_spl_,
    g720_n
  );


  buf

  (
    g950_n_spl_,
    g950_n
  );


  buf

  (
    g595_n_spl_,
    g595_n
  );


  buf

  (
    g595_n_spl_0,
    g595_n_spl_
  );


  buf

  (
    g875_n_spl_,
    g875_n
  );


  buf

  (
    g972_n_spl_,
    g972_n
  );


  buf

  (
    g876_n_spl_,
    g876_n
  );


  buf

  (
    ffc_313_p_spl_,
    ffc_313_p
  );


  buf

  (
    ffc_313_p_spl_0,
    ffc_313_p_spl_
  );


  buf

  (
    g1082_p_spl_,
    g1082_p
  );


  buf

  (
    g1082_p_spl_0,
    g1082_p_spl_
  );


  buf

  (
    g1082_p_spl_1,
    g1082_p_spl_
  );


  buf

  (
    g666_p_spl_,
    g666_p
  );


  buf

  (
    g1086_n_spl_,
    g1086_n
  );


  buf

  (
    g1088_p_spl_,
    g1088_p
  );


  buf

  (
    g665_n_spl_,
    g665_n
  );


  buf

  (
    ffc_352_p_spl_,
    ffc_352_p
  );


  buf

  (
    ffc_302_p_spl_,
    ffc_302_p
  );


  buf

  (
    ffc_304_n_spl_,
    ffc_304_n
  );


  buf

  (
    ffc_304_n_spl_0,
    ffc_304_n_spl_
  );


  buf

  (
    ffc_304_p_spl_,
    ffc_304_p
  );


  buf

  (
    ffc_304_p_spl_0,
    ffc_304_p_spl_
  );


  buf

  (
    g1108_n_spl_,
    g1108_n
  );


  buf

  (
    g663_p_spl_,
    g663_p
  );


  buf

  (
    g660_p_spl_,
    g660_p
  );


  buf

  (
    g990_p_spl_,
    g990_p
  );


  buf

  (
    g701_n_spl_,
    g701_n
  );


  buf

  (
    g992_n_spl_,
    g992_n
  );


  buf

  (
    g995_p_spl_,
    g995_p
  );


  buf

  (
    g998_p_spl_,
    g998_p
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_00,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_000,
    G4_p_spl_00
  );


  buf

  (
    G4_p_spl_001,
    G4_p_spl_00
  );


  buf

  (
    G4_p_spl_01,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_10,
    G4_p_spl_1
  );


  buf

  (
    G4_p_spl_11,
    G4_p_spl_1
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_1,
    G12_p_spl_
  );


  buf

  (
    G13_p_spl_,
    G13_p
  );


  buf

  (
    G13_p_spl_0,
    G13_p_spl_
  );


  buf

  (
    ffc_22_p_spl_,
    ffc_22_p
  );


  buf

  (
    g667_n_spl_,
    g667_n
  );


  buf

  (
    ffc_23_p_spl_,
    ffc_23_p
  );


  buf

  (
    g686_p_spl_,
    g686_p
  );


  buf

  (
    ffc_351_p_spl_,
    ffc_351_p
  );


  buf

  (
    ffc_351_p_spl_0,
    ffc_351_p_spl_
  );


  buf

  (
    ffc_243_p_spl_,
    ffc_243_p
  );


  buf

  (
    ffc_243_p_spl_0,
    ffc_243_p_spl_
  );


  buf

  (
    ffc_243_p_spl_00,
    ffc_243_p_spl_0
  );


  buf

  (
    ffc_243_p_spl_1,
    ffc_243_p_spl_
  );


  buf

  (
    ffc_27_p_spl_,
    ffc_27_p
  );


  buf

  (
    ffc_243_n_spl_,
    ffc_243_n
  );


  buf

  (
    ffc_243_n_spl_0,
    ffc_243_n_spl_
  );


  buf

  (
    ffc_243_n_spl_1,
    ffc_243_n_spl_
  );


  buf

  (
    g1108_p_spl_,
    g1108_p
  );


  buf

  (
    ffc_359_p_spl_,
    ffc_359_p
  );


  buf

  (
    g691_p_spl_,
    g691_p
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G3_p_spl_0,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_00,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_1,
    G3_p_spl_
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    G4_n_spl_0,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_00,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_1,
    G4_n_spl_
  );


  buf

  (
    G3_n_spl_,
    G3_n
  );


  buf

  (
    g1034_n_spl_,
    g1034_n
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G5_p_spl_0,
    G5_p_spl_
  );


  buf

  (
    ffc_325_n_spl_,
    ffc_325_n
  );


  buf

  (
    ffc_359_n_spl_,
    ffc_359_n
  );


  buf

  (
    g691_n_spl_,
    g691_n
  );


  buf

  (
    g658_n_spl_,
    g658_n
  );


  buf

  (
    g658_n_spl_0,
    g658_n_spl_
  );


  buf

  (
    g1179_p_spl_,
    g1179_p
  );


  buf

  (
    g1085_n_spl_,
    g1085_n
  );


  buf

  (
    g1085_n_spl_0,
    g1085_n_spl_
  );


  buf

  (
    g1190_p_spl_,
    g1190_p
  );


  buf

  (
    g1098_n_spl_,
    g1098_n
  );


  buf

  (
    g1098_n_spl_0,
    g1098_n_spl_
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    g1197_n_spl_,
    g1197_n
  );


  buf

  (
    g1035_n_spl_,
    g1035_n
  );


  buf

  (
    g1035_n_spl_0,
    g1035_n_spl_
  );


  buf

  (
    g1074_n_spl_,
    g1074_n
  );


  buf

  (
    g985_n_spl_,
    g985_n
  );


  buf

  (
    g1110_n_spl_,
    g1110_n
  );


  buf

  (
    g1120_p_spl_,
    g1120_p
  );


  buf

  (
    g1121_p_spl_,
    g1121_p
  );


  buf

  (
    G13_n_spl_,
    G13_n
  );


  buf

  (
    g1124_n_spl_,
    g1124_n
  );


  buf

  (
    g1123_n_spl_,
    g1123_n
  );


  buf

  (
    g1208_p_spl_,
    g1208_p
  );


  buf

  (
    G41_p_spl_,
    G41_p
  );


  buf

  (
    g1162_n_spl_,
    g1162_n
  );


  buf

  (
    g1162_n_spl_0,
    g1162_n_spl_
  );


  buf

  (
    g1162_n_spl_1,
    g1162_n_spl_
  );


  buf

  (
    G34_n_spl_,
    G34_n
  );


  buf

  (
    g1122_n_spl_,
    g1122_n
  );


  buf

  (
    g1122_n_spl_0,
    g1122_n_spl_
  );


  buf

  (
    g1122_n_spl_1,
    g1122_n_spl_
  );


  buf

  (
    g1164_p_spl_,
    g1164_p
  );


  buf

  (
    G35_p_spl_,
    G35_p
  );


  buf

  (
    G35_p_spl_0,
    G35_p_spl_
  );


  buf

  (
    g1201_n_spl_,
    g1201_n
  );


  buf

  (
    g1163_n_spl_,
    g1163_n
  );


  buf

  (
    g1200_p_spl_,
    g1200_p
  );


  buf

  (
    G40_p_spl_,
    G40_p
  );


  buf

  (
    G33_p_spl_,
    G33_p
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G34_p_spl_,
    G34_p
  );


  buf

  (
    g1210_n_spl_,
    g1210_n
  );


endmodule
