// Benchmark "c1908" written by ABC on Sun Oct 29 22:18:02 2023

module c1908 ( 
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33,
    G1884, G1885, G1886, G1887, G1888, G1889, G1890, G1891, G1892, G1893,
    G1894, G1895, G1896, G1897, G1898, G1899, G1900, G1901, G1902, G1903,
    G1904, G1905, G1906, G1907, G1908  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33;
  output G1884, G1885, G1886, G1887, G1888, G1889, G1890, G1891, G1892, G1893,
    G1894, G1895, G1896, G1897, G1898, G1899, G1900, G1901, G1902, G1903,
    G1904, G1905, G1906, G1907, G1908;
  wire new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n237_, new_n238_, new_n240_,
    new_n241_, new_n243_, new_n244_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n253_, new_n254_, new_n256_,
    new_n257_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n265_, new_n266_, new_n268_, new_n269_, new_n271_, new_n272_,
    new_n274_, new_n275_, new_n276_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n285_, new_n286_, new_n288_,
    new_n289_, new_n291_, new_n292_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n314_, new_n315_, new_n316_, new_n318_,
    new_n319_, new_n320_, new_n322_, new_n323_, new_n324_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n347_, new_n348_, new_n349_;
  nor1 g000(.dina(G29), .dinb(G33), .dout(new_n59_));
  anb2 g001(.dina(G23), .dinb(G24), .dout(new_n60_));
  anb2 g002(.dina(G31), .dinb(new_n60_), .dout(new_n61_));
  nab2 g003(.dina(new_n59_), .dinb(new_n61_), .dout(new_n62_));
  and2 g004(.dina(G32), .dinb(G33), .dout(new_n63_));
  anb1 g005(.dina(new_n60_), .dinb(new_n63_), .dout(new_n64_));
  anb1 g006(.dina(new_n62_), .dinb(new_n64_), .dout(new_n65_));
  nor1 g007(.dina(G23), .dinb(G31), .dout(new_n66_));
  anb1 g008(.dina(G20), .dinb(new_n66_), .dout(new_n67_));
  anb2 g009(.dina(G33), .dinb(G22), .dout(new_n68_));
  nor1 g010(.dina(G4), .dinb(G14), .dout(new_n69_));
  nor2 g011(.dina(G4), .dinb(G14), .dout(new_n70_));
  anb2 g012(.dina(new_n69_), .dinb(new_n70_), .dout(new_n71_));
  anb2 g013(.dina(new_n68_), .dinb(new_n71_), .dout(new_n72_));
  anb1 g014(.dina(new_n68_), .dinb(new_n71_), .dout(new_n73_));
  anb1 g015(.dina(new_n72_), .dinb(new_n73_), .dout(new_n74_));
  and2 g016(.dina(G12), .dinb(G13), .dout(new_n75_));
  and1 g017(.dina(G12), .dinb(G13), .dout(new_n76_));
  anb1 g018(.dina(new_n75_), .dinb(new_n76_), .dout(new_n77_));
  anb1 g019(.dina(G11), .dinb(new_n77_), .dout(new_n78_));
  anb2 g020(.dina(G11), .dinb(new_n77_), .dout(new_n79_));
  anb2 g021(.dina(new_n78_), .dinb(new_n79_), .dout(new_n80_));
  anb2 g022(.dina(G15), .dinb(G10), .dout(new_n81_));
  anb1 g023(.dina(G15), .dinb(G10), .dout(new_n82_));
  anb1 g024(.dina(new_n81_), .dinb(new_n82_), .dout(new_n83_));
  anb2 g025(.dina(new_n83_), .dinb(G16), .dout(new_n84_));
  anb1 g026(.dina(new_n83_), .dinb(G16), .dout(new_n85_));
  anb1 g027(.dina(new_n84_), .dinb(new_n85_), .dout(new_n86_));
  anb1 g028(.dina(new_n80_), .dinb(new_n86_), .dout(new_n87_));
  anb2 g029(.dina(new_n80_), .dinb(new_n86_), .dout(new_n88_));
  anb2 g030(.dina(new_n87_), .dinb(new_n88_), .dout(new_n89_));
  and2 g031(.dina(G2), .dinb(G3), .dout(new_n90_));
  and1 g032(.dina(G2), .dinb(G3), .dout(new_n91_));
  anb1 g033(.dina(new_n90_), .dinb(new_n91_), .dout(new_n92_));
  anb1 g034(.dina(G1), .dinb(new_n92_), .dout(new_n93_));
  anb2 g035(.dina(G1), .dinb(new_n92_), .dout(new_n94_));
  anb2 g036(.dina(new_n93_), .dinb(new_n94_), .dout(new_n95_));
  anb2 g037(.dina(new_n89_), .dinb(new_n95_), .dout(new_n96_));
  anb1 g038(.dina(new_n89_), .dinb(new_n95_), .dout(new_n97_));
  anb1 g039(.dina(new_n96_), .dinb(new_n97_), .dout(new_n98_));
  anb2 g040(.dina(new_n74_), .dinb(new_n98_), .dout(new_n99_));
  anb1 g041(.dina(new_n74_), .dinb(new_n98_), .dout(new_n100_));
  anb1 g042(.dina(new_n99_), .dinb(new_n100_), .dout(new_n101_));
  nor1 g043(.dina(G31), .dinb(new_n101_), .dout(new_n102_));
  anb2 g044(.dina(G25), .dinb(new_n102_), .dout(new_n103_));
  anb1 g045(.dina(G25), .dinb(new_n102_), .dout(new_n104_));
  anb1 g046(.dina(new_n103_), .dinb(new_n104_), .dout(new_n105_));
  anb1 g047(.dina(new_n67_), .dinb(new_n105_), .dout(new_n106_));
  anb1 g048(.dina(G18), .dinb(G24), .dout(new_n107_));
  anb1 g049(.dina(new_n107_), .dinb(G33), .dout(new_n108_));
  anb1 g050(.dina(G15), .dinb(new_n108_), .dout(new_n109_));
  anb2 g051(.dina(G15), .dinb(new_n108_), .dout(new_n110_));
  anb2 g052(.dina(new_n109_), .dinb(new_n110_), .dout(new_n111_));
  anb2 g053(.dina(G11), .dinb(new_n111_), .dout(new_n112_));
  anb1 g054(.dina(G11), .dinb(new_n111_), .dout(new_n113_));
  anb1 g055(.dina(new_n112_), .dinb(new_n113_), .dout(new_n114_));
  and2 g056(.dina(G9), .dinb(G14), .dout(new_n115_));
  and1 g057(.dina(G9), .dinb(G14), .dout(new_n116_));
  anb1 g058(.dina(new_n115_), .dinb(new_n116_), .dout(new_n117_));
  anb2 g059(.dina(new_n117_), .dinb(G16), .dout(new_n118_));
  anb1 g060(.dina(new_n117_), .dinb(G16), .dout(new_n119_));
  anb1 g061(.dina(new_n118_), .dinb(new_n119_), .dout(new_n120_));
  anb1 g062(.dina(new_n114_), .dinb(new_n120_), .dout(new_n121_));
  anb2 g063(.dina(new_n114_), .dinb(new_n120_), .dout(new_n122_));
  anb2 g064(.dina(new_n121_), .dinb(new_n122_), .dout(new_n123_));
  anb1 g065(.dina(G5), .dinb(G8), .dout(new_n124_));
  anb2 g066(.dina(G5), .dinb(G8), .dout(new_n125_));
  anb2 g067(.dina(new_n124_), .dinb(new_n125_), .dout(new_n126_));
  nab1 g068(.dina(G2), .dinb(new_n126_), .dout(new_n127_));
  nab2 g069(.dina(G2), .dinb(new_n126_), .dout(new_n128_));
  anb2 g070(.dina(new_n127_), .dinb(new_n128_), .dout(new_n129_));
  anb1 g071(.dina(new_n123_), .dinb(new_n129_), .dout(new_n130_));
  anb2 g072(.dina(new_n123_), .dinb(new_n129_), .dout(new_n131_));
  anb2 g073(.dina(new_n130_), .dinb(new_n131_), .dout(new_n132_));
  nab1 g074(.dina(G31), .dinb(new_n132_), .dout(new_n133_));
  anb2 g075(.dina(G27), .dinb(new_n133_), .dout(new_n134_));
  anb1 g076(.dina(G6), .dinb(G8), .dout(new_n135_));
  anb2 g077(.dina(G6), .dinb(G8), .dout(new_n136_));
  anb2 g078(.dina(new_n135_), .dinb(new_n136_), .dout(new_n137_));
  nab1 g079(.dina(G3), .dinb(new_n137_), .dout(new_n138_));
  nab2 g080(.dina(G3), .dinb(new_n137_), .dout(new_n139_));
  anb2 g081(.dina(new_n138_), .dinb(new_n139_), .dout(new_n140_));
  nor1 g082(.dina(G12), .dinb(new_n83_), .dout(new_n141_));
  nor2 g083(.dina(G12), .dinb(new_n83_), .dout(new_n142_));
  anb2 g084(.dina(new_n141_), .dinb(new_n142_), .dout(new_n143_));
  anb1 g085(.dina(new_n140_), .dinb(new_n143_), .dout(new_n144_));
  anb2 g086(.dina(new_n140_), .dinb(new_n143_), .dout(new_n145_));
  anb2 g087(.dina(new_n144_), .dinb(new_n145_), .dout(new_n146_));
  anb1 g088(.dina(G19), .dinb(G23), .dout(new_n147_));
  anb1 g089(.dina(new_n147_), .dinb(G33), .dout(new_n148_));
  anb1 g090(.dina(new_n146_), .dinb(new_n148_), .dout(new_n149_));
  anb2 g091(.dina(new_n146_), .dinb(new_n148_), .dout(new_n150_));
  anb2 g092(.dina(new_n149_), .dinb(new_n150_), .dout(new_n151_));
  nab1 g093(.dina(G31), .dinb(new_n151_), .dout(new_n152_));
  anb1 g094(.dina(new_n152_), .dinb(G28), .dout(new_n153_));
  anb2 g095(.dina(new_n152_), .dinb(G28), .dout(new_n154_));
  anb2 g096(.dina(new_n153_), .dinb(new_n154_), .dout(new_n155_));
  anb1 g097(.dina(G7), .dinb(G10), .dout(new_n156_));
  anb2 g098(.dina(G7), .dinb(G10), .dout(new_n157_));
  anb2 g099(.dina(new_n156_), .dinb(new_n157_), .dout(new_n158_));
  anb2 g100(.dina(G4), .dinb(new_n158_), .dout(new_n159_));
  anb1 g101(.dina(G4), .dinb(new_n158_), .dout(new_n160_));
  anb1 g102(.dina(new_n159_), .dinb(new_n160_), .dout(new_n161_));
  anb1 g103(.dina(new_n120_), .dinb(new_n161_), .dout(new_n162_));
  anb2 g104(.dina(new_n120_), .dinb(new_n161_), .dout(new_n163_));
  anb2 g105(.dina(new_n162_), .dinb(new_n163_), .dout(new_n164_));
  anb1 g106(.dina(G20), .dinb(G23), .dout(new_n165_));
  anb1 g107(.dina(new_n165_), .dinb(G33), .dout(new_n166_));
  anb2 g108(.dina(G13), .dinb(new_n166_), .dout(new_n167_));
  anb1 g109(.dina(G13), .dinb(new_n166_), .dout(new_n168_));
  anb1 g110(.dina(new_n167_), .dinb(new_n168_), .dout(new_n169_));
  anb1 g111(.dina(new_n164_), .dinb(new_n169_), .dout(new_n170_));
  anb2 g112(.dina(new_n164_), .dinb(new_n169_), .dout(new_n171_));
  anb2 g113(.dina(new_n170_), .dinb(new_n171_), .dout(new_n172_));
  nab1 g114(.dina(G31), .dinb(new_n172_), .dout(new_n173_));
  anb1 g115(.dina(G19), .dinb(new_n66_), .dout(new_n174_));
  anb2 g116(.dina(new_n174_), .dinb(new_n173_), .dout(new_n175_));
  anb1 g117(.dina(new_n174_), .dinb(new_n173_), .dout(new_n176_));
  anb1 g118(.dina(new_n175_), .dinb(new_n176_), .dout(new_n177_));
  anb2 g119(.dina(new_n155_), .dinb(new_n177_), .dout(new_n178_));
  anb1 g120(.dina(new_n134_), .dinb(new_n178_), .dout(new_n179_));
  anb1 g121(.dina(G17), .dinb(G24), .dout(new_n180_));
  anb2 g122(.dina(G33), .dinb(new_n180_), .dout(new_n181_));
  nab2 g123(.dina(G1), .dinb(new_n181_), .dout(new_n182_));
  nab1 g124(.dina(G1), .dinb(new_n181_), .dout(new_n183_));
  anb1 g125(.dina(new_n182_), .dinb(new_n183_), .dout(new_n184_));
  and2 g126(.dina(G6), .dinb(G7), .dout(new_n185_));
  and1 g127(.dina(G6), .dinb(G7), .dout(new_n186_));
  anb1 g128(.dina(new_n185_), .dinb(new_n186_), .dout(new_n187_));
  anb1 g129(.dina(G5), .dinb(new_n187_), .dout(new_n188_));
  anb2 g130(.dina(G5), .dinb(new_n187_), .dout(new_n189_));
  anb2 g131(.dina(new_n188_), .dinb(new_n189_), .dout(new_n190_));
  anb2 g132(.dina(new_n89_), .dinb(new_n190_), .dout(new_n191_));
  anb1 g133(.dina(new_n89_), .dinb(new_n190_), .dout(new_n192_));
  anb1 g134(.dina(new_n191_), .dinb(new_n192_), .dout(new_n193_));
  anb1 g135(.dina(new_n184_), .dinb(new_n193_), .dout(new_n194_));
  anb2 g136(.dina(new_n184_), .dinb(new_n193_), .dout(new_n195_));
  anb2 g137(.dina(new_n194_), .dinb(new_n195_), .dout(new_n196_));
  nab1 g138(.dina(G31), .dinb(new_n196_), .dout(new_n197_));
  anb1 g139(.dina(G26), .dinb(new_n197_), .dout(new_n198_));
  anb2 g140(.dina(G26), .dinb(new_n197_), .dout(new_n199_));
  anb1 g141(.dina(G27), .dinb(new_n133_), .dout(new_n200_));
  anb1 g142(.dina(new_n199_), .dinb(new_n200_), .dout(new_n201_));
  anb2 g143(.dina(new_n198_), .dinb(new_n201_), .dout(new_n202_));
  anb1 g144(.dina(new_n179_), .dinb(new_n202_), .dout(new_n203_));
  nor1 g145(.dina(G24), .dinb(G31), .dout(new_n204_));
  anb2 g146(.dina(new_n204_), .dinb(G18), .dout(new_n205_));
  anb2 g147(.dina(G33), .dinb(G21), .dout(new_n206_));
  anb1 g148(.dina(G9), .dinb(new_n86_), .dout(new_n207_));
  anb2 g149(.dina(G9), .dinb(new_n86_), .dout(new_n208_));
  anb2 g150(.dina(new_n207_), .dinb(new_n208_), .dout(new_n209_));
  anb2 g151(.dina(new_n206_), .dinb(new_n209_), .dout(new_n210_));
  anb1 g152(.dina(new_n206_), .dinb(new_n209_), .dout(new_n211_));
  anb1 g153(.dina(new_n210_), .dinb(new_n211_), .dout(new_n212_));
  and1 g154(.dina(new_n95_), .dinb(new_n190_), .dout(new_n213_));
  and2 g155(.dina(new_n95_), .dinb(new_n190_), .dout(new_n214_));
  nab1 g156(.dina(new_n213_), .dinb(new_n214_), .dout(new_n215_));
  anb2 g157(.dina(G8), .dinb(G4), .dout(new_n216_));
  anb1 g158(.dina(G8), .dinb(G4), .dout(new_n217_));
  anb1 g159(.dina(new_n216_), .dinb(new_n217_), .dout(new_n218_));
  anb2 g160(.dina(new_n215_), .dinb(new_n218_), .dout(new_n219_));
  anb1 g161(.dina(new_n215_), .dinb(new_n218_), .dout(new_n220_));
  anb1 g162(.dina(new_n219_), .dinb(new_n220_), .dout(new_n221_));
  anb1 g163(.dina(new_n212_), .dinb(new_n221_), .dout(new_n222_));
  anb2 g164(.dina(new_n212_), .dinb(new_n221_), .dout(new_n223_));
  anb2 g165(.dina(new_n222_), .dinb(new_n223_), .dout(new_n224_));
  nor1 g166(.dina(G31), .dinb(new_n224_), .dout(new_n225_));
  anb1 g167(.dina(G17), .dinb(new_n204_), .dout(new_n226_));
  anb1 g168(.dina(new_n225_), .dinb(new_n226_), .dout(new_n227_));
  anb2 g169(.dina(new_n225_), .dinb(new_n226_), .dout(new_n228_));
  anb2 g170(.dina(new_n227_), .dinb(new_n228_), .dout(new_n229_));
  anb1 g171(.dina(new_n229_), .dinb(new_n205_), .dout(new_n230_));
  anb1 g172(.dina(new_n203_), .dinb(new_n230_), .dout(new_n231_));
  anb1 g173(.dina(new_n231_), .dinb(new_n106_), .dout(new_n232_));
  anb2 g174(.dina(new_n65_), .dinb(new_n232_), .dout(new_n233_));
  nab1 g175(.dina(G1), .dinb(new_n233_), .dout(new_n234_));
  nab2 g176(.dina(G1), .dinb(new_n233_), .dout(new_n235_));
  anb2 g177(.dina(new_n234_), .dinb(new_n235_), .dout(G1884));
  nab1 g178(.dina(G2), .dinb(new_n233_), .dout(new_n237_));
  nab2 g179(.dina(G2), .dinb(new_n233_), .dout(new_n238_));
  anb2 g180(.dina(new_n237_), .dinb(new_n238_), .dout(G1885));
  nab1 g181(.dina(G3), .dinb(new_n233_), .dout(new_n240_));
  nab2 g182(.dina(G3), .dinb(new_n233_), .dout(new_n241_));
  anb2 g183(.dina(new_n240_), .dinb(new_n241_), .dout(G1886));
  nab1 g184(.dina(G4), .dinb(new_n233_), .dout(new_n243_));
  nab2 g185(.dina(G4), .dinb(new_n233_), .dout(new_n244_));
  anb2 g186(.dina(new_n243_), .dinb(new_n244_), .dout(G1887));
  nor1 g187(.dina(G30), .dinb(G33), .dout(new_n246_));
  anb2 g188(.dina(new_n61_), .dinb(new_n246_), .dout(new_n247_));
  anb2 g189(.dina(new_n64_), .dinb(new_n247_), .dout(new_n248_));
  nor2 g190(.dina(new_n232_), .dinb(new_n248_), .dout(new_n249_));
  nab1 g191(.dina(G10), .dinb(new_n249_), .dout(new_n250_));
  nab2 g192(.dina(G10), .dinb(new_n249_), .dout(new_n251_));
  anb2 g193(.dina(new_n250_), .dinb(new_n251_), .dout(G1888));
  nab1 g194(.dina(G15), .dinb(new_n249_), .dout(new_n253_));
  nab2 g195(.dina(G15), .dinb(new_n249_), .dout(new_n254_));
  anb2 g196(.dina(new_n253_), .dinb(new_n254_), .dout(G1889));
  nab1 g197(.dina(G16), .dinb(new_n249_), .dout(new_n256_));
  nab2 g198(.dina(G16), .dinb(new_n249_), .dout(new_n257_));
  anb2 g199(.dina(new_n256_), .dinb(new_n257_), .dout(G1890));
  nor2 g200(.dina(new_n67_), .dinb(new_n105_), .dout(new_n259_));
  anb1 g201(.dina(new_n231_), .dinb(new_n259_), .dout(new_n260_));
  anb2 g202(.dina(new_n65_), .dinb(new_n260_), .dout(new_n261_));
  nab1 g203(.dina(G5), .dinb(new_n261_), .dout(new_n262_));
  nab2 g204(.dina(G5), .dinb(new_n261_), .dout(new_n263_));
  anb2 g205(.dina(new_n262_), .dinb(new_n263_), .dout(G1891));
  nab1 g206(.dina(G6), .dinb(new_n261_), .dout(new_n265_));
  nab2 g207(.dina(G6), .dinb(new_n261_), .dout(new_n266_));
  anb2 g208(.dina(new_n265_), .dinb(new_n266_), .dout(G1892));
  nab1 g209(.dina(G7), .dinb(new_n261_), .dout(new_n268_));
  nab2 g210(.dina(G7), .dinb(new_n261_), .dout(new_n269_));
  anb2 g211(.dina(new_n268_), .dinb(new_n269_), .dout(G1893));
  nab1 g212(.dina(G8), .dinb(new_n261_), .dout(new_n271_));
  nab2 g213(.dina(G8), .dinb(new_n261_), .dout(new_n272_));
  anb2 g214(.dina(new_n271_), .dinb(new_n272_), .dout(G1894));
  nor2 g215(.dina(new_n248_), .dinb(new_n260_), .dout(new_n274_));
  anb1 g216(.dina(G9), .dinb(new_n274_), .dout(new_n275_));
  anb2 g217(.dina(G9), .dinb(new_n274_), .dout(new_n276_));
  anb2 g218(.dina(new_n275_), .dinb(new_n276_), .dout(G1895));
  anb1 g219(.dina(new_n248_), .dinb(new_n205_), .dout(new_n278_));
  nab1 g220(.dina(new_n229_), .dinb(new_n278_), .dout(new_n279_));
  anb2 g221(.dina(new_n106_), .dinb(new_n279_), .dout(new_n280_));
  anb1 g222(.dina(new_n203_), .dinb(new_n280_), .dout(new_n281_));
  anb2 g223(.dina(new_n281_), .dinb(G11), .dout(new_n282_));
  anb1 g224(.dina(new_n281_), .dinb(G11), .dout(new_n283_));
  anb1 g225(.dina(new_n282_), .dinb(new_n283_), .dout(G1896));
  anb2 g226(.dina(new_n281_), .dinb(G12), .dout(new_n285_));
  anb1 g227(.dina(new_n281_), .dinb(G12), .dout(new_n286_));
  anb1 g228(.dina(new_n285_), .dinb(new_n286_), .dout(G1897));
  anb2 g229(.dina(new_n281_), .dinb(G13), .dout(new_n288_));
  anb1 g230(.dina(new_n281_), .dinb(G13), .dout(new_n289_));
  anb1 g231(.dina(new_n288_), .dinb(new_n289_), .dout(G1898));
  anb2 g232(.dina(new_n281_), .dinb(G14), .dout(new_n291_));
  anb1 g233(.dina(new_n281_), .dinb(G14), .dout(new_n292_));
  anb1 g234(.dina(new_n291_), .dinb(new_n292_), .dout(G1899));
  and1 g235(.dina(new_n233_), .dinb(new_n249_), .dout(new_n294_));
  anb1 g236(.dina(G32), .dinb(new_n294_), .dout(new_n295_));
  anb2 g237(.dina(new_n67_), .dinb(new_n205_), .dout(new_n296_));
  anb1 g238(.dina(new_n105_), .dinb(new_n296_), .dout(new_n297_));
  anb2 g239(.dina(new_n229_), .dinb(new_n297_), .dout(new_n298_));
  nab2 g240(.dina(new_n203_), .dinb(new_n298_), .dout(new_n299_));
  nab1 g241(.dina(G33), .dinb(new_n299_), .dout(new_n300_));
  anb2 g242(.dina(new_n295_), .dinb(new_n300_), .dout(G1900));
  anb1 g243(.dina(new_n226_), .dinb(G31), .dout(new_n302_));
  anb2 g244(.dina(new_n294_), .dinb(new_n302_), .dout(new_n303_));
  anb2 g245(.dina(new_n224_), .dinb(new_n303_), .dout(new_n304_));
  anb1 g246(.dina(new_n224_), .dinb(new_n303_), .dout(new_n305_));
  anb1 g247(.dina(new_n304_), .dinb(new_n305_), .dout(new_n306_));
  anb1 g248(.dina(new_n63_), .dinb(new_n306_), .dout(G1901));
  anb1 g249(.dina(G25), .dinb(G31), .dout(new_n308_));
  anb2 g250(.dina(new_n294_), .dinb(new_n308_), .dout(new_n309_));
  anb2 g251(.dina(new_n101_), .dinb(new_n309_), .dout(new_n310_));
  anb1 g252(.dina(new_n101_), .dinb(new_n309_), .dout(new_n311_));
  anb1 g253(.dina(new_n310_), .dinb(new_n311_), .dout(new_n312_));
  anb1 g254(.dina(new_n63_), .dinb(new_n312_), .dout(G1902));
  anb1 g255(.dina(G27), .dinb(G31), .dout(new_n314_));
  anb1 g256(.dina(new_n314_), .dinb(new_n294_), .dout(new_n315_));
  anb1 g257(.dina(new_n132_), .dinb(new_n315_), .dout(new_n316_));
  anb1 g258(.dina(new_n63_), .dinb(new_n316_), .dout(G1903));
  anb1 g259(.dina(G28), .dinb(G31), .dout(new_n318_));
  anb1 g260(.dina(new_n318_), .dinb(new_n294_), .dout(new_n319_));
  anb1 g261(.dina(new_n151_), .dinb(new_n319_), .dout(new_n320_));
  anb1 g262(.dina(new_n63_), .dinb(new_n320_), .dout(G1904));
  anb1 g263(.dina(new_n174_), .dinb(G31), .dout(new_n322_));
  anb1 g264(.dina(new_n322_), .dinb(new_n294_), .dout(new_n323_));
  anb1 g265(.dina(new_n172_), .dinb(new_n323_), .dout(new_n324_));
  anb1 g266(.dina(new_n63_), .dinb(new_n324_), .dout(G1905));
  nor2 g267(.dina(G21), .dinb(G29), .dout(new_n326_));
  anb2 g268(.dina(G33), .dinb(new_n326_), .dout(new_n327_));
  anb2 g269(.dina(new_n59_), .dinb(new_n221_), .dout(new_n328_));
  anb2 g270(.dina(new_n233_), .dinb(new_n328_), .dout(new_n329_));
  anb1 g271(.dina(new_n233_), .dinb(new_n328_), .dout(new_n330_));
  anb1 g272(.dina(new_n329_), .dinb(new_n330_), .dout(new_n331_));
  anb1 g273(.dina(new_n327_), .dinb(new_n331_), .dout(new_n332_));
  anb2 g274(.dina(new_n327_), .dinb(new_n331_), .dout(new_n333_));
  anb2 g275(.dina(new_n332_), .dinb(new_n333_), .dout(G1906));
  nor2 g276(.dina(G22), .dinb(G30), .dout(new_n335_));
  anb2 g277(.dina(G33), .dinb(new_n335_), .dout(new_n336_));
  anb1 g278(.dina(new_n89_), .dinb(new_n117_), .dout(new_n337_));
  anb2 g279(.dina(new_n89_), .dinb(new_n117_), .dout(new_n338_));
  anb2 g280(.dina(new_n337_), .dinb(new_n338_), .dout(new_n339_));
  anb2 g281(.dina(new_n246_), .dinb(new_n339_), .dout(new_n340_));
  anb2 g282(.dina(new_n249_), .dinb(new_n340_), .dout(new_n341_));
  anb1 g283(.dina(new_n249_), .dinb(new_n340_), .dout(new_n342_));
  anb1 g284(.dina(new_n341_), .dinb(new_n342_), .dout(new_n343_));
  anb1 g285(.dina(new_n336_), .dinb(new_n343_), .dout(new_n344_));
  anb2 g286(.dina(new_n336_), .dinb(new_n343_), .dout(new_n345_));
  anb2 g287(.dina(new_n344_), .dinb(new_n345_), .dout(G1907));
  anb1 g288(.dina(G26), .dinb(G31), .dout(new_n347_));
  anb1 g289(.dina(new_n347_), .dinb(new_n294_), .dout(new_n348_));
  anb1 g290(.dina(new_n196_), .dinb(new_n348_), .dout(new_n349_));
  and1 g291(.dina(new_n63_), .dinb(new_n349_), .dout(G1908));
endmodule


