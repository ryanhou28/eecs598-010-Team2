// Benchmark "mymod" written by ABC on Sun Oct 29 19:32:01 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32,
    G6257, G6258, G6259, G6260, G6261, G6262, G6263, G6264, G6265, G6266,
    G6267, G6268, G6269, G6270, G6271, G6272, G6273, G6274, G6275, G6276,
    G6277, G6278, G6279, G6280, G6281, G6282, G6283, G6284, G6285, G6286,
    G6287, G6288  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32;
  output G6257, G6258, G6259, G6260, G6261, G6262, G6263, G6264, G6265, G6266,
    G6267, G6268, G6269, G6270, G6271, G6272, G6273, G6274, G6275, G6276,
    G6277, G6278, G6279, G6280, G6281, G6282, G6283, G6284, G6285, G6286,
    G6287, G6288;
  reg n2491_lo, n2575_lo, n2587_lo, n2599_lo, n2611_lo, n2623_lo, n2635_lo,
    n2647_lo, n2659_lo, n2671_lo, n2683_lo, n2734_lo, n2746_lo, n2758_lo,
    n2770_lo, n2782_lo, n2785_lo, n2794_lo, n2797_lo, n2806_lo, n2809_lo,
    n2818_lo, n2821_lo, n2830_lo, n2833_lo, n2836_lo, n2839_lo, n2842_lo,
    n2845_lo, n2848_lo, n2851_lo, n2854_lo, n2857_lo, n2860_lo, n2863_lo,
    n4871_o2, n4893_o2, n4938_o2, n5056_o2, n5100_o2, n5122_o2, n5254_o2,
    n5276_o2, n5316_o2, n5434_o2, n5473_o2, n5494_o2, n5620_o2, n5643_o2,
    n5682_o2, n5798_o2, n5839_o2, n5867_o2, n6052_o2, n6087_o2, n6153_o2,
    n6408_o2, n6454_o2, n6509_o2, n6775_o2, n6818_o2, n6892_o2, n5779_o2,
    n5780_o2, n7156_o2, n5792_o2, n7205_o2, n5842_o2, n5863_o2, n7263_o2,
    n5881_o2, n5930_o2, n5959_o2, n5981_o2, n6042_o2, n6075_o2, n6103_o2,
    n7610_o2, n6169_o2, n7665_o2, n6205_o2, n6239_o2, n7788_o2, n6309_o2,
    n6461_o2, n6476_o2, n325_inv, n6545_o2, G578_o2, G5106_o2, n6713_o2,
    G5164_o2, n343_inv, n6810_o2, n6973_o2, n352_inv, n7053_o2, G581_o2,
    G5467_o2, n7231_o2, G5527_o2, n370_inv, n7304_o2, n7530_o2, n379_inv,
    n7653_o2, G584_o2, G5820_o2, n7148_o2, n7149_o2, n7224_o2, n7916_o2,
    G5868_o2, n406_inv, n7280_o2, n7313_o2, n8056_o2, n7323_o2, n7398_o2,
    n7459_o2, n7501_o2, n7518_o2, G563_o2, n7606_o2, n439_inv, n7675_o2,
    G3410_o2, n7722_o2, n7747_o2, n7835_o2, G587_o2, G6046_o2, n7909_o2,
    G566_o2, G6070_o2, n472_inv, n8086_o2, n8093_o2, G3752_o2, n484_inv,
    n8199_o2, n2800_lo_buf_o2, G548_o2, n496_inv, G569_o2, G1761_o2,
    n505_inv, G4101_o2, G551_o2, n514_inv, G4743_o2, G5271_o2, G5790_o2,
    G6122_o2, G2082_o2, n2812_lo_buf_o2, n2668_lo_buf_o2, n2680_lo_buf_o2,
    G572_o2, G6125_o2, n547_inv, n2656_lo_buf_o2, G554_o2, G4452_o2,
    n559_inv, n2644_lo_buf_o2, G2410_o2, n2632_lo_buf_o2, n2620_lo_buf_o2,
    G6131_o2, G4693_o2, G5209_o2, G5741_o2, G6082_o2, G6119_o2,
    n2608_lo_buf_o2, n2596_lo_buf_o2, n2584_lo_buf_o2, n2572_lo_buf_o2,
    n2704_lo_buf_o2, G557_o2, G5936_o2, G5442_o2, G4926_o2, G6134_o2,
    G3929_o2, G4425_o2, G4947_o2, n2764_lo_buf_o2, n634_inv,
    n2560_lo_buf_o2, n2824_lo_buf_o2, G575_o2, G2740_o2, n649_inv,
    n2548_lo_buf_o2, n2536_lo_buf_o2, n2524_lo_buf_o2, G875_o2, G1064_o2,
    G1253_o2, G6140_o2, G5151_o2, G5686_o2, G6061_o2, G4803_o2, G5332_o2,
    G5844_o2, G6114_o2, G4806_o2, G3881_o2, G4370_o2, G4896_o2, G5001_o2,
    G3121_o2, n2512_lo_buf_o2, G4085_o2, G4605_o2, G5118_o2, G4997_o2,
    n2500_lo_buf_o2, n2716_lo_buf_o2, G560_o2, G1895_o2, G3064_o2,
    G3269_o2, G3569_o2, n748_inv, G1196_o2, G1007_o2, G818_o2, G674_o2,
    G5041_o2, G5562_o2, G6005_o2, G5214_o2, G5746_o2, G6087_o2, G6086_o2,
    G5745_o2, G5213_o2, G5893_o2, G5391_o2, G4864_o2, G6143_o2, G6008_o2,
    G5565_o2, G5044_o2, G3813_o2, G4325_o2, G4834_o2, G4993_o2, G3989_o2,
    G4490_o2, G5011_o2, G5112_o2, n2776_lo_buf_o2, G3298_o2, G3073_o2,
    G3265_o2, G3624_o2, G1642_o2, G1980_o2, n2488_lo_buf_o2, G626_o2,
    G1139_o2, G950_o2, G707_o2, G545_o2, G4217_o2, G4716_o2, G5244_o2,
    G3136_o2, G3499_o2, G3885_o2, G5243_o2, G3886_o2, G4375_o2, G4901_o2,
    G5054_o2, G4374_o2, G4900_o2, G5053_o2, G5242_o2, G4034_o2, G4556_o2,
    G5064_o2, G5172_o2, G2030_o2, G3016_o2, G3520_o2, G3261_o2, G3620_o2,
    G4220_o2, G4719_o2, G5247_o2, G5109_o2, G1638_o2, G1976_o2, G3560_o2,
    G3205_o2, G3193_o2, G3367_o2, G3670_o2, n979_inv, G1280_o2, G902_o2,
    G659_o2, G983_o2, G740_o2, G2917_o2, G3391_o2, G3494_o2, G1512_o2,
    G1854_o2, G2203_o2, G3493_o2, G3069_o2, G3574_o2, G3319_o2, G3667_o2,
    G3068_o2, G3573_o2, G3666_o2, G3318_o2, G3492_o2, G3241_o2, G3722_o2,
    G3422_o2, G1445_o2, G3257_o2, G3616_o2, G1634_o2, G1972_o2, G2256_o2,
    G3394_o2, G3557_o2, G3364_o2, G3719_o2, G2253_o2, G1583_o2, G1917_o2,
    G1727_o2, G2061_o2, G935_o2, G692_o2, G2136_o2, G1507_o2, G1849_o2,
    G2198_o2, G2197_o2, G1848_o2, G1689_o2, G2016_o2, G2314_o2, G2313_o2,
    G1688_o2, G2015_o2, G1847_o2, G2196_o2, G2118_o2, G1777_o2, G1630_o2,
    G1968_o2, G2309_o2, G2139_o2, G1580_o2, G2250_o2, G1914_o2, G1724_o2,
    G2058_o2, n2728_lo_buf_o2;
  wire new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n853_, new_n855_, new_n857_, new_n859_, new_n861_, new_n863_,
    new_n865_, new_n867_, new_n869_, new_n871_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n929_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n937_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n946_, new_n947_, new_n949_,
    new_n952_, new_n953_, new_n955_, new_n958_, new_n959_, new_n961_,
    new_n964_, new_n965_, new_n967_, new_n970_, new_n971_, new_n973_,
    new_n976_, new_n977_, new_n979_, new_n982_, new_n983_, new_n985_,
    new_n988_, new_n989_, new_n991_, new_n994_, new_n995_, new_n997_,
    new_n998_, new_n999_, new_n1001_, new_n1003_, new_n1004_, new_n1006_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1029_, new_n1030_, new_n1032_, new_n1033_,
    new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1045_, new_n1047_, new_n1049_,
    new_n1052_, new_n1053_, new_n1055_, new_n1057_, new_n1059_, new_n1061_,
    new_n1063_, new_n1065_, new_n1067_, new_n1070_, new_n1071_, new_n1073_,
    new_n1075_, new_n1077_, new_n1079_, new_n1081_, new_n1083_, new_n1085_,
    new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1093_, new_n1094_,
    new_n1095_, new_n1097_, new_n1099_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1119_, new_n1120_, new_n1121_, new_n1123_, new_n1124_,
    new_n1125_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1141_, new_n1143_, new_n1145_, new_n1146_, new_n1147_, new_n1149_,
    new_n1151_, new_n1153_, new_n1155_, new_n1156_, new_n1157_, new_n1159_,
    new_n1161_, new_n1163_, new_n1165_, new_n1167_, new_n1169_, new_n1171_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1180_, new_n1181_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1189_, new_n1191_, new_n1193_, new_n1195_, new_n1196_,
    new_n1197_, new_n1199_, new_n1201_, new_n1203_, new_n1204_, new_n1205_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1213_,
    new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_,
    new_n1220_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1259_, new_n1261_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1290_, new_n1291_, new_n1293_, new_n1294_, new_n1295_,
    new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_,
    new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_,
    new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_,
    new_n1407_, new_n1408_, new_n1409_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1483_, new_n1484_, new_n1485_, new_n1486_,
    new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_,
    new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_,
    new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_,
    new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_,
    new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_,
    new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_,
    new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_,
    new_n1529_, new_n1530_, new_n1531_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_,
    new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_,
    new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_,
    new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_,
    new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_,
    new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_,
    new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_,
    new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_,
    new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_,
    new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_,
    new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_,
    new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_,
    new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_,
    new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_,
    new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_,
    new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_,
    new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_,
    new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_,
    new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_,
    new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_,
    new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_,
    new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_,
    new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_,
    new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_,
    new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_,
    new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_,
    new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_,
    new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_,
    new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_,
    new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_,
    new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_,
    new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_,
    new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_,
    new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_,
    new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_,
    new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_,
    new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_,
    new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_,
    new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_,
    new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_,
    new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_,
    new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_,
    new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_,
    new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_,
    new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_,
    new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_,
    new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_,
    new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_,
    new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_,
    new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_,
    new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_,
    new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_,
    new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_,
    new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_,
    new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_,
    new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_,
    new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_,
    new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_,
    new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_,
    new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_,
    new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_,
    new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_,
    new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_,
    new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_,
    new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_,
    new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_,
    new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_,
    new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_,
    new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_,
    new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_,
    new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_,
    new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_,
    new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_,
    new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_,
    new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_,
    new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_,
    new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_,
    new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_,
    new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_,
    new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_,
    new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_,
    new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_,
    new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_,
    new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_,
    new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_,
    new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_,
    new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_,
    new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_,
    new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_,
    new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_,
    new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_,
    new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_,
    new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_,
    new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_,
    new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_,
    new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_,
    new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_,
    new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_,
    new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_,
    new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_,
    new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_,
    new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_,
    new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_,
    new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_,
    new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_,
    new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_,
    new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_,
    new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_,
    new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_,
    new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_,
    new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_,
    new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_,
    new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_,
    new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_,
    new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_,
    new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_,
    new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_,
    new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_,
    new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_,
    new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_,
    new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_,
    new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_,
    new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_,
    new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_,
    new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_,
    new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_,
    new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_,
    new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_,
    new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_,
    new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_,
    new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_,
    new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_,
    new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_,
    new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_,
    new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_,
    new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_,
    new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_,
    new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_,
    new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_,
    new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_,
    new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_,
    new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_,
    new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_,
    new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_,
    new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_,
    new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_,
    new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_,
    new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_,
    new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_,
    new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_,
    new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_,
    new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_,
    new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_,
    new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_,
    new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_,
    new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_,
    new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_,
    new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_,
    new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_,
    new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_,
    new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_,
    new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_,
    new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_,
    new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_,
    new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_,
    new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_,
    new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_,
    new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_,
    new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_,
    new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_,
    new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_,
    new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_,
    new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_,
    new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_,
    new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_,
    new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_,
    new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_,
    new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_,
    new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_,
    new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_,
    new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_,
    new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_,
    new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_,
    new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_,
    new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_,
    new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_,
    new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_,
    new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_,
    new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_,
    new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_,
    new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_,
    new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_,
    new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_,
    new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_,
    new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_,
    new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_,
    new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_,
    new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_,
    new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_,
    new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_,
    new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_,
    new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_,
    new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_,
    new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_,
    new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_,
    new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_,
    new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_,
    new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_,
    new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_,
    new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_,
    new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_,
    new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_,
    new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_,
    new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_,
    new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_,
    new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_,
    new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_,
    new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_,
    new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_,
    new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_,
    new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_,
    new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_,
    new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_,
    new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_,
    new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_,
    new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_,
    new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_,
    new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_,
    new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_,
    new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_,
    new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_,
    new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_,
    new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_,
    new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_,
    new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_,
    new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_,
    new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_,
    new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_,
    new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_,
    new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_,
    new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_,
    new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_,
    new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_,
    new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_,
    new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_,
    new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_,
    new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_,
    new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_,
    new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_,
    new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_,
    new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_,
    new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_,
    new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_,
    new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_,
    new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_,
    new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_,
    new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_,
    new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_,
    new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_,
    new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_,
    new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_,
    new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_,
    new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_,
    new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_,
    new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_,
    new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_,
    new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_,
    new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_,
    new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_,
    new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_,
    new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_,
    new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_,
    new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_,
    new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_,
    new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_,
    new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_,
    new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_,
    new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_,
    new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_,
    new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_,
    new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_,
    new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_,
    new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_,
    new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_,
    new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_,
    new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_,
    new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_,
    new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_,
    new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_,
    new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_,
    new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_,
    new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_,
    new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_,
    new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_,
    new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_,
    new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_,
    new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_,
    new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_,
    new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_,
    new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_,
    new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_,
    new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_,
    new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_,
    new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_,
    new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_,
    new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_,
    new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_,
    new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_,
    new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_,
    new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_,
    new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_,
    new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_,
    new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_,
    new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_,
    new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_,
    new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_,
    new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_,
    new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_,
    new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_,
    new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_,
    new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_,
    new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_,
    new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_,
    new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_,
    new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_,
    new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_,
    new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_,
    new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_,
    new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_,
    new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_,
    new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_,
    new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_,
    new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_,
    new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_,
    new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_,
    new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_,
    new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_,
    new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_,
    new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_,
    new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_,
    new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_,
    new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_,
    new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_,
    new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_,
    new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_,
    new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_,
    new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_,
    new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_,
    new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_,
    new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_,
    new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_,
    new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_,
    new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_,
    new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_,
    new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_,
    new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_,
    new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_,
    new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_,
    new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_,
    new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_,
    new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_,
    new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_,
    new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_,
    new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_,
    new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_,
    new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_,
    new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_,
    new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_,
    new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_,
    new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_,
    new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_,
    new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_,
    new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_,
    new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_,
    new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_,
    new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_,
    new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_,
    new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_,
    new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_,
    new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_,
    new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_,
    new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_,
    new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_,
    new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_,
    new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_,
    new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_,
    new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_,
    new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_,
    new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_,
    new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_,
    new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_,
    new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_,
    new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_,
    new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_,
    new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_,
    new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_,
    new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_,
    new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_,
    new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_,
    new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_,
    new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_,
    new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_,
    new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_,
    new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_,
    new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_,
    new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_,
    new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_,
    new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_,
    new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_,
    new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_,
    new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_,
    new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_,
    new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_,
    new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_,
    new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_,
    new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_,
    new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_,
    new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_,
    new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_,
    new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_,
    new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_,
    new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_,
    new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_,
    new_n4614_, new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_,
    new_n4620_, new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_,
    new_n4626_, new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_,
    new_n4632_, new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_,
    new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_,
    new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_,
    new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_,
    new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_,
    new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_,
    new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_,
    new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4679_,
    new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_,
    new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_,
    new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_,
    new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_, new_n4703_,
    new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_, new_n4709_,
    new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_,
    new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_,
    new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_,
    new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_,
    new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_,
    new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_,
    new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_,
    new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_,
    new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_,
    new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_,
    new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_,
    new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_,
    new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_,
    new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_,
    new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_,
    new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_,
    new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_,
    new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_,
    new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_,
    new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_,
    new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_,
    new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_,
    new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_,
    new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_,
    new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_,
    new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_,
    new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_,
    new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_,
    new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_,
    new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_,
    new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_,
    new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_,
    new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_,
    new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_,
    new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_,
    new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_,
    new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_,
    new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_,
    new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_,
    new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_,
    new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_,
    new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_,
    new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_,
    new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_,
    new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_,
    new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_,
    new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_,
    new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_,
    new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_,
    new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_,
    new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_,
    new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_,
    new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_,
    new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_,
    new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_,
    new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_,
    new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_,
    new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_,
    new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_,
    new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_,
    new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_,
    new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_,
    new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_,
    new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_,
    new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_,
    new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_,
    new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_,
    new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_,
    new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_,
    new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_,
    new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_,
    new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_,
    new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_,
    new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_,
    new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_,
    new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_,
    new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_,
    new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_,
    new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_,
    new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_,
    new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_,
    new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_,
    new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_,
    new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_,
    new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_,
    new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_,
    new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_,
    new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_,
    new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_,
    new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_,
    new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_,
    new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_,
    new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_,
    new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_,
    new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_,
    new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_,
    new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_,
    new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_,
    new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_,
    new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_,
    new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_,
    new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_,
    new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_,
    new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_,
    new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_,
    new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_,
    new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_,
    new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_,
    new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_,
    new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_,
    new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_,
    new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_,
    new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_,
    new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_,
    new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_,
    new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_,
    new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_,
    new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_,
    new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_,
    new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_,
    new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_,
    new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_,
    new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_,
    new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_,
    new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_,
    new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_,
    new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_,
    new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_,
    new_n5490_, new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_,
    new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_,
    new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_,
    new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_,
    new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_,
    new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_,
    new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_,
    new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_,
    new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_,
    new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_,
    new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_,
    new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_,
    new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_,
    new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_,
    new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_,
    new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_,
    new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5591_,
    new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_,
    new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_,
    new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_,
    new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_,
    new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_,
    new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_,
    new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_,
    new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_,
    new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_,
    new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_,
    new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_,
    new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_,
    new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_,
    new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_,
    new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_,
    new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_,
    new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_,
    new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_,
    new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_,
    new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_,
    new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_,
    new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_,
    new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_,
    new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_,
    new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_,
    new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_,
    new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_,
    new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_,
    new_n5760_, new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_,
    new_n5766_, new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_,
    new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_,
    new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_,
    new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_,
    new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_,
    new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_,
    new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_,
    new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_,
    new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_,
    new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_,
    new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_,
    new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_,
    new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_,
    new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_,
    new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_,
    new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_,
    new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_,
    new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_,
    new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_,
    new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_,
    new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_,
    new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_,
    new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_,
    new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_,
    new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_,
    new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_,
    new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_,
    new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_,
    new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_,
    new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_,
    new_n5946_, new_n5947_, new_n6352_, new_n6353_, new_n6354_, new_n6355_,
    new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_, new_n6361_,
    new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_,
    new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_,
    new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_,
    new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_,
    new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_,
    new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_,
    new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_, new_n6403_,
    new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_,
    new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_,
    new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_,
    new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_,
    new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_,
    new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_,
    new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_,
    new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_,
    new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_,
    new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_,
    new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_,
    new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_,
    new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_,
    new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_,
    new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_,
    new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_,
    new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_,
    new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_,
    new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_,
    new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_, new_n6523_,
    new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_, new_n6529_,
    new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_, new_n6535_,
    new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_, new_n6541_,
    new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_, new_n6547_,
    new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_, new_n6553_,
    new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_, new_n6559_,
    new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_, new_n6565_,
    new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_, new_n6571_,
    new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_, new_n6577_,
    new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_, new_n6583_,
    new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_, new_n6589_,
    new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_, new_n6595_,
    new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_, new_n6601_,
    new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_, new_n6607_,
    new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_, new_n6613_,
    new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_, new_n6619_,
    new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_, new_n6625_,
    new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_, new_n6631_,
    new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_, new_n6637_,
    new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_, new_n6643_,
    new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_, new_n6649_,
    new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_, new_n6655_,
    new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_,
    new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_,
    new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_, new_n6673_,
    new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_, new_n6679_,
    new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_, new_n6685_,
    new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_, new_n6691_,
    new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_, new_n6697_,
    new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_,
    new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_,
    new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_,
    new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_,
    new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_,
    new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_,
    new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_, new_n6739_,
    new_n6740_, new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_,
    new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_,
    new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_,
    new_n6758_, new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_,
    new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_,
    new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n6775_,
    new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_, new_n6781_,
    new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_, new_n6787_,
    new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_,
    new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_,
    new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_,
    new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_,
    new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_,
    new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_,
    new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_,
    new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_,
    new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_,
    new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_,
    new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_,
    new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_,
    new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_,
    new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_,
    new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_,
    new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_,
    new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_,
    new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_,
    new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_,
    new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_,
    new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_,
    new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_,
    new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_,
    new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_,
    new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_,
    new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_,
    new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_,
    new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_,
    new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_,
    new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_,
    new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_,
    new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_,
    new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_,
    new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_,
    new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_,
    new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_,
    new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_,
    new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_,
    new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_,
    new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_,
    new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_,
    new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_,
    new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_,
    new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_,
    new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_,
    new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_,
    new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_,
    new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_,
    new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_,
    new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_,
    new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_,
    new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_,
    new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_,
    new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_,
    new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_,
    new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_,
    new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_,
    new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_,
    new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_,
    new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_,
    new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_,
    new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_,
    new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_,
    new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_,
    new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_,
    new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_,
    new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_,
    new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_,
    new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_,
    new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_,
    new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_,
    new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_,
    new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_,
    new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_,
    new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_,
    new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_,
    new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_,
    new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_,
    new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_,
    new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_,
    new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_,
    new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_,
    new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_,
    new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_,
    new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_,
    new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_,
    new_n7304_, new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_,
    new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_,
    new_n7316_, new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_,
    new_n7322_, new_n7323_, new_n7324_, new_n7325_, new_n7326_, new_n7327_,
    new_n7328_, new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_,
    new_n7334_, new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_,
    new_n7340_, new_n7341_, new_n7342_, new_n7343_, new_n7344_, new_n7345_,
    new_n7346_, new_n7347_, new_n7348_, new_n7349_, new_n7350_, new_n7351_,
    new_n7352_, new_n7353_, new_n7354_, new_n7355_, new_n7356_, new_n7357_,
    new_n7358_, new_n7359_, new_n7360_, new_n7361_, new_n7362_, new_n7363_,
    new_n7364_, new_n7365_, new_n7366_, new_n7367_, new_n7368_, new_n7369_,
    new_n7370_, new_n7371_, new_n7372_, new_n7373_, new_n7374_, new_n7375_,
    new_n7376_, new_n7377_, new_n7378_, new_n7379_, new_n7380_, new_n7381_,
    new_n7382_, new_n7383_, new_n7384_, new_n7385_, new_n7386_, new_n7387_,
    new_n7388_, new_n7389_, new_n7390_, new_n7391_, new_n7392_, new_n7393_,
    new_n7394_, new_n7395_, new_n7396_, new_n7397_, new_n7398_, new_n7399_,
    new_n7400_, new_n7401_, new_n7402_, new_n7403_, new_n7404_, new_n7405_,
    new_n7406_, new_n7407_, new_n7408_, new_n7409_, new_n7410_, new_n7411_,
    new_n7412_, new_n7413_, new_n7414_, new_n7415_, new_n7416_, new_n7417_,
    new_n7418_, new_n7419_, new_n7420_, new_n7421_, new_n7422_, new_n7423_,
    new_n7424_, new_n7425_, new_n7426_, new_n7427_, new_n7428_, new_n7429_,
    new_n7430_, new_n7431_, new_n7432_, new_n7433_, new_n7434_, new_n7435_,
    new_n7436_, new_n7437_, new_n7438_, new_n7439_, new_n7440_, new_n7441_,
    new_n7442_, new_n7443_, new_n7444_, new_n7445_, new_n7446_, new_n7447_,
    new_n7448_, new_n7449_, new_n7450_, new_n7451_, new_n7452_, new_n7453_,
    new_n7454_, new_n7455_, new_n7456_, new_n7457_, new_n7458_, new_n7459_,
    new_n7460_, new_n7461_, new_n7462_, new_n7463_, new_n7464_, new_n7465_,
    new_n7466_, new_n7467_, new_n7468_, new_n7469_, new_n7470_, new_n7471_,
    new_n7472_, new_n7473_, new_n7474_, new_n7475_, new_n7476_, new_n7477_,
    new_n7478_, new_n7479_, new_n7480_, new_n7481_, new_n7482_, new_n7483_,
    new_n7484_, new_n7485_, new_n7486_, new_n7487_, new_n7488_, new_n7489_,
    new_n7490_, new_n7491_, new_n7492_, new_n7493_, new_n7494_, new_n7495_,
    new_n7496_, new_n7497_, new_n7498_, new_n7499_, new_n7500_, new_n7501_,
    new_n7502_, new_n7503_, new_n7504_, new_n7505_, new_n7506_, new_n7507_,
    new_n7508_, new_n7509_, new_n7510_, new_n7511_, new_n7512_, new_n7513_,
    new_n7514_, new_n7515_, new_n7516_, new_n7517_, new_n7518_, new_n7519_,
    new_n7520_, new_n7521_, new_n7522_, new_n7523_, new_n7524_, new_n7525_,
    new_n7526_, new_n7527_, new_n7528_, new_n7529_, new_n7530_, new_n7531_,
    new_n7532_, new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_,
    new_n7538_, new_n7539_, new_n7540_, new_n7541_, new_n7542_, new_n7543_,
    new_n7544_, new_n7545_, new_n7546_, new_n7547_, new_n7548_, new_n7549_,
    new_n7550_, new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_,
    new_n7556_, new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_,
    new_n7562_, new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_,
    new_n7568_, new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_,
    new_n7574_, new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_,
    new_n7580_, new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_,
    new_n7586_, new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_,
    new_n7592_, new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_,
    new_n7598_, new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_,
    new_n7604_, new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_,
    new_n7610_, new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_,
    new_n7616_, new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_,
    new_n7622_, new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_,
    new_n7628_, new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_,
    new_n7634_, new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7639_,
    new_n7640_, new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_,
    new_n7646_, new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_,
    new_n7652_, new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_,
    new_n7658_, new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_,
    new_n7664_, new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_,
    new_n7670_, new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_,
    new_n7676_, new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_,
    new_n7682_, new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_,
    new_n7688_, new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_,
    new_n7694_, new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_,
    new_n7700_, new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_,
    new_n7706_, new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_,
    new_n7712_, new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_,
    new_n7718_, new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_,
    new_n7724_, new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_,
    new_n7730_, new_n7731_, new_n7732_, new_n7733_, new_n7734_, new_n7735_,
    new_n7736_, new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_,
    new_n7742_, new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_,
    new_n7748_, new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_,
    new_n7754_, new_n7755_, new_n7756_, new_n7757_, new_n7758_, new_n7759_,
    new_n7760_, new_n7761_, new_n7762_, new_n7763_, new_n7764_, new_n7765_,
    new_n7766_, new_n7767_, new_n7768_, new_n7769_, new_n7770_, new_n7771_,
    new_n7772_, new_n7773_, new_n7774_, new_n7775_, new_n7776_, new_n7777_,
    new_n7778_, new_n7779_, new_n7780_, new_n7781_, new_n7782_, new_n7783_,
    new_n7784_, new_n7785_, new_n7786_, new_n7787_, new_n7788_, new_n7789_,
    new_n7790_, new_n7791_, new_n7792_, new_n7793_, new_n7794_, new_n7795_,
    new_n7796_, new_n7797_, new_n7798_, new_n7799_, new_n7800_, new_n7801_,
    new_n7802_, new_n7803_, new_n7804_, new_n7805_, new_n7806_, new_n7807_,
    new_n7808_, new_n7809_, new_n7810_, new_n7811_, new_n7812_, new_n7813_,
    new_n7814_, new_n7815_, new_n7816_, new_n7817_, new_n7818_, new_n7819_,
    new_n7820_, new_n7821_, new_n7822_, new_n7823_, new_n7824_, new_n7825_,
    new_n7826_, new_n7827_, new_n7828_, new_n7829_, new_n7830_, new_n7831_,
    new_n7832_, new_n7833_, new_n7834_, new_n7835_, new_n7836_, new_n7837_,
    new_n7838_, new_n7839_, new_n7840_, new_n7841_, new_n7842_, new_n7843_,
    new_n7844_, new_n7845_, new_n7846_, new_n7847_, new_n7848_, new_n7849_,
    new_n7850_, new_n7851_, new_n7852_, new_n7853_, new_n7854_, new_n7855_,
    new_n7856_, new_n7857_, new_n7858_, new_n7859_, new_n7860_, new_n7861_,
    new_n7862_, new_n7863_, new_n7864_, new_n7865_, new_n7866_, new_n7867_,
    new_n7868_, new_n7869_, new_n7870_, new_n7871_, new_n7872_, new_n7873_,
    new_n7874_, new_n7875_, new_n7876_, new_n7877_, new_n7878_, new_n7879_,
    new_n7880_, new_n7881_, new_n7882_, new_n7883_, new_n7884_, new_n7885_,
    new_n7886_, new_n7887_, new_n7888_, new_n7889_, new_n7890_, new_n7891_,
    new_n7892_, new_n7893_, new_n7894_, new_n7895_, new_n7896_, new_n7897_,
    new_n7898_, new_n7899_, new_n7900_, new_n7901_, new_n7902_, new_n7903_,
    new_n7904_, new_n7905_, new_n7906_, new_n7907_, new_n7908_, new_n7909_,
    new_n7910_, new_n7911_, new_n7912_, new_n7913_, new_n7914_, new_n7915_,
    new_n7916_, new_n7917_, new_n7918_, new_n7919_, new_n7920_, new_n7921_,
    new_n7922_, new_n7923_, new_n7924_, new_n7925_, new_n7926_, new_n7927_,
    new_n7928_, new_n7929_, new_n7930_, new_n7931_, new_n7932_, new_n7933_,
    new_n7934_, new_n7935_, new_n7936_, new_n7937_, new_n7938_, new_n7939_,
    new_n7940_, new_n7941_, new_n7942_, new_n7943_, new_n7944_, new_n7945_,
    new_n7946_, new_n7947_, new_n7948_, new_n7949_, new_n7950_, new_n7951_,
    new_n7952_, new_n7953_, new_n7954_, new_n7955_, new_n7956_, new_n7957_,
    new_n7958_, new_n7959_, new_n7960_, new_n7961_, new_n7962_, new_n7963_,
    new_n7964_, new_n7965_, new_n7966_, new_n7967_, new_n7968_, new_n7969_,
    new_n7970_, new_n7971_, new_n7972_, new_n7973_, new_n7974_, new_n7975_,
    new_n7976_, new_n7977_, new_n7978_, new_n7979_, new_n7980_, new_n7981_,
    new_n7982_, new_n7983_, new_n7984_, new_n7985_, new_n7986_, new_n7987_,
    new_n7988_, new_n7989_, new_n7990_, new_n7991_, new_n7992_, new_n7993_,
    new_n7994_, new_n7995_, new_n7996_, new_n7997_, new_n7998_, new_n7999_,
    new_n8000_, new_n8001_, new_n8002_, new_n8003_, new_n8004_, new_n8005_,
    new_n8006_, new_n8007_, new_n8008_, new_n8009_, new_n8010_, new_n8011_,
    new_n8012_, new_n8013_, new_n8014_, new_n8015_, new_n8016_, new_n8017_,
    new_n8018_, new_n8019_, new_n8020_, new_n8021_, new_n8022_, new_n8023_,
    new_n8024_, new_n8025_, new_n8026_, new_n8027_, new_n8028_, new_n8029_,
    new_n8030_, new_n8031_, new_n8032_, new_n8033_, new_n8034_, new_n8035_,
    new_n8036_, new_n8037_, new_n8038_, new_n8039_, new_n8040_, new_n8041_,
    new_n8042_, new_n8043_, new_n8044_, new_n8045_, new_n8046_, new_n8047_,
    new_n8048_, new_n8049_, new_n8050_, new_n8051_, new_n8052_, new_n8053_,
    new_n8054_, new_n8055_, new_n8056_, new_n8057_, new_n8058_, new_n8059_,
    new_n8060_, new_n8061_, new_n8062_, new_n8063_, new_n8064_, new_n8065_,
    new_n8066_, new_n8067_, new_n8068_, new_n8069_, new_n8070_, new_n8071_,
    new_n8072_, new_n8073_, new_n8074_, new_n8075_, new_n8076_, new_n8077_,
    new_n8078_, new_n8079_, new_n8080_, new_n8081_, new_n8082_, new_n8083_,
    new_n8084_, new_n8085_, new_n8086_, new_n8087_, new_n8088_, new_n8089_,
    new_n8090_, new_n8091_, new_n8092_, new_n8093_, new_n8094_, new_n8095_,
    new_n8096_, new_n8097_, new_n8098_, new_n8099_, new_n8100_, new_n8101_,
    new_n8102_, new_n8103_, new_n8104_, new_n8105_, new_n8106_, new_n8107_,
    new_n8108_, new_n8109_, new_n8110_, new_n8111_, new_n8112_, new_n8113_,
    new_n8114_, new_n8115_, new_n8116_, new_n8117_, new_n8118_, new_n8119_,
    new_n8120_, new_n8121_, new_n8122_, new_n8123_, new_n8124_, new_n8125_,
    new_n8126_, new_n8127_, new_n8128_, new_n8129_, new_n8130_, new_n8131_,
    new_n8132_, new_n8133_, new_n8134_, new_n8135_, new_n8136_, new_n8137_,
    new_n8138_, new_n8139_, new_n8140_, new_n8141_, new_n8142_, new_n8143_,
    new_n8144_, new_n8145_, new_n8146_, new_n8147_, new_n8148_, new_n8149_,
    new_n8150_, new_n8151_, new_n8152_, new_n8153_, new_n8154_, new_n8155_,
    new_n8156_, new_n8157_, new_n8158_, new_n8159_, new_n8160_, new_n8161_,
    new_n8162_, new_n8163_, new_n8164_, new_n8165_, new_n8166_, new_n8167_,
    new_n8168_, new_n8169_, new_n8170_, new_n8171_, new_n8172_, new_n8173_,
    new_n8174_, new_n8175_, new_n8176_, new_n8177_, new_n8178_, new_n8179_,
    new_n8180_, new_n8181_, new_n8182_, new_n8183_, new_n8184_, new_n8185_,
    new_n8186_, new_n8187_, new_n8188_, new_n8189_, new_n8190_, new_n8191_,
    new_n8192_, new_n8193_, new_n8194_, new_n8195_, new_n8196_, new_n8197_,
    new_n8198_, new_n8199_, new_n8200_, new_n8201_, new_n8202_, new_n8203_,
    new_n8204_, new_n8205_, new_n8206_, new_n8207_, new_n8208_, new_n8209_,
    new_n8210_, new_n8211_, new_n8212_, new_n8213_, new_n8214_, new_n8215_,
    new_n8216_, new_n8217_, new_n8218_, new_n8219_, new_n8220_, new_n8221_,
    new_n8222_, new_n8223_, new_n8224_, new_n8225_, new_n8226_, new_n8227_,
    new_n8228_, new_n8229_, new_n8230_, new_n8231_, new_n8232_, new_n8233_,
    new_n8234_, new_n8235_, new_n8236_, new_n8237_, new_n8238_, new_n8239_,
    new_n8240_, new_n8241_, new_n8242_, new_n8243_, new_n8244_, new_n8245_,
    new_n8246_, new_n8247_, new_n8248_, new_n8249_, new_n8250_, new_n8251_,
    new_n8252_, new_n8253_, new_n8254_, new_n8255_, new_n8256_, new_n8257_,
    new_n8258_, new_n8259_, new_n8260_, new_n8261_, new_n8262_, new_n8263_,
    new_n8264_, new_n8265_, new_n8266_, new_n8267_, new_n8268_, new_n8269_,
    new_n8270_, new_n8271_, new_n8272_, new_n8273_, new_n8274_, new_n8275_,
    new_n8276_, new_n8277_, new_n8278_, new_n8279_, new_n8280_, new_n8281_,
    new_n8282_, new_n8283_, new_n8284_, new_n8285_, new_n8286_, new_n8287_,
    new_n8288_, new_n8289_, new_n8290_, new_n8291_, new_n8292_, new_n8293_,
    new_n8294_, new_n8295_, new_n8296_, new_n8297_, new_n8298_, new_n8299_,
    new_n8300_, new_n8301_, new_n8302_, new_n8303_, new_n8304_, new_n8305_,
    new_n8306_, new_n8307_, new_n8308_, new_n8309_, new_n8310_, new_n8311_,
    new_n8312_, new_n8313_, new_n8314_, new_n8315_, new_n8316_, new_n8317_,
    new_n8318_, new_n8319_, new_n8320_, new_n8321_, new_n8322_, new_n8323_,
    new_n8324_, new_n8325_, new_n8326_, new_n8327_, new_n8328_, new_n8329_,
    new_n8330_, new_n8331_, new_n8332_, new_n8333_, new_n8334_, new_n8335_,
    new_n8336_, new_n8337_, new_n8338_, new_n8339_, new_n8340_, new_n8341_,
    new_n8342_, new_n8343_, new_n8344_, new_n8345_, new_n8346_, new_n8347_,
    new_n8348_, new_n8349_, new_n8350_, new_n8351_, new_n8352_, new_n8353_,
    new_n8354_, new_n8355_, new_n8356_, new_n8357_, new_n8358_, new_n8359_,
    new_n8360_, new_n8361_, new_n8362_, new_n8363_, new_n8364_, new_n8365_,
    new_n8366_, new_n8367_, new_n8368_, new_n8369_, new_n8370_, new_n8371_,
    new_n8372_, new_n8373_, new_n8374_, new_n8375_, new_n8376_, new_n8377_,
    new_n8378_, new_n8379_, new_n8380_, new_n8381_, new_n8382_, new_n8383_,
    new_n8384_, new_n8385_, new_n8386_, new_n8387_, new_n8388_, new_n8389_,
    new_n8390_, new_n8391_, new_n8392_, new_n8393_, new_n8394_, new_n8395_,
    new_n8396_, new_n8397_, new_n8398_, new_n8399_, new_n8400_, new_n8401_,
    new_n8402_, new_n8403_, new_n8404_, new_n8405_, new_n8406_, new_n8407_,
    new_n8408_, new_n8409_, new_n8410_, new_n8411_, new_n8412_, new_n8413_,
    new_n8414_, new_n8415_, new_n8416_, new_n8417_, new_n8418_, new_n8419_,
    new_n8420_, new_n8421_, new_n8422_, new_n8423_, new_n8424_, new_n8425_,
    new_n8426_, new_n8427_, new_n8428_, new_n8429_, new_n8430_, new_n8431_,
    new_n8432_, new_n8433_, new_n8434_, new_n8435_, new_n8436_, new_n8437_,
    new_n8438_, new_n8439_, new_n8440_, new_n8441_, new_n8442_, new_n8443_,
    new_n8444_, new_n8445_, new_n8446_, new_n8447_, new_n8448_, new_n8449_,
    new_n8450_, new_n8451_, new_n8452_, new_n8453_, new_n8454_, new_n8455_,
    new_n8456_, new_n8457_, new_n8458_, new_n8459_, new_n8460_, new_n8461_,
    new_n8462_, new_n8463_, new_n8464_, new_n8465_, new_n8466_, new_n8467_,
    new_n8468_, new_n8469_, new_n8470_, new_n8471_, new_n8472_, new_n8473_,
    new_n8474_, new_n8475_, new_n8476_, new_n8477_, new_n8478_, new_n8479_,
    new_n8480_, new_n8481_, new_n8482_, new_n8483_, new_n8484_, new_n8485_,
    new_n8486_, new_n8487_, new_n8488_, new_n8489_, new_n8490_, new_n8491_,
    new_n8492_, new_n8493_, new_n8494_, new_n8495_, new_n8496_, new_n8497_,
    new_n8498_, new_n8499_, new_n8500_, new_n8501_, new_n8502_, new_n8503_,
    new_n8504_, new_n8505_, new_n8506_, new_n8507_, new_n8508_, new_n8509_,
    new_n8510_, new_n8511_, new_n8512_, new_n8513_, new_n8514_, new_n8515_,
    new_n8516_, new_n8517_, new_n8518_, new_n8519_, new_n8520_, new_n8521_,
    new_n8522_, new_n8523_, new_n8524_, new_n8525_, new_n8526_, new_n8527_,
    new_n8528_, new_n8529_, new_n8530_, new_n8531_, new_n8532_, new_n8533_,
    new_n8534_, new_n8535_, new_n8536_, new_n8537_, new_n8538_, new_n8539_,
    new_n8540_, new_n8541_, new_n8542_, new_n8543_, new_n8544_, new_n8545_,
    new_n8546_, new_n8547_, new_n8548_, new_n8549_, new_n8550_, new_n8551_,
    new_n8552_, new_n8553_, new_n8554_, new_n8555_, new_n8556_, new_n8557_,
    new_n8558_, new_n8559_, new_n8560_, new_n8561_, new_n8562_, new_n8563_,
    new_n8564_, new_n8565_, new_n8566_, new_n8567_, new_n8568_, new_n8569_,
    new_n8570_, new_n8571_, new_n8572_, new_n8573_, new_n8574_, new_n8575_,
    new_n8576_, new_n8577_, new_n8578_, new_n8579_, new_n8580_, new_n8581_,
    new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_, new_n8587_,
    new_n8588_, new_n8589_, new_n8590_, new_n8591_, new_n8592_, new_n8593_,
    new_n8594_, new_n8595_, new_n8596_, new_n8597_, new_n8598_, new_n8599_,
    new_n8600_, new_n8601_, new_n8602_, new_n8603_, new_n8604_, new_n8605_,
    new_n8606_, new_n8607_, new_n8608_, new_n8609_, new_n8610_, new_n8611_,
    new_n8612_, new_n8613_, new_n8614_, new_n8615_, new_n8616_, new_n8617_,
    new_n8618_, new_n8619_, new_n8620_, new_n8621_, new_n8622_, new_n8623_,
    new_n8624_, new_n8625_, new_n8626_, new_n8627_, new_n8628_, new_n8629_,
    new_n8630_, new_n8631_, new_n8632_, new_n8633_, new_n8634_, new_n8635_,
    new_n8636_, new_n8637_, new_n8638_, new_n8639_, new_n8640_, new_n8641_,
    new_n8642_, new_n8643_, new_n8644_, new_n8645_, new_n8646_, new_n8647_,
    new_n8648_, new_n8649_, new_n8650_, new_n8651_, new_n8652_, new_n8653_,
    new_n8654_, new_n8655_, new_n8656_, new_n8657_, new_n8658_, new_n8659_,
    new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8664_, new_n8665_,
    new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_, new_n8671_,
    new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8676_, new_n8677_,
    new_n8678_, new_n8679_, new_n8680_, new_n8681_, new_n8682_, new_n8683_,
    new_n8684_, new_n8685_, new_n8686_, new_n8687_, new_n8688_, new_n8689_,
    new_n8690_, new_n8691_, new_n8692_, new_n8693_, new_n8694_, new_n8695_,
    new_n8696_, new_n8697_, new_n8698_, new_n8699_, new_n8700_, new_n8701_,
    new_n8702_, new_n8703_, new_n8704_, new_n8705_, new_n8706_, new_n8707_,
    new_n8708_, new_n8709_, new_n8710_, new_n8711_, new_n8712_, new_n8713_,
    new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_, new_n8719_,
    new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_, new_n8725_,
    new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_, new_n8731_,
    new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_, new_n8737_,
    new_n8738_, new_n8739_, new_n8740_, new_n8741_, new_n8742_, new_n8743_,
    new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_, new_n8749_,
    new_n8750_, new_n8751_, new_n8752_, new_n8753_, new_n8754_, new_n8755_,
    new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_, new_n8761_,
    new_n8762_, new_n8763_, new_n8764_, new_n8765_, new_n8766_, new_n8767_,
    new_n8768_, new_n8769_, new_n8770_, new_n8771_, new_n8772_, new_n8773_,
    new_n8774_, new_n8775_, new_n8776_, new_n8777_, new_n8778_, new_n8779_,
    new_n8780_, new_n8781_, new_n8782_, new_n8783_, new_n8784_, new_n8785_,
    new_n8786_, new_n8787_, new_n8788_, new_n8789_, new_n8790_, new_n8791_,
    new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_, new_n8797_,
    new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_, new_n8803_,
    new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_, new_n8809_,
    new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_, new_n8815_,
    new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_, new_n8821_,
    new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_, new_n8827_,
    new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_, new_n8833_,
    new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_, new_n8839_,
    new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_, new_n8845_,
    new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_, new_n8851_,
    new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_, new_n8857_,
    new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_, new_n8863_,
    new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_, new_n8869_,
    new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_, new_n8875_,
    new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_, new_n8881_,
    new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_, new_n8887_,
    new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_, new_n8893_,
    new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_, new_n8899_,
    new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_, new_n8905_,
    new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_, new_n8911_,
    new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_, new_n8917_,
    new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_, new_n8923_,
    new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_, new_n8929_,
    new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_, new_n8935_,
    new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_, new_n8941_,
    new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_, new_n8947_,
    new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_, new_n8953_,
    new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_, new_n8959_,
    new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_, new_n8965_,
    new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_,
    new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_,
    new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_,
    new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_, new_n8989_,
    new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_, new_n8995_,
    new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_, new_n9001_,
    new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_, new_n9007_,
    new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_, new_n9013_,
    new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_,
    new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9024_, new_n9025_,
    new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_,
    new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_,
    new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_,
    new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_,
    new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_,
    new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_,
    new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_,
    new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_,
    new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_,
    new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_, new_n9085_,
    new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_, new_n9091_,
    new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_,
    new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_,
    new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9109_,
    new_n9110_, new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_,
    new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_,
    new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_,
    new_n9128_, new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_,
    new_n9134_, new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_,
    new_n9140_, new_n9141_, new_n9142_, new_n9143_, new_n9144_, new_n9145_,
    new_n9146_, new_n9147_, new_n9148_, new_n9149_, new_n9150_, new_n9151_,
    new_n9152_, new_n9153_, new_n9154_, new_n9155_, new_n9156_, new_n9157_,
    new_n9158_, new_n9159_, new_n9160_, new_n9161_, new_n9162_, new_n9163_,
    new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_, new_n9169_,
    new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_, new_n9175_,
    new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_, new_n9181_,
    new_n9182_, new_n9183_, new_n9184_, new_n9185_, new_n9186_, new_n9187_,
    new_n9188_, new_n9189_, new_n9190_, new_n9191_, new_n9192_, new_n9193_,
    new_n9194_, new_n9195_, new_n9196_, new_n9197_, new_n9198_, new_n9199_,
    new_n9200_, new_n9201_, new_n9202_, new_n9203_, new_n9204_, new_n9205_,
    new_n9206_, new_n9207_, new_n9208_, new_n9209_, new_n9210_, new_n9211_,
    new_n9212_, new_n9213_, new_n9214_, new_n9215_, new_n9216_, new_n9217_,
    new_n9218_, new_n9219_, new_n9220_, new_n9221_, new_n9222_, new_n9223_,
    new_n9224_, new_n9225_, new_n9226_, new_n9227_, new_n9228_, new_n9229_,
    new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_, new_n9235_,
    new_n9236_, new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_,
    new_n9242_, new_n9243_, new_n9244_, new_n9245_, new_n9246_, new_n9247_,
    new_n9248_, new_n9249_, new_n9250_, new_n9251_, new_n9252_, new_n9253_,
    new_n9254_, new_n9255_, new_n9256_, new_n9257_, new_n9258_, new_n9259_,
    new_n9260_, new_n9261_, new_n9262_, new_n9263_, new_n9264_, new_n9265_,
    new_n9266_, new_n9267_, new_n9268_, new_n9269_, new_n9270_, new_n9271_,
    new_n9272_, new_n9273_, new_n9274_, new_n9275_, new_n9276_, new_n9277_,
    new_n9278_, new_n9279_, new_n9280_, new_n9281_, new_n9282_, new_n9283_,
    new_n9284_, new_n9285_, new_n9286_, new_n9287_, new_n9288_, new_n9289_,
    new_n9290_, new_n9291_, new_n9292_, new_n9293_, new_n9294_, new_n9295_,
    new_n9296_, new_n9297_, new_n9298_, new_n9299_, new_n9300_, new_n9301_,
    new_n9302_, new_n9303_, new_n9304_, new_n9305_, new_n9306_, new_n9307_,
    new_n9308_, new_n9309_, new_n9310_, new_n9311_, new_n9312_, new_n9313_,
    new_n9314_, new_n9315_, new_n9316_, new_n9317_, new_n9318_, new_n9319_,
    new_n9320_, new_n9321_, new_n9322_, new_n9323_, new_n9324_, new_n9325_,
    new_n9326_, new_n9327_, new_n9328_, new_n9329_, new_n9330_, new_n9331_,
    new_n9332_, new_n9333_, new_n9334_, new_n9335_, new_n9336_, new_n9337_,
    new_n9338_, new_n9339_, new_n9340_, new_n9341_, new_n9342_, new_n9343_,
    new_n9344_, new_n9345_, new_n9346_, new_n9347_, new_n9348_, new_n9349_,
    new_n9350_, new_n9351_, new_n9352_, new_n9353_, new_n9354_, new_n9355_,
    new_n9356_, new_n9357_, new_n9358_, new_n9359_, new_n9360_, new_n9361_,
    new_n9362_, new_n9363_, new_n9364_, new_n9365_, new_n9366_, new_n9367_,
    new_n9368_, new_n9369_, new_n9370_, new_n9371_, new_n9372_, new_n9373_,
    new_n9374_, new_n9375_, new_n9376_, new_n9377_, new_n9378_, new_n9379_,
    new_n9380_, new_n9381_, new_n9382_, new_n9383_, new_n9384_, new_n9385_,
    new_n9386_, new_n9387_, new_n9388_, new_n9389_, new_n9390_, new_n9391_,
    new_n9392_, new_n9393_, new_n9394_, new_n9395_, new_n9396_, new_n9397_,
    new_n9398_, new_n9399_, new_n9400_, new_n9401_, new_n9402_, new_n9403_,
    new_n9404_, new_n9405_, new_n9406_, new_n9407_, new_n9408_, new_n9409_,
    new_n9410_, new_n9411_, new_n9412_, new_n9413_, new_n9414_, new_n9415_,
    new_n9416_, new_n9417_, new_n9418_, new_n9419_, new_n9420_, new_n9421_,
    new_n9422_, new_n9423_, new_n9424_, new_n9425_, new_n9426_, new_n9427_,
    new_n9428_, new_n9429_, new_n9430_, new_n9431_, new_n9432_, new_n9433_,
    new_n9434_, new_n9435_, new_n9436_, new_n9437_, new_n9438_, new_n9439_,
    new_n9440_, new_n9441_, new_n9442_, new_n9443_, new_n9444_, new_n9445_,
    new_n9446_, new_n9447_, new_n9448_, new_n9449_, new_n9450_, new_n9451_,
    new_n9452_, new_n9453_, new_n9454_, new_n9455_, new_n9456_, new_n9457_,
    new_n9458_, new_n9459_, new_n9460_, new_n9461_, new_n9462_, new_n9463_,
    new_n9464_, new_n9465_, new_n9466_, new_n9467_, new_n9468_, new_n9469_,
    new_n9470_, new_n9471_, new_n9472_, new_n9473_, new_n9474_, new_n9475_,
    new_n9476_, new_n9477_, new_n9478_, new_n9479_, new_n9480_, new_n9481_,
    new_n9482_, new_n9483_, new_n9484_, new_n9485_, new_n9486_, new_n9487_,
    new_n9488_, new_n9489_, new_n9490_, new_n9491_, new_n9492_, new_n9493_,
    new_n9494_, new_n9495_, new_n9496_, new_n9497_, new_n9498_, new_n9499_,
    new_n9500_, new_n9501_, new_n9502_, new_n9503_, new_n9504_, new_n9505_,
    new_n9506_, new_n9507_, new_n9508_, new_n9509_, new_n9510_, new_n9511_,
    new_n9512_, new_n9513_, new_n9514_, new_n9515_, new_n9516_, new_n9517_,
    new_n9518_, new_n9519_, new_n9520_, new_n9521_, new_n9522_, new_n9523_,
    new_n9524_, new_n9525_, new_n9526_, new_n9527_, new_n9528_, new_n9529_,
    new_n9530_, new_n9531_, new_n9532_, new_n9533_, new_n9534_, new_n9535_,
    new_n9536_, new_n9537_, new_n9538_, new_n9539_, new_n9540_, new_n9541_,
    new_n9542_, new_n9543_, new_n9544_, new_n9545_, new_n9546_, new_n9547_,
    new_n9548_, new_n9549_, new_n9550_, new_n9551_, new_n9552_, new_n9553_,
    new_n9554_, new_n9555_, new_n9556_, new_n9557_, new_n9558_, new_n9559_,
    new_n9560_, new_n9561_, new_n9562_, new_n9563_, new_n9564_, new_n9565_,
    new_n9566_, new_n9567_, new_n9568_, new_n9569_, new_n9570_, new_n9571_,
    new_n9572_, new_n9573_, new_n9574_, new_n9575_, new_n9576_, new_n9577_,
    new_n9578_, new_n9579_, new_n9580_, new_n9581_, new_n9582_, new_n9583_,
    new_n9584_, new_n9585_, new_n9586_, new_n9587_, new_n9588_, new_n9589_,
    new_n9590_, new_n9591_, new_n9592_, new_n9593_, new_n9594_, new_n9595_,
    new_n9596_, new_n9597_, new_n9598_, new_n9599_, new_n9600_, new_n9601_,
    new_n9602_, new_n9603_, new_n9604_, new_n9605_, new_n9606_, new_n9607_,
    new_n9608_, new_n9609_, new_n9610_, new_n9611_, new_n9612_, new_n9613_,
    new_n9614_, new_n9615_, new_n9616_, new_n9617_, new_n9618_, new_n9619_,
    new_n9620_, new_n9621_, new_n9622_, new_n9623_, new_n9624_, new_n9625_,
    new_n9626_, new_n9627_, new_n9628_, new_n9629_, new_n9630_, new_n9631_,
    new_n9632_, new_n9633_, new_n9634_, new_n9635_, new_n9636_, new_n9637_,
    new_n9638_, new_n9639_, new_n9640_, new_n9641_, new_n9642_, new_n9643_,
    new_n9644_, new_n9645_, new_n9646_, new_n9647_, new_n9648_, new_n9649_,
    new_n9650_, new_n9651_, new_n9652_, new_n9653_, new_n9654_, new_n9655_,
    new_n9656_, new_n9657_, new_n9658_, new_n9659_, new_n9660_, new_n9661_,
    new_n9662_, new_n9663_, new_n9664_, new_n9665_, new_n9666_, new_n9667_,
    new_n9668_, new_n9669_, new_n9670_, new_n9671_, new_n9672_, new_n9673_,
    new_n9674_, new_n9675_, new_n9676_, new_n9677_, new_n9678_, new_n9679_,
    new_n9680_, new_n9681_, new_n9682_, new_n9683_, new_n9684_, new_n9685_,
    new_n9686_, new_n9687_, new_n9688_, new_n9689_, new_n9690_, new_n9691_,
    new_n9692_, new_n9693_, new_n9694_, new_n9695_, new_n9696_, new_n9697_,
    new_n9698_, new_n9699_, new_n9700_, new_n9701_, new_n9702_, new_n9703_,
    new_n9704_, new_n9705_, new_n9706_, new_n9707_, new_n9708_, new_n9709_,
    new_n9710_, new_n9711_, new_n9712_, new_n9713_, new_n9714_, new_n9715_,
    new_n9716_, new_n9717_, new_n9718_, new_n9719_, new_n9720_, new_n9721_,
    new_n9722_, new_n9723_, new_n9724_, new_n9725_, new_n9726_, new_n9727_,
    new_n9728_, new_n9729_, new_n9730_, new_n9731_, new_n9732_, new_n9733_,
    new_n9734_, new_n9735_, new_n9736_, new_n9737_, new_n9738_, new_n9739_,
    new_n9740_, new_n9741_, new_n9742_, new_n9743_, new_n9744_, new_n9745_,
    new_n9746_, new_n9747_, new_n9748_, new_n9749_, new_n9750_, new_n9751_,
    new_n9752_, new_n9753_, new_n9754_, new_n9755_, new_n9756_, new_n9757_,
    new_n9758_, new_n9759_, new_n9760_, new_n9761_, new_n9762_, new_n9763_,
    new_n9764_, new_n9765_, new_n9766_, new_n9767_, new_n9768_, new_n9769_,
    new_n9770_, new_n9771_, new_n9772_, new_n9773_, new_n9774_, new_n9775_,
    new_n9776_, new_n9777_, new_n9778_, new_n9779_, new_n9780_, new_n9781_,
    new_n9782_, new_n9783_, new_n9784_, new_n9785_, new_n9786_, new_n9787_,
    new_n9788_, new_n9789_, new_n9790_, new_n9791_, new_n9792_, new_n9793_,
    new_n9794_, new_n9795_, new_n9796_, new_n9797_, new_n9798_, new_n9799_,
    new_n9800_, new_n9801_, new_n9802_, new_n9803_, new_n9804_, new_n9805_,
    new_n9806_, new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_,
    new_n9812_, new_n9813_, new_n9814_, new_n9815_, new_n9816_, new_n9817_,
    new_n9818_, new_n9819_, new_n9820_, new_n9821_, new_n9822_, new_n9823_,
    new_n9824_, new_n9825_, new_n9826_, new_n9827_, new_n9828_, new_n9829_,
    new_n9830_, new_n9831_, new_n9832_, new_n9833_, new_n9834_, new_n9835_,
    new_n9836_, new_n9837_, new_n9838_, new_n9839_, new_n9840_, new_n9841_,
    new_n9842_, new_n9843_, new_n9844_, new_n9845_, new_n9846_, new_n9847_,
    new_n9848_, new_n9849_, new_n9850_, new_n9851_, new_n9852_, new_n9853_,
    new_n9854_, new_n9855_, new_n9856_, new_n9857_, new_n9858_, new_n9859_,
    new_n9860_, new_n9861_, new_n9862_, new_n9863_, new_n9864_, new_n9865_,
    new_n9866_, new_n9867_, new_n9868_, new_n9869_, new_n9870_, new_n9871_,
    new_n9872_, new_n9873_, new_n9874_, new_n9875_, new_n9876_, new_n9877_,
    new_n9878_, new_n9879_, new_n9880_, new_n9881_, new_n9882_, new_n9883_,
    new_n9884_, new_n9885_, new_n9886_, new_n9887_, new_n9888_, new_n9889_,
    new_n9890_, new_n9891_, new_n9892_, new_n9893_, new_n9894_, new_n9895_,
    new_n9896_, new_n9897_, new_n9898_, new_n9899_, new_n9900_, new_n9901_,
    new_n9902_, new_n9903_, new_n9904_, new_n9905_, new_n9906_, new_n9907_,
    new_n9908_, new_n9909_, new_n9910_, new_n9911_, new_n9912_, new_n9913_,
    new_n9914_, new_n9915_, new_n9916_, new_n9917_, new_n9918_, new_n9919_,
    new_n9920_, new_n9921_, new_n9922_, new_n9923_, new_n9924_, new_n9925_,
    new_n9926_, new_n9927_, new_n9928_, new_n9929_, new_n9930_, new_n9931_,
    new_n9932_, new_n9933_, new_n9934_, new_n9935_, new_n9936_, new_n9937_,
    new_n9938_, new_n9939_, new_n9940_, new_n9941_, new_n9942_, new_n9943_,
    new_n9944_, new_n9945_, new_n9946_, new_n9947_, new_n9948_, new_n9949_,
    new_n9950_, new_n9951_, new_n9952_, new_n9953_, new_n9954_, new_n9955_,
    new_n9956_, new_n9957_, new_n9958_, new_n9959_, new_n9960_, new_n9961_,
    new_n9962_, new_n9963_, new_n9964_, new_n9965_, new_n9966_, new_n9967_,
    new_n9968_, new_n9969_, new_n9970_, new_n9971_, new_n9972_, new_n9973_,
    new_n9974_, new_n9975_, new_n9976_, new_n9977_, new_n9978_, new_n9979_,
    new_n9980_, new_n9981_, new_n9982_, new_n9983_, new_n9984_, new_n9985_,
    new_n9986_, new_n9987_, new_n9988_, new_n9989_, new_n9990_, new_n9991_,
    new_n9992_, new_n9993_, new_n9994_, new_n9995_, new_n9996_, new_n9997_,
    new_n9998_, new_n9999_, new_n10000_, new_n10001_, new_n10002_,
    new_n10003_, new_n10004_, new_n10005_, new_n10006_, new_n10007_,
    new_n10008_, new_n10009_, new_n10010_, new_n10011_, new_n10012_,
    new_n10013_, new_n10014_, new_n10015_, new_n10016_, new_n10017_,
    new_n10018_, new_n10019_, new_n10020_, new_n10021_, new_n10022_,
    new_n10023_, new_n10024_, new_n10025_, new_n10026_, new_n10027_,
    new_n10028_, new_n10029_, new_n10030_, new_n10031_, new_n10032_,
    new_n10033_, new_n10034_, new_n10035_, new_n10036_, new_n10037_,
    new_n10038_, new_n10039_, new_n10040_, new_n10041_, new_n10042_,
    new_n10043_, new_n10044_, new_n10045_, new_n10046_, new_n10047_,
    new_n10048_, new_n10049_, new_n10050_, new_n10051_, new_n10052_,
    new_n10053_, new_n10054_, new_n10055_, new_n10056_, new_n10057_,
    new_n10058_, new_n10059_, new_n10060_, new_n10061_, new_n10062_,
    new_n10063_, new_n10064_, new_n10065_, new_n10066_, new_n10067_,
    new_n10068_, new_n10069_, new_n10070_, new_n10071_, new_n10072_,
    new_n10073_, new_n10074_, new_n10075_, new_n10076_, new_n10077_,
    new_n10078_, new_n10079_, new_n10080_, new_n10081_, new_n10082_,
    new_n10083_, new_n10084_, new_n10085_, new_n10086_, new_n10087_,
    new_n10088_, new_n10089_, new_n10090_, new_n10091_, new_n10092_,
    new_n10093_, new_n10094_, new_n10095_, new_n10096_, new_n10097_,
    new_n10098_, new_n10099_, new_n10100_, new_n10101_, new_n10102_,
    new_n10103_, new_n10104_, new_n10105_, new_n10106_, new_n10107_,
    new_n10108_, new_n10109_, new_n10110_, new_n10111_, new_n10112_,
    new_n10113_, new_n10114_, new_n10115_, new_n10116_, new_n10117_,
    new_n10118_, new_n10119_, new_n10120_, new_n10121_, new_n10122_,
    new_n10123_, new_n10124_, new_n10125_, new_n10126_, new_n10127_,
    new_n10128_, new_n10129_, new_n10130_, new_n10131_, new_n10132_,
    new_n10133_, new_n10134_, new_n10135_, new_n10136_, new_n10137_,
    new_n10138_, new_n10139_, new_n10140_, new_n10141_, new_n10142_,
    new_n10143_, new_n10144_, new_n10145_, new_n10146_, new_n10147_,
    new_n10148_, new_n10149_, new_n10150_, new_n10151_, new_n10152_,
    new_n10153_, new_n10154_, new_n10155_, new_n10156_, new_n10157_,
    new_n10158_, new_n10159_, new_n10160_, new_n10161_, new_n10162_,
    new_n10163_, new_n10164_, new_n10165_, new_n10166_, new_n10167_,
    new_n10168_, new_n10169_, new_n10170_, new_n10171_, new_n10172_,
    new_n10173_, new_n10174_, new_n10175_, new_n10176_, new_n10177_,
    new_n10178_, new_n10179_, new_n10180_, new_n10181_, new_n10182_,
    new_n10183_, new_n10184_, new_n10185_, new_n10186_, new_n10187_,
    new_n10188_, new_n10189_, new_n10190_, new_n10191_, new_n10192_,
    new_n10193_, new_n10194_, new_n10195_, new_n10196_, new_n10197_,
    new_n10198_, new_n10199_, new_n10200_, new_n10201_, new_n10202_,
    new_n10203_, new_n10204_, new_n10205_, new_n10206_, new_n10207_,
    new_n10208_, new_n10209_, new_n10210_, new_n10211_, new_n10212_,
    new_n10213_, new_n10214_, new_n10215_, new_n10216_, new_n10217_,
    new_n10218_, new_n10219_, new_n10220_, new_n10221_, new_n10222_,
    new_n10223_, new_n10224_, new_n10225_, new_n10226_, new_n10227_,
    new_n10228_, new_n10229_, new_n10230_, new_n10231_, new_n10232_,
    new_n10233_, new_n10234_, new_n10235_, new_n10236_, new_n10237_,
    new_n10238_, new_n10239_, new_n10240_, new_n10241_, new_n10242_,
    new_n10243_, new_n10244_, new_n10245_, new_n10246_, new_n10247_,
    new_n10248_, new_n10249_, new_n10250_, new_n10251_, new_n10252_,
    new_n10253_, new_n10254_, new_n10255_, new_n10256_, new_n10257_,
    new_n10258_, new_n10259_, new_n10260_, new_n10261_, new_n10262_,
    new_n10263_, new_n10264_, new_n10265_, new_n10266_, new_n10267_,
    new_n10268_, new_n10269_, new_n10270_, new_n10271_, new_n10272_,
    new_n10273_, new_n10274_, new_n10275_, new_n10276_, new_n10277_,
    new_n10278_, new_n10279_, new_n10280_, new_n10281_, new_n10282_,
    new_n10283_, new_n10284_, new_n10285_, new_n10286_, new_n10287_,
    new_n10288_, new_n10289_, new_n10290_, new_n10291_, new_n10292_,
    new_n10293_, new_n10294_, new_n10295_, new_n10296_, new_n10297_,
    new_n10298_, new_n10299_, new_n10300_, new_n10301_, new_n10302_,
    new_n10303_, new_n10304_, new_n10305_, new_n10306_, new_n10307_,
    new_n10308_, new_n10309_, new_n10310_, new_n10311_, new_n10312_,
    new_n10313_, new_n10314_, new_n10315_, new_n10316_, new_n10317_,
    new_n10318_, new_n10319_, new_n10320_, new_n10321_, new_n10322_,
    new_n10323_, new_n10324_, new_n10325_, new_n10326_, new_n10327_,
    new_n10328_, new_n10329_, new_n10330_, new_n10331_, new_n10332_,
    new_n10333_, new_n10334_, new_n10335_, new_n10336_, new_n10337_,
    new_n10338_, new_n10339_, new_n10340_, new_n10341_, new_n10342_,
    new_n10343_, new_n10344_, new_n10345_, new_n10346_, new_n10347_,
    new_n10348_, new_n10349_, new_n10350_, new_n10351_, new_n10352_,
    new_n10353_, new_n10354_, new_n10355_, new_n10356_, new_n10357_,
    new_n10358_, new_n10359_, new_n10360_, new_n10361_, new_n10362_,
    new_n10363_, new_n10364_, new_n10365_, new_n10366_, new_n10367_,
    new_n10368_, new_n10369_, new_n10370_, new_n10371_, new_n10372_,
    new_n10373_, new_n10374_, new_n10375_, new_n10376_, new_n10377_,
    new_n10378_, new_n10379_, new_n10380_, new_n10381_, new_n10382_,
    new_n10383_, new_n10384_, new_n10385_, new_n10386_, new_n10387_,
    new_n10388_, new_n10389_, new_n10390_, new_n10391_, new_n10392_,
    new_n10393_, new_n10394_, new_n10395_, new_n10396_, new_n10397_,
    new_n10398_, new_n10399_, new_n10400_, new_n10401_, new_n10402_,
    new_n10403_, new_n10404_, new_n10405_, new_n10406_, new_n10407_,
    new_n10408_, new_n10409_, new_n10410_, new_n10411_, n2491_li, n2575_li,
    n2587_li, n2599_li, n2611_li, n2623_li, n2635_li, n2647_li, n2659_li,
    n2671_li, n2683_li, n2734_li, n2746_li, n2758_li, n2770_li, n2782_li,
    n2785_li, n2794_li, n2797_li, n2806_li, n2809_li, n2818_li, n2821_li,
    n2830_li, n2833_li, n2836_li, n2839_li, n2842_li, n2845_li, n2848_li,
    n2851_li, n2854_li, n2857_li, n2860_li, n2863_li, n4871_i2, n4893_i2,
    n4938_i2, n5056_i2, n5100_i2, n5122_i2, n5254_i2, n5276_i2, n5316_i2,
    n5434_i2, n5473_i2, n5494_i2, n5620_i2, n5643_i2, n5682_i2, n5798_i2,
    n5839_i2, n5867_i2, n6052_i2, n6087_i2, n6153_i2, n6408_i2, n6454_i2,
    n6509_i2, n6775_i2, n6818_i2, n6892_i2, n5779_i2, n5780_i2, n7156_i2,
    n5792_i2, n7205_i2, n5842_i2, n5863_i2, n7263_i2, n5881_i2, n5930_i2,
    n5959_i2, n5981_i2, n6042_i2, n6075_i2, n6103_i2, n7610_i2, n6169_i2,
    n7665_i2, n6205_i2, n6239_i2, n7788_i2, n6309_i2, n6461_i2, n6476_i2,
    n6521_i2, n6545_i2, G578_i2, G5106_i2, n6713_i2, G5164_i2, n6771_i2,
    n6810_i2, n6973_i2, n6995_i2, n7053_i2, G581_i2, G5467_i2, n7231_i2,
    G5527_i2, n7277_i2, n7304_i2, n7530_i2, n7595_i2, n7653_i2, G584_i2,
    G5820_i2, n7148_i2, n7149_i2, n7224_i2, n7916_i2, G5868_i2, n7958_i2,
    n7280_i2, n7313_i2, n8056_i2, n7323_i2, n7398_i2, n7459_i2, n7501_i2,
    n7518_i2, G563_i2, n7606_i2, G3358_i2, n7675_i2, G3410_i2, n7722_i2,
    n7747_i2, n7835_i2, G587_i2, G6046_i2, n7909_i2, G566_i2, G6070_i2,
    G3698_i2, n8086_i2, n8093_i2, G3752_i2, n8156_i2, n8199_i2,
    n2800_lo_buf_i2, G548_i2, G1715_i2, G569_i2, G1761_i2, G4043_i2,
    G4101_i2, G551_i2, G2034_i2, G4743_i2, G5271_i2, G5790_i2, G6122_i2,
    G2082_i2, n2812_lo_buf_i2, n2668_lo_buf_i2, n2680_lo_buf_i2, G572_i2,
    G6125_i2, G4395_i2, n2656_lo_buf_i2, G554_i2, G4452_i2, G2358_i2,
    n2644_lo_buf_i2, G2410_i2, n2632_lo_buf_i2, n2620_lo_buf_i2, G6131_i2,
    G4693_i2, G5209_i2, G5741_i2, G6082_i2, G6119_i2, n2608_lo_buf_i2,
    n2596_lo_buf_i2, n2584_lo_buf_i2, n2572_lo_buf_i2, n2704_lo_buf_i2,
    G557_i2, G5936_i2, G5442_i2, G4926_i2, G6134_i2, G3929_i2, G4425_i2,
    G4947_i2, n2764_lo_buf_i2, G2689_i2, n2560_lo_buf_i2, n2824_lo_buf_i2,
    G575_i2, G2740_i2, G4749_i2, n2548_lo_buf_i2, n2536_lo_buf_i2,
    n2524_lo_buf_i2, G875_i2, G1064_i2, G1253_i2, G6140_i2, G5151_i2,
    G5686_i2, G6061_i2, G4803_i2, G5332_i2, G5844_i2, G6114_i2, G4806_i2,
    G3881_i2, G4370_i2, G4896_i2, G5001_i2, G3121_i2, n2512_lo_buf_i2,
    G4085_i2, G4605_i2, G5118_i2, G4997_i2, n2500_lo_buf_i2,
    n2716_lo_buf_i2, G560_i2, G1895_i2, G3064_i2, G3269_i2, G3569_i2,
    G3022_i2, G1196_i2, G1007_i2, G818_i2, G674_i2, G5041_i2, G5562_i2,
    G6005_i2, G5214_i2, G5746_i2, G6087_i2, G6086_i2, G5745_i2, G5213_i2,
    G5893_i2, G5391_i2, G4864_i2, G6143_i2, G6008_i2, G5565_i2, G5044_i2,
    G3813_i2, G4325_i2, G4834_i2, G4993_i2, G3989_i2, G4490_i2, G5011_i2,
    G5112_i2, n2776_lo_buf_i2, G3298_i2, G3073_i2, G3265_i2, G3624_i2,
    G1642_i2, G1980_i2, n2488_lo_buf_i2, G626_i2, G1139_i2, G950_i2,
    G707_i2, G545_i2, G4217_i2, G4716_i2, G5244_i2, G3136_i2, G3499_i2,
    G3885_i2, G5243_i2, G3886_i2, G4375_i2, G4901_i2, G5054_i2, G4374_i2,
    G4900_i2, G5053_i2, G5242_i2, G4034_i2, G4556_i2, G5064_i2, G5172_i2,
    G2030_i2, G3016_i2, G3520_i2, G3261_i2, G3620_i2, G4220_i2, G4719_i2,
    G5247_i2, G5109_i2, G1638_i2, G1976_i2, G3560_i2, G3205_i2, G3193_i2,
    G3367_i2, G3670_i2, G1400_i2, G1280_i2, G902_i2, G659_i2, G983_i2,
    G740_i2, G2917_i2, G3391_i2, G3494_i2, G1512_i2, G1854_i2, G2203_i2,
    G3493_i2, G3069_i2, G3574_i2, G3319_i2, G3667_i2, G3068_i2, G3573_i2,
    G3666_i2, G3318_i2, G3492_i2, G3241_i2, G3722_i2, G3422_i2, G1445_i2,
    G3257_i2, G3616_i2, G1634_i2, G1972_i2, G2256_i2, G3394_i2, G3557_i2,
    G3364_i2, G3719_i2, G2253_i2, G1583_i2, G1917_i2, G1727_i2, G2061_i2,
    G935_i2, G692_i2, G2136_i2, G1507_i2, G1849_i2, G2198_i2, G2197_i2,
    G1848_i2, G1689_i2, G2016_i2, G2314_i2, G2313_i2, G1688_i2, G2015_i2,
    G1847_i2, G2196_i2, G2118_i2, G1777_i2, G1630_i2, G1968_i2, G2309_i2,
    G2139_i2, G1580_i2, G2250_i2, G1914_i2, G1724_i2, G2058_i2,
    n2728_lo_buf_i2;
  assign new_n809_ = G1;
  assign new_n810_ = ~G1;
  assign new_n811_ = G2;
  assign new_n812_ = ~G2;
  assign new_n813_ = G3;
  assign new_n814_ = ~G3;
  assign new_n815_ = G4;
  assign new_n816_ = ~G4;
  assign new_n817_ = G5;
  assign new_n818_ = ~G5;
  assign new_n819_ = G6;
  assign new_n820_ = ~G6;
  assign new_n821_ = G7;
  assign new_n822_ = ~G7;
  assign new_n823_ = G8;
  assign new_n824_ = ~G8;
  assign new_n825_ = G9;
  assign new_n826_ = ~G9;
  assign new_n827_ = G10;
  assign new_n828_ = ~G10;
  assign new_n829_ = G11;
  assign new_n830_ = ~G11;
  assign new_n831_ = G12;
  assign new_n832_ = ~G12;
  assign new_n833_ = G13;
  assign new_n834_ = ~G13;
  assign new_n835_ = G14;
  assign new_n836_ = ~G14;
  assign new_n837_ = G15;
  assign new_n838_ = ~G15;
  assign new_n839_ = G16;
  assign new_n840_ = ~G16;
  assign new_n841_ = G17;
  assign new_n842_ = ~G17;
  assign new_n843_ = G18;
  assign new_n844_ = ~G18;
  assign new_n845_ = G19;
  assign new_n846_ = ~G19;
  assign new_n847_ = G20;
  assign new_n848_ = ~G20;
  assign new_n849_ = G21;
  assign new_n851_ = G22;
  assign new_n853_ = G23;
  assign new_n855_ = G24;
  assign new_n857_ = G25;
  assign new_n859_ = G26;
  assign new_n861_ = G27;
  assign new_n863_ = G28;
  assign new_n865_ = G29;
  assign new_n867_ = G30;
  assign new_n869_ = G31;
  assign new_n871_ = G32;
  assign new_n873_ = n2491_lo;
  assign new_n875_ = n2575_lo;
  assign new_n876_ = ~n2575_lo;
  assign new_n877_ = n2587_lo;
  assign new_n878_ = ~n2587_lo;
  assign new_n879_ = n2599_lo;
  assign new_n880_ = ~n2599_lo;
  assign new_n881_ = n2611_lo;
  assign new_n882_ = ~n2611_lo;
  assign new_n883_ = n2623_lo;
  assign new_n884_ = ~n2623_lo;
  assign new_n885_ = n2635_lo;
  assign new_n886_ = ~n2635_lo;
  assign new_n887_ = n2647_lo;
  assign new_n888_ = ~n2647_lo;
  assign new_n889_ = n2659_lo;
  assign new_n890_ = ~n2659_lo;
  assign new_n891_ = n2671_lo;
  assign new_n892_ = ~n2671_lo;
  assign new_n893_ = n2683_lo;
  assign new_n895_ = n2734_lo;
  assign new_n896_ = ~n2734_lo;
  assign new_n897_ = n2746_lo;
  assign new_n898_ = ~n2746_lo;
  assign new_n899_ = n2758_lo;
  assign new_n900_ = ~n2758_lo;
  assign new_n901_ = n2770_lo;
  assign new_n902_ = ~n2770_lo;
  assign new_n903_ = n2782_lo;
  assign new_n905_ = n2785_lo;
  assign new_n906_ = ~n2785_lo;
  assign new_n907_ = n2794_lo;
  assign new_n909_ = n2797_lo;
  assign new_n910_ = ~n2797_lo;
  assign new_n911_ = n2806_lo;
  assign new_n913_ = n2809_lo;
  assign new_n914_ = ~n2809_lo;
  assign new_n915_ = n2818_lo;
  assign new_n917_ = n2821_lo;
  assign new_n918_ = ~n2821_lo;
  assign new_n919_ = n2830_lo;
  assign new_n921_ = n2833_lo;
  assign new_n923_ = n2836_lo;
  assign new_n924_ = ~n2836_lo;
  assign new_n925_ = n2839_lo;
  assign new_n926_ = ~n2839_lo;
  assign new_n927_ = n2842_lo;
  assign new_n929_ = n2845_lo;
  assign new_n931_ = n2848_lo;
  assign new_n932_ = ~n2848_lo;
  assign new_n933_ = n2851_lo;
  assign new_n934_ = ~n2851_lo;
  assign new_n935_ = n2854_lo;
  assign new_n937_ = n2857_lo;
  assign new_n939_ = n2860_lo;
  assign new_n940_ = ~n2860_lo;
  assign new_n941_ = n2863_lo;
  assign new_n942_ = ~n2863_lo;
  assign new_n943_ = n4871_o2;
  assign new_n946_ = ~n4893_o2;
  assign new_n947_ = n4938_o2;
  assign new_n949_ = n5056_o2;
  assign new_n952_ = ~n5100_o2;
  assign new_n953_ = n5122_o2;
  assign new_n955_ = n5254_o2;
  assign new_n958_ = ~n5276_o2;
  assign new_n959_ = n5316_o2;
  assign new_n961_ = n5434_o2;
  assign new_n964_ = ~n5473_o2;
  assign new_n965_ = n5494_o2;
  assign new_n967_ = n5620_o2;
  assign new_n970_ = ~n5643_o2;
  assign new_n971_ = n5682_o2;
  assign new_n973_ = n5798_o2;
  assign new_n976_ = ~n5839_o2;
  assign new_n977_ = n5867_o2;
  assign new_n979_ = n6052_o2;
  assign new_n982_ = ~n6087_o2;
  assign new_n983_ = n6153_o2;
  assign new_n985_ = n6408_o2;
  assign new_n988_ = ~n6454_o2;
  assign new_n989_ = n6509_o2;
  assign new_n991_ = n6775_o2;
  assign new_n994_ = ~n6818_o2;
  assign new_n995_ = n6892_o2;
  assign new_n997_ = n5779_o2;
  assign new_n998_ = ~n5779_o2;
  assign new_n999_ = n5780_o2;
  assign new_n1001_ = n7156_o2;
  assign new_n1003_ = n5792_o2;
  assign new_n1004_ = ~n5792_o2;
  assign new_n1006_ = ~n7205_o2;
  assign new_n1007_ = n5842_o2;
  assign new_n1008_ = ~n5842_o2;
  assign new_n1009_ = n5863_o2;
  assign new_n1010_ = ~n5863_o2;
  assign new_n1011_ = n7263_o2;
  assign new_n1013_ = n5881_o2;
  assign new_n1014_ = ~n5881_o2;
  assign new_n1015_ = n5930_o2;
  assign new_n1016_ = ~n5930_o2;
  assign new_n1017_ = n5959_o2;
  assign new_n1018_ = ~n5959_o2;
  assign new_n1019_ = n5981_o2;
  assign new_n1020_ = ~n5981_o2;
  assign new_n1021_ = n6042_o2;
  assign new_n1022_ = ~n6042_o2;
  assign new_n1023_ = n6075_o2;
  assign new_n1024_ = ~n6075_o2;
  assign new_n1025_ = n6103_o2;
  assign new_n1026_ = ~n6103_o2;
  assign new_n1027_ = n7610_o2;
  assign new_n1029_ = n6169_o2;
  assign new_n1030_ = ~n6169_o2;
  assign new_n1032_ = ~n7665_o2;
  assign new_n1033_ = n6205_o2;
  assign new_n1034_ = ~n6205_o2;
  assign new_n1035_ = n6239_o2;
  assign new_n1036_ = ~n6239_o2;
  assign new_n1037_ = n7788_o2;
  assign new_n1039_ = n6309_o2;
  assign new_n1040_ = ~n6309_o2;
  assign new_n1041_ = n6461_o2;
  assign new_n1042_ = ~n6461_o2;
  assign new_n1043_ = n6476_o2;
  assign new_n1045_ = n325_inv;
  assign new_n1047_ = n6545_o2;
  assign new_n1049_ = G578_o2;
  assign new_n1052_ = ~G5106_o2;
  assign new_n1053_ = n6713_o2;
  assign new_n1055_ = G5164_o2;
  assign new_n1057_ = n343_inv;
  assign new_n1059_ = n6810_o2;
  assign new_n1061_ = n6973_o2;
  assign new_n1063_ = n352_inv;
  assign new_n1065_ = n7053_o2;
  assign new_n1067_ = G581_o2;
  assign new_n1070_ = ~G5467_o2;
  assign new_n1071_ = n7231_o2;
  assign new_n1073_ = G5527_o2;
  assign new_n1075_ = n370_inv;
  assign new_n1077_ = n7304_o2;
  assign new_n1079_ = n7530_o2;
  assign new_n1081_ = n379_inv;
  assign new_n1083_ = n7653_o2;
  assign new_n1085_ = G584_o2;
  assign new_n1088_ = ~G5820_o2;
  assign new_n1089_ = n7148_o2;
  assign new_n1090_ = ~n7148_o2;
  assign new_n1091_ = n7149_o2;
  assign new_n1093_ = n7224_o2;
  assign new_n1094_ = ~n7224_o2;
  assign new_n1095_ = n7916_o2;
  assign new_n1097_ = G5868_o2;
  assign new_n1099_ = n406_inv;
  assign new_n1101_ = n7280_o2;
  assign new_n1102_ = ~n7280_o2;
  assign new_n1103_ = n7313_o2;
  assign new_n1104_ = ~n7313_o2;
  assign new_n1105_ = n8056_o2;
  assign new_n1107_ = n7323_o2;
  assign new_n1108_ = ~n7323_o2;
  assign new_n1109_ = n7398_o2;
  assign new_n1110_ = ~n7398_o2;
  assign new_n1111_ = n7459_o2;
  assign new_n1112_ = ~n7459_o2;
  assign new_n1113_ = n7501_o2;
  assign new_n1114_ = ~n7501_o2;
  assign new_n1115_ = n7518_o2;
  assign new_n1116_ = ~n7518_o2;
  assign new_n1117_ = G563_o2;
  assign new_n1119_ = n7606_o2;
  assign new_n1120_ = ~n7606_o2;
  assign new_n1121_ = n439_inv;
  assign new_n1123_ = n7675_o2;
  assign new_n1124_ = ~n7675_o2;
  assign new_n1125_ = G3410_o2;
  assign new_n1127_ = n7722_o2;
  assign new_n1128_ = ~n7722_o2;
  assign new_n1129_ = n7747_o2;
  assign new_n1130_ = ~n7747_o2;
  assign new_n1131_ = n7835_o2;
  assign new_n1132_ = ~n7835_o2;
  assign new_n1133_ = G587_o2;
  assign new_n1136_ = ~G6046_o2;
  assign new_n1137_ = n7909_o2;
  assign new_n1138_ = ~n7909_o2;
  assign new_n1139_ = G566_o2;
  assign new_n1141_ = G6070_o2;
  assign new_n1143_ = n472_inv;
  assign new_n1145_ = n8086_o2;
  assign new_n1146_ = ~n8086_o2;
  assign new_n1147_ = n8093_o2;
  assign new_n1149_ = G3752_o2;
  assign new_n1151_ = n484_inv;
  assign new_n1153_ = n8199_o2;
  assign new_n1155_ = n2800_lo_buf_o2;
  assign new_n1156_ = ~n2800_lo_buf_o2;
  assign new_n1157_ = G548_o2;
  assign new_n1159_ = n496_inv;
  assign new_n1161_ = G569_o2;
  assign new_n1163_ = G1761_o2;
  assign new_n1165_ = n505_inv;
  assign new_n1167_ = G4101_o2;
  assign new_n1169_ = G551_o2;
  assign new_n1171_ = n514_inv;
  assign new_n1173_ = G4743_o2;
  assign new_n1174_ = ~G4743_o2;
  assign new_n1175_ = G5271_o2;
  assign new_n1176_ = ~G5271_o2;
  assign new_n1177_ = G5790_o2;
  assign new_n1178_ = ~G5790_o2;
  assign new_n1180_ = ~G6122_o2;
  assign new_n1181_ = G2082_o2;
  assign new_n1183_ = n2812_lo_buf_o2;
  assign new_n1184_ = ~n2812_lo_buf_o2;
  assign new_n1185_ = n2668_lo_buf_o2;
  assign new_n1186_ = ~n2668_lo_buf_o2;
  assign new_n1187_ = n2680_lo_buf_o2;
  assign new_n1189_ = G572_o2;
  assign new_n1191_ = G6125_o2;
  assign new_n1193_ = n547_inv;
  assign new_n1195_ = n2656_lo_buf_o2;
  assign new_n1196_ = ~n2656_lo_buf_o2;
  assign new_n1197_ = G554_o2;
  assign new_n1199_ = G4452_o2;
  assign new_n1201_ = n559_inv;
  assign new_n1203_ = n2644_lo_buf_o2;
  assign new_n1204_ = ~n2644_lo_buf_o2;
  assign new_n1205_ = G2410_o2;
  assign new_n1207_ = n2632_lo_buf_o2;
  assign new_n1208_ = ~n2632_lo_buf_o2;
  assign new_n1209_ = n2620_lo_buf_o2;
  assign new_n1210_ = ~n2620_lo_buf_o2;
  assign new_n1211_ = G6131_o2;
  assign new_n1213_ = G4693_o2;
  assign new_n1214_ = ~G4693_o2;
  assign new_n1215_ = G5209_o2;
  assign new_n1216_ = ~G5209_o2;
  assign new_n1217_ = G5741_o2;
  assign new_n1218_ = ~G5741_o2;
  assign new_n1219_ = G6082_o2;
  assign new_n1220_ = ~G6082_o2;
  assign new_n1222_ = ~G6119_o2;
  assign new_n1223_ = n2608_lo_buf_o2;
  assign new_n1224_ = ~n2608_lo_buf_o2;
  assign new_n1225_ = n2596_lo_buf_o2;
  assign new_n1226_ = ~n2596_lo_buf_o2;
  assign new_n1227_ = n2584_lo_buf_o2;
  assign new_n1228_ = ~n2584_lo_buf_o2;
  assign new_n1229_ = n2572_lo_buf_o2;
  assign new_n1230_ = ~n2572_lo_buf_o2;
  assign new_n1231_ = n2704_lo_buf_o2;
  assign new_n1232_ = ~n2704_lo_buf_o2;
  assign new_n1233_ = G557_o2;
  assign new_n1235_ = G5936_o2;
  assign new_n1236_ = ~G5936_o2;
  assign new_n1237_ = G5442_o2;
  assign new_n1238_ = ~G5442_o2;
  assign new_n1239_ = G4926_o2;
  assign new_n1240_ = ~G4926_o2;
  assign new_n1241_ = G6134_o2;
  assign new_n1243_ = G3929_o2;
  assign new_n1244_ = ~G3929_o2;
  assign new_n1245_ = G4425_o2;
  assign new_n1246_ = ~G4425_o2;
  assign new_n1247_ = G4947_o2;
  assign new_n1248_ = ~G4947_o2;
  assign new_n1249_ = n2764_lo_buf_o2;
  assign new_n1250_ = ~n2764_lo_buf_o2;
  assign new_n1251_ = n634_inv;
  assign new_n1253_ = n2560_lo_buf_o2;
  assign new_n1254_ = ~n2560_lo_buf_o2;
  assign new_n1255_ = n2824_lo_buf_o2;
  assign new_n1256_ = ~n2824_lo_buf_o2;
  assign new_n1257_ = G575_o2;
  assign new_n1259_ = G2740_o2;
  assign new_n1261_ = n649_inv;
  assign new_n1263_ = n2548_lo_buf_o2;
  assign new_n1264_ = ~n2548_lo_buf_o2;
  assign new_n1265_ = n2536_lo_buf_o2;
  assign new_n1266_ = ~n2536_lo_buf_o2;
  assign new_n1267_ = n2524_lo_buf_o2;
  assign new_n1268_ = ~n2524_lo_buf_o2;
  assign new_n1269_ = G875_o2;
  assign new_n1270_ = ~G875_o2;
  assign new_n1271_ = G1064_o2;
  assign new_n1272_ = ~G1064_o2;
  assign new_n1273_ = G1253_o2;
  assign new_n1274_ = ~G1253_o2;
  assign new_n1275_ = G6140_o2;
  assign new_n1277_ = G5151_o2;
  assign new_n1278_ = ~G5151_o2;
  assign new_n1279_ = G5686_o2;
  assign new_n1280_ = ~G5686_o2;
  assign new_n1281_ = G6061_o2;
  assign new_n1282_ = ~G6061_o2;
  assign new_n1283_ = G4803_o2;
  assign new_n1284_ = ~G4803_o2;
  assign new_n1285_ = G5332_o2;
  assign new_n1286_ = ~G5332_o2;
  assign new_n1287_ = G5844_o2;
  assign new_n1288_ = ~G5844_o2;
  assign new_n1290_ = ~G6114_o2;
  assign new_n1291_ = G4806_o2;
  assign new_n1293_ = G3881_o2;
  assign new_n1294_ = ~G3881_o2;
  assign new_n1295_ = G4370_o2;
  assign new_n1296_ = ~G4370_o2;
  assign new_n1297_ = G4896_o2;
  assign new_n1298_ = ~G4896_o2;
  assign new_n1299_ = G5001_o2;
  assign new_n1300_ = ~G5001_o2;
  assign new_n1301_ = G3121_o2;
  assign new_n1302_ = ~G3121_o2;
  assign new_n1303_ = n2512_lo_buf_o2;
  assign new_n1304_ = ~n2512_lo_buf_o2;
  assign new_n1305_ = G4085_o2;
  assign new_n1306_ = ~G4085_o2;
  assign new_n1307_ = G4605_o2;
  assign new_n1308_ = ~G4605_o2;
  assign new_n1309_ = G5118_o2;
  assign new_n1310_ = ~G5118_o2;
  assign new_n1311_ = G4997_o2;
  assign new_n1312_ = ~G4997_o2;
  assign new_n1313_ = n2500_lo_buf_o2;
  assign new_n1314_ = ~n2500_lo_buf_o2;
  assign new_n1315_ = n2716_lo_buf_o2;
  assign new_n1316_ = ~n2716_lo_buf_o2;
  assign new_n1317_ = G560_o2;
  assign new_n1319_ = G1895_o2;
  assign new_n1320_ = ~G1895_o2;
  assign new_n1321_ = G3064_o2;
  assign new_n1322_ = ~G3064_o2;
  assign new_n1323_ = G3269_o2;
  assign new_n1324_ = ~G3269_o2;
  assign new_n1325_ = G3569_o2;
  assign new_n1326_ = ~G3569_o2;
  assign new_n1327_ = n748_inv;
  assign new_n1329_ = G1196_o2;
  assign new_n1330_ = ~G1196_o2;
  assign new_n1331_ = G1007_o2;
  assign new_n1332_ = ~G1007_o2;
  assign new_n1333_ = G818_o2;
  assign new_n1334_ = ~G818_o2;
  assign new_n1335_ = G674_o2;
  assign new_n1336_ = ~G674_o2;
  assign new_n1337_ = G5041_o2;
  assign new_n1338_ = ~G5041_o2;
  assign new_n1339_ = G5562_o2;
  assign new_n1340_ = ~G5562_o2;
  assign new_n1341_ = G6005_o2;
  assign new_n1342_ = ~G6005_o2;
  assign new_n1343_ = G5214_o2;
  assign new_n1344_ = ~G5214_o2;
  assign new_n1345_ = G5746_o2;
  assign new_n1346_ = ~G5746_o2;
  assign new_n1347_ = G6087_o2;
  assign new_n1348_ = ~G6087_o2;
  assign new_n1349_ = G6086_o2;
  assign new_n1350_ = ~G6086_o2;
  assign new_n1351_ = G5745_o2;
  assign new_n1352_ = ~G5745_o2;
  assign new_n1353_ = G5213_o2;
  assign new_n1354_ = ~G5213_o2;
  assign new_n1355_ = G5893_o2;
  assign new_n1356_ = ~G5893_o2;
  assign new_n1357_ = G5391_o2;
  assign new_n1358_ = ~G5391_o2;
  assign new_n1359_ = G4864_o2;
  assign new_n1360_ = ~G4864_o2;
  assign new_n1361_ = G6143_o2;
  assign new_n1362_ = ~G6143_o2;
  assign new_n1363_ = G6008_o2;
  assign new_n1364_ = ~G6008_o2;
  assign new_n1365_ = G5565_o2;
  assign new_n1366_ = ~G5565_o2;
  assign new_n1367_ = G5044_o2;
  assign new_n1368_ = ~G5044_o2;
  assign new_n1369_ = G3813_o2;
  assign new_n1370_ = ~G3813_o2;
  assign new_n1371_ = G4325_o2;
  assign new_n1372_ = ~G4325_o2;
  assign new_n1373_ = G4834_o2;
  assign new_n1374_ = ~G4834_o2;
  assign new_n1375_ = G4993_o2;
  assign new_n1376_ = ~G4993_o2;
  assign new_n1377_ = G3989_o2;
  assign new_n1378_ = ~G3989_o2;
  assign new_n1379_ = G4490_o2;
  assign new_n1380_ = ~G4490_o2;
  assign new_n1381_ = G5011_o2;
  assign new_n1382_ = ~G5011_o2;
  assign new_n1383_ = G5112_o2;
  assign new_n1384_ = ~G5112_o2;
  assign new_n1385_ = n2776_lo_buf_o2;
  assign new_n1386_ = ~n2776_lo_buf_o2;
  assign new_n1387_ = G3298_o2;
  assign new_n1388_ = ~G3298_o2;
  assign new_n1389_ = G3073_o2;
  assign new_n1391_ = G3265_o2;
  assign new_n1392_ = ~G3265_o2;
  assign new_n1393_ = G3624_o2;
  assign new_n1394_ = ~G3624_o2;
  assign new_n1395_ = G1642_o2;
  assign new_n1396_ = ~G1642_o2;
  assign new_n1397_ = G1980_o2;
  assign new_n1398_ = ~G1980_o2;
  assign new_n1399_ = n2488_lo_buf_o2;
  assign new_n1400_ = ~n2488_lo_buf_o2;
  assign new_n1401_ = G626_o2;
  assign new_n1402_ = ~G626_o2;
  assign new_n1403_ = G1139_o2;
  assign new_n1404_ = ~G1139_o2;
  assign new_n1405_ = G950_o2;
  assign new_n1406_ = ~G950_o2;
  assign new_n1407_ = G707_o2;
  assign new_n1408_ = ~G707_o2;
  assign new_n1409_ = G545_o2;
  assign new_n1411_ = G4217_o2;
  assign new_n1412_ = ~G4217_o2;
  assign new_n1413_ = G4716_o2;
  assign new_n1414_ = ~G4716_o2;
  assign new_n1415_ = G5244_o2;
  assign new_n1416_ = ~G5244_o2;
  assign new_n1417_ = G3136_o2;
  assign new_n1418_ = ~G3136_o2;
  assign new_n1419_ = G3499_o2;
  assign new_n1420_ = ~G3499_o2;
  assign new_n1421_ = G3885_o2;
  assign new_n1422_ = ~G3885_o2;
  assign new_n1423_ = G5243_o2;
  assign new_n1424_ = ~G5243_o2;
  assign new_n1425_ = G3886_o2;
  assign new_n1426_ = ~G3886_o2;
  assign new_n1427_ = G4375_o2;
  assign new_n1428_ = ~G4375_o2;
  assign new_n1429_ = G4901_o2;
  assign new_n1430_ = ~G4901_o2;
  assign new_n1431_ = G5054_o2;
  assign new_n1432_ = ~G5054_o2;
  assign new_n1433_ = G4374_o2;
  assign new_n1434_ = ~G4374_o2;
  assign new_n1435_ = G4900_o2;
  assign new_n1436_ = ~G4900_o2;
  assign new_n1437_ = G5053_o2;
  assign new_n1438_ = ~G5053_o2;
  assign new_n1439_ = G5242_o2;
  assign new_n1440_ = ~G5242_o2;
  assign new_n1441_ = G4034_o2;
  assign new_n1442_ = ~G4034_o2;
  assign new_n1443_ = G4556_o2;
  assign new_n1444_ = ~G4556_o2;
  assign new_n1445_ = G5064_o2;
  assign new_n1446_ = ~G5064_o2;
  assign new_n1447_ = G5172_o2;
  assign new_n1448_ = ~G5172_o2;
  assign new_n1449_ = G2030_o2;
  assign new_n1450_ = ~G2030_o2;
  assign new_n1451_ = G3016_o2;
  assign new_n1452_ = ~G3016_o2;
  assign new_n1453_ = G3520_o2;
  assign new_n1454_ = ~G3520_o2;
  assign new_n1455_ = G3261_o2;
  assign new_n1456_ = ~G3261_o2;
  assign new_n1457_ = G3620_o2;
  assign new_n1458_ = ~G3620_o2;
  assign new_n1459_ = G4220_o2;
  assign new_n1460_ = ~G4220_o2;
  assign new_n1461_ = G4719_o2;
  assign new_n1462_ = ~G4719_o2;
  assign new_n1463_ = G5247_o2;
  assign new_n1464_ = ~G5247_o2;
  assign new_n1465_ = G5109_o2;
  assign new_n1466_ = ~G5109_o2;
  assign new_n1467_ = G1638_o2;
  assign new_n1468_ = ~G1638_o2;
  assign new_n1469_ = G1976_o2;
  assign new_n1470_ = ~G1976_o2;
  assign new_n1471_ = G3560_o2;
  assign new_n1472_ = ~G3560_o2;
  assign new_n1473_ = G3205_o2;
  assign new_n1474_ = ~G3205_o2;
  assign new_n1475_ = G3193_o2;
  assign new_n1476_ = ~G3193_o2;
  assign new_n1477_ = G3367_o2;
  assign new_n1478_ = ~G3367_o2;
  assign new_n1479_ = G3670_o2;
  assign new_n1480_ = ~G3670_o2;
  assign new_n1481_ = n979_inv;
  assign new_n1483_ = G1280_o2;
  assign new_n1484_ = ~G1280_o2;
  assign new_n1485_ = G902_o2;
  assign new_n1486_ = ~G902_o2;
  assign new_n1487_ = G659_o2;
  assign new_n1488_ = ~G659_o2;
  assign new_n1489_ = G983_o2;
  assign new_n1490_ = ~G983_o2;
  assign new_n1491_ = G740_o2;
  assign new_n1492_ = ~G740_o2;
  assign new_n1493_ = G2917_o2;
  assign new_n1494_ = ~G2917_o2;
  assign new_n1495_ = G3391_o2;
  assign new_n1496_ = ~G3391_o2;
  assign new_n1497_ = G3494_o2;
  assign new_n1498_ = ~G3494_o2;
  assign new_n1499_ = G1512_o2;
  assign new_n1500_ = ~G1512_o2;
  assign new_n1501_ = G1854_o2;
  assign new_n1502_ = ~G1854_o2;
  assign new_n1503_ = G2203_o2;
  assign new_n1504_ = ~G2203_o2;
  assign new_n1505_ = G3493_o2;
  assign new_n1506_ = ~G3493_o2;
  assign new_n1507_ = G3069_o2;
  assign new_n1508_ = ~G3069_o2;
  assign new_n1509_ = G3574_o2;
  assign new_n1510_ = ~G3574_o2;
  assign new_n1511_ = G3319_o2;
  assign new_n1512_ = ~G3319_o2;
  assign new_n1513_ = G3667_o2;
  assign new_n1514_ = ~G3667_o2;
  assign new_n1515_ = G3068_o2;
  assign new_n1516_ = ~G3068_o2;
  assign new_n1517_ = G3573_o2;
  assign new_n1518_ = ~G3573_o2;
  assign new_n1519_ = G3666_o2;
  assign new_n1520_ = ~G3666_o2;
  assign new_n1521_ = G3318_o2;
  assign new_n1522_ = ~G3318_o2;
  assign new_n1523_ = G3492_o2;
  assign new_n1524_ = ~G3492_o2;
  assign new_n1525_ = G3241_o2;
  assign new_n1526_ = ~G3241_o2;
  assign new_n1527_ = G3722_o2;
  assign new_n1528_ = ~G3722_o2;
  assign new_n1529_ = G3422_o2;
  assign new_n1530_ = ~G3422_o2;
  assign new_n1531_ = G1445_o2;
  assign new_n1533_ = G3257_o2;
  assign new_n1534_ = ~G3257_o2;
  assign new_n1535_ = G3616_o2;
  assign new_n1536_ = ~G3616_o2;
  assign new_n1537_ = G1634_o2;
  assign new_n1538_ = ~G1634_o2;
  assign new_n1539_ = G1972_o2;
  assign new_n1540_ = ~G1972_o2;
  assign new_n1541_ = G2256_o2;
  assign new_n1542_ = ~G2256_o2;
  assign new_n1543_ = G3394_o2;
  assign new_n1544_ = ~G3394_o2;
  assign new_n1545_ = G3557_o2;
  assign new_n1546_ = ~G3557_o2;
  assign new_n1547_ = G3364_o2;
  assign new_n1548_ = ~G3364_o2;
  assign new_n1549_ = G3719_o2;
  assign new_n1550_ = ~G3719_o2;
  assign new_n1551_ = G2253_o2;
  assign new_n1552_ = ~G2253_o2;
  assign new_n1553_ = G1583_o2;
  assign new_n1554_ = ~G1583_o2;
  assign new_n1555_ = G1917_o2;
  assign new_n1556_ = ~G1917_o2;
  assign new_n1557_ = G1727_o2;
  assign new_n1558_ = ~G1727_o2;
  assign new_n1559_ = G2061_o2;
  assign new_n1560_ = ~G2061_o2;
  assign new_n1561_ = G935_o2;
  assign new_n1562_ = ~G935_o2;
  assign new_n1563_ = G692_o2;
  assign new_n1564_ = ~G692_o2;
  assign new_n1565_ = G2136_o2;
  assign new_n1566_ = ~G2136_o2;
  assign new_n1567_ = G1507_o2;
  assign new_n1568_ = ~G1507_o2;
  assign new_n1569_ = G1849_o2;
  assign new_n1570_ = ~G1849_o2;
  assign new_n1571_ = G2198_o2;
  assign new_n1572_ = ~G2198_o2;
  assign new_n1573_ = G2197_o2;
  assign new_n1574_ = ~G2197_o2;
  assign new_n1575_ = G1848_o2;
  assign new_n1576_ = ~G1848_o2;
  assign new_n1577_ = G1689_o2;
  assign new_n1578_ = ~G1689_o2;
  assign new_n1579_ = G2016_o2;
  assign new_n1580_ = ~G2016_o2;
  assign new_n1581_ = G2314_o2;
  assign new_n1582_ = ~G2314_o2;
  assign new_n1583_ = G2313_o2;
  assign new_n1584_ = ~G2313_o2;
  assign new_n1585_ = G1688_o2;
  assign new_n1586_ = ~G1688_o2;
  assign new_n1587_ = G2015_o2;
  assign new_n1588_ = ~G2015_o2;
  assign new_n1589_ = G1847_o2;
  assign new_n1590_ = ~G1847_o2;
  assign new_n1591_ = G2196_o2;
  assign new_n1592_ = ~G2196_o2;
  assign new_n1593_ = G2118_o2;
  assign new_n1594_ = ~G2118_o2;
  assign new_n1595_ = G1777_o2;
  assign new_n1596_ = ~G1777_o2;
  assign new_n1597_ = G1630_o2;
  assign new_n1598_ = ~G1630_o2;
  assign new_n1599_ = G1968_o2;
  assign new_n1600_ = ~G1968_o2;
  assign new_n1601_ = G2309_o2;
  assign new_n1602_ = ~G2309_o2;
  assign new_n1603_ = G2139_o2;
  assign new_n1604_ = ~G2139_o2;
  assign new_n1605_ = G1580_o2;
  assign new_n1606_ = ~G1580_o2;
  assign new_n1607_ = G2250_o2;
  assign new_n1608_ = ~G2250_o2;
  assign new_n1609_ = G1914_o2;
  assign new_n1610_ = ~G1914_o2;
  assign new_n1611_ = G1724_o2;
  assign new_n1612_ = ~G1724_o2;
  assign new_n1613_ = G2058_o2;
  assign new_n1614_ = ~G2058_o2;
  assign new_n1615_ = n2728_lo_buf_o2;
  assign new_n1616_ = ~n2728_lo_buf_o2;
  assign new_n1617_ = new_n893_ & new_n873_;
  assign new_n1618_ = new_n6352_ | new_n946_;
  assign new_n1619_ = new_n6352_ | new_n943_;
  assign new_n1620_ = new_n1619_ & new_n1618_;
  assign new_n1621_ = new_n6353_ | new_n952_;
  assign new_n1622_ = new_n6353_ | new_n949_;
  assign new_n1623_ = new_n1622_ & new_n1621_;
  assign new_n1624_ = new_n6354_ | new_n958_;
  assign new_n1625_ = new_n6354_ | new_n955_;
  assign new_n1626_ = new_n1625_ & new_n1624_;
  assign new_n1627_ = new_n6355_ | new_n964_;
  assign new_n1628_ = new_n6355_ | new_n961_;
  assign new_n1629_ = new_n1628_ & new_n1627_;
  assign new_n1630_ = new_n6356_ | new_n970_;
  assign new_n1631_ = new_n6356_ | new_n967_;
  assign new_n1632_ = new_n1631_ & new_n1630_;
  assign new_n1633_ = new_n6357_ | new_n976_;
  assign new_n1634_ = new_n6357_ | new_n973_;
  assign new_n1635_ = new_n1634_ & new_n1633_;
  assign new_n1636_ = new_n6358_ | new_n982_;
  assign new_n1637_ = new_n6358_ | new_n979_;
  assign new_n1638_ = new_n1637_ & new_n1636_;
  assign new_n1639_ = new_n6359_ | new_n988_;
  assign new_n1640_ = new_n6359_ | new_n985_;
  assign new_n1641_ = new_n1640_ & new_n1639_;
  assign new_n1642_ = new_n6360_ | new_n994_;
  assign new_n1643_ = new_n6360_ | new_n991_;
  assign new_n1644_ = new_n1643_ & new_n1642_;
  assign new_n1645_ = new_n6361_ | new_n1006_;
  assign new_n1646_ = new_n6361_ | new_n1001_;
  assign new_n1647_ = new_n1646_ & new_n1645_;
  assign new_n1648_ = new_n6362_ | new_n1032_;
  assign new_n1649_ = new_n6362_ | new_n1027_;
  assign new_n1650_ = new_n1649_ & new_n1648_;
  assign new_n1651_ = new_n6363_ | new_n1052_;
  assign new_n1652_ = new_n6363_ | new_n1049_;
  assign new_n1653_ = new_n1652_ & new_n1651_;
  assign new_n1654_ = new_n6364_ | new_n1070_;
  assign new_n1655_ = new_n6364_ | new_n1067_;
  assign new_n1656_ = new_n1655_ & new_n1654_;
  assign new_n1657_ = new_n6365_ | new_n1088_;
  assign new_n1658_ = new_n6365_ | new_n1085_;
  assign new_n1659_ = new_n1658_ & new_n1657_;
  assign new_n1660_ = new_n6366_ | new_n1136_;
  assign new_n1661_ = new_n6366_ | new_n1133_;
  assign new_n1662_ = new_n1661_ & new_n1660_;
  assign new_n1663_ = new_n6367_ | new_n1180_;
  assign new_n1664_ = new_n1663_ & new_n6367_;
  assign new_n1665_ = new_n6368_ | new_n1222_;
  assign new_n1666_ = new_n6368_ | new_n1211_;
  assign new_n1667_ = new_n1666_ & new_n1665_;
  assign new_n1668_ = new_n6370_ | new_n1290_;
  assign new_n1669_ = new_n6370_ | new_n1275_;
  assign new_n1670_ = new_n1669_ & new_n1668_;
  assign new_n1671_ = new_n1350_ & new_n1348_;
  assign new_n1672_ = new_n1349_ | new_n1347_;
  assign new_n1673_ = new_n1362_ & new_n1219_;
  assign new_n1674_ = new_n6369_ | new_n1220_;
  assign new_n1675_ = new_n1674_ & new_n1672_;
  assign new_n1676_ = new_n6371_ | new_n6372_;
  assign new_n1677_ = new_n6374_ | new_n6372_;
  assign new_n1678_ = new_n6374_ | new_n6371_;
  assign new_n1679_ = new_n1678_ & new_n1677_;
  assign new_n1680_ = new_n6375_ & new_n6376_;
  assign new_n1681_ = new_n6377_ | new_n6378_;
  assign new_n1682_ = new_n6380_ & new_n6375_;
  assign new_n1683_ = new_n6382_ | new_n6377_;
  assign new_n1684_ = new_n6380_ & new_n6376_;
  assign new_n1685_ = new_n6382_ | new_n6378_;
  assign new_n1686_ = new_n1685_ & new_n1683_;
  assign new_n1687_ = new_n1684_ | new_n1682_;
  assign new_n1688_ = new_n1676_ & new_n1281_;
  assign new_n1689_ = new_n6373_ | new_n1282_;
  assign new_n1690_ = new_n1689_ & new_n1687_;
  assign new_n1691_ = new_n6383_ | new_n6384_;
  assign new_n1692_ = new_n6386_ | new_n6384_;
  assign new_n1693_ = new_n6386_ | new_n6383_;
  assign new_n1694_ = new_n1693_ & new_n1692_;
  assign new_n1695_ = new_n6388_ & new_n1287_;
  assign new_n1696_ = new_n6390_ | new_n1288_;
  assign new_n1697_ = new_n6388_ & new_n1270_;
  assign new_n1698_ = new_n6390_ | new_n1269_;
  assign new_n1699_ = new_n1698_ & new_n1696_;
  assign new_n1700_ = new_n1697_ | new_n1695_;
  assign new_n1701_ = new_n1236_ & new_n1177_;
  assign new_n1702_ = new_n1235_ | new_n1178_;
  assign new_n1703_ = new_n6391_ & new_n6392_;
  assign new_n1704_ = new_n6393_ | new_n6394_;
  assign new_n1705_ = new_n6396_ & new_n6392_;
  assign new_n1706_ = new_n6398_ | new_n6394_;
  assign new_n1707_ = new_n6396_ & new_n6391_;
  assign new_n1708_ = new_n6398_ | new_n6393_;
  assign new_n1709_ = new_n1708_ & new_n1706_;
  assign new_n1710_ = new_n1707_ | new_n1705_;
  assign new_n1711_ = new_n1691_ & new_n6379_;
  assign new_n1712_ = new_n6385_ | new_n6381_;
  assign new_n1713_ = new_n1712_ & new_n1710_;
  assign new_n1714_ = new_n6399_ | new_n6400_;
  assign new_n1715_ = new_n6402_ | new_n6400_;
  assign new_n1716_ = new_n6402_ | new_n6399_;
  assign new_n1717_ = new_n1716_ & new_n1715_;
  assign new_n1718_ = new_n1352_ & new_n1346_;
  assign new_n1719_ = new_n1351_ | new_n1345_;
  assign new_n1720_ = new_n6406_ & new_n875_;
  assign new_n1721_ = new_n6414_ | new_n876_;
  assign new_n1722_ = new_n6419_ & new_n6420_;
  assign new_n1723_ = new_n6421_ | new_n6422_;
  assign new_n1724_ = new_n6424_ & new_n6420_;
  assign new_n1725_ = new_n6426_ | new_n6422_;
  assign new_n1726_ = new_n6424_ & new_n6419_;
  assign new_n1727_ = new_n6426_ | new_n6421_;
  assign new_n1728_ = new_n1727_ & new_n1725_;
  assign new_n1729_ = new_n1726_ | new_n1724_;
  assign new_n1730_ = new_n6387_ & new_n1217_;
  assign new_n1731_ = new_n6389_ | new_n1218_;
  assign new_n1732_ = new_n6427_ & new_n6428_;
  assign new_n1733_ = new_n6429_ | new_n6430_;
  assign new_n1734_ = new_n6432_ & new_n6428_;
  assign new_n1735_ = new_n6434_ | new_n6430_;
  assign new_n1736_ = new_n6432_ & new_n6427_;
  assign new_n1737_ = new_n6434_ | new_n6429_;
  assign new_n1738_ = new_n1737_ & new_n1735_;
  assign new_n1739_ = new_n1736_ | new_n1734_;
  assign new_n1740_ = new_n1714_ & new_n6395_;
  assign new_n1741_ = new_n6401_ | new_n6397_;
  assign new_n1742_ = new_n1741_ & new_n1739_;
  assign new_n1743_ = new_n6435_ | new_n6436_;
  assign new_n1744_ = new_n6438_ | new_n6436_;
  assign new_n1745_ = new_n6438_ | new_n6435_;
  assign new_n1746_ = new_n1745_ & new_n1744_;
  assign new_n1747_ = new_n6439_ & new_n6440_;
  assign new_n1748_ = new_n6441_ | new_n6442_;
  assign new_n1749_ = new_n6444_ & new_n6439_;
  assign new_n1750_ = new_n6446_ | new_n6441_;
  assign new_n1751_ = new_n6444_ & new_n6440_;
  assign new_n1752_ = new_n6446_ | new_n6442_;
  assign new_n1753_ = new_n1752_ & new_n1750_;
  assign new_n1754_ = new_n1751_ | new_n1749_;
  assign new_n1755_ = new_n6406_ & new_n877_;
  assign new_n1756_ = new_n6414_ | new_n878_;
  assign new_n1757_ = new_n6447_ & new_n6448_;
  assign new_n1758_ = new_n6449_ | new_n6450_;
  assign new_n1759_ = new_n6452_ & new_n6448_;
  assign new_n1760_ = new_n6454_ | new_n6450_;
  assign new_n1761_ = new_n6452_ & new_n6447_;
  assign new_n1762_ = new_n6454_ | new_n6449_;
  assign new_n1763_ = new_n1762_ & new_n1760_;
  assign new_n1764_ = new_n1761_ | new_n1759_;
  assign new_n1765_ = new_n6423_ & new_n1279_;
  assign new_n1766_ = new_n6425_ | new_n1280_;
  assign new_n1767_ = new_n6455_ & new_n6456_;
  assign new_n1768_ = new_n6457_ | new_n6458_;
  assign new_n1769_ = new_n6460_ & new_n6456_;
  assign new_n1770_ = new_n6462_ | new_n6458_;
  assign new_n1771_ = new_n6460_ & new_n6455_;
  assign new_n1772_ = new_n6462_ | new_n6457_;
  assign new_n1773_ = new_n1772_ & new_n1770_;
  assign new_n1774_ = new_n1771_ | new_n1769_;
  assign new_n1775_ = new_n1743_ & new_n6431_;
  assign new_n1776_ = new_n6437_ | new_n6433_;
  assign new_n1777_ = new_n1776_ & new_n1774_;
  assign new_n1778_ = new_n6463_ | new_n6464_;
  assign new_n1779_ = new_n6466_ | new_n6464_;
  assign new_n1780_ = new_n6466_ | new_n6463_;
  assign new_n1781_ = new_n1780_ & new_n1779_;
  assign new_n1782_ = new_n6468_ & new_n1285_;
  assign new_n1783_ = new_n6470_ | new_n1286_;
  assign new_n1784_ = new_n6468_ & new_n1272_;
  assign new_n1785_ = new_n6470_ | new_n1271_;
  assign new_n1786_ = new_n1785_ & new_n1783_;
  assign new_n1787_ = new_n1784_ | new_n1782_;
  assign new_n1788_ = new_n1238_ & new_n1175_;
  assign new_n1789_ = new_n1237_ | new_n1176_;
  assign new_n1790_ = new_n6471_ & new_n6472_;
  assign new_n1791_ = new_n6473_ | new_n6474_;
  assign new_n1792_ = new_n6476_ & new_n6472_;
  assign new_n1793_ = new_n6478_ | new_n6474_;
  assign new_n1794_ = new_n6476_ & new_n6471_;
  assign new_n1795_ = new_n6478_ | new_n6473_;
  assign new_n1796_ = new_n1795_ & new_n1793_;
  assign new_n1797_ = new_n1794_ | new_n1792_;
  assign new_n1798_ = new_n6405_ & new_n879_;
  assign new_n1799_ = new_n6413_ | new_n880_;
  assign new_n1800_ = new_n6479_ & new_n6480_;
  assign new_n1801_ = new_n6481_ | new_n6482_;
  assign new_n1802_ = new_n6484_ & new_n6480_;
  assign new_n1803_ = new_n6486_ | new_n6482_;
  assign new_n1804_ = new_n6484_ & new_n6479_;
  assign new_n1805_ = new_n6486_ | new_n6481_;
  assign new_n1806_ = new_n1805_ & new_n1803_;
  assign new_n1807_ = new_n1804_ | new_n1802_;
  assign new_n1808_ = new_n6451_ & new_n6443_;
  assign new_n1809_ = new_n6453_ | new_n6445_;
  assign new_n1810_ = new_n6487_ & new_n6488_;
  assign new_n1811_ = new_n6489_ | new_n6490_;
  assign new_n1812_ = new_n6492_ & new_n6488_;
  assign new_n1813_ = new_n6494_ | new_n6490_;
  assign new_n1814_ = new_n6492_ & new_n6487_;
  assign new_n1815_ = new_n6494_ | new_n6489_;
  assign new_n1816_ = new_n1815_ & new_n1813_;
  assign new_n1817_ = new_n1814_ | new_n1812_;
  assign new_n1818_ = new_n1778_ & new_n6459_;
  assign new_n1819_ = new_n6465_ | new_n6461_;
  assign new_n1820_ = new_n1819_ & new_n1817_;
  assign new_n1821_ = new_n6495_ | new_n6496_;
  assign new_n1822_ = new_n6498_ | new_n6496_;
  assign new_n1823_ = new_n6498_ | new_n6495_;
  assign new_n1824_ = new_n1823_ & new_n1822_;
  assign new_n1825_ = new_n1354_ & new_n1344_;
  assign new_n1826_ = new_n1353_ | new_n1343_;
  assign new_n1827_ = new_n6501_ & new_n6503_;
  assign new_n1828_ = new_n6506_ | new_n6508_;
  assign new_n1829_ = new_n6509_ & new_n6510_;
  assign new_n1830_ = new_n6511_ | new_n6512_;
  assign new_n1831_ = new_n6514_ & new_n6510_;
  assign new_n1832_ = new_n6516_ | new_n6512_;
  assign new_n1833_ = new_n6514_ & new_n6509_;
  assign new_n1834_ = new_n6516_ | new_n6511_;
  assign new_n1835_ = new_n1834_ & new_n1832_;
  assign new_n1836_ = new_n1833_ | new_n1831_;
  assign new_n1837_ = new_n6467_ & new_n1215_;
  assign new_n1838_ = new_n6469_ | new_n1216_;
  assign new_n1839_ = new_n6517_ & new_n6518_;
  assign new_n1840_ = new_n6519_ | new_n6520_;
  assign new_n1841_ = new_n6522_ & new_n6518_;
  assign new_n1842_ = new_n6524_ | new_n6520_;
  assign new_n1843_ = new_n6522_ & new_n6517_;
  assign new_n1844_ = new_n6524_ | new_n6519_;
  assign new_n1845_ = new_n1844_ & new_n1842_;
  assign new_n1846_ = new_n1843_ | new_n1841_;
  assign new_n1847_ = new_n6407_ & new_n881_;
  assign new_n1848_ = new_n6415_ | new_n882_;
  assign new_n1849_ = new_n6525_ & new_n6526_;
  assign new_n1850_ = new_n6527_ | new_n6528_;
  assign new_n1851_ = new_n6530_ & new_n6526_;
  assign new_n1852_ = new_n6532_ | new_n6528_;
  assign new_n1853_ = new_n6530_ & new_n6525_;
  assign new_n1854_ = new_n6532_ | new_n6527_;
  assign new_n1855_ = new_n1854_ & new_n1852_;
  assign new_n1856_ = new_n1853_ | new_n1851_;
  assign new_n1857_ = new_n6483_ & new_n6475_;
  assign new_n1858_ = new_n6485_ | new_n6477_;
  assign new_n1859_ = new_n6533_ & new_n6534_;
  assign new_n1860_ = new_n6535_ | new_n6536_;
  assign new_n1861_ = new_n6538_ & new_n6534_;
  assign new_n1862_ = new_n6540_ | new_n6536_;
  assign new_n1863_ = new_n6538_ & new_n6533_;
  assign new_n1864_ = new_n6540_ | new_n6535_;
  assign new_n1865_ = new_n1864_ & new_n1862_;
  assign new_n1866_ = new_n1863_ | new_n1861_;
  assign new_n1867_ = new_n1821_ & new_n6491_;
  assign new_n1868_ = new_n6497_ | new_n6493_;
  assign new_n1869_ = new_n1868_ & new_n1866_;
  assign new_n1870_ = new_n6541_ | new_n6542_;
  assign new_n1871_ = new_n6544_ | new_n6542_;
  assign new_n1872_ = new_n6544_ | new_n6541_;
  assign new_n1873_ = new_n1872_ & new_n1871_;
  assign new_n1874_ = new_n6545_ & new_n6546_;
  assign new_n1875_ = new_n6547_ | new_n6548_;
  assign new_n1876_ = new_n6550_ & new_n6545_;
  assign new_n1877_ = new_n6552_ | new_n6547_;
  assign new_n1878_ = new_n6550_ & new_n6546_;
  assign new_n1879_ = new_n6552_ | new_n6548_;
  assign new_n1880_ = new_n1879_ & new_n1877_;
  assign new_n1881_ = new_n1878_ | new_n1876_;
  assign new_n1882_ = new_n6501_ & new_n6553_;
  assign new_n1883_ = new_n6506_ | new_n6554_;
  assign new_n1884_ = new_n6555_ & new_n6556_;
  assign new_n1885_ = new_n6557_ | new_n6558_;
  assign new_n1886_ = new_n6560_ & new_n6556_;
  assign new_n1887_ = new_n6562_ | new_n6558_;
  assign new_n1888_ = new_n6560_ & new_n6555_;
  assign new_n1889_ = new_n6562_ | new_n6557_;
  assign new_n1890_ = new_n1889_ & new_n1887_;
  assign new_n1891_ = new_n1888_ | new_n1886_;
  assign new_n1892_ = new_n6513_ & new_n1277_;
  assign new_n1893_ = new_n6515_ | new_n1278_;
  assign new_n1894_ = new_n6563_ & new_n6564_;
  assign new_n1895_ = new_n6565_ | new_n6566_;
  assign new_n1896_ = new_n6568_ & new_n6564_;
  assign new_n1897_ = new_n6570_ | new_n6566_;
  assign new_n1898_ = new_n6568_ & new_n6563_;
  assign new_n1899_ = new_n6570_ | new_n6565_;
  assign new_n1900_ = new_n1899_ & new_n1897_;
  assign new_n1901_ = new_n1898_ | new_n1896_;
  assign new_n1902_ = new_n6407_ & new_n6503_;
  assign new_n1903_ = new_n6415_ | new_n6508_;
  assign new_n1904_ = new_n6571_ & new_n6572_;
  assign new_n1905_ = new_n6573_ | new_n6574_;
  assign new_n1906_ = new_n6576_ & new_n6572_;
  assign new_n1907_ = new_n6578_ | new_n6574_;
  assign new_n1908_ = new_n6576_ & new_n6571_;
  assign new_n1909_ = new_n6578_ | new_n6573_;
  assign new_n1910_ = new_n1909_ & new_n1907_;
  assign new_n1911_ = new_n1908_ | new_n1906_;
  assign new_n1912_ = new_n6529_ & new_n6521_;
  assign new_n1913_ = new_n6531_ | new_n6523_;
  assign new_n1914_ = new_n6579_ & new_n6580_;
  assign new_n1915_ = new_n6581_ | new_n6582_;
  assign new_n1916_ = new_n6584_ & new_n6580_;
  assign new_n1917_ = new_n6586_ | new_n6582_;
  assign new_n1918_ = new_n6584_ & new_n6579_;
  assign new_n1919_ = new_n6586_ | new_n6581_;
  assign new_n1920_ = new_n1919_ & new_n1917_;
  assign new_n1921_ = new_n1918_ | new_n1916_;
  assign new_n1922_ = new_n1870_ & new_n6537_;
  assign new_n1923_ = new_n6543_ | new_n6539_;
  assign new_n1924_ = new_n1923_ & new_n1921_;
  assign new_n1925_ = new_n6587_ | new_n6588_;
  assign new_n1926_ = new_n6590_ | new_n6588_;
  assign new_n1927_ = new_n6590_ | new_n6587_;
  assign new_n1928_ = new_n1927_ & new_n1926_;
  assign new_n1929_ = new_n6592_ & new_n1283_;
  assign new_n1930_ = new_n6594_ | new_n1284_;
  assign new_n1931_ = new_n6592_ & new_n1274_;
  assign new_n1932_ = new_n6594_ | new_n1273_;
  assign new_n1933_ = new_n1932_ & new_n1930_;
  assign new_n1934_ = new_n1931_ | new_n1929_;
  assign new_n1935_ = new_n1240_ & new_n1173_;
  assign new_n1936_ = new_n1239_ | new_n1174_;
  assign new_n1937_ = new_n6595_ & new_n6596_;
  assign new_n1938_ = new_n6597_ | new_n6598_;
  assign new_n1939_ = new_n6600_ & new_n6596_;
  assign new_n1940_ = new_n6602_ | new_n6598_;
  assign new_n1941_ = new_n6600_ & new_n6595_;
  assign new_n1942_ = new_n6602_ | new_n6597_;
  assign new_n1943_ = new_n1942_ & new_n1940_;
  assign new_n1944_ = new_n1941_ | new_n1939_;
  assign new_n1945_ = new_n6500_ & new_n6603_;
  assign new_n1946_ = new_n6505_ | new_n6604_;
  assign new_n1947_ = new_n6605_ & new_n6606_;
  assign new_n1948_ = new_n6607_ | new_n6608_;
  assign new_n1949_ = new_n6610_ & new_n6606_;
  assign new_n1950_ = new_n6612_ | new_n6608_;
  assign new_n1951_ = new_n6610_ & new_n6605_;
  assign new_n1952_ = new_n6612_ | new_n6607_;
  assign new_n1953_ = new_n1952_ & new_n1950_;
  assign new_n1954_ = new_n1951_ | new_n1949_;
  assign new_n1955_ = new_n6559_ & new_n6549_;
  assign new_n1956_ = new_n6561_ | new_n6551_;
  assign new_n1957_ = new_n6613_ & new_n6614_;
  assign new_n1958_ = new_n6615_ | new_n6616_;
  assign new_n1959_ = new_n6618_ & new_n6614_;
  assign new_n1960_ = new_n6620_ | new_n6616_;
  assign new_n1961_ = new_n6618_ & new_n6613_;
  assign new_n1962_ = new_n6620_ | new_n6615_;
  assign new_n1963_ = new_n1962_ & new_n1960_;
  assign new_n1964_ = new_n1961_ | new_n1959_;
  assign new_n1965_ = new_n6409_ & new_n6553_;
  assign new_n1966_ = new_n6417_ | new_n6554_;
  assign new_n1967_ = new_n6621_ & new_n6622_;
  assign new_n1968_ = new_n6623_ | new_n6624_;
  assign new_n1969_ = new_n6626_ & new_n6622_;
  assign new_n1970_ = new_n6628_ | new_n6624_;
  assign new_n1971_ = new_n6626_ & new_n6621_;
  assign new_n1972_ = new_n6628_ | new_n6623_;
  assign new_n1973_ = new_n1972_ & new_n1970_;
  assign new_n1974_ = new_n1971_ | new_n1969_;
  assign new_n1975_ = new_n6575_ & new_n6567_;
  assign new_n1976_ = new_n6577_ | new_n6569_;
  assign new_n1977_ = new_n6629_ & new_n6630_;
  assign new_n1978_ = new_n6631_ | new_n6632_;
  assign new_n1979_ = new_n6634_ & new_n6630_;
  assign new_n1980_ = new_n6636_ | new_n6632_;
  assign new_n1981_ = new_n6634_ & new_n6629_;
  assign new_n1982_ = new_n6636_ | new_n6631_;
  assign new_n1983_ = new_n1982_ & new_n1980_;
  assign new_n1984_ = new_n1981_ | new_n1979_;
  assign new_n1985_ = new_n1925_ & new_n6583_;
  assign new_n1986_ = new_n6589_ | new_n6585_;
  assign new_n1987_ = new_n1986_ & new_n1984_;
  assign new_n1988_ = new_n6637_ | new_n6638_;
  assign new_n1989_ = new_n6640_ | new_n6638_;
  assign new_n1990_ = new_n6640_ | new_n6637_;
  assign new_n1991_ = new_n1990_ & new_n1989_;
  assign new_n1992_ = new_n925_ & new_n6642_;
  assign new_n1993_ = new_n926_ | new_n6644_;
  assign new_n1994_ = new_n6591_ & new_n1213_;
  assign new_n1995_ = new_n6593_ | new_n1214_;
  assign new_n1996_ = new_n6645_ & new_n6646_;
  assign new_n1997_ = new_n6647_ | new_n6648_;
  assign new_n1998_ = new_n6650_ & new_n6646_;
  assign new_n1999_ = new_n6652_ | new_n6648_;
  assign new_n2000_ = new_n6650_ & new_n6645_;
  assign new_n2001_ = new_n6652_ | new_n6647_;
  assign new_n2002_ = new_n2001_ & new_n1999_;
  assign new_n2003_ = new_n2000_ | new_n1998_;
  assign new_n2004_ = new_n6502_ & new_n6653_;
  assign new_n2005_ = new_n6507_ | new_n6654_;
  assign new_n2006_ = new_n6655_ & new_n6656_;
  assign new_n2007_ = new_n6657_ | new_n6658_;
  assign new_n2008_ = new_n6660_ & new_n6656_;
  assign new_n2009_ = new_n6662_ | new_n6658_;
  assign new_n2010_ = new_n6660_ & new_n6655_;
  assign new_n2011_ = new_n6662_ | new_n6657_;
  assign new_n2012_ = new_n2011_ & new_n2009_;
  assign new_n2013_ = new_n2010_ | new_n2008_;
  assign new_n2014_ = new_n6609_ & new_n6599_;
  assign new_n2015_ = new_n6611_ | new_n6601_;
  assign new_n2016_ = new_n6663_ & new_n6664_;
  assign new_n2017_ = new_n6665_ | new_n6666_;
  assign new_n2018_ = new_n6668_ & new_n6664_;
  assign new_n2019_ = new_n6670_ | new_n6666_;
  assign new_n2020_ = new_n6668_ & new_n6663_;
  assign new_n2021_ = new_n6670_ | new_n6665_;
  assign new_n2022_ = new_n2021_ & new_n2019_;
  assign new_n2023_ = new_n2020_ | new_n2018_;
  assign new_n2024_ = new_n6409_ & new_n6603_;
  assign new_n2025_ = new_n6417_ | new_n6604_;
  assign new_n2026_ = new_n6671_ & new_n6672_;
  assign new_n2027_ = new_n6673_ | new_n6674_;
  assign new_n2028_ = new_n6676_ & new_n6672_;
  assign new_n2029_ = new_n6678_ | new_n6674_;
  assign new_n2030_ = new_n6676_ & new_n6671_;
  assign new_n2031_ = new_n6678_ | new_n6673_;
  assign new_n2032_ = new_n2031_ & new_n2029_;
  assign new_n2033_ = new_n2030_ | new_n2028_;
  assign new_n2034_ = new_n6625_ & new_n6617_;
  assign new_n2035_ = new_n6627_ | new_n6619_;
  assign new_n2036_ = new_n6679_ & new_n6680_;
  assign new_n2037_ = new_n6681_ | new_n6682_;
  assign new_n2038_ = new_n6684_ & new_n6680_;
  assign new_n2039_ = new_n6686_ | new_n6682_;
  assign new_n2040_ = new_n6684_ & new_n6679_;
  assign new_n2041_ = new_n6686_ | new_n6681_;
  assign new_n2042_ = new_n2041_ & new_n2039_;
  assign new_n2043_ = new_n2040_ | new_n2038_;
  assign new_n2044_ = new_n1988_ & new_n6633_;
  assign new_n2045_ = new_n6639_ | new_n6635_;
  assign new_n2046_ = new_n2045_ & new_n2043_;
  assign new_n2047_ = new_n6687_ | new_n6688_;
  assign new_n2048_ = new_n6690_ | new_n6688_;
  assign new_n2049_ = new_n6690_ | new_n6687_;
  assign new_n2050_ = new_n2049_ & new_n2048_;
  assign new_n2051_ = new_n6502_ & new_n6642_;
  assign new_n2052_ = new_n6507_ | new_n6644_;
  assign new_n2053_ = new_n6659_ & new_n6649_;
  assign new_n2054_ = new_n6661_ | new_n6651_;
  assign new_n2055_ = new_n6691_ & new_n6692_;
  assign new_n2056_ = new_n6693_ | new_n6694_;
  assign new_n2057_ = new_n6696_ & new_n6692_;
  assign new_n2058_ = new_n6698_ | new_n6694_;
  assign new_n2059_ = new_n6696_ & new_n6691_;
  assign new_n2060_ = new_n6698_ | new_n6693_;
  assign new_n2061_ = new_n2060_ & new_n2058_;
  assign new_n2062_ = new_n2059_ | new_n2057_;
  assign new_n2063_ = new_n6410_ & new_n6653_;
  assign new_n2064_ = new_n6418_ | new_n6654_;
  assign new_n2065_ = new_n6699_ & new_n6700_;
  assign new_n2066_ = new_n6701_ | new_n6702_;
  assign new_n2067_ = new_n6704_ & new_n6700_;
  assign new_n2068_ = new_n6706_ | new_n6702_;
  assign new_n2069_ = new_n6704_ & new_n6699_;
  assign new_n2070_ = new_n6706_ | new_n6701_;
  assign new_n2071_ = new_n2070_ & new_n2068_;
  assign new_n2072_ = new_n2069_ | new_n2067_;
  assign new_n2073_ = new_n6675_ & new_n6667_;
  assign new_n2074_ = new_n6677_ | new_n6669_;
  assign new_n2075_ = new_n6707_ & new_n6708_;
  assign new_n2076_ = new_n6709_ | new_n6710_;
  assign new_n2077_ = new_n6712_ & new_n6708_;
  assign new_n2078_ = new_n6714_ | new_n6710_;
  assign new_n2079_ = new_n6712_ & new_n6707_;
  assign new_n2080_ = new_n6714_ | new_n6709_;
  assign new_n2081_ = new_n2080_ & new_n2078_;
  assign new_n2082_ = new_n2079_ | new_n2077_;
  assign new_n2083_ = new_n2047_ & new_n6683_;
  assign new_n2084_ = new_n6689_ | new_n6685_;
  assign new_n2085_ = new_n2084_ & new_n2082_;
  assign new_n2086_ = new_n6715_ | new_n6716_;
  assign new_n2087_ = new_n6718_ | new_n6716_;
  assign new_n2088_ = new_n6718_ | new_n6715_;
  assign new_n2089_ = new_n2088_ & new_n2087_;
  assign new_n2090_ = new_n6410_ & new_n6641_;
  assign new_n2091_ = new_n6418_ | new_n6643_;
  assign new_n2092_ = new_n6703_ & new_n6695_;
  assign new_n2093_ = new_n6705_ | new_n6697_;
  assign new_n2094_ = new_n6719_ & new_n6720_;
  assign new_n2095_ = new_n6721_ | new_n6722_;
  assign new_n2096_ = new_n6724_ & new_n6720_;
  assign new_n2097_ = new_n6725_ | new_n6722_;
  assign new_n2098_ = new_n6724_ & new_n6719_;
  assign new_n2099_ = new_n6725_ | new_n6721_;
  assign new_n2100_ = new_n2099_ & new_n2097_;
  assign new_n2101_ = new_n2098_ | new_n2096_;
  assign new_n2102_ = new_n2086_ & new_n6711_;
  assign new_n2103_ = new_n6717_ | new_n6713_;
  assign new_n2104_ = new_n2102_ | new_n2100_;
  assign new_n2105_ = new_n6727_ & new_n6723_;
  assign new_n2106_ = new_n6727_ & new_n2101_;
  assign new_n2107_ = new_n6726_ & new_n2103_;
  assign new_n2108_ = new_n2107_ | new_n2106_;
  assign new_n2109_ = new_n6731_ & new_n6740_;
  assign new_n2110_ = new_n6745_ | new_n6753_;
  assign new_n2111_ = new_n1438_ & new_n1432_;
  assign new_n2112_ = new_n1437_ | new_n1431_;
  assign new_n2113_ = new_n6755_ & new_n2110_;
  assign new_n2114_ = new_n2111_ | new_n6756_;
  assign new_n2115_ = new_n6740_ & new_n6760_;
  assign new_n2116_ = new_n6753_ | new_n6774_;
  assign new_n2117_ = new_n6785_ & new_n6786_;
  assign new_n2118_ = new_n6787_ | new_n6788_;
  assign new_n2119_ = new_n6790_ & new_n6785_;
  assign new_n2120_ = new_n6792_ | new_n6787_;
  assign new_n2121_ = new_n6790_ & new_n6786_;
  assign new_n2122_ = new_n6792_ | new_n6788_;
  assign new_n2123_ = new_n2122_ & new_n2120_;
  assign new_n2124_ = new_n2121_ | new_n2119_;
  assign new_n2125_ = new_n2114_ & new_n1375_;
  assign new_n2126_ = new_n6793_ | new_n1376_;
  assign new_n2127_ = new_n6794_ & new_n6795_;
  assign new_n2128_ = new_n6796_ | new_n6797_;
  assign new_n2129_ = new_n6799_ & new_n6795_;
  assign new_n2130_ = new_n6801_ | new_n6797_;
  assign new_n2131_ = new_n6799_ & new_n6794_;
  assign new_n2132_ = new_n6801_ | new_n6796_;
  assign new_n2133_ = new_n2132_ & new_n2130_;
  assign new_n2134_ = new_n2131_ | new_n2129_;
  assign new_n2135_ = new_n6802_ & new_n2116_;
  assign new_n2136_ = new_n2133_ | new_n6803_;
  assign new_n2137_ = new_n6739_ & new_n6807_;
  assign new_n2138_ = new_n6754_ | new_n6817_;
  assign new_n2139_ = new_n6825_ & new_n1383_;
  assign new_n2140_ = new_n6827_ | new_n1384_;
  assign new_n2141_ = new_n6825_ & new_n1336_;
  assign new_n2142_ = new_n6827_ | new_n1335_;
  assign new_n2143_ = new_n2142_ & new_n2140_;
  assign new_n2144_ = new_n2141_ | new_n2139_;
  assign new_n2145_ = new_n6789_ & new_n1311_;
  assign new_n2146_ = new_n6791_ | new_n1312_;
  assign new_n2147_ = new_n6828_ & new_n6829_;
  assign new_n2148_ = new_n6830_ | new_n6831_;
  assign new_n2149_ = new_n6833_ & new_n6829_;
  assign new_n2150_ = new_n6835_ | new_n6831_;
  assign new_n2151_ = new_n6833_ & new_n6828_;
  assign new_n2152_ = new_n6835_ | new_n6830_;
  assign new_n2153_ = new_n2152_ & new_n2150_;
  assign new_n2154_ = new_n2151_ | new_n2149_;
  assign new_n2155_ = new_n6837_ & new_n6760_;
  assign new_n2156_ = new_n6839_ | new_n6774_;
  assign new_n2157_ = new_n6840_ & new_n6841_;
  assign new_n2158_ = new_n6842_ | new_n6843_;
  assign new_n2159_ = new_n6845_ & new_n6841_;
  assign new_n2160_ = new_n6847_ | new_n6843_;
  assign new_n2161_ = new_n6845_ & new_n6840_;
  assign new_n2162_ = new_n6847_ | new_n6842_;
  assign new_n2163_ = new_n2162_ & new_n2160_;
  assign new_n2164_ = new_n2161_ | new_n2159_;
  assign new_n2165_ = new_n2136_ & new_n6798_;
  assign new_n2166_ = new_n6848_ | new_n6800_;
  assign new_n2167_ = new_n6849_ & new_n6850_;
  assign new_n2168_ = new_n6851_ | new_n6852_;
  assign new_n2169_ = new_n6854_ & new_n6850_;
  assign new_n2170_ = new_n6856_ | new_n6852_;
  assign new_n2171_ = new_n6854_ & new_n6849_;
  assign new_n2172_ = new_n6856_ | new_n6851_;
  assign new_n2173_ = new_n2172_ & new_n2170_;
  assign new_n2174_ = new_n2171_ | new_n2169_;
  assign new_n2175_ = new_n6857_ & new_n2138_;
  assign new_n2176_ = new_n2173_ | new_n6858_;
  assign new_n2177_ = new_n6861_ & new_n6865_;
  assign new_n2178_ = new_n6870_ | new_n6874_;
  assign new_n2179_ = new_n6877_ & new_n1474_;
  assign new_n2180_ = new_n6879_ | new_n1473_;
  assign new_n2181_ = new_n6877_ & new_n1418_;
  assign new_n2182_ = new_n6879_ | new_n1417_;
  assign new_n2183_ = new_n2182_ & new_n2180_;
  assign new_n2184_ = new_n2181_ | new_n2179_;
  assign new_n2185_ = new_n6880_ & new_n2178_;
  assign new_n2186_ = new_n2183_ | new_n6881_;
  assign new_n2187_ = new_n6741_ & new_n6884_;
  assign new_n2188_ = new_n6754_ | new_n6890_;
  assign new_n2189_ = new_n1440_ & new_n1423_;
  assign new_n2190_ = new_n1439_ | new_n1424_;
  assign new_n2191_ = new_n6824_ & new_n1299_;
  assign new_n2192_ = new_n6826_ | new_n1300_;
  assign new_n2193_ = new_n6894_ & new_n6895_;
  assign new_n2194_ = new_n6896_ | new_n6897_;
  assign new_n2195_ = new_n6899_ & new_n6895_;
  assign new_n2196_ = new_n6901_ | new_n6897_;
  assign new_n2197_ = new_n6899_ & new_n6894_;
  assign new_n2198_ = new_n6901_ | new_n6896_;
  assign new_n2199_ = new_n2198_ & new_n2196_;
  assign new_n2200_ = new_n2197_ | new_n2195_;
  assign new_n2201_ = new_n6903_ & new_n6761_;
  assign new_n2202_ = new_n6905_ | new_n6775_;
  assign new_n2203_ = new_n6906_ & new_n6907_;
  assign new_n2204_ = new_n6908_ | new_n6909_;
  assign new_n2205_ = new_n6911_ & new_n6907_;
  assign new_n2206_ = new_n6913_ | new_n6909_;
  assign new_n2207_ = new_n6911_ & new_n6906_;
  assign new_n2208_ = new_n6913_ | new_n6908_;
  assign new_n2209_ = new_n2208_ & new_n2206_;
  assign new_n2210_ = new_n2207_ | new_n2205_;
  assign new_n2211_ = new_n6844_ & new_n6832_;
  assign new_n2212_ = new_n6846_ | new_n6834_;
  assign new_n2213_ = new_n6914_ & new_n6915_;
  assign new_n2214_ = new_n6916_ | new_n6917_;
  assign new_n2215_ = new_n6919_ & new_n6915_;
  assign new_n2216_ = new_n6921_ | new_n6917_;
  assign new_n2217_ = new_n6919_ & new_n6914_;
  assign new_n2218_ = new_n6921_ | new_n6916_;
  assign new_n2219_ = new_n2218_ & new_n2216_;
  assign new_n2220_ = new_n2217_ | new_n2215_;
  assign new_n2221_ = new_n6837_ & new_n6807_;
  assign new_n2222_ = new_n6839_ | new_n6817_;
  assign new_n2223_ = new_n6922_ & new_n6923_;
  assign new_n2224_ = new_n6924_ | new_n6925_;
  assign new_n2225_ = new_n6927_ & new_n6923_;
  assign new_n2226_ = new_n6929_ | new_n6925_;
  assign new_n2227_ = new_n6927_ & new_n6922_;
  assign new_n2228_ = new_n6929_ | new_n6924_;
  assign new_n2229_ = new_n2228_ & new_n2226_;
  assign new_n2230_ = new_n2227_ | new_n2225_;
  assign new_n2231_ = new_n2176_ & new_n6853_;
  assign new_n2232_ = new_n6930_ | new_n6855_;
  assign new_n2233_ = new_n6931_ & new_n6932_;
  assign new_n2234_ = new_n6933_ | new_n6934_;
  assign new_n2235_ = new_n6936_ & new_n6932_;
  assign new_n2236_ = new_n6938_ | new_n6934_;
  assign new_n2237_ = new_n6936_ & new_n6931_;
  assign new_n2238_ = new_n6938_ | new_n6933_;
  assign new_n2239_ = new_n2238_ & new_n2236_;
  assign new_n2240_ = new_n2237_ | new_n2235_;
  assign new_n2241_ = new_n6942_ & new_n6865_;
  assign new_n2242_ = new_n6955_ | new_n6874_;
  assign new_n2243_ = new_n6965_ & new_n2188_;
  assign new_n2244_ = new_n2239_ | new_n6966_;
  assign new_n2245_ = new_n1522_ & new_n1512_;
  assign new_n2246_ = new_n1521_ | new_n1511_;
  assign new_n2247_ = new_n6861_ & new_n6969_;
  assign new_n2248_ = new_n6870_ | new_n6975_;
  assign new_n2249_ = new_n6977_ & new_n6978_;
  assign new_n2250_ = new_n6979_ | new_n6980_;
  assign new_n2251_ = new_n6982_ & new_n6978_;
  assign new_n2252_ = new_n6984_ | new_n6980_;
  assign new_n2253_ = new_n6982_ & new_n6977_;
  assign new_n2254_ = new_n6984_ | new_n6979_;
  assign new_n2255_ = new_n2254_ & new_n2252_;
  assign new_n2256_ = new_n2253_ | new_n2251_;
  assign new_n2257_ = new_n2186_ & new_n6876_;
  assign new_n2258_ = new_n6985_ | new_n6878_;
  assign new_n2259_ = new_n6986_ & new_n6987_;
  assign new_n2260_ = new_n6988_ | new_n6989_;
  assign new_n2261_ = new_n6991_ & new_n6987_;
  assign new_n2262_ = new_n6993_ | new_n6989_;
  assign new_n2263_ = new_n6991_ & new_n6986_;
  assign new_n2264_ = new_n6993_ | new_n6988_;
  assign new_n2265_ = new_n2264_ & new_n2262_;
  assign new_n2266_ = new_n2263_ | new_n2261_;
  assign new_n2267_ = new_n6994_ & new_n2242_;
  assign new_n2268_ = new_n2265_ | new_n6995_;
  assign new_n2269_ = new_n6998_ & new_n7001_;
  assign new_n2270_ = new_n7004_ | new_n7007_;
  assign new_n2271_ = new_n7008_ & new_n7009_;
  assign new_n2272_ = new_n7010_ | new_n7011_;
  assign new_n2273_ = new_n7013_ & new_n7008_;
  assign new_n2274_ = new_n7015_ | new_n7010_;
  assign new_n2275_ = new_n7013_ & new_n7009_;
  assign new_n2276_ = new_n7015_ | new_n7011_;
  assign new_n2277_ = new_n2276_ & new_n2274_;
  assign new_n2278_ = new_n2275_ | new_n2273_;
  assign new_n2279_ = new_n6866_ & new_n7019_;
  assign new_n2280_ = new_n6873_ | new_n7034_;
  assign new_n2281_ = new_n7046_ & new_n2270_;
  assign new_n2282_ = new_n2277_ | new_n7047_;
  assign new_n2283_ = new_n7048_ & new_n7049_;
  assign new_n2284_ = new_n7050_ | new_n7051_;
  assign new_n2285_ = new_n7053_ & new_n7048_;
  assign new_n2286_ = new_n7055_ | new_n7050_;
  assign new_n2287_ = new_n7053_ & new_n7049_;
  assign new_n2288_ = new_n7055_ | new_n7051_;
  assign new_n2289_ = new_n2288_ & new_n2286_;
  assign new_n2290_ = new_n2287_ | new_n2285_;
  assign new_n2291_ = new_n6981_ & new_n1455_;
  assign new_n2292_ = new_n6983_ | new_n1456_;
  assign new_n2293_ = new_n7056_ & new_n7057_;
  assign new_n2294_ = new_n7058_ | new_n7059_;
  assign new_n2295_ = new_n7061_ & new_n7057_;
  assign new_n2296_ = new_n7063_ | new_n7059_;
  assign new_n2297_ = new_n7061_ & new_n7056_;
  assign new_n2298_ = new_n7063_ | new_n7058_;
  assign new_n2299_ = new_n2298_ & new_n2296_;
  assign new_n2300_ = new_n2297_ | new_n2295_;
  assign new_n2301_ = new_n6942_ & new_n6969_;
  assign new_n2302_ = new_n6955_ | new_n6975_;
  assign new_n2303_ = new_n7064_ & new_n7065_;
  assign new_n2304_ = new_n7066_ | new_n7067_;
  assign new_n2305_ = new_n7069_ & new_n7065_;
  assign new_n2306_ = new_n7071_ | new_n7067_;
  assign new_n2307_ = new_n7069_ & new_n7064_;
  assign new_n2308_ = new_n7071_ | new_n7066_;
  assign new_n2309_ = new_n2308_ & new_n2306_;
  assign new_n2310_ = new_n2307_ | new_n2305_;
  assign new_n2311_ = new_n2268_ & new_n6990_;
  assign new_n2312_ = new_n7072_ | new_n6992_;
  assign new_n2313_ = new_n7073_ & new_n7074_;
  assign new_n2314_ = new_n7075_ | new_n7076_;
  assign new_n2315_ = new_n7078_ & new_n7074_;
  assign new_n2316_ = new_n7080_ | new_n7076_;
  assign new_n2317_ = new_n7078_ & new_n7073_;
  assign new_n2318_ = new_n7080_ | new_n7075_;
  assign new_n2319_ = new_n2318_ & new_n2316_;
  assign new_n2320_ = new_n2317_ | new_n2315_;
  assign new_n2321_ = new_n7081_ & new_n2280_;
  assign new_n2322_ = new_n2319_ | new_n7082_;
  assign new_n2323_ = new_n6998_ & new_n7086_;
  assign new_n2324_ = new_n7004_ | new_n7094_;
  assign new_n2325_ = new_n7100_ & new_n1554_;
  assign new_n2326_ = new_n7102_ | new_n1553_;
  assign new_n2327_ = new_n7100_ & new_n1500_;
  assign new_n2328_ = new_n7102_ | new_n1499_;
  assign new_n2329_ = new_n2328_ & new_n2326_;
  assign new_n2330_ = new_n2327_ | new_n2325_;
  assign new_n2331_ = new_n7105_ & new_n7001_;
  assign new_n2332_ = new_n7110_ | new_n7007_;
  assign new_n2333_ = new_n7112_ & new_n7113_;
  assign new_n2334_ = new_n7114_ | new_n7115_;
  assign new_n2335_ = new_n7117_ & new_n7113_;
  assign new_n2336_ = new_n7119_ | new_n7115_;
  assign new_n2337_ = new_n7117_ & new_n7112_;
  assign new_n2338_ = new_n7119_ | new_n7114_;
  assign new_n2339_ = new_n2338_ & new_n2336_;
  assign new_n2340_ = new_n2337_ | new_n2335_;
  assign new_n2341_ = new_n2282_ & new_n7012_;
  assign new_n2342_ = new_n7120_ | new_n7014_;
  assign new_n2343_ = new_n7121_ & new_n7122_;
  assign new_n2344_ = new_n7123_ | new_n7124_;
  assign new_n2345_ = new_n7126_ & new_n7122_;
  assign new_n2346_ = new_n7128_ | new_n7124_;
  assign new_n2347_ = new_n7126_ & new_n7121_;
  assign new_n2348_ = new_n7128_ | new_n7123_;
  assign new_n2349_ = new_n2348_ & new_n2346_;
  assign new_n2350_ = new_n2347_ | new_n2345_;
  assign new_n2351_ = new_n7131_ & new_n7135_;
  assign new_n2352_ = new_n7139_ | new_n7143_;
  assign new_n2353_ = new_n7144_ & new_n7135_;
  assign new_n2354_ = new_n7145_ | new_n7143_;
  assign new_n2355_ = new_n1426_ & new_n1422_;
  assign new_n2356_ = new_n1425_ | new_n1421_;
  assign new_n2357_ = new_n7144_ & new_n7147_;
  assign new_n2358_ = new_n7145_ | new_n7150_;
  assign new_n2359_ = new_n7152_ & new_n7153_;
  assign new_n2360_ = new_n7154_ | new_n7155_;
  assign new_n2361_ = new_n7157_ & new_n1369_;
  assign new_n2362_ = new_n7159_ | new_n1370_;
  assign new_n2363_ = new_n7160_ & new_n7161_;
  assign new_n2364_ = new_n7162_ | new_n7163_;
  assign new_n2365_ = new_n7165_ & new_n7161_;
  assign new_n2366_ = new_n7167_ | new_n7163_;
  assign new_n2367_ = new_n7165_ & new_n7160_;
  assign new_n2368_ = new_n7167_ | new_n7162_;
  assign new_n2369_ = new_n2368_ & new_n2366_;
  assign new_n2370_ = new_n2367_ | new_n2365_;
  assign new_n2371_ = new_n7131_ & new_n7147_;
  assign new_n2372_ = new_n7139_ | new_n7150_;
  assign new_n2373_ = new_n7168_ & new_n7169_;
  assign new_n2374_ = new_n7170_ | new_n7171_;
  assign new_n2375_ = new_n7173_ & new_n7164_;
  assign new_n2376_ = new_n7175_ | new_n7166_;
  assign new_n2377_ = new_n7176_ & new_n7177_;
  assign new_n2378_ = new_n7178_ | new_n7179_;
  assign new_n2379_ = new_n7181_ & new_n7177_;
  assign new_n2380_ = new_n7183_ | new_n7179_;
  assign new_n2381_ = new_n7181_ & new_n7176_;
  assign new_n2382_ = new_n7183_ | new_n7178_;
  assign new_n2383_ = new_n2382_ & new_n2380_;
  assign new_n2384_ = new_n2381_ | new_n2379_;
  assign new_n2385_ = new_n6731_ & new_n7148_;
  assign new_n2386_ = new_n6745_ | new_n7151_;
  assign new_n2387_ = new_n7184_ & new_n7185_;
  assign new_n2388_ = new_n7186_ | new_n7187_;
  assign new_n2389_ = new_n7189_ & new_n7185_;
  assign new_n2390_ = new_n7191_ | new_n7187_;
  assign new_n2391_ = new_n7189_ & new_n7184_;
  assign new_n2392_ = new_n7191_ | new_n7186_;
  assign new_n2393_ = new_n2392_ & new_n2390_;
  assign new_n2394_ = new_n2391_ | new_n2389_;
  assign new_n2395_ = new_n7173_ & new_n7169_;
  assign new_n2396_ = new_n7175_ | new_n7171_;
  assign new_n2397_ = new_n7172_ & new_n7168_;
  assign new_n2398_ = new_n7174_ | new_n7170_;
  assign new_n2399_ = new_n2398_ & new_n2396_;
  assign new_n2400_ = new_n2397_ | new_n2395_;
  assign new_n2401_ = new_n7157_ & new_n7153_;
  assign new_n2402_ = new_n7159_ | new_n7155_;
  assign new_n2403_ = new_n7156_ & new_n7152_;
  assign new_n2404_ = new_n7158_ | new_n7154_;
  assign new_n2405_ = new_n2404_ & new_n2402_;
  assign new_n2406_ = new_n2403_ | new_n2401_;
  assign new_n2407_ = new_n7193_ & new_n1293_;
  assign new_n2408_ = new_n7195_ | new_n1294_;
  assign new_n2409_ = new_n7196_ & new_n7197_;
  assign new_n2410_ = new_n7198_ | new_n7199_;
  assign new_n2411_ = new_n7201_ & new_n7197_;
  assign new_n2412_ = new_n7203_ | new_n7199_;
  assign new_n2413_ = new_n7201_ & new_n7196_;
  assign new_n2414_ = new_n7203_ | new_n7198_;
  assign new_n2415_ = new_n2414_ & new_n2412_;
  assign new_n2416_ = new_n2413_ | new_n2411_;
  assign new_n2417_ = new_n7132_ & new_n7205_;
  assign new_n2418_ = new_n7140_ | new_n7208_;
  assign new_n2419_ = new_n7209_ & new_n7210_;
  assign new_n2420_ = new_n7211_ | new_n7212_;
  assign new_n2421_ = new_n7214_ & new_n7200_;
  assign new_n2422_ = new_n7216_ | new_n7202_;
  assign new_n2423_ = new_n7217_ & new_n7218_;
  assign new_n2424_ = new_n7219_ | new_n7220_;
  assign new_n2425_ = new_n7222_ & new_n7218_;
  assign new_n2426_ = new_n7224_ | new_n7220_;
  assign new_n2427_ = new_n7222_ & new_n7217_;
  assign new_n2428_ = new_n7224_ | new_n7219_;
  assign new_n2429_ = new_n2428_ & new_n2426_;
  assign new_n2430_ = new_n2427_ | new_n2425_;
  assign new_n2431_ = new_n6732_ & new_n7205_;
  assign new_n2432_ = new_n6746_ | new_n7208_;
  assign new_n2433_ = new_n7225_ & new_n7226_;
  assign new_n2434_ = new_n7227_ | new_n7228_;
  assign new_n2435_ = new_n7230_ & new_n7221_;
  assign new_n2436_ = new_n7232_ | new_n7223_;
  assign new_n2437_ = new_n7233_ & new_n7234_;
  assign new_n2438_ = new_n7235_ | new_n7236_;
  assign new_n2439_ = new_n7193_ & new_n1377_;
  assign new_n2440_ = new_n7195_ | new_n1378_;
  assign new_n2441_ = new_n7192_ & new_n1330_;
  assign new_n2442_ = new_n7194_ | new_n1329_;
  assign new_n2443_ = new_n2442_ & new_n2440_;
  assign new_n2444_ = new_n2441_ | new_n2439_;
  assign new_n2445_ = new_n1306_ & new_n1243_;
  assign new_n2446_ = new_n1305_ | new_n1244_;
  assign new_n2447_ = new_n7237_ & new_n7238_;
  assign new_n2448_ = new_n7239_ | new_n7240_;
  assign new_n2449_ = new_n7242_ & new_n7238_;
  assign new_n2450_ = new_n7244_ | new_n7240_;
  assign new_n2451_ = new_n7242_ & new_n7237_;
  assign new_n2452_ = new_n7244_ | new_n7239_;
  assign new_n2453_ = new_n2452_ & new_n2450_;
  assign new_n2454_ = new_n2451_ | new_n2449_;
  assign new_n2455_ = new_n7132_ & new_n7246_;
  assign new_n2456_ = new_n7140_ | new_n7249_;
  assign new_n2457_ = new_n7250_ & new_n7251_;
  assign new_n2458_ = new_n7252_ | new_n7253_;
  assign new_n2459_ = new_n7255_ & new_n7251_;
  assign new_n2460_ = new_n7257_ | new_n7253_;
  assign new_n2461_ = new_n7255_ & new_n7250_;
  assign new_n2462_ = new_n7257_ | new_n7252_;
  assign new_n2463_ = new_n2462_ & new_n2460_;
  assign new_n2464_ = new_n2461_ | new_n2459_;
  assign new_n2465_ = new_n7258_ & new_n7259_;
  assign new_n2466_ = new_n7260_ | new_n7261_;
  assign new_n2467_ = new_n7263_ & new_n7258_;
  assign new_n2468_ = new_n7265_ | new_n7260_;
  assign new_n2469_ = new_n7263_ & new_n7259_;
  assign new_n2470_ = new_n7265_ | new_n7261_;
  assign new_n2471_ = new_n2470_ & new_n2468_;
  assign new_n2472_ = new_n2469_ | new_n2467_;
  assign new_n2473_ = new_n7133_ & new_n7267_;
  assign new_n2474_ = new_n7141_ | new_n7270_;
  assign new_n2475_ = new_n7271_ & new_n7272_;
  assign new_n2476_ = new_n7273_ | new_n7274_;
  assign new_n2477_ = new_n7276_ & new_n7262_;
  assign new_n2478_ = new_n7278_ | new_n7264_;
  assign new_n2479_ = new_n7279_ & new_n7280_;
  assign new_n2480_ = new_n7281_ | new_n7282_;
  assign new_n2481_ = new_n7284_ & new_n7280_;
  assign new_n2482_ = new_n7286_ | new_n7282_;
  assign new_n2483_ = new_n7284_ & new_n7279_;
  assign new_n2484_ = new_n7286_ | new_n7281_;
  assign new_n2485_ = new_n2484_ & new_n2482_;
  assign new_n2486_ = new_n2483_ | new_n2481_;
  assign new_n2487_ = new_n6732_ & new_n7267_;
  assign new_n2488_ = new_n6746_ | new_n7270_;
  assign new_n2489_ = new_n7287_ & new_n7288_;
  assign new_n2490_ = new_n7289_ | new_n7290_;
  assign new_n2491_ = new_n7292_ & new_n7288_;
  assign new_n2492_ = new_n7294_ | new_n7290_;
  assign new_n2493_ = new_n7292_ & new_n7287_;
  assign new_n2494_ = new_n7294_ | new_n7289_;
  assign new_n2495_ = new_n2494_ & new_n2492_;
  assign new_n2496_ = new_n2493_ | new_n2491_;
  assign new_n2497_ = new_n7276_ & new_n7272_;
  assign new_n2498_ = new_n7278_ | new_n7274_;
  assign new_n2499_ = new_n7275_ & new_n7271_;
  assign new_n2500_ = new_n7277_ | new_n7273_;
  assign new_n2501_ = new_n2500_ & new_n2498_;
  assign new_n2502_ = new_n2499_ | new_n2497_;
  assign new_n2503_ = new_n1434_ & new_n1428_;
  assign new_n2504_ = new_n1433_ | new_n1427_;
  assign new_n2505_ = new_n7133_ & new_n7296_;
  assign new_n2506_ = new_n7141_ | new_n7299_;
  assign new_n2507_ = new_n7301_ & new_n7302_;
  assign new_n2508_ = new_n7303_ | new_n7304_;
  assign new_n2509_ = new_n7306_ & new_n1371_;
  assign new_n2510_ = new_n7308_ | new_n1372_;
  assign new_n2511_ = new_n7309_ & new_n7310_;
  assign new_n2512_ = new_n7311_ | new_n7312_;
  assign new_n2513_ = new_n7314_ & new_n7310_;
  assign new_n2514_ = new_n7316_ | new_n7312_;
  assign new_n2515_ = new_n7314_ & new_n7309_;
  assign new_n2516_ = new_n7316_ | new_n7311_;
  assign new_n2517_ = new_n2516_ & new_n2514_;
  assign new_n2518_ = new_n2515_ | new_n2513_;
  assign new_n2519_ = new_n6734_ & new_n7296_;
  assign new_n2520_ = new_n6748_ | new_n7299_;
  assign new_n2521_ = new_n7317_ & new_n7318_;
  assign new_n2522_ = new_n7319_ | new_n7320_;
  assign new_n2523_ = new_n7322_ & new_n7313_;
  assign new_n2524_ = new_n7324_ | new_n7315_;
  assign new_n2525_ = new_n7325_ & new_n7326_;
  assign new_n2526_ = new_n7327_ | new_n7328_;
  assign new_n2527_ = new_n7330_ & new_n7326_;
  assign new_n2528_ = new_n7332_ | new_n7328_;
  assign new_n2529_ = new_n7330_ & new_n7325_;
  assign new_n2530_ = new_n7332_ | new_n7327_;
  assign new_n2531_ = new_n2530_ & new_n2528_;
  assign new_n2532_ = new_n2529_ | new_n2527_;
  assign new_n2533_ = new_n7297_ & new_n6761_;
  assign new_n2534_ = new_n7300_ | new_n6775_;
  assign new_n2535_ = new_n7333_ & new_n7334_;
  assign new_n2536_ = new_n7335_ | new_n7336_;
  assign new_n2537_ = new_n7338_ & new_n7334_;
  assign new_n2538_ = new_n7340_ | new_n7336_;
  assign new_n2539_ = new_n7338_ & new_n7333_;
  assign new_n2540_ = new_n7340_ | new_n7335_;
  assign new_n2541_ = new_n2540_ & new_n2538_;
  assign new_n2542_ = new_n2539_ | new_n2537_;
  assign new_n2543_ = new_n7322_ & new_n7318_;
  assign new_n2544_ = new_n7324_ | new_n7320_;
  assign new_n2545_ = new_n7321_ & new_n7317_;
  assign new_n2546_ = new_n7323_ | new_n7319_;
  assign new_n2547_ = new_n2546_ & new_n2544_;
  assign new_n2548_ = new_n2545_ | new_n2543_;
  assign new_n2549_ = new_n7306_ & new_n7302_;
  assign new_n2550_ = new_n7308_ | new_n7304_;
  assign new_n2551_ = new_n7305_ & new_n7301_;
  assign new_n2552_ = new_n7307_ | new_n7303_;
  assign new_n2553_ = new_n2552_ & new_n2550_;
  assign new_n2554_ = new_n2551_ | new_n2549_;
  assign new_n2555_ = new_n7342_ & new_n1295_;
  assign new_n2556_ = new_n7344_ | new_n1296_;
  assign new_n2557_ = new_n7345_ & new_n7346_;
  assign new_n2558_ = new_n7347_ | new_n7348_;
  assign new_n2559_ = new_n7350_ & new_n7346_;
  assign new_n2560_ = new_n7352_ | new_n7348_;
  assign new_n2561_ = new_n7350_ & new_n7345_;
  assign new_n2562_ = new_n7352_ | new_n7347_;
  assign new_n2563_ = new_n2562_ & new_n2560_;
  assign new_n2564_ = new_n2561_ | new_n2559_;
  assign new_n2565_ = new_n6734_ & new_n7354_;
  assign new_n2566_ = new_n6748_ | new_n7357_;
  assign new_n2567_ = new_n7358_ & new_n7359_;
  assign new_n2568_ = new_n7360_ | new_n7361_;
  assign new_n2569_ = new_n7363_ & new_n7349_;
  assign new_n2570_ = new_n7365_ | new_n7351_;
  assign new_n2571_ = new_n7366_ & new_n7367_;
  assign new_n2572_ = new_n7368_ | new_n7369_;
  assign new_n2573_ = new_n7371_ & new_n7367_;
  assign new_n2574_ = new_n7373_ | new_n7369_;
  assign new_n2575_ = new_n7371_ & new_n7366_;
  assign new_n2576_ = new_n7373_ | new_n7368_;
  assign new_n2577_ = new_n2576_ & new_n2574_;
  assign new_n2578_ = new_n2575_ | new_n2573_;
  assign new_n2579_ = new_n7354_ & new_n6763_;
  assign new_n2580_ = new_n7357_ | new_n6777_;
  assign new_n2581_ = new_n7374_ & new_n7375_;
  assign new_n2582_ = new_n7376_ | new_n7377_;
  assign new_n2583_ = new_n7379_ & new_n7370_;
  assign new_n2584_ = new_n7381_ | new_n7372_;
  assign new_n2585_ = new_n7382_ & new_n7383_;
  assign new_n2586_ = new_n7384_ | new_n7385_;
  assign new_n2587_ = new_n7342_ & new_n1379_;
  assign new_n2588_ = new_n7344_ | new_n1380_;
  assign new_n2589_ = new_n7341_ & new_n1332_;
  assign new_n2590_ = new_n7343_ | new_n1331_;
  assign new_n2591_ = new_n2590_ & new_n2588_;
  assign new_n2592_ = new_n2589_ | new_n2587_;
  assign new_n2593_ = new_n1308_ & new_n1245_;
  assign new_n2594_ = new_n1307_ | new_n1246_;
  assign new_n2595_ = new_n7386_ & new_n7387_;
  assign new_n2596_ = new_n7388_ | new_n7389_;
  assign new_n2597_ = new_n7391_ & new_n7387_;
  assign new_n2598_ = new_n7393_ | new_n7389_;
  assign new_n2599_ = new_n7391_ & new_n7386_;
  assign new_n2600_ = new_n7393_ | new_n7388_;
  assign new_n2601_ = new_n2600_ & new_n2598_;
  assign new_n2602_ = new_n2599_ | new_n2597_;
  assign new_n2603_ = new_n6733_ & new_n7395_;
  assign new_n2604_ = new_n6747_ | new_n7398_;
  assign new_n2605_ = new_n7399_ & new_n7400_;
  assign new_n2606_ = new_n7401_ | new_n7402_;
  assign new_n2607_ = new_n7404_ & new_n7400_;
  assign new_n2608_ = new_n7406_ | new_n7402_;
  assign new_n2609_ = new_n7404_ & new_n7399_;
  assign new_n2610_ = new_n7406_ | new_n7401_;
  assign new_n2611_ = new_n2610_ & new_n2608_;
  assign new_n2612_ = new_n2609_ | new_n2607_;
  assign new_n2613_ = new_n7407_ & new_n7408_;
  assign new_n2614_ = new_n7409_ | new_n7410_;
  assign new_n2615_ = new_n7412_ & new_n7407_;
  assign new_n2616_ = new_n7414_ | new_n7409_;
  assign new_n2617_ = new_n7412_ & new_n7408_;
  assign new_n2618_ = new_n7414_ | new_n7410_;
  assign new_n2619_ = new_n2618_ & new_n2616_;
  assign new_n2620_ = new_n2617_ | new_n2615_;
  assign new_n2621_ = new_n6736_ & new_n7416_;
  assign new_n2622_ = new_n6750_ | new_n7419_;
  assign new_n2623_ = new_n7420_ & new_n7421_;
  assign new_n2624_ = new_n7422_ | new_n7423_;
  assign new_n2625_ = new_n7425_ & new_n7411_;
  assign new_n2626_ = new_n7427_ | new_n7413_;
  assign new_n2627_ = new_n7428_ & new_n7429_;
  assign new_n2628_ = new_n7430_ | new_n7431_;
  assign new_n2629_ = new_n7433_ & new_n7429_;
  assign new_n2630_ = new_n7435_ | new_n7431_;
  assign new_n2631_ = new_n7433_ & new_n7428_;
  assign new_n2632_ = new_n7435_ | new_n7430_;
  assign new_n2633_ = new_n2632_ & new_n2630_;
  assign new_n2634_ = new_n2631_ | new_n2629_;
  assign new_n2635_ = new_n7416_ & new_n6763_;
  assign new_n2636_ = new_n7419_ | new_n6777_;
  assign new_n2637_ = new_n7436_ & new_n7437_;
  assign new_n2638_ = new_n7438_ | new_n7439_;
  assign new_n2639_ = new_n7441_ & new_n7437_;
  assign new_n2640_ = new_n7443_ | new_n7439_;
  assign new_n2641_ = new_n7441_ & new_n7436_;
  assign new_n2642_ = new_n7443_ | new_n7438_;
  assign new_n2643_ = new_n2642_ & new_n2640_;
  assign new_n2644_ = new_n2641_ | new_n2639_;
  assign new_n2645_ = new_n7425_ & new_n7421_;
  assign new_n2646_ = new_n7427_ | new_n7423_;
  assign new_n2647_ = new_n7424_ & new_n7420_;
  assign new_n2648_ = new_n7426_ | new_n7422_;
  assign new_n2649_ = new_n2648_ & new_n2646_;
  assign new_n2650_ = new_n2647_ | new_n2645_;
  assign new_n2651_ = new_n1436_ & new_n1430_;
  assign new_n2652_ = new_n1435_ | new_n1429_;
  assign new_n2653_ = new_n6736_ & new_n7445_;
  assign new_n2654_ = new_n6750_ | new_n7447_;
  assign new_n2655_ = new_n7449_ & new_n7450_;
  assign new_n2656_ = new_n7451_ | new_n7452_;
  assign new_n2657_ = new_n7454_ & new_n1373_;
  assign new_n2658_ = new_n7456_ | new_n1374_;
  assign new_n2659_ = new_n7457_ & new_n7458_;
  assign new_n2660_ = new_n7459_ | new_n7460_;
  assign new_n2661_ = new_n7462_ & new_n7458_;
  assign new_n2662_ = new_n7464_ | new_n7460_;
  assign new_n2663_ = new_n7462_ & new_n7457_;
  assign new_n2664_ = new_n7464_ | new_n7459_;
  assign new_n2665_ = new_n2664_ & new_n2662_;
  assign new_n2666_ = new_n2663_ | new_n2661_;
  assign new_n2667_ = new_n7445_ & new_n6764_;
  assign new_n2668_ = new_n7447_ | new_n6778_;
  assign new_n2669_ = new_n7465_ & new_n7466_;
  assign new_n2670_ = new_n7467_ | new_n7468_;
  assign new_n2671_ = new_n7470_ & new_n7461_;
  assign new_n2672_ = new_n7472_ | new_n7463_;
  assign new_n2673_ = new_n7473_ & new_n7474_;
  assign new_n2674_ = new_n7475_ | new_n7476_;
  assign new_n2675_ = new_n7478_ & new_n7474_;
  assign new_n2676_ = new_n7480_ | new_n7476_;
  assign new_n2677_ = new_n7478_ & new_n7473_;
  assign new_n2678_ = new_n7480_ | new_n7475_;
  assign new_n2679_ = new_n2678_ & new_n2676_;
  assign new_n2680_ = new_n2677_ | new_n2675_;
  assign new_n2681_ = new_n7444_ & new_n6808_;
  assign new_n2682_ = new_n7448_ | new_n6818_;
  assign new_n2683_ = new_n7481_ & new_n7482_;
  assign new_n2684_ = new_n7483_ | new_n7484_;
  assign new_n2685_ = new_n7486_ & new_n7482_;
  assign new_n2686_ = new_n7488_ | new_n7484_;
  assign new_n2687_ = new_n7486_ & new_n7481_;
  assign new_n2688_ = new_n7488_ | new_n7483_;
  assign new_n2689_ = new_n2688_ & new_n2686_;
  assign new_n2690_ = new_n2687_ | new_n2685_;
  assign new_n2691_ = new_n7470_ & new_n7466_;
  assign new_n2692_ = new_n7472_ | new_n7468_;
  assign new_n2693_ = new_n7469_ & new_n7465_;
  assign new_n2694_ = new_n7471_ | new_n7467_;
  assign new_n2695_ = new_n2694_ & new_n2692_;
  assign new_n2696_ = new_n2693_ | new_n2691_;
  assign new_n2697_ = new_n7454_ & new_n7450_;
  assign new_n2698_ = new_n7456_ | new_n7452_;
  assign new_n2699_ = new_n7453_ & new_n7449_;
  assign new_n2700_ = new_n7455_ | new_n7451_;
  assign new_n2701_ = new_n2700_ & new_n2698_;
  assign new_n2702_ = new_n2699_ | new_n2697_;
  assign new_n2703_ = new_n7490_ & new_n1297_;
  assign new_n2704_ = new_n7492_ | new_n1298_;
  assign new_n2705_ = new_n7493_ & new_n7494_;
  assign new_n2706_ = new_n7495_ | new_n7496_;
  assign new_n2707_ = new_n7498_ & new_n7494_;
  assign new_n2708_ = new_n7500_ | new_n7496_;
  assign new_n2709_ = new_n7498_ & new_n7493_;
  assign new_n2710_ = new_n7500_ | new_n7495_;
  assign new_n2711_ = new_n2710_ & new_n2708_;
  assign new_n2712_ = new_n2709_ | new_n2707_;
  assign new_n2713_ = new_n7502_ & new_n6764_;
  assign new_n2714_ = new_n7504_ | new_n6778_;
  assign new_n2715_ = new_n7505_ & new_n7506_;
  assign new_n2716_ = new_n7507_ | new_n7508_;
  assign new_n2717_ = new_n7510_ & new_n7497_;
  assign new_n2718_ = new_n7512_ | new_n7499_;
  assign new_n2719_ = new_n7513_ & new_n7514_;
  assign new_n2720_ = new_n7515_ | new_n7516_;
  assign new_n2721_ = new_n7518_ & new_n7514_;
  assign new_n2722_ = new_n7520_ | new_n7516_;
  assign new_n2723_ = new_n7518_ & new_n7513_;
  assign new_n2724_ = new_n7520_ | new_n7515_;
  assign new_n2725_ = new_n2724_ & new_n2722_;
  assign new_n2726_ = new_n2723_ | new_n2721_;
  assign new_n2727_ = new_n7502_ & new_n6808_;
  assign new_n2728_ = new_n7504_ | new_n6818_;
  assign new_n2729_ = new_n7521_ & new_n7522_;
  assign new_n2730_ = new_n7523_ | new_n7524_;
  assign new_n2731_ = new_n7526_ & new_n7517_;
  assign new_n2732_ = new_n7528_ | new_n7519_;
  assign new_n2733_ = new_n7529_ & new_n7530_;
  assign new_n2734_ = new_n7531_ | new_n7532_;
  assign new_n2735_ = new_n7533_ & new_n7534_;
  assign new_n2736_ = new_n7535_ | new_n7536_;
  assign new_n2737_ = new_n7538_ & new_n7533_;
  assign new_n2738_ = new_n7540_ | new_n7535_;
  assign new_n2739_ = new_n7538_ & new_n7534_;
  assign new_n2740_ = new_n7540_ | new_n7536_;
  assign new_n2741_ = new_n2740_ & new_n2738_;
  assign new_n2742_ = new_n2739_ | new_n2737_;
  assign new_n2743_ = new_n7542_ & new_n6767_;
  assign new_n2744_ = new_n7544_ | new_n6781_;
  assign new_n2745_ = new_n7545_ & new_n7546_;
  assign new_n2746_ = new_n7547_ | new_n7548_;
  assign new_n2747_ = new_n7550_ & new_n7546_;
  assign new_n2748_ = new_n7552_ | new_n7548_;
  assign new_n2749_ = new_n7550_ & new_n7545_;
  assign new_n2750_ = new_n7552_ | new_n7547_;
  assign new_n2751_ = new_n2750_ & new_n2748_;
  assign new_n2752_ = new_n2749_ | new_n2747_;
  assign new_n2753_ = new_n6910_ & new_n6898_;
  assign new_n2754_ = new_n6912_ | new_n6900_;
  assign new_n2755_ = new_n7553_ & new_n7554_;
  assign new_n2756_ = new_n7555_ | new_n7556_;
  assign new_n2757_ = new_n7558_ & new_n7554_;
  assign new_n2758_ = new_n7560_ | new_n7556_;
  assign new_n2759_ = new_n7558_ & new_n7553_;
  assign new_n2760_ = new_n7560_ | new_n7555_;
  assign new_n2761_ = new_n2760_ & new_n2758_;
  assign new_n2762_ = new_n2759_ | new_n2757_;
  assign new_n2763_ = new_n6903_ & new_n6810_;
  assign new_n2764_ = new_n6905_ | new_n6820_;
  assign new_n2765_ = new_n7561_ & new_n7562_;
  assign new_n2766_ = new_n7563_ | new_n7564_;
  assign new_n2767_ = new_n7566_ & new_n7562_;
  assign new_n2768_ = new_n7568_ | new_n7564_;
  assign new_n2769_ = new_n7566_ & new_n7561_;
  assign new_n2770_ = new_n7568_ | new_n7563_;
  assign new_n2771_ = new_n2770_ & new_n2768_;
  assign new_n2772_ = new_n2769_ | new_n2767_;
  assign new_n2773_ = new_n6926_ & new_n6918_;
  assign new_n2774_ = new_n6928_ | new_n6920_;
  assign new_n2775_ = new_n7569_ & new_n7570_;
  assign new_n2776_ = new_n7571_ | new_n7572_;
  assign new_n2777_ = new_n7574_ & new_n7570_;
  assign new_n2778_ = new_n7576_ | new_n7572_;
  assign new_n2779_ = new_n7574_ & new_n7569_;
  assign new_n2780_ = new_n7576_ | new_n7571_;
  assign new_n2781_ = new_n2780_ & new_n2778_;
  assign new_n2782_ = new_n2779_ | new_n2777_;
  assign new_n2783_ = new_n6836_ & new_n6884_;
  assign new_n2784_ = new_n6838_ | new_n6890_;
  assign new_n2785_ = new_n7577_ & new_n7578_;
  assign new_n2786_ = new_n7579_ | new_n7580_;
  assign new_n2787_ = new_n7582_ & new_n7578_;
  assign new_n2788_ = new_n7584_ | new_n7580_;
  assign new_n2789_ = new_n7582_ & new_n7577_;
  assign new_n2790_ = new_n7584_ | new_n7579_;
  assign new_n2791_ = new_n2790_ & new_n2788_;
  assign new_n2792_ = new_n2789_ | new_n2787_;
  assign new_n2793_ = new_n2244_ & new_n6935_;
  assign new_n2794_ = new_n7585_ | new_n6937_;
  assign new_n2795_ = new_n7586_ & new_n7587_;
  assign new_n2796_ = new_n2793_ | new_n2791_;
  assign new_n2797_ = new_n7588_ & new_n7587_;
  assign new_n2798_ = new_n7588_ & new_n7586_;
  assign new_n2799_ = new_n2798_ | new_n2797_;
  assign new_n2800_ = new_n7589_ & new_n2324_;
  assign new_n2801_ = new_n2349_ | new_n7590_;
  assign new_n2802_ = new_n6866_ & new_n7594_;
  assign new_n2803_ = new_n6875_ | new_n7607_;
  assign new_n2804_ = new_n7618_ & new_n1477_;
  assign new_n2805_ = new_n7620_ | new_n1478_;
  assign new_n2806_ = new_n7618_ & new_n1408_;
  assign new_n2807_ = new_n7620_ | new_n1407_;
  assign new_n2808_ = new_n2807_ & new_n2805_;
  assign new_n2809_ = new_n2806_ | new_n2804_;
  assign new_n2810_ = new_n7052_ & new_n1391_;
  assign new_n2811_ = new_n7054_ | new_n1392_;
  assign new_n2812_ = new_n7621_ & new_n7622_;
  assign new_n2813_ = new_n7623_ | new_n7624_;
  assign new_n2814_ = new_n7626_ & new_n7622_;
  assign new_n2815_ = new_n7628_ | new_n7624_;
  assign new_n2816_ = new_n7626_ & new_n7621_;
  assign new_n2817_ = new_n7628_ | new_n7623_;
  assign new_n2818_ = new_n2817_ & new_n2815_;
  assign new_n2819_ = new_n2816_ | new_n2814_;
  assign new_n2820_ = new_n6943_ & new_n7631_;
  assign new_n2821_ = new_n6956_ | new_n7635_;
  assign new_n2822_ = new_n7637_ & new_n7638_;
  assign new_n2823_ = new_n7639_ | new_n7640_;
  assign new_n2824_ = new_n7642_ & new_n7638_;
  assign new_n2825_ = new_n7644_ | new_n7640_;
  assign new_n2826_ = new_n7642_ & new_n7637_;
  assign new_n2827_ = new_n7644_ | new_n7639_;
  assign new_n2828_ = new_n2827_ & new_n2825_;
  assign new_n2829_ = new_n2826_ | new_n2824_;
  assign new_n2830_ = new_n7068_ & new_n7060_;
  assign new_n2831_ = new_n7070_ | new_n7062_;
  assign new_n2832_ = new_n7645_ & new_n7646_;
  assign new_n2833_ = new_n7647_ | new_n7648_;
  assign new_n2834_ = new_n7650_ & new_n7646_;
  assign new_n2835_ = new_n7652_ | new_n7648_;
  assign new_n2836_ = new_n7650_ & new_n7645_;
  assign new_n2837_ = new_n7652_ | new_n7647_;
  assign new_n2838_ = new_n2837_ & new_n2835_;
  assign new_n2839_ = new_n2836_ | new_n2834_;
  assign new_n2840_ = new_n6970_ & new_n7019_;
  assign new_n2841_ = new_n6974_ | new_n7034_;
  assign new_n2842_ = new_n7653_ & new_n7654_;
  assign new_n2843_ = new_n7655_ | new_n7656_;
  assign new_n2844_ = new_n7658_ & new_n7654_;
  assign new_n2845_ = new_n7660_ | new_n7656_;
  assign new_n2846_ = new_n7658_ & new_n7653_;
  assign new_n2847_ = new_n7660_ | new_n7655_;
  assign new_n2848_ = new_n2847_ & new_n2845_;
  assign new_n2849_ = new_n2846_ | new_n2844_;
  assign new_n2850_ = new_n2322_ & new_n7077_;
  assign new_n2851_ = new_n7661_ | new_n7079_;
  assign new_n2852_ = new_n7662_ & new_n7663_;
  assign new_n2853_ = new_n7664_ | new_n7665_;
  assign new_n2854_ = new_n7667_ & new_n7663_;
  assign new_n2855_ = new_n7669_ | new_n7665_;
  assign new_n2856_ = new_n7667_ & new_n7662_;
  assign new_n2857_ = new_n7669_ | new_n7664_;
  assign new_n2858_ = new_n2857_ & new_n2855_;
  assign new_n2859_ = new_n2856_ | new_n2854_;
  assign new_n2860_ = new_n7673_ & new_n6997_;
  assign new_n2861_ = new_n7688_ | new_n7003_;
  assign new_n2862_ = new_n7700_ & new_n2803_;
  assign new_n2863_ = new_n2858_ | new_n7701_;
  assign new_n2864_ = new_n1586_ & new_n1578_;
  assign new_n2865_ = new_n1585_ | new_n1577_;
  assign new_n2866_ = new_n7704_ & new_n7000_;
  assign new_n2867_ = new_n7710_ | new_n7006_;
  assign new_n2868_ = new_n7712_ & new_n7713_;
  assign new_n2869_ = new_n7714_ | new_n7715_;
  assign new_n2870_ = new_n7717_ & new_n7713_;
  assign new_n2871_ = new_n7719_ | new_n7715_;
  assign new_n2872_ = new_n7717_ & new_n7712_;
  assign new_n2873_ = new_n7719_ | new_n7714_;
  assign new_n2874_ = new_n2873_ & new_n2871_;
  assign new_n2875_ = new_n2872_ | new_n2870_;
  assign new_n2876_ = new_n7116_ & new_n7099_;
  assign new_n2877_ = new_n7118_ | new_n7101_;
  assign new_n2878_ = new_n7720_ & new_n7721_;
  assign new_n2879_ = new_n7722_ | new_n7723_;
  assign new_n2880_ = new_n7725_ & new_n7721_;
  assign new_n2881_ = new_n7727_ | new_n7723_;
  assign new_n2882_ = new_n7725_ & new_n7720_;
  assign new_n2883_ = new_n7727_ | new_n7722_;
  assign new_n2884_ = new_n2883_ & new_n2881_;
  assign new_n2885_ = new_n2882_ | new_n2880_;
  assign new_n2886_ = new_n7086_ & new_n7105_;
  assign new_n2887_ = new_n7094_ | new_n7110_;
  assign new_n2888_ = new_n7728_ & new_n7729_;
  assign new_n2889_ = new_n7730_ | new_n7731_;
  assign new_n2890_ = new_n7733_ & new_n7729_;
  assign new_n2891_ = new_n7735_ | new_n7731_;
  assign new_n2892_ = new_n7733_ & new_n7728_;
  assign new_n2893_ = new_n7735_ | new_n7730_;
  assign new_n2894_ = new_n2893_ & new_n2891_;
  assign new_n2895_ = new_n2892_ | new_n2890_;
  assign new_n2896_ = new_n2801_ & new_n7125_;
  assign new_n2897_ = new_n7736_ | new_n7127_;
  assign new_n2898_ = new_n7737_ & new_n7738_;
  assign new_n2899_ = new_n7739_ | new_n7740_;
  assign new_n2900_ = new_n7742_ & new_n7738_;
  assign new_n2901_ = new_n7744_ | new_n7740_;
  assign new_n2902_ = new_n7742_ & new_n7737_;
  assign new_n2903_ = new_n7744_ | new_n7739_;
  assign new_n2904_ = new_n2903_ & new_n2901_;
  assign new_n2905_ = new_n2902_ | new_n2900_;
  assign new_n2906_ = new_n7745_ & new_n2861_;
  assign new_n2907_ = new_n2904_ | new_n7746_;
  assign new_n2908_ = new_n7748_ | new_n2795_;
  assign new_n2909_ = new_n6737_ & new_n7136_;
  assign new_n2910_ = new_n6751_ | new_n7142_;
  assign new_n2911_ = new_n7188_ & new_n7180_;
  assign new_n2912_ = new_n7190_ | new_n7182_;
  assign new_n2913_ = new_n2911_ | new_n2909_;
  assign new_n2914_ = new_n7214_ & new_n7210_;
  assign new_n2915_ = new_n7216_ | new_n7212_;
  assign new_n2916_ = new_n7213_ & new_n7209_;
  assign new_n2917_ = new_n7215_ | new_n7211_;
  assign new_n2918_ = new_n2917_ & new_n2915_;
  assign new_n2919_ = new_n2916_ | new_n2914_;
  assign new_n2920_ = new_n7254_ & new_n7241_;
  assign new_n2921_ = new_n7256_ | new_n7243_;
  assign new_n2922_ = new_n7749_ & new_n7750_;
  assign new_n2923_ = new_n7751_ | new_n7752_;
  assign new_n2924_ = new_n7754_ & new_n7750_;
  assign new_n2925_ = new_n7756_ | new_n7752_;
  assign new_n2926_ = new_n7754_ & new_n7749_;
  assign new_n2927_ = new_n7756_ | new_n7751_;
  assign new_n2928_ = new_n2927_ & new_n2925_;
  assign new_n2929_ = new_n2926_ | new_n2924_;
  assign new_n2930_ = new_n6737_ & new_n7246_;
  assign new_n2931_ = new_n6751_ | new_n7249_;
  assign new_n2932_ = new_n7757_ & new_n7758_;
  assign new_n2933_ = new_n7759_ | new_n7760_;
  assign new_n2934_ = new_n7762_ & new_n7758_;
  assign new_n2935_ = new_n7764_ | new_n7760_;
  assign new_n2936_ = new_n7762_ & new_n7757_;
  assign new_n2937_ = new_n7764_ | new_n7759_;
  assign new_n2938_ = new_n2937_ & new_n2935_;
  assign new_n2939_ = new_n2936_ | new_n2934_;
  assign new_n2940_ = new_n7291_ & new_n7283_;
  assign new_n2941_ = new_n7293_ | new_n7285_;
  assign new_n2942_ = new_n7765_ & new_n7766_;
  assign new_n2943_ = new_n7767_ | new_n7768_;
  assign new_n2944_ = new_n7770_ & new_n7766_;
  assign new_n2945_ = new_n7772_ | new_n7768_;
  assign new_n2946_ = new_n7770_ & new_n7765_;
  assign new_n2947_ = new_n7772_ | new_n7767_;
  assign new_n2948_ = new_n2947_ & new_n2945_;
  assign new_n2949_ = new_n2946_ | new_n2944_;
  assign new_n2950_ = new_n7268_ & new_n6767_;
  assign new_n2951_ = new_n7269_ | new_n6781_;
  assign new_n2952_ = new_n7773_ & new_n7774_;
  assign new_n2953_ = new_n7775_ | new_n7776_;
  assign new_n2954_ = new_n7778_ & new_n7774_;
  assign new_n2955_ = new_n7780_ | new_n7776_;
  assign new_n2956_ = new_n7778_ & new_n7773_;
  assign new_n2957_ = new_n7780_ | new_n7775_;
  assign new_n2958_ = new_n2957_ & new_n2955_;
  assign new_n2959_ = new_n2956_ | new_n2954_;
  assign new_n2960_ = new_n7337_ & new_n7329_;
  assign new_n2961_ = new_n7339_ | new_n7331_;
  assign new_n2962_ = new_n2960_ | new_n2958_;
  assign new_n2963_ = new_n7363_ & new_n7359_;
  assign new_n2964_ = new_n7365_ | new_n7361_;
  assign new_n2965_ = new_n7362_ & new_n7358_;
  assign new_n2966_ = new_n7364_ | new_n7360_;
  assign new_n2967_ = new_n2966_ & new_n2964_;
  assign new_n2968_ = new_n2965_ | new_n2963_;
  assign new_n2969_ = new_n7403_ & new_n7390_;
  assign new_n2970_ = new_n7405_ | new_n7392_;
  assign new_n2971_ = new_n7781_ & new_n7782_;
  assign new_n2972_ = new_n7783_ | new_n7784_;
  assign new_n2973_ = new_n7786_ & new_n7782_;
  assign new_n2974_ = new_n7788_ | new_n7784_;
  assign new_n2975_ = new_n7786_ & new_n7781_;
  assign new_n2976_ = new_n7788_ | new_n7783_;
  assign new_n2977_ = new_n2976_ & new_n2974_;
  assign new_n2978_ = new_n2975_ | new_n2973_;
  assign new_n2979_ = new_n7395_ & new_n6768_;
  assign new_n2980_ = new_n7398_ | new_n6782_;
  assign new_n2981_ = new_n7789_ & new_n7790_;
  assign new_n2982_ = new_n7791_ | new_n7792_;
  assign new_n2983_ = new_n7794_ & new_n7790_;
  assign new_n2984_ = new_n7796_ | new_n7792_;
  assign new_n2985_ = new_n7794_ & new_n7789_;
  assign new_n2986_ = new_n7796_ | new_n7791_;
  assign new_n2987_ = new_n2986_ & new_n2984_;
  assign new_n2988_ = new_n2985_ | new_n2983_;
  assign new_n2989_ = new_n7440_ & new_n7432_;
  assign new_n2990_ = new_n7442_ | new_n7434_;
  assign new_n2991_ = new_n7797_ & new_n7798_;
  assign new_n2992_ = new_n7799_ | new_n7800_;
  assign new_n2993_ = new_n7802_ & new_n7798_;
  assign new_n2994_ = new_n7804_ | new_n7800_;
  assign new_n2995_ = new_n7802_ & new_n7797_;
  assign new_n2996_ = new_n7804_ | new_n7799_;
  assign new_n2997_ = new_n2996_ & new_n2994_;
  assign new_n2998_ = new_n2995_ | new_n2993_;
  assign new_n2999_ = new_n7417_ & new_n6810_;
  assign new_n3000_ = new_n7418_ | new_n6820_;
  assign new_n3001_ = new_n7805_ & new_n7806_;
  assign new_n3002_ = new_n7807_ | new_n7808_;
  assign new_n3003_ = new_n7810_ & new_n7806_;
  assign new_n3004_ = new_n7812_ | new_n7808_;
  assign new_n3005_ = new_n7810_ & new_n7805_;
  assign new_n3006_ = new_n7812_ | new_n7807_;
  assign new_n3007_ = new_n3006_ & new_n3004_;
  assign new_n3008_ = new_n3005_ | new_n3003_;
  assign new_n3009_ = new_n7485_ & new_n7477_;
  assign new_n3010_ = new_n7487_ | new_n7479_;
  assign new_n3011_ = new_n3009_ | new_n3007_;
  assign new_n3012_ = new_n7510_ & new_n7506_;
  assign new_n3013_ = new_n7512_ | new_n7508_;
  assign new_n3014_ = new_n7509_ & new_n7505_;
  assign new_n3015_ = new_n7511_ | new_n7507_;
  assign new_n3016_ = new_n3015_ & new_n3013_;
  assign new_n3017_ = new_n3014_ | new_n3012_;
  assign new_n3018_ = new_n7490_ & new_n1381_;
  assign new_n3019_ = new_n7492_ | new_n1382_;
  assign new_n3020_ = new_n7489_ & new_n1334_;
  assign new_n3021_ = new_n7491_ | new_n1333_;
  assign new_n3022_ = new_n3021_ & new_n3019_;
  assign new_n3023_ = new_n3020_ | new_n3018_;
  assign new_n3024_ = new_n1310_ & new_n1247_;
  assign new_n3025_ = new_n1309_ | new_n1248_;
  assign new_n3026_ = new_n7813_ & new_n7814_;
  assign new_n3027_ = new_n7815_ | new_n7816_;
  assign new_n3028_ = new_n7818_ & new_n7814_;
  assign new_n3029_ = new_n7820_ | new_n7816_;
  assign new_n3030_ = new_n7818_ & new_n7813_;
  assign new_n3031_ = new_n7820_ | new_n7815_;
  assign new_n3032_ = new_n3031_ & new_n3029_;
  assign new_n3033_ = new_n3030_ | new_n3028_;
  assign new_n3034_ = new_n7822_ & new_n6768_;
  assign new_n3035_ = new_n7824_ | new_n6782_;
  assign new_n3036_ = new_n7825_ & new_n7826_;
  assign new_n3037_ = new_n7827_ | new_n7828_;
  assign new_n3038_ = new_n7830_ & new_n7817_;
  assign new_n3039_ = new_n7832_ | new_n7819_;
  assign new_n3040_ = new_n7833_ & new_n7834_;
  assign new_n3041_ = new_n7835_ | new_n7836_;
  assign new_n3042_ = new_n7838_ & new_n7834_;
  assign new_n3043_ = new_n7840_ | new_n7836_;
  assign new_n3044_ = new_n7838_ & new_n7833_;
  assign new_n3045_ = new_n7840_ | new_n7835_;
  assign new_n3046_ = new_n3045_ & new_n3043_;
  assign new_n3047_ = new_n3044_ | new_n3042_;
  assign new_n3048_ = new_n7822_ & new_n6809_;
  assign new_n3049_ = new_n7824_ | new_n6819_;
  assign new_n3050_ = new_n7841_ & new_n7842_;
  assign new_n3051_ = new_n7843_ | new_n7844_;
  assign new_n3052_ = new_n7846_ & new_n7842_;
  assign new_n3053_ = new_n7848_ | new_n7844_;
  assign new_n3054_ = new_n7846_ & new_n7841_;
  assign new_n3055_ = new_n7848_ | new_n7843_;
  assign new_n3056_ = new_n3055_ & new_n3053_;
  assign new_n3057_ = new_n3054_ | new_n3052_;
  assign new_n3058_ = new_n7830_ & new_n7826_;
  assign new_n3059_ = new_n7832_ | new_n7828_;
  assign new_n3060_ = new_n7829_ & new_n7825_;
  assign new_n3061_ = new_n7831_ | new_n7827_;
  assign new_n3062_ = new_n3061_ & new_n3059_;
  assign new_n3063_ = new_n3060_ | new_n3058_;
  assign new_n3064_ = new_n7549_ & new_n7537_;
  assign new_n3065_ = new_n7551_ | new_n7539_;
  assign new_n3066_ = new_n7849_ & new_n7850_;
  assign new_n3067_ = new_n7851_ | new_n7852_;
  assign new_n3068_ = new_n7854_ & new_n7850_;
  assign new_n3069_ = new_n7856_ | new_n7852_;
  assign new_n3070_ = new_n7854_ & new_n7849_;
  assign new_n3071_ = new_n7856_ | new_n7851_;
  assign new_n3072_ = new_n3071_ & new_n3069_;
  assign new_n3073_ = new_n3070_ | new_n3068_;
  assign new_n3074_ = new_n7542_ & new_n6812_;
  assign new_n3075_ = new_n7544_ | new_n6822_;
  assign new_n3076_ = new_n7857_ & new_n7858_;
  assign new_n3077_ = new_n7859_ | new_n7860_;
  assign new_n3078_ = new_n7862_ & new_n7853_;
  assign new_n3079_ = new_n7864_ | new_n7855_;
  assign new_n3080_ = new_n7865_ & new_n7866_;
  assign new_n3081_ = new_n7867_ | new_n7868_;
  assign new_n3082_ = new_n7870_ & new_n7866_;
  assign new_n3083_ = new_n7872_ | new_n7868_;
  assign new_n3084_ = new_n7870_ & new_n7865_;
  assign new_n3085_ = new_n7872_ | new_n7867_;
  assign new_n3086_ = new_n3085_ & new_n3083_;
  assign new_n3087_ = new_n3084_ | new_n3082_;
  assign new_n3088_ = new_n7541_ & new_n6885_;
  assign new_n3089_ = new_n7543_ | new_n6891_;
  assign new_n3090_ = new_n7873_ & new_n7874_;
  assign new_n3091_ = new_n7875_ | new_n7876_;
  assign new_n3092_ = new_n7878_ & new_n7874_;
  assign new_n3093_ = new_n7880_ | new_n7876_;
  assign new_n3094_ = new_n7878_ & new_n7873_;
  assign new_n3095_ = new_n7880_ | new_n7875_;
  assign new_n3096_ = new_n3095_ & new_n3093_;
  assign new_n3097_ = new_n3094_ | new_n3092_;
  assign new_n3098_ = new_n7862_ & new_n7858_;
  assign new_n3099_ = new_n7864_ | new_n7860_;
  assign new_n3100_ = new_n7861_ & new_n7857_;
  assign new_n3101_ = new_n7863_ | new_n7859_;
  assign new_n3102_ = new_n3101_ & new_n3099_;
  assign new_n3103_ = new_n3100_ | new_n3098_;
  assign new_n3104_ = new_n7565_ & new_n7557_;
  assign new_n3105_ = new_n7567_ | new_n7559_;
  assign new_n3106_ = new_n7881_ & new_n7882_;
  assign new_n3107_ = new_n7883_ | new_n7884_;
  assign new_n3108_ = new_n7886_ & new_n7882_;
  assign new_n3109_ = new_n7888_ | new_n7884_;
  assign new_n3110_ = new_n7886_ & new_n7881_;
  assign new_n3111_ = new_n7888_ | new_n7883_;
  assign new_n3112_ = new_n3111_ & new_n3109_;
  assign new_n3113_ = new_n3110_ | new_n3108_;
  assign new_n3114_ = new_n6902_ & new_n6885_;
  assign new_n3115_ = new_n6904_ | new_n6891_;
  assign new_n3116_ = new_n7889_ & new_n7890_;
  assign new_n3117_ = new_n7891_ | new_n7892_;
  assign new_n3118_ = new_n7894_ & new_n7885_;
  assign new_n3119_ = new_n7896_ | new_n7887_;
  assign new_n3120_ = new_n3118_ | new_n3096_;
  assign new_n3121_ = new_n7894_ & new_n7890_;
  assign new_n3122_ = new_n7896_ | new_n7892_;
  assign new_n3123_ = new_n7893_ & new_n7889_;
  assign new_n3124_ = new_n7895_ | new_n7891_;
  assign new_n3125_ = new_n3124_ & new_n3122_;
  assign new_n3126_ = new_n3123_ | new_n3121_;
  assign new_n3127_ = new_n7581_ & new_n7573_;
  assign new_n3128_ = new_n7583_ | new_n7575_;
  assign new_n3129_ = new_n7897_ & new_n7898_;
  assign new_n3130_ = new_n3127_ | new_n3125_;
  assign new_n3131_ = new_n7899_ & new_n7898_;
  assign new_n3132_ = new_n7899_ & new_n7897_;
  assign new_n3133_ = new_n3132_ | new_n3131_;
  assign new_n3134_ = new_n6999_ & new_n7903_;
  assign new_n3135_ = new_n7005_ | new_n7918_;
  assign new_n3136_ = new_n7931_ & new_n7530_;
  assign new_n3137_ = new_n7932_ | new_n7532_;
  assign new_n3138_ = new_n7931_ & new_n7529_;
  assign new_n3139_ = new_n7932_ | new_n7531_;
  assign new_n3140_ = new_n3139_ & new_n3137_;
  assign new_n3141_ = new_n3138_ | new_n3136_;
  assign new_n3142_ = new_n7501_ & new_n6887_;
  assign new_n3143_ = new_n7503_ | new_n6893_;
  assign new_n3144_ = new_n3142_ | new_n3140_;
  assign new_n3145_ = new_n7934_ & new_n7383_;
  assign new_n3146_ = new_n7935_ | new_n7385_;
  assign new_n3147_ = new_n7934_ & new_n7382_;
  assign new_n3148_ = new_n7935_ | new_n7384_;
  assign new_n3149_ = new_n3148_ & new_n3146_;
  assign new_n3150_ = new_n3147_ | new_n3145_;
  assign new_n3151_ = new_n7355_ & new_n6812_;
  assign new_n3152_ = new_n7356_ | new_n6822_;
  assign new_n3153_ = new_n3151_ | new_n3149_;
  assign new_n3154_ = new_n7937_ & new_n7234_;
  assign new_n3155_ = new_n7938_ | new_n7236_;
  assign new_n3156_ = new_n7937_ & new_n7233_;
  assign new_n3157_ = new_n7938_ | new_n7235_;
  assign new_n3158_ = new_n3157_ & new_n3155_;
  assign new_n3159_ = new_n3156_ | new_n3154_;
  assign new_n3160_ = new_n7206_ & new_n6770_;
  assign new_n3161_ = new_n7207_ | new_n6784_;
  assign new_n3162_ = new_n3160_ | new_n3158_;
  assign new_n3163_ = new_n7939_ & new_n7940_;
  assign new_n3164_ = new_n6860_ & new_n7942_;
  assign new_n3165_ = new_n6869_ | new_n7945_;
  assign new_n3166_ = new_n7946_ & new_n7947_;
  assign new_n3167_ = new_n7948_ | new_n7949_;
  assign new_n3168_ = new_n7951_ & new_n7947_;
  assign new_n3169_ = new_n7953_ | new_n7949_;
  assign new_n3170_ = new_n7951_ & new_n7946_;
  assign new_n3171_ = new_n7953_ | new_n7948_;
  assign new_n3172_ = new_n3171_ & new_n3169_;
  assign new_n3173_ = new_n3170_ | new_n3168_;
  assign new_n3174_ = new_n6862_ & new_n7955_;
  assign new_n3175_ = new_n6871_ | new_n7958_;
  assign new_n3176_ = new_n7959_ & new_n7960_;
  assign new_n3177_ = new_n7961_ | new_n7962_;
  assign new_n3178_ = new_n7964_ & new_n7950_;
  assign new_n3179_ = new_n7966_ | new_n7952_;
  assign new_n3180_ = new_n7967_ & new_n7968_;
  assign new_n3181_ = new_n7969_ | new_n7970_;
  assign new_n3182_ = new_n7972_ & new_n7968_;
  assign new_n3183_ = new_n7974_ | new_n7970_;
  assign new_n3184_ = new_n7972_ & new_n7967_;
  assign new_n3185_ = new_n7974_ | new_n7969_;
  assign new_n3186_ = new_n3185_ & new_n3183_;
  assign new_n3187_ = new_n3184_ | new_n3182_;
  assign new_n3188_ = new_n6943_ & new_n7955_;
  assign new_n3189_ = new_n6956_ | new_n7958_;
  assign new_n3190_ = new_n7975_ & new_n7976_;
  assign new_n3191_ = new_n7977_ | new_n7978_;
  assign new_n3192_ = new_n7980_ & new_n7976_;
  assign new_n3193_ = new_n7982_ | new_n7978_;
  assign new_n3194_ = new_n7980_ & new_n7975_;
  assign new_n3195_ = new_n7982_ | new_n7977_;
  assign new_n3196_ = new_n3195_ & new_n3193_;
  assign new_n3197_ = new_n3194_ | new_n3192_;
  assign new_n3198_ = new_n7964_ & new_n7960_;
  assign new_n3199_ = new_n7966_ | new_n7962_;
  assign new_n3200_ = new_n7963_ & new_n7959_;
  assign new_n3201_ = new_n7965_ | new_n7961_;
  assign new_n3202_ = new_n3201_ & new_n3199_;
  assign new_n3203_ = new_n3200_ | new_n3198_;
  assign new_n3204_ = new_n1516_ & new_n1508_;
  assign new_n3205_ = new_n1515_ | new_n1507_;
  assign new_n3206_ = new_n6862_ & new_n7984_;
  assign new_n3207_ = new_n6871_ | new_n7987_;
  assign new_n3208_ = new_n7989_ & new_n7990_;
  assign new_n3209_ = new_n7991_ | new_n7992_;
  assign new_n3210_ = new_n7994_ & new_n1451_;
  assign new_n3211_ = new_n7996_ | new_n1452_;
  assign new_n3212_ = new_n7997_ & new_n7998_;
  assign new_n3213_ = new_n7999_ | new_n8000_;
  assign new_n3214_ = new_n8002_ & new_n7998_;
  assign new_n3215_ = new_n8004_ | new_n8000_;
  assign new_n3216_ = new_n8002_ & new_n7997_;
  assign new_n3217_ = new_n8004_ | new_n7999_;
  assign new_n3218_ = new_n3217_ & new_n3215_;
  assign new_n3219_ = new_n3216_ | new_n3214_;
  assign new_n3220_ = new_n6945_ & new_n7984_;
  assign new_n3221_ = new_n6958_ | new_n7987_;
  assign new_n3222_ = new_n8005_ & new_n8006_;
  assign new_n3223_ = new_n8007_ | new_n8008_;
  assign new_n3224_ = new_n8010_ & new_n8001_;
  assign new_n3225_ = new_n8012_ | new_n8003_;
  assign new_n3226_ = new_n8013_ & new_n8014_;
  assign new_n3227_ = new_n8015_ | new_n8016_;
  assign new_n3228_ = new_n8018_ & new_n8014_;
  assign new_n3229_ = new_n8020_ | new_n8016_;
  assign new_n3230_ = new_n8018_ & new_n8013_;
  assign new_n3231_ = new_n8020_ | new_n8015_;
  assign new_n3232_ = new_n3231_ & new_n3229_;
  assign new_n3233_ = new_n3230_ | new_n3228_;
  assign new_n3234_ = new_n7985_ & new_n7020_;
  assign new_n3235_ = new_n7988_ | new_n7035_;
  assign new_n3236_ = new_n8021_ & new_n8022_;
  assign new_n3237_ = new_n8023_ | new_n8024_;
  assign new_n3238_ = new_n8026_ & new_n8022_;
  assign new_n3239_ = new_n8028_ | new_n8024_;
  assign new_n3240_ = new_n8026_ & new_n8021_;
  assign new_n3241_ = new_n8028_ | new_n8023_;
  assign new_n3242_ = new_n3241_ & new_n3239_;
  assign new_n3243_ = new_n3240_ | new_n3238_;
  assign new_n3244_ = new_n8010_ & new_n8006_;
  assign new_n3245_ = new_n8012_ | new_n8008_;
  assign new_n3246_ = new_n8009_ & new_n8005_;
  assign new_n3247_ = new_n8011_ | new_n8007_;
  assign new_n3248_ = new_n3247_ & new_n3245_;
  assign new_n3249_ = new_n3246_ | new_n3244_;
  assign new_n3250_ = new_n7994_ & new_n7990_;
  assign new_n3251_ = new_n7996_ | new_n7992_;
  assign new_n3252_ = new_n7993_ & new_n7989_;
  assign new_n3253_ = new_n7995_ | new_n7991_;
  assign new_n3254_ = new_n3253_ & new_n3251_;
  assign new_n3255_ = new_n3252_ | new_n3250_;
  assign new_n3256_ = new_n8030_ & new_n1321_;
  assign new_n3257_ = new_n8032_ | new_n1322_;
  assign new_n3258_ = new_n8033_ & new_n8034_;
  assign new_n3259_ = new_n8035_ | new_n8036_;
  assign new_n3260_ = new_n8038_ & new_n8034_;
  assign new_n3261_ = new_n8040_ | new_n8036_;
  assign new_n3262_ = new_n8038_ & new_n8033_;
  assign new_n3263_ = new_n8040_ | new_n8035_;
  assign new_n3264_ = new_n3263_ & new_n3261_;
  assign new_n3265_ = new_n3262_ | new_n3260_;
  assign new_n3266_ = new_n6945_ & new_n8042_;
  assign new_n3267_ = new_n6958_ | new_n8045_;
  assign new_n3268_ = new_n8046_ & new_n8047_;
  assign new_n3269_ = new_n8048_ | new_n8049_;
  assign new_n3270_ = new_n8051_ & new_n8037_;
  assign new_n3271_ = new_n8053_ | new_n8039_;
  assign new_n3272_ = new_n8054_ & new_n8055_;
  assign new_n3273_ = new_n8056_ | new_n8057_;
  assign new_n3274_ = new_n8059_ & new_n8055_;
  assign new_n3275_ = new_n8061_ | new_n8057_;
  assign new_n3276_ = new_n8059_ & new_n8054_;
  assign new_n3277_ = new_n8061_ | new_n8056_;
  assign new_n3278_ = new_n3277_ & new_n3275_;
  assign new_n3279_ = new_n3276_ | new_n3274_;
  assign new_n3280_ = new_n8042_ & new_n7020_;
  assign new_n3281_ = new_n8045_ | new_n7035_;
  assign new_n3282_ = new_n8062_ & new_n8063_;
  assign new_n3283_ = new_n8064_ | new_n8065_;
  assign new_n3284_ = new_n8067_ & new_n8058_;
  assign new_n3285_ = new_n8069_ | new_n8060_;
  assign new_n3286_ = new_n8070_ & new_n8071_;
  assign new_n3287_ = new_n8072_ | new_n8073_;
  assign new_n3288_ = new_n8030_ & new_n1475_;
  assign new_n3289_ = new_n8032_ | new_n1476_;
  assign new_n3290_ = new_n8029_ & new_n1404_;
  assign new_n3291_ = new_n8031_ | new_n1403_;
  assign new_n3292_ = new_n3291_ & new_n3289_;
  assign new_n3293_ = new_n3290_ | new_n3288_;
  assign new_n3294_ = new_n1388_ & new_n1301_;
  assign new_n3295_ = new_n1387_ | new_n1302_;
  assign new_n3296_ = new_n8074_ & new_n8075_;
  assign new_n3297_ = new_n8076_ | new_n8077_;
  assign new_n3298_ = new_n8079_ & new_n8075_;
  assign new_n3299_ = new_n8081_ | new_n8077_;
  assign new_n3300_ = new_n8079_ & new_n8074_;
  assign new_n3301_ = new_n8081_ | new_n8076_;
  assign new_n3302_ = new_n3301_ & new_n3299_;
  assign new_n3303_ = new_n3300_ | new_n3298_;
  assign new_n3304_ = new_n6946_ & new_n8083_;
  assign new_n3305_ = new_n6959_ | new_n8086_;
  assign new_n3306_ = new_n8087_ & new_n8088_;
  assign new_n3307_ = new_n8089_ | new_n8090_;
  assign new_n3308_ = new_n8092_ & new_n8088_;
  assign new_n3309_ = new_n8094_ | new_n8090_;
  assign new_n3310_ = new_n8092_ & new_n8087_;
  assign new_n3311_ = new_n8094_ | new_n8089_;
  assign new_n3312_ = new_n3311_ & new_n3309_;
  assign new_n3313_ = new_n3310_ | new_n3308_;
  assign new_n3314_ = new_n8095_ & new_n8096_;
  assign new_n3315_ = new_n8097_ | new_n8098_;
  assign new_n3316_ = new_n8100_ & new_n8095_;
  assign new_n3317_ = new_n8102_ | new_n8097_;
  assign new_n3318_ = new_n8100_ & new_n8096_;
  assign new_n3319_ = new_n8102_ | new_n8098_;
  assign new_n3320_ = new_n3319_ & new_n3317_;
  assign new_n3321_ = new_n3318_ | new_n3316_;
  assign new_n3322_ = new_n6946_ & new_n8104_;
  assign new_n3323_ = new_n6959_ | new_n8107_;
  assign new_n3324_ = new_n8108_ & new_n8109_;
  assign new_n3325_ = new_n8110_ | new_n8111_;
  assign new_n3326_ = new_n8113_ & new_n8099_;
  assign new_n3327_ = new_n8115_ | new_n8101_;
  assign new_n3328_ = new_n8116_ & new_n8117_;
  assign new_n3329_ = new_n8118_ | new_n8119_;
  assign new_n3330_ = new_n8121_ & new_n8117_;
  assign new_n3331_ = new_n8123_ | new_n8119_;
  assign new_n3332_ = new_n8121_ & new_n8116_;
  assign new_n3333_ = new_n8123_ | new_n8118_;
  assign new_n3334_ = new_n3333_ & new_n3331_;
  assign new_n3335_ = new_n3332_ | new_n3330_;
  assign new_n3336_ = new_n8104_ & new_n7022_;
  assign new_n3337_ = new_n8107_ | new_n7037_;
  assign new_n3338_ = new_n8124_ & new_n8125_;
  assign new_n3339_ = new_n8126_ | new_n8127_;
  assign new_n3340_ = new_n8129_ & new_n8125_;
  assign new_n3341_ = new_n8131_ | new_n8127_;
  assign new_n3342_ = new_n8129_ & new_n8124_;
  assign new_n3343_ = new_n8131_ | new_n8126_;
  assign new_n3344_ = new_n3343_ & new_n3341_;
  assign new_n3345_ = new_n3342_ | new_n3340_;
  assign new_n3346_ = new_n8113_ & new_n8109_;
  assign new_n3347_ = new_n8115_ | new_n8111_;
  assign new_n3348_ = new_n8112_ & new_n8108_;
  assign new_n3349_ = new_n8114_ | new_n8110_;
  assign new_n3350_ = new_n3349_ & new_n3347_;
  assign new_n3351_ = new_n3348_ | new_n3346_;
  assign new_n3352_ = new_n1518_ & new_n1510_;
  assign new_n3353_ = new_n1517_ | new_n1509_;
  assign new_n3354_ = new_n6949_ & new_n8133_;
  assign new_n3355_ = new_n6962_ | new_n8136_;
  assign new_n3356_ = new_n8138_ & new_n8139_;
  assign new_n3357_ = new_n8140_ | new_n8141_;
  assign new_n3358_ = new_n8143_ & new_n1453_;
  assign new_n3359_ = new_n8145_ | new_n1454_;
  assign new_n3360_ = new_n8146_ & new_n8147_;
  assign new_n3361_ = new_n8148_ | new_n8149_;
  assign new_n3362_ = new_n8151_ & new_n8147_;
  assign new_n3363_ = new_n8153_ | new_n8149_;
  assign new_n3364_ = new_n8151_ & new_n8146_;
  assign new_n3365_ = new_n8153_ | new_n8148_;
  assign new_n3366_ = new_n3365_ & new_n3363_;
  assign new_n3367_ = new_n3364_ | new_n3362_;
  assign new_n3368_ = new_n8133_ & new_n7022_;
  assign new_n3369_ = new_n8136_ | new_n7037_;
  assign new_n3370_ = new_n8154_ & new_n8155_;
  assign new_n3371_ = new_n8156_ | new_n8157_;
  assign new_n3372_ = new_n8159_ & new_n8150_;
  assign new_n3373_ = new_n8161_ | new_n8152_;
  assign new_n3374_ = new_n8162_ & new_n8163_;
  assign new_n3375_ = new_n8164_ | new_n8165_;
  assign new_n3376_ = new_n8167_ & new_n8163_;
  assign new_n3377_ = new_n8169_ | new_n8165_;
  assign new_n3378_ = new_n8167_ & new_n8162_;
  assign new_n3379_ = new_n8169_ | new_n8164_;
  assign new_n3380_ = new_n3379_ & new_n3377_;
  assign new_n3381_ = new_n3378_ | new_n3376_;
  assign new_n3382_ = new_n8134_ & new_n7594_;
  assign new_n3383_ = new_n8137_ | new_n7607_;
  assign new_n3384_ = new_n8170_ & new_n8171_;
  assign new_n3385_ = new_n8172_ | new_n8173_;
  assign new_n3386_ = new_n8175_ & new_n8171_;
  assign new_n3387_ = new_n8177_ | new_n8173_;
  assign new_n3388_ = new_n8175_ & new_n8170_;
  assign new_n3389_ = new_n8177_ | new_n8172_;
  assign new_n3390_ = new_n3389_ & new_n3387_;
  assign new_n3391_ = new_n3388_ | new_n3386_;
  assign new_n3392_ = new_n8159_ & new_n8155_;
  assign new_n3393_ = new_n8161_ | new_n8157_;
  assign new_n3394_ = new_n8158_ & new_n8154_;
  assign new_n3395_ = new_n8160_ | new_n8156_;
  assign new_n3396_ = new_n3395_ & new_n3393_;
  assign new_n3397_ = new_n3394_ | new_n3392_;
  assign new_n3398_ = new_n8143_ & new_n8139_;
  assign new_n3399_ = new_n8145_ | new_n8141_;
  assign new_n3400_ = new_n8142_ & new_n8138_;
  assign new_n3401_ = new_n8144_ | new_n8140_;
  assign new_n3402_ = new_n3401_ & new_n3399_;
  assign new_n3403_ = new_n3400_ | new_n3398_;
  assign new_n3404_ = new_n8179_ & new_n1325_;
  assign new_n3405_ = new_n8181_ | new_n1326_;
  assign new_n3406_ = new_n8182_ & new_n8183_;
  assign new_n3407_ = new_n8184_ | new_n8185_;
  assign new_n3408_ = new_n8187_ & new_n8183_;
  assign new_n3409_ = new_n8189_ | new_n8185_;
  assign new_n3410_ = new_n8187_ & new_n8182_;
  assign new_n3411_ = new_n8189_ | new_n8184_;
  assign new_n3412_ = new_n3411_ & new_n3409_;
  assign new_n3413_ = new_n3410_ | new_n3408_;
  assign new_n3414_ = new_n8191_ & new_n7023_;
  assign new_n3415_ = new_n8194_ | new_n7038_;
  assign new_n3416_ = new_n8195_ & new_n8196_;
  assign new_n3417_ = new_n8197_ | new_n8198_;
  assign new_n3418_ = new_n8200_ & new_n8186_;
  assign new_n3419_ = new_n8202_ | new_n8188_;
  assign new_n3420_ = new_n8203_ & new_n8204_;
  assign new_n3421_ = new_n8205_ | new_n8206_;
  assign new_n3422_ = new_n8208_ & new_n8204_;
  assign new_n3423_ = new_n8210_ | new_n8206_;
  assign new_n3424_ = new_n8208_ & new_n8203_;
  assign new_n3425_ = new_n8210_ | new_n8205_;
  assign new_n3426_ = new_n3425_ & new_n3423_;
  assign new_n3427_ = new_n3424_ | new_n3422_;
  assign new_n3428_ = new_n8191_ & new_n7595_;
  assign new_n3429_ = new_n8194_ | new_n7608_;
  assign new_n3430_ = new_n8211_ & new_n8212_;
  assign new_n3431_ = new_n8213_ | new_n8214_;
  assign new_n3432_ = new_n8216_ & new_n8207_;
  assign new_n3433_ = new_n8218_ | new_n8209_;
  assign new_n3434_ = new_n8219_ & new_n8220_;
  assign new_n3435_ = new_n8221_ | new_n8222_;
  assign new_n3436_ = new_n8179_ & new_n1479_;
  assign new_n3437_ = new_n8181_ | new_n1480_;
  assign new_n3438_ = new_n8178_ & new_n1406_;
  assign new_n3439_ = new_n8180_ | new_n1405_;
  assign new_n3440_ = new_n3439_ & new_n3437_;
  assign new_n3441_ = new_n3438_ | new_n3436_;
  assign new_n3442_ = new_n8223_ & new_n8224_;
  assign new_n3443_ = new_n8225_ | new_n8226_;
  assign new_n3444_ = new_n8228_ & new_n1393_;
  assign new_n3445_ = new_n8230_ | new_n1394_;
  assign new_n3446_ = new_n8231_ & new_n8232_;
  assign new_n3447_ = new_n8233_ | new_n8234_;
  assign new_n3448_ = new_n8236_ & new_n8232_;
  assign new_n3449_ = new_n8238_ | new_n8234_;
  assign new_n3450_ = new_n8236_ & new_n8231_;
  assign new_n3451_ = new_n8238_ | new_n8233_;
  assign new_n3452_ = new_n3451_ & new_n3449_;
  assign new_n3453_ = new_n3450_ | new_n3448_;
  assign new_n3454_ = new_n8240_ & new_n7023_;
  assign new_n3455_ = new_n8243_ | new_n7038_;
  assign new_n3456_ = new_n8244_ & new_n8245_;
  assign new_n3457_ = new_n8246_ | new_n8247_;
  assign new_n3458_ = new_n8249_ & new_n8245_;
  assign new_n3459_ = new_n8251_ | new_n8247_;
  assign new_n3460_ = new_n8249_ & new_n8244_;
  assign new_n3461_ = new_n8251_ | new_n8246_;
  assign new_n3462_ = new_n3461_ & new_n3459_;
  assign new_n3463_ = new_n3460_ | new_n3458_;
  assign new_n3464_ = new_n8228_ & new_n8223_;
  assign new_n3465_ = new_n8230_ | new_n8225_;
  assign new_n3466_ = new_n8227_ & new_n8224_;
  assign new_n3467_ = new_n8229_ | new_n8226_;
  assign new_n3468_ = new_n3467_ & new_n3465_;
  assign new_n3469_ = new_n3466_ | new_n3464_;
  assign new_n3470_ = new_n1520_ & new_n1514_;
  assign new_n3471_ = new_n1519_ | new_n1513_;
  assign new_n3472_ = new_n6949_ & new_n8254_;
  assign new_n3473_ = new_n6962_ | new_n8257_;
  assign new_n3474_ = new_n8259_ & new_n8260_;
  assign new_n3475_ = new_n8261_ | new_n8262_;
  assign new_n3476_ = new_n8264_ & new_n1457_;
  assign new_n3477_ = new_n8266_ | new_n1458_;
  assign new_n3478_ = new_n8267_ & new_n8268_;
  assign new_n3479_ = new_n8269_ | new_n8270_;
  assign new_n3480_ = new_n8272_ & new_n8268_;
  assign new_n3481_ = new_n8274_ | new_n8270_;
  assign new_n3482_ = new_n8272_ & new_n8267_;
  assign new_n3483_ = new_n8274_ | new_n8269_;
  assign new_n3484_ = new_n3483_ & new_n3481_;
  assign new_n3485_ = new_n3482_ | new_n3480_;
  assign new_n3486_ = new_n8254_ & new_n7026_;
  assign new_n3487_ = new_n8257_ | new_n7041_;
  assign new_n3488_ = new_n8275_ & new_n8276_;
  assign new_n3489_ = new_n8277_ | new_n8278_;
  assign new_n3490_ = new_n8280_ & new_n8271_;
  assign new_n3491_ = new_n8282_ | new_n8273_;
  assign new_n3492_ = new_n8283_ & new_n8284_;
  assign new_n3493_ = new_n8285_ | new_n8286_;
  assign new_n3494_ = new_n8288_ & new_n8284_;
  assign new_n3495_ = new_n8290_ | new_n8286_;
  assign new_n3496_ = new_n8288_ & new_n8283_;
  assign new_n3497_ = new_n8290_ | new_n8285_;
  assign new_n3498_ = new_n3497_ & new_n3495_;
  assign new_n3499_ = new_n3496_ | new_n3494_;
  assign new_n3500_ = new_n8253_ & new_n7595_;
  assign new_n3501_ = new_n8258_ | new_n7608_;
  assign new_n3502_ = new_n8291_ & new_n8292_;
  assign new_n3503_ = new_n8293_ | new_n8294_;
  assign new_n3504_ = new_n8296_ & new_n8292_;
  assign new_n3505_ = new_n8298_ | new_n8294_;
  assign new_n3506_ = new_n8296_ & new_n8291_;
  assign new_n3507_ = new_n8298_ | new_n8293_;
  assign new_n3508_ = new_n3507_ & new_n3505_;
  assign new_n3509_ = new_n3506_ | new_n3504_;
  assign new_n3510_ = new_n8280_ & new_n8276_;
  assign new_n3511_ = new_n8282_ | new_n8278_;
  assign new_n3512_ = new_n8279_ & new_n8275_;
  assign new_n3513_ = new_n8281_ | new_n8277_;
  assign new_n3514_ = new_n3513_ & new_n3511_;
  assign new_n3515_ = new_n3512_ | new_n3510_;
  assign new_n3516_ = new_n8264_ & new_n8260_;
  assign new_n3517_ = new_n8266_ | new_n8262_;
  assign new_n3518_ = new_n8263_ & new_n8259_;
  assign new_n3519_ = new_n8265_ | new_n8261_;
  assign new_n3520_ = new_n3519_ & new_n3517_;
  assign new_n3521_ = new_n3518_ | new_n3516_;
  assign new_n3522_ = new_n8300_ & new_n1472_;
  assign new_n3523_ = new_n8302_ | new_n1471_;
  assign new_n3524_ = new_n8300_ & new_n1420_;
  assign new_n3525_ = new_n8302_ | new_n1419_;
  assign new_n3526_ = new_n3525_ & new_n3523_;
  assign new_n3527_ = new_n3524_ | new_n3522_;
  assign new_n3528_ = new_n6950_ & new_n8305_;
  assign new_n3529_ = new_n6963_ | new_n8309_;
  assign new_n3530_ = new_n8311_ & new_n8312_;
  assign new_n3531_ = new_n8313_ | new_n8314_;
  assign new_n3532_ = new_n8316_ & new_n8299_;
  assign new_n3533_ = new_n8318_ | new_n8301_;
  assign new_n3534_ = new_n8319_ & new_n8320_;
  assign new_n3535_ = new_n8321_ | new_n8322_;
  assign new_n3536_ = new_n8324_ & new_n8320_;
  assign new_n3537_ = new_n8326_ | new_n8322_;
  assign new_n3538_ = new_n8324_ & new_n8319_;
  assign new_n3539_ = new_n8326_ | new_n8321_;
  assign new_n3540_ = new_n3539_ & new_n3537_;
  assign new_n3541_ = new_n3538_ | new_n3536_;
  assign new_n3542_ = new_n8305_ & new_n7026_;
  assign new_n3543_ = new_n8309_ | new_n7041_;
  assign new_n3544_ = new_n8327_ & new_n8328_;
  assign new_n3545_ = new_n8329_ | new_n8330_;
  assign new_n3546_ = new_n8332_ & new_n8323_;
  assign new_n3547_ = new_n8334_ | new_n8325_;
  assign new_n3548_ = new_n8335_ & new_n8336_;
  assign new_n3549_ = new_n8337_ | new_n8338_;
  assign new_n3550_ = new_n8340_ & new_n8336_;
  assign new_n3551_ = new_n8342_ | new_n8338_;
  assign new_n3552_ = new_n8340_ & new_n8335_;
  assign new_n3553_ = new_n8342_ | new_n8337_;
  assign new_n3554_ = new_n3553_ & new_n3551_;
  assign new_n3555_ = new_n3552_ | new_n3550_;
  assign new_n3556_ = new_n8304_ & new_n7597_;
  assign new_n3557_ = new_n8308_ | new_n7610_;
  assign new_n3558_ = new_n8343_ & new_n8344_;
  assign new_n3559_ = new_n8345_ | new_n8346_;
  assign new_n3560_ = new_n8348_ & new_n8339_;
  assign new_n3561_ = new_n8350_ | new_n8341_;
  assign new_n3562_ = new_n8351_ & new_n8352_;
  assign new_n3563_ = new_n8353_ | new_n8354_;
  assign new_n3564_ = new_n8356_ & new_n8352_;
  assign new_n3565_ = new_n8358_ | new_n8354_;
  assign new_n3566_ = new_n8356_ & new_n8351_;
  assign new_n3567_ = new_n8358_ | new_n8353_;
  assign new_n3568_ = new_n3567_ & new_n3565_;
  assign new_n3569_ = new_n3566_ | new_n3564_;
  assign new_n3570_ = new_n8306_ & new_n8362_;
  assign new_n3571_ = new_n8310_ | new_n8371_;
  assign new_n3572_ = new_n8377_ & new_n8378_;
  assign new_n3573_ = new_n8379_ | new_n8380_;
  assign new_n3574_ = new_n8382_ & new_n8378_;
  assign new_n3575_ = new_n8384_ | new_n8380_;
  assign new_n3576_ = new_n8382_ & new_n8377_;
  assign new_n3577_ = new_n8384_ | new_n8379_;
  assign new_n3578_ = new_n3577_ & new_n3575_;
  assign new_n3579_ = new_n3576_ | new_n3574_;
  assign new_n3580_ = new_n8348_ & new_n8344_;
  assign new_n3581_ = new_n8350_ | new_n8346_;
  assign new_n3582_ = new_n8347_ & new_n8343_;
  assign new_n3583_ = new_n8349_ | new_n8345_;
  assign new_n3584_ = new_n3583_ & new_n3581_;
  assign new_n3585_ = new_n3582_ | new_n3580_;
  assign new_n3586_ = new_n8332_ & new_n8328_;
  assign new_n3587_ = new_n8334_ | new_n8330_;
  assign new_n3588_ = new_n8331_ & new_n8327_;
  assign new_n3589_ = new_n8333_ | new_n8329_;
  assign new_n3590_ = new_n3589_ & new_n3587_;
  assign new_n3591_ = new_n3588_ | new_n3586_;
  assign new_n3592_ = new_n8316_ & new_n8312_;
  assign new_n3593_ = new_n8318_ | new_n8314_;
  assign new_n3594_ = new_n8315_ & new_n8311_;
  assign new_n3595_ = new_n8317_ | new_n8313_;
  assign new_n3596_ = new_n3595_ & new_n3593_;
  assign new_n3597_ = new_n3594_ | new_n3592_;
  assign new_n3598_ = new_n8385_ & new_n8386_;
  assign new_n3599_ = new_n8387_ | new_n8388_;
  assign new_n3600_ = new_n8390_ & new_n8385_;
  assign new_n3601_ = new_n8392_ | new_n8387_;
  assign new_n3602_ = new_n8390_ & new_n8386_;
  assign new_n3603_ = new_n8392_ | new_n8388_;
  assign new_n3604_ = new_n3603_ & new_n3601_;
  assign new_n3605_ = new_n3602_ | new_n3600_;
  assign new_n3606_ = new_n6950_ & new_n8395_;
  assign new_n3607_ = new_n6963_ | new_n8400_;
  assign new_n3608_ = new_n8402_ & new_n8403_;
  assign new_n3609_ = new_n8404_ | new_n8405_;
  assign new_n3610_ = new_n8407_ & new_n8389_;
  assign new_n3611_ = new_n8409_ | new_n8391_;
  assign new_n3612_ = new_n8410_ & new_n8411_;
  assign new_n3613_ = new_n8412_ | new_n8413_;
  assign new_n3614_ = new_n8415_ & new_n8411_;
  assign new_n3615_ = new_n8417_ | new_n8413_;
  assign new_n3616_ = new_n8415_ & new_n8410_;
  assign new_n3617_ = new_n8417_ | new_n8412_;
  assign new_n3618_ = new_n3617_ & new_n3615_;
  assign new_n3619_ = new_n3616_ | new_n3614_;
  assign new_n3620_ = new_n8395_ & new_n7027_;
  assign new_n3621_ = new_n8400_ | new_n7042_;
  assign new_n3622_ = new_n8418_ & new_n8419_;
  assign new_n3623_ = new_n8420_ | new_n8421_;
  assign new_n3624_ = new_n8423_ & new_n8414_;
  assign new_n3625_ = new_n8425_ | new_n8416_;
  assign new_n3626_ = new_n8426_ & new_n8427_;
  assign new_n3627_ = new_n8428_ | new_n8429_;
  assign new_n3628_ = new_n8431_ & new_n8427_;
  assign new_n3629_ = new_n8433_ | new_n8429_;
  assign new_n3630_ = new_n8431_ & new_n8426_;
  assign new_n3631_ = new_n8433_ | new_n8428_;
  assign new_n3632_ = new_n3631_ & new_n3629_;
  assign new_n3633_ = new_n3630_ | new_n3628_;
  assign new_n3634_ = new_n8396_ & new_n7597_;
  assign new_n3635_ = new_n8399_ | new_n7610_;
  assign new_n3636_ = new_n8434_ & new_n8435_;
  assign new_n3637_ = new_n8436_ | new_n8437_;
  assign new_n3638_ = new_n8439_ & new_n8430_;
  assign new_n3639_ = new_n8441_ | new_n8432_;
  assign new_n3640_ = new_n8442_ & new_n8443_;
  assign new_n3641_ = new_n8444_ | new_n8445_;
  assign new_n3642_ = new_n8447_ & new_n8443_;
  assign new_n3643_ = new_n8449_ | new_n8445_;
  assign new_n3644_ = new_n8447_ & new_n8442_;
  assign new_n3645_ = new_n8449_ | new_n8444_;
  assign new_n3646_ = new_n3645_ & new_n3643_;
  assign new_n3647_ = new_n3644_ | new_n3642_;
  assign new_n3648_ = new_n8396_ & new_n8362_;
  assign new_n3649_ = new_n8401_ | new_n8371_;
  assign new_n3650_ = new_n8450_ & new_n8451_;
  assign new_n3651_ = new_n8452_ | new_n8453_;
  assign new_n3652_ = new_n8455_ & new_n8446_;
  assign new_n3653_ = new_n8457_ | new_n8448_;
  assign new_n3654_ = new_n8458_ & new_n8459_;
  assign new_n3655_ = new_n8460_ | new_n8461_;
  assign new_n3656_ = new_n8462_ & new_n8463_;
  assign new_n3657_ = new_n8464_ | new_n8465_;
  assign new_n3658_ = new_n8467_ & new_n8462_;
  assign new_n3659_ = new_n8469_ | new_n8464_;
  assign new_n3660_ = new_n8467_ & new_n8463_;
  assign new_n3661_ = new_n8469_ | new_n8465_;
  assign new_n3662_ = new_n3661_ & new_n3659_;
  assign new_n3663_ = new_n3660_ | new_n3658_;
  assign new_n3664_ = new_n7716_ & new_n1537_;
  assign new_n3665_ = new_n7718_ | new_n1538_;
  assign new_n3666_ = new_n8470_ & new_n8471_;
  assign new_n3667_ = new_n8472_ | new_n8473_;
  assign new_n3668_ = new_n8475_ & new_n8471_;
  assign new_n3669_ = new_n8477_ | new_n8473_;
  assign new_n3670_ = new_n8475_ & new_n8470_;
  assign new_n3671_ = new_n8477_ | new_n8472_;
  assign new_n3672_ = new_n3671_ & new_n3669_;
  assign new_n3673_ = new_n3670_ | new_n3668_;
  assign new_n3674_ = new_n7085_ & new_n7704_;
  assign new_n3675_ = new_n7093_ | new_n7710_;
  assign new_n3676_ = new_n8478_ & new_n8479_;
  assign new_n3677_ = new_n8480_ | new_n8481_;
  assign new_n3678_ = new_n8483_ & new_n8479_;
  assign new_n3679_ = new_n8485_ | new_n8481_;
  assign new_n3680_ = new_n8483_ & new_n8478_;
  assign new_n3681_ = new_n8485_ | new_n8480_;
  assign new_n3682_ = new_n3681_ & new_n3679_;
  assign new_n3683_ = new_n3680_ | new_n3678_;
  assign new_n3684_ = new_n7732_ & new_n7724_;
  assign new_n3685_ = new_n7734_ | new_n7726_;
  assign new_n3686_ = new_n8486_ & new_n8487_;
  assign new_n3687_ = new_n8488_ | new_n8489_;
  assign new_n3688_ = new_n8491_ & new_n8487_;
  assign new_n3689_ = new_n8493_ | new_n8489_;
  assign new_n3690_ = new_n8491_ & new_n8486_;
  assign new_n3691_ = new_n8493_ | new_n8488_;
  assign new_n3692_ = new_n3691_ & new_n3689_;
  assign new_n3693_ = new_n3690_ | new_n3688_;
  assign new_n3694_ = new_n7673_ & new_n7106_;
  assign new_n3695_ = new_n7688_ | new_n7109_;
  assign new_n3696_ = new_n8494_ & new_n8495_;
  assign new_n3697_ = new_n8496_ | new_n8497_;
  assign new_n3698_ = new_n8499_ & new_n8495_;
  assign new_n3699_ = new_n8501_ | new_n8497_;
  assign new_n3700_ = new_n8499_ & new_n8494_;
  assign new_n3701_ = new_n8501_ | new_n8496_;
  assign new_n3702_ = new_n3701_ & new_n3699_;
  assign new_n3703_ = new_n3700_ | new_n3698_;
  assign new_n3704_ = new_n2907_ & new_n7741_;
  assign new_n3705_ = new_n8502_ | new_n7743_;
  assign new_n3706_ = new_n8503_ & new_n8504_;
  assign new_n3707_ = new_n8505_ | new_n8506_;
  assign new_n3708_ = new_n8508_ & new_n8504_;
  assign new_n3709_ = new_n8510_ | new_n8506_;
  assign new_n3710_ = new_n8508_ & new_n8503_;
  assign new_n3711_ = new_n8510_ | new_n8505_;
  assign new_n3712_ = new_n3711_ & new_n3709_;
  assign new_n3713_ = new_n3710_ | new_n3708_;
  assign new_n3714_ = new_n6867_ & new_n8363_;
  assign new_n3715_ = new_n6875_ | new_n8372_;
  assign new_n3716_ = new_n8511_ & new_n3135_;
  assign new_n3717_ = new_n3712_ | new_n8512_;
  assign new_n3718_ = new_n1524_ & new_n1505_;
  assign new_n3719_ = new_n1523_ | new_n1506_;
  assign new_n3720_ = new_n7617_ & new_n1323_;
  assign new_n3721_ = new_n7619_ | new_n1324_;
  assign new_n3722_ = new_n8513_ & new_n8514_;
  assign new_n3723_ = new_n8515_ | new_n8516_;
  assign new_n3724_ = new_n8518_ & new_n8514_;
  assign new_n3725_ = new_n8520_ | new_n8516_;
  assign new_n3726_ = new_n8518_ & new_n8513_;
  assign new_n3727_ = new_n8520_ | new_n8515_;
  assign new_n3728_ = new_n3727_ & new_n3725_;
  assign new_n3729_ = new_n3726_ | new_n3724_;
  assign new_n3730_ = new_n6951_ & new_n8523_;
  assign new_n3731_ = new_n6964_ | new_n8528_;
  assign new_n3732_ = new_n8530_ & new_n8531_;
  assign new_n3733_ = new_n8532_ | new_n8533_;
  assign new_n3734_ = new_n8535_ & new_n8531_;
  assign new_n3735_ = new_n8537_ | new_n8533_;
  assign new_n3736_ = new_n8535_ & new_n8530_;
  assign new_n3737_ = new_n8537_ | new_n8532_;
  assign new_n3738_ = new_n3737_ & new_n3735_;
  assign new_n3739_ = new_n3736_ | new_n3734_;
  assign new_n3740_ = new_n7641_ & new_n7625_;
  assign new_n3741_ = new_n7643_ | new_n7627_;
  assign new_n3742_ = new_n8538_ & new_n8539_;
  assign new_n3743_ = new_n8540_ | new_n8541_;
  assign new_n3744_ = new_n8543_ & new_n8539_;
  assign new_n3745_ = new_n8545_ | new_n8541_;
  assign new_n3746_ = new_n8543_ & new_n8538_;
  assign new_n3747_ = new_n8545_ | new_n8540_;
  assign new_n3748_ = new_n3747_ & new_n3745_;
  assign new_n3749_ = new_n3746_ | new_n3744_;
  assign new_n3750_ = new_n7631_ & new_n7027_;
  assign new_n3751_ = new_n7635_ | new_n7042_;
  assign new_n3752_ = new_n8546_ & new_n8547_;
  assign new_n3753_ = new_n8548_ | new_n8549_;
  assign new_n3754_ = new_n8551_ & new_n8547_;
  assign new_n3755_ = new_n8553_ | new_n8549_;
  assign new_n3756_ = new_n8551_ & new_n8546_;
  assign new_n3757_ = new_n8553_ | new_n8548_;
  assign new_n3758_ = new_n3757_ & new_n3755_;
  assign new_n3759_ = new_n3756_ | new_n3754_;
  assign new_n3760_ = new_n7657_ & new_n7649_;
  assign new_n3761_ = new_n7659_ | new_n7651_;
  assign new_n3762_ = new_n8554_ & new_n8555_;
  assign new_n3763_ = new_n8556_ | new_n8557_;
  assign new_n3764_ = new_n8559_ & new_n8555_;
  assign new_n3765_ = new_n8561_ | new_n8557_;
  assign new_n3766_ = new_n8559_ & new_n8554_;
  assign new_n3767_ = new_n8561_ | new_n8556_;
  assign new_n3768_ = new_n3767_ & new_n3765_;
  assign new_n3769_ = new_n3766_ | new_n3764_;
  assign new_n3770_ = new_n6970_ & new_n7598_;
  assign new_n3771_ = new_n6976_ | new_n7611_;
  assign new_n3772_ = new_n8562_ & new_n8563_;
  assign new_n3773_ = new_n8564_ | new_n8565_;
  assign new_n3774_ = new_n8567_ & new_n8563_;
  assign new_n3775_ = new_n8569_ | new_n8565_;
  assign new_n3776_ = new_n8567_ & new_n8562_;
  assign new_n3777_ = new_n8569_ | new_n8564_;
  assign new_n3778_ = new_n3777_ & new_n3775_;
  assign new_n3779_ = new_n3776_ | new_n3774_;
  assign new_n3780_ = new_n2863_ & new_n7666_;
  assign new_n3781_ = new_n8570_ | new_n7668_;
  assign new_n3782_ = new_n8571_ & new_n8572_;
  assign new_n3783_ = new_n8573_ | new_n8574_;
  assign new_n3784_ = new_n8576_ & new_n8572_;
  assign new_n3785_ = new_n8578_ | new_n8574_;
  assign new_n3786_ = new_n8576_ & new_n8571_;
  assign new_n3787_ = new_n8578_ | new_n8573_;
  assign new_n3788_ = new_n3787_ & new_n3785_;
  assign new_n3789_ = new_n3786_ | new_n3784_;
  assign new_n3790_ = new_n7448_ | new_n6893_;
  assign new_n3791_ = new_n7300_ | new_n6823_;
  assign new_n3792_ = new_n7151_ | new_n6784_;
  assign new_n3793_ = new_n8579_ | new_n3129_;
  assign new_n3794_ = new_n7230_ & new_n7226_;
  assign new_n3795_ = new_n7232_ | new_n7228_;
  assign new_n3796_ = new_n7229_ & new_n7225_;
  assign new_n3797_ = new_n7231_ | new_n7227_;
  assign new_n3798_ = new_n3797_ & new_n3795_;
  assign new_n3799_ = new_n3796_ | new_n3794_;
  assign new_n3800_ = new_n7761_ & new_n7753_;
  assign new_n3801_ = new_n7763_ | new_n7755_;
  assign new_n3802_ = new_n8580_ & new_n8581_;
  assign new_n3803_ = new_n8582_ | new_n8583_;
  assign new_n3804_ = new_n8585_ & new_n8581_;
  assign new_n3805_ = new_n8586_ | new_n8583_;
  assign new_n3806_ = new_n8585_ & new_n8580_;
  assign new_n3807_ = new_n8586_ | new_n8582_;
  assign new_n3808_ = new_n3807_ & new_n3805_;
  assign new_n3809_ = new_n3806_ | new_n3804_;
  assign new_n3810_ = new_n7247_ & new_n6770_;
  assign new_n3811_ = new_n7248_ | new_n6783_;
  assign new_n3812_ = new_n8587_ & new_n8588_;
  assign new_n3813_ = new_n8589_ | new_n8590_;
  assign new_n3814_ = new_n8592_ & new_n8588_;
  assign new_n3815_ = new_n8593_ | new_n8590_;
  assign new_n3816_ = new_n8592_ & new_n8587_;
  assign new_n3817_ = new_n8593_ | new_n8589_;
  assign new_n3818_ = new_n3817_ & new_n3815_;
  assign new_n3819_ = new_n3816_ | new_n3814_;
  assign new_n3820_ = new_n7777_ & new_n7769_;
  assign new_n3821_ = new_n7779_ | new_n7771_;
  assign new_n3822_ = new_n3820_ | new_n3818_;
  assign new_n3823_ = new_n7379_ & new_n7375_;
  assign new_n3824_ = new_n7381_ | new_n7377_;
  assign new_n3825_ = new_n7378_ & new_n7374_;
  assign new_n3826_ = new_n7380_ | new_n7376_;
  assign new_n3827_ = new_n3826_ & new_n3824_;
  assign new_n3828_ = new_n3825_ | new_n3823_;
  assign new_n3829_ = new_n7793_ & new_n7785_;
  assign new_n3830_ = new_n7795_ | new_n7787_;
  assign new_n3831_ = new_n8594_ & new_n8595_;
  assign new_n3832_ = new_n8596_ | new_n8597_;
  assign new_n3833_ = new_n8599_ & new_n8595_;
  assign new_n3834_ = new_n8600_ | new_n8597_;
  assign new_n3835_ = new_n8599_ & new_n8594_;
  assign new_n3836_ = new_n8600_ | new_n8596_;
  assign new_n3837_ = new_n3836_ & new_n3834_;
  assign new_n3838_ = new_n3835_ | new_n3833_;
  assign new_n3839_ = new_n7396_ & new_n6813_;
  assign new_n3840_ = new_n7397_ | new_n6823_;
  assign new_n3841_ = new_n8601_ & new_n8602_;
  assign new_n3842_ = new_n8603_ | new_n8604_;
  assign new_n3843_ = new_n8606_ & new_n8602_;
  assign new_n3844_ = new_n8607_ | new_n8604_;
  assign new_n3845_ = new_n8606_ & new_n8601_;
  assign new_n3846_ = new_n8607_ | new_n8603_;
  assign new_n3847_ = new_n3846_ & new_n3844_;
  assign new_n3848_ = new_n3845_ | new_n3843_;
  assign new_n3849_ = new_n7809_ & new_n7801_;
  assign new_n3850_ = new_n7811_ | new_n7803_;
  assign new_n3851_ = new_n3849_ | new_n3847_;
  assign new_n3852_ = new_n7526_ & new_n7522_;
  assign new_n3853_ = new_n7528_ | new_n7524_;
  assign new_n3854_ = new_n7525_ & new_n7521_;
  assign new_n3855_ = new_n7527_ | new_n7523_;
  assign new_n3856_ = new_n3855_ & new_n3853_;
  assign new_n3857_ = new_n3854_ | new_n3852_;
  assign new_n3858_ = new_n7845_ & new_n7837_;
  assign new_n3859_ = new_n7847_ | new_n7839_;
  assign new_n3860_ = new_n8608_ & new_n8609_;
  assign new_n3861_ = new_n8610_ | new_n8611_;
  assign new_n3862_ = new_n8613_ & new_n8609_;
  assign new_n3863_ = new_n8614_ | new_n8611_;
  assign new_n3864_ = new_n8613_ & new_n8608_;
  assign new_n3865_ = new_n8614_ | new_n8610_;
  assign new_n3866_ = new_n3865_ & new_n3863_;
  assign new_n3867_ = new_n3864_ | new_n3862_;
  assign new_n3868_ = new_n7821_ & new_n6887_;
  assign new_n3869_ = new_n7823_ | new_n6892_;
  assign new_n3870_ = new_n8615_ & new_n8616_;
  assign new_n3871_ = new_n8617_ | new_n8618_;
  assign new_n3872_ = new_n8620_ & new_n8616_;
  assign new_n3873_ = new_n8621_ | new_n8618_;
  assign new_n3874_ = new_n8620_ & new_n8615_;
  assign new_n3875_ = new_n8621_ | new_n8617_;
  assign new_n3876_ = new_n3875_ & new_n3873_;
  assign new_n3877_ = new_n3874_ | new_n3872_;
  assign new_n3878_ = new_n7877_ & new_n7869_;
  assign new_n3879_ = new_n7879_ | new_n7871_;
  assign new_n3880_ = new_n3878_ | new_n3876_;
  assign new_n3881_ = new_n8623_ & new_n2910_;
  assign new_n3882_ = new_n8623_ & new_n2912_;
  assign new_n3883_ = new_n3882_ | new_n3881_;
  assign new_n3884_ = new_n8625_ & new_n2959_;
  assign new_n3885_ = new_n8625_ & new_n2961_;
  assign new_n3886_ = new_n3885_ | new_n3884_;
  assign new_n3887_ = new_n8627_ & new_n3008_;
  assign new_n3888_ = new_n8627_ & new_n3010_;
  assign new_n3889_ = new_n3888_ | new_n3887_;
  assign new_n3890_ = new_n8629_ & new_n3097_;
  assign new_n3891_ = new_n8629_ & new_n3119_;
  assign new_n3892_ = new_n3891_ | new_n3890_;
  assign new_n3893_ = new_n8630_ & new_n3715_;
  assign new_n3894_ = new_n3788_ | new_n8631_;
  assign new_n3895_ = new_n6951_ & new_n7942_;
  assign new_n3896_ = new_n6964_ | new_n7945_;
  assign new_n3897_ = new_n7979_ & new_n7971_;
  assign new_n3898_ = new_n7981_ | new_n7973_;
  assign new_n3899_ = new_n8632_ & new_n8633_;
  assign new_n3900_ = new_n8634_ | new_n8635_;
  assign new_n3901_ = new_n8637_ & new_n8633_;
  assign new_n3902_ = new_n8639_ | new_n8635_;
  assign new_n3903_ = new_n8637_ & new_n8632_;
  assign new_n3904_ = new_n8639_ | new_n8634_;
  assign new_n3905_ = new_n3904_ & new_n3902_;
  assign new_n3906_ = new_n3903_ | new_n3901_;
  assign new_n3907_ = new_n7956_ & new_n7029_;
  assign new_n3908_ = new_n7957_ | new_n7044_;
  assign new_n3909_ = new_n8640_ & new_n8641_;
  assign new_n3910_ = new_n8642_ | new_n8643_;
  assign new_n3911_ = new_n8645_ & new_n8641_;
  assign new_n3912_ = new_n8647_ | new_n8643_;
  assign new_n3913_ = new_n8645_ & new_n8640_;
  assign new_n3914_ = new_n8647_ | new_n8642_;
  assign new_n3915_ = new_n3914_ & new_n3912_;
  assign new_n3916_ = new_n3913_ | new_n3911_;
  assign new_n3917_ = new_n8025_ & new_n8017_;
  assign new_n3918_ = new_n8027_ | new_n8019_;
  assign new_n3919_ = new_n3917_ | new_n3915_;
  assign new_n3920_ = new_n8051_ & new_n8047_;
  assign new_n3921_ = new_n8053_ | new_n8049_;
  assign new_n3922_ = new_n8050_ & new_n8046_;
  assign new_n3923_ = new_n8052_ | new_n8048_;
  assign new_n3924_ = new_n3923_ & new_n3921_;
  assign new_n3925_ = new_n3922_ | new_n3920_;
  assign new_n3926_ = new_n8091_ & new_n8078_;
  assign new_n3927_ = new_n8093_ | new_n8080_;
  assign new_n3928_ = new_n8648_ & new_n8649_;
  assign new_n3929_ = new_n8650_ | new_n8651_;
  assign new_n3930_ = new_n8653_ & new_n8649_;
  assign new_n3931_ = new_n8655_ | new_n8651_;
  assign new_n3932_ = new_n8653_ & new_n8648_;
  assign new_n3933_ = new_n8655_ | new_n8650_;
  assign new_n3934_ = new_n3933_ & new_n3931_;
  assign new_n3935_ = new_n3932_ | new_n3930_;
  assign new_n3936_ = new_n8083_ & new_n7029_;
  assign new_n3937_ = new_n8086_ | new_n7044_;
  assign new_n3938_ = new_n8656_ & new_n8657_;
  assign new_n3939_ = new_n8658_ | new_n8659_;
  assign new_n3940_ = new_n8661_ & new_n8657_;
  assign new_n3941_ = new_n8663_ | new_n8659_;
  assign new_n3942_ = new_n8661_ & new_n8656_;
  assign new_n3943_ = new_n8663_ | new_n8658_;
  assign new_n3944_ = new_n3943_ & new_n3941_;
  assign new_n3945_ = new_n3942_ | new_n3940_;
  assign new_n3946_ = new_n8128_ & new_n8120_;
  assign new_n3947_ = new_n8130_ | new_n8122_;
  assign new_n3948_ = new_n8664_ & new_n8665_;
  assign new_n3949_ = new_n8666_ | new_n8667_;
  assign new_n3950_ = new_n8669_ & new_n8665_;
  assign new_n3951_ = new_n8671_ | new_n8667_;
  assign new_n3952_ = new_n8669_ & new_n8664_;
  assign new_n3953_ = new_n8671_ | new_n8666_;
  assign new_n3954_ = new_n3953_ & new_n3951_;
  assign new_n3955_ = new_n3952_ | new_n3950_;
  assign new_n3956_ = new_n8105_ & new_n7598_;
  assign new_n3957_ = new_n8106_ | new_n7611_;
  assign new_n3958_ = new_n8672_ & new_n8673_;
  assign new_n3959_ = new_n8674_ | new_n8675_;
  assign new_n3960_ = new_n8677_ & new_n8673_;
  assign new_n3961_ = new_n8679_ | new_n8675_;
  assign new_n3962_ = new_n8677_ & new_n8672_;
  assign new_n3963_ = new_n8679_ | new_n8674_;
  assign new_n3964_ = new_n3963_ & new_n3961_;
  assign new_n3965_ = new_n3962_ | new_n3960_;
  assign new_n3966_ = new_n8174_ & new_n8166_;
  assign new_n3967_ = new_n8176_ | new_n8168_;
  assign new_n3968_ = new_n3966_ | new_n3964_;
  assign new_n3969_ = new_n8200_ & new_n8196_;
  assign new_n3970_ = new_n8202_ | new_n8198_;
  assign new_n3971_ = new_n8199_ & new_n8195_;
  assign new_n3972_ = new_n8201_ | new_n8197_;
  assign new_n3973_ = new_n3972_ & new_n3970_;
  assign new_n3974_ = new_n3971_ | new_n3969_;
  assign new_n3975_ = new_n8248_ & new_n8235_;
  assign new_n3976_ = new_n8250_ | new_n8237_;
  assign new_n3977_ = new_n8680_ & new_n8681_;
  assign new_n3978_ = new_n8682_ | new_n8683_;
  assign new_n3979_ = new_n8685_ & new_n8681_;
  assign new_n3980_ = new_n8687_ | new_n8683_;
  assign new_n3981_ = new_n8685_ & new_n8680_;
  assign new_n3982_ = new_n8687_ | new_n8682_;
  assign new_n3983_ = new_n3982_ & new_n3980_;
  assign new_n3984_ = new_n3981_ | new_n3979_;
  assign new_n3985_ = new_n8240_ & new_n7601_;
  assign new_n3986_ = new_n8243_ | new_n7614_;
  assign new_n3987_ = new_n8688_ & new_n8689_;
  assign new_n3988_ = new_n8690_ | new_n8691_;
  assign new_n3989_ = new_n8693_ & new_n8689_;
  assign new_n3990_ = new_n8695_ | new_n8691_;
  assign new_n3991_ = new_n8693_ & new_n8688_;
  assign new_n3992_ = new_n8695_ | new_n8690_;
  assign new_n3993_ = new_n3992_ & new_n3990_;
  assign new_n3994_ = new_n3991_ | new_n3989_;
  assign new_n3995_ = new_n8295_ & new_n8287_;
  assign new_n3996_ = new_n8297_ | new_n8289_;
  assign new_n3997_ = new_n8696_ & new_n8697_;
  assign new_n3998_ = new_n8698_ | new_n8699_;
  assign new_n3999_ = new_n8701_ & new_n8697_;
  assign new_n4000_ = new_n8703_ | new_n8699_;
  assign new_n4001_ = new_n8701_ & new_n8696_;
  assign new_n4002_ = new_n8703_ | new_n8698_;
  assign new_n4003_ = new_n4002_ & new_n4000_;
  assign new_n4004_ = new_n4001_ | new_n3999_;
  assign new_n4005_ = new_n8255_ & new_n8363_;
  assign new_n4006_ = new_n8258_ | new_n8372_;
  assign new_n4007_ = new_n8704_ & new_n8705_;
  assign new_n4008_ = new_n8706_ | new_n8707_;
  assign new_n4009_ = new_n8709_ & new_n8705_;
  assign new_n4010_ = new_n8711_ | new_n8707_;
  assign new_n4011_ = new_n8709_ & new_n8704_;
  assign new_n4012_ = new_n8711_ | new_n8706_;
  assign new_n4013_ = new_n4012_ & new_n4010_;
  assign new_n4014_ = new_n4011_ | new_n4009_;
  assign new_n4015_ = new_n8381_ & new_n8355_;
  assign new_n4016_ = new_n8383_ | new_n8357_;
  assign new_n4017_ = new_n4015_ | new_n4013_;
  assign new_n4018_ = new_n8439_ & new_n8435_;
  assign new_n4019_ = new_n8441_ | new_n8437_;
  assign new_n4020_ = new_n8438_ & new_n8434_;
  assign new_n4021_ = new_n8440_ | new_n8436_;
  assign new_n4022_ = new_n4021_ & new_n4019_;
  assign new_n4023_ = new_n4020_ | new_n4018_;
  assign new_n4024_ = new_n8423_ & new_n8419_;
  assign new_n4025_ = new_n8425_ | new_n8421_;
  assign new_n4026_ = new_n8422_ & new_n8418_;
  assign new_n4027_ = new_n8424_ | new_n8420_;
  assign new_n4028_ = new_n4027_ & new_n4025_;
  assign new_n4029_ = new_n4026_ | new_n4024_;
  assign new_n4030_ = new_n8407_ & new_n8403_;
  assign new_n4031_ = new_n8409_ | new_n8405_;
  assign new_n4032_ = new_n8406_ & new_n8402_;
  assign new_n4033_ = new_n8408_ | new_n8404_;
  assign new_n4034_ = new_n4033_ & new_n4031_;
  assign new_n4035_ = new_n4032_ | new_n4030_;
  assign new_n4036_ = new_n8534_ & new_n8517_;
  assign new_n4037_ = new_n8536_ | new_n8519_;
  assign new_n4038_ = new_n8712_ & new_n8713_;
  assign new_n4039_ = new_n8714_ | new_n8715_;
  assign new_n4040_ = new_n8717_ & new_n8713_;
  assign new_n4041_ = new_n8719_ | new_n8715_;
  assign new_n4042_ = new_n8717_ & new_n8712_;
  assign new_n4043_ = new_n8719_ | new_n8714_;
  assign new_n4044_ = new_n4043_ & new_n4041_;
  assign new_n4045_ = new_n4042_ | new_n4040_;
  assign new_n4046_ = new_n8523_ & new_n7030_;
  assign new_n4047_ = new_n8528_ | new_n7045_;
  assign new_n4048_ = new_n8720_ & new_n8721_;
  assign new_n4049_ = new_n8722_ | new_n8723_;
  assign new_n4050_ = new_n8725_ & new_n8716_;
  assign new_n4051_ = new_n8727_ | new_n8718_;
  assign new_n4052_ = new_n8728_ & new_n8729_;
  assign new_n4053_ = new_n8730_ | new_n8731_;
  assign new_n4054_ = new_n8733_ & new_n8729_;
  assign new_n4055_ = new_n8735_ | new_n8731_;
  assign new_n4056_ = new_n8733_ & new_n8728_;
  assign new_n4057_ = new_n8735_ | new_n8730_;
  assign new_n4058_ = new_n4057_ & new_n4055_;
  assign new_n4059_ = new_n4056_ | new_n4054_;
  assign new_n4060_ = new_n8524_ & new_n7601_;
  assign new_n4061_ = new_n8527_ | new_n7614_;
  assign new_n4062_ = new_n8736_ & new_n8737_;
  assign new_n4063_ = new_n8738_ | new_n8739_;
  assign new_n4064_ = new_n8741_ & new_n8732_;
  assign new_n4065_ = new_n8743_ | new_n8734_;
  assign new_n4066_ = new_n8744_ & new_n8745_;
  assign new_n4067_ = new_n8746_ | new_n8747_;
  assign new_n4068_ = new_n8749_ & new_n8745_;
  assign new_n4069_ = new_n8751_ | new_n8747_;
  assign new_n4070_ = new_n8749_ & new_n8744_;
  assign new_n4071_ = new_n8751_ | new_n8746_;
  assign new_n4072_ = new_n4071_ & new_n4069_;
  assign new_n4073_ = new_n4070_ | new_n4068_;
  assign new_n4074_ = new_n8524_ & new_n8364_;
  assign new_n4075_ = new_n8529_ | new_n8373_;
  assign new_n4076_ = new_n8752_ & new_n8753_;
  assign new_n4077_ = new_n8754_ | new_n8755_;
  assign new_n4078_ = new_n8757_ & new_n8753_;
  assign new_n4079_ = new_n8759_ | new_n8755_;
  assign new_n4080_ = new_n8757_ & new_n8752_;
  assign new_n4081_ = new_n8759_ | new_n8754_;
  assign new_n4082_ = new_n4081_ & new_n4079_;
  assign new_n4083_ = new_n4080_ | new_n4078_;
  assign new_n4084_ = new_n8741_ & new_n8737_;
  assign new_n4085_ = new_n8743_ | new_n8739_;
  assign new_n4086_ = new_n8740_ & new_n8736_;
  assign new_n4087_ = new_n8742_ | new_n8738_;
  assign new_n4088_ = new_n4087_ & new_n4085_;
  assign new_n4089_ = new_n4086_ | new_n4084_;
  assign new_n4090_ = new_n8725_ & new_n8721_;
  assign new_n4091_ = new_n8727_ | new_n8723_;
  assign new_n4092_ = new_n8724_ & new_n8720_;
  assign new_n4093_ = new_n8726_ | new_n8722_;
  assign new_n4094_ = new_n4093_ & new_n4091_;
  assign new_n4095_ = new_n4092_ | new_n4090_;
  assign new_n4096_ = new_n8550_ & new_n8542_;
  assign new_n4097_ = new_n8552_ | new_n8544_;
  assign new_n4098_ = new_n8760_ & new_n8761_;
  assign new_n4099_ = new_n8762_ | new_n8763_;
  assign new_n4100_ = new_n8765_ & new_n8761_;
  assign new_n4101_ = new_n8767_ | new_n8763_;
  assign new_n4102_ = new_n8765_ & new_n8760_;
  assign new_n4103_ = new_n8767_ | new_n8762_;
  assign new_n4104_ = new_n4103_ & new_n4101_;
  assign new_n4105_ = new_n4102_ | new_n4100_;
  assign new_n4106_ = new_n7630_ & new_n7602_;
  assign new_n4107_ = new_n7634_ | new_n7615_;
  assign new_n4108_ = new_n8768_ & new_n8769_;
  assign new_n4109_ = new_n8770_ | new_n8771_;
  assign new_n4110_ = new_n8773_ & new_n8764_;
  assign new_n4111_ = new_n8775_ | new_n8766_;
  assign new_n4112_ = new_n8776_ & new_n8777_;
  assign new_n4113_ = new_n8778_ | new_n8779_;
  assign new_n4114_ = new_n8781_ & new_n8777_;
  assign new_n4115_ = new_n8783_ | new_n8779_;
  assign new_n4116_ = new_n8781_ & new_n8776_;
  assign new_n4117_ = new_n8783_ | new_n8778_;
  assign new_n4118_ = new_n4117_ & new_n4115_;
  assign new_n4119_ = new_n4116_ | new_n4114_;
  assign new_n4120_ = new_n7632_ & new_n8364_;
  assign new_n4121_ = new_n7636_ | new_n8373_;
  assign new_n4122_ = new_n8784_ & new_n8785_;
  assign new_n4123_ = new_n8786_ | new_n8787_;
  assign new_n4124_ = new_n8789_ & new_n8780_;
  assign new_n4125_ = new_n8791_ | new_n8782_;
  assign new_n4126_ = new_n4124_ | new_n4082_;
  assign new_n4127_ = new_n7087_ & new_n8794_;
  assign new_n4128_ = new_n7095_ | new_n8797_;
  assign new_n4129_ = new_n1450_ & new_n1319_;
  assign new_n4130_ = new_n1449_ | new_n1320_;
  assign new_n4131_ = new_n8798_ & new_n8799_;
  assign new_n4132_ = new_n8800_ | new_n8801_;
  assign new_n4133_ = new_n8803_ & new_n8799_;
  assign new_n4134_ = new_n8805_ | new_n8801_;
  assign new_n4135_ = new_n8803_ & new_n8798_;
  assign new_n4136_ = new_n8805_ | new_n8800_;
  assign new_n4137_ = new_n4136_ & new_n4134_;
  assign new_n4138_ = new_n4135_ | new_n4133_;
  assign new_n4139_ = new_n7674_ & new_n8807_;
  assign new_n4140_ = new_n7689_ | new_n8810_;
  assign new_n4141_ = new_n8811_ & new_n8812_;
  assign new_n4142_ = new_n8813_ | new_n8814_;
  assign new_n4143_ = new_n8816_ & new_n8812_;
  assign new_n4144_ = new_n8818_ | new_n8814_;
  assign new_n4145_ = new_n8816_ & new_n8811_;
  assign new_n4146_ = new_n8818_ | new_n8813_;
  assign new_n4147_ = new_n4146_ & new_n4144_;
  assign new_n4148_ = new_n4145_ | new_n4143_;
  assign new_n4149_ = new_n8819_ & new_n8820_;
  assign new_n4150_ = new_n8821_ | new_n8822_;
  assign new_n4151_ = new_n8824_ & new_n8819_;
  assign new_n4152_ = new_n8826_ | new_n8821_;
  assign new_n4153_ = new_n8824_ & new_n8820_;
  assign new_n4154_ = new_n8826_ | new_n8822_;
  assign new_n4155_ = new_n4154_ & new_n4152_;
  assign new_n4156_ = new_n4153_ | new_n4151_;
  assign new_n4157_ = new_n7674_ & new_n8828_;
  assign new_n4158_ = new_n7689_ | new_n8831_;
  assign new_n4159_ = new_n8832_ & new_n8833_;
  assign new_n4160_ = new_n8834_ | new_n8835_;
  assign new_n4161_ = new_n8837_ & new_n8823_;
  assign new_n4162_ = new_n8839_ | new_n8825_;
  assign new_n4163_ = new_n8840_ & new_n8841_;
  assign new_n4164_ = new_n8842_ | new_n8843_;
  assign new_n4165_ = new_n8845_ & new_n8841_;
  assign new_n4166_ = new_n8847_ | new_n8843_;
  assign new_n4167_ = new_n8845_ & new_n8840_;
  assign new_n4168_ = new_n8847_ | new_n8842_;
  assign new_n4169_ = new_n4168_ & new_n4166_;
  assign new_n4170_ = new_n4167_ | new_n4165_;
  assign new_n4171_ = new_n8828_ & new_n7903_;
  assign new_n4172_ = new_n8831_ | new_n7918_;
  assign new_n4173_ = new_n8848_ & new_n8849_;
  assign new_n4174_ = new_n8850_ | new_n8851_;
  assign new_n4175_ = new_n8853_ & new_n8849_;
  assign new_n4176_ = new_n8855_ | new_n8851_;
  assign new_n4177_ = new_n8853_ & new_n8848_;
  assign new_n4178_ = new_n8855_ | new_n8850_;
  assign new_n4179_ = new_n4178_ & new_n4176_;
  assign new_n4180_ = new_n4177_ | new_n4175_;
  assign new_n4181_ = new_n8837_ & new_n8833_;
  assign new_n4182_ = new_n8839_ | new_n8835_;
  assign new_n4183_ = new_n8836_ & new_n8832_;
  assign new_n4184_ = new_n8838_ | new_n8834_;
  assign new_n4185_ = new_n4184_ & new_n4182_;
  assign new_n4186_ = new_n4183_ | new_n4181_;
  assign new_n4187_ = new_n1584_ & new_n1582_;
  assign new_n4188_ = new_n1583_ | new_n1581_;
  assign new_n4189_ = new_n7676_ & new_n8857_;
  assign new_n4190_ = new_n7691_ | new_n8860_;
  assign new_n4191_ = new_n8862_ & new_n8863_;
  assign new_n4192_ = new_n8864_ | new_n8865_;
  assign new_n4193_ = new_n8867_ & new_n1541_;
  assign new_n4194_ = new_n8869_ | new_n1542_;
  assign new_n4195_ = new_n8870_ & new_n8871_;
  assign new_n4196_ = new_n8872_ | new_n8873_;
  assign new_n4197_ = new_n8875_ & new_n8871_;
  assign new_n4198_ = new_n8877_ | new_n8873_;
  assign new_n4199_ = new_n8875_ & new_n8870_;
  assign new_n4200_ = new_n8877_ | new_n8872_;
  assign new_n4201_ = new_n4200_ & new_n4198_;
  assign new_n4202_ = new_n4199_ | new_n4197_;
  assign new_n4203_ = new_n8857_ & new_n7904_;
  assign new_n4204_ = new_n8860_ | new_n7919_;
  assign new_n4205_ = new_n8878_ & new_n8879_;
  assign new_n4206_ = new_n8880_ | new_n8881_;
  assign new_n4207_ = new_n8883_ & new_n8874_;
  assign new_n4208_ = new_n8885_ | new_n8876_;
  assign new_n4209_ = new_n8886_ & new_n8887_;
  assign new_n4210_ = new_n8888_ | new_n8889_;
  assign new_n4211_ = new_n8891_ & new_n8887_;
  assign new_n4212_ = new_n8893_ | new_n8889_;
  assign new_n4213_ = new_n8891_ & new_n8886_;
  assign new_n4214_ = new_n8893_ | new_n8888_;
  assign new_n4215_ = new_n4214_ & new_n4212_;
  assign new_n4216_ = new_n4213_ | new_n4211_;
  assign new_n4217_ = new_n8858_ & new_n8897_;
  assign new_n4218_ = new_n8861_ | new_n8911_;
  assign new_n4219_ = new_n8922_ & new_n8923_;
  assign new_n4220_ = new_n8924_ | new_n8925_;
  assign new_n4221_ = new_n8927_ & new_n8923_;
  assign new_n4222_ = new_n8929_ | new_n8925_;
  assign new_n4223_ = new_n8927_ & new_n8922_;
  assign new_n4224_ = new_n8929_ | new_n8924_;
  assign new_n4225_ = new_n4224_ & new_n4222_;
  assign new_n4226_ = new_n4223_ | new_n4221_;
  assign new_n4227_ = new_n8883_ & new_n8879_;
  assign new_n4228_ = new_n8885_ | new_n8881_;
  assign new_n4229_ = new_n8882_ & new_n8878_;
  assign new_n4230_ = new_n8884_ | new_n8880_;
  assign new_n4231_ = new_n4230_ & new_n4228_;
  assign new_n4232_ = new_n4229_ | new_n4227_;
  assign new_n4233_ = new_n8867_ & new_n8863_;
  assign new_n4234_ = new_n8869_ | new_n8865_;
  assign new_n4235_ = new_n8866_ & new_n8862_;
  assign new_n4236_ = new_n8868_ | new_n8864_;
  assign new_n4237_ = new_n4236_ & new_n4234_;
  assign new_n4238_ = new_n4235_ | new_n4233_;
  assign new_n4239_ = new_n8931_ & new_n1552_;
  assign new_n4240_ = new_n8933_ | new_n1551_;
  assign new_n4241_ = new_n8931_ & new_n1504_;
  assign new_n4242_ = new_n8933_ | new_n1503_;
  assign new_n4243_ = new_n4242_ & new_n4240_;
  assign new_n4244_ = new_n4241_ | new_n4239_;
  assign new_n4245_ = new_n7676_ & new_n8936_;
  assign new_n4246_ = new_n7691_ | new_n8939_;
  assign new_n4247_ = new_n8941_ & new_n8942_;
  assign new_n4248_ = new_n8943_ | new_n8944_;
  assign new_n4249_ = new_n8946_ & new_n8930_;
  assign new_n4250_ = new_n8948_ | new_n8932_;
  assign new_n4251_ = new_n8949_ & new_n8950_;
  assign new_n4252_ = new_n8951_ | new_n8952_;
  assign new_n4253_ = new_n8954_ & new_n8950_;
  assign new_n4254_ = new_n8956_ | new_n8952_;
  assign new_n4255_ = new_n8954_ & new_n8949_;
  assign new_n4256_ = new_n8956_ | new_n8951_;
  assign new_n4257_ = new_n4256_ & new_n4254_;
  assign new_n4258_ = new_n4255_ | new_n4253_;
  assign new_n4259_ = new_n8936_ & new_n7904_;
  assign new_n4260_ = new_n8939_ | new_n7919_;
  assign new_n4261_ = new_n8957_ & new_n8958_;
  assign new_n4262_ = new_n8959_ | new_n8960_;
  assign new_n4263_ = new_n8962_ & new_n8953_;
  assign new_n4264_ = new_n8964_ | new_n8955_;
  assign new_n4265_ = new_n8965_ & new_n8966_;
  assign new_n4266_ = new_n8967_ | new_n8968_;
  assign new_n4267_ = new_n8970_ & new_n8966_;
  assign new_n4268_ = new_n8972_ | new_n8968_;
  assign new_n4269_ = new_n8970_ & new_n8965_;
  assign new_n4270_ = new_n8972_ | new_n8967_;
  assign new_n4271_ = new_n4270_ & new_n4268_;
  assign new_n4272_ = new_n4269_ | new_n4267_;
  assign new_n4273_ = new_n8935_ & new_n8897_;
  assign new_n4274_ = new_n8940_ | new_n8911_;
  assign new_n4275_ = new_n8973_ & new_n8974_;
  assign new_n4276_ = new_n8975_ | new_n8976_;
  assign new_n4277_ = new_n8978_ & new_n8969_;
  assign new_n4278_ = new_n8980_ | new_n8971_;
  assign new_n4279_ = new_n8981_ & new_n8982_;
  assign new_n4280_ = new_n8983_ | new_n8984_;
  assign new_n4281_ = new_n8986_ & new_n8071_;
  assign new_n4282_ = new_n8987_ | new_n8073_;
  assign new_n4283_ = new_n8986_ & new_n8070_;
  assign new_n4284_ = new_n8987_ | new_n8072_;
  assign new_n4285_ = new_n4284_ & new_n4282_;
  assign new_n4286_ = new_n4283_ | new_n4281_;
  assign new_n4287_ = new_n8043_ & new_n7602_;
  assign new_n4288_ = new_n8044_ | new_n7615_;
  assign new_n4289_ = new_n4287_ | new_n4285_;
  assign new_n4290_ = new_n8989_ & new_n8220_;
  assign new_n4291_ = new_n8990_ | new_n8222_;
  assign new_n4292_ = new_n8989_ & new_n8219_;
  assign new_n4293_ = new_n8990_ | new_n8221_;
  assign new_n4294_ = new_n4293_ & new_n4291_;
  assign new_n4295_ = new_n4292_ | new_n4290_;
  assign new_n4296_ = new_n8192_ & new_n8366_;
  assign new_n4297_ = new_n8193_ | new_n8375_;
  assign new_n4298_ = new_n4296_ | new_n4294_;
  assign new_n4299_ = new_n8992_ & new_n8459_;
  assign new_n4300_ = new_n8993_ | new_n8461_;
  assign new_n4301_ = new_n8992_ & new_n8458_;
  assign new_n4302_ = new_n8993_ | new_n8460_;
  assign new_n4303_ = new_n4302_ & new_n4300_;
  assign new_n4304_ = new_n4301_ | new_n4299_;
  assign new_n4305_ = new_n8397_ & new_n8995_;
  assign new_n4306_ = new_n8401_ | new_n8998_;
  assign new_n4307_ = new_n4305_ | new_n4303_;
  assign new_n4308_ = new_n8789_ & new_n8785_;
  assign new_n4309_ = new_n8791_ | new_n8787_;
  assign new_n4310_ = new_n8788_ & new_n8784_;
  assign new_n4311_ = new_n8790_ | new_n8786_;
  assign new_n4312_ = new_n4311_ & new_n4309_;
  assign new_n4313_ = new_n4310_ | new_n4308_;
  assign new_n4314_ = new_n8773_ & new_n8769_;
  assign new_n4315_ = new_n8775_ | new_n8771_;
  assign new_n4316_ = new_n8772_ & new_n8768_;
  assign new_n4317_ = new_n8774_ | new_n8770_;
  assign new_n4318_ = new_n4317_ & new_n4315_;
  assign new_n4319_ = new_n4316_ | new_n4314_;
  assign new_n4320_ = new_n8566_ & new_n8558_;
  assign new_n4321_ = new_n8568_ | new_n8560_;
  assign new_n4322_ = new_n9000_ & new_n9001_;
  assign new_n4323_ = new_n9002_ | new_n9003_;
  assign new_n4324_ = new_n9005_ & new_n9001_;
  assign new_n4325_ = new_n9007_ | new_n9003_;
  assign new_n4326_ = new_n9005_ & new_n9000_;
  assign new_n4327_ = new_n9007_ | new_n9002_;
  assign new_n4328_ = new_n4327_ & new_n4325_;
  assign new_n4329_ = new_n4326_ | new_n4324_;
  assign new_n4330_ = new_n6972_ & new_n8366_;
  assign new_n4331_ = new_n6976_ | new_n8375_;
  assign new_n4332_ = new_n9008_ & new_n9009_;
  assign new_n4333_ = new_n9010_ | new_n9011_;
  assign new_n4334_ = new_n9013_ & new_n9004_;
  assign new_n4335_ = new_n9015_ | new_n9006_;
  assign new_n4336_ = new_n4334_ | new_n4312_;
  assign new_n4337_ = new_n7005_ | new_n8912_;
  assign new_n4338_ = new_n9019_ & new_n9029_;
  assign new_n4339_ = new_n9034_ | new_n9043_;
  assign new_n4340_ = new_n9047_ & new_n9029_;
  assign new_n4341_ = new_n9061_ | new_n9043_;
  assign new_n4342_ = new_n9076_ & new_n9030_;
  assign new_n4343_ = new_n9091_ | new_n9042_;
  assign new_n4344_ = new_n9047_ & new_n9104_;
  assign new_n4345_ = new_n9061_ | new_n9107_;
  assign new_n4346_ = new_n9109_ & new_n9110_;
  assign new_n4347_ = new_n9111_ | new_n9112_;
  assign new_n4348_ = new_n9113_ & new_n9110_;
  assign new_n4349_ = new_n9114_ | new_n9112_;
  assign new_n4350_ = new_n9116_ & new_n9117_;
  assign new_n4351_ = new_n9119_ | new_n9120_;
  assign new_n4352_ = new_n9122_ & new_n9117_;
  assign new_n4353_ = new_n9124_ | new_n9120_;
  assign new_n4354_ = new_n9122_ & new_n9116_;
  assign new_n4355_ = new_n9124_ | new_n9119_;
  assign new_n4356_ = new_n4355_ & new_n4353_;
  assign new_n4357_ = new_n4354_ | new_n4352_;
  assign new_n4358_ = new_n9019_ & new_n9104_;
  assign new_n4359_ = new_n9034_ | new_n9107_;
  assign new_n4360_ = new_n9125_ & new_n9126_;
  assign new_n4361_ = new_n9127_ | new_n9128_;
  assign new_n4362_ = new_n9130_ & new_n9121_;
  assign new_n4363_ = new_n9132_ | new_n9123_;
  assign new_n4364_ = new_n9133_ & new_n9134_;
  assign new_n4365_ = new_n9135_ | new_n9136_;
  assign new_n4366_ = new_n7677_ & new_n8794_;
  assign new_n4367_ = new_n7692_ | new_n8797_;
  assign new_n4368_ = new_n8815_ & new_n8802_;
  assign new_n4369_ = new_n8817_ | new_n8804_;
  assign new_n4370_ = new_n9137_ & new_n9138_;
  assign new_n4371_ = new_n9139_ | new_n9140_;
  assign new_n4372_ = new_n9142_ & new_n9138_;
  assign new_n4373_ = new_n9144_ | new_n9140_;
  assign new_n4374_ = new_n9142_ & new_n9137_;
  assign new_n4375_ = new_n9144_ | new_n9139_;
  assign new_n4376_ = new_n4375_ & new_n4373_;
  assign new_n4377_ = new_n4374_ | new_n4372_;
  assign new_n4378_ = new_n8807_ & new_n7906_;
  assign new_n4379_ = new_n8810_ | new_n7921_;
  assign new_n4380_ = new_n9145_ & new_n9146_;
  assign new_n4381_ = new_n9147_ | new_n9148_;
  assign new_n4382_ = new_n9150_ & new_n9146_;
  assign new_n4383_ = new_n9152_ | new_n9148_;
  assign new_n4384_ = new_n9150_ & new_n9145_;
  assign new_n4385_ = new_n9152_ | new_n9147_;
  assign new_n4386_ = new_n4385_ & new_n4383_;
  assign new_n4387_ = new_n4384_ | new_n4382_;
  assign new_n4388_ = new_n8852_ & new_n8844_;
  assign new_n4389_ = new_n8854_ | new_n8846_;
  assign new_n4390_ = new_n9153_ & new_n9154_;
  assign new_n4391_ = new_n9155_ | new_n9156_;
  assign new_n4392_ = new_n9158_ & new_n9154_;
  assign new_n4393_ = new_n9160_ | new_n9156_;
  assign new_n4394_ = new_n9158_ & new_n9153_;
  assign new_n4395_ = new_n9160_ | new_n9155_;
  assign new_n4396_ = new_n4395_ & new_n4393_;
  assign new_n4397_ = new_n4394_ | new_n4392_;
  assign new_n4398_ = new_n8829_ & new_n8898_;
  assign new_n4399_ = new_n8830_ | new_n8912_;
  assign new_n4400_ = new_n9161_ & new_n9162_;
  assign new_n4401_ = new_n9163_ | new_n9164_;
  assign new_n4402_ = new_n9166_ & new_n9162_;
  assign new_n4403_ = new_n9168_ | new_n9164_;
  assign new_n4404_ = new_n9166_ & new_n9161_;
  assign new_n4405_ = new_n9168_ | new_n9163_;
  assign new_n4406_ = new_n4405_ & new_n4403_;
  assign new_n4407_ = new_n4404_ | new_n4402_;
  assign new_n4408_ = new_n8926_ & new_n8890_;
  assign new_n4409_ = new_n8928_ | new_n8892_;
  assign new_n4410_ = new_n4408_ | new_n4406_;
  assign new_n4411_ = new_n1588_ & new_n1580_;
  assign new_n4412_ = new_n1587_ | new_n1579_;
  assign new_n4413_ = new_n7087_ & new_n9171_;
  assign new_n4414_ = new_n7095_ | new_n9177_;
  assign new_n4415_ = new_n9179_ & new_n9180_;
  assign new_n4416_ = new_n9181_ | new_n9182_;
  assign new_n4417_ = new_n9184_ & new_n9180_;
  assign new_n4418_ = new_n9186_ | new_n9182_;
  assign new_n4419_ = new_n9184_ & new_n9179_;
  assign new_n4420_ = new_n9186_ | new_n9181_;
  assign new_n4421_ = new_n4420_ & new_n4418_;
  assign new_n4422_ = new_n4419_ | new_n4417_;
  assign new_n4423_ = new_n9188_ & new_n1556_;
  assign new_n4424_ = new_n9190_ | new_n1555_;
  assign new_n4425_ = new_n9188_ & new_n1502_;
  assign new_n4426_ = new_n9190_ | new_n1501_;
  assign new_n4427_ = new_n4426_ & new_n4424_;
  assign new_n4428_ = new_n4425_ | new_n4423_;
  assign new_n4429_ = new_n7089_ & new_n9193_;
  assign new_n4430_ = new_n7097_ | new_n9198_;
  assign new_n4431_ = new_n9200_ & new_n9201_;
  assign new_n4432_ = new_n9202_ | new_n9203_;
  assign new_n4433_ = new_n9205_ & new_n9187_;
  assign new_n4434_ = new_n9207_ | new_n9189_;
  assign new_n4435_ = new_n9208_ & new_n9209_;
  assign new_n4436_ = new_n9210_ | new_n9211_;
  assign new_n4437_ = new_n9213_ & new_n9209_;
  assign new_n4438_ = new_n9215_ | new_n9211_;
  assign new_n4439_ = new_n9213_ & new_n9208_;
  assign new_n4440_ = new_n9215_ | new_n9210_;
  assign new_n4441_ = new_n4440_ & new_n4438_;
  assign new_n4442_ = new_n4439_ | new_n4437_;
  assign new_n4443_ = new_n7677_ & new_n9193_;
  assign new_n4444_ = new_n7692_ | new_n9198_;
  assign new_n4445_ = new_n9216_ & new_n9217_;
  assign new_n4446_ = new_n9218_ | new_n9219_;
  assign new_n4447_ = new_n9221_ & new_n9217_;
  assign new_n4448_ = new_n9223_ | new_n9219_;
  assign new_n4449_ = new_n9221_ & new_n9216_;
  assign new_n4450_ = new_n9223_ | new_n9218_;
  assign new_n4451_ = new_n4450_ & new_n4448_;
  assign new_n4452_ = new_n4449_ | new_n4447_;
  assign new_n4453_ = new_n9205_ & new_n9201_;
  assign new_n4454_ = new_n9207_ | new_n9203_;
  assign new_n4455_ = new_n9204_ & new_n9200_;
  assign new_n4456_ = new_n9206_ | new_n9202_;
  assign new_n4457_ = new_n4456_ & new_n4454_;
  assign new_n4458_ = new_n4455_ | new_n4453_;
  assign new_n4459_ = new_n9224_ & new_n9225_;
  assign new_n4460_ = new_n9226_ | new_n9227_;
  assign new_n4461_ = new_n9229_ & new_n9224_;
  assign new_n4462_ = new_n9231_ | new_n9226_;
  assign new_n4463_ = new_n9229_ & new_n9225_;
  assign new_n4464_ = new_n9231_ | new_n9227_;
  assign new_n4465_ = new_n4464_ & new_n4462_;
  assign new_n4466_ = new_n4463_ | new_n4461_;
  assign new_n4467_ = new_n7089_ & new_n9234_;
  assign new_n4468_ = new_n7097_ | new_n9239_;
  assign new_n4469_ = new_n9241_ & new_n9242_;
  assign new_n4470_ = new_n9243_ | new_n9244_;
  assign new_n4471_ = new_n9246_ & new_n9228_;
  assign new_n4472_ = new_n9248_ | new_n9230_;
  assign new_n4473_ = new_n9249_ & new_n9250_;
  assign new_n4474_ = new_n9251_ | new_n9252_;
  assign new_n4475_ = new_n9254_ & new_n9250_;
  assign new_n4476_ = new_n9256_ | new_n9252_;
  assign new_n4477_ = new_n9254_ & new_n9249_;
  assign new_n4478_ = new_n9256_ | new_n9251_;
  assign new_n4479_ = new_n4478_ & new_n4476_;
  assign new_n4480_ = new_n4477_ | new_n4475_;
  assign new_n4481_ = new_n7680_ & new_n9234_;
  assign new_n4482_ = new_n7695_ | new_n9239_;
  assign new_n4483_ = new_n9257_ & new_n9258_;
  assign new_n4484_ = new_n9259_ | new_n9260_;
  assign new_n4485_ = new_n9262_ & new_n9253_;
  assign new_n4486_ = new_n9264_ | new_n9255_;
  assign new_n4487_ = new_n9265_ & new_n9266_;
  assign new_n4488_ = new_n9267_ | new_n9268_;
  assign new_n4489_ = new_n9270_ & new_n9266_;
  assign new_n4490_ = new_n9272_ | new_n9268_;
  assign new_n4491_ = new_n9270_ & new_n9265_;
  assign new_n4492_ = new_n9272_ | new_n9267_;
  assign new_n4493_ = new_n4492_ & new_n4490_;
  assign new_n4494_ = new_n4491_ | new_n4489_;
  assign new_n4495_ = new_n9235_ & new_n7906_;
  assign new_n4496_ = new_n9238_ | new_n7921_;
  assign new_n4497_ = new_n9273_ & new_n9274_;
  assign new_n4498_ = new_n9275_ | new_n9276_;
  assign new_n4499_ = new_n9278_ & new_n9274_;
  assign new_n4500_ = new_n9280_ | new_n9276_;
  assign new_n4501_ = new_n9278_ & new_n9273_;
  assign new_n4502_ = new_n9280_ | new_n9275_;
  assign new_n4503_ = new_n4502_ & new_n4500_;
  assign new_n4504_ = new_n4501_ | new_n4499_;
  assign new_n4505_ = new_n9262_ & new_n9258_;
  assign new_n4506_ = new_n9264_ | new_n9260_;
  assign new_n4507_ = new_n9261_ & new_n9257_;
  assign new_n4508_ = new_n9263_ | new_n9259_;
  assign new_n4509_ = new_n4508_ & new_n4506_;
  assign new_n4510_ = new_n4507_ | new_n4505_;
  assign new_n4511_ = new_n9246_ & new_n9242_;
  assign new_n4512_ = new_n9248_ | new_n9244_;
  assign new_n4513_ = new_n9245_ & new_n9241_;
  assign new_n4514_ = new_n9247_ | new_n9243_;
  assign new_n4515_ = new_n4514_ & new_n4512_;
  assign new_n4516_ = new_n4513_ | new_n4511_;
  assign new_n4517_ = new_n1590_ & new_n1575_;
  assign new_n4518_ = new_n1589_ | new_n1576_;
  assign new_n4519_ = new_n9282_ & new_n1395_;
  assign new_n4520_ = new_n9284_ | new_n1396_;
  assign new_n4521_ = new_n9285_ & new_n9286_;
  assign new_n4522_ = new_n9287_ | new_n9288_;
  assign new_n4523_ = new_n9290_ & new_n9286_;
  assign new_n4524_ = new_n9292_ | new_n9288_;
  assign new_n4525_ = new_n9290_ & new_n9285_;
  assign new_n4526_ = new_n9292_ | new_n9287_;
  assign new_n4527_ = new_n4526_ & new_n4524_;
  assign new_n4528_ = new_n4525_ | new_n4523_;
  assign new_n4529_ = new_n7090_ & new_n9295_;
  assign new_n4530_ = new_n7098_ | new_n9300_;
  assign new_n4531_ = new_n9302_ & new_n9303_;
  assign new_n4532_ = new_n9304_ | new_n9305_;
  assign new_n4533_ = new_n9307_ & new_n9289_;
  assign new_n4534_ = new_n9309_ | new_n9291_;
  assign new_n4535_ = new_n9310_ & new_n9311_;
  assign new_n4536_ = new_n9312_ | new_n9313_;
  assign new_n4537_ = new_n9315_ & new_n9311_;
  assign new_n4538_ = new_n9317_ | new_n9313_;
  assign new_n4539_ = new_n9315_ & new_n9310_;
  assign new_n4540_ = new_n9317_ | new_n9312_;
  assign new_n4541_ = new_n4540_ & new_n4538_;
  assign new_n4542_ = new_n4539_ | new_n4537_;
  assign new_n4543_ = new_n7680_ & new_n9295_;
  assign new_n4544_ = new_n7695_ | new_n9300_;
  assign new_n4545_ = new_n9318_ & new_n9319_;
  assign new_n4546_ = new_n9320_ | new_n9321_;
  assign new_n4547_ = new_n9323_ & new_n9314_;
  assign new_n4548_ = new_n9325_ | new_n9316_;
  assign new_n4549_ = new_n9326_ & new_n9327_;
  assign new_n4550_ = new_n9328_ | new_n9329_;
  assign new_n4551_ = new_n9331_ & new_n9327_;
  assign new_n4552_ = new_n9333_ | new_n9329_;
  assign new_n4553_ = new_n9331_ & new_n9326_;
  assign new_n4554_ = new_n9333_ | new_n9328_;
  assign new_n4555_ = new_n4554_ & new_n4552_;
  assign new_n4556_ = new_n4553_ | new_n4551_;
  assign new_n4557_ = new_n9296_ & new_n7907_;
  assign new_n4558_ = new_n9299_ | new_n7922_;
  assign new_n4559_ = new_n9334_ & new_n9335_;
  assign new_n4560_ = new_n9336_ | new_n9337_;
  assign new_n4561_ = new_n9339_ & new_n9330_;
  assign new_n4562_ = new_n9341_ | new_n9332_;
  assign new_n4563_ = new_n9342_ & new_n9343_;
  assign new_n4564_ = new_n9344_ | new_n9345_;
  assign new_n4565_ = new_n9347_ & new_n9343_;
  assign new_n4566_ = new_n9349_ | new_n9345_;
  assign new_n4567_ = new_n9347_ & new_n9342_;
  assign new_n4568_ = new_n9349_ | new_n9344_;
  assign new_n4569_ = new_n4568_ & new_n4566_;
  assign new_n4570_ = new_n4567_ | new_n4565_;
  assign new_n4571_ = new_n9296_ & new_n8898_;
  assign new_n4572_ = new_n9301_ | new_n8914_;
  assign new_n4573_ = new_n9350_ & new_n9351_;
  assign new_n4574_ = new_n9352_ | new_n9353_;
  assign new_n4575_ = new_n9355_ & new_n9351_;
  assign new_n4576_ = new_n9357_ | new_n9353_;
  assign new_n4577_ = new_n9355_ & new_n9350_;
  assign new_n4578_ = new_n9357_ | new_n9352_;
  assign new_n4579_ = new_n4578_ & new_n4576_;
  assign new_n4580_ = new_n4577_ | new_n4575_;
  assign new_n4581_ = new_n9339_ & new_n9335_;
  assign new_n4582_ = new_n9341_ | new_n9337_;
  assign new_n4583_ = new_n9338_ & new_n9334_;
  assign new_n4584_ = new_n9340_ | new_n9336_;
  assign new_n4585_ = new_n4584_ & new_n4582_;
  assign new_n4586_ = new_n4583_ | new_n4581_;
  assign new_n4587_ = new_n9323_ & new_n9319_;
  assign new_n4588_ = new_n9325_ | new_n9321_;
  assign new_n4589_ = new_n9322_ & new_n9318_;
  assign new_n4590_ = new_n9324_ | new_n9320_;
  assign new_n4591_ = new_n4590_ & new_n4588_;
  assign new_n4592_ = new_n4589_ | new_n4587_;
  assign new_n4593_ = new_n9307_ & new_n9303_;
  assign new_n4594_ = new_n9309_ | new_n9305_;
  assign new_n4595_ = new_n9306_ & new_n9302_;
  assign new_n4596_ = new_n9308_ | new_n9304_;
  assign new_n4597_ = new_n4596_ & new_n4594_;
  assign new_n4598_ = new_n4595_ | new_n4593_;
  assign new_n4599_ = new_n9282_ & new_n1557_;
  assign new_n4600_ = new_n9284_ | new_n1558_;
  assign new_n4601_ = new_n9281_ & new_n1492_;
  assign new_n4602_ = new_n9283_ | new_n1491_;
  assign new_n4603_ = new_n4602_ & new_n4600_;
  assign new_n4604_ = new_n4601_ | new_n4599_;
  assign new_n4605_ = new_n8466_ & new_n1467_;
  assign new_n4606_ = new_n8468_ | new_n1468_;
  assign new_n4607_ = new_n9358_ & new_n9359_;
  assign new_n4608_ = new_n9360_ | new_n9361_;
  assign new_n4609_ = new_n9363_ & new_n9359_;
  assign new_n4610_ = new_n9365_ | new_n9361_;
  assign new_n4611_ = new_n9363_ & new_n9358_;
  assign new_n4612_ = new_n9365_ | new_n9360_;
  assign new_n4613_ = new_n4612_ & new_n4610_;
  assign new_n4614_ = new_n4611_ | new_n4609_;
  assign new_n4615_ = new_n7090_ & new_n9368_;
  assign new_n4616_ = new_n7098_ | new_n9372_;
  assign new_n4617_ = new_n9374_ & new_n9375_;
  assign new_n4618_ = new_n9376_ | new_n9377_;
  assign new_n4619_ = new_n9379_ & new_n9362_;
  assign new_n4620_ = new_n9381_ | new_n9364_;
  assign new_n4621_ = new_n9382_ & new_n9383_;
  assign new_n4622_ = new_n9384_ | new_n9385_;
  assign new_n4623_ = new_n9387_ & new_n9383_;
  assign new_n4624_ = new_n9389_ | new_n9385_;
  assign new_n4625_ = new_n9387_ & new_n9382_;
  assign new_n4626_ = new_n9389_ | new_n9384_;
  assign new_n4627_ = new_n4626_ & new_n4624_;
  assign new_n4628_ = new_n4625_ | new_n4623_;
  assign new_n4629_ = new_n7681_ & new_n9368_;
  assign new_n4630_ = new_n7696_ | new_n9372_;
  assign new_n4631_ = new_n9390_ & new_n9391_;
  assign new_n4632_ = new_n9392_ | new_n9393_;
  assign new_n4633_ = new_n9395_ & new_n9386_;
  assign new_n4634_ = new_n9397_ | new_n9388_;
  assign new_n4635_ = new_n9398_ & new_n9399_;
  assign new_n4636_ = new_n9400_ | new_n9401_;
  assign new_n4637_ = new_n9403_ & new_n9399_;
  assign new_n4638_ = new_n9405_ | new_n9401_;
  assign new_n4639_ = new_n9403_ & new_n9398_;
  assign new_n4640_ = new_n9405_ | new_n9400_;
  assign new_n4641_ = new_n4640_ & new_n4638_;
  assign new_n4642_ = new_n4639_ | new_n4637_;
  assign new_n4643_ = new_n9367_ & new_n7907_;
  assign new_n4644_ = new_n9371_ | new_n7922_;
  assign new_n4645_ = new_n9406_ & new_n9407_;
  assign new_n4646_ = new_n9408_ | new_n9409_;
  assign new_n4647_ = new_n9411_ & new_n9402_;
  assign new_n4648_ = new_n9413_ | new_n9404_;
  assign new_n4649_ = new_n9414_ & new_n9415_;
  assign new_n4650_ = new_n9416_ | new_n9417_;
  assign new_n4651_ = new_n9419_ & new_n9415_;
  assign new_n4652_ = new_n9421_ | new_n9417_;
  assign new_n4653_ = new_n9419_ & new_n9414_;
  assign new_n4654_ = new_n9421_ | new_n9416_;
  assign new_n4655_ = new_n4654_ & new_n4652_;
  assign new_n4656_ = new_n4653_ | new_n4651_;
  assign new_n4657_ = new_n9369_ & new_n8900_;
  assign new_n4658_ = new_n9373_ | new_n8914_;
  assign new_n4659_ = new_n9422_ & new_n9423_;
  assign new_n4660_ = new_n9424_ | new_n9425_;
  assign new_n4661_ = new_n9427_ & new_n9418_;
  assign new_n4662_ = new_n9429_ | new_n9420_;
  assign new_n4663_ = new_n4661_ | new_n4579_;
  assign new_n4664_ = new_n8962_ & new_n8958_;
  assign new_n4665_ = new_n8964_ | new_n8960_;
  assign new_n4666_ = new_n8961_ & new_n8957_;
  assign new_n4667_ = new_n8963_ | new_n8959_;
  assign new_n4668_ = new_n4667_ & new_n4665_;
  assign new_n4669_ = new_n4666_ | new_n4664_;
  assign new_n4670_ = new_n8946_ & new_n8942_;
  assign new_n4671_ = new_n8948_ | new_n8944_;
  assign new_n4672_ = new_n8945_ & new_n8941_;
  assign new_n4673_ = new_n8947_ | new_n8943_;
  assign new_n4674_ = new_n4673_ & new_n4671_;
  assign new_n4675_ = new_n4672_ | new_n4670_;
  assign new_n4676_ = new_n9430_ & new_n9431_;
  assign new_n4677_ = new_n9432_ | new_n9433_;
  assign new_n4678_ = new_n9435_ & new_n9430_;
  assign new_n4679_ = new_n9437_ | new_n9432_;
  assign new_n4680_ = new_n9435_ & new_n9431_;
  assign new_n4681_ = new_n9437_ | new_n9433_;
  assign new_n4682_ = new_n4681_ & new_n4679_;
  assign new_n4683_ = new_n4680_ | new_n4678_;
  assign new_n4684_ = new_n7681_ & new_n9440_;
  assign new_n4685_ = new_n7696_ | new_n9443_;
  assign new_n4686_ = new_n9445_ & new_n9446_;
  assign new_n4687_ = new_n9447_ | new_n9448_;
  assign new_n4688_ = new_n9450_ & new_n9434_;
  assign new_n4689_ = new_n9452_ | new_n9436_;
  assign new_n4690_ = new_n9453_ & new_n9454_;
  assign new_n4691_ = new_n9455_ | new_n9456_;
  assign new_n4692_ = new_n9458_ & new_n9454_;
  assign new_n4693_ = new_n9460_ | new_n9456_;
  assign new_n4694_ = new_n9458_ & new_n9453_;
  assign new_n4695_ = new_n9460_ | new_n9455_;
  assign new_n4696_ = new_n4695_ & new_n4693_;
  assign new_n4697_ = new_n4694_ | new_n4692_;
  assign new_n4698_ = new_n9440_ & new_n7910_;
  assign new_n4699_ = new_n9443_ | new_n7925_;
  assign new_n4700_ = new_n9461_ & new_n9462_;
  assign new_n4701_ = new_n9463_ | new_n9464_;
  assign new_n4702_ = new_n9466_ & new_n9457_;
  assign new_n4703_ = new_n9468_ | new_n9459_;
  assign new_n4704_ = new_n9469_ & new_n9470_;
  assign new_n4705_ = new_n9471_ | new_n9472_;
  assign new_n4706_ = new_n9474_ & new_n9470_;
  assign new_n4707_ = new_n9476_ | new_n9472_;
  assign new_n4708_ = new_n9474_ & new_n9469_;
  assign new_n4709_ = new_n9476_ | new_n9471_;
  assign new_n4710_ = new_n4709_ & new_n4707_;
  assign new_n4711_ = new_n4708_ | new_n4706_;
  assign new_n4712_ = new_n9439_ & new_n8900_;
  assign new_n4713_ = new_n9444_ | new_n8915_;
  assign new_n4714_ = new_n9477_ & new_n9478_;
  assign new_n4715_ = new_n9479_ | new_n9480_;
  assign new_n4716_ = new_n9482_ & new_n9478_;
  assign new_n4717_ = new_n9484_ | new_n9480_;
  assign new_n4718_ = new_n9482_ & new_n9477_;
  assign new_n4719_ = new_n9484_ | new_n9479_;
  assign new_n4720_ = new_n4719_ & new_n4717_;
  assign new_n4721_ = new_n4718_ | new_n4716_;
  assign new_n4722_ = new_n9466_ & new_n9462_;
  assign new_n4723_ = new_n9468_ | new_n9464_;
  assign new_n4724_ = new_n9465_ & new_n9461_;
  assign new_n4725_ = new_n9467_ | new_n9463_;
  assign new_n4726_ = new_n4725_ & new_n4723_;
  assign new_n4727_ = new_n4724_ | new_n4722_;
  assign new_n4728_ = new_n9450_ & new_n9446_;
  assign new_n4729_ = new_n9452_ | new_n9448_;
  assign new_n4730_ = new_n9449_ & new_n9445_;
  assign new_n4731_ = new_n9451_ | new_n9447_;
  assign new_n4732_ = new_n4731_ & new_n4729_;
  assign new_n4733_ = new_n4730_ | new_n4728_;
  assign new_n4734_ = new_n1592_ & new_n1573_;
  assign new_n4735_ = new_n1591_ | new_n1574_;
  assign new_n4736_ = new_n9486_ & new_n1397_;
  assign new_n4737_ = new_n9488_ | new_n1398_;
  assign new_n4738_ = new_n9489_ & new_n9490_;
  assign new_n4739_ = new_n9491_ | new_n9492_;
  assign new_n4740_ = new_n9494_ & new_n9490_;
  assign new_n4741_ = new_n9496_ | new_n9492_;
  assign new_n4742_ = new_n9494_ & new_n9489_;
  assign new_n4743_ = new_n9496_ | new_n9491_;
  assign new_n4744_ = new_n4743_ & new_n4741_;
  assign new_n4745_ = new_n4742_ | new_n4740_;
  assign new_n4746_ = new_n7683_ & new_n9499_;
  assign new_n4747_ = new_n7698_ | new_n9502_;
  assign new_n4748_ = new_n9504_ & new_n9505_;
  assign new_n4749_ = new_n9506_ | new_n9507_;
  assign new_n4750_ = new_n9509_ & new_n9493_;
  assign new_n4751_ = new_n9511_ | new_n9495_;
  assign new_n4752_ = new_n9512_ & new_n9513_;
  assign new_n4753_ = new_n9514_ | new_n9515_;
  assign new_n4754_ = new_n9517_ & new_n9513_;
  assign new_n4755_ = new_n9519_ | new_n9515_;
  assign new_n4756_ = new_n9517_ & new_n9512_;
  assign new_n4757_ = new_n9519_ | new_n9514_;
  assign new_n4758_ = new_n4757_ & new_n4755_;
  assign new_n4759_ = new_n4756_ | new_n4754_;
  assign new_n4760_ = new_n9499_ & new_n7910_;
  assign new_n4761_ = new_n9502_ | new_n7925_;
  assign new_n4762_ = new_n9520_ & new_n9521_;
  assign new_n4763_ = new_n9522_ | new_n9523_;
  assign new_n4764_ = new_n9525_ & new_n9516_;
  assign new_n4765_ = new_n9527_ | new_n9518_;
  assign new_n4766_ = new_n9528_ & new_n9529_;
  assign new_n4767_ = new_n9530_ | new_n9531_;
  assign new_n4768_ = new_n9533_ & new_n9529_;
  assign new_n4769_ = new_n9535_ | new_n9531_;
  assign new_n4770_ = new_n9533_ & new_n9528_;
  assign new_n4771_ = new_n9535_ | new_n9530_;
  assign new_n4772_ = new_n4771_ & new_n4769_;
  assign new_n4773_ = new_n4770_ | new_n4768_;
  assign new_n4774_ = new_n9498_ & new_n8901_;
  assign new_n4775_ = new_n9503_ | new_n8915_;
  assign new_n4776_ = new_n9536_ & new_n9537_;
  assign new_n4777_ = new_n9538_ | new_n9539_;
  assign new_n4778_ = new_n9541_ & new_n9532_;
  assign new_n4779_ = new_n9543_ | new_n9534_;
  assign new_n4780_ = new_n9544_ & new_n9545_;
  assign new_n4781_ = new_n9546_ | new_n9547_;
  assign new_n4782_ = new_n9549_ & new_n9545_;
  assign new_n4783_ = new_n9551_ | new_n9547_;
  assign new_n4784_ = new_n9549_ & new_n9544_;
  assign new_n4785_ = new_n9551_ | new_n9546_;
  assign new_n4786_ = new_n4785_ & new_n4783_;
  assign new_n4787_ = new_n4784_ | new_n4782_;
  assign new_n4788_ = new_n9500_ & new_n9555_;
  assign new_n4789_ = new_n9503_ | new_n9564_;
  assign new_n4790_ = new_n9570_ & new_n9571_;
  assign new_n4791_ = new_n9572_ | new_n9573_;
  assign new_n4792_ = new_n9575_ & new_n9571_;
  assign new_n4793_ = new_n9577_ | new_n9573_;
  assign new_n4794_ = new_n9575_ & new_n9570_;
  assign new_n4795_ = new_n9577_ | new_n9572_;
  assign new_n4796_ = new_n4795_ & new_n4793_;
  assign new_n4797_ = new_n4794_ | new_n4792_;
  assign new_n4798_ = new_n9541_ & new_n9537_;
  assign new_n4799_ = new_n9543_ | new_n9539_;
  assign new_n4800_ = new_n9540_ & new_n9536_;
  assign new_n4801_ = new_n9542_ | new_n9538_;
  assign new_n4802_ = new_n4801_ & new_n4799_;
  assign new_n4803_ = new_n4800_ | new_n4798_;
  assign new_n4804_ = new_n9525_ & new_n9521_;
  assign new_n4805_ = new_n9527_ | new_n9523_;
  assign new_n4806_ = new_n9524_ & new_n9520_;
  assign new_n4807_ = new_n9526_ | new_n9522_;
  assign new_n4808_ = new_n4807_ & new_n4805_;
  assign new_n4809_ = new_n4806_ | new_n4804_;
  assign new_n4810_ = new_n9509_ & new_n9505_;
  assign new_n4811_ = new_n9511_ | new_n9507_;
  assign new_n4812_ = new_n9508_ & new_n9504_;
  assign new_n4813_ = new_n9510_ | new_n9506_;
  assign new_n4814_ = new_n4813_ & new_n4811_;
  assign new_n4815_ = new_n4812_ | new_n4810_;
  assign new_n4816_ = new_n9486_ & new_n1559_;
  assign new_n4817_ = new_n9488_ | new_n1560_;
  assign new_n4818_ = new_n9485_ & new_n1490_;
  assign new_n4819_ = new_n9487_ | new_n1489_;
  assign new_n4820_ = new_n4819_ & new_n4817_;
  assign new_n4821_ = new_n4818_ | new_n4816_;
  assign new_n4822_ = new_n9578_ & new_n9579_;
  assign new_n4823_ = new_n9580_ | new_n9581_;
  assign new_n4824_ = new_n9583_ & new_n1469_;
  assign new_n4825_ = new_n9585_ | new_n1470_;
  assign new_n4826_ = new_n9586_ & new_n9587_;
  assign new_n4827_ = new_n9588_ | new_n9589_;
  assign new_n4828_ = new_n9591_ & new_n9587_;
  assign new_n4829_ = new_n9593_ | new_n9589_;
  assign new_n4830_ = new_n9591_ & new_n9586_;
  assign new_n4831_ = new_n9593_ | new_n9588_;
  assign new_n4832_ = new_n4831_ & new_n4829_;
  assign new_n4833_ = new_n4830_ | new_n4828_;
  assign new_n4834_ = new_n7683_ & new_n9596_;
  assign new_n4835_ = new_n7698_ | new_n9600_;
  assign new_n4836_ = new_n9602_ & new_n9603_;
  assign new_n4837_ = new_n9604_ | new_n9605_;
  assign new_n4838_ = new_n9607_ & new_n9590_;
  assign new_n4839_ = new_n9609_ | new_n9592_;
  assign new_n4840_ = new_n9610_ & new_n9611_;
  assign new_n4841_ = new_n9612_ | new_n9613_;
  assign new_n4842_ = new_n9615_ & new_n9611_;
  assign new_n4843_ = new_n9617_ | new_n9613_;
  assign new_n4844_ = new_n9615_ & new_n9610_;
  assign new_n4845_ = new_n9617_ | new_n9612_;
  assign new_n4846_ = new_n4845_ & new_n4843_;
  assign new_n4847_ = new_n4844_ | new_n4842_;
  assign new_n4848_ = new_n9596_ & new_n7911_;
  assign new_n4849_ = new_n9600_ | new_n7926_;
  assign new_n4850_ = new_n9618_ & new_n9619_;
  assign new_n4851_ = new_n9620_ | new_n9621_;
  assign new_n4852_ = new_n9623_ & new_n9614_;
  assign new_n4853_ = new_n9625_ | new_n9616_;
  assign new_n4854_ = new_n9626_ & new_n9627_;
  assign new_n4855_ = new_n9628_ | new_n9629_;
  assign new_n4856_ = new_n9631_ & new_n9627_;
  assign new_n4857_ = new_n9633_ | new_n9629_;
  assign new_n4858_ = new_n9631_ & new_n9626_;
  assign new_n4859_ = new_n9633_ | new_n9628_;
  assign new_n4860_ = new_n4859_ & new_n4857_;
  assign new_n4861_ = new_n4858_ | new_n4856_;
  assign new_n4862_ = new_n9595_ & new_n8901_;
  assign new_n4863_ = new_n9599_ | new_n8918_;
  assign new_n4864_ = new_n9634_ & new_n9635_;
  assign new_n4865_ = new_n9636_ | new_n9637_;
  assign new_n4866_ = new_n9639_ & new_n9630_;
  assign new_n4867_ = new_n9641_ | new_n9632_;
  assign new_n4868_ = new_n9642_ & new_n9643_;
  assign new_n4869_ = new_n9644_ | new_n9645_;
  assign new_n4870_ = new_n9647_ & new_n9643_;
  assign new_n4871_ = new_n9649_ | new_n9645_;
  assign new_n4872_ = new_n9647_ & new_n9642_;
  assign new_n4873_ = new_n9649_ | new_n9644_;
  assign new_n4874_ = new_n4873_ & new_n4871_;
  assign new_n4875_ = new_n4872_ | new_n4870_;
  assign new_n4876_ = new_n9597_ & new_n9555_;
  assign new_n4877_ = new_n9601_ | new_n9564_;
  assign new_n4878_ = new_n9650_ & new_n9651_;
  assign new_n4879_ = new_n9652_ | new_n9653_;
  assign new_n4880_ = new_n9655_ & new_n9646_;
  assign new_n4881_ = new_n9657_ | new_n9648_;
  assign new_n4882_ = new_n4880_ | new_n4796_;
  assign new_n4883_ = new_n9379_ & new_n9375_;
  assign new_n4884_ = new_n9381_ | new_n9377_;
  assign new_n4885_ = new_n9378_ & new_n9374_;
  assign new_n4886_ = new_n9380_ | new_n9376_;
  assign new_n4887_ = new_n4886_ & new_n4884_;
  assign new_n4888_ = new_n4885_ | new_n4883_;
  assign new_n4889_ = new_n8482_ & new_n8474_;
  assign new_n4890_ = new_n8484_ | new_n8476_;
  assign new_n4891_ = new_n9658_ & new_n9659_;
  assign new_n4892_ = new_n9660_ | new_n9661_;
  assign new_n4893_ = new_n9663_ & new_n9659_;
  assign new_n4894_ = new_n9665_ | new_n9661_;
  assign new_n4895_ = new_n9663_ & new_n9658_;
  assign new_n4896_ = new_n9665_ | new_n9660_;
  assign new_n4897_ = new_n4896_ & new_n4894_;
  assign new_n4898_ = new_n4895_ | new_n4893_;
  assign new_n4899_ = new_n7684_ & new_n7705_;
  assign new_n4900_ = new_n7699_ | new_n7709_;
  assign new_n4901_ = new_n9666_ & new_n9667_;
  assign new_n4902_ = new_n9668_ | new_n9669_;
  assign new_n4903_ = new_n9671_ & new_n9667_;
  assign new_n4904_ = new_n9673_ | new_n9669_;
  assign new_n4905_ = new_n9671_ & new_n9666_;
  assign new_n4906_ = new_n9673_ | new_n9668_;
  assign new_n4907_ = new_n4906_ & new_n4904_;
  assign new_n4908_ = new_n4905_ | new_n4903_;
  assign new_n4909_ = new_n8498_ & new_n8490_;
  assign new_n4910_ = new_n8500_ | new_n8492_;
  assign new_n4911_ = new_n9674_ & new_n9675_;
  assign new_n4912_ = new_n9676_ | new_n9677_;
  assign new_n4913_ = new_n9679_ & new_n9675_;
  assign new_n4914_ = new_n9681_ | new_n9677_;
  assign new_n4915_ = new_n9679_ & new_n9674_;
  assign new_n4916_ = new_n9681_ | new_n9676_;
  assign new_n4917_ = new_n4916_ & new_n4914_;
  assign new_n4918_ = new_n4915_ | new_n4913_;
  assign new_n4919_ = new_n7106_ & new_n7911_;
  assign new_n4920_ = new_n7111_ | new_n7926_;
  assign new_n4921_ = new_n9682_ & new_n9683_;
  assign new_n4922_ = new_n9684_ | new_n9685_;
  assign new_n4923_ = new_n9687_ & new_n9683_;
  assign new_n4924_ = new_n9689_ | new_n9685_;
  assign new_n4925_ = new_n9687_ & new_n9682_;
  assign new_n4926_ = new_n9689_ | new_n9684_;
  assign new_n4927_ = new_n4926_ & new_n4924_;
  assign new_n4928_ = new_n4925_ | new_n4923_;
  assign new_n4929_ = new_n3717_ & new_n8507_;
  assign new_n4930_ = new_n9690_ | new_n8509_;
  assign new_n4931_ = new_n9691_ & new_n9692_;
  assign new_n4932_ = new_n4929_ | new_n4927_;
  assign new_n4933_ = new_n9693_ & new_n9692_;
  assign new_n4934_ = new_n9693_ & new_n9691_;
  assign new_n4935_ = new_n4934_ | new_n4933_;
  assign new_n4936_ = new_n7988_ | new_n7616_;
  assign new_n4937_ = new_n8137_ | new_n8376_;
  assign new_n4938_ = new_n8310_ | new_n8998_;
  assign new_n4939_ = new_n7636_ | new_n8999_;
  assign new_n4940_ = new_n8591_ & new_n8584_;
  assign new_n4941_ = new_n8605_ & new_n8598_;
  assign new_n4942_ = new_n8619_ & new_n8612_;
  assign new_n4943_ = new_n9695_ & new_n3821_;
  assign new_n4944_ = new_n9697_ & new_n3850_;
  assign new_n4945_ = new_n9699_ & new_n3879_;
  assign new_n4946_ = new_n9699_ & new_n3877_;
  assign new_n4947_ = new_n9697_ & new_n3848_;
  assign new_n4948_ = new_n9695_ & new_n3819_;
  assign new_n4949_ = new_n9700_ & new_n9701_;
  assign new_n4950_ = new_n9702_ & new_n9703_;
  assign new_n4951_ = new_n9704_ & new_n9705_;
  assign new_n4952_ = new_n9706_ & new_n9707_;
  assign new_n4953_ = new_n9709_ & new_n3141_;
  assign new_n4954_ = new_n9709_ & new_n3143_;
  assign new_n4955_ = new_n4954_ | new_n4953_;
  assign new_n4956_ = new_n9711_ & new_n3150_;
  assign new_n4957_ = new_n9711_ & new_n3152_;
  assign new_n4958_ = new_n4957_ | new_n4956_;
  assign new_n4959_ = new_n9713_ & new_n3159_;
  assign new_n4960_ = new_n9713_ & new_n3161_;
  assign new_n4961_ = new_n4960_ | new_n4959_;
  assign new_n4962_ = new_n7943_ & new_n7030_;
  assign new_n4963_ = new_n7944_ | new_n7045_;
  assign new_n4964_ = new_n8644_ & new_n8636_;
  assign new_n4965_ = new_n8646_ | new_n8638_;
  assign new_n4966_ = new_n4964_ | new_n4962_;
  assign new_n4967_ = new_n8067_ & new_n8063_;
  assign new_n4968_ = new_n8069_ | new_n8065_;
  assign new_n4969_ = new_n8066_ & new_n8062_;
  assign new_n4970_ = new_n8068_ | new_n8064_;
  assign new_n4971_ = new_n4970_ & new_n4968_;
  assign new_n4972_ = new_n4969_ | new_n4967_;
  assign new_n4973_ = new_n8660_ & new_n8652_;
  assign new_n4974_ = new_n8662_ | new_n8654_;
  assign new_n4975_ = new_n9714_ & new_n9715_;
  assign new_n4976_ = new_n9716_ | new_n9717_;
  assign new_n4977_ = new_n9719_ & new_n9715_;
  assign new_n4978_ = new_n9720_ | new_n9717_;
  assign new_n4979_ = new_n9719_ & new_n9714_;
  assign new_n4980_ = new_n9720_ | new_n9716_;
  assign new_n4981_ = new_n4980_ & new_n4978_;
  assign new_n4982_ = new_n4979_ | new_n4977_;
  assign new_n4983_ = new_n8084_ & new_n7603_;
  assign new_n4984_ = new_n8085_ | new_n7616_;
  assign new_n4985_ = new_n9721_ & new_n9722_;
  assign new_n4986_ = new_n9723_ | new_n9724_;
  assign new_n4987_ = new_n9726_ & new_n9722_;
  assign new_n4988_ = new_n9727_ | new_n9724_;
  assign new_n4989_ = new_n9726_ & new_n9721_;
  assign new_n4990_ = new_n9727_ | new_n9723_;
  assign new_n4991_ = new_n4990_ & new_n4988_;
  assign new_n4992_ = new_n4989_ | new_n4987_;
  assign new_n4993_ = new_n8676_ & new_n8668_;
  assign new_n4994_ = new_n8678_ | new_n8670_;
  assign new_n4995_ = new_n4993_ | new_n4991_;
  assign new_n4996_ = new_n8216_ & new_n8212_;
  assign new_n4997_ = new_n8218_ | new_n8214_;
  assign new_n4998_ = new_n8215_ & new_n8211_;
  assign new_n4999_ = new_n8217_ | new_n8213_;
  assign new_n5000_ = new_n4999_ & new_n4997_;
  assign new_n5001_ = new_n4998_ | new_n4996_;
  assign new_n5002_ = new_n8692_ & new_n8684_;
  assign new_n5003_ = new_n8694_ | new_n8686_;
  assign new_n5004_ = new_n9728_ & new_n9729_;
  assign new_n5005_ = new_n9730_ | new_n9731_;
  assign new_n5006_ = new_n9733_ & new_n9729_;
  assign new_n5007_ = new_n9734_ | new_n9731_;
  assign new_n5008_ = new_n9733_ & new_n9728_;
  assign new_n5009_ = new_n9734_ | new_n9730_;
  assign new_n5010_ = new_n5009_ & new_n5007_;
  assign new_n5011_ = new_n5008_ | new_n5006_;
  assign new_n5012_ = new_n8241_ & new_n8367_;
  assign new_n5013_ = new_n8242_ | new_n8376_;
  assign new_n5014_ = new_n9735_ & new_n9736_;
  assign new_n5015_ = new_n9737_ | new_n9738_;
  assign new_n5016_ = new_n9740_ & new_n9736_;
  assign new_n5017_ = new_n9741_ | new_n9738_;
  assign new_n5018_ = new_n9740_ & new_n9735_;
  assign new_n5019_ = new_n9741_ | new_n9737_;
  assign new_n5020_ = new_n5019_ & new_n5017_;
  assign new_n5021_ = new_n5018_ | new_n5016_;
  assign new_n5022_ = new_n8708_ & new_n8700_;
  assign new_n5023_ = new_n8710_ | new_n8702_;
  assign new_n5024_ = new_n5022_ | new_n5020_;
  assign new_n5025_ = new_n9013_ & new_n9009_;
  assign new_n5026_ = new_n9015_ | new_n9011_;
  assign new_n5027_ = new_n9012_ & new_n9008_;
  assign new_n5028_ = new_n9014_ | new_n9010_;
  assign new_n5029_ = new_n5028_ & new_n5026_;
  assign new_n5030_ = new_n5027_ | new_n5025_;
  assign new_n5031_ = new_n3894_ & new_n8575_;
  assign new_n5032_ = new_n9742_ | new_n8577_;
  assign new_n5033_ = new_n5031_ | new_n5029_;
  assign new_n5034_ = new_n9744_ & new_n3916_;
  assign new_n5035_ = new_n9744_ & new_n3918_;
  assign new_n5036_ = new_n5035_ | new_n5034_;
  assign new_n5037_ = new_n9746_ & new_n3965_;
  assign new_n5038_ = new_n9746_ & new_n3967_;
  assign new_n5039_ = new_n5038_ | new_n5037_;
  assign new_n5040_ = new_n9748_ & new_n4014_;
  assign new_n5041_ = new_n9748_ & new_n4016_;
  assign new_n5042_ = new_n5041_ | new_n5040_;
  assign new_n5043_ = new_n9750_ & new_n4083_;
  assign new_n5044_ = new_n9750_ & new_n4125_;
  assign new_n5045_ = new_n5044_ | new_n5043_;
  assign new_n5046_ = new_n9752_ & new_n8982_;
  assign new_n5047_ = new_n9753_ | new_n8984_;
  assign new_n5048_ = new_n9752_ & new_n8981_;
  assign new_n5049_ = new_n9753_ | new_n8983_;
  assign new_n5050_ = new_n5049_ & new_n5047_;
  assign new_n5051_ = new_n5048_ | new_n5046_;
  assign new_n5052_ = new_n8937_ & new_n9556_;
  assign new_n5053_ = new_n8940_ | new_n9565_;
  assign new_n5054_ = new_n5052_ | new_n5050_;
  assign new_n5055_ = new_n9754_ & new_n9755_;
  assign new_n5056_ = new_n9427_ & new_n9423_;
  assign new_n5057_ = new_n9429_ | new_n9425_;
  assign new_n5058_ = new_n9426_ & new_n9422_;
  assign new_n5059_ = new_n9428_ | new_n9424_;
  assign new_n5060_ = new_n5059_ & new_n5057_;
  assign new_n5061_ = new_n5058_ | new_n5056_;
  assign new_n5062_ = new_n9411_ & new_n9407_;
  assign new_n5063_ = new_n9413_ | new_n9409_;
  assign new_n5064_ = new_n9410_ & new_n9406_;
  assign new_n5065_ = new_n9412_ | new_n9408_;
  assign new_n5066_ = new_n5065_ & new_n5063_;
  assign new_n5067_ = new_n5064_ | new_n5062_;
  assign new_n5068_ = new_n9395_ & new_n9391_;
  assign new_n5069_ = new_n9397_ | new_n9393_;
  assign new_n5070_ = new_n9394_ & new_n9390_;
  assign new_n5071_ = new_n9396_ | new_n9392_;
  assign new_n5072_ = new_n5071_ & new_n5069_;
  assign new_n5073_ = new_n5070_ | new_n5068_;
  assign new_n5074_ = new_n9670_ & new_n9662_;
  assign new_n5075_ = new_n9672_ | new_n9664_;
  assign new_n5076_ = new_n9756_ & new_n9757_;
  assign new_n5077_ = new_n9758_ | new_n9759_;
  assign new_n5078_ = new_n9761_ & new_n9757_;
  assign new_n5079_ = new_n9763_ | new_n9759_;
  assign new_n5080_ = new_n9761_ & new_n9756_;
  assign new_n5081_ = new_n9763_ | new_n9758_;
  assign new_n5082_ = new_n5081_ & new_n5079_;
  assign new_n5083_ = new_n5080_ | new_n5078_;
  assign new_n5084_ = new_n7705_ & new_n7913_;
  assign new_n5085_ = new_n7711_ | new_n7928_;
  assign new_n5086_ = new_n9764_ & new_n9765_;
  assign new_n5087_ = new_n9766_ | new_n9767_;
  assign new_n5088_ = new_n9769_ & new_n9760_;
  assign new_n5089_ = new_n9771_ | new_n9762_;
  assign new_n5090_ = new_n9772_ & new_n9773_;
  assign new_n5091_ = new_n9774_ | new_n9775_;
  assign new_n5092_ = new_n9777_ & new_n9773_;
  assign new_n5093_ = new_n9779_ | new_n9775_;
  assign new_n5094_ = new_n9777_ & new_n9772_;
  assign new_n5095_ = new_n9779_ | new_n9774_;
  assign new_n5096_ = new_n5095_ & new_n5093_;
  assign new_n5097_ = new_n5094_ | new_n5092_;
  assign new_n5098_ = new_n7707_ & new_n8904_;
  assign new_n5099_ = new_n7711_ | new_n8918_;
  assign new_n5100_ = new_n9780_ & new_n9781_;
  assign new_n5101_ = new_n9782_ | new_n9783_;
  assign new_n5102_ = new_n9785_ & new_n9776_;
  assign new_n5103_ = new_n9787_ | new_n9778_;
  assign new_n5104_ = new_n5102_ | new_n5060_;
  assign new_n5105_ = new_n9655_ & new_n9651_;
  assign new_n5106_ = new_n9657_ | new_n9653_;
  assign new_n5107_ = new_n9654_ & new_n9650_;
  assign new_n5108_ = new_n9656_ | new_n9652_;
  assign new_n5109_ = new_n5108_ & new_n5106_;
  assign new_n5110_ = new_n5107_ | new_n5105_;
  assign new_n5111_ = new_n9639_ & new_n9635_;
  assign new_n5112_ = new_n9641_ | new_n9637_;
  assign new_n5113_ = new_n9638_ & new_n9634_;
  assign new_n5114_ = new_n9640_ | new_n9636_;
  assign new_n5115_ = new_n5114_ & new_n5112_;
  assign new_n5116_ = new_n5113_ | new_n5111_;
  assign new_n5117_ = new_n9623_ & new_n9619_;
  assign new_n5118_ = new_n9625_ | new_n9621_;
  assign new_n5119_ = new_n9622_ & new_n9618_;
  assign new_n5120_ = new_n9624_ | new_n9620_;
  assign new_n5121_ = new_n5120_ & new_n5118_;
  assign new_n5122_ = new_n5119_ | new_n5117_;
  assign new_n5123_ = new_n9607_ & new_n9603_;
  assign new_n5124_ = new_n9609_ | new_n9605_;
  assign new_n5125_ = new_n9606_ & new_n9602_;
  assign new_n5126_ = new_n9608_ | new_n9604_;
  assign new_n5127_ = new_n5126_ & new_n5124_;
  assign new_n5128_ = new_n5125_ | new_n5123_;
  assign new_n5129_ = new_n9583_ & new_n9578_;
  assign new_n5130_ = new_n9585_ | new_n9580_;
  assign new_n5131_ = new_n9582_ & new_n9579_;
  assign new_n5132_ = new_n9584_ | new_n9581_;
  assign new_n5133_ = new_n5132_ & new_n5130_;
  assign new_n5134_ = new_n5131_ | new_n5129_;
  assign new_n5135_ = new_n9183_ & new_n1539_;
  assign new_n5136_ = new_n9185_ | new_n1540_;
  assign new_n5137_ = new_n9788_ & new_n9789_;
  assign new_n5138_ = new_n9790_ | new_n9791_;
  assign new_n5139_ = new_n9793_ & new_n9789_;
  assign new_n5140_ = new_n9795_ | new_n9791_;
  assign new_n5141_ = new_n9793_ & new_n9788_;
  assign new_n5142_ = new_n9795_ | new_n9790_;
  assign new_n5143_ = new_n5142_ & new_n5140_;
  assign new_n5144_ = new_n5141_ | new_n5139_;
  assign new_n5145_ = new_n7684_ & new_n9171_;
  assign new_n5146_ = new_n7699_ | new_n9177_;
  assign new_n5147_ = new_n9796_ & new_n9797_;
  assign new_n5148_ = new_n9798_ | new_n9799_;
  assign new_n5149_ = new_n9801_ & new_n9792_;
  assign new_n5150_ = new_n9803_ | new_n9794_;
  assign new_n5151_ = new_n9804_ & new_n9805_;
  assign new_n5152_ = new_n9806_ | new_n9807_;
  assign new_n5153_ = new_n9809_ & new_n9805_;
  assign new_n5154_ = new_n9811_ | new_n9807_;
  assign new_n5155_ = new_n9809_ & new_n9804_;
  assign new_n5156_ = new_n9811_ | new_n9806_;
  assign new_n5157_ = new_n5156_ & new_n5154_;
  assign new_n5158_ = new_n5155_ | new_n5153_;
  assign new_n5159_ = new_n9172_ & new_n7913_;
  assign new_n5160_ = new_n9176_ | new_n7928_;
  assign new_n5161_ = new_n9812_ & new_n9813_;
  assign new_n5162_ = new_n9814_ | new_n9815_;
  assign new_n5163_ = new_n9817_ & new_n9808_;
  assign new_n5164_ = new_n9819_ | new_n9810_;
  assign new_n5165_ = new_n9820_ & new_n9821_;
  assign new_n5166_ = new_n9822_ | new_n9823_;
  assign new_n5167_ = new_n9825_ & new_n9821_;
  assign new_n5168_ = new_n9827_ | new_n9823_;
  assign new_n5169_ = new_n9825_ & new_n9820_;
  assign new_n5170_ = new_n9827_ | new_n9822_;
  assign new_n5171_ = new_n5170_ & new_n5168_;
  assign new_n5172_ = new_n5169_ | new_n5167_;
  assign new_n5173_ = new_n9172_ & new_n8904_;
  assign new_n5174_ = new_n9178_ | new_n8919_;
  assign new_n5175_ = new_n9828_ & new_n9829_;
  assign new_n5176_ = new_n9830_ | new_n9831_;
  assign new_n5177_ = new_n9833_ & new_n9824_;
  assign new_n5178_ = new_n9835_ | new_n9826_;
  assign new_n5179_ = new_n9836_ & new_n9837_;
  assign new_n5180_ = new_n9838_ | new_n9839_;
  assign new_n5181_ = new_n9841_ & new_n9837_;
  assign new_n5182_ = new_n9843_ | new_n9839_;
  assign new_n5183_ = new_n9841_ & new_n9836_;
  assign new_n5184_ = new_n9843_ | new_n9838_;
  assign new_n5185_ = new_n5184_ & new_n5182_;
  assign new_n5186_ = new_n5183_ | new_n5181_;
  assign new_n5187_ = new_n9174_ & new_n9556_;
  assign new_n5188_ = new_n9178_ | new_n9565_;
  assign new_n5189_ = new_n9844_ & new_n9845_;
  assign new_n5190_ = new_n9846_ | new_n9847_;
  assign new_n5191_ = new_n9849_ & new_n9840_;
  assign new_n5192_ = new_n9851_ | new_n9842_;
  assign new_n5193_ = new_n5191_ | new_n5109_;
  assign new_n5194_ = new_n9076_ & new_n9853_;
  assign new_n5195_ = new_n9091_ | new_n9856_;
  assign new_n5196_ = new_n9048_ & new_n9858_;
  assign new_n5197_ = new_n9062_ | new_n9861_;
  assign new_n5198_ = new_n9862_ & new_n9863_;
  assign new_n5199_ = new_n9864_ | new_n9865_;
  assign new_n5200_ = new_n9866_ & new_n9863_;
  assign new_n5201_ = new_n9867_ | new_n9865_;
  assign new_n5202_ = new_n9866_ & new_n9862_;
  assign new_n5203_ = new_n9867_ | new_n9864_;
  assign new_n5204_ = new_n5203_ & new_n9869_;
  assign new_n5205_ = new_n5202_ | new_n9871_;
  assign new_n5206_ = new_n9077_ & new_n9858_;
  assign new_n5207_ = new_n9092_ | new_n9861_;
  assign new_n5208_ = new_n9048_ & new_n9873_;
  assign new_n5209_ = new_n9062_ | new_n9875_;
  assign new_n5210_ = new_n9876_ & new_n9877_;
  assign new_n5211_ = new_n9878_ | new_n9879_;
  assign new_n5212_ = new_n9880_ & new_n9877_;
  assign new_n5213_ = new_n9881_ | new_n9879_;
  assign new_n5214_ = new_n9882_ | new_n5204_;
  assign new_n5215_ = new_n9077_ & new_n9885_;
  assign new_n5216_ = new_n9092_ | new_n9888_;
  assign new_n5217_ = new_n9050_ & new_n9892_;
  assign new_n5218_ = new_n9064_ | new_n9895_;
  assign new_n5219_ = new_n9897_ & new_n9898_;
  assign new_n5220_ = new_n9899_ | new_n9900_;
  assign new_n5221_ = new_n9901_ & new_n9898_;
  assign new_n5222_ = new_n9902_ | new_n9900_;
  assign new_n5223_ = new_n9901_ & new_n9897_;
  assign new_n5224_ = new_n9902_ | new_n9899_;
  assign new_n5225_ = new_n5224_ & new_n9904_;
  assign new_n5226_ = new_n5223_ | new_n9906_;
  assign new_n5227_ = new_n9079_ & new_n9892_;
  assign new_n5228_ = new_n9094_ | new_n9895_;
  assign new_n5229_ = new_n9050_ & new_n9909_;
  assign new_n5230_ = new_n9064_ | new_n9912_;
  assign new_n5231_ = new_n9914_ & new_n9915_;
  assign new_n5232_ = new_n9916_ | new_n9917_;
  assign new_n5233_ = new_n9918_ & new_n9915_;
  assign new_n5234_ = new_n9919_ | new_n9917_;
  assign new_n5235_ = new_n9921_ & new_n9922_;
  assign new_n5236_ = new_n9924_ | new_n9925_;
  assign new_n5237_ = new_n9927_ & new_n9922_;
  assign new_n5238_ = new_n9929_ | new_n9925_;
  assign new_n5239_ = new_n9927_ & new_n9921_;
  assign new_n5240_ = new_n9929_ | new_n9924_;
  assign new_n5241_ = new_n5240_ & new_n5238_;
  assign new_n5242_ = new_n5239_ | new_n5237_;
  assign new_n5243_ = new_n9020_ & new_n9909_;
  assign new_n5244_ = new_n9035_ | new_n9912_;
  assign new_n5245_ = new_n9930_ & new_n9931_;
  assign new_n5246_ = new_n9932_ | new_n9933_;
  assign new_n5247_ = new_n9935_ & new_n9931_;
  assign new_n5248_ = new_n9937_ | new_n9933_;
  assign new_n5249_ = new_n9935_ & new_n9930_;
  assign new_n5250_ = new_n9937_ | new_n9932_;
  assign new_n5251_ = new_n5250_ & new_n5248_;
  assign new_n5252_ = new_n5249_ | new_n5247_;
  assign new_n5253_ = new_n9918_ & new_n9914_;
  assign new_n5254_ = new_n9919_ | new_n9916_;
  assign new_n5255_ = new_n5254_ & new_n9920_;
  assign new_n5256_ = new_n5253_ | new_n9923_;
  assign new_n5257_ = new_n9079_ & new_n9908_;
  assign new_n5258_ = new_n9094_ | new_n9913_;
  assign new_n5259_ = new_n9051_ & new_n9939_;
  assign new_n5260_ = new_n9065_ | new_n9942_;
  assign new_n5261_ = new_n9944_ & new_n9945_;
  assign new_n5262_ = new_n9946_ | new_n9947_;
  assign new_n5263_ = new_n9948_ & new_n9945_;
  assign new_n5264_ = new_n9949_ | new_n9947_;
  assign new_n5265_ = new_n9951_ & new_n9952_;
  assign new_n5266_ = new_n9954_ | new_n9955_;
  assign new_n5267_ = new_n9957_ & new_n9952_;
  assign new_n5268_ = new_n9959_ | new_n9955_;
  assign new_n5269_ = new_n9957_ & new_n9951_;
  assign new_n5270_ = new_n9959_ | new_n9954_;
  assign new_n5271_ = new_n5270_ & new_n5268_;
  assign new_n5272_ = new_n5269_ | new_n5267_;
  assign new_n5273_ = new_n9020_ & new_n9939_;
  assign new_n5274_ = new_n9035_ | new_n9942_;
  assign new_n5275_ = new_n9960_ & new_n9961_;
  assign new_n5276_ = new_n9962_ | new_n9963_;
  assign new_n5277_ = new_n9965_ & new_n9956_;
  assign new_n5278_ = new_n9967_ | new_n9958_;
  assign new_n5279_ = new_n5277_ | new_n5251_;
  assign new_n5280_ = new_n6972_ & new_n8995_;
  assign new_n5281_ = new_n8861_ | new_n9566_;
  assign new_n5282_ = new_n9601_ | new_n902_;
  assign new_n5283_ = new_n9373_ | new_n9566_;
  assign new_n5284_ = new_n9065_ | new_n810_;
  assign new_n5285_ = new_n9725_ & new_n9718_;
  assign new_n5286_ = new_n9739_ & new_n9732_;
  assign new_n5287_ = new_n8455_ & new_n8451_;
  assign new_n5288_ = new_n8457_ | new_n8453_;
  assign new_n5289_ = new_n8454_ & new_n8450_;
  assign new_n5290_ = new_n8456_ | new_n8452_;
  assign new_n5291_ = new_n5290_ & new_n5288_;
  assign new_n5292_ = new_n5289_ | new_n5287_;
  assign new_n5293_ = new_n8756_ & new_n8748_;
  assign new_n5294_ = new_n8758_ | new_n8750_;
  assign new_n5295_ = new_n9968_ & new_n9969_;
  assign new_n5296_ = new_n9970_ | new_n9971_;
  assign new_n5297_ = new_n9973_ & new_n9969_;
  assign new_n5298_ = new_n9974_ | new_n9971_;
  assign new_n5299_ = new_n9973_ & new_n9968_;
  assign new_n5300_ = new_n9974_ | new_n9970_;
  assign new_n5301_ = new_n5300_ & new_n5298_;
  assign new_n5302_ = new_n5299_ | new_n5297_;
  assign new_n5303_ = new_n8525_ & new_n8996_;
  assign new_n5304_ = new_n8529_ | new_n8999_;
  assign new_n5305_ = new_n5303_ | new_n5301_;
  assign new_n5306_ = new_n9976_ & new_n9972_;
  assign new_n5307_ = new_n9977_ | new_n4931_;
  assign new_n5308_ = new_n9817_ & new_n9813_;
  assign new_n5309_ = new_n9819_ | new_n9815_;
  assign new_n5310_ = new_n9816_ & new_n9812_;
  assign new_n5311_ = new_n9818_ | new_n9814_;
  assign new_n5312_ = new_n5311_ & new_n5309_;
  assign new_n5313_ = new_n5310_ | new_n5308_;
  assign new_n5314_ = new_n9801_ & new_n9797_;
  assign new_n5315_ = new_n9803_ | new_n9799_;
  assign new_n5316_ = new_n9800_ & new_n9796_;
  assign new_n5317_ = new_n9802_ | new_n9798_;
  assign new_n5318_ = new_n5317_ & new_n5315_;
  assign new_n5319_ = new_n5316_ | new_n5314_;
  assign new_n5320_ = new_n9220_ & new_n9212_;
  assign new_n5321_ = new_n9222_ | new_n9214_;
  assign new_n5322_ = new_n9978_ & new_n9979_;
  assign new_n5323_ = new_n9980_ | new_n9981_;
  assign new_n5324_ = new_n9983_ & new_n9979_;
  assign new_n5325_ = new_n9985_ | new_n9981_;
  assign new_n5326_ = new_n9983_ & new_n9978_;
  assign new_n5327_ = new_n9985_ | new_n9980_;
  assign new_n5328_ = new_n5327_ & new_n5325_;
  assign new_n5329_ = new_n5326_ | new_n5324_;
  assign new_n5330_ = new_n9194_ & new_n7914_;
  assign new_n5331_ = new_n9197_ | new_n7929_;
  assign new_n5332_ = new_n9986_ & new_n9987_;
  assign new_n5333_ = new_n9988_ | new_n9989_;
  assign new_n5334_ = new_n9991_ & new_n9982_;
  assign new_n5335_ = new_n9993_ | new_n9984_;
  assign new_n5336_ = new_n9994_ & new_n9995_;
  assign new_n5337_ = new_n9996_ | new_n9997_;
  assign new_n5338_ = new_n9999_ & new_n9995_;
  assign new_n5339_ = new_n10001_ | new_n9997_;
  assign new_n5340_ = new_n9999_ & new_n9994_;
  assign new_n5341_ = new_n10001_ | new_n9996_;
  assign new_n5342_ = new_n5341_ & new_n5339_;
  assign new_n5343_ = new_n5340_ | new_n5338_;
  assign new_n5344_ = new_n9194_ & new_n8905_;
  assign new_n5345_ = new_n9199_ | new_n8919_;
  assign new_n5346_ = new_n10002_ & new_n10003_;
  assign new_n5347_ = new_n10004_ | new_n10005_;
  assign new_n5348_ = new_n10007_ & new_n10003_;
  assign new_n5349_ = new_n10009_ | new_n10005_;
  assign new_n5350_ = new_n10007_ & new_n10002_;
  assign new_n5351_ = new_n10009_ | new_n10004_;
  assign new_n5352_ = new_n5351_ & new_n5349_;
  assign new_n5353_ = new_n5350_ | new_n5348_;
  assign new_n5354_ = new_n9991_ & new_n9987_;
  assign new_n5355_ = new_n9993_ | new_n9989_;
  assign new_n5356_ = new_n9990_ & new_n9986_;
  assign new_n5357_ = new_n9992_ | new_n9988_;
  assign new_n5358_ = new_n5357_ & new_n5355_;
  assign new_n5359_ = new_n5356_ | new_n5354_;
  assign new_n5360_ = new_n9277_ & new_n9269_;
  assign new_n5361_ = new_n9279_ | new_n9271_;
  assign new_n5362_ = new_n10010_ & new_n10011_;
  assign new_n5363_ = new_n10012_ | new_n10013_;
  assign new_n5364_ = new_n10015_ & new_n10011_;
  assign new_n5365_ = new_n10017_ | new_n10013_;
  assign new_n5366_ = new_n10015_ & new_n10010_;
  assign new_n5367_ = new_n10017_ | new_n10012_;
  assign new_n5368_ = new_n5367_ & new_n5365_;
  assign new_n5369_ = new_n5366_ | new_n5364_;
  assign new_n5370_ = new_n9235_ & new_n8905_;
  assign new_n5371_ = new_n9240_ | new_n8921_;
  assign new_n5372_ = new_n10018_ & new_n10019_;
  assign new_n5373_ = new_n10020_ | new_n10021_;
  assign new_n5374_ = new_n10023_ & new_n10014_;
  assign new_n5375_ = new_n10025_ | new_n10016_;
  assign new_n5376_ = new_n10026_ & new_n10027_;
  assign new_n5377_ = new_n10028_ | new_n10029_;
  assign new_n5378_ = new_n10031_ & new_n10027_;
  assign new_n5379_ = new_n10032_ | new_n10029_;
  assign new_n5380_ = new_n10031_ & new_n10026_;
  assign new_n5381_ = new_n10032_ | new_n10028_;
  assign new_n5382_ = new_n5381_ & new_n5379_;
  assign new_n5383_ = new_n5380_ | new_n5378_;
  assign new_n5384_ = new_n9236_ & new_n9557_;
  assign new_n5385_ = new_n9240_ | new_n9568_;
  assign new_n5386_ = new_n5384_ | new_n5382_;
  assign new_n5387_ = new_n10034_ & new_n10030_;
  assign new_n5388_ = new_n10036_ & new_n4963_;
  assign new_n5389_ = new_n9976_ & new_n5304_;
  assign new_n5390_ = new_n10036_ & new_n4965_;
  assign new_n5391_ = new_n10038_ & new_n4994_;
  assign new_n5392_ = new_n10040_ & new_n5023_;
  assign new_n5393_ = new_n10042_ & new_n5032_;
  assign new_n5394_ = new_n10038_ & new_n4992_;
  assign new_n5395_ = new_n10040_ & new_n5021_;
  assign new_n5396_ = new_n10042_ & new_n5030_;
  assign new_n5397_ = new_n9975_ & new_n5302_;
  assign new_n5398_ = new_n10043_ & new_n10044_;
  assign new_n5399_ = new_n10045_ & new_n10046_;
  assign new_n5400_ = new_n10047_ & new_n10048_;
  assign new_n5401_ = new_n10049_ & new_n10050_;
  assign new_n5402_ = new_n10052_ & new_n9134_;
  assign new_n5403_ = new_n10053_ | new_n9136_;
  assign new_n5404_ = new_n10052_ & new_n9133_;
  assign new_n5405_ = new_n10053_ | new_n9135_;
  assign new_n5406_ = new_n5405_ & new_n5403_;
  assign new_n5407_ = new_n5404_ | new_n5402_;
  assign new_n5408_ = new_n10056_ & new_n9103_;
  assign new_n5409_ = new_n10062_ | new_n9108_;
  assign new_n5410_ = new_n5408_ | new_n5406_;
  assign new_n5411_ = new_n8793_ & new_n7914_;
  assign new_n5412_ = new_n8796_ | new_n7929_;
  assign new_n5413_ = new_n9149_ & new_n9141_;
  assign new_n5414_ = new_n9151_ | new_n9143_;
  assign new_n5415_ = new_n10065_ & new_n10066_;
  assign new_n5416_ = new_n10067_ | new_n10068_;
  assign new_n5417_ = new_n10070_ & new_n10066_;
  assign new_n5418_ = new_n10071_ | new_n10068_;
  assign new_n5419_ = new_n10070_ & new_n10065_;
  assign new_n5420_ = new_n10071_ | new_n10067_;
  assign new_n5421_ = new_n5420_ & new_n5418_;
  assign new_n5422_ = new_n5419_ | new_n5417_;
  assign new_n5423_ = new_n8808_ & new_n8907_;
  assign new_n5424_ = new_n8809_ | new_n8921_;
  assign new_n5425_ = new_n10072_ & new_n10073_;
  assign new_n5426_ = new_n10074_ | new_n10075_;
  assign new_n5427_ = new_n10077_ & new_n10073_;
  assign new_n5428_ = new_n10078_ | new_n10075_;
  assign new_n5429_ = new_n10077_ & new_n10072_;
  assign new_n5430_ = new_n10078_ | new_n10074_;
  assign new_n5431_ = new_n5430_ & new_n5428_;
  assign new_n5432_ = new_n5429_ | new_n5427_;
  assign new_n5433_ = new_n9165_ & new_n9157_;
  assign new_n5434_ = new_n9167_ | new_n9159_;
  assign new_n5435_ = new_n5433_ | new_n5431_;
  assign new_n5436_ = new_n8978_ & new_n8974_;
  assign new_n5437_ = new_n8980_ | new_n8976_;
  assign new_n5438_ = new_n8977_ & new_n8973_;
  assign new_n5439_ = new_n8979_ | new_n8975_;
  assign new_n5440_ = new_n5439_ & new_n5437_;
  assign new_n5441_ = new_n5438_ | new_n5436_;
  assign new_n5442_ = new_n9481_ & new_n9473_;
  assign new_n5443_ = new_n9483_ | new_n9475_;
  assign new_n5444_ = new_n10079_ & new_n10080_;
  assign new_n5445_ = new_n10081_ | new_n10082_;
  assign new_n5446_ = new_n10084_ & new_n10080_;
  assign new_n5447_ = new_n10085_ | new_n10082_;
  assign new_n5448_ = new_n10084_ & new_n10079_;
  assign new_n5449_ = new_n10085_ | new_n10081_;
  assign new_n5450_ = new_n5449_ & new_n5447_;
  assign new_n5451_ = new_n5448_ | new_n5446_;
  assign new_n5452_ = new_n9441_ & new_n9557_;
  assign new_n5453_ = new_n9444_ | new_n9568_;
  assign new_n5454_ = new_n10086_ & new_n10087_;
  assign new_n5455_ = new_n10088_ | new_n10089_;
  assign new_n5456_ = new_n10091_ & new_n10087_;
  assign new_n5457_ = new_n10092_ | new_n10089_;
  assign new_n5458_ = new_n10091_ & new_n10086_;
  assign new_n5459_ = new_n10092_ | new_n10088_;
  assign new_n5460_ = new_n5459_ & new_n5457_;
  assign new_n5461_ = new_n5458_ | new_n5456_;
  assign new_n5462_ = new_n9574_ & new_n9548_;
  assign new_n5463_ = new_n9576_ | new_n9550_;
  assign new_n5464_ = new_n5462_ | new_n5460_;
  assign new_n5465_ = new_n9785_ & new_n9781_;
  assign new_n5466_ = new_n9787_ | new_n9783_;
  assign new_n5467_ = new_n9784_ & new_n9780_;
  assign new_n5468_ = new_n9786_ | new_n9782_;
  assign new_n5469_ = new_n5468_ & new_n5466_;
  assign new_n5470_ = new_n5467_ | new_n5465_;
  assign new_n5471_ = new_n9769_ & new_n9765_;
  assign new_n5472_ = new_n9771_ | new_n9767_;
  assign new_n5473_ = new_n9768_ & new_n9764_;
  assign new_n5474_ = new_n9770_ | new_n9766_;
  assign new_n5475_ = new_n5474_ & new_n5472_;
  assign new_n5476_ = new_n5473_ | new_n5471_;
  assign new_n5477_ = new_n9686_ & new_n9678_;
  assign new_n5478_ = new_n9688_ | new_n9680_;
  assign new_n5479_ = new_n10093_ & new_n10094_;
  assign new_n5480_ = new_n10095_ | new_n10096_;
  assign new_n5481_ = new_n10098_ & new_n10094_;
  assign new_n5482_ = new_n10100_ | new_n10096_;
  assign new_n5483_ = new_n10098_ & new_n10093_;
  assign new_n5484_ = new_n10100_ | new_n10095_;
  assign new_n5485_ = new_n5484_ & new_n5482_;
  assign new_n5486_ = new_n5483_ | new_n5481_;
  assign new_n5487_ = new_n7107_ & new_n8907_;
  assign new_n5488_ = new_n7111_ | new_n8920_;
  assign new_n5489_ = new_n10101_ & new_n10102_;
  assign new_n5490_ = new_n5487_ | new_n5485_;
  assign new_n5491_ = new_n10104_ & new_n10097_;
  assign new_n5492_ = new_n5489_ | new_n10099_;
  assign new_n5493_ = new_n5491_ | new_n5469_;
  assign new_n5494_ = new_n9849_ & new_n9845_;
  assign new_n5495_ = new_n9851_ | new_n9847_;
  assign new_n5496_ = new_n9848_ & new_n9844_;
  assign new_n5497_ = new_n9850_ | new_n9846_;
  assign new_n5498_ = new_n5497_ & new_n5495_;
  assign new_n5499_ = new_n5496_ | new_n5494_;
  assign new_n5500_ = new_n9833_ & new_n9829_;
  assign new_n5501_ = new_n9835_ | new_n9831_;
  assign new_n5502_ = new_n9832_ & new_n9828_;
  assign new_n5503_ = new_n9834_ | new_n9830_;
  assign new_n5504_ = new_n5503_ & new_n5501_;
  assign new_n5505_ = new_n5502_ | new_n5500_;
  assign new_n5506_ = new_n10006_ & new_n9998_;
  assign new_n5507_ = new_n10008_ | new_n10000_;
  assign new_n5508_ = new_n10105_ & new_n10106_;
  assign new_n5509_ = new_n10107_ | new_n10108_;
  assign new_n5510_ = new_n10110_ & new_n10106_;
  assign new_n5511_ = new_n10112_ | new_n10108_;
  assign new_n5512_ = new_n10110_ & new_n10105_;
  assign new_n5513_ = new_n10112_ | new_n10107_;
  assign new_n5514_ = new_n5513_ & new_n5511_;
  assign new_n5515_ = new_n5512_ | new_n5510_;
  assign new_n5516_ = new_n9195_ & new_n9559_;
  assign new_n5517_ = new_n9199_ | new_n9569_;
  assign new_n5518_ = new_n5517_ & new_n5515_;
  assign new_n5519_ = new_n10113_ | new_n10114_;
  assign new_n5520_ = new_n5519_ & new_n10109_;
  assign new_n5521_ = new_n10116_ | new_n10111_;
  assign new_n5522_ = new_n5520_ | new_n5498_;
  assign new_n5523_ = new_n10118_ & new_n4286_;
  assign new_n5524_ = new_n10118_ & new_n4288_;
  assign new_n5525_ = new_n5524_ | new_n5523_;
  assign new_n5526_ = new_n10120_ & new_n4295_;
  assign new_n5527_ = new_n10120_ & new_n4297_;
  assign new_n5528_ = new_n5527_ | new_n5526_;
  assign new_n5529_ = new_n10122_ & new_n4304_;
  assign new_n5530_ = new_n10122_ & new_n4306_;
  assign new_n5531_ = new_n5530_ | new_n5529_;
  assign new_n5532_ = new_n10124_ & new_n4313_;
  assign new_n5533_ = new_n10124_ & new_n4335_;
  assign new_n5534_ = new_n5533_ | new_n5532_;
  assign new_n5535_ = new_n9880_ & new_n9876_;
  assign new_n5536_ = new_n9881_ | new_n9878_;
  assign new_n5537_ = new_n5536_ & new_n10125_;
  assign new_n5538_ = new_n5535_ | new_n9882_;
  assign new_n5539_ = new_n9080_ & new_n9873_;
  assign new_n5540_ = new_n9095_ | new_n9875_;
  assign new_n5541_ = new_n9051_ & new_n10127_;
  assign new_n5542_ = new_n9068_ | new_n10129_;
  assign new_n5543_ = new_n10130_ & new_n10131_;
  assign new_n5544_ = new_n10132_ | new_n10133_;
  assign new_n5545_ = new_n10134_ & new_n10131_;
  assign new_n5546_ = new_n10135_ | new_n10133_;
  assign new_n5547_ = new_n10136_ | new_n5537_;
  assign new_n5548_ = new_n9965_ & new_n9961_;
  assign new_n5549_ = new_n9967_ | new_n9963_;
  assign new_n5550_ = new_n9964_ & new_n9960_;
  assign new_n5551_ = new_n9966_ | new_n9962_;
  assign new_n5552_ = new_n5551_ & new_n5549_;
  assign new_n5553_ = new_n5550_ | new_n5548_;
  assign new_n5554_ = new_n9948_ & new_n9944_;
  assign new_n5555_ = new_n9949_ | new_n9946_;
  assign new_n5556_ = new_n5555_ & new_n9950_;
  assign new_n5557_ = new_n5554_ | new_n9953_;
  assign new_n5558_ = new_n9080_ & new_n9940_;
  assign new_n5559_ = new_n9095_ | new_n9943_;
  assign new_n5560_ = new_n9054_ & new_n10139_;
  assign new_n5561_ = new_n9068_ | new_n10142_;
  assign new_n5562_ = new_n10143_ & new_n10144_;
  assign new_n5563_ = new_n10145_ | new_n10146_;
  assign new_n5564_ = new_n10147_ & new_n10144_;
  assign new_n5565_ = new_n10148_ | new_n10146_;
  assign new_n5566_ = new_n10150_ & new_n10151_;
  assign new_n5567_ = new_n10153_ | new_n10154_;
  assign new_n5568_ = new_n10156_ & new_n10151_;
  assign new_n5569_ = new_n10158_ | new_n10154_;
  assign new_n5570_ = new_n10156_ & new_n10150_;
  assign new_n5571_ = new_n10158_ | new_n10153_;
  assign new_n5572_ = new_n5571_ & new_n5569_;
  assign new_n5573_ = new_n5570_ | new_n5568_;
  assign new_n5574_ = new_n9022_ & new_n10139_;
  assign new_n5575_ = new_n9037_ | new_n10142_;
  assign new_n5576_ = new_n10159_ & new_n10160_;
  assign new_n5577_ = new_n10161_ | new_n10162_;
  assign new_n5578_ = new_n10164_ & new_n10155_;
  assign new_n5579_ = new_n10166_ | new_n10157_;
  assign new_n5580_ = new_n5578_ | new_n5552_;
  assign new_n5581_ = new_n10116_ | new_n10114_;
  assign new_n5582_ = new_n10115_ | new_n10113_;
  assign new_n5583_ = new_n5582_ & new_n5581_;
  assign new_n5584_ = new_n10104_ & new_n10102_;
  assign new_n5585_ = new_n10103_ & new_n10101_;
  assign new_n5586_ = new_n5585_ | new_n5584_;
  assign new_n5587_ = new_n10168_ & new_n4407_;
  assign new_n5588_ = new_n10168_ & new_n4409_;
  assign new_n5589_ = new_n5588_ | new_n5587_;
  assign new_n5590_ = new_n10170_ & new_n4580_;
  assign new_n5591_ = new_n10170_ & new_n4662_;
  assign new_n5592_ = new_n5591_ | new_n5590_;
  assign new_n5593_ = new_n10172_ & new_n4797_;
  assign new_n5594_ = new_n10172_ & new_n4881_;
  assign new_n5595_ = new_n5594_ | new_n5593_;
  assign new_n5596_ = new_n9083_ & new_n10174_;
  assign new_n5597_ = new_n9098_ | new_n10175_;
  assign new_n5598_ = new_n8795_ & new_n8906_;
  assign new_n5599_ = new_n9174_ & new_n10176_;
  assign new_n5600_ = new_n7707_ & new_n9559_;
  assign new_n5601_ = new_n10062_ | new_n9943_;
  assign new_n5602_ = new_n9037_ | new_n9874_;
  assign new_n5603_ = new_n10076_ & new_n10069_;
  assign new_n5604_ = new_n10090_ & new_n10083_;
  assign new_n5605_ = new_n10023_ & new_n10019_;
  assign new_n5606_ = new_n10025_ | new_n10021_;
  assign new_n5607_ = new_n10022_ & new_n10018_;
  assign new_n5608_ = new_n10024_ | new_n10020_;
  assign new_n5609_ = new_n5608_ & new_n5606_;
  assign new_n5610_ = new_n5607_ | new_n5605_;
  assign new_n5611_ = new_n9354_ & new_n9346_;
  assign new_n5612_ = new_n9356_ | new_n9348_;
  assign new_n5613_ = new_n10177_ & new_n10178_;
  assign new_n5614_ = new_n10179_ | new_n10180_;
  assign new_n5615_ = new_n10182_ & new_n10178_;
  assign new_n5616_ = new_n10183_ | new_n10180_;
  assign new_n5617_ = new_n10182_ & new_n10177_;
  assign new_n5618_ = new_n10183_ | new_n10179_;
  assign new_n5619_ = new_n5618_ & new_n5616_;
  assign new_n5620_ = new_n5617_ | new_n5615_;
  assign new_n5621_ = new_n9297_ & new_n9560_;
  assign new_n5622_ = new_n9301_ | new_n9569_;
  assign new_n5623_ = new_n5621_ | new_n5619_;
  assign new_n5624_ = new_n10185_ & new_n10181_;
  assign new_n5625_ = new_n9083_ & new_n10187_;
  assign new_n5626_ = new_n9098_ | new_n10188_;
  assign new_n5627_ = new_n9054_ & new_n10174_;
  assign new_n5628_ = new_n9069_ | new_n10175_;
  assign new_n5629_ = new_n5628_ & new_n5625_;
  assign new_n5630_ = new_n10189_ | new_n5626_;
  assign new_n5631_ = new_n9084_ & new_n10138_;
  assign new_n5632_ = new_n9099_ | new_n10141_;
  assign new_n5633_ = new_n9055_ & new_n10191_;
  assign new_n5634_ = new_n9069_ | new_n10194_;
  assign new_n5635_ = new_n10195_ & new_n10196_;
  assign new_n5636_ = new_n10197_ | new_n10198_;
  assign new_n5637_ = new_n10199_ & new_n10196_;
  assign new_n5638_ = new_n10200_ | new_n10198_;
  assign new_n5639_ = new_n10199_ & new_n10195_;
  assign new_n5640_ = new_n10200_ | new_n10197_;
  assign new_n5641_ = new_n5640_ & new_n10202_;
  assign new_n5642_ = new_n5639_ | new_n10204_;
  assign new_n5643_ = new_n9084_ & new_n10191_;
  assign new_n5644_ = new_n9099_ | new_n10194_;
  assign new_n5645_ = new_n9055_ & new_n9853_;
  assign new_n5646_ = new_n9071_ | new_n9856_;
  assign new_n5647_ = new_n10205_ & new_n10206_;
  assign new_n5648_ = new_n10207_ | new_n10208_;
  assign new_n5649_ = new_n10209_ & new_n10206_;
  assign new_n5650_ = new_n10210_ | new_n10208_;
  assign new_n5651_ = new_n10212_ & new_n10213_;
  assign new_n5652_ = new_n10215_ | new_n10216_;
  assign new_n5653_ = new_n10218_ & new_n10213_;
  assign new_n5654_ = new_n10219_ | new_n10216_;
  assign new_n5655_ = new_n10218_ & new_n10212_;
  assign new_n5656_ = new_n10219_ | new_n10215_;
  assign new_n5657_ = new_n5656_ & new_n5654_;
  assign new_n5658_ = new_n5655_ | new_n5653_;
  assign new_n5659_ = new_n9022_ & new_n9854_;
  assign new_n5660_ = new_n9038_ | new_n9855_;
  assign new_n5661_ = new_n5659_ | new_n5657_;
  assign new_n5662_ = new_n10221_ & new_n10217_;
  assign new_n5663_ = new_n9086_ & new_n9105_;
  assign new_n5664_ = new_n9101_ | new_n9108_;
  assign new_n5665_ = new_n9057_ & new_n10224_;
  assign new_n5666_ = new_n9071_ | new_n10227_;
  assign new_n5667_ = new_n10229_ & new_n10230_;
  assign new_n5668_ = new_n10231_ | new_n10232_;
  assign new_n5669_ = new_n10233_ & new_n10230_;
  assign new_n5670_ = new_n10234_ | new_n10232_;
  assign new_n5671_ = new_n10233_ & new_n10229_;
  assign new_n5672_ = new_n10234_ | new_n10231_;
  assign new_n5673_ = new_n5672_ & new_n10236_;
  assign new_n5674_ = new_n5671_ | new_n10238_;
  assign new_n5675_ = new_n9086_ & new_n10224_;
  assign new_n5676_ = new_n9101_ | new_n10227_;
  assign new_n5677_ = new_n9057_ & new_n9885_;
  assign new_n5678_ = new_n9072_ | new_n9888_;
  assign new_n5679_ = new_n10239_ & new_n10240_;
  assign new_n5680_ = new_n10241_ | new_n10242_;
  assign new_n5681_ = new_n10243_ & new_n10240_;
  assign new_n5682_ = new_n10244_ | new_n10242_;
  assign new_n5683_ = new_n10246_ & new_n10247_;
  assign new_n5684_ = new_n10249_ | new_n10250_;
  assign new_n5685_ = new_n10252_ & new_n10247_;
  assign new_n5686_ = new_n10254_ | new_n10250_;
  assign new_n5687_ = new_n10252_ & new_n10246_;
  assign new_n5688_ = new_n10254_ | new_n10249_;
  assign new_n5689_ = new_n5688_ & new_n5686_;
  assign new_n5690_ = new_n5687_ | new_n5685_;
  assign new_n5691_ = new_n9023_ & new_n9884_;
  assign new_n5692_ = new_n9038_ | new_n9889_;
  assign new_n5693_ = new_n10255_ & new_n10256_;
  assign new_n5694_ = new_n10257_ | new_n10258_;
  assign new_n5695_ = new_n10260_ & new_n10256_;
  assign new_n5696_ = new_n10262_ | new_n10258_;
  assign new_n5697_ = new_n10260_ & new_n10255_;
  assign new_n5698_ = new_n10262_ | new_n10257_;
  assign new_n5699_ = new_n5698_ & new_n5696_;
  assign new_n5700_ = new_n5697_ | new_n5695_;
  assign new_n5701_ = new_n10243_ & new_n10239_;
  assign new_n5702_ = new_n10244_ | new_n10241_;
  assign new_n5703_ = new_n5702_ & new_n10245_;
  assign new_n5704_ = new_n5701_ | new_n10248_;
  assign new_n5705_ = new_n10263_ & new_n9904_;
  assign new_n5706_ = new_n10264_ | new_n9906_;
  assign new_n5707_ = new_n10266_ & new_n10263_;
  assign new_n5708_ = new_n10268_ | new_n10264_;
  assign new_n5709_ = new_n10266_ & new_n9903_;
  assign new_n5710_ = new_n10268_ | new_n9905_;
  assign new_n5711_ = new_n5710_ & new_n5708_;
  assign new_n5712_ = new_n5709_ | new_n5707_;
  assign new_n5713_ = new_n9023_ & new_n9891_;
  assign new_n5714_ = new_n9040_ | new_n9896_;
  assign new_n5715_ = new_n10269_ & new_n10270_;
  assign new_n5716_ = new_n10271_ | new_n10272_;
  assign new_n5717_ = new_n10274_ & new_n10265_;
  assign new_n5718_ = new_n10276_ | new_n10267_;
  assign new_n5719_ = new_n10277_ & new_n10278_;
  assign new_n5720_ = new_n10279_ | new_n10280_;
  assign new_n5721_ = new_n10282_ & new_n10278_;
  assign new_n5722_ = new_n10283_ | new_n10280_;
  assign new_n5723_ = new_n10282_ & new_n10277_;
  assign new_n5724_ = new_n10283_ | new_n10279_;
  assign new_n5725_ = new_n5724_ & new_n5722_;
  assign new_n5726_ = new_n5723_ | new_n5721_;
  assign new_n5727_ = new_n10056_ & new_n9893_;
  assign new_n5728_ = new_n10063_ | new_n9896_;
  assign new_n5729_ = new_n5727_ | new_n5725_;
  assign new_n5730_ = new_n10285_ & new_n10281_;
  assign new_n5731_ = new_n10185_ & new_n5622_;
  assign new_n5732_ = new_n10287_ & new_n5434_;
  assign new_n5733_ = new_n10289_ & new_n5463_;
  assign new_n5734_ = new_n10291_ & new_n5492_;
  assign new_n5735_ = new_n10293_ & new_n5521_;
  assign new_n5736_ = new_n10287_ & new_n5432_;
  assign new_n5737_ = new_n10289_ & new_n5461_;
  assign new_n5738_ = new_n10293_ & new_n5499_;
  assign new_n5739_ = new_n10291_ & new_n5470_;
  assign new_n5740_ = new_n10184_ & new_n5620_;
  assign new_n5741_ = new_n10294_ & new_n10295_;
  assign new_n5742_ = new_n10296_ & new_n10297_;
  assign new_n5743_ = new_n10298_ & new_n10299_;
  assign new_n5744_ = new_n10300_ & new_n10301_;
  assign new_n5745_ = new_n10302_ & new_n10303_;
  assign new_n5746_ = new_n10304_ | new_n10305_;
  assign new_n5747_ = new_n10134_ & new_n10130_;
  assign new_n5748_ = new_n10135_ | new_n10132_;
  assign new_n5749_ = new_n5748_ & new_n10306_;
  assign new_n5750_ = new_n5747_ | new_n10136_;
  assign new_n5751_ = new_n9087_ & new_n10127_;
  assign new_n5752_ = new_n9100_ | new_n10129_;
  assign new_n5753_ = new_n9056_ & new_n10187_;
  assign new_n5754_ = new_n9072_ | new_n10188_;
  assign new_n5755_ = new_n10307_ & new_n10308_;
  assign new_n5756_ = new_n5753_ | new_n10309_;
  assign new_n5757_ = new_n10310_ & new_n10308_;
  assign new_n5758_ = new_n5755_ | new_n10309_;
  assign new_n5759_ = new_n10311_ | new_n5749_;
  assign new_n5760_ = new_n10164_ & new_n10160_;
  assign new_n5761_ = new_n10166_ | new_n10162_;
  assign new_n5762_ = new_n10163_ & new_n10159_;
  assign new_n5763_ = new_n10165_ | new_n10161_;
  assign new_n5764_ = new_n5763_ & new_n5761_;
  assign new_n5765_ = new_n5762_ | new_n5760_;
  assign new_n5766_ = new_n10147_ & new_n10143_;
  assign new_n5767_ = new_n10148_ | new_n10145_;
  assign new_n5768_ = new_n5767_ & new_n10149_;
  assign new_n5769_ = new_n5766_ | new_n10152_;
  assign new_n5770_ = new_n10312_ & new_n10202_;
  assign new_n5771_ = new_n10313_ | new_n10204_;
  assign new_n5772_ = new_n10315_ & new_n10312_;
  assign new_n5773_ = new_n10317_ | new_n10313_;
  assign new_n5774_ = new_n10315_ & new_n10201_;
  assign new_n5775_ = new_n10317_ | new_n10203_;
  assign new_n5776_ = new_n5775_ & new_n5773_;
  assign new_n5777_ = new_n5774_ | new_n5772_;
  assign new_n5778_ = new_n9026_ & new_n10192_;
  assign new_n5779_ = new_n9040_ | new_n10193_;
  assign new_n5780_ = new_n5779_ & new_n5777_;
  assign new_n5781_ = new_n10318_ | new_n10319_;
  assign new_n5782_ = new_n5781_ & new_n10314_;
  assign new_n5783_ = new_n10321_ | new_n10316_;
  assign new_n5784_ = new_n5782_ | new_n5764_;
  assign new_n5785_ = new_n9130_ & new_n9126_;
  assign new_n5786_ = new_n9132_ | new_n9128_;
  assign new_n5787_ = new_n9129_ & new_n9125_;
  assign new_n5788_ = new_n9131_ | new_n9127_;
  assign new_n5789_ = new_n5788_ & new_n5786_;
  assign new_n5790_ = new_n5787_ | new_n5785_;
  assign new_n5791_ = new_n9113_ & new_n9109_;
  assign new_n5792_ = new_n9114_ | new_n9111_;
  assign new_n5793_ = new_n5792_ & new_n9115_;
  assign new_n5794_ = new_n5791_ | new_n9118_;
  assign new_n5795_ = new_n10322_ & new_n10236_;
  assign new_n5796_ = new_n10323_ | new_n10238_;
  assign new_n5797_ = new_n10325_ & new_n10322_;
  assign new_n5798_ = new_n10327_ | new_n10323_;
  assign new_n5799_ = new_n10325_ & new_n10235_;
  assign new_n5800_ = new_n10327_ | new_n10237_;
  assign new_n5801_ = new_n5800_ & new_n5798_;
  assign new_n5802_ = new_n5799_ | new_n5797_;
  assign new_n5803_ = new_n9026_ & new_n10223_;
  assign new_n5804_ = new_n9041_ | new_n10228_;
  assign new_n5805_ = new_n10328_ & new_n10329_;
  assign new_n5806_ = new_n10330_ | new_n10331_;
  assign new_n5807_ = new_n10333_ & new_n10324_;
  assign new_n5808_ = new_n10335_ | new_n10326_;
  assign new_n5809_ = new_n10336_ & new_n10337_;
  assign new_n5810_ = new_n10338_ | new_n10339_;
  assign new_n5811_ = new_n10341_ & new_n10337_;
  assign new_n5812_ = new_n10342_ | new_n10339_;
  assign new_n5813_ = new_n10341_ & new_n10336_;
  assign new_n5814_ = new_n10342_ | new_n10338_;
  assign new_n5815_ = new_n5814_ & new_n5812_;
  assign new_n5816_ = new_n5813_ | new_n5811_;
  assign new_n5817_ = new_n10057_ & new_n10225_;
  assign new_n5818_ = new_n10063_ | new_n10228_;
  assign new_n5819_ = new_n10343_ & new_n10344_;
  assign new_n5820_ = new_n10345_ | new_n10346_;
  assign new_n5821_ = new_n10348_ & new_n10344_;
  assign new_n5822_ = new_n10349_ | new_n10346_;
  assign new_n5823_ = new_n10348_ & new_n10343_;
  assign new_n5824_ = new_n10349_ | new_n10345_;
  assign new_n5825_ = new_n5824_ & new_n5822_;
  assign new_n5826_ = new_n5823_ | new_n5821_;
  assign new_n5827_ = new_n10333_ & new_n10329_;
  assign new_n5828_ = new_n10335_ | new_n10331_;
  assign new_n5829_ = new_n10332_ & new_n10328_;
  assign new_n5830_ = new_n10334_ | new_n10330_;
  assign new_n5831_ = new_n5830_ & new_n5828_;
  assign new_n5832_ = new_n5829_ | new_n5827_;
  assign new_n5833_ = new_n10259_ & new_n10251_;
  assign new_n5834_ = new_n10261_ | new_n10253_;
  assign new_n5835_ = new_n10350_ & new_n10351_;
  assign new_n5836_ = new_n10352_ | new_n10353_;
  assign new_n5837_ = new_n10355_ & new_n10351_;
  assign new_n5838_ = new_n10357_ | new_n10353_;
  assign new_n5839_ = new_n10355_ & new_n10350_;
  assign new_n5840_ = new_n10357_ | new_n10352_;
  assign new_n5841_ = new_n5840_ & new_n5838_;
  assign new_n5842_ = new_n5839_ | new_n5837_;
  assign new_n5843_ = new_n10057_ & new_n9886_;
  assign new_n5844_ = new_n10064_ | new_n9889_;
  assign new_n5845_ = new_n5844_ & new_n5842_;
  assign new_n5846_ = new_n10358_ | new_n10359_;
  assign new_n5847_ = new_n5846_ & new_n10354_;
  assign new_n5848_ = new_n10361_ | new_n10356_;
  assign new_n5849_ = new_n5847_ | new_n5825_;
  assign new_n5850_ = new_n10363_ & new_n5051_;
  assign new_n5851_ = new_n10363_ & new_n5053_;
  assign new_n5852_ = new_n5851_ | new_n5850_;
  assign new_n5853_ = new_n10034_ & new_n5383_;
  assign new_n5854_ = new_n10033_ & new_n5385_;
  assign new_n5855_ = new_n5854_ | new_n5853_;
  assign new_n5856_ = new_n10365_ & new_n5061_;
  assign new_n5857_ = new_n10365_ & new_n5103_;
  assign new_n5858_ = new_n5857_ | new_n5856_;
  assign new_n5859_ = new_n10367_ & new_n5110_;
  assign new_n5860_ = new_n10367_ & new_n5192_;
  assign new_n5861_ = new_n5860_ | new_n5859_;
  assign new_n5862_ = new_n10361_ | new_n10359_;
  assign new_n5863_ = new_n10360_ | new_n10358_;
  assign new_n5864_ = new_n5863_ & new_n5862_;
  assign new_n5865_ = new_n10310_ & new_n10307_;
  assign new_n5866_ = new_n5865_ | new_n10311_;
  assign new_n5867_ = new_n10321_ | new_n10319_;
  assign new_n5868_ = new_n10320_ | new_n10318_;
  assign new_n5869_ = new_n5868_ & new_n5867_;
  assign new_n5870_ = new_n10369_ & new_n5205_;
  assign new_n5871_ = new_n10369_ & new_n10125_;
  assign new_n5872_ = new_n5871_ | new_n5870_;
  assign new_n5873_ = new_n10371_ & new_n5252_;
  assign new_n5874_ = new_n10371_ & new_n5278_;
  assign new_n5875_ = new_n5874_ | new_n5873_;
  assign new_n5876_ = new_n10059_ & new_n10140_;
  assign new_n5877_ = new_n9025_ & new_n10128_;
  assign new_n5878_ = new_n10347_ & new_n10340_;
  assign new_n5879_ = new_n10372_ | new_n5597_;
  assign new_n5880_ = new_n10209_ & new_n10205_;
  assign new_n5881_ = new_n10210_ | new_n10207_;
  assign new_n5882_ = new_n5881_ & new_n10211_;
  assign new_n5883_ = new_n5880_ | new_n10214_;
  assign new_n5884_ = new_n10373_ & new_n9869_;
  assign new_n5885_ = new_n10374_ | new_n9871_;
  assign new_n5886_ = new_n10376_ & new_n10373_;
  assign new_n5887_ = new_n10377_ | new_n10374_;
  assign new_n5888_ = new_n10376_ & new_n9868_;
  assign new_n5889_ = new_n10377_ | new_n9870_;
  assign new_n5890_ = new_n5889_ & new_n5887_;
  assign new_n5891_ = new_n5888_ | new_n5886_;
  assign new_n5892_ = new_n9027_ & new_n9859_;
  assign new_n5893_ = new_n9041_ | new_n9860_;
  assign new_n5894_ = new_n5892_ | new_n5890_;
  assign new_n5895_ = new_n10379_ & new_n10375_;
  assign new_n5896_ = new_n10274_ & new_n10270_;
  assign new_n5897_ = new_n10276_ | new_n10272_;
  assign new_n5898_ = new_n10273_ & new_n10269_;
  assign new_n5899_ = new_n10275_ | new_n10271_;
  assign new_n5900_ = new_n5899_ & new_n5897_;
  assign new_n5901_ = new_n5898_ | new_n5896_;
  assign new_n5902_ = new_n9934_ & new_n9926_;
  assign new_n5903_ = new_n9936_ | new_n9928_;
  assign new_n5904_ = new_n10380_ & new_n10381_;
  assign new_n5905_ = new_n10382_ | new_n10383_;
  assign new_n5906_ = new_n10385_ & new_n10381_;
  assign new_n5907_ = new_n10386_ | new_n10383_;
  assign new_n5908_ = new_n10385_ & new_n10380_;
  assign new_n5909_ = new_n10386_ | new_n10382_;
  assign new_n5910_ = new_n5909_ & new_n5907_;
  assign new_n5911_ = new_n5908_ | new_n5906_;
  assign new_n5912_ = new_n10059_ & new_n9910_;
  assign new_n5913_ = new_n10064_ | new_n9913_;
  assign new_n5914_ = new_n5912_ | new_n5910_;
  assign new_n5915_ = new_n10388_ & new_n10384_;
  assign new_n5916_ = new_n10388_ & new_n5913_;
  assign new_n5917_ = new_n10379_ & new_n5893_;
  assign new_n5918_ = new_n10390_ & new_n5758_;
  assign new_n5919_ = new_n10392_ & new_n5783_;
  assign new_n5920_ = new_n10394_ & new_n5848_;
  assign new_n5921_ = new_n10394_ & new_n5826_;
  assign new_n5922_ = new_n10390_ & new_n5750_;
  assign new_n5923_ = new_n10392_ & new_n5765_;
  assign new_n5924_ = new_n10378_ & new_n5891_;
  assign new_n5925_ = new_n10387_ & new_n5911_;
  assign new_n5926_ = new_n10395_ & new_n10396_;
  assign new_n5927_ = new_n10397_ & new_n10398_;
  assign new_n5928_ = new_n10399_ & new_n10401_;
  assign new_n5929_ = new_n10402_ | new_n10403_;
  assign new_n5930_ = new_n10404_ | new_n10405_;
  assign new_n5931_ = new_n10407_ & new_n5407_;
  assign new_n5932_ = new_n10407_ & new_n5409_;
  assign new_n5933_ = new_n5932_ | new_n5931_;
  assign new_n5934_ = new_n10189_ | new_n5627_;
  assign new_n5935_ = new_n5934_ & new_n10401_;
  assign new_n5936_ = new_n10285_ & new_n5726_;
  assign new_n5937_ = new_n10284_ & new_n5728_;
  assign new_n5938_ = new_n5937_ | new_n5936_;
  assign new_n5939_ = new_n10221_ & new_n5658_;
  assign new_n5940_ = new_n10220_ & new_n5660_;
  assign new_n5941_ = new_n5940_ | new_n5939_;
  assign new_n5942_ = new_n10409_ & new_n5538_;
  assign new_n5943_ = new_n10409_ & new_n10306_;
  assign new_n5944_ = new_n5943_ | new_n5942_;
  assign new_n5945_ = new_n10411_ & new_n5553_;
  assign new_n5946_ = new_n10411_ & new_n5579_;
  assign new_n5947_ = new_n5946_ | new_n5945_;
  assign G6257 = new_n1617_;
  assign G6258 = new_n1620_;
  assign G6259 = new_n1623_;
  assign G6260 = new_n1626_;
  assign G6261 = new_n1629_;
  assign G6262 = new_n1632_;
  assign G6263 = new_n1635_;
  assign G6264 = new_n1638_;
  assign G6265 = new_n1641_;
  assign G6266 = new_n1644_;
  assign G6267 = new_n1647_;
  assign G6268 = new_n1650_;
  assign G6269 = new_n1653_;
  assign G6270 = new_n1656_;
  assign G6271 = new_n1659_;
  assign G6272 = new_n1662_;
  assign G6273 = new_n1664_;
  assign G6274 = new_n1667_;
  assign G6275 = new_n1670_;
  assign G6276 = new_n1679_;
  assign G6277 = new_n1694_;
  assign G6278 = new_n1717_;
  assign G6279 = new_n1746_;
  assign G6280 = new_n1781_;
  assign G6281 = new_n1824_;
  assign G6282 = new_n1873_;
  assign G6283 = new_n1928_;
  assign G6284 = new_n1991_;
  assign G6285 = new_n2050_;
  assign G6286 = new_n2089_;
  assign G6287 = new_n2105_;
  assign G6288 = ~new_n2108_;
  assign n2491_li = new_n6741_;
  assign n2575_li = new_n7417_;
  assign n2587_li = new_n7396_;
  assign n2599_li = new_n7355_;
  assign n2611_li = new_n7297_;
  assign n2623_li = new_n7268_;
  assign n2635_li = new_n7247_;
  assign n2647_li = new_n7206_;
  assign n2659_li = new_n7148_;
  assign n2671_li = new_n7136_;
  assign n2683_li = new_n999_;
  assign n2734_li = new_n851_;
  assign n2746_li = new_n853_;
  assign n2758_li = new_n855_;
  assign n2770_li = new_n857_;
  assign n2782_li = new_n859_;
  assign n2785_li = new_n903_;
  assign n2794_li = new_n861_;
  assign n2797_li = new_n907_;
  assign n2806_li = new_n863_;
  assign n2809_li = new_n911_;
  assign n2818_li = new_n865_;
  assign n2821_li = new_n915_;
  assign n2830_li = new_n867_;
  assign n2833_li = new_n919_;
  assign n2836_li = new_n921_;
  assign n2839_li = new_n6769_;
  assign n2842_li = new_n869_;
  assign n2845_li = new_n927_;
  assign n2848_li = new_n929_;
  assign n2851_li = new_n6813_;
  assign n2854_li = new_n871_;
  assign n2857_li = new_n935_;
  assign n2860_li = new_n937_;
  assign n2863_li = new_n6886_;
  assign n4871_i2 = new_n1043_;
  assign n4893_i2 = new_n1045_;
  assign n4938_i2 = new_n1047_;
  assign n5056_i2 = new_n1053_;
  assign n5100_i2 = new_n1057_;
  assign n5122_i2 = new_n1059_;
  assign n5254_i2 = new_n1061_;
  assign n5276_i2 = new_n1063_;
  assign n5316_i2 = new_n1065_;
  assign n5434_i2 = new_n1071_;
  assign n5473_i2 = new_n1075_;
  assign n5494_i2 = new_n1077_;
  assign n5620_i2 = new_n1079_;
  assign n5643_i2 = new_n1081_;
  assign n5682_i2 = new_n1083_;
  assign n5798_i2 = new_n1095_;
  assign n5839_i2 = new_n1099_;
  assign n5867_i2 = new_n1105_;
  assign n6052_i2 = new_n1117_;
  assign n6087_i2 = new_n1121_;
  assign n6153_i2 = new_n1125_;
  assign n6408_i2 = new_n1139_;
  assign n6454_i2 = new_n1143_;
  assign n6509_i2 = new_n1149_;
  assign n6775_i2 = new_n1161_;
  assign n6818_i2 = new_n1165_;
  assign n6892_i2 = new_n1167_;
  assign n5779_i2 = new_n7943_;
  assign n5780_i2 = new_n1091_;
  assign n7156_i2 = new_n1189_;
  assign n5792_i2 = new_n7956_;
  assign n7205_i2 = new_n1193_;
  assign n5842_i2 = new_n7985_;
  assign n5863_i2 = new_n8043_;
  assign n7263_i2 = new_n1199_;
  assign n5881_i2 = new_n8084_;
  assign n5930_i2 = new_n8105_;
  assign n5959_i2 = new_n8134_;
  assign n5981_i2 = new_n8192_;
  assign n6042_i2 = new_n8241_;
  assign n6075_i2 = new_n8255_;
  assign n6103_i2 = new_n8306_;
  assign n7610_i2 = new_n1257_;
  assign n6169_i2 = new_n8397_;
  assign n7665_i2 = new_n1261_;
  assign n6205_i2 = new_n8525_;
  assign n6239_i2 = new_n7632_;
  assign n7788_i2 = new_n1291_;
  assign n6309_i2 = new_n6971_;
  assign n6461_i2 = new_n6867_;
  assign n6476_i2 = new_n1147_;
  assign n6521_i2 = new_n1151_;
  assign n6545_i2 = new_n1153_;
  assign G578_i2 = new_n6756_;
  assign G5106_i2 = new_n6755_;
  assign n6713_i2 = new_n1157_;
  assign G5164_i2 = new_n6793_;
  assign n6771_i2 = new_n1159_;
  assign n6810_i2 = new_n1163_;
  assign n6973_i2 = new_n1169_;
  assign n6995_i2 = new_n1171_;
  assign n7053_i2 = new_n1181_;
  assign G581_i2 = new_n6803_;
  assign G5467_i2 = new_n6802_;
  assign n7231_i2 = new_n1197_;
  assign G5527_i2 = new_n6848_;
  assign n7277_i2 = new_n1201_;
  assign n7304_i2 = new_n1205_;
  assign n7530_i2 = new_n1233_;
  assign n7595_i2 = new_n1251_;
  assign n7653_i2 = new_n1259_;
  assign G584_i2 = new_n6858_;
  assign G5820_i2 = new_n6857_;
  assign n7148_i2 = new_n8795_;
  assign n7149_i2 = new_n1187_;
  assign n7224_i2 = new_n8808_;
  assign n7916_i2 = new_n1317_;
  assign G5868_i2 = new_n6930_;
  assign n7958_i2 = new_n1327_;
  assign n7280_i2 = new_n8829_;
  assign n7313_i2 = new_n8858_;
  assign n8056_i2 = new_n1389_;
  assign n7323_i2 = new_n8937_;
  assign n7398_i2 = new_n9441_;
  assign n7459_i2 = new_n9500_;
  assign n7501_i2 = new_n9597_;
  assign n7518_i2 = new_n9173_;
  assign G563_i2 = new_n6881_;
  assign n7606_i2 = new_n9195_;
  assign G3358_i2 = new_n6880_;
  assign n7675_i2 = new_n9236_;
  assign G3410_i2 = new_n6985_;
  assign n7722_i2 = new_n9297_;
  assign n7747_i2 = new_n9369_;
  assign n7835_i2 = new_n7706_;
  assign G587_i2 = new_n6966_;
  assign G6046_i2 = new_n6965_;
  assign n7909_i2 = new_n7107_;
  assign G566_i2 = new_n6995_;
  assign G6070_i2 = new_n7585_;
  assign G3698_i2 = new_n6994_;
  assign n8086_i2 = new_n6999_;
  assign n8093_i2 = new_n1409_;
  assign G3752_i2 = new_n7072_;
  assign n8156_i2 = new_n1481_;
  assign n8199_i2 = new_n1531_;
  assign n2800_lo_buf_i2 = new_n7603_;
  assign G548_i2 = new_n7047_;
  assign G1715_i2 = new_n7046_;
  assign G569_i2 = new_n7082_;
  assign G1761_i2 = new_n7120_;
  assign G4043_i2 = new_n7081_;
  assign G4101_i2 = new_n7661_;
  assign G551_i2 = new_n7590_;
  assign G2034_i2 = new_n7589_;
  assign G4743_i2 = new_n7936_;
  assign G5271_i2 = new_n7933_;
  assign G5790_i2 = new_n7930_;
  assign G6122_i2 = new_n7748_;
  assign G2082_i2 = new_n7736_;
  assign n2812_lo_buf_i2 = new_n8367_;
  assign n2668_lo_buf_i2 = new_n9030_;
  assign n2680_lo_buf_i2 = new_n9087_;
  assign G572_i2 = new_n7701_;
  assign G6125_i2 = new_n7747_;
  assign G4395_i2 = new_n7700_;
  assign n2656_lo_buf_i2 = new_n9105_;
  assign G554_i2 = new_n7746_;
  assign G4452_i2 = new_n8570_;
  assign G2358_i2 = new_n7745_;
  assign n2644_lo_buf_i2 = new_n10225_;
  assign G2410_i2 = new_n8502_;
  assign n2632_lo_buf_i2 = new_n9886_;
  assign n2620_lo_buf_i2 = new_n9893_;
  assign G6131_i2 = ~new_n7940_;
  assign G4693_i2 = new_n8622_;
  assign G5209_i2 = new_n8624_;
  assign G5741_i2 = new_n8626_;
  assign G6082_i2 = new_n8628_;
  assign G6119_i2 = new_n7939_;
  assign n2608_lo_buf_i2 = new_n9910_;
  assign n2596_lo_buf_i2 = new_n9940_;
  assign n2584_lo_buf_i2 = new_n10140_;
  assign n2572_lo_buf_i2 = new_n10192_;
  assign n2704_lo_buf_i2 = new_n9027_;
  assign G557_i2 = new_n8512_;
  assign G5936_i2 = ~new_n9708_;
  assign G5442_i2 = ~new_n9710_;
  assign G4926_i2 = ~new_n9712_;
  assign G6134_i2 = new_n8579_;
  assign G3929_i2 = new_n8985_;
  assign G4425_i2 = new_n8988_;
  assign G4947_i2 = new_n8991_;
  assign n2764_lo_buf_i2 = new_n9560_;
  assign G2689_i2 = new_n8511_;
  assign n2560_lo_buf_i2 = new_n9854_;
  assign n2824_lo_buf_i2 = new_n8996_;
  assign G575_i2 = new_n8631_;
  assign G2740_i2 = new_n9690_;
  assign G4749_i2 = new_n8630_;
  assign n2548_lo_buf_i2 = new_n9859_;
  assign n2536_lo_buf_i2 = new_n9872_;
  assign n2524_lo_buf_i2 = new_n10128_;
  assign G875_i2 = ~new_n9701_;
  assign G1064_i2 = ~new_n9703_;
  assign G1253_i2 = ~new_n9705_;
  assign G6140_i2 = ~new_n9707_;
  assign G5151_i2 = new_n9694_;
  assign G5686_i2 = new_n9696_;
  assign G6061_i2 = new_n9698_;
  assign G4803_i2 = new_n9704_;
  assign G5332_i2 = new_n9702_;
  assign G5844_i2 = new_n9700_;
  assign G6114_i2 = new_n9706_;
  assign G4806_i2 = new_n9742_;
  assign G3881_i2 = new_n9743_;
  assign G4370_i2 = new_n9745_;
  assign G4896_i2 = new_n9747_;
  assign G5001_i2 = new_n9749_;
  assign G3121_i2 = new_n9751_;
  assign n2512_lo_buf_i2 = new_n10186_;
  assign G4085_i2 = ~new_n10117_;
  assign G4605_i2 = ~new_n10119_;
  assign G5118_i2 = ~new_n10121_;
  assign G4997_i2 = new_n10123_;
  assign n2500_lo_buf_i2 = new_n10173_;
  assign n2716_lo_buf_i2 = new_n10058_;
  assign G560_i2 = ~new_n9755_;
  assign G1895_i2 = new_n10051_;
  assign G3064_i2 = new_n10167_;
  assign G3269_i2 = new_n10169_;
  assign G3569_i2 = new_n10171_;
  assign G3022_i2 = new_n9754_;
  assign G1196_i2 = ~new_n10044_;
  assign G1007_i2 = ~new_n10046_;
  assign G818_i2 = ~new_n10048_;
  assign G674_i2 = ~new_n10050_;
  assign G5041_i2 = new_n4940_;
  assign G5562_i2 = new_n4941_;
  assign G6005_i2 = new_n4942_;
  assign G5214_i2 = new_n4943_;
  assign G5746_i2 = new_n4944_;
  assign G6087_i2 = new_n4945_;
  assign G6086_i2 = new_n4946_;
  assign G5745_i2 = new_n4947_;
  assign G5213_i2 = new_n4948_;
  assign G5893_i2 = new_n4949_;
  assign G5391_i2 = new_n4950_;
  assign G4864_i2 = new_n4951_;
  assign G6143_i2 = new_n4952_;
  assign G6008_i2 = ~new_n4955_;
  assign G5565_i2 = ~new_n4958_;
  assign G5044_i2 = ~new_n4961_;
  assign G3813_i2 = new_n10035_;
  assign G4325_i2 = new_n10037_;
  assign G4834_i2 = new_n10039_;
  assign G4993_i2 = new_n10041_;
  assign G3989_i2 = new_n10043_;
  assign G4490_i2 = new_n10045_;
  assign G5011_i2 = new_n10047_;
  assign G5112_i2 = new_n10049_;
  assign n2776_lo_buf_i2 = new_n10176_;
  assign G3298_i2 = ~new_n10362_;
  assign G3073_i2 = new_n9977_;
  assign G3265_i2 = new_n10364_;
  assign G3624_i2 = new_n10366_;
  assign G1642_i2 = new_n10368_;
  assign G1980_i2 = new_n10370_;
  assign n2488_lo_buf_i2 = new_n809_;
  assign G626_i2 = new_n5280_;
  assign G1139_i2 = ~new_n10295_;
  assign G950_i2 = ~new_n10297_;
  assign G707_i2 = ~new_n10299_;
  assign G545_i2 = ~new_n10301_;
  assign G4217_i2 = new_n5285_;
  assign G4716_i2 = new_n5286_;
  assign G5244_i2 = new_n5306_;
  assign G3136_i2 = ~new_n10303_;
  assign G3499_i2 = new_n10305_;
  assign G3885_i2 = new_n5388_;
  assign G5243_i2 = ~new_n5389_;
  assign G3886_i2 = new_n5390_;
  assign G4375_i2 = new_n5391_;
  assign G4901_i2 = new_n5392_;
  assign G5054_i2 = new_n5393_;
  assign G4374_i2 = new_n5394_;
  assign G4900_i2 = new_n5395_;
  assign G5053_i2 = new_n5396_;
  assign G5242_i2 = new_n5397_;
  assign G4034_i2 = new_n5398_;
  assign G4556_i2 = new_n5399_;
  assign G5064_i2 = new_n5400_;
  assign G5172_i2 = new_n5401_;
  assign G2030_i2 = ~new_n10406_;
  assign G3016_i2 = new_n10286_;
  assign G3520_i2 = new_n10288_;
  assign G3261_i2 = new_n10290_;
  assign G3620_i2 = new_n10292_;
  assign G4220_i2 = ~new_n5525_;
  assign G4719_i2 = ~new_n5528_;
  assign G5247_i2 = ~new_n5531_;
  assign G5109_i2 = new_n5534_;
  assign G1638_i2 = new_n10408_;
  assign G1976_i2 = new_n10410_;
  assign G3560_i2 = new_n10304_;
  assign G3205_i2 = ~new_n10302_;
  assign G3193_i2 = new_n10294_;
  assign G3367_i2 = new_n10298_;
  assign G3670_i2 = new_n10296_;
  assign G1400_i2 = new_n10300_;
  assign G1280_i2 = new_n5598_;
  assign G902_i2 = new_n5599_;
  assign G659_i2 = new_n5600_;
  assign G983_i2 = ~new_n10396_;
  assign G740_i2 = ~new_n10398_;
  assign G2917_i2 = new_n5603_;
  assign G3391_i2 = new_n5604_;
  assign G3494_i2 = new_n5624_;
  assign G1512_i2 = ~new_n10400_;
  assign G1854_i2 = new_n10403_;
  assign G2203_i2 = new_n10405_;
  assign G3493_i2 = ~new_n5731_;
  assign G3069_i2 = new_n5732_;
  assign G3574_i2 = new_n5733_;
  assign G3319_i2 = new_n5734_;
  assign G3667_i2 = new_n5735_;
  assign G3068_i2 = new_n5736_;
  assign G3573_i2 = new_n5737_;
  assign G3666_i2 = new_n5738_;
  assign G3318_i2 = new_n5739_;
  assign G3492_i2 = new_n5740_;
  assign G3241_i2 = new_n5741_;
  assign G3722_i2 = new_n5742_;
  assign G3422_i2 = new_n5743_;
  assign G1445_i2 = new_n10372_;
  assign G3257_i2 = ~new_n5745_;
  assign G3616_i2 = new_n5746_;
  assign G1634_i2 = new_n10389_;
  assign G1972_i2 = new_n10391_;
  assign G2256_i2 = new_n10393_;
  assign G3394_i2 = ~new_n5852_;
  assign G3557_i2 = ~new_n5855_;
  assign G3364_i2 = new_n5858_;
  assign G3719_i2 = new_n5861_;
  assign G2253_i2 = new_n10404_;
  assign G1583_i2 = ~new_n10399_;
  assign G1917_i2 = new_n10402_;
  assign G1727_i2 = new_n10397_;
  assign G2061_i2 = new_n10395_;
  assign G935_i2 = new_n5876_;
  assign G692_i2 = new_n5877_;
  assign G2136_i2 = new_n5878_;
  assign G1507_i2 = ~new_n5879_;
  assign G1849_i2 = new_n5895_;
  assign G2198_i2 = new_n5915_;
  assign G2197_i2 = ~new_n5916_;
  assign G1848_i2 = ~new_n5917_;
  assign G1689_i2 = new_n5918_;
  assign G2016_i2 = new_n5919_;
  assign G2314_i2 = new_n5920_;
  assign G2313_i2 = new_n5921_;
  assign G1688_i2 = new_n5922_;
  assign G2015_i2 = new_n5923_;
  assign G1847_i2 = new_n5924_;
  assign G2196_i2 = new_n5925_;
  assign G2118_i2 = new_n5926_;
  assign G1777_i2 = new_n5927_;
  assign G1630_i2 = ~new_n5928_;
  assign G1968_i2 = new_n5929_;
  assign G2309_i2 = new_n5930_;
  assign G2139_i2 = ~new_n5933_;
  assign G1580_i2 = new_n5935_;
  assign G2250_i2 = ~new_n5938_;
  assign G1914_i2 = ~new_n5941_;
  assign G1724_i2 = new_n5944_;
  assign G2058_i2 = new_n5947_;
  assign n2728_lo_buf_i2 = new_n849_;
  assign new_n6352_ = new_n947_;
  assign new_n6353_ = new_n953_;
  assign new_n6354_ = new_n959_;
  assign new_n6355_ = new_n965_;
  assign new_n6356_ = new_n971_;
  assign new_n6357_ = new_n977_;
  assign new_n6358_ = new_n983_;
  assign new_n6359_ = new_n989_;
  assign new_n6360_ = new_n995_;
  assign new_n6361_ = new_n1011_;
  assign new_n6362_ = new_n1037_;
  assign new_n6363_ = new_n1055_;
  assign new_n6364_ = new_n1073_;
  assign new_n6365_ = new_n1097_;
  assign new_n6366_ = new_n1141_;
  assign new_n6367_ = new_n1191_;
  assign new_n6368_ = new_n1241_;
  assign new_n6369_ = new_n1361_;
  assign new_n6370_ = new_n6369_;
  assign new_n6371_ = new_n1673_;
  assign new_n6372_ = new_n1671_;
  assign new_n6373_ = new_n1675_;
  assign new_n6374_ = new_n6373_;
  assign new_n6375_ = new_n1364_;
  assign new_n6376_ = new_n1342_;
  assign new_n6377_ = new_n1363_;
  assign new_n6378_ = new_n1341_;
  assign new_n6379_ = new_n1681_;
  assign new_n6380_ = new_n6379_;
  assign new_n6381_ = new_n1680_;
  assign new_n6382_ = new_n6381_;
  assign new_n6383_ = new_n1688_;
  assign new_n6384_ = new_n1686_;
  assign new_n6385_ = new_n1690_;
  assign new_n6386_ = new_n6385_;
  assign new_n6387_ = new_n1356_;
  assign new_n6388_ = new_n6387_;
  assign new_n6389_ = new_n1355_;
  assign new_n6390_ = new_n6389_;
  assign new_n6391_ = new_n1702_;
  assign new_n6392_ = new_n1700_;
  assign new_n6393_ = new_n1701_;
  assign new_n6394_ = new_n1699_;
  assign new_n6395_ = new_n1704_;
  assign new_n6396_ = new_n6395_;
  assign new_n6397_ = new_n1703_;
  assign new_n6398_ = new_n6397_;
  assign new_n6399_ = new_n1711_;
  assign new_n6400_ = new_n1709_;
  assign new_n6401_ = new_n1713_;
  assign new_n6402_ = new_n6401_;
  assign new_n6403_ = new_n941_;
  assign new_n6404_ = new_n6403_;
  assign new_n6405_ = new_n6404_;
  assign new_n6406_ = new_n6405_;
  assign new_n6407_ = new_n6404_;
  assign new_n6408_ = new_n6403_;
  assign new_n6409_ = new_n6408_;
  assign new_n6410_ = new_n6408_;
  assign new_n6411_ = new_n942_;
  assign new_n6412_ = new_n6411_;
  assign new_n6413_ = new_n6412_;
  assign new_n6414_ = new_n6413_;
  assign new_n6415_ = new_n6412_;
  assign new_n6416_ = new_n6411_;
  assign new_n6417_ = new_n6416_;
  assign new_n6418_ = new_n6416_;
  assign new_n6419_ = new_n1721_;
  assign new_n6420_ = new_n1719_;
  assign new_n6421_ = new_n1720_;
  assign new_n6422_ = new_n1718_;
  assign new_n6423_ = new_n1723_;
  assign new_n6424_ = new_n6423_;
  assign new_n6425_ = new_n1722_;
  assign new_n6426_ = new_n6425_;
  assign new_n6427_ = new_n1731_;
  assign new_n6428_ = new_n1729_;
  assign new_n6429_ = new_n1730_;
  assign new_n6430_ = new_n1728_;
  assign new_n6431_ = new_n1733_;
  assign new_n6432_ = new_n6431_;
  assign new_n6433_ = new_n1732_;
  assign new_n6434_ = new_n6433_;
  assign new_n6435_ = new_n1740_;
  assign new_n6436_ = new_n1738_;
  assign new_n6437_ = new_n1742_;
  assign new_n6438_ = new_n6437_;
  assign new_n6439_ = new_n1366_;
  assign new_n6440_ = new_n1340_;
  assign new_n6441_ = new_n1365_;
  assign new_n6442_ = new_n1339_;
  assign new_n6443_ = new_n1748_;
  assign new_n6444_ = new_n6443_;
  assign new_n6445_ = new_n1747_;
  assign new_n6446_ = new_n6445_;
  assign new_n6447_ = new_n1756_;
  assign new_n6448_ = new_n1754_;
  assign new_n6449_ = new_n1755_;
  assign new_n6450_ = new_n1753_;
  assign new_n6451_ = new_n1758_;
  assign new_n6452_ = new_n6451_;
  assign new_n6453_ = new_n1757_;
  assign new_n6454_ = new_n6453_;
  assign new_n6455_ = new_n1766_;
  assign new_n6456_ = new_n1764_;
  assign new_n6457_ = new_n1765_;
  assign new_n6458_ = new_n1763_;
  assign new_n6459_ = new_n1768_;
  assign new_n6460_ = new_n6459_;
  assign new_n6461_ = new_n1767_;
  assign new_n6462_ = new_n6461_;
  assign new_n6463_ = new_n1775_;
  assign new_n6464_ = new_n1773_;
  assign new_n6465_ = new_n1777_;
  assign new_n6466_ = new_n6465_;
  assign new_n6467_ = new_n1358_;
  assign new_n6468_ = new_n6467_;
  assign new_n6469_ = new_n1357_;
  assign new_n6470_ = new_n6469_;
  assign new_n6471_ = new_n1789_;
  assign new_n6472_ = new_n1787_;
  assign new_n6473_ = new_n1788_;
  assign new_n6474_ = new_n1786_;
  assign new_n6475_ = new_n1791_;
  assign new_n6476_ = new_n6475_;
  assign new_n6477_ = new_n1790_;
  assign new_n6478_ = new_n6477_;
  assign new_n6479_ = new_n1799_;
  assign new_n6480_ = new_n1797_;
  assign new_n6481_ = new_n1798_;
  assign new_n6482_ = new_n1796_;
  assign new_n6483_ = new_n1801_;
  assign new_n6484_ = new_n6483_;
  assign new_n6485_ = new_n1800_;
  assign new_n6486_ = new_n6485_;
  assign new_n6487_ = new_n1809_;
  assign new_n6488_ = new_n1807_;
  assign new_n6489_ = new_n1808_;
  assign new_n6490_ = new_n1806_;
  assign new_n6491_ = new_n1811_;
  assign new_n6492_ = new_n6491_;
  assign new_n6493_ = new_n1810_;
  assign new_n6494_ = new_n6493_;
  assign new_n6495_ = new_n1818_;
  assign new_n6496_ = new_n1816_;
  assign new_n6497_ = new_n1820_;
  assign new_n6498_ = new_n6497_;
  assign new_n6499_ = new_n933_;
  assign new_n6500_ = new_n6499_;
  assign new_n6501_ = new_n6500_;
  assign new_n6502_ = new_n6499_;
  assign new_n6503_ = new_n883_;
  assign new_n6504_ = new_n934_;
  assign new_n6505_ = new_n6504_;
  assign new_n6506_ = new_n6505_;
  assign new_n6507_ = new_n6504_;
  assign new_n6508_ = new_n884_;
  assign new_n6509_ = new_n1828_;
  assign new_n6510_ = new_n1826_;
  assign new_n6511_ = new_n1827_;
  assign new_n6512_ = new_n1825_;
  assign new_n6513_ = new_n1830_;
  assign new_n6514_ = new_n6513_;
  assign new_n6515_ = new_n1829_;
  assign new_n6516_ = new_n6515_;
  assign new_n6517_ = new_n1838_;
  assign new_n6518_ = new_n1836_;
  assign new_n6519_ = new_n1837_;
  assign new_n6520_ = new_n1835_;
  assign new_n6521_ = new_n1840_;
  assign new_n6522_ = new_n6521_;
  assign new_n6523_ = new_n1839_;
  assign new_n6524_ = new_n6523_;
  assign new_n6525_ = new_n1848_;
  assign new_n6526_ = new_n1846_;
  assign new_n6527_ = new_n1847_;
  assign new_n6528_ = new_n1845_;
  assign new_n6529_ = new_n1850_;
  assign new_n6530_ = new_n6529_;
  assign new_n6531_ = new_n1849_;
  assign new_n6532_ = new_n6531_;
  assign new_n6533_ = new_n1858_;
  assign new_n6534_ = new_n1856_;
  assign new_n6535_ = new_n1857_;
  assign new_n6536_ = new_n1855_;
  assign new_n6537_ = new_n1860_;
  assign new_n6538_ = new_n6537_;
  assign new_n6539_ = new_n1859_;
  assign new_n6540_ = new_n6539_;
  assign new_n6541_ = new_n1867_;
  assign new_n6542_ = new_n1865_;
  assign new_n6543_ = new_n1869_;
  assign new_n6544_ = new_n6543_;
  assign new_n6545_ = new_n1368_;
  assign new_n6546_ = new_n1338_;
  assign new_n6547_ = new_n1367_;
  assign new_n6548_ = new_n1337_;
  assign new_n6549_ = new_n1875_;
  assign new_n6550_ = new_n6549_;
  assign new_n6551_ = new_n1874_;
  assign new_n6552_ = new_n6551_;
  assign new_n6553_ = new_n885_;
  assign new_n6554_ = new_n886_;
  assign new_n6555_ = new_n1883_;
  assign new_n6556_ = new_n1881_;
  assign new_n6557_ = new_n1882_;
  assign new_n6558_ = new_n1880_;
  assign new_n6559_ = new_n1885_;
  assign new_n6560_ = new_n6559_;
  assign new_n6561_ = new_n1884_;
  assign new_n6562_ = new_n6561_;
  assign new_n6563_ = new_n1893_;
  assign new_n6564_ = new_n1891_;
  assign new_n6565_ = new_n1892_;
  assign new_n6566_ = new_n1890_;
  assign new_n6567_ = new_n1895_;
  assign new_n6568_ = new_n6567_;
  assign new_n6569_ = new_n1894_;
  assign new_n6570_ = new_n6569_;
  assign new_n6571_ = new_n1903_;
  assign new_n6572_ = new_n1901_;
  assign new_n6573_ = new_n1902_;
  assign new_n6574_ = new_n1900_;
  assign new_n6575_ = new_n1905_;
  assign new_n6576_ = new_n6575_;
  assign new_n6577_ = new_n1904_;
  assign new_n6578_ = new_n6577_;
  assign new_n6579_ = new_n1913_;
  assign new_n6580_ = new_n1911_;
  assign new_n6581_ = new_n1912_;
  assign new_n6582_ = new_n1910_;
  assign new_n6583_ = new_n1915_;
  assign new_n6584_ = new_n6583_;
  assign new_n6585_ = new_n1914_;
  assign new_n6586_ = new_n6585_;
  assign new_n6587_ = new_n1922_;
  assign new_n6588_ = new_n1920_;
  assign new_n6589_ = new_n1924_;
  assign new_n6590_ = new_n6589_;
  assign new_n6591_ = new_n1360_;
  assign new_n6592_ = new_n6591_;
  assign new_n6593_ = new_n1359_;
  assign new_n6594_ = new_n6593_;
  assign new_n6595_ = new_n1936_;
  assign new_n6596_ = new_n1934_;
  assign new_n6597_ = new_n1935_;
  assign new_n6598_ = new_n1933_;
  assign new_n6599_ = new_n1938_;
  assign new_n6600_ = new_n6599_;
  assign new_n6601_ = new_n1937_;
  assign new_n6602_ = new_n6601_;
  assign new_n6603_ = new_n887_;
  assign new_n6604_ = new_n888_;
  assign new_n6605_ = new_n1946_;
  assign new_n6606_ = new_n1944_;
  assign new_n6607_ = new_n1945_;
  assign new_n6608_ = new_n1943_;
  assign new_n6609_ = new_n1948_;
  assign new_n6610_ = new_n6609_;
  assign new_n6611_ = new_n1947_;
  assign new_n6612_ = new_n6611_;
  assign new_n6613_ = new_n1956_;
  assign new_n6614_ = new_n1954_;
  assign new_n6615_ = new_n1955_;
  assign new_n6616_ = new_n1953_;
  assign new_n6617_ = new_n1958_;
  assign new_n6618_ = new_n6617_;
  assign new_n6619_ = new_n1957_;
  assign new_n6620_ = new_n6619_;
  assign new_n6621_ = new_n1966_;
  assign new_n6622_ = new_n1964_;
  assign new_n6623_ = new_n1965_;
  assign new_n6624_ = new_n1963_;
  assign new_n6625_ = new_n1968_;
  assign new_n6626_ = new_n6625_;
  assign new_n6627_ = new_n1967_;
  assign new_n6628_ = new_n6627_;
  assign new_n6629_ = new_n1976_;
  assign new_n6630_ = new_n1974_;
  assign new_n6631_ = new_n1975_;
  assign new_n6632_ = new_n1973_;
  assign new_n6633_ = new_n1978_;
  assign new_n6634_ = new_n6633_;
  assign new_n6635_ = new_n1977_;
  assign new_n6636_ = new_n6635_;
  assign new_n6637_ = new_n1985_;
  assign new_n6638_ = new_n1983_;
  assign new_n6639_ = new_n1987_;
  assign new_n6640_ = new_n6639_;
  assign new_n6641_ = new_n891_;
  assign new_n6642_ = new_n6641_;
  assign new_n6643_ = new_n892_;
  assign new_n6644_ = new_n6643_;
  assign new_n6645_ = new_n1995_;
  assign new_n6646_ = new_n1993_;
  assign new_n6647_ = new_n1994_;
  assign new_n6648_ = new_n1992_;
  assign new_n6649_ = new_n1997_;
  assign new_n6650_ = new_n6649_;
  assign new_n6651_ = new_n1996_;
  assign new_n6652_ = new_n6651_;
  assign new_n6653_ = new_n889_;
  assign new_n6654_ = new_n890_;
  assign new_n6655_ = new_n2005_;
  assign new_n6656_ = new_n2003_;
  assign new_n6657_ = new_n2004_;
  assign new_n6658_ = new_n2002_;
  assign new_n6659_ = new_n2007_;
  assign new_n6660_ = new_n6659_;
  assign new_n6661_ = new_n2006_;
  assign new_n6662_ = new_n6661_;
  assign new_n6663_ = new_n2015_;
  assign new_n6664_ = new_n2013_;
  assign new_n6665_ = new_n2014_;
  assign new_n6666_ = new_n2012_;
  assign new_n6667_ = new_n2017_;
  assign new_n6668_ = new_n6667_;
  assign new_n6669_ = new_n2016_;
  assign new_n6670_ = new_n6669_;
  assign new_n6671_ = new_n2025_;
  assign new_n6672_ = new_n2023_;
  assign new_n6673_ = new_n2024_;
  assign new_n6674_ = new_n2022_;
  assign new_n6675_ = new_n2027_;
  assign new_n6676_ = new_n6675_;
  assign new_n6677_ = new_n2026_;
  assign new_n6678_ = new_n6677_;
  assign new_n6679_ = new_n2035_;
  assign new_n6680_ = new_n2033_;
  assign new_n6681_ = new_n2034_;
  assign new_n6682_ = new_n2032_;
  assign new_n6683_ = new_n2037_;
  assign new_n6684_ = new_n6683_;
  assign new_n6685_ = new_n2036_;
  assign new_n6686_ = new_n6685_;
  assign new_n6687_ = new_n2044_;
  assign new_n6688_ = new_n2042_;
  assign new_n6689_ = new_n2046_;
  assign new_n6690_ = new_n6689_;
  assign new_n6691_ = new_n2054_;
  assign new_n6692_ = new_n2052_;
  assign new_n6693_ = new_n2053_;
  assign new_n6694_ = new_n2051_;
  assign new_n6695_ = new_n2056_;
  assign new_n6696_ = new_n6695_;
  assign new_n6697_ = new_n2055_;
  assign new_n6698_ = new_n6697_;
  assign new_n6699_ = new_n2064_;
  assign new_n6700_ = new_n2062_;
  assign new_n6701_ = new_n2063_;
  assign new_n6702_ = new_n2061_;
  assign new_n6703_ = new_n2066_;
  assign new_n6704_ = new_n6703_;
  assign new_n6705_ = new_n2065_;
  assign new_n6706_ = new_n6705_;
  assign new_n6707_ = new_n2074_;
  assign new_n6708_ = new_n2072_;
  assign new_n6709_ = new_n2073_;
  assign new_n6710_ = new_n2071_;
  assign new_n6711_ = new_n2076_;
  assign new_n6712_ = new_n6711_;
  assign new_n6713_ = new_n2075_;
  assign new_n6714_ = new_n6713_;
  assign new_n6715_ = new_n2083_;
  assign new_n6716_ = new_n2081_;
  assign new_n6717_ = new_n2085_;
  assign new_n6718_ = new_n6717_;
  assign new_n6719_ = new_n2093_;
  assign new_n6720_ = new_n2091_;
  assign new_n6721_ = new_n2092_;
  assign new_n6722_ = new_n2090_;
  assign new_n6723_ = new_n2095_;
  assign new_n6724_ = new_n6723_;
  assign new_n6725_ = new_n2094_;
  assign new_n6726_ = new_n2104_;
  assign new_n6727_ = new_n6726_;
  assign new_n6728_ = new_n1255_;
  assign new_n6729_ = new_n6728_;
  assign new_n6730_ = new_n6729_;
  assign new_n6731_ = new_n6730_;
  assign new_n6732_ = new_n6730_;
  assign new_n6733_ = new_n6729_;
  assign new_n6734_ = new_n6733_;
  assign new_n6735_ = new_n6728_;
  assign new_n6736_ = new_n6735_;
  assign new_n6737_ = new_n6735_;
  assign new_n6738_ = new_n1041_;
  assign new_n6739_ = new_n6738_;
  assign new_n6740_ = new_n6739_;
  assign new_n6741_ = new_n6738_;
  assign new_n6742_ = new_n1256_;
  assign new_n6743_ = new_n6742_;
  assign new_n6744_ = new_n6743_;
  assign new_n6745_ = new_n6744_;
  assign new_n6746_ = new_n6744_;
  assign new_n6747_ = new_n6743_;
  assign new_n6748_ = new_n6747_;
  assign new_n6749_ = new_n6742_;
  assign new_n6750_ = new_n6749_;
  assign new_n6751_ = new_n6749_;
  assign new_n6752_ = new_n1042_;
  assign new_n6753_ = new_n6752_;
  assign new_n6754_ = new_n6752_;
  assign new_n6755_ = new_n2112_;
  assign new_n6756_ = new_n2109_;
  assign new_n6757_ = new_n923_;
  assign new_n6758_ = new_n6757_;
  assign new_n6759_ = new_n6758_;
  assign new_n6760_ = new_n6759_;
  assign new_n6761_ = new_n6759_;
  assign new_n6762_ = new_n6758_;
  assign new_n6763_ = new_n6762_;
  assign new_n6764_ = new_n6762_;
  assign new_n6765_ = new_n6757_;
  assign new_n6766_ = new_n6765_;
  assign new_n6767_ = new_n6766_;
  assign new_n6768_ = new_n6766_;
  assign new_n6769_ = new_n6765_;
  assign new_n6770_ = new_n6769_;
  assign new_n6771_ = new_n924_;
  assign new_n6772_ = new_n6771_;
  assign new_n6773_ = new_n6772_;
  assign new_n6774_ = new_n6773_;
  assign new_n6775_ = new_n6773_;
  assign new_n6776_ = new_n6772_;
  assign new_n6777_ = new_n6776_;
  assign new_n6778_ = new_n6776_;
  assign new_n6779_ = new_n6771_;
  assign new_n6780_ = new_n6779_;
  assign new_n6781_ = new_n6780_;
  assign new_n6782_ = new_n6780_;
  assign new_n6783_ = new_n6779_;
  assign new_n6784_ = new_n6783_;
  assign new_n6785_ = new_n1465_;
  assign new_n6786_ = new_n1402_;
  assign new_n6787_ = new_n1466_;
  assign new_n6788_ = new_n1401_;
  assign new_n6789_ = new_n2118_;
  assign new_n6790_ = new_n6789_;
  assign new_n6791_ = new_n2117_;
  assign new_n6792_ = new_n6791_;
  assign new_n6793_ = new_n2113_;
  assign new_n6794_ = new_n2126_;
  assign new_n6795_ = new_n2124_;
  assign new_n6796_ = new_n2125_;
  assign new_n6797_ = new_n2123_;
  assign new_n6798_ = new_n2128_;
  assign new_n6799_ = new_n6798_;
  assign new_n6800_ = new_n2127_;
  assign new_n6801_ = new_n6800_;
  assign new_n6802_ = new_n2134_;
  assign new_n6803_ = new_n2115_;
  assign new_n6804_ = new_n931_;
  assign new_n6805_ = new_n6804_;
  assign new_n6806_ = new_n6805_;
  assign new_n6807_ = new_n6806_;
  assign new_n6808_ = new_n6806_;
  assign new_n6809_ = new_n6805_;
  assign new_n6810_ = new_n6809_;
  assign new_n6811_ = new_n6804_;
  assign new_n6812_ = new_n6811_;
  assign new_n6813_ = new_n6811_;
  assign new_n6814_ = new_n932_;
  assign new_n6815_ = new_n6814_;
  assign new_n6816_ = new_n6815_;
  assign new_n6817_ = new_n6816_;
  assign new_n6818_ = new_n6816_;
  assign new_n6819_ = new_n6815_;
  assign new_n6820_ = new_n6819_;
  assign new_n6821_ = new_n6814_;
  assign new_n6822_ = new_n6821_;
  assign new_n6823_ = new_n6821_;
  assign new_n6824_ = new_n1448_;
  assign new_n6825_ = new_n6824_;
  assign new_n6826_ = new_n1447_;
  assign new_n6827_ = new_n6826_;
  assign new_n6828_ = new_n2146_;
  assign new_n6829_ = new_n2144_;
  assign new_n6830_ = new_n2145_;
  assign new_n6831_ = new_n2143_;
  assign new_n6832_ = new_n2148_;
  assign new_n6833_ = new_n6832_;
  assign new_n6834_ = new_n2147_;
  assign new_n6835_ = new_n6834_;
  assign new_n6836_ = new_n1039_;
  assign new_n6837_ = new_n6836_;
  assign new_n6838_ = new_n1040_;
  assign new_n6839_ = new_n6838_;
  assign new_n6840_ = new_n2156_;
  assign new_n6841_ = new_n2154_;
  assign new_n6842_ = new_n2155_;
  assign new_n6843_ = new_n2153_;
  assign new_n6844_ = new_n2158_;
  assign new_n6845_ = new_n6844_;
  assign new_n6846_ = new_n2157_;
  assign new_n6847_ = new_n6846_;
  assign new_n6848_ = new_n2135_;
  assign new_n6849_ = new_n2166_;
  assign new_n6850_ = new_n2164_;
  assign new_n6851_ = new_n2165_;
  assign new_n6852_ = new_n2163_;
  assign new_n6853_ = new_n2168_;
  assign new_n6854_ = new_n6853_;
  assign new_n6855_ = new_n2167_;
  assign new_n6856_ = new_n6855_;
  assign new_n6857_ = new_n2174_;
  assign new_n6858_ = new_n2137_;
  assign new_n6859_ = new_n1249_;
  assign new_n6860_ = new_n6859_;
  assign new_n6861_ = new_n6860_;
  assign new_n6862_ = new_n6859_;
  assign new_n6863_ = new_n1145_;
  assign new_n6864_ = new_n6863_;
  assign new_n6865_ = new_n6864_;
  assign new_n6866_ = new_n6864_;
  assign new_n6867_ = new_n6863_;
  assign new_n6868_ = new_n1250_;
  assign new_n6869_ = new_n6868_;
  assign new_n6870_ = new_n6869_;
  assign new_n6871_ = new_n6868_;
  assign new_n6872_ = new_n1146_;
  assign new_n6873_ = new_n6872_;
  assign new_n6874_ = new_n6873_;
  assign new_n6875_ = new_n6872_;
  assign new_n6876_ = new_n1533_;
  assign new_n6877_ = new_n6876_;
  assign new_n6878_ = new_n1534_;
  assign new_n6879_ = new_n6878_;
  assign new_n6880_ = new_n2184_;
  assign new_n6881_ = new_n2177_;
  assign new_n6882_ = new_n939_;
  assign new_n6883_ = new_n6882_;
  assign new_n6884_ = new_n6883_;
  assign new_n6885_ = new_n6883_;
  assign new_n6886_ = new_n6882_;
  assign new_n6887_ = new_n6886_;
  assign new_n6888_ = new_n940_;
  assign new_n6889_ = new_n6888_;
  assign new_n6890_ = new_n6889_;
  assign new_n6891_ = new_n6889_;
  assign new_n6892_ = new_n6888_;
  assign new_n6893_ = new_n6892_;
  assign new_n6894_ = new_n2192_;
  assign new_n6895_ = new_n2190_;
  assign new_n6896_ = new_n2191_;
  assign new_n6897_ = new_n2189_;
  assign new_n6898_ = new_n2194_;
  assign new_n6899_ = new_n6898_;
  assign new_n6900_ = new_n2193_;
  assign new_n6901_ = new_n6900_;
  assign new_n6902_ = new_n1035_;
  assign new_n6903_ = new_n6902_;
  assign new_n6904_ = new_n1036_;
  assign new_n6905_ = new_n6904_;
  assign new_n6906_ = new_n2202_;
  assign new_n6907_ = new_n2200_;
  assign new_n6908_ = new_n2201_;
  assign new_n6909_ = new_n2199_;
  assign new_n6910_ = new_n2204_;
  assign new_n6911_ = new_n6910_;
  assign new_n6912_ = new_n2203_;
  assign new_n6913_ = new_n6912_;
  assign new_n6914_ = new_n2212_;
  assign new_n6915_ = new_n2210_;
  assign new_n6916_ = new_n2211_;
  assign new_n6917_ = new_n2209_;
  assign new_n6918_ = new_n2214_;
  assign new_n6919_ = new_n6918_;
  assign new_n6920_ = new_n2213_;
  assign new_n6921_ = new_n6920_;
  assign new_n6922_ = new_n2222_;
  assign new_n6923_ = new_n2220_;
  assign new_n6924_ = new_n2221_;
  assign new_n6925_ = new_n2219_;
  assign new_n6926_ = new_n2224_;
  assign new_n6927_ = new_n6926_;
  assign new_n6928_ = new_n2223_;
  assign new_n6929_ = new_n6928_;
  assign new_n6930_ = new_n2175_;
  assign new_n6931_ = new_n2232_;
  assign new_n6932_ = new_n2230_;
  assign new_n6933_ = new_n2231_;
  assign new_n6934_ = new_n2229_;
  assign new_n6935_ = new_n2234_;
  assign new_n6936_ = new_n6935_;
  assign new_n6937_ = new_n2233_;
  assign new_n6938_ = new_n6937_;
  assign new_n6939_ = new_n1385_;
  assign new_n6940_ = new_n6939_;
  assign new_n6941_ = new_n6940_;
  assign new_n6942_ = new_n6941_;
  assign new_n6943_ = new_n6941_;
  assign new_n6944_ = new_n6940_;
  assign new_n6945_ = new_n6944_;
  assign new_n6946_ = new_n6944_;
  assign new_n6947_ = new_n6939_;
  assign new_n6948_ = new_n6947_;
  assign new_n6949_ = new_n6948_;
  assign new_n6950_ = new_n6948_;
  assign new_n6951_ = new_n6947_;
  assign new_n6952_ = new_n1386_;
  assign new_n6953_ = new_n6952_;
  assign new_n6954_ = new_n6953_;
  assign new_n6955_ = new_n6954_;
  assign new_n6956_ = new_n6954_;
  assign new_n6957_ = new_n6953_;
  assign new_n6958_ = new_n6957_;
  assign new_n6959_ = new_n6957_;
  assign new_n6960_ = new_n6952_;
  assign new_n6961_ = new_n6960_;
  assign new_n6962_ = new_n6961_;
  assign new_n6963_ = new_n6961_;
  assign new_n6964_ = new_n6960_;
  assign new_n6965_ = new_n2240_;
  assign new_n6966_ = new_n2187_;
  assign new_n6967_ = new_n1137_;
  assign new_n6968_ = new_n6967_;
  assign new_n6969_ = new_n6968_;
  assign new_n6970_ = new_n6968_;
  assign new_n6971_ = new_n6967_;
  assign new_n6972_ = new_n6971_;
  assign new_n6973_ = new_n1138_;
  assign new_n6974_ = new_n6973_;
  assign new_n6975_ = new_n6974_;
  assign new_n6976_ = new_n6973_;
  assign new_n6977_ = new_n2248_;
  assign new_n6978_ = new_n2246_;
  assign new_n6979_ = new_n2247_;
  assign new_n6980_ = new_n2245_;
  assign new_n6981_ = new_n2250_;
  assign new_n6982_ = new_n6981_;
  assign new_n6983_ = new_n2249_;
  assign new_n6984_ = new_n6983_;
  assign new_n6985_ = new_n2185_;
  assign new_n6986_ = new_n2258_;
  assign new_n6987_ = new_n2256_;
  assign new_n6988_ = new_n2257_;
  assign new_n6989_ = new_n2255_;
  assign new_n6990_ = new_n2260_;
  assign new_n6991_ = new_n6990_;
  assign new_n6992_ = new_n2259_;
  assign new_n6993_ = new_n6992_;
  assign new_n6994_ = new_n2266_;
  assign new_n6995_ = new_n2241_;
  assign new_n6996_ = new_n1399_;
  assign new_n6997_ = new_n6996_;
  assign new_n6998_ = new_n6997_;
  assign new_n6999_ = new_n6996_;
  assign new_n7000_ = new_n1231_;
  assign new_n7001_ = new_n7000_;
  assign new_n7002_ = new_n1400_;
  assign new_n7003_ = new_n7002_;
  assign new_n7004_ = new_n7003_;
  assign new_n7005_ = new_n7002_;
  assign new_n7006_ = new_n1232_;
  assign new_n7007_ = new_n7006_;
  assign new_n7008_ = new_n1606_;
  assign new_n7009_ = new_n1568_;
  assign new_n7010_ = new_n1605_;
  assign new_n7011_ = new_n1567_;
  assign new_n7012_ = new_n2272_;
  assign new_n7013_ = new_n7012_;
  assign new_n7014_ = new_n2271_;
  assign new_n7015_ = new_n7014_;
  assign new_n7016_ = new_n905_;
  assign new_n7017_ = new_n7016_;
  assign new_n7018_ = new_n7017_;
  assign new_n7019_ = new_n7018_;
  assign new_n7020_ = new_n7018_;
  assign new_n7021_ = new_n7017_;
  assign new_n7022_ = new_n7021_;
  assign new_n7023_ = new_n7021_;
  assign new_n7024_ = new_n7016_;
  assign new_n7025_ = new_n7024_;
  assign new_n7026_ = new_n7025_;
  assign new_n7027_ = new_n7025_;
  assign new_n7028_ = new_n7024_;
  assign new_n7029_ = new_n7028_;
  assign new_n7030_ = new_n7028_;
  assign new_n7031_ = new_n906_;
  assign new_n7032_ = new_n7031_;
  assign new_n7033_ = new_n7032_;
  assign new_n7034_ = new_n7033_;
  assign new_n7035_ = new_n7033_;
  assign new_n7036_ = new_n7032_;
  assign new_n7037_ = new_n7036_;
  assign new_n7038_ = new_n7036_;
  assign new_n7039_ = new_n7031_;
  assign new_n7040_ = new_n7039_;
  assign new_n7041_ = new_n7040_;
  assign new_n7042_ = new_n7040_;
  assign new_n7043_ = new_n7039_;
  assign new_n7044_ = new_n7043_;
  assign new_n7045_ = new_n7043_;
  assign new_n7046_ = new_n2278_;
  assign new_n7047_ = new_n2269_;
  assign new_n7048_ = new_n1547_;
  assign new_n7049_ = new_n1488_;
  assign new_n7050_ = new_n1548_;
  assign new_n7051_ = new_n1487_;
  assign new_n7052_ = new_n2284_;
  assign new_n7053_ = new_n7052_;
  assign new_n7054_ = new_n2283_;
  assign new_n7055_ = new_n7054_;
  assign new_n7056_ = new_n2292_;
  assign new_n7057_ = new_n2290_;
  assign new_n7058_ = new_n2291_;
  assign new_n7059_ = new_n2289_;
  assign new_n7060_ = new_n2294_;
  assign new_n7061_ = new_n7060_;
  assign new_n7062_ = new_n2293_;
  assign new_n7063_ = new_n7062_;
  assign new_n7064_ = new_n2302_;
  assign new_n7065_ = new_n2300_;
  assign new_n7066_ = new_n2301_;
  assign new_n7067_ = new_n2299_;
  assign new_n7068_ = new_n2304_;
  assign new_n7069_ = new_n7068_;
  assign new_n7070_ = new_n2303_;
  assign new_n7071_ = new_n7070_;
  assign new_n7072_ = new_n2267_;
  assign new_n7073_ = new_n2312_;
  assign new_n7074_ = new_n2310_;
  assign new_n7075_ = new_n2311_;
  assign new_n7076_ = new_n2309_;
  assign new_n7077_ = new_n2314_;
  assign new_n7078_ = new_n7077_;
  assign new_n7079_ = new_n2313_;
  assign new_n7080_ = new_n7079_;
  assign new_n7081_ = new_n2320_;
  assign new_n7082_ = new_n2279_;
  assign new_n7083_ = new_n1315_;
  assign new_n7084_ = new_n7083_;
  assign new_n7085_ = new_n7084_;
  assign new_n7086_ = new_n7085_;
  assign new_n7087_ = new_n7084_;
  assign new_n7088_ = new_n7083_;
  assign new_n7089_ = new_n7088_;
  assign new_n7090_ = new_n7088_;
  assign new_n7091_ = new_n1316_;
  assign new_n7092_ = new_n7091_;
  assign new_n7093_ = new_n7092_;
  assign new_n7094_ = new_n7093_;
  assign new_n7095_ = new_n7092_;
  assign new_n7096_ = new_n7091_;
  assign new_n7097_ = new_n7096_;
  assign new_n7098_ = new_n7096_;
  assign new_n7099_ = new_n1597_;
  assign new_n7100_ = new_n7099_;
  assign new_n7101_ = new_n1598_;
  assign new_n7102_ = new_n7101_;
  assign new_n7103_ = new_n1313_;
  assign new_n7104_ = new_n7103_;
  assign new_n7105_ = new_n7104_;
  assign new_n7106_ = new_n7104_;
  assign new_n7107_ = new_n7103_;
  assign new_n7108_ = new_n1314_;
  assign new_n7109_ = new_n7108_;
  assign new_n7110_ = new_n7109_;
  assign new_n7111_ = new_n7108_;
  assign new_n7112_ = new_n2332_;
  assign new_n7113_ = new_n2330_;
  assign new_n7114_ = new_n2331_;
  assign new_n7115_ = new_n2329_;
  assign new_n7116_ = new_n2334_;
  assign new_n7117_ = new_n7116_;
  assign new_n7118_ = new_n2333_;
  assign new_n7119_ = new_n7118_;
  assign new_n7120_ = new_n2281_;
  assign new_n7121_ = new_n2342_;
  assign new_n7122_ = new_n2340_;
  assign new_n7123_ = new_n2341_;
  assign new_n7124_ = new_n2339_;
  assign new_n7125_ = new_n2344_;
  assign new_n7126_ = new_n7125_;
  assign new_n7127_ = new_n2343_;
  assign new_n7128_ = new_n7127_;
  assign new_n7129_ = new_n1183_;
  assign new_n7130_ = new_n7129_;
  assign new_n7131_ = new_n7130_;
  assign new_n7132_ = new_n7130_;
  assign new_n7133_ = new_n7129_;
  assign new_n7134_ = new_n997_;
  assign new_n7135_ = new_n7134_;
  assign new_n7136_ = new_n7134_;
  assign new_n7137_ = new_n1184_;
  assign new_n7138_ = new_n7137_;
  assign new_n7139_ = new_n7138_;
  assign new_n7140_ = new_n7138_;
  assign new_n7141_ = new_n7137_;
  assign new_n7142_ = new_n998_;
  assign new_n7143_ = new_n7142_;
  assign new_n7144_ = new_n1155_;
  assign new_n7145_ = new_n1156_;
  assign new_n7146_ = new_n1003_;
  assign new_n7147_ = new_n7146_;
  assign new_n7148_ = new_n7146_;
  assign new_n7149_ = new_n1004_;
  assign new_n7150_ = new_n7149_;
  assign new_n7151_ = new_n7149_;
  assign new_n7152_ = new_n2358_;
  assign new_n7153_ = new_n2356_;
  assign new_n7154_ = new_n2357_;
  assign new_n7155_ = new_n2355_;
  assign new_n7156_ = new_n2360_;
  assign new_n7157_ = new_n7156_;
  assign new_n7158_ = new_n2359_;
  assign new_n7159_ = new_n7158_;
  assign new_n7160_ = new_n2362_;
  assign new_n7161_ = new_n2354_;
  assign new_n7162_ = new_n2361_;
  assign new_n7163_ = new_n2353_;
  assign new_n7164_ = new_n2364_;
  assign new_n7165_ = new_n7164_;
  assign new_n7166_ = new_n2363_;
  assign new_n7167_ = new_n7166_;
  assign new_n7168_ = new_n2372_;
  assign new_n7169_ = new_n2370_;
  assign new_n7170_ = new_n2371_;
  assign new_n7171_ = new_n2369_;
  assign new_n7172_ = new_n2374_;
  assign new_n7173_ = new_n7172_;
  assign new_n7174_ = new_n2373_;
  assign new_n7175_ = new_n7174_;
  assign new_n7176_ = new_n2376_;
  assign new_n7177_ = new_n2352_;
  assign new_n7178_ = new_n2375_;
  assign new_n7179_ = new_n2351_;
  assign new_n7180_ = new_n2378_;
  assign new_n7181_ = new_n7180_;
  assign new_n7182_ = new_n2377_;
  assign new_n7183_ = new_n7182_;
  assign new_n7184_ = new_n2386_;
  assign new_n7185_ = new_n2384_;
  assign new_n7186_ = new_n2385_;
  assign new_n7187_ = new_n2383_;
  assign new_n7188_ = new_n2388_;
  assign new_n7189_ = new_n7188_;
  assign new_n7190_ = new_n2387_;
  assign new_n7191_ = new_n7190_;
  assign new_n7192_ = new_n1442_;
  assign new_n7193_ = new_n7192_;
  assign new_n7194_ = new_n1441_;
  assign new_n7195_ = new_n7194_;
  assign new_n7196_ = new_n2408_;
  assign new_n7197_ = new_n2406_;
  assign new_n7198_ = new_n2407_;
  assign new_n7199_ = new_n2405_;
  assign new_n7200_ = new_n2410_;
  assign new_n7201_ = new_n7200_;
  assign new_n7202_ = new_n2409_;
  assign new_n7203_ = new_n7202_;
  assign new_n7204_ = new_n1007_;
  assign new_n7205_ = new_n7204_;
  assign new_n7206_ = new_n7204_;
  assign new_n7207_ = new_n1008_;
  assign new_n7208_ = new_n7207_;
  assign new_n7209_ = new_n2418_;
  assign new_n7210_ = new_n2416_;
  assign new_n7211_ = new_n2417_;
  assign new_n7212_ = new_n2415_;
  assign new_n7213_ = new_n2420_;
  assign new_n7214_ = new_n7213_;
  assign new_n7215_ = new_n2419_;
  assign new_n7216_ = new_n7215_;
  assign new_n7217_ = new_n2422_;
  assign new_n7218_ = new_n2400_;
  assign new_n7219_ = new_n2421_;
  assign new_n7220_ = new_n2399_;
  assign new_n7221_ = new_n2424_;
  assign new_n7222_ = new_n7221_;
  assign new_n7223_ = new_n2423_;
  assign new_n7224_ = new_n7223_;
  assign new_n7225_ = new_n2432_;
  assign new_n7226_ = new_n2430_;
  assign new_n7227_ = new_n2431_;
  assign new_n7228_ = new_n2429_;
  assign new_n7229_ = new_n2434_;
  assign new_n7230_ = new_n7229_;
  assign new_n7231_ = new_n2433_;
  assign new_n7232_ = new_n7231_;
  assign new_n7233_ = new_n2436_;
  assign new_n7234_ = new_n2394_;
  assign new_n7235_ = new_n2435_;
  assign new_n7236_ = new_n2393_;
  assign new_n7237_ = new_n2446_;
  assign new_n7238_ = new_n2444_;
  assign new_n7239_ = new_n2445_;
  assign new_n7240_ = new_n2443_;
  assign new_n7241_ = new_n2448_;
  assign new_n7242_ = new_n7241_;
  assign new_n7243_ = new_n2447_;
  assign new_n7244_ = new_n7243_;
  assign new_n7245_ = new_n1009_;
  assign new_n7246_ = new_n7245_;
  assign new_n7247_ = new_n7245_;
  assign new_n7248_ = new_n1010_;
  assign new_n7249_ = new_n7248_;
  assign new_n7250_ = new_n2456_;
  assign new_n7251_ = new_n2454_;
  assign new_n7252_ = new_n2455_;
  assign new_n7253_ = new_n2453_;
  assign new_n7254_ = new_n2458_;
  assign new_n7255_ = new_n7254_;
  assign new_n7256_ = new_n2457_;
  assign new_n7257_ = new_n7256_;
  assign new_n7258_ = new_n1460_;
  assign new_n7259_ = new_n1412_;
  assign new_n7260_ = new_n1459_;
  assign new_n7261_ = new_n1411_;
  assign new_n7262_ = new_n2466_;
  assign new_n7263_ = new_n7262_;
  assign new_n7264_ = new_n2465_;
  assign new_n7265_ = new_n7264_;
  assign new_n7266_ = new_n1013_;
  assign new_n7267_ = new_n7266_;
  assign new_n7268_ = new_n7266_;
  assign new_n7269_ = new_n1014_;
  assign new_n7270_ = new_n7269_;
  assign new_n7271_ = new_n2474_;
  assign new_n7272_ = new_n2472_;
  assign new_n7273_ = new_n2473_;
  assign new_n7274_ = new_n2471_;
  assign new_n7275_ = new_n2476_;
  assign new_n7276_ = new_n7275_;
  assign new_n7277_ = new_n2475_;
  assign new_n7278_ = new_n7277_;
  assign new_n7279_ = new_n2478_;
  assign new_n7280_ = new_n2464_;
  assign new_n7281_ = new_n2477_;
  assign new_n7282_ = new_n2463_;
  assign new_n7283_ = new_n2480_;
  assign new_n7284_ = new_n7283_;
  assign new_n7285_ = new_n2479_;
  assign new_n7286_ = new_n7285_;
  assign new_n7287_ = new_n2488_;
  assign new_n7288_ = new_n2486_;
  assign new_n7289_ = new_n2487_;
  assign new_n7290_ = new_n2485_;
  assign new_n7291_ = new_n2490_;
  assign new_n7292_ = new_n7291_;
  assign new_n7293_ = new_n2489_;
  assign new_n7294_ = new_n7293_;
  assign new_n7295_ = new_n1015_;
  assign new_n7296_ = new_n7295_;
  assign new_n7297_ = new_n7295_;
  assign new_n7298_ = new_n1016_;
  assign new_n7299_ = new_n7298_;
  assign new_n7300_ = new_n7298_;
  assign new_n7301_ = new_n2506_;
  assign new_n7302_ = new_n2504_;
  assign new_n7303_ = new_n2505_;
  assign new_n7304_ = new_n2503_;
  assign new_n7305_ = new_n2508_;
  assign new_n7306_ = new_n7305_;
  assign new_n7307_ = new_n2507_;
  assign new_n7308_ = new_n7307_;
  assign new_n7309_ = new_n2510_;
  assign new_n7310_ = new_n2502_;
  assign new_n7311_ = new_n2509_;
  assign new_n7312_ = new_n2501_;
  assign new_n7313_ = new_n2512_;
  assign new_n7314_ = new_n7313_;
  assign new_n7315_ = new_n2511_;
  assign new_n7316_ = new_n7315_;
  assign new_n7317_ = new_n2520_;
  assign new_n7318_ = new_n2518_;
  assign new_n7319_ = new_n2519_;
  assign new_n7320_ = new_n2517_;
  assign new_n7321_ = new_n2522_;
  assign new_n7322_ = new_n7321_;
  assign new_n7323_ = new_n2521_;
  assign new_n7324_ = new_n7323_;
  assign new_n7325_ = new_n2524_;
  assign new_n7326_ = new_n2496_;
  assign new_n7327_ = new_n2523_;
  assign new_n7328_ = new_n2495_;
  assign new_n7329_ = new_n2526_;
  assign new_n7330_ = new_n7329_;
  assign new_n7331_ = new_n2525_;
  assign new_n7332_ = new_n7331_;
  assign new_n7333_ = new_n2534_;
  assign new_n7334_ = new_n2532_;
  assign new_n7335_ = new_n2533_;
  assign new_n7336_ = new_n2531_;
  assign new_n7337_ = new_n2536_;
  assign new_n7338_ = new_n7337_;
  assign new_n7339_ = new_n2535_;
  assign new_n7340_ = new_n7339_;
  assign new_n7341_ = new_n1444_;
  assign new_n7342_ = new_n7341_;
  assign new_n7343_ = new_n1443_;
  assign new_n7344_ = new_n7343_;
  assign new_n7345_ = new_n2556_;
  assign new_n7346_ = new_n2554_;
  assign new_n7347_ = new_n2555_;
  assign new_n7348_ = new_n2553_;
  assign new_n7349_ = new_n2558_;
  assign new_n7350_ = new_n7349_;
  assign new_n7351_ = new_n2557_;
  assign new_n7352_ = new_n7351_;
  assign new_n7353_ = new_n1017_;
  assign new_n7354_ = new_n7353_;
  assign new_n7355_ = new_n7353_;
  assign new_n7356_ = new_n1018_;
  assign new_n7357_ = new_n7356_;
  assign new_n7358_ = new_n2566_;
  assign new_n7359_ = new_n2564_;
  assign new_n7360_ = new_n2565_;
  assign new_n7361_ = new_n2563_;
  assign new_n7362_ = new_n2568_;
  assign new_n7363_ = new_n7362_;
  assign new_n7364_ = new_n2567_;
  assign new_n7365_ = new_n7364_;
  assign new_n7366_ = new_n2570_;
  assign new_n7367_ = new_n2548_;
  assign new_n7368_ = new_n2569_;
  assign new_n7369_ = new_n2547_;
  assign new_n7370_ = new_n2572_;
  assign new_n7371_ = new_n7370_;
  assign new_n7372_ = new_n2571_;
  assign new_n7373_ = new_n7372_;
  assign new_n7374_ = new_n2580_;
  assign new_n7375_ = new_n2578_;
  assign new_n7376_ = new_n2579_;
  assign new_n7377_ = new_n2577_;
  assign new_n7378_ = new_n2582_;
  assign new_n7379_ = new_n7378_;
  assign new_n7380_ = new_n2581_;
  assign new_n7381_ = new_n7380_;
  assign new_n7382_ = new_n2584_;
  assign new_n7383_ = new_n2542_;
  assign new_n7384_ = new_n2583_;
  assign new_n7385_ = new_n2541_;
  assign new_n7386_ = new_n2594_;
  assign new_n7387_ = new_n2592_;
  assign new_n7388_ = new_n2593_;
  assign new_n7389_ = new_n2591_;
  assign new_n7390_ = new_n2596_;
  assign new_n7391_ = new_n7390_;
  assign new_n7392_ = new_n2595_;
  assign new_n7393_ = new_n7392_;
  assign new_n7394_ = new_n1019_;
  assign new_n7395_ = new_n7394_;
  assign new_n7396_ = new_n7394_;
  assign new_n7397_ = new_n1020_;
  assign new_n7398_ = new_n7397_;
  assign new_n7399_ = new_n2604_;
  assign new_n7400_ = new_n2602_;
  assign new_n7401_ = new_n2603_;
  assign new_n7402_ = new_n2601_;
  assign new_n7403_ = new_n2606_;
  assign new_n7404_ = new_n7403_;
  assign new_n7405_ = new_n2605_;
  assign new_n7406_ = new_n7405_;
  assign new_n7407_ = new_n1462_;
  assign new_n7408_ = new_n1414_;
  assign new_n7409_ = new_n1461_;
  assign new_n7410_ = new_n1413_;
  assign new_n7411_ = new_n2614_;
  assign new_n7412_ = new_n7411_;
  assign new_n7413_ = new_n2613_;
  assign new_n7414_ = new_n7413_;
  assign new_n7415_ = new_n1021_;
  assign new_n7416_ = new_n7415_;
  assign new_n7417_ = new_n7415_;
  assign new_n7418_ = new_n1022_;
  assign new_n7419_ = new_n7418_;
  assign new_n7420_ = new_n2622_;
  assign new_n7421_ = new_n2620_;
  assign new_n7422_ = new_n2621_;
  assign new_n7423_ = new_n2619_;
  assign new_n7424_ = new_n2624_;
  assign new_n7425_ = new_n7424_;
  assign new_n7426_ = new_n2623_;
  assign new_n7427_ = new_n7426_;
  assign new_n7428_ = new_n2626_;
  assign new_n7429_ = new_n2612_;
  assign new_n7430_ = new_n2625_;
  assign new_n7431_ = new_n2611_;
  assign new_n7432_ = new_n2628_;
  assign new_n7433_ = new_n7432_;
  assign new_n7434_ = new_n2627_;
  assign new_n7435_ = new_n7434_;
  assign new_n7436_ = new_n2636_;
  assign new_n7437_ = new_n2634_;
  assign new_n7438_ = new_n2635_;
  assign new_n7439_ = new_n2633_;
  assign new_n7440_ = new_n2638_;
  assign new_n7441_ = new_n7440_;
  assign new_n7442_ = new_n2637_;
  assign new_n7443_ = new_n7442_;
  assign new_n7444_ = new_n1023_;
  assign new_n7445_ = new_n7444_;
  assign new_n7446_ = new_n1024_;
  assign new_n7447_ = new_n7446_;
  assign new_n7448_ = new_n7446_;
  assign new_n7449_ = new_n2654_;
  assign new_n7450_ = new_n2652_;
  assign new_n7451_ = new_n2653_;
  assign new_n7452_ = new_n2651_;
  assign new_n7453_ = new_n2656_;
  assign new_n7454_ = new_n7453_;
  assign new_n7455_ = new_n2655_;
  assign new_n7456_ = new_n7455_;
  assign new_n7457_ = new_n2658_;
  assign new_n7458_ = new_n2650_;
  assign new_n7459_ = new_n2657_;
  assign new_n7460_ = new_n2649_;
  assign new_n7461_ = new_n2660_;
  assign new_n7462_ = new_n7461_;
  assign new_n7463_ = new_n2659_;
  assign new_n7464_ = new_n7463_;
  assign new_n7465_ = new_n2668_;
  assign new_n7466_ = new_n2666_;
  assign new_n7467_ = new_n2667_;
  assign new_n7468_ = new_n2665_;
  assign new_n7469_ = new_n2670_;
  assign new_n7470_ = new_n7469_;
  assign new_n7471_ = new_n2669_;
  assign new_n7472_ = new_n7471_;
  assign new_n7473_ = new_n2672_;
  assign new_n7474_ = new_n2644_;
  assign new_n7475_ = new_n2671_;
  assign new_n7476_ = new_n2643_;
  assign new_n7477_ = new_n2674_;
  assign new_n7478_ = new_n7477_;
  assign new_n7479_ = new_n2673_;
  assign new_n7480_ = new_n7479_;
  assign new_n7481_ = new_n2682_;
  assign new_n7482_ = new_n2680_;
  assign new_n7483_ = new_n2681_;
  assign new_n7484_ = new_n2679_;
  assign new_n7485_ = new_n2684_;
  assign new_n7486_ = new_n7485_;
  assign new_n7487_ = new_n2683_;
  assign new_n7488_ = new_n7487_;
  assign new_n7489_ = new_n1446_;
  assign new_n7490_ = new_n7489_;
  assign new_n7491_ = new_n1445_;
  assign new_n7492_ = new_n7491_;
  assign new_n7493_ = new_n2704_;
  assign new_n7494_ = new_n2702_;
  assign new_n7495_ = new_n2703_;
  assign new_n7496_ = new_n2701_;
  assign new_n7497_ = new_n2706_;
  assign new_n7498_ = new_n7497_;
  assign new_n7499_ = new_n2705_;
  assign new_n7500_ = new_n7499_;
  assign new_n7501_ = new_n1025_;
  assign new_n7502_ = new_n7501_;
  assign new_n7503_ = new_n1026_;
  assign new_n7504_ = new_n7503_;
  assign new_n7505_ = new_n2714_;
  assign new_n7506_ = new_n2712_;
  assign new_n7507_ = new_n2713_;
  assign new_n7508_ = new_n2711_;
  assign new_n7509_ = new_n2716_;
  assign new_n7510_ = new_n7509_;
  assign new_n7511_ = new_n2715_;
  assign new_n7512_ = new_n7511_;
  assign new_n7513_ = new_n2718_;
  assign new_n7514_ = new_n2696_;
  assign new_n7515_ = new_n2717_;
  assign new_n7516_ = new_n2695_;
  assign new_n7517_ = new_n2720_;
  assign new_n7518_ = new_n7517_;
  assign new_n7519_ = new_n2719_;
  assign new_n7520_ = new_n7519_;
  assign new_n7521_ = new_n2728_;
  assign new_n7522_ = new_n2726_;
  assign new_n7523_ = new_n2727_;
  assign new_n7524_ = new_n2725_;
  assign new_n7525_ = new_n2730_;
  assign new_n7526_ = new_n7525_;
  assign new_n7527_ = new_n2729_;
  assign new_n7528_ = new_n7527_;
  assign new_n7529_ = new_n2732_;
  assign new_n7530_ = new_n2690_;
  assign new_n7531_ = new_n2731_;
  assign new_n7532_ = new_n2689_;
  assign new_n7533_ = new_n1464_;
  assign new_n7534_ = new_n1416_;
  assign new_n7535_ = new_n1463_;
  assign new_n7536_ = new_n1415_;
  assign new_n7537_ = new_n2736_;
  assign new_n7538_ = new_n7537_;
  assign new_n7539_ = new_n2735_;
  assign new_n7540_ = new_n7539_;
  assign new_n7541_ = new_n1033_;
  assign new_n7542_ = new_n7541_;
  assign new_n7543_ = new_n1034_;
  assign new_n7544_ = new_n7543_;
  assign new_n7545_ = new_n2744_;
  assign new_n7546_ = new_n2742_;
  assign new_n7547_ = new_n2743_;
  assign new_n7548_ = new_n2741_;
  assign new_n7549_ = new_n2746_;
  assign new_n7550_ = new_n7549_;
  assign new_n7551_ = new_n2745_;
  assign new_n7552_ = new_n7551_;
  assign new_n7553_ = new_n2754_;
  assign new_n7554_ = new_n2752_;
  assign new_n7555_ = new_n2753_;
  assign new_n7556_ = new_n2751_;
  assign new_n7557_ = new_n2756_;
  assign new_n7558_ = new_n7557_;
  assign new_n7559_ = new_n2755_;
  assign new_n7560_ = new_n7559_;
  assign new_n7561_ = new_n2764_;
  assign new_n7562_ = new_n2762_;
  assign new_n7563_ = new_n2763_;
  assign new_n7564_ = new_n2761_;
  assign new_n7565_ = new_n2766_;
  assign new_n7566_ = new_n7565_;
  assign new_n7567_ = new_n2765_;
  assign new_n7568_ = new_n7567_;
  assign new_n7569_ = new_n2774_;
  assign new_n7570_ = new_n2772_;
  assign new_n7571_ = new_n2773_;
  assign new_n7572_ = new_n2771_;
  assign new_n7573_ = new_n2776_;
  assign new_n7574_ = new_n7573_;
  assign new_n7575_ = new_n2775_;
  assign new_n7576_ = new_n7575_;
  assign new_n7577_ = new_n2784_;
  assign new_n7578_ = new_n2782_;
  assign new_n7579_ = new_n2783_;
  assign new_n7580_ = new_n2781_;
  assign new_n7581_ = new_n2786_;
  assign new_n7582_ = new_n7581_;
  assign new_n7583_ = new_n2785_;
  assign new_n7584_ = new_n7583_;
  assign new_n7585_ = new_n2243_;
  assign new_n7586_ = new_n2794_;
  assign new_n7587_ = new_n2792_;
  assign new_n7588_ = new_n2796_;
  assign new_n7589_ = new_n2350_;
  assign new_n7590_ = new_n2323_;
  assign new_n7591_ = new_n909_;
  assign new_n7592_ = new_n7591_;
  assign new_n7593_ = new_n7592_;
  assign new_n7594_ = new_n7593_;
  assign new_n7595_ = new_n7593_;
  assign new_n7596_ = new_n7592_;
  assign new_n7597_ = new_n7596_;
  assign new_n7598_ = new_n7596_;
  assign new_n7599_ = new_n7591_;
  assign new_n7600_ = new_n7599_;
  assign new_n7601_ = new_n7600_;
  assign new_n7602_ = new_n7600_;
  assign new_n7603_ = new_n7599_;
  assign new_n7604_ = new_n910_;
  assign new_n7605_ = new_n7604_;
  assign new_n7606_ = new_n7605_;
  assign new_n7607_ = new_n7606_;
  assign new_n7608_ = new_n7606_;
  assign new_n7609_ = new_n7605_;
  assign new_n7610_ = new_n7609_;
  assign new_n7611_ = new_n7609_;
  assign new_n7612_ = new_n7604_;
  assign new_n7613_ = new_n7612_;
  assign new_n7614_ = new_n7613_;
  assign new_n7615_ = new_n7613_;
  assign new_n7616_ = new_n7612_;
  assign new_n7617_ = new_n1530_;
  assign new_n7618_ = new_n7617_;
  assign new_n7619_ = new_n1529_;
  assign new_n7620_ = new_n7619_;
  assign new_n7621_ = new_n2811_;
  assign new_n7622_ = new_n2809_;
  assign new_n7623_ = new_n2810_;
  assign new_n7624_ = new_n2808_;
  assign new_n7625_ = new_n2813_;
  assign new_n7626_ = new_n7625_;
  assign new_n7627_ = new_n2812_;
  assign new_n7628_ = new_n7627_;
  assign new_n7629_ = new_n1131_;
  assign new_n7630_ = new_n7629_;
  assign new_n7631_ = new_n7630_;
  assign new_n7632_ = new_n7629_;
  assign new_n7633_ = new_n1132_;
  assign new_n7634_ = new_n7633_;
  assign new_n7635_ = new_n7634_;
  assign new_n7636_ = new_n7633_;
  assign new_n7637_ = new_n2821_;
  assign new_n7638_ = new_n2819_;
  assign new_n7639_ = new_n2820_;
  assign new_n7640_ = new_n2818_;
  assign new_n7641_ = new_n2823_;
  assign new_n7642_ = new_n7641_;
  assign new_n7643_ = new_n2822_;
  assign new_n7644_ = new_n7643_;
  assign new_n7645_ = new_n2831_;
  assign new_n7646_ = new_n2829_;
  assign new_n7647_ = new_n2830_;
  assign new_n7648_ = new_n2828_;
  assign new_n7649_ = new_n2833_;
  assign new_n7650_ = new_n7649_;
  assign new_n7651_ = new_n2832_;
  assign new_n7652_ = new_n7651_;
  assign new_n7653_ = new_n2841_;
  assign new_n7654_ = new_n2839_;
  assign new_n7655_ = new_n2840_;
  assign new_n7656_ = new_n2838_;
  assign new_n7657_ = new_n2843_;
  assign new_n7658_ = new_n7657_;
  assign new_n7659_ = new_n2842_;
  assign new_n7660_ = new_n7659_;
  assign new_n7661_ = new_n2321_;
  assign new_n7662_ = new_n2851_;
  assign new_n7663_ = new_n2849_;
  assign new_n7664_ = new_n2850_;
  assign new_n7665_ = new_n2848_;
  assign new_n7666_ = new_n2853_;
  assign new_n7667_ = new_n7666_;
  assign new_n7668_ = new_n2852_;
  assign new_n7669_ = new_n7668_;
  assign new_n7670_ = new_n1615_;
  assign new_n7671_ = new_n7670_;
  assign new_n7672_ = new_n7671_;
  assign new_n7673_ = new_n7672_;
  assign new_n7674_ = new_n7672_;
  assign new_n7675_ = new_n7671_;
  assign new_n7676_ = new_n7675_;
  assign new_n7677_ = new_n7675_;
  assign new_n7678_ = new_n7670_;
  assign new_n7679_ = new_n7678_;
  assign new_n7680_ = new_n7679_;
  assign new_n7681_ = new_n7679_;
  assign new_n7682_ = new_n7678_;
  assign new_n7683_ = new_n7682_;
  assign new_n7684_ = new_n7682_;
  assign new_n7685_ = new_n1616_;
  assign new_n7686_ = new_n7685_;
  assign new_n7687_ = new_n7686_;
  assign new_n7688_ = new_n7687_;
  assign new_n7689_ = new_n7687_;
  assign new_n7690_ = new_n7686_;
  assign new_n7691_ = new_n7690_;
  assign new_n7692_ = new_n7690_;
  assign new_n7693_ = new_n7685_;
  assign new_n7694_ = new_n7693_;
  assign new_n7695_ = new_n7694_;
  assign new_n7696_ = new_n7694_;
  assign new_n7697_ = new_n7693_;
  assign new_n7698_ = new_n7697_;
  assign new_n7699_ = new_n7697_;
  assign new_n7700_ = new_n2859_;
  assign new_n7701_ = new_n2802_;
  assign new_n7702_ = new_n1303_;
  assign new_n7703_ = new_n7702_;
  assign new_n7704_ = new_n7703_;
  assign new_n7705_ = new_n7703_;
  assign new_n7706_ = new_n7702_;
  assign new_n7707_ = new_n7706_;
  assign new_n7708_ = new_n1304_;
  assign new_n7709_ = new_n7708_;
  assign new_n7710_ = new_n7709_;
  assign new_n7711_ = new_n7708_;
  assign new_n7712_ = new_n2867_;
  assign new_n7713_ = new_n2865_;
  assign new_n7714_ = new_n2866_;
  assign new_n7715_ = new_n2864_;
  assign new_n7716_ = new_n2869_;
  assign new_n7717_ = new_n7716_;
  assign new_n7718_ = new_n2868_;
  assign new_n7719_ = new_n7718_;
  assign new_n7720_ = new_n2877_;
  assign new_n7721_ = new_n2875_;
  assign new_n7722_ = new_n2876_;
  assign new_n7723_ = new_n2874_;
  assign new_n7724_ = new_n2879_;
  assign new_n7725_ = new_n7724_;
  assign new_n7726_ = new_n2878_;
  assign new_n7727_ = new_n7726_;
  assign new_n7728_ = new_n2887_;
  assign new_n7729_ = new_n2885_;
  assign new_n7730_ = new_n2886_;
  assign new_n7731_ = new_n2884_;
  assign new_n7732_ = new_n2889_;
  assign new_n7733_ = new_n7732_;
  assign new_n7734_ = new_n2888_;
  assign new_n7735_ = new_n7734_;
  assign new_n7736_ = new_n2800_;
  assign new_n7737_ = new_n2897_;
  assign new_n7738_ = new_n2895_;
  assign new_n7739_ = new_n2896_;
  assign new_n7740_ = new_n2894_;
  assign new_n7741_ = new_n2899_;
  assign new_n7742_ = new_n7741_;
  assign new_n7743_ = new_n2898_;
  assign new_n7744_ = new_n7743_;
  assign new_n7745_ = new_n2905_;
  assign new_n7746_ = new_n2860_;
  assign new_n7747_ = new_n2799_;
  assign new_n7748_ = new_n7747_;
  assign new_n7749_ = new_n2921_;
  assign new_n7750_ = new_n2919_;
  assign new_n7751_ = new_n2920_;
  assign new_n7752_ = new_n2918_;
  assign new_n7753_ = new_n2923_;
  assign new_n7754_ = new_n7753_;
  assign new_n7755_ = new_n2922_;
  assign new_n7756_ = new_n7755_;
  assign new_n7757_ = new_n2931_;
  assign new_n7758_ = new_n2929_;
  assign new_n7759_ = new_n2930_;
  assign new_n7760_ = new_n2928_;
  assign new_n7761_ = new_n2933_;
  assign new_n7762_ = new_n7761_;
  assign new_n7763_ = new_n2932_;
  assign new_n7764_ = new_n7763_;
  assign new_n7765_ = new_n2941_;
  assign new_n7766_ = new_n2939_;
  assign new_n7767_ = new_n2940_;
  assign new_n7768_ = new_n2938_;
  assign new_n7769_ = new_n2943_;
  assign new_n7770_ = new_n7769_;
  assign new_n7771_ = new_n2942_;
  assign new_n7772_ = new_n7771_;
  assign new_n7773_ = new_n2951_;
  assign new_n7774_ = new_n2949_;
  assign new_n7775_ = new_n2950_;
  assign new_n7776_ = new_n2948_;
  assign new_n7777_ = new_n2953_;
  assign new_n7778_ = new_n7777_;
  assign new_n7779_ = new_n2952_;
  assign new_n7780_ = new_n7779_;
  assign new_n7781_ = new_n2970_;
  assign new_n7782_ = new_n2968_;
  assign new_n7783_ = new_n2969_;
  assign new_n7784_ = new_n2967_;
  assign new_n7785_ = new_n2972_;
  assign new_n7786_ = new_n7785_;
  assign new_n7787_ = new_n2971_;
  assign new_n7788_ = new_n7787_;
  assign new_n7789_ = new_n2980_;
  assign new_n7790_ = new_n2978_;
  assign new_n7791_ = new_n2979_;
  assign new_n7792_ = new_n2977_;
  assign new_n7793_ = new_n2982_;
  assign new_n7794_ = new_n7793_;
  assign new_n7795_ = new_n2981_;
  assign new_n7796_ = new_n7795_;
  assign new_n7797_ = new_n2990_;
  assign new_n7798_ = new_n2988_;
  assign new_n7799_ = new_n2989_;
  assign new_n7800_ = new_n2987_;
  assign new_n7801_ = new_n2992_;
  assign new_n7802_ = new_n7801_;
  assign new_n7803_ = new_n2991_;
  assign new_n7804_ = new_n7803_;
  assign new_n7805_ = new_n3000_;
  assign new_n7806_ = new_n2998_;
  assign new_n7807_ = new_n2999_;
  assign new_n7808_ = new_n2997_;
  assign new_n7809_ = new_n3002_;
  assign new_n7810_ = new_n7809_;
  assign new_n7811_ = new_n3001_;
  assign new_n7812_ = new_n7811_;
  assign new_n7813_ = new_n3025_;
  assign new_n7814_ = new_n3023_;
  assign new_n7815_ = new_n3024_;
  assign new_n7816_ = new_n3022_;
  assign new_n7817_ = new_n3027_;
  assign new_n7818_ = new_n7817_;
  assign new_n7819_ = new_n3026_;
  assign new_n7820_ = new_n7819_;
  assign new_n7821_ = new_n1029_;
  assign new_n7822_ = new_n7821_;
  assign new_n7823_ = new_n1030_;
  assign new_n7824_ = new_n7823_;
  assign new_n7825_ = new_n3035_;
  assign new_n7826_ = new_n3033_;
  assign new_n7827_ = new_n3034_;
  assign new_n7828_ = new_n3032_;
  assign new_n7829_ = new_n3037_;
  assign new_n7830_ = new_n7829_;
  assign new_n7831_ = new_n3036_;
  assign new_n7832_ = new_n7831_;
  assign new_n7833_ = new_n3039_;
  assign new_n7834_ = new_n3017_;
  assign new_n7835_ = new_n3038_;
  assign new_n7836_ = new_n3016_;
  assign new_n7837_ = new_n3041_;
  assign new_n7838_ = new_n7837_;
  assign new_n7839_ = new_n3040_;
  assign new_n7840_ = new_n7839_;
  assign new_n7841_ = new_n3049_;
  assign new_n7842_ = new_n3047_;
  assign new_n7843_ = new_n3048_;
  assign new_n7844_ = new_n3046_;
  assign new_n7845_ = new_n3051_;
  assign new_n7846_ = new_n7845_;
  assign new_n7847_ = new_n3050_;
  assign new_n7848_ = new_n7847_;
  assign new_n7849_ = new_n3065_;
  assign new_n7850_ = new_n3063_;
  assign new_n7851_ = new_n3064_;
  assign new_n7852_ = new_n3062_;
  assign new_n7853_ = new_n3067_;
  assign new_n7854_ = new_n7853_;
  assign new_n7855_ = new_n3066_;
  assign new_n7856_ = new_n7855_;
  assign new_n7857_ = new_n3075_;
  assign new_n7858_ = new_n3073_;
  assign new_n7859_ = new_n3074_;
  assign new_n7860_ = new_n3072_;
  assign new_n7861_ = new_n3077_;
  assign new_n7862_ = new_n7861_;
  assign new_n7863_ = new_n3076_;
  assign new_n7864_ = new_n7863_;
  assign new_n7865_ = new_n3079_;
  assign new_n7866_ = new_n3057_;
  assign new_n7867_ = new_n3078_;
  assign new_n7868_ = new_n3056_;
  assign new_n7869_ = new_n3081_;
  assign new_n7870_ = new_n7869_;
  assign new_n7871_ = new_n3080_;
  assign new_n7872_ = new_n7871_;
  assign new_n7873_ = new_n3089_;
  assign new_n7874_ = new_n3087_;
  assign new_n7875_ = new_n3088_;
  assign new_n7876_ = new_n3086_;
  assign new_n7877_ = new_n3091_;
  assign new_n7878_ = new_n7877_;
  assign new_n7879_ = new_n3090_;
  assign new_n7880_ = new_n7879_;
  assign new_n7881_ = new_n3105_;
  assign new_n7882_ = new_n3103_;
  assign new_n7883_ = new_n3104_;
  assign new_n7884_ = new_n3102_;
  assign new_n7885_ = new_n3107_;
  assign new_n7886_ = new_n7885_;
  assign new_n7887_ = new_n3106_;
  assign new_n7888_ = new_n7887_;
  assign new_n7889_ = new_n3115_;
  assign new_n7890_ = new_n3113_;
  assign new_n7891_ = new_n3114_;
  assign new_n7892_ = new_n3112_;
  assign new_n7893_ = new_n3117_;
  assign new_n7894_ = new_n7893_;
  assign new_n7895_ = new_n3116_;
  assign new_n7896_ = new_n7895_;
  assign new_n7897_ = new_n3128_;
  assign new_n7898_ = new_n3126_;
  assign new_n7899_ = new_n3130_;
  assign new_n7900_ = new_n895_;
  assign new_n7901_ = new_n7900_;
  assign new_n7902_ = new_n7901_;
  assign new_n7903_ = new_n7902_;
  assign new_n7904_ = new_n7902_;
  assign new_n7905_ = new_n7901_;
  assign new_n7906_ = new_n7905_;
  assign new_n7907_ = new_n7905_;
  assign new_n7908_ = new_n7900_;
  assign new_n7909_ = new_n7908_;
  assign new_n7910_ = new_n7909_;
  assign new_n7911_ = new_n7909_;
  assign new_n7912_ = new_n7908_;
  assign new_n7913_ = new_n7912_;
  assign new_n7914_ = new_n7912_;
  assign new_n7915_ = new_n896_;
  assign new_n7916_ = new_n7915_;
  assign new_n7917_ = new_n7916_;
  assign new_n7918_ = new_n7917_;
  assign new_n7919_ = new_n7917_;
  assign new_n7920_ = new_n7916_;
  assign new_n7921_ = new_n7920_;
  assign new_n7922_ = new_n7920_;
  assign new_n7923_ = new_n7915_;
  assign new_n7924_ = new_n7923_;
  assign new_n7925_ = new_n7924_;
  assign new_n7926_ = new_n7924_;
  assign new_n7927_ = new_n7923_;
  assign new_n7928_ = new_n7927_;
  assign new_n7929_ = new_n7927_;
  assign new_n7930_ = new_n2734_;
  assign new_n7931_ = new_n7930_;
  assign new_n7932_ = new_n2733_;
  assign new_n7933_ = new_n2586_;
  assign new_n7934_ = new_n7933_;
  assign new_n7935_ = new_n2585_;
  assign new_n7936_ = new_n2438_;
  assign new_n7937_ = new_n7936_;
  assign new_n7938_ = new_n2437_;
  assign new_n7939_ = new_n3133_;
  assign new_n7940_ = new_n2908_;
  assign new_n7941_ = new_n1089_;
  assign new_n7942_ = new_n7941_;
  assign new_n7943_ = new_n7941_;
  assign new_n7944_ = new_n1090_;
  assign new_n7945_ = new_n7944_;
  assign new_n7946_ = new_n1494_;
  assign new_n7947_ = new_n1484_;
  assign new_n7948_ = new_n1493_;
  assign new_n7949_ = new_n1483_;
  assign new_n7950_ = new_n3167_;
  assign new_n7951_ = new_n7950_;
  assign new_n7952_ = new_n3166_;
  assign new_n7953_ = new_n7952_;
  assign new_n7954_ = new_n1093_;
  assign new_n7955_ = new_n7954_;
  assign new_n7956_ = new_n7954_;
  assign new_n7957_ = new_n1094_;
  assign new_n7958_ = new_n7957_;
  assign new_n7959_ = new_n3175_;
  assign new_n7960_ = new_n3173_;
  assign new_n7961_ = new_n3174_;
  assign new_n7962_ = new_n3172_;
  assign new_n7963_ = new_n3177_;
  assign new_n7964_ = new_n7963_;
  assign new_n7965_ = new_n3176_;
  assign new_n7966_ = new_n7965_;
  assign new_n7967_ = new_n3179_;
  assign new_n7968_ = new_n3165_;
  assign new_n7969_ = new_n3178_;
  assign new_n7970_ = new_n3164_;
  assign new_n7971_ = new_n3181_;
  assign new_n7972_ = new_n7971_;
  assign new_n7973_ = new_n3180_;
  assign new_n7974_ = new_n7973_;
  assign new_n7975_ = new_n3189_;
  assign new_n7976_ = new_n3187_;
  assign new_n7977_ = new_n3188_;
  assign new_n7978_ = new_n3186_;
  assign new_n7979_ = new_n3191_;
  assign new_n7980_ = new_n7979_;
  assign new_n7981_ = new_n3190_;
  assign new_n7982_ = new_n7981_;
  assign new_n7983_ = new_n1101_;
  assign new_n7984_ = new_n7983_;
  assign new_n7985_ = new_n7983_;
  assign new_n7986_ = new_n1102_;
  assign new_n7987_ = new_n7986_;
  assign new_n7988_ = new_n7986_;
  assign new_n7989_ = new_n3207_;
  assign new_n7990_ = new_n3205_;
  assign new_n7991_ = new_n3206_;
  assign new_n7992_ = new_n3204_;
  assign new_n7993_ = new_n3209_;
  assign new_n7994_ = new_n7993_;
  assign new_n7995_ = new_n3208_;
  assign new_n7996_ = new_n7995_;
  assign new_n7997_ = new_n3211_;
  assign new_n7998_ = new_n3203_;
  assign new_n7999_ = new_n3210_;
  assign new_n8000_ = new_n3202_;
  assign new_n8001_ = new_n3213_;
  assign new_n8002_ = new_n8001_;
  assign new_n8003_ = new_n3212_;
  assign new_n8004_ = new_n8003_;
  assign new_n8005_ = new_n3221_;
  assign new_n8006_ = new_n3219_;
  assign new_n8007_ = new_n3220_;
  assign new_n8008_ = new_n3218_;
  assign new_n8009_ = new_n3223_;
  assign new_n8010_ = new_n8009_;
  assign new_n8011_ = new_n3222_;
  assign new_n8012_ = new_n8011_;
  assign new_n8013_ = new_n3225_;
  assign new_n8014_ = new_n3197_;
  assign new_n8015_ = new_n3224_;
  assign new_n8016_ = new_n3196_;
  assign new_n8017_ = new_n3227_;
  assign new_n8018_ = new_n8017_;
  assign new_n8019_ = new_n3226_;
  assign new_n8020_ = new_n8019_;
  assign new_n8021_ = new_n3235_;
  assign new_n8022_ = new_n3233_;
  assign new_n8023_ = new_n3234_;
  assign new_n8024_ = new_n3232_;
  assign new_n8025_ = new_n3237_;
  assign new_n8026_ = new_n8025_;
  assign new_n8027_ = new_n3236_;
  assign new_n8028_ = new_n8027_;
  assign new_n8029_ = new_n1526_;
  assign new_n8030_ = new_n8029_;
  assign new_n8031_ = new_n1525_;
  assign new_n8032_ = new_n8031_;
  assign new_n8033_ = new_n3257_;
  assign new_n8034_ = new_n3255_;
  assign new_n8035_ = new_n3256_;
  assign new_n8036_ = new_n3254_;
  assign new_n8037_ = new_n3259_;
  assign new_n8038_ = new_n8037_;
  assign new_n8039_ = new_n3258_;
  assign new_n8040_ = new_n8039_;
  assign new_n8041_ = new_n1103_;
  assign new_n8042_ = new_n8041_;
  assign new_n8043_ = new_n8041_;
  assign new_n8044_ = new_n1104_;
  assign new_n8045_ = new_n8044_;
  assign new_n8046_ = new_n3267_;
  assign new_n8047_ = new_n3265_;
  assign new_n8048_ = new_n3266_;
  assign new_n8049_ = new_n3264_;
  assign new_n8050_ = new_n3269_;
  assign new_n8051_ = new_n8050_;
  assign new_n8052_ = new_n3268_;
  assign new_n8053_ = new_n8052_;
  assign new_n8054_ = new_n3271_;
  assign new_n8055_ = new_n3249_;
  assign new_n8056_ = new_n3270_;
  assign new_n8057_ = new_n3248_;
  assign new_n8058_ = new_n3273_;
  assign new_n8059_ = new_n8058_;
  assign new_n8060_ = new_n3272_;
  assign new_n8061_ = new_n8060_;
  assign new_n8062_ = new_n3281_;
  assign new_n8063_ = new_n3279_;
  assign new_n8064_ = new_n3280_;
  assign new_n8065_ = new_n3278_;
  assign new_n8066_ = new_n3283_;
  assign new_n8067_ = new_n8066_;
  assign new_n8068_ = new_n3282_;
  assign new_n8069_ = new_n8068_;
  assign new_n8070_ = new_n3285_;
  assign new_n8071_ = new_n3243_;
  assign new_n8072_ = new_n3284_;
  assign new_n8073_ = new_n3242_;
  assign new_n8074_ = new_n3295_;
  assign new_n8075_ = new_n3293_;
  assign new_n8076_ = new_n3294_;
  assign new_n8077_ = new_n3292_;
  assign new_n8078_ = new_n3297_;
  assign new_n8079_ = new_n8078_;
  assign new_n8080_ = new_n3296_;
  assign new_n8081_ = new_n8080_;
  assign new_n8082_ = new_n1107_;
  assign new_n8083_ = new_n8082_;
  assign new_n8084_ = new_n8082_;
  assign new_n8085_ = new_n1108_;
  assign new_n8086_ = new_n8085_;
  assign new_n8087_ = new_n3305_;
  assign new_n8088_ = new_n3303_;
  assign new_n8089_ = new_n3304_;
  assign new_n8090_ = new_n3302_;
  assign new_n8091_ = new_n3307_;
  assign new_n8092_ = new_n8091_;
  assign new_n8093_ = new_n3306_;
  assign new_n8094_ = new_n8093_;
  assign new_n8095_ = new_n1544_;
  assign new_n8096_ = new_n1496_;
  assign new_n8097_ = new_n1543_;
  assign new_n8098_ = new_n1495_;
  assign new_n8099_ = new_n3315_;
  assign new_n8100_ = new_n8099_;
  assign new_n8101_ = new_n3314_;
  assign new_n8102_ = new_n8101_;
  assign new_n8103_ = new_n1109_;
  assign new_n8104_ = new_n8103_;
  assign new_n8105_ = new_n8103_;
  assign new_n8106_ = new_n1110_;
  assign new_n8107_ = new_n8106_;
  assign new_n8108_ = new_n3323_;
  assign new_n8109_ = new_n3321_;
  assign new_n8110_ = new_n3322_;
  assign new_n8111_ = new_n3320_;
  assign new_n8112_ = new_n3325_;
  assign new_n8113_ = new_n8112_;
  assign new_n8114_ = new_n3324_;
  assign new_n8115_ = new_n8114_;
  assign new_n8116_ = new_n3327_;
  assign new_n8117_ = new_n3313_;
  assign new_n8118_ = new_n3326_;
  assign new_n8119_ = new_n3312_;
  assign new_n8120_ = new_n3329_;
  assign new_n8121_ = new_n8120_;
  assign new_n8122_ = new_n3328_;
  assign new_n8123_ = new_n8122_;
  assign new_n8124_ = new_n3337_;
  assign new_n8125_ = new_n3335_;
  assign new_n8126_ = new_n3336_;
  assign new_n8127_ = new_n3334_;
  assign new_n8128_ = new_n3339_;
  assign new_n8129_ = new_n8128_;
  assign new_n8130_ = new_n3338_;
  assign new_n8131_ = new_n8130_;
  assign new_n8132_ = new_n1111_;
  assign new_n8133_ = new_n8132_;
  assign new_n8134_ = new_n8132_;
  assign new_n8135_ = new_n1112_;
  assign new_n8136_ = new_n8135_;
  assign new_n8137_ = new_n8135_;
  assign new_n8138_ = new_n3355_;
  assign new_n8139_ = new_n3353_;
  assign new_n8140_ = new_n3354_;
  assign new_n8141_ = new_n3352_;
  assign new_n8142_ = new_n3357_;
  assign new_n8143_ = new_n8142_;
  assign new_n8144_ = new_n3356_;
  assign new_n8145_ = new_n8144_;
  assign new_n8146_ = new_n3359_;
  assign new_n8147_ = new_n3351_;
  assign new_n8148_ = new_n3358_;
  assign new_n8149_ = new_n3350_;
  assign new_n8150_ = new_n3361_;
  assign new_n8151_ = new_n8150_;
  assign new_n8152_ = new_n3360_;
  assign new_n8153_ = new_n8152_;
  assign new_n8154_ = new_n3369_;
  assign new_n8155_ = new_n3367_;
  assign new_n8156_ = new_n3368_;
  assign new_n8157_ = new_n3366_;
  assign new_n8158_ = new_n3371_;
  assign new_n8159_ = new_n8158_;
  assign new_n8160_ = new_n3370_;
  assign new_n8161_ = new_n8160_;
  assign new_n8162_ = new_n3373_;
  assign new_n8163_ = new_n3345_;
  assign new_n8164_ = new_n3372_;
  assign new_n8165_ = new_n3344_;
  assign new_n8166_ = new_n3375_;
  assign new_n8167_ = new_n8166_;
  assign new_n8168_ = new_n3374_;
  assign new_n8169_ = new_n8168_;
  assign new_n8170_ = new_n3383_;
  assign new_n8171_ = new_n3381_;
  assign new_n8172_ = new_n3382_;
  assign new_n8173_ = new_n3380_;
  assign new_n8174_ = new_n3385_;
  assign new_n8175_ = new_n8174_;
  assign new_n8176_ = new_n3384_;
  assign new_n8177_ = new_n8176_;
  assign new_n8178_ = new_n1528_;
  assign new_n8179_ = new_n8178_;
  assign new_n8180_ = new_n1527_;
  assign new_n8181_ = new_n8180_;
  assign new_n8182_ = new_n3405_;
  assign new_n8183_ = new_n3403_;
  assign new_n8184_ = new_n3404_;
  assign new_n8185_ = new_n3402_;
  assign new_n8186_ = new_n3407_;
  assign new_n8187_ = new_n8186_;
  assign new_n8188_ = new_n3406_;
  assign new_n8189_ = new_n8188_;
  assign new_n8190_ = new_n1113_;
  assign new_n8191_ = new_n8190_;
  assign new_n8192_ = new_n8190_;
  assign new_n8193_ = new_n1114_;
  assign new_n8194_ = new_n8193_;
  assign new_n8195_ = new_n3415_;
  assign new_n8196_ = new_n3413_;
  assign new_n8197_ = new_n3414_;
  assign new_n8198_ = new_n3412_;
  assign new_n8199_ = new_n3417_;
  assign new_n8200_ = new_n8199_;
  assign new_n8201_ = new_n3416_;
  assign new_n8202_ = new_n8201_;
  assign new_n8203_ = new_n3419_;
  assign new_n8204_ = new_n3397_;
  assign new_n8205_ = new_n3418_;
  assign new_n8206_ = new_n3396_;
  assign new_n8207_ = new_n3421_;
  assign new_n8208_ = new_n8207_;
  assign new_n8209_ = new_n3420_;
  assign new_n8210_ = new_n8209_;
  assign new_n8211_ = new_n3429_;
  assign new_n8212_ = new_n3427_;
  assign new_n8213_ = new_n3428_;
  assign new_n8214_ = new_n3426_;
  assign new_n8215_ = new_n3431_;
  assign new_n8216_ = new_n8215_;
  assign new_n8217_ = new_n3430_;
  assign new_n8218_ = new_n8217_;
  assign new_n8219_ = new_n3433_;
  assign new_n8220_ = new_n3391_;
  assign new_n8221_ = new_n3432_;
  assign new_n8222_ = new_n3390_;
  assign new_n8223_ = new_n1549_;
  assign new_n8224_ = new_n1486_;
  assign new_n8225_ = new_n1550_;
  assign new_n8226_ = new_n1485_;
  assign new_n8227_ = new_n3443_;
  assign new_n8228_ = new_n8227_;
  assign new_n8229_ = new_n3442_;
  assign new_n8230_ = new_n8229_;
  assign new_n8231_ = new_n3445_;
  assign new_n8232_ = new_n3441_;
  assign new_n8233_ = new_n3444_;
  assign new_n8234_ = new_n3440_;
  assign new_n8235_ = new_n3447_;
  assign new_n8236_ = new_n8235_;
  assign new_n8237_ = new_n3446_;
  assign new_n8238_ = new_n8237_;
  assign new_n8239_ = new_n1115_;
  assign new_n8240_ = new_n8239_;
  assign new_n8241_ = new_n8239_;
  assign new_n8242_ = new_n1116_;
  assign new_n8243_ = new_n8242_;
  assign new_n8244_ = new_n3455_;
  assign new_n8245_ = new_n3453_;
  assign new_n8246_ = new_n3454_;
  assign new_n8247_ = new_n3452_;
  assign new_n8248_ = new_n3457_;
  assign new_n8249_ = new_n8248_;
  assign new_n8250_ = new_n3456_;
  assign new_n8251_ = new_n8250_;
  assign new_n8252_ = new_n1119_;
  assign new_n8253_ = new_n8252_;
  assign new_n8254_ = new_n8253_;
  assign new_n8255_ = new_n8252_;
  assign new_n8256_ = new_n1120_;
  assign new_n8257_ = new_n8256_;
  assign new_n8258_ = new_n8256_;
  assign new_n8259_ = new_n3473_;
  assign new_n8260_ = new_n3471_;
  assign new_n8261_ = new_n3472_;
  assign new_n8262_ = new_n3470_;
  assign new_n8263_ = new_n3475_;
  assign new_n8264_ = new_n8263_;
  assign new_n8265_ = new_n3474_;
  assign new_n8266_ = new_n8265_;
  assign new_n8267_ = new_n3477_;
  assign new_n8268_ = new_n3469_;
  assign new_n8269_ = new_n3476_;
  assign new_n8270_ = new_n3468_;
  assign new_n8271_ = new_n3479_;
  assign new_n8272_ = new_n8271_;
  assign new_n8273_ = new_n3478_;
  assign new_n8274_ = new_n8273_;
  assign new_n8275_ = new_n3487_;
  assign new_n8276_ = new_n3485_;
  assign new_n8277_ = new_n3486_;
  assign new_n8278_ = new_n3484_;
  assign new_n8279_ = new_n3489_;
  assign new_n8280_ = new_n8279_;
  assign new_n8281_ = new_n3488_;
  assign new_n8282_ = new_n8281_;
  assign new_n8283_ = new_n3491_;
  assign new_n8284_ = new_n3463_;
  assign new_n8285_ = new_n3490_;
  assign new_n8286_ = new_n3462_;
  assign new_n8287_ = new_n3493_;
  assign new_n8288_ = new_n8287_;
  assign new_n8289_ = new_n3492_;
  assign new_n8290_ = new_n8289_;
  assign new_n8291_ = new_n3501_;
  assign new_n8292_ = new_n3499_;
  assign new_n8293_ = new_n3500_;
  assign new_n8294_ = new_n3498_;
  assign new_n8295_ = new_n3503_;
  assign new_n8296_ = new_n8295_;
  assign new_n8297_ = new_n3502_;
  assign new_n8298_ = new_n8297_;
  assign new_n8299_ = new_n1535_;
  assign new_n8300_ = new_n8299_;
  assign new_n8301_ = new_n1536_;
  assign new_n8302_ = new_n8301_;
  assign new_n8303_ = new_n1123_;
  assign new_n8304_ = new_n8303_;
  assign new_n8305_ = new_n8304_;
  assign new_n8306_ = new_n8303_;
  assign new_n8307_ = new_n1124_;
  assign new_n8308_ = new_n8307_;
  assign new_n8309_ = new_n8308_;
  assign new_n8310_ = new_n8307_;
  assign new_n8311_ = new_n3529_;
  assign new_n8312_ = new_n3527_;
  assign new_n8313_ = new_n3528_;
  assign new_n8314_ = new_n3526_;
  assign new_n8315_ = new_n3531_;
  assign new_n8316_ = new_n8315_;
  assign new_n8317_ = new_n3530_;
  assign new_n8318_ = new_n8317_;
  assign new_n8319_ = new_n3533_;
  assign new_n8320_ = new_n3521_;
  assign new_n8321_ = new_n3532_;
  assign new_n8322_ = new_n3520_;
  assign new_n8323_ = new_n3535_;
  assign new_n8324_ = new_n8323_;
  assign new_n8325_ = new_n3534_;
  assign new_n8326_ = new_n8325_;
  assign new_n8327_ = new_n3543_;
  assign new_n8328_ = new_n3541_;
  assign new_n8329_ = new_n3542_;
  assign new_n8330_ = new_n3540_;
  assign new_n8331_ = new_n3545_;
  assign new_n8332_ = new_n8331_;
  assign new_n8333_ = new_n3544_;
  assign new_n8334_ = new_n8333_;
  assign new_n8335_ = new_n3547_;
  assign new_n8336_ = new_n3515_;
  assign new_n8337_ = new_n3546_;
  assign new_n8338_ = new_n3514_;
  assign new_n8339_ = new_n3549_;
  assign new_n8340_ = new_n8339_;
  assign new_n8341_ = new_n3548_;
  assign new_n8342_ = new_n8341_;
  assign new_n8343_ = new_n3557_;
  assign new_n8344_ = new_n3555_;
  assign new_n8345_ = new_n3556_;
  assign new_n8346_ = new_n3554_;
  assign new_n8347_ = new_n3559_;
  assign new_n8348_ = new_n8347_;
  assign new_n8349_ = new_n3558_;
  assign new_n8350_ = new_n8349_;
  assign new_n8351_ = new_n3561_;
  assign new_n8352_ = new_n3509_;
  assign new_n8353_ = new_n3560_;
  assign new_n8354_ = new_n3508_;
  assign new_n8355_ = new_n3563_;
  assign new_n8356_ = new_n8355_;
  assign new_n8357_ = new_n3562_;
  assign new_n8358_ = new_n8357_;
  assign new_n8359_ = new_n913_;
  assign new_n8360_ = new_n8359_;
  assign new_n8361_ = new_n8360_;
  assign new_n8362_ = new_n8361_;
  assign new_n8363_ = new_n8361_;
  assign new_n8364_ = new_n8360_;
  assign new_n8365_ = new_n8359_;
  assign new_n8366_ = new_n8365_;
  assign new_n8367_ = new_n8365_;
  assign new_n8368_ = new_n914_;
  assign new_n8369_ = new_n8368_;
  assign new_n8370_ = new_n8369_;
  assign new_n8371_ = new_n8370_;
  assign new_n8372_ = new_n8370_;
  assign new_n8373_ = new_n8369_;
  assign new_n8374_ = new_n8368_;
  assign new_n8375_ = new_n8374_;
  assign new_n8376_ = new_n8374_;
  assign new_n8377_ = new_n3571_;
  assign new_n8378_ = new_n3569_;
  assign new_n8379_ = new_n3570_;
  assign new_n8380_ = new_n3568_;
  assign new_n8381_ = new_n3573_;
  assign new_n8382_ = new_n8381_;
  assign new_n8383_ = new_n3572_;
  assign new_n8384_ = new_n8383_;
  assign new_n8385_ = new_n1546_;
  assign new_n8386_ = new_n1498_;
  assign new_n8387_ = new_n1545_;
  assign new_n8388_ = new_n1497_;
  assign new_n8389_ = new_n3599_;
  assign new_n8390_ = new_n8389_;
  assign new_n8391_ = new_n3598_;
  assign new_n8392_ = new_n8391_;
  assign new_n8393_ = new_n1127_;
  assign new_n8394_ = new_n8393_;
  assign new_n8395_ = new_n8394_;
  assign new_n8396_ = new_n8394_;
  assign new_n8397_ = new_n8393_;
  assign new_n8398_ = new_n1128_;
  assign new_n8399_ = new_n8398_;
  assign new_n8400_ = new_n8399_;
  assign new_n8401_ = new_n8398_;
  assign new_n8402_ = new_n3607_;
  assign new_n8403_ = new_n3605_;
  assign new_n8404_ = new_n3606_;
  assign new_n8405_ = new_n3604_;
  assign new_n8406_ = new_n3609_;
  assign new_n8407_ = new_n8406_;
  assign new_n8408_ = new_n3608_;
  assign new_n8409_ = new_n8408_;
  assign new_n8410_ = new_n3611_;
  assign new_n8411_ = new_n3597_;
  assign new_n8412_ = new_n3610_;
  assign new_n8413_ = new_n3596_;
  assign new_n8414_ = new_n3613_;
  assign new_n8415_ = new_n8414_;
  assign new_n8416_ = new_n3612_;
  assign new_n8417_ = new_n8416_;
  assign new_n8418_ = new_n3621_;
  assign new_n8419_ = new_n3619_;
  assign new_n8420_ = new_n3620_;
  assign new_n8421_ = new_n3618_;
  assign new_n8422_ = new_n3623_;
  assign new_n8423_ = new_n8422_;
  assign new_n8424_ = new_n3622_;
  assign new_n8425_ = new_n8424_;
  assign new_n8426_ = new_n3625_;
  assign new_n8427_ = new_n3591_;
  assign new_n8428_ = new_n3624_;
  assign new_n8429_ = new_n3590_;
  assign new_n8430_ = new_n3627_;
  assign new_n8431_ = new_n8430_;
  assign new_n8432_ = new_n3626_;
  assign new_n8433_ = new_n8432_;
  assign new_n8434_ = new_n3635_;
  assign new_n8435_ = new_n3633_;
  assign new_n8436_ = new_n3634_;
  assign new_n8437_ = new_n3632_;
  assign new_n8438_ = new_n3637_;
  assign new_n8439_ = new_n8438_;
  assign new_n8440_ = new_n3636_;
  assign new_n8441_ = new_n8440_;
  assign new_n8442_ = new_n3639_;
  assign new_n8443_ = new_n3585_;
  assign new_n8444_ = new_n3638_;
  assign new_n8445_ = new_n3584_;
  assign new_n8446_ = new_n3641_;
  assign new_n8447_ = new_n8446_;
  assign new_n8448_ = new_n3640_;
  assign new_n8449_ = new_n8448_;
  assign new_n8450_ = new_n3649_;
  assign new_n8451_ = new_n3647_;
  assign new_n8452_ = new_n3648_;
  assign new_n8453_ = new_n3646_;
  assign new_n8454_ = new_n3651_;
  assign new_n8455_ = new_n8454_;
  assign new_n8456_ = new_n3650_;
  assign new_n8457_ = new_n8456_;
  assign new_n8458_ = new_n3653_;
  assign new_n8459_ = new_n3579_;
  assign new_n8460_ = new_n3652_;
  assign new_n8461_ = new_n3578_;
  assign new_n8462_ = new_n1611_;
  assign new_n8463_ = new_n1564_;
  assign new_n8464_ = new_n1612_;
  assign new_n8465_ = new_n1563_;
  assign new_n8466_ = new_n3657_;
  assign new_n8467_ = new_n8466_;
  assign new_n8468_ = new_n3656_;
  assign new_n8469_ = new_n8468_;
  assign new_n8470_ = new_n3665_;
  assign new_n8471_ = new_n3663_;
  assign new_n8472_ = new_n3664_;
  assign new_n8473_ = new_n3662_;
  assign new_n8474_ = new_n3667_;
  assign new_n8475_ = new_n8474_;
  assign new_n8476_ = new_n3666_;
  assign new_n8477_ = new_n8476_;
  assign new_n8478_ = new_n3675_;
  assign new_n8479_ = new_n3673_;
  assign new_n8480_ = new_n3674_;
  assign new_n8481_ = new_n3672_;
  assign new_n8482_ = new_n3677_;
  assign new_n8483_ = new_n8482_;
  assign new_n8484_ = new_n3676_;
  assign new_n8485_ = new_n8484_;
  assign new_n8486_ = new_n3685_;
  assign new_n8487_ = new_n3683_;
  assign new_n8488_ = new_n3684_;
  assign new_n8489_ = new_n3682_;
  assign new_n8490_ = new_n3687_;
  assign new_n8491_ = new_n8490_;
  assign new_n8492_ = new_n3686_;
  assign new_n8493_ = new_n8492_;
  assign new_n8494_ = new_n3695_;
  assign new_n8495_ = new_n3693_;
  assign new_n8496_ = new_n3694_;
  assign new_n8497_ = new_n3692_;
  assign new_n8498_ = new_n3697_;
  assign new_n8499_ = new_n8498_;
  assign new_n8500_ = new_n3696_;
  assign new_n8501_ = new_n8500_;
  assign new_n8502_ = new_n2906_;
  assign new_n8503_ = new_n3705_;
  assign new_n8504_ = new_n3703_;
  assign new_n8505_ = new_n3704_;
  assign new_n8506_ = new_n3702_;
  assign new_n8507_ = new_n3707_;
  assign new_n8508_ = new_n8507_;
  assign new_n8509_ = new_n3706_;
  assign new_n8510_ = new_n8509_;
  assign new_n8511_ = new_n3713_;
  assign new_n8512_ = new_n3134_;
  assign new_n8513_ = new_n3721_;
  assign new_n8514_ = new_n3719_;
  assign new_n8515_ = new_n3720_;
  assign new_n8516_ = new_n3718_;
  assign new_n8517_ = new_n3723_;
  assign new_n8518_ = new_n8517_;
  assign new_n8519_ = new_n3722_;
  assign new_n8520_ = new_n8519_;
  assign new_n8521_ = new_n1129_;
  assign new_n8522_ = new_n8521_;
  assign new_n8523_ = new_n8522_;
  assign new_n8524_ = new_n8522_;
  assign new_n8525_ = new_n8521_;
  assign new_n8526_ = new_n1130_;
  assign new_n8527_ = new_n8526_;
  assign new_n8528_ = new_n8527_;
  assign new_n8529_ = new_n8526_;
  assign new_n8530_ = new_n3731_;
  assign new_n8531_ = new_n3729_;
  assign new_n8532_ = new_n3730_;
  assign new_n8533_ = new_n3728_;
  assign new_n8534_ = new_n3733_;
  assign new_n8535_ = new_n8534_;
  assign new_n8536_ = new_n3732_;
  assign new_n8537_ = new_n8536_;
  assign new_n8538_ = new_n3741_;
  assign new_n8539_ = new_n3739_;
  assign new_n8540_ = new_n3740_;
  assign new_n8541_ = new_n3738_;
  assign new_n8542_ = new_n3743_;
  assign new_n8543_ = new_n8542_;
  assign new_n8544_ = new_n3742_;
  assign new_n8545_ = new_n8544_;
  assign new_n8546_ = new_n3751_;
  assign new_n8547_ = new_n3749_;
  assign new_n8548_ = new_n3750_;
  assign new_n8549_ = new_n3748_;
  assign new_n8550_ = new_n3753_;
  assign new_n8551_ = new_n8550_;
  assign new_n8552_ = new_n3752_;
  assign new_n8553_ = new_n8552_;
  assign new_n8554_ = new_n3761_;
  assign new_n8555_ = new_n3759_;
  assign new_n8556_ = new_n3760_;
  assign new_n8557_ = new_n3758_;
  assign new_n8558_ = new_n3763_;
  assign new_n8559_ = new_n8558_;
  assign new_n8560_ = new_n3762_;
  assign new_n8561_ = new_n8560_;
  assign new_n8562_ = new_n3771_;
  assign new_n8563_ = new_n3769_;
  assign new_n8564_ = new_n3770_;
  assign new_n8565_ = new_n3768_;
  assign new_n8566_ = new_n3773_;
  assign new_n8567_ = new_n8566_;
  assign new_n8568_ = new_n3772_;
  assign new_n8569_ = new_n8568_;
  assign new_n8570_ = new_n2862_;
  assign new_n8571_ = new_n3781_;
  assign new_n8572_ = new_n3779_;
  assign new_n8573_ = new_n3780_;
  assign new_n8574_ = new_n3778_;
  assign new_n8575_ = new_n3783_;
  assign new_n8576_ = new_n8575_;
  assign new_n8577_ = new_n3782_;
  assign new_n8578_ = new_n8577_;
  assign new_n8579_ = new_n3163_;
  assign new_n8580_ = new_n3801_;
  assign new_n8581_ = new_n3799_;
  assign new_n8582_ = new_n3800_;
  assign new_n8583_ = new_n3798_;
  assign new_n8584_ = new_n3803_;
  assign new_n8585_ = new_n8584_;
  assign new_n8586_ = new_n3802_;
  assign new_n8587_ = new_n3811_;
  assign new_n8588_ = new_n3809_;
  assign new_n8589_ = new_n3810_;
  assign new_n8590_ = new_n3808_;
  assign new_n8591_ = new_n3813_;
  assign new_n8592_ = new_n8591_;
  assign new_n8593_ = new_n3812_;
  assign new_n8594_ = new_n3830_;
  assign new_n8595_ = new_n3828_;
  assign new_n8596_ = new_n3829_;
  assign new_n8597_ = new_n3827_;
  assign new_n8598_ = new_n3832_;
  assign new_n8599_ = new_n8598_;
  assign new_n8600_ = new_n3831_;
  assign new_n8601_ = new_n3840_;
  assign new_n8602_ = new_n3838_;
  assign new_n8603_ = new_n3839_;
  assign new_n8604_ = new_n3837_;
  assign new_n8605_ = new_n3842_;
  assign new_n8606_ = new_n8605_;
  assign new_n8607_ = new_n3841_;
  assign new_n8608_ = new_n3859_;
  assign new_n8609_ = new_n3857_;
  assign new_n8610_ = new_n3858_;
  assign new_n8611_ = new_n3856_;
  assign new_n8612_ = new_n3861_;
  assign new_n8613_ = new_n8612_;
  assign new_n8614_ = new_n3860_;
  assign new_n8615_ = new_n3869_;
  assign new_n8616_ = new_n3867_;
  assign new_n8617_ = new_n3868_;
  assign new_n8618_ = new_n3866_;
  assign new_n8619_ = new_n3871_;
  assign new_n8620_ = new_n8619_;
  assign new_n8621_ = new_n3870_;
  assign new_n8622_ = new_n2913_;
  assign new_n8623_ = new_n8622_;
  assign new_n8624_ = new_n2962_;
  assign new_n8625_ = new_n8624_;
  assign new_n8626_ = new_n3011_;
  assign new_n8627_ = new_n8626_;
  assign new_n8628_ = new_n3120_;
  assign new_n8629_ = new_n8628_;
  assign new_n8630_ = new_n3789_;
  assign new_n8631_ = new_n3714_;
  assign new_n8632_ = new_n3898_;
  assign new_n8633_ = new_n3896_;
  assign new_n8634_ = new_n3897_;
  assign new_n8635_ = new_n3895_;
  assign new_n8636_ = new_n3900_;
  assign new_n8637_ = new_n8636_;
  assign new_n8638_ = new_n3899_;
  assign new_n8639_ = new_n8638_;
  assign new_n8640_ = new_n3908_;
  assign new_n8641_ = new_n3906_;
  assign new_n8642_ = new_n3907_;
  assign new_n8643_ = new_n3905_;
  assign new_n8644_ = new_n3910_;
  assign new_n8645_ = new_n8644_;
  assign new_n8646_ = new_n3909_;
  assign new_n8647_ = new_n8646_;
  assign new_n8648_ = new_n3927_;
  assign new_n8649_ = new_n3925_;
  assign new_n8650_ = new_n3926_;
  assign new_n8651_ = new_n3924_;
  assign new_n8652_ = new_n3929_;
  assign new_n8653_ = new_n8652_;
  assign new_n8654_ = new_n3928_;
  assign new_n8655_ = new_n8654_;
  assign new_n8656_ = new_n3937_;
  assign new_n8657_ = new_n3935_;
  assign new_n8658_ = new_n3936_;
  assign new_n8659_ = new_n3934_;
  assign new_n8660_ = new_n3939_;
  assign new_n8661_ = new_n8660_;
  assign new_n8662_ = new_n3938_;
  assign new_n8663_ = new_n8662_;
  assign new_n8664_ = new_n3947_;
  assign new_n8665_ = new_n3945_;
  assign new_n8666_ = new_n3946_;
  assign new_n8667_ = new_n3944_;
  assign new_n8668_ = new_n3949_;
  assign new_n8669_ = new_n8668_;
  assign new_n8670_ = new_n3948_;
  assign new_n8671_ = new_n8670_;
  assign new_n8672_ = new_n3957_;
  assign new_n8673_ = new_n3955_;
  assign new_n8674_ = new_n3956_;
  assign new_n8675_ = new_n3954_;
  assign new_n8676_ = new_n3959_;
  assign new_n8677_ = new_n8676_;
  assign new_n8678_ = new_n3958_;
  assign new_n8679_ = new_n8678_;
  assign new_n8680_ = new_n3976_;
  assign new_n8681_ = new_n3974_;
  assign new_n8682_ = new_n3975_;
  assign new_n8683_ = new_n3973_;
  assign new_n8684_ = new_n3978_;
  assign new_n8685_ = new_n8684_;
  assign new_n8686_ = new_n3977_;
  assign new_n8687_ = new_n8686_;
  assign new_n8688_ = new_n3986_;
  assign new_n8689_ = new_n3984_;
  assign new_n8690_ = new_n3985_;
  assign new_n8691_ = new_n3983_;
  assign new_n8692_ = new_n3988_;
  assign new_n8693_ = new_n8692_;
  assign new_n8694_ = new_n3987_;
  assign new_n8695_ = new_n8694_;
  assign new_n8696_ = new_n3996_;
  assign new_n8697_ = new_n3994_;
  assign new_n8698_ = new_n3995_;
  assign new_n8699_ = new_n3993_;
  assign new_n8700_ = new_n3998_;
  assign new_n8701_ = new_n8700_;
  assign new_n8702_ = new_n3997_;
  assign new_n8703_ = new_n8702_;
  assign new_n8704_ = new_n4006_;
  assign new_n8705_ = new_n4004_;
  assign new_n8706_ = new_n4005_;
  assign new_n8707_ = new_n4003_;
  assign new_n8708_ = new_n4008_;
  assign new_n8709_ = new_n8708_;
  assign new_n8710_ = new_n4007_;
  assign new_n8711_ = new_n8710_;
  assign new_n8712_ = new_n4037_;
  assign new_n8713_ = new_n4035_;
  assign new_n8714_ = new_n4036_;
  assign new_n8715_ = new_n4034_;
  assign new_n8716_ = new_n4039_;
  assign new_n8717_ = new_n8716_;
  assign new_n8718_ = new_n4038_;
  assign new_n8719_ = new_n8718_;
  assign new_n8720_ = new_n4047_;
  assign new_n8721_ = new_n4045_;
  assign new_n8722_ = new_n4046_;
  assign new_n8723_ = new_n4044_;
  assign new_n8724_ = new_n4049_;
  assign new_n8725_ = new_n8724_;
  assign new_n8726_ = new_n4048_;
  assign new_n8727_ = new_n8726_;
  assign new_n8728_ = new_n4051_;
  assign new_n8729_ = new_n4029_;
  assign new_n8730_ = new_n4050_;
  assign new_n8731_ = new_n4028_;
  assign new_n8732_ = new_n4053_;
  assign new_n8733_ = new_n8732_;
  assign new_n8734_ = new_n4052_;
  assign new_n8735_ = new_n8734_;
  assign new_n8736_ = new_n4061_;
  assign new_n8737_ = new_n4059_;
  assign new_n8738_ = new_n4060_;
  assign new_n8739_ = new_n4058_;
  assign new_n8740_ = new_n4063_;
  assign new_n8741_ = new_n8740_;
  assign new_n8742_ = new_n4062_;
  assign new_n8743_ = new_n8742_;
  assign new_n8744_ = new_n4065_;
  assign new_n8745_ = new_n4023_;
  assign new_n8746_ = new_n4064_;
  assign new_n8747_ = new_n4022_;
  assign new_n8748_ = new_n4067_;
  assign new_n8749_ = new_n8748_;
  assign new_n8750_ = new_n4066_;
  assign new_n8751_ = new_n8750_;
  assign new_n8752_ = new_n4075_;
  assign new_n8753_ = new_n4073_;
  assign new_n8754_ = new_n4074_;
  assign new_n8755_ = new_n4072_;
  assign new_n8756_ = new_n4077_;
  assign new_n8757_ = new_n8756_;
  assign new_n8758_ = new_n4076_;
  assign new_n8759_ = new_n8758_;
  assign new_n8760_ = new_n4097_;
  assign new_n8761_ = new_n4095_;
  assign new_n8762_ = new_n4096_;
  assign new_n8763_ = new_n4094_;
  assign new_n8764_ = new_n4099_;
  assign new_n8765_ = new_n8764_;
  assign new_n8766_ = new_n4098_;
  assign new_n8767_ = new_n8766_;
  assign new_n8768_ = new_n4107_;
  assign new_n8769_ = new_n4105_;
  assign new_n8770_ = new_n4106_;
  assign new_n8771_ = new_n4104_;
  assign new_n8772_ = new_n4109_;
  assign new_n8773_ = new_n8772_;
  assign new_n8774_ = new_n4108_;
  assign new_n8775_ = new_n8774_;
  assign new_n8776_ = new_n4111_;
  assign new_n8777_ = new_n4089_;
  assign new_n8778_ = new_n4110_;
  assign new_n8779_ = new_n4088_;
  assign new_n8780_ = new_n4113_;
  assign new_n8781_ = new_n8780_;
  assign new_n8782_ = new_n4112_;
  assign new_n8783_ = new_n8782_;
  assign new_n8784_ = new_n4121_;
  assign new_n8785_ = new_n4119_;
  assign new_n8786_ = new_n4120_;
  assign new_n8787_ = new_n4118_;
  assign new_n8788_ = new_n4123_;
  assign new_n8789_ = new_n8788_;
  assign new_n8790_ = new_n4122_;
  assign new_n8791_ = new_n8790_;
  assign new_n8792_ = new_n1185_;
  assign new_n8793_ = new_n8792_;
  assign new_n8794_ = new_n8793_;
  assign new_n8795_ = new_n8792_;
  assign new_n8796_ = new_n1186_;
  assign new_n8797_ = new_n8796_;
  assign new_n8798_ = new_n4130_;
  assign new_n8799_ = new_n4128_;
  assign new_n8800_ = new_n4129_;
  assign new_n8801_ = new_n4127_;
  assign new_n8802_ = new_n4132_;
  assign new_n8803_ = new_n8802_;
  assign new_n8804_ = new_n4131_;
  assign new_n8805_ = new_n8804_;
  assign new_n8806_ = new_n1195_;
  assign new_n8807_ = new_n8806_;
  assign new_n8808_ = new_n8806_;
  assign new_n8809_ = new_n1196_;
  assign new_n8810_ = new_n8809_;
  assign new_n8811_ = new_n4140_;
  assign new_n8812_ = new_n4138_;
  assign new_n8813_ = new_n4139_;
  assign new_n8814_ = new_n4137_;
  assign new_n8815_ = new_n4142_;
  assign new_n8816_ = new_n8815_;
  assign new_n8817_ = new_n4141_;
  assign new_n8818_ = new_n8817_;
  assign new_n8819_ = new_n1604_;
  assign new_n8820_ = new_n1566_;
  assign new_n8821_ = new_n1603_;
  assign new_n8822_ = new_n1565_;
  assign new_n8823_ = new_n4150_;
  assign new_n8824_ = new_n8823_;
  assign new_n8825_ = new_n4149_;
  assign new_n8826_ = new_n8825_;
  assign new_n8827_ = new_n1203_;
  assign new_n8828_ = new_n8827_;
  assign new_n8829_ = new_n8827_;
  assign new_n8830_ = new_n1204_;
  assign new_n8831_ = new_n8830_;
  assign new_n8832_ = new_n4158_;
  assign new_n8833_ = new_n4156_;
  assign new_n8834_ = new_n4157_;
  assign new_n8835_ = new_n4155_;
  assign new_n8836_ = new_n4160_;
  assign new_n8837_ = new_n8836_;
  assign new_n8838_ = new_n4159_;
  assign new_n8839_ = new_n8838_;
  assign new_n8840_ = new_n4162_;
  assign new_n8841_ = new_n4148_;
  assign new_n8842_ = new_n4161_;
  assign new_n8843_ = new_n4147_;
  assign new_n8844_ = new_n4164_;
  assign new_n8845_ = new_n8844_;
  assign new_n8846_ = new_n4163_;
  assign new_n8847_ = new_n8846_;
  assign new_n8848_ = new_n4172_;
  assign new_n8849_ = new_n4170_;
  assign new_n8850_ = new_n4171_;
  assign new_n8851_ = new_n4169_;
  assign new_n8852_ = new_n4174_;
  assign new_n8853_ = new_n8852_;
  assign new_n8854_ = new_n4173_;
  assign new_n8855_ = new_n8854_;
  assign new_n8856_ = new_n1207_;
  assign new_n8857_ = new_n8856_;
  assign new_n8858_ = new_n8856_;
  assign new_n8859_ = new_n1208_;
  assign new_n8860_ = new_n8859_;
  assign new_n8861_ = new_n8859_;
  assign new_n8862_ = new_n4190_;
  assign new_n8863_ = new_n4188_;
  assign new_n8864_ = new_n4189_;
  assign new_n8865_ = new_n4187_;
  assign new_n8866_ = new_n4192_;
  assign new_n8867_ = new_n8866_;
  assign new_n8868_ = new_n4191_;
  assign new_n8869_ = new_n8868_;
  assign new_n8870_ = new_n4194_;
  assign new_n8871_ = new_n4186_;
  assign new_n8872_ = new_n4193_;
  assign new_n8873_ = new_n4185_;
  assign new_n8874_ = new_n4196_;
  assign new_n8875_ = new_n8874_;
  assign new_n8876_ = new_n4195_;
  assign new_n8877_ = new_n8876_;
  assign new_n8878_ = new_n4204_;
  assign new_n8879_ = new_n4202_;
  assign new_n8880_ = new_n4203_;
  assign new_n8881_ = new_n4201_;
  assign new_n8882_ = new_n4206_;
  assign new_n8883_ = new_n8882_;
  assign new_n8884_ = new_n4205_;
  assign new_n8885_ = new_n8884_;
  assign new_n8886_ = new_n4208_;
  assign new_n8887_ = new_n4180_;
  assign new_n8888_ = new_n4207_;
  assign new_n8889_ = new_n4179_;
  assign new_n8890_ = new_n4210_;
  assign new_n8891_ = new_n8890_;
  assign new_n8892_ = new_n4209_;
  assign new_n8893_ = new_n8892_;
  assign new_n8894_ = new_n897_;
  assign new_n8895_ = new_n8894_;
  assign new_n8896_ = new_n8895_;
  assign new_n8897_ = new_n8896_;
  assign new_n8898_ = new_n8896_;
  assign new_n8899_ = new_n8895_;
  assign new_n8900_ = new_n8899_;
  assign new_n8901_ = new_n8899_;
  assign new_n8902_ = new_n8894_;
  assign new_n8903_ = new_n8902_;
  assign new_n8904_ = new_n8903_;
  assign new_n8905_ = new_n8903_;
  assign new_n8906_ = new_n8902_;
  assign new_n8907_ = new_n8906_;
  assign new_n8908_ = new_n898_;
  assign new_n8909_ = new_n8908_;
  assign new_n8910_ = new_n8909_;
  assign new_n8911_ = new_n8910_;
  assign new_n8912_ = new_n8910_;
  assign new_n8913_ = new_n8909_;
  assign new_n8914_ = new_n8913_;
  assign new_n8915_ = new_n8913_;
  assign new_n8916_ = new_n8908_;
  assign new_n8917_ = new_n8916_;
  assign new_n8918_ = new_n8917_;
  assign new_n8919_ = new_n8917_;
  assign new_n8920_ = new_n8916_;
  assign new_n8921_ = new_n8920_;
  assign new_n8922_ = new_n4218_;
  assign new_n8923_ = new_n4216_;
  assign new_n8924_ = new_n4217_;
  assign new_n8925_ = new_n4215_;
  assign new_n8926_ = new_n4220_;
  assign new_n8927_ = new_n8926_;
  assign new_n8928_ = new_n4219_;
  assign new_n8929_ = new_n8928_;
  assign new_n8930_ = new_n1601_;
  assign new_n8931_ = new_n8930_;
  assign new_n8932_ = new_n1602_;
  assign new_n8933_ = new_n8932_;
  assign new_n8934_ = new_n1209_;
  assign new_n8935_ = new_n8934_;
  assign new_n8936_ = new_n8935_;
  assign new_n8937_ = new_n8934_;
  assign new_n8938_ = new_n1210_;
  assign new_n8939_ = new_n8938_;
  assign new_n8940_ = new_n8938_;
  assign new_n8941_ = new_n4246_;
  assign new_n8942_ = new_n4244_;
  assign new_n8943_ = new_n4245_;
  assign new_n8944_ = new_n4243_;
  assign new_n8945_ = new_n4248_;
  assign new_n8946_ = new_n8945_;
  assign new_n8947_ = new_n4247_;
  assign new_n8948_ = new_n8947_;
  assign new_n8949_ = new_n4250_;
  assign new_n8950_ = new_n4238_;
  assign new_n8951_ = new_n4249_;
  assign new_n8952_ = new_n4237_;
  assign new_n8953_ = new_n4252_;
  assign new_n8954_ = new_n8953_;
  assign new_n8955_ = new_n4251_;
  assign new_n8956_ = new_n8955_;
  assign new_n8957_ = new_n4260_;
  assign new_n8958_ = new_n4258_;
  assign new_n8959_ = new_n4259_;
  assign new_n8960_ = new_n4257_;
  assign new_n8961_ = new_n4262_;
  assign new_n8962_ = new_n8961_;
  assign new_n8963_ = new_n4261_;
  assign new_n8964_ = new_n8963_;
  assign new_n8965_ = new_n4264_;
  assign new_n8966_ = new_n4232_;
  assign new_n8967_ = new_n4263_;
  assign new_n8968_ = new_n4231_;
  assign new_n8969_ = new_n4266_;
  assign new_n8970_ = new_n8969_;
  assign new_n8971_ = new_n4265_;
  assign new_n8972_ = new_n8971_;
  assign new_n8973_ = new_n4274_;
  assign new_n8974_ = new_n4272_;
  assign new_n8975_ = new_n4273_;
  assign new_n8976_ = new_n4271_;
  assign new_n8977_ = new_n4276_;
  assign new_n8978_ = new_n8977_;
  assign new_n8979_ = new_n4275_;
  assign new_n8980_ = new_n8979_;
  assign new_n8981_ = new_n4278_;
  assign new_n8982_ = new_n4226_;
  assign new_n8983_ = new_n4277_;
  assign new_n8984_ = new_n4225_;
  assign new_n8985_ = new_n3287_;
  assign new_n8986_ = new_n8985_;
  assign new_n8987_ = new_n3286_;
  assign new_n8988_ = new_n3435_;
  assign new_n8989_ = new_n8988_;
  assign new_n8990_ = new_n3434_;
  assign new_n8991_ = new_n3655_;
  assign new_n8992_ = new_n8991_;
  assign new_n8993_ = new_n3654_;
  assign new_n8994_ = new_n917_;
  assign new_n8995_ = new_n8994_;
  assign new_n8996_ = new_n8994_;
  assign new_n8997_ = new_n918_;
  assign new_n8998_ = new_n8997_;
  assign new_n8999_ = new_n8997_;
  assign new_n9000_ = new_n4321_;
  assign new_n9001_ = new_n4319_;
  assign new_n9002_ = new_n4320_;
  assign new_n9003_ = new_n4318_;
  assign new_n9004_ = new_n4323_;
  assign new_n9005_ = new_n9004_;
  assign new_n9006_ = new_n4322_;
  assign new_n9007_ = new_n9006_;
  assign new_n9008_ = new_n4331_;
  assign new_n9009_ = new_n4329_;
  assign new_n9010_ = new_n4330_;
  assign new_n9011_ = new_n4328_;
  assign new_n9012_ = new_n4333_;
  assign new_n9013_ = new_n9012_;
  assign new_n9014_ = new_n4332_;
  assign new_n9015_ = new_n9014_;
  assign new_n9016_ = new_n845_;
  assign new_n9017_ = new_n9016_;
  assign new_n9018_ = new_n9017_;
  assign new_n9019_ = new_n9018_;
  assign new_n9020_ = new_n9018_;
  assign new_n9021_ = new_n9017_;
  assign new_n9022_ = new_n9021_;
  assign new_n9023_ = new_n9021_;
  assign new_n9024_ = new_n9016_;
  assign new_n9025_ = new_n9024_;
  assign new_n9026_ = new_n9025_;
  assign new_n9027_ = new_n9024_;
  assign new_n9028_ = new_n839_;
  assign new_n9029_ = new_n9028_;
  assign new_n9030_ = new_n9028_;
  assign new_n9031_ = new_n846_;
  assign new_n9032_ = new_n9031_;
  assign new_n9033_ = new_n9032_;
  assign new_n9034_ = new_n9033_;
  assign new_n9035_ = new_n9033_;
  assign new_n9036_ = new_n9032_;
  assign new_n9037_ = new_n9036_;
  assign new_n9038_ = new_n9036_;
  assign new_n9039_ = new_n9031_;
  assign new_n9040_ = new_n9039_;
  assign new_n9041_ = new_n9039_;
  assign new_n9042_ = new_n840_;
  assign new_n9043_ = new_n9042_;
  assign new_n9044_ = new_n843_;
  assign new_n9045_ = new_n9044_;
  assign new_n9046_ = new_n9045_;
  assign new_n9047_ = new_n9046_;
  assign new_n9048_ = new_n9046_;
  assign new_n9049_ = new_n9045_;
  assign new_n9050_ = new_n9049_;
  assign new_n9051_ = new_n9049_;
  assign new_n9052_ = new_n9044_;
  assign new_n9053_ = new_n9052_;
  assign new_n9054_ = new_n9053_;
  assign new_n9055_ = new_n9053_;
  assign new_n9056_ = new_n9052_;
  assign new_n9057_ = new_n9056_;
  assign new_n9058_ = new_n844_;
  assign new_n9059_ = new_n9058_;
  assign new_n9060_ = new_n9059_;
  assign new_n9061_ = new_n9060_;
  assign new_n9062_ = new_n9060_;
  assign new_n9063_ = new_n9059_;
  assign new_n9064_ = new_n9063_;
  assign new_n9065_ = new_n9063_;
  assign new_n9066_ = new_n9058_;
  assign new_n9067_ = new_n9066_;
  assign new_n9068_ = new_n9067_;
  assign new_n9069_ = new_n9067_;
  assign new_n9070_ = new_n9066_;
  assign new_n9071_ = new_n9070_;
  assign new_n9072_ = new_n9070_;
  assign new_n9073_ = new_n841_;
  assign new_n9074_ = new_n9073_;
  assign new_n9075_ = new_n9074_;
  assign new_n9076_ = new_n9075_;
  assign new_n9077_ = new_n9075_;
  assign new_n9078_ = new_n9074_;
  assign new_n9079_ = new_n9078_;
  assign new_n9080_ = new_n9078_;
  assign new_n9081_ = new_n9073_;
  assign new_n9082_ = new_n9081_;
  assign new_n9083_ = new_n9082_;
  assign new_n9084_ = new_n9082_;
  assign new_n9085_ = new_n9081_;
  assign new_n9086_ = new_n9085_;
  assign new_n9087_ = new_n9085_;
  assign new_n9088_ = new_n842_;
  assign new_n9089_ = new_n9088_;
  assign new_n9090_ = new_n9089_;
  assign new_n9091_ = new_n9090_;
  assign new_n9092_ = new_n9090_;
  assign new_n9093_ = new_n9089_;
  assign new_n9094_ = new_n9093_;
  assign new_n9095_ = new_n9093_;
  assign new_n9096_ = new_n9088_;
  assign new_n9097_ = new_n9096_;
  assign new_n9098_ = new_n9097_;
  assign new_n9099_ = new_n9097_;
  assign new_n9100_ = new_n9096_;
  assign new_n9101_ = new_n9100_;
  assign new_n9102_ = new_n837_;
  assign new_n9103_ = new_n9102_;
  assign new_n9104_ = new_n9103_;
  assign new_n9105_ = new_n9102_;
  assign new_n9106_ = new_n838_;
  assign new_n9107_ = new_n9106_;
  assign new_n9108_ = new_n9106_;
  assign new_n9109_ = new_n4345_;
  assign new_n9110_ = new_n4342_;
  assign new_n9111_ = new_n4344_;
  assign new_n9112_ = new_n4343_;
  assign new_n9113_ = new_n4347_;
  assign new_n9114_ = new_n4346_;
  assign new_n9115_ = new_n4349_;
  assign new_n9116_ = new_n9115_;
  assign new_n9117_ = new_n4341_;
  assign new_n9118_ = new_n4348_;
  assign new_n9119_ = new_n9118_;
  assign new_n9120_ = new_n4340_;
  assign new_n9121_ = new_n4351_;
  assign new_n9122_ = new_n9121_;
  assign new_n9123_ = new_n4350_;
  assign new_n9124_ = new_n9123_;
  assign new_n9125_ = new_n4359_;
  assign new_n9126_ = new_n4357_;
  assign new_n9127_ = new_n4358_;
  assign new_n9128_ = new_n4356_;
  assign new_n9129_ = new_n4361_;
  assign new_n9130_ = new_n9129_;
  assign new_n9131_ = new_n4360_;
  assign new_n9132_ = new_n9131_;
  assign new_n9133_ = new_n4363_;
  assign new_n9134_ = new_n4339_;
  assign new_n9135_ = new_n4362_;
  assign new_n9136_ = new_n4338_;
  assign new_n9137_ = new_n4369_;
  assign new_n9138_ = new_n4367_;
  assign new_n9139_ = new_n4368_;
  assign new_n9140_ = new_n4366_;
  assign new_n9141_ = new_n4371_;
  assign new_n9142_ = new_n9141_;
  assign new_n9143_ = new_n4370_;
  assign new_n9144_ = new_n9143_;
  assign new_n9145_ = new_n4379_;
  assign new_n9146_ = new_n4377_;
  assign new_n9147_ = new_n4378_;
  assign new_n9148_ = new_n4376_;
  assign new_n9149_ = new_n4381_;
  assign new_n9150_ = new_n9149_;
  assign new_n9151_ = new_n4380_;
  assign new_n9152_ = new_n9151_;
  assign new_n9153_ = new_n4389_;
  assign new_n9154_ = new_n4387_;
  assign new_n9155_ = new_n4388_;
  assign new_n9156_ = new_n4386_;
  assign new_n9157_ = new_n4391_;
  assign new_n9158_ = new_n9157_;
  assign new_n9159_ = new_n4390_;
  assign new_n9160_ = new_n9159_;
  assign new_n9161_ = new_n4399_;
  assign new_n9162_ = new_n4397_;
  assign new_n9163_ = new_n4398_;
  assign new_n9164_ = new_n4396_;
  assign new_n9165_ = new_n4401_;
  assign new_n9166_ = new_n9165_;
  assign new_n9167_ = new_n4400_;
  assign new_n9168_ = new_n9167_;
  assign new_n9169_ = new_n1229_;
  assign new_n9170_ = new_n9169_;
  assign new_n9171_ = new_n9170_;
  assign new_n9172_ = new_n9170_;
  assign new_n9173_ = new_n9169_;
  assign new_n9174_ = new_n9173_;
  assign new_n9175_ = new_n1230_;
  assign new_n9176_ = new_n9175_;
  assign new_n9177_ = new_n9176_;
  assign new_n9178_ = new_n9175_;
  assign new_n9179_ = new_n4414_;
  assign new_n9180_ = new_n4412_;
  assign new_n9181_ = new_n4413_;
  assign new_n9182_ = new_n4411_;
  assign new_n9183_ = new_n4416_;
  assign new_n9184_ = new_n9183_;
  assign new_n9185_ = new_n4415_;
  assign new_n9186_ = new_n9185_;
  assign new_n9187_ = new_n1599_;
  assign new_n9188_ = new_n9187_;
  assign new_n9189_ = new_n1600_;
  assign new_n9190_ = new_n9189_;
  assign new_n9191_ = new_n1253_;
  assign new_n9192_ = new_n9191_;
  assign new_n9193_ = new_n9192_;
  assign new_n9194_ = new_n9192_;
  assign new_n9195_ = new_n9191_;
  assign new_n9196_ = new_n1254_;
  assign new_n9197_ = new_n9196_;
  assign new_n9198_ = new_n9197_;
  assign new_n9199_ = new_n9196_;
  assign new_n9200_ = new_n4430_;
  assign new_n9201_ = new_n4428_;
  assign new_n9202_ = new_n4429_;
  assign new_n9203_ = new_n4427_;
  assign new_n9204_ = new_n4432_;
  assign new_n9205_ = new_n9204_;
  assign new_n9206_ = new_n4431_;
  assign new_n9207_ = new_n9206_;
  assign new_n9208_ = new_n4434_;
  assign new_n9209_ = new_n4422_;
  assign new_n9210_ = new_n4433_;
  assign new_n9211_ = new_n4421_;
  assign new_n9212_ = new_n4436_;
  assign new_n9213_ = new_n9212_;
  assign new_n9214_ = new_n4435_;
  assign new_n9215_ = new_n9214_;
  assign new_n9216_ = new_n4444_;
  assign new_n9217_ = new_n4442_;
  assign new_n9218_ = new_n4443_;
  assign new_n9219_ = new_n4441_;
  assign new_n9220_ = new_n4446_;
  assign new_n9221_ = new_n9220_;
  assign new_n9222_ = new_n4445_;
  assign new_n9223_ = new_n9222_;
  assign new_n9224_ = new_n1610_;
  assign new_n9225_ = new_n1570_;
  assign new_n9226_ = new_n1609_;
  assign new_n9227_ = new_n1569_;
  assign new_n9228_ = new_n4460_;
  assign new_n9229_ = new_n9228_;
  assign new_n9230_ = new_n4459_;
  assign new_n9231_ = new_n9230_;
  assign new_n9232_ = new_n1263_;
  assign new_n9233_ = new_n9232_;
  assign new_n9234_ = new_n9233_;
  assign new_n9235_ = new_n9233_;
  assign new_n9236_ = new_n9232_;
  assign new_n9237_ = new_n1264_;
  assign new_n9238_ = new_n9237_;
  assign new_n9239_ = new_n9238_;
  assign new_n9240_ = new_n9237_;
  assign new_n9241_ = new_n4468_;
  assign new_n9242_ = new_n4466_;
  assign new_n9243_ = new_n4467_;
  assign new_n9244_ = new_n4465_;
  assign new_n9245_ = new_n4470_;
  assign new_n9246_ = new_n9245_;
  assign new_n9247_ = new_n4469_;
  assign new_n9248_ = new_n9247_;
  assign new_n9249_ = new_n4472_;
  assign new_n9250_ = new_n4458_;
  assign new_n9251_ = new_n4471_;
  assign new_n9252_ = new_n4457_;
  assign new_n9253_ = new_n4474_;
  assign new_n9254_ = new_n9253_;
  assign new_n9255_ = new_n4473_;
  assign new_n9256_ = new_n9255_;
  assign new_n9257_ = new_n4482_;
  assign new_n9258_ = new_n4480_;
  assign new_n9259_ = new_n4481_;
  assign new_n9260_ = new_n4479_;
  assign new_n9261_ = new_n4484_;
  assign new_n9262_ = new_n9261_;
  assign new_n9263_ = new_n4483_;
  assign new_n9264_ = new_n9263_;
  assign new_n9265_ = new_n4486_;
  assign new_n9266_ = new_n4452_;
  assign new_n9267_ = new_n4485_;
  assign new_n9268_ = new_n4451_;
  assign new_n9269_ = new_n4488_;
  assign new_n9270_ = new_n9269_;
  assign new_n9271_ = new_n4487_;
  assign new_n9272_ = new_n9271_;
  assign new_n9273_ = new_n4496_;
  assign new_n9274_ = new_n4494_;
  assign new_n9275_ = new_n4495_;
  assign new_n9276_ = new_n4493_;
  assign new_n9277_ = new_n4498_;
  assign new_n9278_ = new_n9277_;
  assign new_n9279_ = new_n4497_;
  assign new_n9280_ = new_n9279_;
  assign new_n9281_ = new_n1596_;
  assign new_n9282_ = new_n9281_;
  assign new_n9283_ = new_n1595_;
  assign new_n9284_ = new_n9283_;
  assign new_n9285_ = new_n4520_;
  assign new_n9286_ = new_n4518_;
  assign new_n9287_ = new_n4519_;
  assign new_n9288_ = new_n4517_;
  assign new_n9289_ = new_n4522_;
  assign new_n9290_ = new_n9289_;
  assign new_n9291_ = new_n4521_;
  assign new_n9292_ = new_n9291_;
  assign new_n9293_ = new_n1265_;
  assign new_n9294_ = new_n9293_;
  assign new_n9295_ = new_n9294_;
  assign new_n9296_ = new_n9294_;
  assign new_n9297_ = new_n9293_;
  assign new_n9298_ = new_n1266_;
  assign new_n9299_ = new_n9298_;
  assign new_n9300_ = new_n9299_;
  assign new_n9301_ = new_n9298_;
  assign new_n9302_ = new_n4530_;
  assign new_n9303_ = new_n4528_;
  assign new_n9304_ = new_n4529_;
  assign new_n9305_ = new_n4527_;
  assign new_n9306_ = new_n4532_;
  assign new_n9307_ = new_n9306_;
  assign new_n9308_ = new_n4531_;
  assign new_n9309_ = new_n9308_;
  assign new_n9310_ = new_n4534_;
  assign new_n9311_ = new_n4516_;
  assign new_n9312_ = new_n4533_;
  assign new_n9313_ = new_n4515_;
  assign new_n9314_ = new_n4536_;
  assign new_n9315_ = new_n9314_;
  assign new_n9316_ = new_n4535_;
  assign new_n9317_ = new_n9316_;
  assign new_n9318_ = new_n4544_;
  assign new_n9319_ = new_n4542_;
  assign new_n9320_ = new_n4543_;
  assign new_n9321_ = new_n4541_;
  assign new_n9322_ = new_n4546_;
  assign new_n9323_ = new_n9322_;
  assign new_n9324_ = new_n4545_;
  assign new_n9325_ = new_n9324_;
  assign new_n9326_ = new_n4548_;
  assign new_n9327_ = new_n4510_;
  assign new_n9328_ = new_n4547_;
  assign new_n9329_ = new_n4509_;
  assign new_n9330_ = new_n4550_;
  assign new_n9331_ = new_n9330_;
  assign new_n9332_ = new_n4549_;
  assign new_n9333_ = new_n9332_;
  assign new_n9334_ = new_n4558_;
  assign new_n9335_ = new_n4556_;
  assign new_n9336_ = new_n4557_;
  assign new_n9337_ = new_n4555_;
  assign new_n9338_ = new_n4560_;
  assign new_n9339_ = new_n9338_;
  assign new_n9340_ = new_n4559_;
  assign new_n9341_ = new_n9340_;
  assign new_n9342_ = new_n4562_;
  assign new_n9343_ = new_n4504_;
  assign new_n9344_ = new_n4561_;
  assign new_n9345_ = new_n4503_;
  assign new_n9346_ = new_n4564_;
  assign new_n9347_ = new_n9346_;
  assign new_n9348_ = new_n4563_;
  assign new_n9349_ = new_n9348_;
  assign new_n9350_ = new_n4572_;
  assign new_n9351_ = new_n4570_;
  assign new_n9352_ = new_n4571_;
  assign new_n9353_ = new_n4569_;
  assign new_n9354_ = new_n4574_;
  assign new_n9355_ = new_n9354_;
  assign new_n9356_ = new_n4573_;
  assign new_n9357_ = new_n9356_;
  assign new_n9358_ = new_n4606_;
  assign new_n9359_ = new_n4604_;
  assign new_n9360_ = new_n4605_;
  assign new_n9361_ = new_n4603_;
  assign new_n9362_ = new_n4608_;
  assign new_n9363_ = new_n9362_;
  assign new_n9364_ = new_n4607_;
  assign new_n9365_ = new_n9364_;
  assign new_n9366_ = new_n1267_;
  assign new_n9367_ = new_n9366_;
  assign new_n9368_ = new_n9367_;
  assign new_n9369_ = new_n9366_;
  assign new_n9370_ = new_n1268_;
  assign new_n9371_ = new_n9370_;
  assign new_n9372_ = new_n9371_;
  assign new_n9373_ = new_n9370_;
  assign new_n9374_ = new_n4616_;
  assign new_n9375_ = new_n4614_;
  assign new_n9376_ = new_n4615_;
  assign new_n9377_ = new_n4613_;
  assign new_n9378_ = new_n4618_;
  assign new_n9379_ = new_n9378_;
  assign new_n9380_ = new_n4617_;
  assign new_n9381_ = new_n9380_;
  assign new_n9382_ = new_n4620_;
  assign new_n9383_ = new_n4598_;
  assign new_n9384_ = new_n4619_;
  assign new_n9385_ = new_n4597_;
  assign new_n9386_ = new_n4622_;
  assign new_n9387_ = new_n9386_;
  assign new_n9388_ = new_n4621_;
  assign new_n9389_ = new_n9388_;
  assign new_n9390_ = new_n4630_;
  assign new_n9391_ = new_n4628_;
  assign new_n9392_ = new_n4629_;
  assign new_n9393_ = new_n4627_;
  assign new_n9394_ = new_n4632_;
  assign new_n9395_ = new_n9394_;
  assign new_n9396_ = new_n4631_;
  assign new_n9397_ = new_n9396_;
  assign new_n9398_ = new_n4634_;
  assign new_n9399_ = new_n4592_;
  assign new_n9400_ = new_n4633_;
  assign new_n9401_ = new_n4591_;
  assign new_n9402_ = new_n4636_;
  assign new_n9403_ = new_n9402_;
  assign new_n9404_ = new_n4635_;
  assign new_n9405_ = new_n9404_;
  assign new_n9406_ = new_n4644_;
  assign new_n9407_ = new_n4642_;
  assign new_n9408_ = new_n4643_;
  assign new_n9409_ = new_n4641_;
  assign new_n9410_ = new_n4646_;
  assign new_n9411_ = new_n9410_;
  assign new_n9412_ = new_n4645_;
  assign new_n9413_ = new_n9412_;
  assign new_n9414_ = new_n4648_;
  assign new_n9415_ = new_n4586_;
  assign new_n9416_ = new_n4647_;
  assign new_n9417_ = new_n4585_;
  assign new_n9418_ = new_n4650_;
  assign new_n9419_ = new_n9418_;
  assign new_n9420_ = new_n4649_;
  assign new_n9421_ = new_n9420_;
  assign new_n9422_ = new_n4658_;
  assign new_n9423_ = new_n4656_;
  assign new_n9424_ = new_n4657_;
  assign new_n9425_ = new_n4655_;
  assign new_n9426_ = new_n4660_;
  assign new_n9427_ = new_n9426_;
  assign new_n9428_ = new_n4659_;
  assign new_n9429_ = new_n9428_;
  assign new_n9430_ = new_n1608_;
  assign new_n9431_ = new_n1572_;
  assign new_n9432_ = new_n1607_;
  assign new_n9433_ = new_n1571_;
  assign new_n9434_ = new_n4677_;
  assign new_n9435_ = new_n9434_;
  assign new_n9436_ = new_n4676_;
  assign new_n9437_ = new_n9436_;
  assign new_n9438_ = new_n1223_;
  assign new_n9439_ = new_n9438_;
  assign new_n9440_ = new_n9439_;
  assign new_n9441_ = new_n9438_;
  assign new_n9442_ = new_n1224_;
  assign new_n9443_ = new_n9442_;
  assign new_n9444_ = new_n9442_;
  assign new_n9445_ = new_n4685_;
  assign new_n9446_ = new_n4683_;
  assign new_n9447_ = new_n4684_;
  assign new_n9448_ = new_n4682_;
  assign new_n9449_ = new_n4687_;
  assign new_n9450_ = new_n9449_;
  assign new_n9451_ = new_n4686_;
  assign new_n9452_ = new_n9451_;
  assign new_n9453_ = new_n4689_;
  assign new_n9454_ = new_n4675_;
  assign new_n9455_ = new_n4688_;
  assign new_n9456_ = new_n4674_;
  assign new_n9457_ = new_n4691_;
  assign new_n9458_ = new_n9457_;
  assign new_n9459_ = new_n4690_;
  assign new_n9460_ = new_n9459_;
  assign new_n9461_ = new_n4699_;
  assign new_n9462_ = new_n4697_;
  assign new_n9463_ = new_n4698_;
  assign new_n9464_ = new_n4696_;
  assign new_n9465_ = new_n4701_;
  assign new_n9466_ = new_n9465_;
  assign new_n9467_ = new_n4700_;
  assign new_n9468_ = new_n9467_;
  assign new_n9469_ = new_n4703_;
  assign new_n9470_ = new_n4669_;
  assign new_n9471_ = new_n4702_;
  assign new_n9472_ = new_n4668_;
  assign new_n9473_ = new_n4705_;
  assign new_n9474_ = new_n9473_;
  assign new_n9475_ = new_n4704_;
  assign new_n9476_ = new_n9475_;
  assign new_n9477_ = new_n4713_;
  assign new_n9478_ = new_n4711_;
  assign new_n9479_ = new_n4712_;
  assign new_n9480_ = new_n4710_;
  assign new_n9481_ = new_n4715_;
  assign new_n9482_ = new_n9481_;
  assign new_n9483_ = new_n4714_;
  assign new_n9484_ = new_n9483_;
  assign new_n9485_ = new_n1594_;
  assign new_n9486_ = new_n9485_;
  assign new_n9487_ = new_n1593_;
  assign new_n9488_ = new_n9487_;
  assign new_n9489_ = new_n4737_;
  assign new_n9490_ = new_n4735_;
  assign new_n9491_ = new_n4736_;
  assign new_n9492_ = new_n4734_;
  assign new_n9493_ = new_n4739_;
  assign new_n9494_ = new_n9493_;
  assign new_n9495_ = new_n4738_;
  assign new_n9496_ = new_n9495_;
  assign new_n9497_ = new_n1225_;
  assign new_n9498_ = new_n9497_;
  assign new_n9499_ = new_n9498_;
  assign new_n9500_ = new_n9497_;
  assign new_n9501_ = new_n1226_;
  assign new_n9502_ = new_n9501_;
  assign new_n9503_ = new_n9501_;
  assign new_n9504_ = new_n4747_;
  assign new_n9505_ = new_n4745_;
  assign new_n9506_ = new_n4746_;
  assign new_n9507_ = new_n4744_;
  assign new_n9508_ = new_n4749_;
  assign new_n9509_ = new_n9508_;
  assign new_n9510_ = new_n4748_;
  assign new_n9511_ = new_n9510_;
  assign new_n9512_ = new_n4751_;
  assign new_n9513_ = new_n4733_;
  assign new_n9514_ = new_n4750_;
  assign new_n9515_ = new_n4732_;
  assign new_n9516_ = new_n4753_;
  assign new_n9517_ = new_n9516_;
  assign new_n9518_ = new_n4752_;
  assign new_n9519_ = new_n9518_;
  assign new_n9520_ = new_n4761_;
  assign new_n9521_ = new_n4759_;
  assign new_n9522_ = new_n4760_;
  assign new_n9523_ = new_n4758_;
  assign new_n9524_ = new_n4763_;
  assign new_n9525_ = new_n9524_;
  assign new_n9526_ = new_n4762_;
  assign new_n9527_ = new_n9526_;
  assign new_n9528_ = new_n4765_;
  assign new_n9529_ = new_n4727_;
  assign new_n9530_ = new_n4764_;
  assign new_n9531_ = new_n4726_;
  assign new_n9532_ = new_n4767_;
  assign new_n9533_ = new_n9532_;
  assign new_n9534_ = new_n4766_;
  assign new_n9535_ = new_n9534_;
  assign new_n9536_ = new_n4775_;
  assign new_n9537_ = new_n4773_;
  assign new_n9538_ = new_n4774_;
  assign new_n9539_ = new_n4772_;
  assign new_n9540_ = new_n4777_;
  assign new_n9541_ = new_n9540_;
  assign new_n9542_ = new_n4776_;
  assign new_n9543_ = new_n9542_;
  assign new_n9544_ = new_n4779_;
  assign new_n9545_ = new_n4721_;
  assign new_n9546_ = new_n4778_;
  assign new_n9547_ = new_n4720_;
  assign new_n9548_ = new_n4781_;
  assign new_n9549_ = new_n9548_;
  assign new_n9550_ = new_n4780_;
  assign new_n9551_ = new_n9550_;
  assign new_n9552_ = new_n899_;
  assign new_n9553_ = new_n9552_;
  assign new_n9554_ = new_n9553_;
  assign new_n9555_ = new_n9554_;
  assign new_n9556_ = new_n9554_;
  assign new_n9557_ = new_n9553_;
  assign new_n9558_ = new_n9552_;
  assign new_n9559_ = new_n9558_;
  assign new_n9560_ = new_n9558_;
  assign new_n9561_ = new_n900_;
  assign new_n9562_ = new_n9561_;
  assign new_n9563_ = new_n9562_;
  assign new_n9564_ = new_n9563_;
  assign new_n9565_ = new_n9563_;
  assign new_n9566_ = new_n9562_;
  assign new_n9567_ = new_n9561_;
  assign new_n9568_ = new_n9567_;
  assign new_n9569_ = new_n9567_;
  assign new_n9570_ = new_n4789_;
  assign new_n9571_ = new_n4787_;
  assign new_n9572_ = new_n4788_;
  assign new_n9573_ = new_n4786_;
  assign new_n9574_ = new_n4791_;
  assign new_n9575_ = new_n9574_;
  assign new_n9576_ = new_n4790_;
  assign new_n9577_ = new_n9576_;
  assign new_n9578_ = new_n1613_;
  assign new_n9579_ = new_n1562_;
  assign new_n9580_ = new_n1614_;
  assign new_n9581_ = new_n1561_;
  assign new_n9582_ = new_n4823_;
  assign new_n9583_ = new_n9582_;
  assign new_n9584_ = new_n4822_;
  assign new_n9585_ = new_n9584_;
  assign new_n9586_ = new_n4825_;
  assign new_n9587_ = new_n4821_;
  assign new_n9588_ = new_n4824_;
  assign new_n9589_ = new_n4820_;
  assign new_n9590_ = new_n4827_;
  assign new_n9591_ = new_n9590_;
  assign new_n9592_ = new_n4826_;
  assign new_n9593_ = new_n9592_;
  assign new_n9594_ = new_n1227_;
  assign new_n9595_ = new_n9594_;
  assign new_n9596_ = new_n9595_;
  assign new_n9597_ = new_n9594_;
  assign new_n9598_ = new_n1228_;
  assign new_n9599_ = new_n9598_;
  assign new_n9600_ = new_n9599_;
  assign new_n9601_ = new_n9598_;
  assign new_n9602_ = new_n4835_;
  assign new_n9603_ = new_n4833_;
  assign new_n9604_ = new_n4834_;
  assign new_n9605_ = new_n4832_;
  assign new_n9606_ = new_n4837_;
  assign new_n9607_ = new_n9606_;
  assign new_n9608_ = new_n4836_;
  assign new_n9609_ = new_n9608_;
  assign new_n9610_ = new_n4839_;
  assign new_n9611_ = new_n4815_;
  assign new_n9612_ = new_n4838_;
  assign new_n9613_ = new_n4814_;
  assign new_n9614_ = new_n4841_;
  assign new_n9615_ = new_n9614_;
  assign new_n9616_ = new_n4840_;
  assign new_n9617_ = new_n9616_;
  assign new_n9618_ = new_n4849_;
  assign new_n9619_ = new_n4847_;
  assign new_n9620_ = new_n4848_;
  assign new_n9621_ = new_n4846_;
  assign new_n9622_ = new_n4851_;
  assign new_n9623_ = new_n9622_;
  assign new_n9624_ = new_n4850_;
  assign new_n9625_ = new_n9624_;
  assign new_n9626_ = new_n4853_;
  assign new_n9627_ = new_n4809_;
  assign new_n9628_ = new_n4852_;
  assign new_n9629_ = new_n4808_;
  assign new_n9630_ = new_n4855_;
  assign new_n9631_ = new_n9630_;
  assign new_n9632_ = new_n4854_;
  assign new_n9633_ = new_n9632_;
  assign new_n9634_ = new_n4863_;
  assign new_n9635_ = new_n4861_;
  assign new_n9636_ = new_n4862_;
  assign new_n9637_ = new_n4860_;
  assign new_n9638_ = new_n4865_;
  assign new_n9639_ = new_n9638_;
  assign new_n9640_ = new_n4864_;
  assign new_n9641_ = new_n9640_;
  assign new_n9642_ = new_n4867_;
  assign new_n9643_ = new_n4803_;
  assign new_n9644_ = new_n4866_;
  assign new_n9645_ = new_n4802_;
  assign new_n9646_ = new_n4869_;
  assign new_n9647_ = new_n9646_;
  assign new_n9648_ = new_n4868_;
  assign new_n9649_ = new_n9648_;
  assign new_n9650_ = new_n4877_;
  assign new_n9651_ = new_n4875_;
  assign new_n9652_ = new_n4876_;
  assign new_n9653_ = new_n4874_;
  assign new_n9654_ = new_n4879_;
  assign new_n9655_ = new_n9654_;
  assign new_n9656_ = new_n4878_;
  assign new_n9657_ = new_n9656_;
  assign new_n9658_ = new_n4890_;
  assign new_n9659_ = new_n4888_;
  assign new_n9660_ = new_n4889_;
  assign new_n9661_ = new_n4887_;
  assign new_n9662_ = new_n4892_;
  assign new_n9663_ = new_n9662_;
  assign new_n9664_ = new_n4891_;
  assign new_n9665_ = new_n9664_;
  assign new_n9666_ = new_n4900_;
  assign new_n9667_ = new_n4898_;
  assign new_n9668_ = new_n4899_;
  assign new_n9669_ = new_n4897_;
  assign new_n9670_ = new_n4902_;
  assign new_n9671_ = new_n9670_;
  assign new_n9672_ = new_n4901_;
  assign new_n9673_ = new_n9672_;
  assign new_n9674_ = new_n4910_;
  assign new_n9675_ = new_n4908_;
  assign new_n9676_ = new_n4909_;
  assign new_n9677_ = new_n4907_;
  assign new_n9678_ = new_n4912_;
  assign new_n9679_ = new_n9678_;
  assign new_n9680_ = new_n4911_;
  assign new_n9681_ = new_n9680_;
  assign new_n9682_ = new_n4920_;
  assign new_n9683_ = new_n4918_;
  assign new_n9684_ = new_n4919_;
  assign new_n9685_ = new_n4917_;
  assign new_n9686_ = new_n4922_;
  assign new_n9687_ = new_n9686_;
  assign new_n9688_ = new_n4921_;
  assign new_n9689_ = new_n9688_;
  assign new_n9690_ = new_n3716_;
  assign new_n9691_ = new_n4930_;
  assign new_n9692_ = new_n4928_;
  assign new_n9693_ = new_n4932_;
  assign new_n9694_ = new_n3822_;
  assign new_n9695_ = new_n9694_;
  assign new_n9696_ = new_n3851_;
  assign new_n9697_ = new_n9696_;
  assign new_n9698_ = new_n3880_;
  assign new_n9699_ = new_n9698_;
  assign new_n9700_ = new_n3889_;
  assign new_n9701_ = new_n3790_;
  assign new_n9702_ = new_n3886_;
  assign new_n9703_ = new_n3791_;
  assign new_n9704_ = new_n3883_;
  assign new_n9705_ = new_n3792_;
  assign new_n9706_ = new_n3892_;
  assign new_n9707_ = new_n3793_;
  assign new_n9708_ = new_n3144_;
  assign new_n9709_ = new_n9708_;
  assign new_n9710_ = new_n3153_;
  assign new_n9711_ = new_n9710_;
  assign new_n9712_ = new_n3162_;
  assign new_n9713_ = new_n9712_;
  assign new_n9714_ = new_n4974_;
  assign new_n9715_ = new_n4972_;
  assign new_n9716_ = new_n4973_;
  assign new_n9717_ = new_n4971_;
  assign new_n9718_ = new_n4976_;
  assign new_n9719_ = new_n9718_;
  assign new_n9720_ = new_n4975_;
  assign new_n9721_ = new_n4984_;
  assign new_n9722_ = new_n4982_;
  assign new_n9723_ = new_n4983_;
  assign new_n9724_ = new_n4981_;
  assign new_n9725_ = new_n4986_;
  assign new_n9726_ = new_n9725_;
  assign new_n9727_ = new_n4985_;
  assign new_n9728_ = new_n5003_;
  assign new_n9729_ = new_n5001_;
  assign new_n9730_ = new_n5002_;
  assign new_n9731_ = new_n5000_;
  assign new_n9732_ = new_n5005_;
  assign new_n9733_ = new_n9732_;
  assign new_n9734_ = new_n5004_;
  assign new_n9735_ = new_n5013_;
  assign new_n9736_ = new_n5011_;
  assign new_n9737_ = new_n5012_;
  assign new_n9738_ = new_n5010_;
  assign new_n9739_ = new_n5015_;
  assign new_n9740_ = new_n9739_;
  assign new_n9741_ = new_n5014_;
  assign new_n9742_ = new_n3893_;
  assign new_n9743_ = new_n3919_;
  assign new_n9744_ = new_n9743_;
  assign new_n9745_ = new_n3968_;
  assign new_n9746_ = new_n9745_;
  assign new_n9747_ = new_n4017_;
  assign new_n9748_ = new_n9747_;
  assign new_n9749_ = new_n4126_;
  assign new_n9750_ = new_n9749_;
  assign new_n9751_ = new_n4280_;
  assign new_n9752_ = new_n9751_;
  assign new_n9753_ = new_n4279_;
  assign new_n9754_ = new_n4935_;
  assign new_n9755_ = new_n4337_;
  assign new_n9756_ = new_n5075_;
  assign new_n9757_ = new_n5073_;
  assign new_n9758_ = new_n5074_;
  assign new_n9759_ = new_n5072_;
  assign new_n9760_ = new_n5077_;
  assign new_n9761_ = new_n9760_;
  assign new_n9762_ = new_n5076_;
  assign new_n9763_ = new_n9762_;
  assign new_n9764_ = new_n5085_;
  assign new_n9765_ = new_n5083_;
  assign new_n9766_ = new_n5084_;
  assign new_n9767_ = new_n5082_;
  assign new_n9768_ = new_n5087_;
  assign new_n9769_ = new_n9768_;
  assign new_n9770_ = new_n5086_;
  assign new_n9771_ = new_n9770_;
  assign new_n9772_ = new_n5089_;
  assign new_n9773_ = new_n5067_;
  assign new_n9774_ = new_n5088_;
  assign new_n9775_ = new_n5066_;
  assign new_n9776_ = new_n5091_;
  assign new_n9777_ = new_n9776_;
  assign new_n9778_ = new_n5090_;
  assign new_n9779_ = new_n9778_;
  assign new_n9780_ = new_n5099_;
  assign new_n9781_ = new_n5097_;
  assign new_n9782_ = new_n5098_;
  assign new_n9783_ = new_n5096_;
  assign new_n9784_ = new_n5101_;
  assign new_n9785_ = new_n9784_;
  assign new_n9786_ = new_n5100_;
  assign new_n9787_ = new_n9786_;
  assign new_n9788_ = new_n5136_;
  assign new_n9789_ = new_n5134_;
  assign new_n9790_ = new_n5135_;
  assign new_n9791_ = new_n5133_;
  assign new_n9792_ = new_n5138_;
  assign new_n9793_ = new_n9792_;
  assign new_n9794_ = new_n5137_;
  assign new_n9795_ = new_n9794_;
  assign new_n9796_ = new_n5146_;
  assign new_n9797_ = new_n5144_;
  assign new_n9798_ = new_n5145_;
  assign new_n9799_ = new_n5143_;
  assign new_n9800_ = new_n5148_;
  assign new_n9801_ = new_n9800_;
  assign new_n9802_ = new_n5147_;
  assign new_n9803_ = new_n9802_;
  assign new_n9804_ = new_n5150_;
  assign new_n9805_ = new_n5128_;
  assign new_n9806_ = new_n5149_;
  assign new_n9807_ = new_n5127_;
  assign new_n9808_ = new_n5152_;
  assign new_n9809_ = new_n9808_;
  assign new_n9810_ = new_n5151_;
  assign new_n9811_ = new_n9810_;
  assign new_n9812_ = new_n5160_;
  assign new_n9813_ = new_n5158_;
  assign new_n9814_ = new_n5159_;
  assign new_n9815_ = new_n5157_;
  assign new_n9816_ = new_n5162_;
  assign new_n9817_ = new_n9816_;
  assign new_n9818_ = new_n5161_;
  assign new_n9819_ = new_n9818_;
  assign new_n9820_ = new_n5164_;
  assign new_n9821_ = new_n5122_;
  assign new_n9822_ = new_n5163_;
  assign new_n9823_ = new_n5121_;
  assign new_n9824_ = new_n5166_;
  assign new_n9825_ = new_n9824_;
  assign new_n9826_ = new_n5165_;
  assign new_n9827_ = new_n9826_;
  assign new_n9828_ = new_n5174_;
  assign new_n9829_ = new_n5172_;
  assign new_n9830_ = new_n5173_;
  assign new_n9831_ = new_n5171_;
  assign new_n9832_ = new_n5176_;
  assign new_n9833_ = new_n9832_;
  assign new_n9834_ = new_n5175_;
  assign new_n9835_ = new_n9834_;
  assign new_n9836_ = new_n5178_;
  assign new_n9837_ = new_n5116_;
  assign new_n9838_ = new_n5177_;
  assign new_n9839_ = new_n5115_;
  assign new_n9840_ = new_n5180_;
  assign new_n9841_ = new_n9840_;
  assign new_n9842_ = new_n5179_;
  assign new_n9843_ = new_n9842_;
  assign new_n9844_ = new_n5188_;
  assign new_n9845_ = new_n5186_;
  assign new_n9846_ = new_n5187_;
  assign new_n9847_ = new_n5185_;
  assign new_n9848_ = new_n5190_;
  assign new_n9849_ = new_n9848_;
  assign new_n9850_ = new_n5189_;
  assign new_n9851_ = new_n9850_;
  assign new_n9852_ = new_n821_;
  assign new_n9853_ = new_n9852_;
  assign new_n9854_ = new_n9852_;
  assign new_n9855_ = new_n822_;
  assign new_n9856_ = new_n9855_;
  assign new_n9857_ = new_n819_;
  assign new_n9858_ = new_n9857_;
  assign new_n9859_ = new_n9857_;
  assign new_n9860_ = new_n820_;
  assign new_n9861_ = new_n9860_;
  assign new_n9862_ = new_n5197_;
  assign new_n9863_ = new_n5194_;
  assign new_n9864_ = new_n5196_;
  assign new_n9865_ = new_n5195_;
  assign new_n9866_ = new_n5199_;
  assign new_n9867_ = new_n5198_;
  assign new_n9868_ = new_n5201_;
  assign new_n9869_ = new_n9868_;
  assign new_n9870_ = new_n5200_;
  assign new_n9871_ = new_n9870_;
  assign new_n9872_ = new_n817_;
  assign new_n9873_ = new_n9872_;
  assign new_n9874_ = new_n818_;
  assign new_n9875_ = new_n9874_;
  assign new_n9876_ = new_n5209_;
  assign new_n9877_ = new_n5206_;
  assign new_n9878_ = new_n5208_;
  assign new_n9879_ = new_n5207_;
  assign new_n9880_ = new_n5211_;
  assign new_n9881_ = new_n5210_;
  assign new_n9882_ = new_n5212_;
  assign new_n9883_ = new_n833_;
  assign new_n9884_ = new_n9883_;
  assign new_n9885_ = new_n9884_;
  assign new_n9886_ = new_n9883_;
  assign new_n9887_ = new_n834_;
  assign new_n9888_ = new_n9887_;
  assign new_n9889_ = new_n9887_;
  assign new_n9890_ = new_n831_;
  assign new_n9891_ = new_n9890_;
  assign new_n9892_ = new_n9891_;
  assign new_n9893_ = new_n9890_;
  assign new_n9894_ = new_n832_;
  assign new_n9895_ = new_n9894_;
  assign new_n9896_ = new_n9894_;
  assign new_n9897_ = new_n5218_;
  assign new_n9898_ = new_n5215_;
  assign new_n9899_ = new_n5217_;
  assign new_n9900_ = new_n5216_;
  assign new_n9901_ = new_n5220_;
  assign new_n9902_ = new_n5219_;
  assign new_n9903_ = new_n5222_;
  assign new_n9904_ = new_n9903_;
  assign new_n9905_ = new_n5221_;
  assign new_n9906_ = new_n9905_;
  assign new_n9907_ = new_n829_;
  assign new_n9908_ = new_n9907_;
  assign new_n9909_ = new_n9908_;
  assign new_n9910_ = new_n9907_;
  assign new_n9911_ = new_n830_;
  assign new_n9912_ = new_n9911_;
  assign new_n9913_ = new_n9911_;
  assign new_n9914_ = new_n5230_;
  assign new_n9915_ = new_n5227_;
  assign new_n9916_ = new_n5229_;
  assign new_n9917_ = new_n5228_;
  assign new_n9918_ = new_n5232_;
  assign new_n9919_ = new_n5231_;
  assign new_n9920_ = new_n5234_;
  assign new_n9921_ = new_n9920_;
  assign new_n9922_ = new_n5226_;
  assign new_n9923_ = new_n5233_;
  assign new_n9924_ = new_n9923_;
  assign new_n9925_ = new_n5225_;
  assign new_n9926_ = new_n5236_;
  assign new_n9927_ = new_n9926_;
  assign new_n9928_ = new_n5235_;
  assign new_n9929_ = new_n9928_;
  assign new_n9930_ = new_n5244_;
  assign new_n9931_ = new_n5242_;
  assign new_n9932_ = new_n5243_;
  assign new_n9933_ = new_n5241_;
  assign new_n9934_ = new_n5246_;
  assign new_n9935_ = new_n9934_;
  assign new_n9936_ = new_n5245_;
  assign new_n9937_ = new_n9936_;
  assign new_n9938_ = new_n827_;
  assign new_n9939_ = new_n9938_;
  assign new_n9940_ = new_n9938_;
  assign new_n9941_ = new_n828_;
  assign new_n9942_ = new_n9941_;
  assign new_n9943_ = new_n9941_;
  assign new_n9944_ = new_n5260_;
  assign new_n9945_ = new_n5257_;
  assign new_n9946_ = new_n5259_;
  assign new_n9947_ = new_n5258_;
  assign new_n9948_ = new_n5262_;
  assign new_n9949_ = new_n5261_;
  assign new_n9950_ = new_n5264_;
  assign new_n9951_ = new_n9950_;
  assign new_n9952_ = new_n5256_;
  assign new_n9953_ = new_n5263_;
  assign new_n9954_ = new_n9953_;
  assign new_n9955_ = new_n5255_;
  assign new_n9956_ = new_n5266_;
  assign new_n9957_ = new_n9956_;
  assign new_n9958_ = new_n5265_;
  assign new_n9959_ = new_n9958_;
  assign new_n9960_ = new_n5274_;
  assign new_n9961_ = new_n5272_;
  assign new_n9962_ = new_n5273_;
  assign new_n9963_ = new_n5271_;
  assign new_n9964_ = new_n5276_;
  assign new_n9965_ = new_n9964_;
  assign new_n9966_ = new_n5275_;
  assign new_n9967_ = new_n9966_;
  assign new_n9968_ = new_n5294_;
  assign new_n9969_ = new_n5292_;
  assign new_n9970_ = new_n5293_;
  assign new_n9971_ = new_n5291_;
  assign new_n9972_ = new_n5296_;
  assign new_n9973_ = new_n9972_;
  assign new_n9974_ = new_n5295_;
  assign new_n9975_ = new_n5305_;
  assign new_n9976_ = new_n9975_;
  assign new_n9977_ = new_n5055_;
  assign new_n9978_ = new_n5321_;
  assign new_n9979_ = new_n5319_;
  assign new_n9980_ = new_n5320_;
  assign new_n9981_ = new_n5318_;
  assign new_n9982_ = new_n5323_;
  assign new_n9983_ = new_n9982_;
  assign new_n9984_ = new_n5322_;
  assign new_n9985_ = new_n9984_;
  assign new_n9986_ = new_n5331_;
  assign new_n9987_ = new_n5329_;
  assign new_n9988_ = new_n5330_;
  assign new_n9989_ = new_n5328_;
  assign new_n9990_ = new_n5333_;
  assign new_n9991_ = new_n9990_;
  assign new_n9992_ = new_n5332_;
  assign new_n9993_ = new_n9992_;
  assign new_n9994_ = new_n5335_;
  assign new_n9995_ = new_n5313_;
  assign new_n9996_ = new_n5334_;
  assign new_n9997_ = new_n5312_;
  assign new_n9998_ = new_n5337_;
  assign new_n9999_ = new_n9998_;
  assign new_n10000_ = new_n5336_;
  assign new_n10001_ = new_n10000_;
  assign new_n10002_ = new_n5345_;
  assign new_n10003_ = new_n5343_;
  assign new_n10004_ = new_n5344_;
  assign new_n10005_ = new_n5342_;
  assign new_n10006_ = new_n5347_;
  assign new_n10007_ = new_n10006_;
  assign new_n10008_ = new_n5346_;
  assign new_n10009_ = new_n10008_;
  assign new_n10010_ = new_n5361_;
  assign new_n10011_ = new_n5359_;
  assign new_n10012_ = new_n5360_;
  assign new_n10013_ = new_n5358_;
  assign new_n10014_ = new_n5363_;
  assign new_n10015_ = new_n10014_;
  assign new_n10016_ = new_n5362_;
  assign new_n10017_ = new_n10016_;
  assign new_n10018_ = new_n5371_;
  assign new_n10019_ = new_n5369_;
  assign new_n10020_ = new_n5370_;
  assign new_n10021_ = new_n5368_;
  assign new_n10022_ = new_n5373_;
  assign new_n10023_ = new_n10022_;
  assign new_n10024_ = new_n5372_;
  assign new_n10025_ = new_n10024_;
  assign new_n10026_ = new_n5375_;
  assign new_n10027_ = new_n5353_;
  assign new_n10028_ = new_n5374_;
  assign new_n10029_ = new_n5352_;
  assign new_n10030_ = new_n5377_;
  assign new_n10031_ = new_n10030_;
  assign new_n10032_ = new_n5376_;
  assign new_n10033_ = new_n5386_;
  assign new_n10034_ = new_n10033_;
  assign new_n10035_ = new_n4966_;
  assign new_n10036_ = new_n10035_;
  assign new_n10037_ = new_n4995_;
  assign new_n10038_ = new_n10037_;
  assign new_n10039_ = new_n5024_;
  assign new_n10040_ = new_n10039_;
  assign new_n10041_ = new_n5033_;
  assign new_n10042_ = new_n10041_;
  assign new_n10043_ = new_n5036_;
  assign new_n10044_ = new_n4936_;
  assign new_n10045_ = new_n5039_;
  assign new_n10046_ = new_n4937_;
  assign new_n10047_ = new_n5042_;
  assign new_n10048_ = new_n4938_;
  assign new_n10049_ = new_n5045_;
  assign new_n10050_ = new_n4939_;
  assign new_n10051_ = new_n4365_;
  assign new_n10052_ = new_n10051_;
  assign new_n10053_ = new_n4364_;
  assign new_n10054_ = new_n847_;
  assign new_n10055_ = new_n10054_;
  assign new_n10056_ = new_n10055_;
  assign new_n10057_ = new_n10055_;
  assign new_n10058_ = new_n10054_;
  assign new_n10059_ = new_n10058_;
  assign new_n10060_ = new_n848_;
  assign new_n10061_ = new_n10060_;
  assign new_n10062_ = new_n10061_;
  assign new_n10063_ = new_n10061_;
  assign new_n10064_ = new_n10060_;
  assign new_n10065_ = new_n5414_;
  assign new_n10066_ = new_n5412_;
  assign new_n10067_ = new_n5413_;
  assign new_n10068_ = new_n5411_;
  assign new_n10069_ = new_n5416_;
  assign new_n10070_ = new_n10069_;
  assign new_n10071_ = new_n5415_;
  assign new_n10072_ = new_n5424_;
  assign new_n10073_ = new_n5422_;
  assign new_n10074_ = new_n5423_;
  assign new_n10075_ = new_n5421_;
  assign new_n10076_ = new_n5426_;
  assign new_n10077_ = new_n10076_;
  assign new_n10078_ = new_n5425_;
  assign new_n10079_ = new_n5443_;
  assign new_n10080_ = new_n5441_;
  assign new_n10081_ = new_n5442_;
  assign new_n10082_ = new_n5440_;
  assign new_n10083_ = new_n5445_;
  assign new_n10084_ = new_n10083_;
  assign new_n10085_ = new_n5444_;
  assign new_n10086_ = new_n5453_;
  assign new_n10087_ = new_n5451_;
  assign new_n10088_ = new_n5452_;
  assign new_n10089_ = new_n5450_;
  assign new_n10090_ = new_n5455_;
  assign new_n10091_ = new_n10090_;
  assign new_n10092_ = new_n5454_;
  assign new_n10093_ = new_n5478_;
  assign new_n10094_ = new_n5476_;
  assign new_n10095_ = new_n5477_;
  assign new_n10096_ = new_n5475_;
  assign new_n10097_ = new_n5480_;
  assign new_n10098_ = new_n10097_;
  assign new_n10099_ = new_n5479_;
  assign new_n10100_ = new_n10099_;
  assign new_n10101_ = new_n5488_;
  assign new_n10102_ = new_n5486_;
  assign new_n10103_ = new_n5490_;
  assign new_n10104_ = new_n10103_;
  assign new_n10105_ = new_n5507_;
  assign new_n10106_ = new_n5505_;
  assign new_n10107_ = new_n5506_;
  assign new_n10108_ = new_n5504_;
  assign new_n10109_ = new_n5509_;
  assign new_n10110_ = new_n10109_;
  assign new_n10111_ = new_n5508_;
  assign new_n10112_ = new_n10111_;
  assign new_n10113_ = new_n5516_;
  assign new_n10114_ = new_n5514_;
  assign new_n10115_ = new_n5518_;
  assign new_n10116_ = new_n10115_;
  assign new_n10117_ = new_n4289_;
  assign new_n10118_ = new_n10117_;
  assign new_n10119_ = new_n4298_;
  assign new_n10120_ = new_n10119_;
  assign new_n10121_ = new_n4307_;
  assign new_n10122_ = new_n10121_;
  assign new_n10123_ = new_n4336_;
  assign new_n10124_ = new_n10123_;
  assign new_n10125_ = new_n5213_;
  assign new_n10126_ = new_n815_;
  assign new_n10127_ = new_n10126_;
  assign new_n10128_ = new_n10126_;
  assign new_n10129_ = new_n816_;
  assign new_n10130_ = new_n5542_;
  assign new_n10131_ = new_n5539_;
  assign new_n10132_ = new_n5541_;
  assign new_n10133_ = new_n5540_;
  assign new_n10134_ = new_n5544_;
  assign new_n10135_ = new_n5543_;
  assign new_n10136_ = new_n5545_;
  assign new_n10137_ = new_n825_;
  assign new_n10138_ = new_n10137_;
  assign new_n10139_ = new_n10138_;
  assign new_n10140_ = new_n10137_;
  assign new_n10141_ = new_n826_;
  assign new_n10142_ = new_n10141_;
  assign new_n10143_ = new_n5561_;
  assign new_n10144_ = new_n5558_;
  assign new_n10145_ = new_n5560_;
  assign new_n10146_ = new_n5559_;
  assign new_n10147_ = new_n5563_;
  assign new_n10148_ = new_n5562_;
  assign new_n10149_ = new_n5565_;
  assign new_n10150_ = new_n10149_;
  assign new_n10151_ = new_n5557_;
  assign new_n10152_ = new_n5564_;
  assign new_n10153_ = new_n10152_;
  assign new_n10154_ = new_n5556_;
  assign new_n10155_ = new_n5567_;
  assign new_n10156_ = new_n10155_;
  assign new_n10157_ = new_n5566_;
  assign new_n10158_ = new_n10157_;
  assign new_n10159_ = new_n5575_;
  assign new_n10160_ = new_n5573_;
  assign new_n10161_ = new_n5574_;
  assign new_n10162_ = new_n5572_;
  assign new_n10163_ = new_n5577_;
  assign new_n10164_ = new_n10163_;
  assign new_n10165_ = new_n5576_;
  assign new_n10166_ = new_n10165_;
  assign new_n10167_ = new_n4410_;
  assign new_n10168_ = new_n10167_;
  assign new_n10169_ = new_n4663_;
  assign new_n10170_ = new_n10169_;
  assign new_n10171_ = new_n4882_;
  assign new_n10172_ = new_n10171_;
  assign new_n10173_ = new_n811_;
  assign new_n10174_ = new_n10173_;
  assign new_n10175_ = new_n812_;
  assign new_n10176_ = new_n901_;
  assign new_n10177_ = new_n5612_;
  assign new_n10178_ = new_n5610_;
  assign new_n10179_ = new_n5611_;
  assign new_n10180_ = new_n5609_;
  assign new_n10181_ = new_n5614_;
  assign new_n10182_ = new_n10181_;
  assign new_n10183_ = new_n5613_;
  assign new_n10184_ = new_n5623_;
  assign new_n10185_ = new_n10184_;
  assign new_n10186_ = new_n813_;
  assign new_n10187_ = new_n10186_;
  assign new_n10188_ = new_n814_;
  assign new_n10189_ = new_n5629_;
  assign new_n10190_ = new_n823_;
  assign new_n10191_ = new_n10190_;
  assign new_n10192_ = new_n10190_;
  assign new_n10193_ = new_n824_;
  assign new_n10194_ = new_n10193_;
  assign new_n10195_ = new_n5634_;
  assign new_n10196_ = new_n5631_;
  assign new_n10197_ = new_n5633_;
  assign new_n10198_ = new_n5632_;
  assign new_n10199_ = new_n5636_;
  assign new_n10200_ = new_n5635_;
  assign new_n10201_ = new_n5638_;
  assign new_n10202_ = new_n10201_;
  assign new_n10203_ = new_n5637_;
  assign new_n10204_ = new_n10203_;
  assign new_n10205_ = new_n5646_;
  assign new_n10206_ = new_n5643_;
  assign new_n10207_ = new_n5645_;
  assign new_n10208_ = new_n5644_;
  assign new_n10209_ = new_n5648_;
  assign new_n10210_ = new_n5647_;
  assign new_n10211_ = new_n5650_;
  assign new_n10212_ = new_n10211_;
  assign new_n10213_ = new_n5642_;
  assign new_n10214_ = new_n5649_;
  assign new_n10215_ = new_n10214_;
  assign new_n10216_ = new_n5641_;
  assign new_n10217_ = new_n5652_;
  assign new_n10218_ = new_n10217_;
  assign new_n10219_ = new_n5651_;
  assign new_n10220_ = new_n5661_;
  assign new_n10221_ = new_n10220_;
  assign new_n10222_ = new_n835_;
  assign new_n10223_ = new_n10222_;
  assign new_n10224_ = new_n10223_;
  assign new_n10225_ = new_n10222_;
  assign new_n10226_ = new_n836_;
  assign new_n10227_ = new_n10226_;
  assign new_n10228_ = new_n10226_;
  assign new_n10229_ = new_n5666_;
  assign new_n10230_ = new_n5663_;
  assign new_n10231_ = new_n5665_;
  assign new_n10232_ = new_n5664_;
  assign new_n10233_ = new_n5668_;
  assign new_n10234_ = new_n5667_;
  assign new_n10235_ = new_n5670_;
  assign new_n10236_ = new_n10235_;
  assign new_n10237_ = new_n5669_;
  assign new_n10238_ = new_n10237_;
  assign new_n10239_ = new_n5678_;
  assign new_n10240_ = new_n5675_;
  assign new_n10241_ = new_n5677_;
  assign new_n10242_ = new_n5676_;
  assign new_n10243_ = new_n5680_;
  assign new_n10244_ = new_n5679_;
  assign new_n10245_ = new_n5682_;
  assign new_n10246_ = new_n10245_;
  assign new_n10247_ = new_n5674_;
  assign new_n10248_ = new_n5681_;
  assign new_n10249_ = new_n10248_;
  assign new_n10250_ = new_n5673_;
  assign new_n10251_ = new_n5684_;
  assign new_n10252_ = new_n10251_;
  assign new_n10253_ = new_n5683_;
  assign new_n10254_ = new_n10253_;
  assign new_n10255_ = new_n5692_;
  assign new_n10256_ = new_n5690_;
  assign new_n10257_ = new_n5691_;
  assign new_n10258_ = new_n5689_;
  assign new_n10259_ = new_n5694_;
  assign new_n10260_ = new_n10259_;
  assign new_n10261_ = new_n5693_;
  assign new_n10262_ = new_n10261_;
  assign new_n10263_ = new_n5704_;
  assign new_n10264_ = new_n5703_;
  assign new_n10265_ = new_n5706_;
  assign new_n10266_ = new_n10265_;
  assign new_n10267_ = new_n5705_;
  assign new_n10268_ = new_n10267_;
  assign new_n10269_ = new_n5714_;
  assign new_n10270_ = new_n5712_;
  assign new_n10271_ = new_n5713_;
  assign new_n10272_ = new_n5711_;
  assign new_n10273_ = new_n5716_;
  assign new_n10274_ = new_n10273_;
  assign new_n10275_ = new_n5715_;
  assign new_n10276_ = new_n10275_;
  assign new_n10277_ = new_n5718_;
  assign new_n10278_ = new_n5700_;
  assign new_n10279_ = new_n5717_;
  assign new_n10280_ = new_n5699_;
  assign new_n10281_ = new_n5720_;
  assign new_n10282_ = new_n10281_;
  assign new_n10283_ = new_n5719_;
  assign new_n10284_ = new_n5729_;
  assign new_n10285_ = new_n10284_;
  assign new_n10286_ = new_n5435_;
  assign new_n10287_ = new_n10286_;
  assign new_n10288_ = new_n5464_;
  assign new_n10289_ = new_n10288_;
  assign new_n10290_ = new_n5493_;
  assign new_n10291_ = new_n10290_;
  assign new_n10292_ = new_n5522_;
  assign new_n10293_ = new_n10292_;
  assign new_n10294_ = new_n5589_;
  assign new_n10295_ = new_n5281_;
  assign new_n10296_ = new_n5595_;
  assign new_n10297_ = new_n5282_;
  assign new_n10298_ = new_n5592_;
  assign new_n10299_ = new_n5283_;
  assign new_n10300_ = new_n5596_;
  assign new_n10301_ = new_n5284_;
  assign new_n10302_ = new_n5586_;
  assign new_n10303_ = new_n5307_;
  assign new_n10304_ = new_n5583_;
  assign new_n10305_ = new_n5387_;
  assign new_n10306_ = new_n5546_;
  assign new_n10307_ = new_n5754_;
  assign new_n10308_ = new_n5751_;
  assign new_n10309_ = new_n5752_;
  assign new_n10310_ = new_n5756_;
  assign new_n10311_ = new_n5757_;
  assign new_n10312_ = new_n5769_;
  assign new_n10313_ = new_n5768_;
  assign new_n10314_ = new_n5771_;
  assign new_n10315_ = new_n10314_;
  assign new_n10316_ = new_n5770_;
  assign new_n10317_ = new_n10316_;
  assign new_n10318_ = new_n5778_;
  assign new_n10319_ = new_n5776_;
  assign new_n10320_ = new_n5780_;
  assign new_n10321_ = new_n10320_;
  assign new_n10322_ = new_n5794_;
  assign new_n10323_ = new_n5793_;
  assign new_n10324_ = new_n5796_;
  assign new_n10325_ = new_n10324_;
  assign new_n10326_ = new_n5795_;
  assign new_n10327_ = new_n10326_;
  assign new_n10328_ = new_n5804_;
  assign new_n10329_ = new_n5802_;
  assign new_n10330_ = new_n5803_;
  assign new_n10331_ = new_n5801_;
  assign new_n10332_ = new_n5806_;
  assign new_n10333_ = new_n10332_;
  assign new_n10334_ = new_n5805_;
  assign new_n10335_ = new_n10334_;
  assign new_n10336_ = new_n5808_;
  assign new_n10337_ = new_n5790_;
  assign new_n10338_ = new_n5807_;
  assign new_n10339_ = new_n5789_;
  assign new_n10340_ = new_n5810_;
  assign new_n10341_ = new_n10340_;
  assign new_n10342_ = new_n5809_;
  assign new_n10343_ = new_n5818_;
  assign new_n10344_ = new_n5816_;
  assign new_n10345_ = new_n5817_;
  assign new_n10346_ = new_n5815_;
  assign new_n10347_ = new_n5820_;
  assign new_n10348_ = new_n10347_;
  assign new_n10349_ = new_n5819_;
  assign new_n10350_ = new_n5834_;
  assign new_n10351_ = new_n5832_;
  assign new_n10352_ = new_n5833_;
  assign new_n10353_ = new_n5831_;
  assign new_n10354_ = new_n5836_;
  assign new_n10355_ = new_n10354_;
  assign new_n10356_ = new_n5835_;
  assign new_n10357_ = new_n10356_;
  assign new_n10358_ = new_n5843_;
  assign new_n10359_ = new_n5841_;
  assign new_n10360_ = new_n5845_;
  assign new_n10361_ = new_n10360_;
  assign new_n10362_ = new_n5054_;
  assign new_n10363_ = new_n10362_;
  assign new_n10364_ = new_n5104_;
  assign new_n10365_ = new_n10364_;
  assign new_n10366_ = new_n5193_;
  assign new_n10367_ = new_n10366_;
  assign new_n10368_ = new_n5214_;
  assign new_n10369_ = new_n10368_;
  assign new_n10370_ = new_n5279_;
  assign new_n10371_ = new_n10370_;
  assign new_n10372_ = new_n5744_;
  assign new_n10373_ = new_n5883_;
  assign new_n10374_ = new_n5882_;
  assign new_n10375_ = new_n5885_;
  assign new_n10376_ = new_n10375_;
  assign new_n10377_ = new_n5884_;
  assign new_n10378_ = new_n5894_;
  assign new_n10379_ = new_n10378_;
  assign new_n10380_ = new_n5903_;
  assign new_n10381_ = new_n5901_;
  assign new_n10382_ = new_n5902_;
  assign new_n10383_ = new_n5900_;
  assign new_n10384_ = new_n5905_;
  assign new_n10385_ = new_n10384_;
  assign new_n10386_ = new_n5904_;
  assign new_n10387_ = new_n5914_;
  assign new_n10388_ = new_n10387_;
  assign new_n10389_ = new_n5759_;
  assign new_n10390_ = new_n10389_;
  assign new_n10391_ = new_n5784_;
  assign new_n10392_ = new_n10391_;
  assign new_n10393_ = new_n5849_;
  assign new_n10394_ = new_n10393_;
  assign new_n10395_ = new_n5875_;
  assign new_n10396_ = new_n5601_;
  assign new_n10397_ = new_n5872_;
  assign new_n10398_ = new_n5602_;
  assign new_n10399_ = new_n5866_;
  assign new_n10400_ = new_n5630_;
  assign new_n10401_ = new_n10400_;
  assign new_n10402_ = new_n5869_;
  assign new_n10403_ = new_n5662_;
  assign new_n10404_ = new_n5864_;
  assign new_n10405_ = new_n5730_;
  assign new_n10406_ = new_n5410_;
  assign new_n10407_ = new_n10406_;
  assign new_n10408_ = new_n5547_;
  assign new_n10409_ = new_n10408_;
  assign new_n10410_ = new_n5580_;
  assign new_n10411_ = new_n10410_;
  always @ (posedge clock) begin
    n2491_lo <= n2491_li;
    n2575_lo <= n2575_li;
    n2587_lo <= n2587_li;
    n2599_lo <= n2599_li;
    n2611_lo <= n2611_li;
    n2623_lo <= n2623_li;
    n2635_lo <= n2635_li;
    n2647_lo <= n2647_li;
    n2659_lo <= n2659_li;
    n2671_lo <= n2671_li;
    n2683_lo <= n2683_li;
    n2734_lo <= n2734_li;
    n2746_lo <= n2746_li;
    n2758_lo <= n2758_li;
    n2770_lo <= n2770_li;
    n2782_lo <= n2782_li;
    n2785_lo <= n2785_li;
    n2794_lo <= n2794_li;
    n2797_lo <= n2797_li;
    n2806_lo <= n2806_li;
    n2809_lo <= n2809_li;
    n2818_lo <= n2818_li;
    n2821_lo <= n2821_li;
    n2830_lo <= n2830_li;
    n2833_lo <= n2833_li;
    n2836_lo <= n2836_li;
    n2839_lo <= n2839_li;
    n2842_lo <= n2842_li;
    n2845_lo <= n2845_li;
    n2848_lo <= n2848_li;
    n2851_lo <= n2851_li;
    n2854_lo <= n2854_li;
    n2857_lo <= n2857_li;
    n2860_lo <= n2860_li;
    n2863_lo <= n2863_li;
    n4871_o2 <= n4871_i2;
    n4893_o2 <= n4893_i2;
    n4938_o2 <= n4938_i2;
    n5056_o2 <= n5056_i2;
    n5100_o2 <= n5100_i2;
    n5122_o2 <= n5122_i2;
    n5254_o2 <= n5254_i2;
    n5276_o2 <= n5276_i2;
    n5316_o2 <= n5316_i2;
    n5434_o2 <= n5434_i2;
    n5473_o2 <= n5473_i2;
    n5494_o2 <= n5494_i2;
    n5620_o2 <= n5620_i2;
    n5643_o2 <= n5643_i2;
    n5682_o2 <= n5682_i2;
    n5798_o2 <= n5798_i2;
    n5839_o2 <= n5839_i2;
    n5867_o2 <= n5867_i2;
    n6052_o2 <= n6052_i2;
    n6087_o2 <= n6087_i2;
    n6153_o2 <= n6153_i2;
    n6408_o2 <= n6408_i2;
    n6454_o2 <= n6454_i2;
    n6509_o2 <= n6509_i2;
    n6775_o2 <= n6775_i2;
    n6818_o2 <= n6818_i2;
    n6892_o2 <= n6892_i2;
    n5779_o2 <= n5779_i2;
    n5780_o2 <= n5780_i2;
    n7156_o2 <= n7156_i2;
    n5792_o2 <= n5792_i2;
    n7205_o2 <= n7205_i2;
    n5842_o2 <= n5842_i2;
    n5863_o2 <= n5863_i2;
    n7263_o2 <= n7263_i2;
    n5881_o2 <= n5881_i2;
    n5930_o2 <= n5930_i2;
    n5959_o2 <= n5959_i2;
    n5981_o2 <= n5981_i2;
    n6042_o2 <= n6042_i2;
    n6075_o2 <= n6075_i2;
    n6103_o2 <= n6103_i2;
    n7610_o2 <= n7610_i2;
    n6169_o2 <= n6169_i2;
    n7665_o2 <= n7665_i2;
    n6205_o2 <= n6205_i2;
    n6239_o2 <= n6239_i2;
    n7788_o2 <= n7788_i2;
    n6309_o2 <= n6309_i2;
    n6461_o2 <= n6461_i2;
    n6476_o2 <= n6476_i2;
    n325_inv <= n6521_i2;
    n6545_o2 <= n6545_i2;
    G578_o2 <= G578_i2;
    G5106_o2 <= G5106_i2;
    n6713_o2 <= n6713_i2;
    G5164_o2 <= G5164_i2;
    n343_inv <= n6771_i2;
    n6810_o2 <= n6810_i2;
    n6973_o2 <= n6973_i2;
    n352_inv <= n6995_i2;
    n7053_o2 <= n7053_i2;
    G581_o2 <= G581_i2;
    G5467_o2 <= G5467_i2;
    n7231_o2 <= n7231_i2;
    G5527_o2 <= G5527_i2;
    n370_inv <= n7277_i2;
    n7304_o2 <= n7304_i2;
    n7530_o2 <= n7530_i2;
    n379_inv <= n7595_i2;
    n7653_o2 <= n7653_i2;
    G584_o2 <= G584_i2;
    G5820_o2 <= G5820_i2;
    n7148_o2 <= n7148_i2;
    n7149_o2 <= n7149_i2;
    n7224_o2 <= n7224_i2;
    n7916_o2 <= n7916_i2;
    G5868_o2 <= G5868_i2;
    n406_inv <= n7958_i2;
    n7280_o2 <= n7280_i2;
    n7313_o2 <= n7313_i2;
    n8056_o2 <= n8056_i2;
    n7323_o2 <= n7323_i2;
    n7398_o2 <= n7398_i2;
    n7459_o2 <= n7459_i2;
    n7501_o2 <= n7501_i2;
    n7518_o2 <= n7518_i2;
    G563_o2 <= G563_i2;
    n7606_o2 <= n7606_i2;
    n439_inv <= G3358_i2;
    n7675_o2 <= n7675_i2;
    G3410_o2 <= G3410_i2;
    n7722_o2 <= n7722_i2;
    n7747_o2 <= n7747_i2;
    n7835_o2 <= n7835_i2;
    G587_o2 <= G587_i2;
    G6046_o2 <= G6046_i2;
    n7909_o2 <= n7909_i2;
    G566_o2 <= G566_i2;
    G6070_o2 <= G6070_i2;
    n472_inv <= G3698_i2;
    n8086_o2 <= n8086_i2;
    n8093_o2 <= n8093_i2;
    G3752_o2 <= G3752_i2;
    n484_inv <= n8156_i2;
    n8199_o2 <= n8199_i2;
    n2800_lo_buf_o2 <= n2800_lo_buf_i2;
    G548_o2 <= G548_i2;
    n496_inv <= G1715_i2;
    G569_o2 <= G569_i2;
    G1761_o2 <= G1761_i2;
    n505_inv <= G4043_i2;
    G4101_o2 <= G4101_i2;
    G551_o2 <= G551_i2;
    n514_inv <= G2034_i2;
    G4743_o2 <= G4743_i2;
    G5271_o2 <= G5271_i2;
    G5790_o2 <= G5790_i2;
    G6122_o2 <= G6122_i2;
    G2082_o2 <= G2082_i2;
    n2812_lo_buf_o2 <= n2812_lo_buf_i2;
    n2668_lo_buf_o2 <= n2668_lo_buf_i2;
    n2680_lo_buf_o2 <= n2680_lo_buf_i2;
    G572_o2 <= G572_i2;
    G6125_o2 <= G6125_i2;
    n547_inv <= G4395_i2;
    n2656_lo_buf_o2 <= n2656_lo_buf_i2;
    G554_o2 <= G554_i2;
    G4452_o2 <= G4452_i2;
    n559_inv <= G2358_i2;
    n2644_lo_buf_o2 <= n2644_lo_buf_i2;
    G2410_o2 <= G2410_i2;
    n2632_lo_buf_o2 <= n2632_lo_buf_i2;
    n2620_lo_buf_o2 <= n2620_lo_buf_i2;
    G6131_o2 <= G6131_i2;
    G4693_o2 <= G4693_i2;
    G5209_o2 <= G5209_i2;
    G5741_o2 <= G5741_i2;
    G6082_o2 <= G6082_i2;
    G6119_o2 <= G6119_i2;
    n2608_lo_buf_o2 <= n2608_lo_buf_i2;
    n2596_lo_buf_o2 <= n2596_lo_buf_i2;
    n2584_lo_buf_o2 <= n2584_lo_buf_i2;
    n2572_lo_buf_o2 <= n2572_lo_buf_i2;
    n2704_lo_buf_o2 <= n2704_lo_buf_i2;
    G557_o2 <= G557_i2;
    G5936_o2 <= G5936_i2;
    G5442_o2 <= G5442_i2;
    G4926_o2 <= G4926_i2;
    G6134_o2 <= G6134_i2;
    G3929_o2 <= G3929_i2;
    G4425_o2 <= G4425_i2;
    G4947_o2 <= G4947_i2;
    n2764_lo_buf_o2 <= n2764_lo_buf_i2;
    n634_inv <= G2689_i2;
    n2560_lo_buf_o2 <= n2560_lo_buf_i2;
    n2824_lo_buf_o2 <= n2824_lo_buf_i2;
    G575_o2 <= G575_i2;
    G2740_o2 <= G2740_i2;
    n649_inv <= G4749_i2;
    n2548_lo_buf_o2 <= n2548_lo_buf_i2;
    n2536_lo_buf_o2 <= n2536_lo_buf_i2;
    n2524_lo_buf_o2 <= n2524_lo_buf_i2;
    G875_o2 <= G875_i2;
    G1064_o2 <= G1064_i2;
    G1253_o2 <= G1253_i2;
    G6140_o2 <= G6140_i2;
    G5151_o2 <= G5151_i2;
    G5686_o2 <= G5686_i2;
    G6061_o2 <= G6061_i2;
    G4803_o2 <= G4803_i2;
    G5332_o2 <= G5332_i2;
    G5844_o2 <= G5844_i2;
    G6114_o2 <= G6114_i2;
    G4806_o2 <= G4806_i2;
    G3881_o2 <= G3881_i2;
    G4370_o2 <= G4370_i2;
    G4896_o2 <= G4896_i2;
    G5001_o2 <= G5001_i2;
    G3121_o2 <= G3121_i2;
    n2512_lo_buf_o2 <= n2512_lo_buf_i2;
    G4085_o2 <= G4085_i2;
    G4605_o2 <= G4605_i2;
    G5118_o2 <= G5118_i2;
    G4997_o2 <= G4997_i2;
    n2500_lo_buf_o2 <= n2500_lo_buf_i2;
    n2716_lo_buf_o2 <= n2716_lo_buf_i2;
    G560_o2 <= G560_i2;
    G1895_o2 <= G1895_i2;
    G3064_o2 <= G3064_i2;
    G3269_o2 <= G3269_i2;
    G3569_o2 <= G3569_i2;
    n748_inv <= G3022_i2;
    G1196_o2 <= G1196_i2;
    G1007_o2 <= G1007_i2;
    G818_o2 <= G818_i2;
    G674_o2 <= G674_i2;
    G5041_o2 <= G5041_i2;
    G5562_o2 <= G5562_i2;
    G6005_o2 <= G6005_i2;
    G5214_o2 <= G5214_i2;
    G5746_o2 <= G5746_i2;
    G6087_o2 <= G6087_i2;
    G6086_o2 <= G6086_i2;
    G5745_o2 <= G5745_i2;
    G5213_o2 <= G5213_i2;
    G5893_o2 <= G5893_i2;
    G5391_o2 <= G5391_i2;
    G4864_o2 <= G4864_i2;
    G6143_o2 <= G6143_i2;
    G6008_o2 <= G6008_i2;
    G5565_o2 <= G5565_i2;
    G5044_o2 <= G5044_i2;
    G3813_o2 <= G3813_i2;
    G4325_o2 <= G4325_i2;
    G4834_o2 <= G4834_i2;
    G4993_o2 <= G4993_i2;
    G3989_o2 <= G3989_i2;
    G4490_o2 <= G4490_i2;
    G5011_o2 <= G5011_i2;
    G5112_o2 <= G5112_i2;
    n2776_lo_buf_o2 <= n2776_lo_buf_i2;
    G3298_o2 <= G3298_i2;
    G3073_o2 <= G3073_i2;
    G3265_o2 <= G3265_i2;
    G3624_o2 <= G3624_i2;
    G1642_o2 <= G1642_i2;
    G1980_o2 <= G1980_i2;
    n2488_lo_buf_o2 <= n2488_lo_buf_i2;
    G626_o2 <= G626_i2;
    G1139_o2 <= G1139_i2;
    G950_o2 <= G950_i2;
    G707_o2 <= G707_i2;
    G545_o2 <= G545_i2;
    G4217_o2 <= G4217_i2;
    G4716_o2 <= G4716_i2;
    G5244_o2 <= G5244_i2;
    G3136_o2 <= G3136_i2;
    G3499_o2 <= G3499_i2;
    G3885_o2 <= G3885_i2;
    G5243_o2 <= G5243_i2;
    G3886_o2 <= G3886_i2;
    G4375_o2 <= G4375_i2;
    G4901_o2 <= G4901_i2;
    G5054_o2 <= G5054_i2;
    G4374_o2 <= G4374_i2;
    G4900_o2 <= G4900_i2;
    G5053_o2 <= G5053_i2;
    G5242_o2 <= G5242_i2;
    G4034_o2 <= G4034_i2;
    G4556_o2 <= G4556_i2;
    G5064_o2 <= G5064_i2;
    G5172_o2 <= G5172_i2;
    G2030_o2 <= G2030_i2;
    G3016_o2 <= G3016_i2;
    G3520_o2 <= G3520_i2;
    G3261_o2 <= G3261_i2;
    G3620_o2 <= G3620_i2;
    G4220_o2 <= G4220_i2;
    G4719_o2 <= G4719_i2;
    G5247_o2 <= G5247_i2;
    G5109_o2 <= G5109_i2;
    G1638_o2 <= G1638_i2;
    G1976_o2 <= G1976_i2;
    G3560_o2 <= G3560_i2;
    G3205_o2 <= G3205_i2;
    G3193_o2 <= G3193_i2;
    G3367_o2 <= G3367_i2;
    G3670_o2 <= G3670_i2;
    n979_inv <= G1400_i2;
    G1280_o2 <= G1280_i2;
    G902_o2 <= G902_i2;
    G659_o2 <= G659_i2;
    G983_o2 <= G983_i2;
    G740_o2 <= G740_i2;
    G2917_o2 <= G2917_i2;
    G3391_o2 <= G3391_i2;
    G3494_o2 <= G3494_i2;
    G1512_o2 <= G1512_i2;
    G1854_o2 <= G1854_i2;
    G2203_o2 <= G2203_i2;
    G3493_o2 <= G3493_i2;
    G3069_o2 <= G3069_i2;
    G3574_o2 <= G3574_i2;
    G3319_o2 <= G3319_i2;
    G3667_o2 <= G3667_i2;
    G3068_o2 <= G3068_i2;
    G3573_o2 <= G3573_i2;
    G3666_o2 <= G3666_i2;
    G3318_o2 <= G3318_i2;
    G3492_o2 <= G3492_i2;
    G3241_o2 <= G3241_i2;
    G3722_o2 <= G3722_i2;
    G3422_o2 <= G3422_i2;
    G1445_o2 <= G1445_i2;
    G3257_o2 <= G3257_i2;
    G3616_o2 <= G3616_i2;
    G1634_o2 <= G1634_i2;
    G1972_o2 <= G1972_i2;
    G2256_o2 <= G2256_i2;
    G3394_o2 <= G3394_i2;
    G3557_o2 <= G3557_i2;
    G3364_o2 <= G3364_i2;
    G3719_o2 <= G3719_i2;
    G2253_o2 <= G2253_i2;
    G1583_o2 <= G1583_i2;
    G1917_o2 <= G1917_i2;
    G1727_o2 <= G1727_i2;
    G2061_o2 <= G2061_i2;
    G935_o2 <= G935_i2;
    G692_o2 <= G692_i2;
    G2136_o2 <= G2136_i2;
    G1507_o2 <= G1507_i2;
    G1849_o2 <= G1849_i2;
    G2198_o2 <= G2198_i2;
    G2197_o2 <= G2197_i2;
    G1848_o2 <= G1848_i2;
    G1689_o2 <= G1689_i2;
    G2016_o2 <= G2016_i2;
    G2314_o2 <= G2314_i2;
    G2313_o2 <= G2313_i2;
    G1688_o2 <= G1688_i2;
    G2015_o2 <= G2015_i2;
    G1847_o2 <= G1847_i2;
    G2196_o2 <= G2196_i2;
    G2118_o2 <= G2118_i2;
    G1777_o2 <= G1777_i2;
    G1630_o2 <= G1630_i2;
    G1968_o2 <= G1968_i2;
    G2309_o2 <= G2309_i2;
    G2139_o2 <= G2139_i2;
    G1580_o2 <= G1580_i2;
    G2250_o2 <= G2250_i2;
    G1914_o2 <= G1914_i2;
    G1724_o2 <= G1724_i2;
    G2058_o2 <= G2058_i2;
    n2728_lo_buf_o2 <= n2728_lo_buf_i2;
  end
  initial begin
    n2491_lo <= 1'b0;
    n2575_lo <= 1'b0;
    n2587_lo <= 1'b0;
    n2599_lo <= 1'b0;
    n2611_lo <= 1'b0;
    n2623_lo <= 1'b0;
    n2635_lo <= 1'b0;
    n2647_lo <= 1'b0;
    n2659_lo <= 1'b0;
    n2671_lo <= 1'b0;
    n2683_lo <= 1'b0;
    n2734_lo <= 1'b0;
    n2746_lo <= 1'b0;
    n2758_lo <= 1'b0;
    n2770_lo <= 1'b0;
    n2782_lo <= 1'b0;
    n2785_lo <= 1'b0;
    n2794_lo <= 1'b0;
    n2797_lo <= 1'b0;
    n2806_lo <= 1'b0;
    n2809_lo <= 1'b0;
    n2818_lo <= 1'b0;
    n2821_lo <= 1'b0;
    n2830_lo <= 1'b0;
    n2833_lo <= 1'b0;
    n2836_lo <= 1'b0;
    n2839_lo <= 1'b0;
    n2842_lo <= 1'b0;
    n2845_lo <= 1'b0;
    n2848_lo <= 1'b0;
    n2851_lo <= 1'b0;
    n2854_lo <= 1'b0;
    n2857_lo <= 1'b0;
    n2860_lo <= 1'b0;
    n2863_lo <= 1'b0;
    n4871_o2 <= 1'b0;
    n4893_o2 <= 1'b0;
    n4938_o2 <= 1'b0;
    n5056_o2 <= 1'b0;
    n5100_o2 <= 1'b0;
    n5122_o2 <= 1'b0;
    n5254_o2 <= 1'b0;
    n5276_o2 <= 1'b0;
    n5316_o2 <= 1'b0;
    n5434_o2 <= 1'b0;
    n5473_o2 <= 1'b0;
    n5494_o2 <= 1'b0;
    n5620_o2 <= 1'b0;
    n5643_o2 <= 1'b0;
    n5682_o2 <= 1'b0;
    n5798_o2 <= 1'b0;
    n5839_o2 <= 1'b0;
    n5867_o2 <= 1'b0;
    n6052_o2 <= 1'b0;
    n6087_o2 <= 1'b0;
    n6153_o2 <= 1'b0;
    n6408_o2 <= 1'b0;
    n6454_o2 <= 1'b0;
    n6509_o2 <= 1'b0;
    n6775_o2 <= 1'b0;
    n6818_o2 <= 1'b0;
    n6892_o2 <= 1'b0;
    n5779_o2 <= 1'b0;
    n5780_o2 <= 1'b0;
    n7156_o2 <= 1'b0;
    n5792_o2 <= 1'b0;
    n7205_o2 <= 1'b0;
    n5842_o2 <= 1'b0;
    n5863_o2 <= 1'b0;
    n7263_o2 <= 1'b0;
    n5881_o2 <= 1'b0;
    n5930_o2 <= 1'b0;
    n5959_o2 <= 1'b0;
    n5981_o2 <= 1'b0;
    n6042_o2 <= 1'b0;
    n6075_o2 <= 1'b0;
    n6103_o2 <= 1'b0;
    n7610_o2 <= 1'b0;
    n6169_o2 <= 1'b0;
    n7665_o2 <= 1'b0;
    n6205_o2 <= 1'b0;
    n6239_o2 <= 1'b0;
    n7788_o2 <= 1'b0;
    n6309_o2 <= 1'b0;
    n6461_o2 <= 1'b0;
    n6476_o2 <= 1'b0;
    n325_inv <= 1'b0;
    n6545_o2 <= 1'b0;
    G578_o2 <= 1'b0;
    G5106_o2 <= 1'b0;
    n6713_o2 <= 1'b0;
    G5164_o2 <= 1'b0;
    n343_inv <= 1'b0;
    n6810_o2 <= 1'b0;
    n6973_o2 <= 1'b0;
    n352_inv <= 1'b0;
    n7053_o2 <= 1'b0;
    G581_o2 <= 1'b0;
    G5467_o2 <= 1'b0;
    n7231_o2 <= 1'b0;
    G5527_o2 <= 1'b0;
    n370_inv <= 1'b0;
    n7304_o2 <= 1'b0;
    n7530_o2 <= 1'b0;
    n379_inv <= 1'b0;
    n7653_o2 <= 1'b0;
    G584_o2 <= 1'b0;
    G5820_o2 <= 1'b0;
    n7148_o2 <= 1'b0;
    n7149_o2 <= 1'b0;
    n7224_o2 <= 1'b0;
    n7916_o2 <= 1'b0;
    G5868_o2 <= 1'b0;
    n406_inv <= 1'b0;
    n7280_o2 <= 1'b0;
    n7313_o2 <= 1'b0;
    n8056_o2 <= 1'b0;
    n7323_o2 <= 1'b0;
    n7398_o2 <= 1'b0;
    n7459_o2 <= 1'b0;
    n7501_o2 <= 1'b0;
    n7518_o2 <= 1'b0;
    G563_o2 <= 1'b0;
    n7606_o2 <= 1'b0;
    n439_inv <= 1'b0;
    n7675_o2 <= 1'b0;
    G3410_o2 <= 1'b0;
    n7722_o2 <= 1'b0;
    n7747_o2 <= 1'b0;
    n7835_o2 <= 1'b0;
    G587_o2 <= 1'b0;
    G6046_o2 <= 1'b0;
    n7909_o2 <= 1'b0;
    G566_o2 <= 1'b0;
    G6070_o2 <= 1'b0;
    n472_inv <= 1'b0;
    n8086_o2 <= 1'b0;
    n8093_o2 <= 1'b0;
    G3752_o2 <= 1'b0;
    n484_inv <= 1'b0;
    n8199_o2 <= 1'b0;
    n2800_lo_buf_o2 <= 1'b0;
    G548_o2 <= 1'b0;
    n496_inv <= 1'b0;
    G569_o2 <= 1'b0;
    G1761_o2 <= 1'b0;
    n505_inv <= 1'b0;
    G4101_o2 <= 1'b0;
    G551_o2 <= 1'b0;
    n514_inv <= 1'b0;
    G4743_o2 <= 1'b0;
    G5271_o2 <= 1'b0;
    G5790_o2 <= 1'b0;
    G6122_o2 <= 1'b0;
    G2082_o2 <= 1'b0;
    n2812_lo_buf_o2 <= 1'b0;
    n2668_lo_buf_o2 <= 1'b0;
    n2680_lo_buf_o2 <= 1'b0;
    G572_o2 <= 1'b0;
    G6125_o2 <= 1'b0;
    n547_inv <= 1'b0;
    n2656_lo_buf_o2 <= 1'b0;
    G554_o2 <= 1'b0;
    G4452_o2 <= 1'b0;
    n559_inv <= 1'b0;
    n2644_lo_buf_o2 <= 1'b0;
    G2410_o2 <= 1'b0;
    n2632_lo_buf_o2 <= 1'b0;
    n2620_lo_buf_o2 <= 1'b0;
    G6131_o2 <= 1'b0;
    G4693_o2 <= 1'b0;
    G5209_o2 <= 1'b0;
    G5741_o2 <= 1'b0;
    G6082_o2 <= 1'b0;
    G6119_o2 <= 1'b0;
    n2608_lo_buf_o2 <= 1'b0;
    n2596_lo_buf_o2 <= 1'b0;
    n2584_lo_buf_o2 <= 1'b0;
    n2572_lo_buf_o2 <= 1'b0;
    n2704_lo_buf_o2 <= 1'b0;
    G557_o2 <= 1'b0;
    G5936_o2 <= 1'b0;
    G5442_o2 <= 1'b0;
    G4926_o2 <= 1'b0;
    G6134_o2 <= 1'b0;
    G3929_o2 <= 1'b0;
    G4425_o2 <= 1'b0;
    G4947_o2 <= 1'b0;
    n2764_lo_buf_o2 <= 1'b0;
    n634_inv <= 1'b0;
    n2560_lo_buf_o2 <= 1'b0;
    n2824_lo_buf_o2 <= 1'b0;
    G575_o2 <= 1'b0;
    G2740_o2 <= 1'b0;
    n649_inv <= 1'b0;
    n2548_lo_buf_o2 <= 1'b0;
    n2536_lo_buf_o2 <= 1'b0;
    n2524_lo_buf_o2 <= 1'b0;
    G875_o2 <= 1'b0;
    G1064_o2 <= 1'b0;
    G1253_o2 <= 1'b0;
    G6140_o2 <= 1'b0;
    G5151_o2 <= 1'b0;
    G5686_o2 <= 1'b0;
    G6061_o2 <= 1'b0;
    G4803_o2 <= 1'b0;
    G5332_o2 <= 1'b0;
    G5844_o2 <= 1'b0;
    G6114_o2 <= 1'b0;
    G4806_o2 <= 1'b0;
    G3881_o2 <= 1'b0;
    G4370_o2 <= 1'b0;
    G4896_o2 <= 1'b0;
    G5001_o2 <= 1'b0;
    G3121_o2 <= 1'b0;
    n2512_lo_buf_o2 <= 1'b0;
    G4085_o2 <= 1'b0;
    G4605_o2 <= 1'b0;
    G5118_o2 <= 1'b0;
    G4997_o2 <= 1'b0;
    n2500_lo_buf_o2 <= 1'b0;
    n2716_lo_buf_o2 <= 1'b0;
    G560_o2 <= 1'b0;
    G1895_o2 <= 1'b0;
    G3064_o2 <= 1'b0;
    G3269_o2 <= 1'b0;
    G3569_o2 <= 1'b0;
    n748_inv <= 1'b0;
    G1196_o2 <= 1'b0;
    G1007_o2 <= 1'b0;
    G818_o2 <= 1'b0;
    G674_o2 <= 1'b0;
    G5041_o2 <= 1'b0;
    G5562_o2 <= 1'b0;
    G6005_o2 <= 1'b0;
    G5214_o2 <= 1'b0;
    G5746_o2 <= 1'b0;
    G6087_o2 <= 1'b0;
    G6086_o2 <= 1'b0;
    G5745_o2 <= 1'b0;
    G5213_o2 <= 1'b0;
    G5893_o2 <= 1'b0;
    G5391_o2 <= 1'b0;
    G4864_o2 <= 1'b0;
    G6143_o2 <= 1'b0;
    G6008_o2 <= 1'b0;
    G5565_o2 <= 1'b0;
    G5044_o2 <= 1'b0;
    G3813_o2 <= 1'b0;
    G4325_o2 <= 1'b0;
    G4834_o2 <= 1'b0;
    G4993_o2 <= 1'b0;
    G3989_o2 <= 1'b0;
    G4490_o2 <= 1'b0;
    G5011_o2 <= 1'b0;
    G5112_o2 <= 1'b0;
    n2776_lo_buf_o2 <= 1'b0;
    G3298_o2 <= 1'b0;
    G3073_o2 <= 1'b0;
    G3265_o2 <= 1'b0;
    G3624_o2 <= 1'b0;
    G1642_o2 <= 1'b0;
    G1980_o2 <= 1'b0;
    n2488_lo_buf_o2 <= 1'b0;
    G626_o2 <= 1'b0;
    G1139_o2 <= 1'b0;
    G950_o2 <= 1'b0;
    G707_o2 <= 1'b0;
    G545_o2 <= 1'b0;
    G4217_o2 <= 1'b0;
    G4716_o2 <= 1'b0;
    G5244_o2 <= 1'b0;
    G3136_o2 <= 1'b0;
    G3499_o2 <= 1'b0;
    G3885_o2 <= 1'b0;
    G5243_o2 <= 1'b0;
    G3886_o2 <= 1'b0;
    G4375_o2 <= 1'b0;
    G4901_o2 <= 1'b0;
    G5054_o2 <= 1'b0;
    G4374_o2 <= 1'b0;
    G4900_o2 <= 1'b0;
    G5053_o2 <= 1'b0;
    G5242_o2 <= 1'b0;
    G4034_o2 <= 1'b0;
    G4556_o2 <= 1'b0;
    G5064_o2 <= 1'b0;
    G5172_o2 <= 1'b0;
    G2030_o2 <= 1'b0;
    G3016_o2 <= 1'b0;
    G3520_o2 <= 1'b0;
    G3261_o2 <= 1'b0;
    G3620_o2 <= 1'b0;
    G4220_o2 <= 1'b0;
    G4719_o2 <= 1'b0;
    G5247_o2 <= 1'b0;
    G5109_o2 <= 1'b0;
    G1638_o2 <= 1'b0;
    G1976_o2 <= 1'b0;
    G3560_o2 <= 1'b0;
    G3205_o2 <= 1'b0;
    G3193_o2 <= 1'b0;
    G3367_o2 <= 1'b0;
    G3670_o2 <= 1'b0;
    n979_inv <= 1'b0;
    G1280_o2 <= 1'b0;
    G902_o2 <= 1'b0;
    G659_o2 <= 1'b0;
    G983_o2 <= 1'b0;
    G740_o2 <= 1'b0;
    G2917_o2 <= 1'b0;
    G3391_o2 <= 1'b0;
    G3494_o2 <= 1'b0;
    G1512_o2 <= 1'b0;
    G1854_o2 <= 1'b0;
    G2203_o2 <= 1'b0;
    G3493_o2 <= 1'b0;
    G3069_o2 <= 1'b0;
    G3574_o2 <= 1'b0;
    G3319_o2 <= 1'b0;
    G3667_o2 <= 1'b0;
    G3068_o2 <= 1'b0;
    G3573_o2 <= 1'b0;
    G3666_o2 <= 1'b0;
    G3318_o2 <= 1'b0;
    G3492_o2 <= 1'b0;
    G3241_o2 <= 1'b0;
    G3722_o2 <= 1'b0;
    G3422_o2 <= 1'b0;
    G1445_o2 <= 1'b0;
    G3257_o2 <= 1'b0;
    G3616_o2 <= 1'b0;
    G1634_o2 <= 1'b0;
    G1972_o2 <= 1'b0;
    G2256_o2 <= 1'b0;
    G3394_o2 <= 1'b0;
    G3557_o2 <= 1'b0;
    G3364_o2 <= 1'b0;
    G3719_o2 <= 1'b0;
    G2253_o2 <= 1'b0;
    G1583_o2 <= 1'b0;
    G1917_o2 <= 1'b0;
    G1727_o2 <= 1'b0;
    G2061_o2 <= 1'b0;
    G935_o2 <= 1'b0;
    G692_o2 <= 1'b0;
    G2136_o2 <= 1'b0;
    G1507_o2 <= 1'b0;
    G1849_o2 <= 1'b0;
    G2198_o2 <= 1'b0;
    G2197_o2 <= 1'b0;
    G1848_o2 <= 1'b0;
    G1689_o2 <= 1'b0;
    G2016_o2 <= 1'b0;
    G2314_o2 <= 1'b0;
    G2313_o2 <= 1'b0;
    G1688_o2 <= 1'b0;
    G2015_o2 <= 1'b0;
    G1847_o2 <= 1'b0;
    G2196_o2 <= 1'b0;
    G2118_o2 <= 1'b0;
    G1777_o2 <= 1'b0;
    G1630_o2 <= 1'b0;
    G1968_o2 <= 1'b0;
    G2309_o2 <= 1'b0;
    G2139_o2 <= 1'b0;
    G1580_o2 <= 1'b0;
    G2250_o2 <= 1'b0;
    G1914_o2 <= 1'b0;
    G1724_o2 <= 1'b0;
    G2058_o2 <= 1'b0;
    n2728_lo_buf_o2 <= 1'b0;
  end
endmodule


