
module mymod
(
  G1_p,
  G1_n,
  G2_p,
  G2_n,
  G3_p,
  G3_n,
  G4_p,
  G4_n,
  G5_p,
  G5_n,
  G6_p,
  G6_n,
  G7_p,
  G7_n,
  G8_p,
  G8_n,
  G9_p,
  G9_n,
  G10_p,
  G10_n,
  G11_p,
  G11_n,
  G12_p,
  G12_n,
  G13_p,
  G13_n,
  G14_p,
  G14_n,
  G15_p,
  G15_n,
  G16_p,
  G16_n,
  G17_p,
  G17_n,
  G18_p,
  G18_n,
  G19_p,
  G19_n,
  G20_p,
  G20_n,
  G21_p,
  G21_n,
  G22_p,
  G22_n,
  G23_p,
  G23_n,
  G24_p,
  G24_n,
  G25_p,
  G25_n,
  G26_p,
  G26_n,
  G27_p,
  G27_n,
  G28_p,
  G28_n,
  G29_p,
  G29_n,
  G30_p,
  G30_n,
  G31_p,
  G31_n,
  G32_p,
  G32_n,
  G33_p,
  G33_n,
  G34_p,
  G34_n,
  G35_p,
  G35_n,
  G36_p,
  G36_n,
  G37_p,
  G37_n,
  G38_p,
  G38_n,
  G39_p,
  G39_n,
  G40_p,
  G40_n,
  G41_p,
  G41_n,
  G468_p,
  G469_p,
  G470_p,
  G471_p,
  G472_p,
  G473_p,
  G474_p,
  G475_p,
  G476_p,
  G477_p,
  G478_p,
  G479_p,
  G480_p,
  G481_p,
  G482_p,
  G483_p,
  G484_p,
  G485_p,
  G486_p,
  G487_p,
  G488_p,
  G489_p,
  G490_p,
  G491_p,
  G492_p,
  G493_p,
  G494_p,
  G495_p,
  G496_p,
  G497_p,
  G498_p,
  G499_p
);

  input G1_p;input G1_n;input G2_p;input G2_n;input G3_p;input G3_n;input G4_p;input G4_n;input G5_p;input G5_n;input G6_p;input G6_n;input G7_p;input G7_n;input G8_p;input G8_n;input G9_p;input G9_n;input G10_p;input G10_n;input G11_p;input G11_n;input G12_p;input G12_n;input G13_p;input G13_n;input G14_p;input G14_n;input G15_p;input G15_n;input G16_p;input G16_n;input G17_p;input G17_n;input G18_p;input G18_n;input G19_p;input G19_n;input G20_p;input G20_n;input G21_p;input G21_n;input G22_p;input G22_n;input G23_p;input G23_n;input G24_p;input G24_n;input G25_p;input G25_n;input G26_p;input G26_n;input G27_p;input G27_n;input G28_p;input G28_n;input G29_p;input G29_n;input G30_p;input G30_n;input G31_p;input G31_n;input G32_p;input G32_n;input G33_p;input G33_n;input G34_p;input G34_n;input G35_p;input G35_n;input G36_p;input G36_n;input G37_p;input G37_n;input G38_p;input G38_n;input G39_p;input G39_n;input G40_p;input G40_n;input G41_p;input G41_n;
  output G468_p;output G469_p;output G470_p;output G471_p;output G472_p;output G473_p;output G474_p;output G475_p;output G476_p;output G477_p;output G478_p;output G479_p;output G480_p;output G481_p;output G482_p;output G483_p;output G484_p;output G485_p;output G486_p;output G487_p;output G488_p;output G489_p;output G490_p;output G491_p;output G492_p;output G493_p;output G494_p;output G495_p;output G496_p;output G497_p;output G498_p;output G499_p;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire ffc_0_p;
  wire ffc_0_n;
  wire ffc_1_p;
  wire ffc_1_n;
  wire ffc_2_p;
  wire ffc_2_n;
  wire ffc_3_p;
  wire ffc_3_n;
  wire ffc_4_p;
  wire ffc_4_n;
  wire ffc_5_p;
  wire ffc_5_n;
  wire ffc_6_p;
  wire ffc_6_n;
  wire ffc_7_p;
  wire ffc_7_n;
  wire ffc_8_p;
  wire ffc_8_n;
  wire ffc_9_p;
  wire ffc_9_n;
  wire ffc_10_p;
  wire ffc_10_n;
  wire ffc_11_p;
  wire ffc_11_n;
  wire ffc_12_p;
  wire ffc_12_n;
  wire ffc_13_p;
  wire ffc_13_n;
  wire ffc_14_p;
  wire ffc_14_n;
  wire ffc_15_p;
  wire ffc_15_n;
  wire ffc_16_p;
  wire ffc_16_n;
  wire ffc_17_p;
  wire ffc_17_n;
  wire ffc_18_p;
  wire ffc_18_n;
  wire ffc_19_p;
  wire ffc_19_n;
  wire ffc_20_p;
  wire ffc_20_n;
  wire ffc_21_p;
  wire ffc_21_n;
  wire ffc_22_p;
  wire ffc_22_n;
  wire ffc_23_p;
  wire ffc_23_n;
  wire ffc_24_p;
  wire ffc_24_n;
  wire ffc_25_p;
  wire ffc_25_n;
  wire ffc_26_p;
  wire ffc_26_n;
  wire ffc_27_p;
  wire ffc_27_n;
  wire ffc_28_p;
  wire ffc_28_n;
  wire ffc_29_p;
  wire ffc_29_n;
  wire ffc_30_p;
  wire ffc_30_n;
  wire ffc_31_p;
  wire ffc_31_n;
  wire ffc_32_p;
  wire ffc_32_n;
  wire ffc_33_p;
  wire ffc_33_n;
  wire ffc_34_p;
  wire ffc_34_n;
  wire ffc_35_p;
  wire ffc_35_n;
  wire ffc_36_p;
  wire ffc_36_n;
  wire ffc_37_p;
  wire ffc_37_n;
  wire ffc_38_p;
  wire ffc_38_n;
  wire ffc_39_p;
  wire ffc_39_n;
  wire ffc_40_p;
  wire ffc_40_n;
  wire ffc_41_p;
  wire ffc_41_n;
  wire ffc_42_p;
  wire ffc_42_n;
  wire ffc_43_p;
  wire ffc_43_n;
  wire ffc_44_p;
  wire ffc_44_n;
  wire ffc_45_p;
  wire ffc_45_n;
  wire ffc_46_p;
  wire ffc_46_n;
  wire ffc_47_p;
  wire ffc_47_n;
  wire ffc_48_p;
  wire ffc_48_n;
  wire ffc_49_p;
  wire ffc_49_n;
  wire ffc_50_p;
  wire ffc_50_n;
  wire ffc_51_p;
  wire ffc_51_n;
  wire ffc_52_p;
  wire ffc_52_n;
  wire ffc_53_p;
  wire ffc_53_n;
  wire ffc_54_p;
  wire ffc_54_n;
  wire ffc_55_p;
  wire ffc_55_n;
  wire ffc_56_p;
  wire ffc_56_n;
  wire ffc_57_p;
  wire ffc_57_n;
  wire ffc_58_p;
  wire ffc_58_n;
  wire ffc_59_p;
  wire ffc_59_n;
  wire ffc_60_p;
  wire ffc_60_n;
  wire ffc_61_p;
  wire ffc_61_n;
  wire ffc_62_p;
  wire ffc_62_n;
  wire ffc_63_p;
  wire ffc_63_n;
  wire ffc_64_p;
  wire ffc_64_n;
  wire ffc_65_p;
  wire ffc_65_n;
  wire ffc_66_p;
  wire ffc_66_n;
  wire ffc_67_p;
  wire ffc_67_n;
  wire ffc_68_p;
  wire ffc_68_n;
  wire ffc_69_p;
  wire ffc_69_n;
  wire ffc_70_p;
  wire ffc_70_n;
  wire ffc_71_p;
  wire ffc_71_n;
  wire ffc_72_p;
  wire ffc_72_n;
  wire ffc_73_p;
  wire ffc_73_n;
  wire ffc_74_p;
  wire ffc_74_n;
  wire ffc_75_p;
  wire ffc_75_n;
  wire ffc_76_p;
  wire ffc_76_n;
  wire ffc_77_p;
  wire ffc_77_n;
  wire ffc_78_p;
  wire ffc_78_n;
  wire ffc_79_p;
  wire ffc_79_n;
  wire ffc_80_p;
  wire ffc_80_n;
  wire ffc_81_p;
  wire ffc_81_n;
  wire ffc_82_p;
  wire ffc_82_n;
  wire ffc_83_p;
  wire ffc_83_n;
  wire ffc_84_p;
  wire ffc_84_n;
  wire ffc_85_p;
  wire ffc_85_n;
  wire ffc_86_p;
  wire ffc_86_n;
  wire ffc_87_p;
  wire ffc_87_n;
  wire ffc_88_p;
  wire ffc_88_n;
  wire ffc_89_p;
  wire ffc_89_n;
  wire ffc_90_p;
  wire ffc_90_n;
  wire ffc_91_p;
  wire ffc_91_n;
  wire ffc_92_p;
  wire ffc_92_n;
  wire ffc_93_p;
  wire ffc_93_n;
  wire ffc_94_p;
  wire ffc_94_n;
  wire ffc_95_p;
  wire ffc_95_n;
  wire ffc_96_p;
  wire ffc_96_n;
  wire ffc_97_p;
  wire ffc_97_n;
  wire ffc_98_p;
  wire ffc_98_n;
  wire ffc_99_p;
  wire ffc_99_n;
  wire ffc_100_p;
  wire ffc_100_n;
  wire ffc_101_p;
  wire ffc_101_n;
  wire ffc_102_p;
  wire ffc_102_n;
  wire ffc_103_p;
  wire ffc_103_n;
  wire ffc_104_p;
  wire ffc_104_n;
  wire ffc_105_p;
  wire ffc_105_n;
  wire ffc_106_p;
  wire ffc_106_n;
  wire ffc_107_p;
  wire ffc_107_n;
  wire ffc_108_p;
  wire ffc_108_n;
  wire ffc_109_p;
  wire ffc_109_n;
  wire ffc_110_p;
  wire ffc_110_n;
  wire ffc_111_p;
  wire ffc_111_n;
  wire ffc_112_p;
  wire ffc_112_n;
  wire ffc_113_p;
  wire ffc_113_n;
  wire ffc_114_p;
  wire ffc_114_n;
  wire ffc_115_p;
  wire ffc_115_n;
  wire ffc_116_p;
  wire ffc_116_n;
  wire ffc_117_p;
  wire ffc_117_n;
  wire ffc_118_p;
  wire ffc_118_n;
  wire ffc_119_p;
  wire ffc_119_n;
  wire ffc_120_p;
  wire ffc_120_n;
  wire ffc_121_p;
  wire ffc_121_n;
  wire ffc_122_p;
  wire ffc_122_n;
  wire ffc_123_p;
  wire ffc_123_n;
  wire ffc_124_p;
  wire ffc_124_n;
  wire ffc_125_p;
  wire ffc_125_n;
  wire ffc_126_p;
  wire ffc_126_n;
  wire ffc_127_p;
  wire ffc_127_n;
  wire ffc_128_p;
  wire ffc_128_n;
  wire ffc_129_p;
  wire ffc_129_n;
  wire ffc_130_p;
  wire ffc_130_n;
  wire ffc_131_p;
  wire ffc_131_n;
  wire ffc_132_p;
  wire ffc_132_n;
  wire ffc_133_p;
  wire ffc_133_n;
  wire ffc_134_p;
  wire ffc_134_n;
  wire ffc_135_p;
  wire ffc_135_n;
  wire ffc_136_p;
  wire ffc_136_n;
  wire ffc_137_p;
  wire ffc_137_n;
  wire ffc_138_p;
  wire ffc_138_n;
  wire ffc_139_p;
  wire ffc_139_n;
  wire ffc_140_p;
  wire ffc_140_n;
  wire ffc_141_p;
  wire ffc_141_n;
  wire ffc_142_p;
  wire ffc_142_n;
  wire ffc_143_p;
  wire ffc_143_n;
  wire ffc_144_p;
  wire ffc_144_n;
  wire ffc_145_p;
  wire ffc_145_n;
  wire ffc_146_p;
  wire ffc_146_n;
  wire ffc_147_p;
  wire ffc_147_n;
  wire ffc_148_p;
  wire ffc_148_n;
  wire ffc_149_p;
  wire ffc_149_n;
  wire ffc_150_p;
  wire ffc_150_n;
  wire ffc_151_p;
  wire ffc_151_n;
  wire ffc_152_p;
  wire ffc_152_n;
  wire ffc_153_p;
  wire ffc_153_n;
  wire ffc_154_p;
  wire ffc_154_n;
  wire ffc_155_p;
  wire ffc_155_n;
  wire ffc_156_p;
  wire ffc_156_n;
  wire ffc_157_p;
  wire ffc_157_n;
  wire ffc_158_p;
  wire ffc_158_n;
  wire ffc_159_p;
  wire ffc_159_n;
  wire ffc_160_p;
  wire ffc_160_n;
  wire ffc_161_p;
  wire ffc_161_n;
  wire ffc_162_p;
  wire ffc_162_n;
  wire ffc_163_p;
  wire ffc_163_n;
  wire ffc_164_p;
  wire ffc_164_n;
  wire ffc_165_p;
  wire ffc_165_n;
  wire ffc_166_p;
  wire ffc_166_n;
  wire ffc_167_p;
  wire ffc_167_n;
  wire ffc_168_p;
  wire ffc_168_n;
  wire ffc_169_p;
  wire ffc_169_n;
  wire ffc_170_p;
  wire ffc_170_n;
  wire ffc_171_p;
  wire ffc_171_n;
  wire ffc_172_p;
  wire ffc_172_n;
  wire ffc_173_p;
  wire ffc_173_n;
  wire ffc_174_p;
  wire ffc_174_n;
  wire ffc_175_p;
  wire ffc_175_n;
  wire ffc_176_p;
  wire ffc_176_n;
  wire ffc_177_p;
  wire ffc_177_n;
  wire ffc_178_p;
  wire ffc_178_n;
  wire ffc_179_p;
  wire ffc_179_n;
  wire ffc_180_p;
  wire ffc_180_n;
  wire ffc_181_p;
  wire ffc_181_n;
  wire ffc_182_p;
  wire ffc_182_n;
  wire ffc_183_p;
  wire ffc_183_n;
  wire ffc_184_p;
  wire ffc_184_n;
  wire ffc_185_p;
  wire ffc_185_n;
  wire ffc_186_p;
  wire ffc_186_n;
  wire ffc_187_p;
  wire ffc_187_n;
  wire ffc_188_p;
  wire ffc_188_n;
  wire ffc_189_p;
  wire ffc_189_n;
  wire ffc_190_p;
  wire ffc_190_n;
  wire ffc_191_p;
  wire ffc_191_n;
  wire ffc_192_p;
  wire ffc_192_n;
  wire ffc_193_p;
  wire ffc_193_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g236_n_spl_;
  wire g236_n_spl_0;
  wire g236_n_spl_1;
  wire g236_p_spl_;
  wire g236_p_spl_0;
  wire g236_p_spl_1;
  wire ffc_73_p_spl_;
  wire ffc_73_p_spl_0;
  wire ffc_73_p_spl_1;
  wire g238_p_spl_;
  wire g238_p_spl_0;
  wire g238_p_spl_1;
  wire ffc_73_n_spl_;
  wire ffc_73_n_spl_0;
  wire ffc_73_n_spl_1;
  wire g238_n_spl_;
  wire g238_n_spl_0;
  wire g238_n_spl_1;
  wire ffc_74_p_spl_;
  wire ffc_74_p_spl_0;
  wire ffc_74_p_spl_00;
  wire ffc_74_p_spl_1;
  wire ffc_74_n_spl_;
  wire ffc_74_n_spl_0;
  wire ffc_74_n_spl_00;
  wire ffc_74_n_spl_1;
  wire ffc_75_p_spl_;
  wire ffc_75_p_spl_0;
  wire ffc_75_p_spl_00;
  wire ffc_75_p_spl_01;
  wire ffc_75_p_spl_1;
  wire ffc_75_n_spl_;
  wire ffc_75_n_spl_0;
  wire ffc_75_n_spl_00;
  wire ffc_75_n_spl_01;
  wire ffc_75_n_spl_1;
  wire ffc_76_p_spl_;
  wire ffc_76_p_spl_0;
  wire ffc_76_p_spl_1;
  wire ffc_76_n_spl_;
  wire ffc_76_n_spl_0;
  wire ffc_76_n_spl_1;
  wire g256_p_spl_;
  wire g256_p_spl_0;
  wire g256_p_spl_1;
  wire g256_n_spl_;
  wire g256_n_spl_0;
  wire g256_n_spl_1;
  wire g274_p_spl_;
  wire g274_p_spl_0;
  wire g274_p_spl_1;
  wire g274_n_spl_;
  wire g274_n_spl_0;
  wire g274_n_spl_1;
  wire g292_p_spl_;
  wire g292_p_spl_0;
  wire g292_p_spl_1;
  wire g292_n_spl_;
  wire g292_n_spl_0;
  wire g292_n_spl_1;
  wire ffc_128_p_spl_;
  wire ffc_128_p_spl_0;
  wire ffc_128_p_spl_1;
  wire ffc_128_n_spl_;
  wire ffc_128_n_spl_0;
  wire ffc_128_n_spl_1;
  wire ffc_77_p_spl_;
  wire ffc_77_p_spl_0;
  wire ffc_77_p_spl_1;
  wire g310_p_spl_;
  wire g310_p_spl_0;
  wire g310_p_spl_1;
  wire ffc_77_n_spl_;
  wire ffc_77_n_spl_0;
  wire ffc_77_n_spl_1;
  wire g310_n_spl_;
  wire g310_n_spl_0;
  wire g310_n_spl_1;
  wire ffc_78_p_spl_;
  wire ffc_78_p_spl_0;
  wire ffc_78_p_spl_1;
  wire ffc_78_n_spl_;
  wire ffc_78_n_spl_0;
  wire ffc_78_n_spl_1;
  wire ffc_79_p_spl_;
  wire ffc_79_p_spl_0;
  wire ffc_79_p_spl_1;
  wire ffc_79_n_spl_;
  wire ffc_79_n_spl_0;
  wire ffc_79_n_spl_1;
  wire ffc_80_p_spl_;
  wire ffc_80_p_spl_0;
  wire ffc_80_p_spl_1;
  wire ffc_80_n_spl_;
  wire ffc_80_n_spl_0;
  wire ffc_80_n_spl_1;
  wire g328_p_spl_;
  wire g328_p_spl_0;
  wire g328_p_spl_1;
  wire g328_n_spl_;
  wire g328_n_spl_0;
  wire g328_n_spl_1;
  wire g346_p_spl_;
  wire g346_p_spl_0;
  wire g346_p_spl_1;
  wire g346_n_spl_;
  wire g346_n_spl_0;
  wire g346_n_spl_1;
  wire g364_p_spl_;
  wire g364_p_spl_0;
  wire g364_p_spl_1;
  wire g364_n_spl_;
  wire g364_n_spl_0;
  wire g364_n_spl_1;
  wire g382_n_spl_;
  wire g382_n_spl_0;
  wire g383_n_spl_;
  wire g383_n_spl_0;
  wire g385_p_spl_;
  wire g385_p_spl_0;
  wire g388_p_spl_;
  wire g388_p_spl_0;
  wire g385_n_spl_;
  wire g385_n_spl_0;
  wire g388_n_spl_;
  wire g388_n_spl_0;
  wire g386_p_spl_;
  wire g386_p_spl_0;
  wire g387_p_spl_;
  wire g387_p_spl_0;
  wire g381_n_spl_;
  wire g381_n_spl_0;
  wire g390_n_spl_;
  wire g384_n_spl_;
  wire g384_n_spl_0;
  wire g395_n_spl_;
  wire g389_n_spl_;
  wire g386_n_spl_;
  wire g386_n_spl_0;
  wire g387_n_spl_;
  wire g387_n_spl_0;
  wire g394_n_spl_;
  wire g396_n_spl_;
  wire g397_n_spl_;
  wire g391_n_spl_;
  wire g392_n_spl_;
  wire g398_n_spl_;
  wire g393_n_spl_;
  wire ffc_90_p_spl_;
  wire ffc_90_p_spl_0;
  wire ffc_94_n_spl_;
  wire ffc_90_n_spl_;
  wire ffc_94_p_spl_;
  wire ffc_94_p_spl_0;
  wire ffc_98_p_spl_;
  wire ffc_98_p_spl_0;
  wire ffc_102_n_spl_;
  wire ffc_98_n_spl_;
  wire ffc_102_p_spl_;
  wire ffc_102_p_spl_0;
  wire ffc_153_p_spl_;
  wire ffc_153_p_spl_0;
  wire ffc_153_p_spl_00;
  wire ffc_153_p_spl_01;
  wire ffc_153_p_spl_1;
  wire ffc_153_p_spl_10;
  wire ffc_153_p_spl_11;
  wire ffc_153_n_spl_;
  wire ffc_153_n_spl_0;
  wire ffc_153_n_spl_00;
  wire ffc_153_n_spl_01;
  wire ffc_153_n_spl_1;
  wire ffc_153_n_spl_10;
  wire ffc_153_n_spl_11;
  wire ffc_158_n_spl_;
  wire ffc_158_n_spl_0;
  wire ffc_158_n_spl_1;
  wire ffc_159_p_spl_;
  wire ffc_159_p_spl_0;
  wire ffc_159_p_spl_1;
  wire ffc_158_p_spl_;
  wire ffc_158_p_spl_0;
  wire ffc_158_p_spl_1;
  wire ffc_159_n_spl_;
  wire ffc_159_n_spl_0;
  wire ffc_159_n_spl_1;
  wire g421_n_spl_;
  wire g428_p_spl_;
  wire ffc_91_p_spl_;
  wire ffc_91_p_spl_0;
  wire ffc_95_n_spl_;
  wire ffc_91_n_spl_;
  wire ffc_95_p_spl_;
  wire ffc_95_p_spl_0;
  wire ffc_99_p_spl_;
  wire ffc_99_p_spl_0;
  wire ffc_103_n_spl_;
  wire ffc_99_n_spl_;
  wire ffc_103_p_spl_;
  wire ffc_103_p_spl_0;
  wire ffc_160_p_spl_;
  wire ffc_160_p_spl_0;
  wire ffc_160_p_spl_1;
  wire ffc_161_n_spl_;
  wire ffc_161_n_spl_0;
  wire ffc_161_n_spl_1;
  wire ffc_160_n_spl_;
  wire ffc_160_n_spl_0;
  wire ffc_160_n_spl_1;
  wire ffc_161_p_spl_;
  wire ffc_161_p_spl_0;
  wire ffc_161_p_spl_1;
  wire g439_n_spl_;
  wire g446_p_spl_;
  wire ffc_92_p_spl_;
  wire ffc_92_p_spl_0;
  wire ffc_96_n_spl_;
  wire ffc_92_n_spl_;
  wire ffc_96_p_spl_;
  wire ffc_96_p_spl_0;
  wire ffc_100_p_spl_;
  wire ffc_100_p_spl_0;
  wire ffc_104_n_spl_;
  wire ffc_100_n_spl_;
  wire ffc_104_p_spl_;
  wire ffc_104_p_spl_0;
  wire g457_n_spl_;
  wire g464_p_spl_;
  wire ffc_93_p_spl_;
  wire ffc_93_p_spl_0;
  wire ffc_97_n_spl_;
  wire ffc_93_n_spl_;
  wire ffc_97_p_spl_;
  wire ffc_97_p_spl_0;
  wire ffc_101_p_spl_;
  wire ffc_101_p_spl_0;
  wire ffc_105_n_spl_;
  wire ffc_101_n_spl_;
  wire ffc_105_p_spl_;
  wire ffc_105_p_spl_0;
  wire g475_n_spl_;
  wire g482_p_spl_;
  wire ffc_106_p_spl_;
  wire ffc_106_p_spl_0;
  wire ffc_110_n_spl_;
  wire ffc_106_n_spl_;
  wire ffc_110_p_spl_;
  wire ffc_110_p_spl_0;
  wire ffc_114_p_spl_;
  wire ffc_114_p_spl_0;
  wire ffc_118_n_spl_;
  wire ffc_114_n_spl_;
  wire ffc_118_p_spl_;
  wire ffc_118_p_spl_0;
  wire ffc_154_n_spl_;
  wire ffc_154_n_spl_0;
  wire ffc_154_n_spl_1;
  wire ffc_155_p_spl_;
  wire ffc_155_p_spl_0;
  wire ffc_155_p_spl_1;
  wire ffc_154_p_spl_;
  wire ffc_154_p_spl_0;
  wire ffc_154_p_spl_1;
  wire ffc_155_n_spl_;
  wire ffc_155_n_spl_0;
  wire ffc_155_n_spl_1;
  wire g493_n_spl_;
  wire g500_p_spl_;
  wire ffc_107_p_spl_;
  wire ffc_107_p_spl_0;
  wire ffc_111_n_spl_;
  wire ffc_107_n_spl_;
  wire ffc_111_p_spl_;
  wire ffc_111_p_spl_0;
  wire ffc_115_p_spl_;
  wire ffc_115_p_spl_0;
  wire ffc_119_n_spl_;
  wire ffc_115_n_spl_;
  wire ffc_119_p_spl_;
  wire ffc_119_p_spl_0;
  wire ffc_156_n_spl_;
  wire ffc_156_n_spl_0;
  wire ffc_156_n_spl_1;
  wire ffc_157_p_spl_;
  wire ffc_157_p_spl_0;
  wire ffc_157_p_spl_1;
  wire ffc_156_p_spl_;
  wire ffc_156_p_spl_0;
  wire ffc_156_p_spl_1;
  wire ffc_157_n_spl_;
  wire ffc_157_n_spl_0;
  wire ffc_157_n_spl_1;
  wire g511_n_spl_;
  wire g518_p_spl_;
  wire ffc_108_p_spl_;
  wire ffc_108_p_spl_0;
  wire ffc_112_n_spl_;
  wire ffc_108_n_spl_;
  wire ffc_112_p_spl_;
  wire ffc_112_p_spl_0;
  wire ffc_116_p_spl_;
  wire ffc_116_p_spl_0;
  wire ffc_120_n_spl_;
  wire ffc_116_n_spl_;
  wire ffc_120_p_spl_;
  wire ffc_120_p_spl_0;
  wire g529_n_spl_;
  wire g536_p_spl_;
  wire ffc_109_p_spl_;
  wire ffc_109_p_spl_0;
  wire ffc_113_n_spl_;
  wire ffc_109_n_spl_;
  wire ffc_113_p_spl_;
  wire ffc_113_p_spl_0;
  wire ffc_117_p_spl_;
  wire ffc_117_p_spl_0;
  wire ffc_121_n_spl_;
  wire ffc_117_n_spl_;
  wire ffc_121_p_spl_;
  wire ffc_121_p_spl_0;
  wire g547_n_spl_;
  wire g554_p_spl_;
  wire ffc_162_p_spl_;
  wire ffc_162_p_spl_0;
  wire ffc_163_n_spl_;
  wire ffc_162_n_spl_;
  wire ffc_163_p_spl_;
  wire ffc_163_p_spl_0;
  wire ffc_164_p_spl_;
  wire ffc_164_p_spl_0;
  wire ffc_165_n_spl_;
  wire ffc_164_n_spl_;
  wire ffc_165_p_spl_;
  wire ffc_165_p_spl_0;
  wire ffc_166_p_spl_;
  wire ffc_166_p_spl_0;
  wire ffc_167_n_spl_;
  wire ffc_166_n_spl_;
  wire ffc_167_p_spl_;
  wire ffc_167_p_spl_0;
  wire ffc_168_p_spl_;
  wire ffc_168_p_spl_0;
  wire ffc_169_n_spl_;
  wire ffc_168_n_spl_;
  wire ffc_169_p_spl_;
  wire ffc_169_p_spl_0;
  wire ffc_170_p_spl_;
  wire ffc_170_p_spl_0;
  wire ffc_171_n_spl_;
  wire ffc_170_n_spl_;
  wire ffc_171_p_spl_;
  wire ffc_171_p_spl_0;
  wire ffc_172_p_spl_;
  wire ffc_172_p_spl_0;
  wire ffc_173_n_spl_;
  wire ffc_172_n_spl_;
  wire ffc_173_p_spl_;
  wire ffc_173_p_spl_0;
  wire ffc_174_p_spl_;
  wire ffc_174_p_spl_0;
  wire ffc_175_n_spl_;
  wire ffc_174_n_spl_;
  wire ffc_175_p_spl_;
  wire ffc_175_p_spl_0;
  wire ffc_176_p_spl_;
  wire ffc_176_p_spl_0;
  wire ffc_177_n_spl_;
  wire ffc_176_n_spl_;
  wire ffc_177_p_spl_;
  wire ffc_177_p_spl_0;
  wire ffc_178_p_spl_;
  wire ffc_178_p_spl_0;
  wire ffc_179_n_spl_;
  wire ffc_178_n_spl_;
  wire ffc_179_p_spl_;
  wire ffc_179_p_spl_0;
  wire ffc_180_p_spl_;
  wire ffc_180_p_spl_0;
  wire ffc_181_n_spl_;
  wire ffc_180_n_spl_;
  wire ffc_181_p_spl_;
  wire ffc_181_p_spl_0;
  wire ffc_182_p_spl_;
  wire ffc_182_p_spl_0;
  wire ffc_183_n_spl_;
  wire ffc_182_n_spl_;
  wire ffc_183_p_spl_;
  wire ffc_183_p_spl_0;
  wire ffc_184_p_spl_;
  wire ffc_184_p_spl_0;
  wire ffc_185_n_spl_;
  wire ffc_184_n_spl_;
  wire ffc_185_p_spl_;
  wire ffc_185_p_spl_0;
  wire ffc_186_p_spl_;
  wire ffc_186_p_spl_0;
  wire ffc_187_n_spl_;
  wire ffc_186_n_spl_;
  wire ffc_187_p_spl_;
  wire ffc_187_p_spl_0;
  wire ffc_188_p_spl_;
  wire ffc_188_p_spl_0;
  wire ffc_189_n_spl_;
  wire ffc_188_n_spl_;
  wire ffc_189_p_spl_;
  wire ffc_189_p_spl_0;
  wire ffc_190_p_spl_;
  wire ffc_190_p_spl_0;
  wire ffc_191_n_spl_;
  wire ffc_190_n_spl_;
  wire ffc_191_p_spl_;
  wire ffc_191_p_spl_0;
  wire ffc_192_p_spl_;
  wire ffc_192_p_spl_0;
  wire ffc_193_n_spl_;
  wire ffc_192_n_spl_;
  wire ffc_193_p_spl_;
  wire ffc_193_p_spl_0;

  andX
  g_g236_p
  (
    .dout(g236_p),
    .din1(ffc_122_n),
    .din2(ffc_123_n)
  );


  orX
  g_g236_n
  (
    .dout(g236_n),
    .din1(ffc_122_p),
    .din2(ffc_123_p)
  );


  andX
  g_g237_p
  (
    .dout(g237_p),
    .din1(ffc_124_p),
    .din2(ffc_126_p)
  );


  orX
  g_g237_n
  (
    .dout(g237_n),
    .din1(ffc_124_n),
    .din2(ffc_126_n)
  );


  andX
  g_g238_p
  (
    .dout(g238_p),
    .din1(g236_n_spl_0),
    .din2(g237_p)
  );


  orX
  g_g238_n
  (
    .dout(g238_n),
    .din1(g236_p_spl_0),
    .din2(g237_n)
  );


  andX
  g_g239_p
  (
    .dout(g239_p),
    .din1(ffc_73_p_spl_0),
    .din2(g238_p_spl_0)
  );


  orX
  g_g239_n
  (
    .dout(g239_n),
    .din1(ffc_73_n_spl_0),
    .din2(g238_n_spl_0)
  );


  andX
  g_g240_p
  (
    .dout(g240_p),
    .din1(ffc_0_n),
    .din2(g239_p)
  );


  andX
  g_g241_p
  (
    .dout(g241_p),
    .din1(ffc_0_p),
    .din2(g239_n)
  );


  orX
  g_g242_n
  (
    .dout(g242_n),
    .din1(g240_p),
    .din2(g241_p)
  );


  andX
  g_g243_p
  (
    .dout(g243_p),
    .din1(ffc_74_p_spl_00),
    .din2(g238_p_spl_0)
  );


  orX
  g_g243_n
  (
    .dout(g243_n),
    .din1(ffc_74_n_spl_00),
    .din2(g238_n_spl_0)
  );


  andX
  g_g244_p
  (
    .dout(g244_p),
    .din1(ffc_1_n),
    .din2(g243_p)
  );


  andX
  g_g245_p
  (
    .dout(g245_p),
    .din1(ffc_1_p),
    .din2(g243_n)
  );


  orX
  g_g246_n
  (
    .dout(g246_n),
    .din1(g244_p),
    .din2(g245_p)
  );


  andX
  g_g247_p
  (
    .dout(g247_p),
    .din1(ffc_75_p_spl_00),
    .din2(g238_p_spl_1)
  );


  orX
  g_g247_n
  (
    .dout(g247_n),
    .din1(ffc_75_n_spl_00),
    .din2(g238_n_spl_1)
  );


  andX
  g_g248_p
  (
    .dout(g248_p),
    .din1(ffc_2_n),
    .din2(g247_p)
  );


  andX
  g_g249_p
  (
    .dout(g249_p),
    .din1(ffc_2_p),
    .din2(g247_n)
  );


  orX
  g_g250_n
  (
    .dout(g250_n),
    .din1(g248_p),
    .din2(g249_p)
  );


  andX
  g_g251_p
  (
    .dout(g251_p),
    .din1(ffc_76_p_spl_0),
    .din2(g238_p_spl_1)
  );


  orX
  g_g251_n
  (
    .dout(g251_n),
    .din1(ffc_76_n_spl_0),
    .din2(g238_n_spl_1)
  );


  andX
  g_g252_p
  (
    .dout(g252_p),
    .din1(ffc_3_n),
    .din2(g251_p)
  );


  andX
  g_g253_p
  (
    .dout(g253_p),
    .din1(ffc_3_p),
    .din2(g251_n)
  );


  orX
  g_g254_n
  (
    .dout(g254_n),
    .din1(g252_p),
    .din2(g253_p)
  );


  andX
  g_g255_p
  (
    .dout(g255_p),
    .din1(ffc_83_p),
    .din2(ffc_89_n)
  );


  orX
  g_g255_n
  (
    .dout(g255_n),
    .din1(ffc_83_n),
    .din2(ffc_89_p)
  );


  andX
  g_g256_p
  (
    .dout(g256_p),
    .din1(g236_n_spl_0),
    .din2(g255_p)
  );


  orX
  g_g256_n
  (
    .dout(g256_n),
    .din1(g236_p_spl_0),
    .din2(g255_n)
  );


  andX
  g_g257_p
  (
    .dout(g257_p),
    .din1(ffc_73_p_spl_0),
    .din2(g256_p_spl_0)
  );


  orX
  g_g257_n
  (
    .dout(g257_n),
    .din1(ffc_73_n_spl_0),
    .din2(g256_n_spl_0)
  );


  andX
  g_g258_p
  (
    .dout(g258_p),
    .din1(ffc_4_n),
    .din2(g257_p)
  );


  andX
  g_g259_p
  (
    .dout(g259_p),
    .din1(ffc_4_p),
    .din2(g257_n)
  );


  orX
  g_g260_n
  (
    .dout(g260_n),
    .din1(g258_p),
    .din2(g259_p)
  );


  andX
  g_g261_p
  (
    .dout(g261_p),
    .din1(ffc_74_p_spl_00),
    .din2(g256_p_spl_0)
  );


  orX
  g_g261_n
  (
    .dout(g261_n),
    .din1(ffc_74_n_spl_00),
    .din2(g256_n_spl_0)
  );


  andX
  g_g262_p
  (
    .dout(g262_p),
    .din1(ffc_5_n),
    .din2(g261_p)
  );


  andX
  g_g263_p
  (
    .dout(g263_p),
    .din1(ffc_5_p),
    .din2(g261_n)
  );


  orX
  g_g264_n
  (
    .dout(g264_n),
    .din1(g262_p),
    .din2(g263_p)
  );


  andX
  g_g265_p
  (
    .dout(g265_p),
    .din1(ffc_75_p_spl_00),
    .din2(g256_p_spl_1)
  );


  orX
  g_g265_n
  (
    .dout(g265_n),
    .din1(ffc_75_n_spl_00),
    .din2(g256_n_spl_1)
  );


  andX
  g_g266_p
  (
    .dout(g266_p),
    .din1(ffc_6_n),
    .din2(g265_p)
  );


  andX
  g_g267_p
  (
    .dout(g267_p),
    .din1(ffc_6_p),
    .din2(g265_n)
  );


  orX
  g_g268_n
  (
    .dout(g268_n),
    .din1(g266_p),
    .din2(g267_p)
  );


  andX
  g_g269_p
  (
    .dout(g269_p),
    .din1(ffc_76_p_spl_0),
    .din2(g256_p_spl_1)
  );


  orX
  g_g269_n
  (
    .dout(g269_n),
    .din1(ffc_76_n_spl_0),
    .din2(g256_n_spl_1)
  );


  andX
  g_g270_p
  (
    .dout(g270_p),
    .din1(ffc_7_n),
    .din2(g269_p)
  );


  andX
  g_g271_p
  (
    .dout(g271_p),
    .din1(ffc_7_p),
    .din2(g269_n)
  );


  orX
  g_g272_n
  (
    .dout(g272_n),
    .din1(g270_p),
    .din2(g271_p)
  );


  andX
  g_g273_p
  (
    .dout(g273_p),
    .din1(ffc_84_n),
    .din2(ffc_85_p)
  );


  orX
  g_g273_n
  (
    .dout(g273_n),
    .din1(ffc_84_p),
    .din2(ffc_85_n)
  );


  andX
  g_g274_p
  (
    .dout(g274_p),
    .din1(g236_n_spl_1),
    .din2(g273_p)
  );


  orX
  g_g274_n
  (
    .dout(g274_n),
    .din1(g236_p_spl_1),
    .din2(g273_n)
  );


  andX
  g_g275_p
  (
    .dout(g275_p),
    .din1(ffc_73_p_spl_1),
    .din2(g274_p_spl_0)
  );


  orX
  g_g275_n
  (
    .dout(g275_n),
    .din1(ffc_73_n_spl_1),
    .din2(g274_n_spl_0)
  );


  andX
  g_g276_p
  (
    .dout(g276_p),
    .din1(ffc_8_n),
    .din2(g275_p)
  );


  andX
  g_g277_p
  (
    .dout(g277_p),
    .din1(ffc_8_p),
    .din2(g275_n)
  );


  orX
  g_g278_n
  (
    .dout(g278_n),
    .din1(g276_p),
    .din2(g277_p)
  );


  andX
  g_g279_p
  (
    .dout(g279_p),
    .din1(ffc_74_p_spl_0),
    .din2(g274_p_spl_0)
  );


  orX
  g_g279_n
  (
    .dout(g279_n),
    .din1(ffc_74_n_spl_0),
    .din2(g274_n_spl_0)
  );


  andX
  g_g280_p
  (
    .dout(g280_p),
    .din1(ffc_9_n),
    .din2(g279_p)
  );


  andX
  g_g281_p
  (
    .dout(g281_p),
    .din1(ffc_9_p),
    .din2(g279_n)
  );


  orX
  g_g282_n
  (
    .dout(g282_n),
    .din1(g280_p),
    .din2(g281_p)
  );


  andX
  g_g283_p
  (
    .dout(g283_p),
    .din1(ffc_75_p_spl_01),
    .din2(g274_p_spl_1)
  );


  orX
  g_g283_n
  (
    .dout(g283_n),
    .din1(ffc_75_n_spl_01),
    .din2(g274_n_spl_1)
  );


  andX
  g_g284_p
  (
    .dout(g284_p),
    .din1(ffc_10_n),
    .din2(g283_p)
  );


  andX
  g_g285_p
  (
    .dout(g285_p),
    .din1(ffc_10_p),
    .din2(g283_n)
  );


  orX
  g_g286_n
  (
    .dout(g286_n),
    .din1(g284_p),
    .din2(g285_p)
  );


  andX
  g_g287_p
  (
    .dout(g287_p),
    .din1(ffc_76_p_spl_1),
    .din2(g274_p_spl_1)
  );


  orX
  g_g287_n
  (
    .dout(g287_n),
    .din1(ffc_76_n_spl_1),
    .din2(g274_n_spl_1)
  );


  andX
  g_g288_p
  (
    .dout(g288_p),
    .din1(ffc_11_n),
    .din2(g287_p)
  );


  andX
  g_g289_p
  (
    .dout(g289_p),
    .din1(ffc_11_p),
    .din2(g287_n)
  );


  orX
  g_g290_n
  (
    .dout(g290_n),
    .din1(g288_p),
    .din2(g289_p)
  );


  andX
  g_g291_p
  (
    .dout(g291_p),
    .din1(ffc_125_p),
    .din2(ffc_127_p)
  );


  orX
  g_g291_n
  (
    .dout(g291_n),
    .din1(ffc_125_n),
    .din2(ffc_127_n)
  );


  andX
  g_g292_p
  (
    .dout(g292_p),
    .din1(g236_n_spl_1),
    .din2(g291_p)
  );


  orX
  g_g292_n
  (
    .dout(g292_n),
    .din1(g236_p_spl_1),
    .din2(g291_n)
  );


  andX
  g_g293_p
  (
    .dout(g293_p),
    .din1(ffc_73_p_spl_1),
    .din2(g292_p_spl_0)
  );


  orX
  g_g293_n
  (
    .dout(g293_n),
    .din1(ffc_73_n_spl_1),
    .din2(g292_n_spl_0)
  );


  andX
  g_g294_p
  (
    .dout(g294_p),
    .din1(ffc_12_n),
    .din2(g293_p)
  );


  andX
  g_g295_p
  (
    .dout(g295_p),
    .din1(ffc_12_p),
    .din2(g293_n)
  );


  orX
  g_g296_n
  (
    .dout(g296_n),
    .din1(g294_p),
    .din2(g295_p)
  );


  andX
  g_g297_p
  (
    .dout(g297_p),
    .din1(ffc_74_p_spl_1),
    .din2(g292_p_spl_0)
  );


  orX
  g_g297_n
  (
    .dout(g297_n),
    .din1(ffc_74_n_spl_1),
    .din2(g292_n_spl_0)
  );


  andX
  g_g298_p
  (
    .dout(g298_p),
    .din1(ffc_13_n),
    .din2(g297_p)
  );


  andX
  g_g299_p
  (
    .dout(g299_p),
    .din1(ffc_13_p),
    .din2(g297_n)
  );


  orX
  g_g300_n
  (
    .dout(g300_n),
    .din1(g298_p),
    .din2(g299_p)
  );


  andX
  g_g301_p
  (
    .dout(g301_p),
    .din1(ffc_75_p_spl_01),
    .din2(g292_p_spl_1)
  );


  orX
  g_g301_n
  (
    .dout(g301_n),
    .din1(ffc_75_n_spl_01),
    .din2(g292_n_spl_1)
  );


  andX
  g_g302_p
  (
    .dout(g302_p),
    .din1(ffc_14_n),
    .din2(g301_p)
  );


  andX
  g_g303_p
  (
    .dout(g303_p),
    .din1(ffc_14_p),
    .din2(g301_n)
  );


  orX
  g_g304_n
  (
    .dout(g304_n),
    .din1(g302_p),
    .din2(g303_p)
  );


  andX
  g_g305_p
  (
    .dout(g305_p),
    .din1(ffc_76_p_spl_1),
    .din2(g292_p_spl_1)
  );


  orX
  g_g305_n
  (
    .dout(g305_n),
    .din1(ffc_76_n_spl_1),
    .din2(g292_n_spl_1)
  );


  andX
  g_g306_p
  (
    .dout(g306_p),
    .din1(ffc_15_n),
    .din2(g305_p)
  );


  andX
  g_g307_p
  (
    .dout(g307_p),
    .din1(ffc_15_p),
    .din2(g305_n)
  );


  orX
  g_g308_n
  (
    .dout(g308_n),
    .din1(g306_p),
    .din2(g307_p)
  );


  andX
  g_g309_p
  (
    .dout(g309_p),
    .din1(ffc_88_p),
    .din2(ffc_128_p_spl_0)
  );


  orX
  g_g309_n
  (
    .dout(g309_n),
    .din1(ffc_88_n),
    .din2(ffc_128_n_spl_0)
  );


  andX
  g_g310_p
  (
    .dout(g310_p),
    .din1(ffc_75_p_spl_1),
    .din2(g309_p)
  );


  orX
  g_g310_n
  (
    .dout(g310_n),
    .din1(ffc_75_n_spl_1),
    .din2(g309_n)
  );


  andX
  g_g311_p
  (
    .dout(g311_p),
    .din1(ffc_77_p_spl_0),
    .din2(g310_p_spl_0)
  );


  orX
  g_g311_n
  (
    .dout(g311_n),
    .din1(ffc_77_n_spl_0),
    .din2(g310_n_spl_0)
  );


  andX
  g_g312_p
  (
    .dout(g312_p),
    .din1(ffc_16_n),
    .din2(g311_p)
  );


  andX
  g_g313_p
  (
    .dout(g313_p),
    .din1(ffc_16_p),
    .din2(g311_n)
  );


  orX
  g_g314_n
  (
    .dout(g314_n),
    .din1(g312_p),
    .din2(g313_p)
  );


  andX
  g_g315_p
  (
    .dout(g315_p),
    .din1(ffc_78_p_spl_0),
    .din2(g310_p_spl_0)
  );


  orX
  g_g315_n
  (
    .dout(g315_n),
    .din1(ffc_78_n_spl_0),
    .din2(g310_n_spl_0)
  );


  andX
  g_g316_p
  (
    .dout(g316_p),
    .din1(ffc_17_n),
    .din2(g315_p)
  );


  andX
  g_g317_p
  (
    .dout(g317_p),
    .din1(ffc_17_p),
    .din2(g315_n)
  );


  orX
  g_g318_n
  (
    .dout(g318_n),
    .din1(g316_p),
    .din2(g317_p)
  );


  andX
  g_g319_p
  (
    .dout(g319_p),
    .din1(ffc_79_p_spl_0),
    .din2(g310_p_spl_1)
  );


  orX
  g_g319_n
  (
    .dout(g319_n),
    .din1(ffc_79_n_spl_0),
    .din2(g310_n_spl_1)
  );


  andX
  g_g320_p
  (
    .dout(g320_p),
    .din1(ffc_18_n),
    .din2(g319_p)
  );


  andX
  g_g321_p
  (
    .dout(g321_p),
    .din1(ffc_18_p),
    .din2(g319_n)
  );


  orX
  g_g322_n
  (
    .dout(g322_n),
    .din1(g320_p),
    .din2(g321_p)
  );


  andX
  g_g323_p
  (
    .dout(g323_p),
    .din1(ffc_80_p_spl_0),
    .din2(g310_p_spl_1)
  );


  orX
  g_g323_n
  (
    .dout(g323_n),
    .din1(ffc_80_n_spl_0),
    .din2(g310_n_spl_1)
  );


  andX
  g_g324_p
  (
    .dout(g324_p),
    .din1(ffc_19_n),
    .din2(g323_p)
  );


  andX
  g_g325_p
  (
    .dout(g325_p),
    .din1(ffc_19_p),
    .din2(g323_n)
  );


  orX
  g_g326_n
  (
    .dout(g326_n),
    .din1(g324_p),
    .din2(g325_p)
  );


  andX
  g_g327_p
  (
    .dout(g327_p),
    .din1(ffc_81_p),
    .din2(ffc_82_p)
  );


  orX
  g_g327_n
  (
    .dout(g327_n),
    .din1(ffc_81_n),
    .din2(ffc_82_n)
  );


  andX
  g_g328_p
  (
    .dout(g328_p),
    .din1(ffc_128_p_spl_0),
    .din2(g327_p)
  );


  orX
  g_g328_n
  (
    .dout(g328_n),
    .din1(ffc_128_n_spl_0),
    .din2(g327_n)
  );


  andX
  g_g329_p
  (
    .dout(g329_p),
    .din1(ffc_77_p_spl_0),
    .din2(g328_p_spl_0)
  );


  orX
  g_g329_n
  (
    .dout(g329_n),
    .din1(ffc_77_n_spl_0),
    .din2(g328_n_spl_0)
  );


  andX
  g_g330_p
  (
    .dout(g330_p),
    .din1(ffc_20_n),
    .din2(g329_p)
  );


  andX
  g_g331_p
  (
    .dout(g331_p),
    .din1(ffc_20_p),
    .din2(g329_n)
  );


  orX
  g_g332_n
  (
    .dout(g332_n),
    .din1(g330_p),
    .din2(g331_p)
  );


  andX
  g_g333_p
  (
    .dout(g333_p),
    .din1(ffc_78_p_spl_0),
    .din2(g328_p_spl_0)
  );


  orX
  g_g333_n
  (
    .dout(g333_n),
    .din1(ffc_78_n_spl_0),
    .din2(g328_n_spl_0)
  );


  andX
  g_g334_p
  (
    .dout(g334_p),
    .din1(ffc_21_n),
    .din2(g333_p)
  );


  andX
  g_g335_p
  (
    .dout(g335_p),
    .din1(ffc_21_p),
    .din2(g333_n)
  );


  orX
  g_g336_n
  (
    .dout(g336_n),
    .din1(g334_p),
    .din2(g335_p)
  );


  andX
  g_g337_p
  (
    .dout(g337_p),
    .din1(ffc_79_p_spl_0),
    .din2(g328_p_spl_1)
  );


  orX
  g_g337_n
  (
    .dout(g337_n),
    .din1(ffc_79_n_spl_0),
    .din2(g328_n_spl_1)
  );


  andX
  g_g338_p
  (
    .dout(g338_p),
    .din1(ffc_22_n),
    .din2(g337_p)
  );


  andX
  g_g339_p
  (
    .dout(g339_p),
    .din1(ffc_22_p),
    .din2(g337_n)
  );


  orX
  g_g340_n
  (
    .dout(g340_n),
    .din1(g338_p),
    .din2(g339_p)
  );


  andX
  g_g341_p
  (
    .dout(g341_p),
    .din1(ffc_80_p_spl_0),
    .din2(g328_p_spl_1)
  );


  orX
  g_g341_n
  (
    .dout(g341_n),
    .din1(ffc_80_n_spl_0),
    .din2(g328_n_spl_1)
  );


  andX
  g_g342_p
  (
    .dout(g342_p),
    .din1(ffc_23_n),
    .din2(g341_p)
  );


  andX
  g_g343_p
  (
    .dout(g343_p),
    .din1(ffc_23_p),
    .din2(g341_n)
  );


  orX
  g_g344_n
  (
    .dout(g344_n),
    .din1(g342_p),
    .din2(g343_p)
  );


  andX
  g_g345_p
  (
    .dout(g345_p),
    .din1(ffc_75_p_spl_1),
    .din2(ffc_87_p)
  );


  orX
  g_g345_n
  (
    .dout(g345_n),
    .din1(ffc_75_n_spl_1),
    .din2(ffc_87_n)
  );


  andX
  g_g346_p
  (
    .dout(g346_p),
    .din1(ffc_128_p_spl_1),
    .din2(g345_p)
  );


  orX
  g_g346_n
  (
    .dout(g346_n),
    .din1(ffc_128_n_spl_1),
    .din2(g345_n)
  );


  andX
  g_g347_p
  (
    .dout(g347_p),
    .din1(ffc_77_p_spl_1),
    .din2(g346_p_spl_0)
  );


  orX
  g_g347_n
  (
    .dout(g347_n),
    .din1(ffc_77_n_spl_1),
    .din2(g346_n_spl_0)
  );


  andX
  g_g348_p
  (
    .dout(g348_p),
    .din1(ffc_24_n),
    .din2(g347_p)
  );


  andX
  g_g349_p
  (
    .dout(g349_p),
    .din1(ffc_24_p),
    .din2(g347_n)
  );


  orX
  g_g350_n
  (
    .dout(g350_n),
    .din1(g348_p),
    .din2(g349_p)
  );


  andX
  g_g351_p
  (
    .dout(g351_p),
    .din1(ffc_78_p_spl_1),
    .din2(g346_p_spl_0)
  );


  orX
  g_g351_n
  (
    .dout(g351_n),
    .din1(ffc_78_n_spl_1),
    .din2(g346_n_spl_0)
  );


  andX
  g_g352_p
  (
    .dout(g352_p),
    .din1(ffc_25_n),
    .din2(g351_p)
  );


  andX
  g_g353_p
  (
    .dout(g353_p),
    .din1(ffc_25_p),
    .din2(g351_n)
  );


  orX
  g_g354_n
  (
    .dout(g354_n),
    .din1(g352_p),
    .din2(g353_p)
  );


  andX
  g_g355_p
  (
    .dout(g355_p),
    .din1(ffc_79_p_spl_1),
    .din2(g346_p_spl_1)
  );


  orX
  g_g355_n
  (
    .dout(g355_n),
    .din1(ffc_79_n_spl_1),
    .din2(g346_n_spl_1)
  );


  andX
  g_g356_p
  (
    .dout(g356_p),
    .din1(ffc_26_n),
    .din2(g355_p)
  );


  andX
  g_g357_p
  (
    .dout(g357_p),
    .din1(ffc_26_p),
    .din2(g355_n)
  );


  orX
  g_g358_n
  (
    .dout(g358_n),
    .din1(g356_p),
    .din2(g357_p)
  );


  andX
  g_g359_p
  (
    .dout(g359_p),
    .din1(ffc_80_p_spl_1),
    .din2(g346_p_spl_1)
  );


  orX
  g_g359_n
  (
    .dout(g359_n),
    .din1(ffc_80_n_spl_1),
    .din2(g346_n_spl_1)
  );


  andX
  g_g360_p
  (
    .dout(g360_p),
    .din1(ffc_27_n),
    .din2(g359_p)
  );


  andX
  g_g361_p
  (
    .dout(g361_p),
    .din1(ffc_27_p),
    .din2(g359_n)
  );


  orX
  g_g362_n
  (
    .dout(g362_n),
    .din1(g360_p),
    .din2(g361_p)
  );


  andX
  g_g363_p
  (
    .dout(g363_p),
    .din1(ffc_74_p_spl_1),
    .din2(ffc_86_p)
  );


  orX
  g_g363_n
  (
    .dout(g363_n),
    .din1(ffc_74_n_spl_1),
    .din2(ffc_86_n)
  );


  andX
  g_g364_p
  (
    .dout(g364_p),
    .din1(ffc_128_p_spl_1),
    .din2(g363_p)
  );


  orX
  g_g364_n
  (
    .dout(g364_n),
    .din1(ffc_128_n_spl_1),
    .din2(g363_n)
  );


  andX
  g_g365_p
  (
    .dout(g365_p),
    .din1(ffc_77_p_spl_1),
    .din2(g364_p_spl_0)
  );


  orX
  g_g365_n
  (
    .dout(g365_n),
    .din1(ffc_77_n_spl_1),
    .din2(g364_n_spl_0)
  );


  andX
  g_g366_p
  (
    .dout(g366_p),
    .din1(ffc_28_n),
    .din2(g365_p)
  );


  andX
  g_g367_p
  (
    .dout(g367_p),
    .din1(ffc_28_p),
    .din2(g365_n)
  );


  orX
  g_g368_n
  (
    .dout(g368_n),
    .din1(g366_p),
    .din2(g367_p)
  );


  andX
  g_g369_p
  (
    .dout(g369_p),
    .din1(ffc_78_p_spl_1),
    .din2(g364_p_spl_0)
  );


  orX
  g_g369_n
  (
    .dout(g369_n),
    .din1(ffc_78_n_spl_1),
    .din2(g364_n_spl_0)
  );


  andX
  g_g370_p
  (
    .dout(g370_p),
    .din1(ffc_29_n),
    .din2(g369_p)
  );


  andX
  g_g371_p
  (
    .dout(g371_p),
    .din1(ffc_29_p),
    .din2(g369_n)
  );


  orX
  g_g372_n
  (
    .dout(g372_n),
    .din1(g370_p),
    .din2(g371_p)
  );


  andX
  g_g373_p
  (
    .dout(g373_p),
    .din1(ffc_79_p_spl_1),
    .din2(g364_p_spl_1)
  );


  orX
  g_g373_n
  (
    .dout(g373_n),
    .din1(ffc_79_n_spl_1),
    .din2(g364_n_spl_1)
  );


  andX
  g_g374_p
  (
    .dout(g374_p),
    .din1(ffc_30_n),
    .din2(g373_p)
  );


  andX
  g_g375_p
  (
    .dout(g375_p),
    .din1(ffc_30_p),
    .din2(g373_n)
  );


  orX
  g_g376_n
  (
    .dout(g376_n),
    .din1(g374_p),
    .din2(g375_p)
  );


  andX
  g_g377_p
  (
    .dout(g377_p),
    .din1(ffc_80_p_spl_1),
    .din2(g364_p_spl_1)
  );


  orX
  g_g377_n
  (
    .dout(g377_n),
    .din1(ffc_80_n_spl_1),
    .din2(g364_n_spl_1)
  );


  andX
  g_g378_p
  (
    .dout(g378_p),
    .din1(ffc_31_n),
    .din2(g377_p)
  );


  andX
  g_g379_p
  (
    .dout(g379_p),
    .din1(ffc_31_p),
    .din2(g377_n)
  );


  orX
  g_g380_n
  (
    .dout(g380_n),
    .din1(g378_p),
    .din2(g379_p)
  );


  andX
  g_g381_p
  (
    .dout(g381_p),
    .din1(ffc_129_n),
    .din2(ffc_130_n)
  );


  orX
  g_g381_n
  (
    .dout(g381_n),
    .din1(ffc_129_p),
    .din2(ffc_130_p)
  );


  andX
  g_g382_p
  (
    .dout(g382_p),
    .din1(ffc_131_n),
    .din2(ffc_132_n)
  );


  orX
  g_g382_n
  (
    .dout(g382_n),
    .din1(ffc_131_p),
    .din2(ffc_132_p)
  );


  andX
  g_g383_p
  (
    .dout(g383_p),
    .din1(ffc_133_n),
    .din2(ffc_134_n)
  );


  orX
  g_g383_n
  (
    .dout(g383_n),
    .din1(ffc_133_p),
    .din2(ffc_134_p)
  );


  andX
  g_g384_p
  (
    .dout(g384_p),
    .din1(ffc_135_n),
    .din2(ffc_136_n)
  );


  orX
  g_g384_n
  (
    .dout(g384_n),
    .din1(ffc_135_p),
    .din2(ffc_136_p)
  );


  andX
  g_g385_p
  (
    .dout(g385_p),
    .din1(ffc_137_n),
    .din2(ffc_138_n)
  );


  orX
  g_g385_n
  (
    .dout(g385_n),
    .din1(ffc_137_p),
    .din2(ffc_138_p)
  );


  andX
  g_g386_p
  (
    .dout(g386_p),
    .din1(ffc_139_n),
    .din2(ffc_140_n)
  );


  orX
  g_g386_n
  (
    .dout(g386_n),
    .din1(ffc_139_p),
    .din2(ffc_140_p)
  );


  andX
  g_g387_p
  (
    .dout(g387_p),
    .din1(ffc_141_n),
    .din2(ffc_142_n)
  );


  orX
  g_g387_n
  (
    .dout(g387_n),
    .din1(ffc_141_p),
    .din2(ffc_142_p)
  );


  andX
  g_g388_p
  (
    .dout(g388_p),
    .din1(ffc_143_n),
    .din2(ffc_144_n)
  );


  orX
  g_g388_n
  (
    .dout(g388_n),
    .din1(ffc_143_p),
    .din2(ffc_144_p)
  );


  orX
  g_g389_n
  (
    .dout(g389_n),
    .din1(g381_p),
    .din2(g382_n_spl_0)
  );


  orX
  g_g390_n
  (
    .dout(g390_n),
    .din1(g383_n_spl_0),
    .din2(g384_p)
  );


  orX
  g_g391_n
  (
    .dout(g391_n),
    .din1(g385_p_spl_0),
    .din2(g388_p_spl_0)
  );


  andX
  g_g392_p
  (
    .dout(g392_p),
    .din1(g385_p_spl_0),
    .din2(g388_p_spl_0)
  );


  orX
  g_g392_n
  (
    .dout(g392_n),
    .din1(g385_n_spl_0),
    .din2(g388_n_spl_0)
  );


  orX
  g_g393_n
  (
    .dout(g393_n),
    .din1(g386_p_spl_0),
    .din2(g387_p_spl_0)
  );


  orX
  g_g394_n
  (
    .dout(g394_n),
    .din1(g381_n_spl_0),
    .din2(g390_n_spl_)
  );


  orX
  g_g395_n
  (
    .dout(g395_n),
    .din1(g381_n_spl_0),
    .din2(g384_n_spl_0)
  );


  orX
  g_g396_n
  (
    .dout(g396_n),
    .din1(g382_p),
    .din2(g395_n_spl_)
  );


  orX
  g_g397_n
  (
    .dout(g397_n),
    .din1(g384_n_spl_0),
    .din2(g389_n_spl_)
  );


  andX
  g_g398_p
  (
    .dout(g398_p),
    .din1(g386_p_spl_0),
    .din2(g387_p_spl_0)
  );


  orX
  g_g398_n
  (
    .dout(g398_n),
    .din1(g386_n_spl_0),
    .din2(g387_n_spl_0)
  );


  orX
  g_g399_n
  (
    .dout(g399_n),
    .din1(g383_p),
    .din2(g395_n_spl_)
  );


  andX
  g_g400_p
  (
    .dout(g400_p),
    .din1(g394_n_spl_),
    .din2(g399_n)
  );


  orX
  g_g401_n
  (
    .dout(g401_n),
    .din1(g382_n_spl_0),
    .din2(g400_p)
  );


  andX
  g_g402_p
  (
    .dout(g402_p),
    .din1(g396_n_spl_),
    .din2(g397_n_spl_)
  );


  orX
  g_g403_n
  (
    .dout(g403_n),
    .din1(g383_n_spl_0),
    .din2(g402_p)
  );


  andX
  g_g404_p
  (
    .dout(g404_p),
    .din1(g385_n_spl_0),
    .din2(g386_p_spl_)
  );


  andX
  g_g405_p
  (
    .dout(g405_p),
    .din1(g385_p_spl_),
    .din2(g386_n_spl_0)
  );


  andX
  g_g406_p
  (
    .dout(g406_p),
    .din1(g387_n_spl_0),
    .din2(g388_p_spl_)
  );


  andX
  g_g407_p
  (
    .dout(g407_p),
    .din1(g387_p_spl_),
    .din2(g388_n_spl_0)
  );


  andX
  g_g408_p
  (
    .dout(g408_p),
    .din1(g391_n_spl_),
    .din2(g392_n_spl_)
  );


  orX
  g_g409_n
  (
    .dout(g409_n),
    .din1(g398_n_spl_),
    .din2(g408_p)
  );


  andX
  g_g410_p
  (
    .dout(g410_p),
    .din1(g392_p),
    .din2(g393_n_spl_)
  );


  orX
  g_g411_n
  (
    .dout(g411_n),
    .din1(g398_p),
    .din2(g410_p)
  );


  andX
  g_g412_p
  (
    .dout(g412_p),
    .din1(g409_n),
    .din2(g411_n)
  );


  andX
  g_g413_p
  (
    .dout(g413_p),
    .din1(ffc_90_p_spl_0),
    .din2(ffc_94_n_spl_)
  );


  orX
  g_g413_n
  (
    .dout(g413_n),
    .din1(ffc_90_n_spl_),
    .din2(ffc_94_p_spl_0)
  );


  andX
  g_g414_p
  (
    .dout(g414_p),
    .din1(ffc_90_n_spl_),
    .din2(ffc_94_p_spl_0)
  );


  orX
  g_g414_n
  (
    .dout(g414_n),
    .din1(ffc_90_p_spl_0),
    .din2(ffc_94_n_spl_)
  );


  andX
  g_g415_p
  (
    .dout(g415_p),
    .din1(g413_n),
    .din2(g414_n)
  );


  orX
  g_g415_n
  (
    .dout(g415_n),
    .din1(g413_p),
    .din2(g414_p)
  );


  andX
  g_g416_p
  (
    .dout(g416_p),
    .din1(ffc_98_p_spl_0),
    .din2(ffc_102_n_spl_)
  );


  orX
  g_g416_n
  (
    .dout(g416_n),
    .din1(ffc_98_n_spl_),
    .din2(ffc_102_p_spl_0)
  );


  andX
  g_g417_p
  (
    .dout(g417_p),
    .din1(ffc_98_n_spl_),
    .din2(ffc_102_p_spl_0)
  );


  orX
  g_g417_n
  (
    .dout(g417_n),
    .din1(ffc_98_p_spl_0),
    .din2(ffc_102_n_spl_)
  );


  andX
  g_g418_p
  (
    .dout(g418_p),
    .din1(g416_n),
    .din2(g417_n)
  );


  orX
  g_g418_n
  (
    .dout(g418_n),
    .din1(g416_p),
    .din2(g417_p)
  );


  andX
  g_g419_p
  (
    .dout(g419_p),
    .din1(g415_p),
    .din2(g418_n)
  );


  andX
  g_g420_p
  (
    .dout(g420_p),
    .din1(g415_n),
    .din2(g418_p)
  );


  orX
  g_g421_n
  (
    .dout(g421_n),
    .din1(g419_p),
    .din2(g420_p)
  );


  andX
  g_g422_p
  (
    .dout(g422_p),
    .din1(ffc_145_p),
    .din2(ffc_153_p_spl_00)
  );


  orX
  g_g422_n
  (
    .dout(g422_n),
    .din1(ffc_145_n),
    .din2(ffc_153_n_spl_00)
  );


  andX
  g_g423_p
  (
    .dout(g423_p),
    .din1(ffc_158_n_spl_0),
    .din2(ffc_159_p_spl_0)
  );


  orX
  g_g423_n
  (
    .dout(g423_n),
    .din1(ffc_158_p_spl_0),
    .din2(ffc_159_n_spl_0)
  );


  andX
  g_g424_p
  (
    .dout(g424_p),
    .din1(ffc_158_p_spl_0),
    .din2(ffc_159_n_spl_0)
  );


  orX
  g_g424_n
  (
    .dout(g424_n),
    .din1(ffc_158_n_spl_0),
    .din2(ffc_159_p_spl_0)
  );


  andX
  g_g425_p
  (
    .dout(g425_p),
    .din1(g423_n),
    .din2(g424_n)
  );


  orX
  g_g425_n
  (
    .dout(g425_n),
    .din1(g423_p),
    .din2(g424_p)
  );


  orX
  g_g426_n
  (
    .dout(g426_n),
    .din1(g422_p),
    .din2(g425_p)
  );


  orX
  g_g427_n
  (
    .dout(g427_n),
    .din1(g422_n),
    .din2(g425_n)
  );


  andX
  g_g428_p
  (
    .dout(g428_p),
    .din1(g426_n),
    .din2(g427_n)
  );


  orX
  g_g429_n
  (
    .dout(g429_n),
    .din1(g421_n_spl_),
    .din2(g428_p_spl_)
  );


  andX
  g_g430_p
  (
    .dout(g430_p),
    .din1(g421_n_spl_),
    .din2(g428_p_spl_)
  );


  andX
  g_g431_p
  (
    .dout(g431_p),
    .din1(ffc_91_p_spl_0),
    .din2(ffc_95_n_spl_)
  );


  orX
  g_g431_n
  (
    .dout(g431_n),
    .din1(ffc_91_n_spl_),
    .din2(ffc_95_p_spl_0)
  );


  andX
  g_g432_p
  (
    .dout(g432_p),
    .din1(ffc_91_n_spl_),
    .din2(ffc_95_p_spl_0)
  );


  orX
  g_g432_n
  (
    .dout(g432_n),
    .din1(ffc_91_p_spl_0),
    .din2(ffc_95_n_spl_)
  );


  andX
  g_g433_p
  (
    .dout(g433_p),
    .din1(g431_n),
    .din2(g432_n)
  );


  orX
  g_g433_n
  (
    .dout(g433_n),
    .din1(g431_p),
    .din2(g432_p)
  );


  andX
  g_g434_p
  (
    .dout(g434_p),
    .din1(ffc_99_p_spl_0),
    .din2(ffc_103_n_spl_)
  );


  orX
  g_g434_n
  (
    .dout(g434_n),
    .din1(ffc_99_n_spl_),
    .din2(ffc_103_p_spl_0)
  );


  andX
  g_g435_p
  (
    .dout(g435_p),
    .din1(ffc_99_n_spl_),
    .din2(ffc_103_p_spl_0)
  );


  orX
  g_g435_n
  (
    .dout(g435_n),
    .din1(ffc_99_p_spl_0),
    .din2(ffc_103_n_spl_)
  );


  andX
  g_g436_p
  (
    .dout(g436_p),
    .din1(g434_n),
    .din2(g435_n)
  );


  orX
  g_g436_n
  (
    .dout(g436_n),
    .din1(g434_p),
    .din2(g435_p)
  );


  andX
  g_g437_p
  (
    .dout(g437_p),
    .din1(g433_p),
    .din2(g436_n)
  );


  andX
  g_g438_p
  (
    .dout(g438_p),
    .din1(g433_n),
    .din2(g436_p)
  );


  orX
  g_g439_n
  (
    .dout(g439_n),
    .din1(g437_p),
    .din2(g438_p)
  );


  andX
  g_g440_p
  (
    .dout(g440_p),
    .din1(ffc_146_p),
    .din2(ffc_153_p_spl_00)
  );


  orX
  g_g440_n
  (
    .dout(g440_n),
    .din1(ffc_146_n),
    .din2(ffc_153_n_spl_00)
  );


  andX
  g_g441_p
  (
    .dout(g441_p),
    .din1(ffc_160_p_spl_0),
    .din2(ffc_161_n_spl_0)
  );


  orX
  g_g441_n
  (
    .dout(g441_n),
    .din1(ffc_160_n_spl_0),
    .din2(ffc_161_p_spl_0)
  );


  andX
  g_g442_p
  (
    .dout(g442_p),
    .din1(ffc_160_n_spl_0),
    .din2(ffc_161_p_spl_0)
  );


  orX
  g_g442_n
  (
    .dout(g442_n),
    .din1(ffc_160_p_spl_0),
    .din2(ffc_161_n_spl_0)
  );


  andX
  g_g443_p
  (
    .dout(g443_p),
    .din1(g441_n),
    .din2(g442_n)
  );


  orX
  g_g443_n
  (
    .dout(g443_n),
    .din1(g441_p),
    .din2(g442_p)
  );


  orX
  g_g444_n
  (
    .dout(g444_n),
    .din1(g440_p),
    .din2(g443_p)
  );


  orX
  g_g445_n
  (
    .dout(g445_n),
    .din1(g440_n),
    .din2(g443_n)
  );


  andX
  g_g446_p
  (
    .dout(g446_p),
    .din1(g444_n),
    .din2(g445_n)
  );


  orX
  g_g447_n
  (
    .dout(g447_n),
    .din1(g439_n_spl_),
    .din2(g446_p_spl_)
  );


  andX
  g_g448_p
  (
    .dout(g448_p),
    .din1(g439_n_spl_),
    .din2(g446_p_spl_)
  );


  andX
  g_g449_p
  (
    .dout(g449_p),
    .din1(ffc_92_p_spl_0),
    .din2(ffc_96_n_spl_)
  );


  orX
  g_g449_n
  (
    .dout(g449_n),
    .din1(ffc_92_n_spl_),
    .din2(ffc_96_p_spl_0)
  );


  andX
  g_g450_p
  (
    .dout(g450_p),
    .din1(ffc_92_n_spl_),
    .din2(ffc_96_p_spl_0)
  );


  orX
  g_g450_n
  (
    .dout(g450_n),
    .din1(ffc_92_p_spl_0),
    .din2(ffc_96_n_spl_)
  );


  andX
  g_g451_p
  (
    .dout(g451_p),
    .din1(g449_n),
    .din2(g450_n)
  );


  orX
  g_g451_n
  (
    .dout(g451_n),
    .din1(g449_p),
    .din2(g450_p)
  );


  andX
  g_g452_p
  (
    .dout(g452_p),
    .din1(ffc_100_p_spl_0),
    .din2(ffc_104_n_spl_)
  );


  orX
  g_g452_n
  (
    .dout(g452_n),
    .din1(ffc_100_n_spl_),
    .din2(ffc_104_p_spl_0)
  );


  andX
  g_g453_p
  (
    .dout(g453_p),
    .din1(ffc_100_n_spl_),
    .din2(ffc_104_p_spl_0)
  );


  orX
  g_g453_n
  (
    .dout(g453_n),
    .din1(ffc_100_p_spl_0),
    .din2(ffc_104_n_spl_)
  );


  andX
  g_g454_p
  (
    .dout(g454_p),
    .din1(g452_n),
    .din2(g453_n)
  );


  orX
  g_g454_n
  (
    .dout(g454_n),
    .din1(g452_p),
    .din2(g453_p)
  );


  andX
  g_g455_p
  (
    .dout(g455_p),
    .din1(g451_p),
    .din2(g454_n)
  );


  andX
  g_g456_p
  (
    .dout(g456_p),
    .din1(g451_n),
    .din2(g454_p)
  );


  orX
  g_g457_n
  (
    .dout(g457_n),
    .din1(g455_p),
    .din2(g456_p)
  );


  andX
  g_g458_p
  (
    .dout(g458_p),
    .din1(ffc_147_p),
    .din2(ffc_153_p_spl_01)
  );


  orX
  g_g458_n
  (
    .dout(g458_n),
    .din1(ffc_147_n),
    .din2(ffc_153_n_spl_01)
  );


  andX
  g_g459_p
  (
    .dout(g459_p),
    .din1(ffc_158_n_spl_1),
    .din2(ffc_160_p_spl_1)
  );


  orX
  g_g459_n
  (
    .dout(g459_n),
    .din1(ffc_158_p_spl_1),
    .din2(ffc_160_n_spl_1)
  );


  andX
  g_g460_p
  (
    .dout(g460_p),
    .din1(ffc_158_p_spl_1),
    .din2(ffc_160_n_spl_1)
  );


  orX
  g_g460_n
  (
    .dout(g460_n),
    .din1(ffc_158_n_spl_1),
    .din2(ffc_160_p_spl_1)
  );


  andX
  g_g461_p
  (
    .dout(g461_p),
    .din1(g459_n),
    .din2(g460_n)
  );


  orX
  g_g461_n
  (
    .dout(g461_n),
    .din1(g459_p),
    .din2(g460_p)
  );


  orX
  g_g462_n
  (
    .dout(g462_n),
    .din1(g458_p),
    .din2(g461_p)
  );


  orX
  g_g463_n
  (
    .dout(g463_n),
    .din1(g458_n),
    .din2(g461_n)
  );


  andX
  g_g464_p
  (
    .dout(g464_p),
    .din1(g462_n),
    .din2(g463_n)
  );


  orX
  g_g465_n
  (
    .dout(g465_n),
    .din1(g457_n_spl_),
    .din2(g464_p_spl_)
  );


  andX
  g_g466_p
  (
    .dout(g466_p),
    .din1(g457_n_spl_),
    .din2(g464_p_spl_)
  );


  andX
  g_g467_p
  (
    .dout(g467_p),
    .din1(ffc_93_p_spl_0),
    .din2(ffc_97_n_spl_)
  );


  orX
  g_g467_n
  (
    .dout(g467_n),
    .din1(ffc_93_n_spl_),
    .din2(ffc_97_p_spl_0)
  );


  andX
  g_g468_p
  (
    .dout(g468_p),
    .din1(ffc_93_n_spl_),
    .din2(ffc_97_p_spl_0)
  );


  orX
  g_g468_n
  (
    .dout(g468_n),
    .din1(ffc_93_p_spl_0),
    .din2(ffc_97_n_spl_)
  );


  andX
  g_g469_p
  (
    .dout(g469_p),
    .din1(g467_n),
    .din2(g468_n)
  );


  orX
  g_g469_n
  (
    .dout(g469_n),
    .din1(g467_p),
    .din2(g468_p)
  );


  andX
  g_g470_p
  (
    .dout(g470_p),
    .din1(ffc_101_p_spl_0),
    .din2(ffc_105_n_spl_)
  );


  orX
  g_g470_n
  (
    .dout(g470_n),
    .din1(ffc_101_n_spl_),
    .din2(ffc_105_p_spl_0)
  );


  andX
  g_g471_p
  (
    .dout(g471_p),
    .din1(ffc_101_n_spl_),
    .din2(ffc_105_p_spl_0)
  );


  orX
  g_g471_n
  (
    .dout(g471_n),
    .din1(ffc_101_p_spl_0),
    .din2(ffc_105_n_spl_)
  );


  andX
  g_g472_p
  (
    .dout(g472_p),
    .din1(g470_n),
    .din2(g471_n)
  );


  orX
  g_g472_n
  (
    .dout(g472_n),
    .din1(g470_p),
    .din2(g471_p)
  );


  andX
  g_g473_p
  (
    .dout(g473_p),
    .din1(g469_p),
    .din2(g472_n)
  );


  andX
  g_g474_p
  (
    .dout(g474_p),
    .din1(g469_n),
    .din2(g472_p)
  );


  orX
  g_g475_n
  (
    .dout(g475_n),
    .din1(g473_p),
    .din2(g474_p)
  );


  andX
  g_g476_p
  (
    .dout(g476_p),
    .din1(ffc_148_p),
    .din2(ffc_153_p_spl_01)
  );


  orX
  g_g476_n
  (
    .dout(g476_n),
    .din1(ffc_148_n),
    .din2(ffc_153_n_spl_01)
  );


  andX
  g_g477_p
  (
    .dout(g477_p),
    .din1(ffc_159_n_spl_1),
    .din2(ffc_161_p_spl_1)
  );


  orX
  g_g477_n
  (
    .dout(g477_n),
    .din1(ffc_159_p_spl_1),
    .din2(ffc_161_n_spl_1)
  );


  andX
  g_g478_p
  (
    .dout(g478_p),
    .din1(ffc_159_p_spl_1),
    .din2(ffc_161_n_spl_1)
  );


  orX
  g_g478_n
  (
    .dout(g478_n),
    .din1(ffc_159_n_spl_1),
    .din2(ffc_161_p_spl_1)
  );


  andX
  g_g479_p
  (
    .dout(g479_p),
    .din1(g477_n),
    .din2(g478_n)
  );


  orX
  g_g479_n
  (
    .dout(g479_n),
    .din1(g477_p),
    .din2(g478_p)
  );


  orX
  g_g480_n
  (
    .dout(g480_n),
    .din1(g476_p),
    .din2(g479_p)
  );


  orX
  g_g481_n
  (
    .dout(g481_n),
    .din1(g476_n),
    .din2(g479_n)
  );


  andX
  g_g482_p
  (
    .dout(g482_p),
    .din1(g480_n),
    .din2(g481_n)
  );


  orX
  g_g483_n
  (
    .dout(g483_n),
    .din1(g475_n_spl_),
    .din2(g482_p_spl_)
  );


  andX
  g_g484_p
  (
    .dout(g484_p),
    .din1(g475_n_spl_),
    .din2(g482_p_spl_)
  );


  andX
  g_g485_p
  (
    .dout(g485_p),
    .din1(ffc_106_p_spl_0),
    .din2(ffc_110_n_spl_)
  );


  orX
  g_g485_n
  (
    .dout(g485_n),
    .din1(ffc_106_n_spl_),
    .din2(ffc_110_p_spl_0)
  );


  andX
  g_g486_p
  (
    .dout(g486_p),
    .din1(ffc_106_n_spl_),
    .din2(ffc_110_p_spl_0)
  );


  orX
  g_g486_n
  (
    .dout(g486_n),
    .din1(ffc_106_p_spl_0),
    .din2(ffc_110_n_spl_)
  );


  andX
  g_g487_p
  (
    .dout(g487_p),
    .din1(g485_n),
    .din2(g486_n)
  );


  orX
  g_g487_n
  (
    .dout(g487_n),
    .din1(g485_p),
    .din2(g486_p)
  );


  andX
  g_g488_p
  (
    .dout(g488_p),
    .din1(ffc_114_p_spl_0),
    .din2(ffc_118_n_spl_)
  );


  orX
  g_g488_n
  (
    .dout(g488_n),
    .din1(ffc_114_n_spl_),
    .din2(ffc_118_p_spl_0)
  );


  andX
  g_g489_p
  (
    .dout(g489_p),
    .din1(ffc_114_n_spl_),
    .din2(ffc_118_p_spl_0)
  );


  orX
  g_g489_n
  (
    .dout(g489_n),
    .din1(ffc_114_p_spl_0),
    .din2(ffc_118_n_spl_)
  );


  andX
  g_g490_p
  (
    .dout(g490_p),
    .din1(g488_n),
    .din2(g489_n)
  );


  orX
  g_g490_n
  (
    .dout(g490_n),
    .din1(g488_p),
    .din2(g489_p)
  );


  andX
  g_g491_p
  (
    .dout(g491_p),
    .din1(g487_p),
    .din2(g490_n)
  );


  andX
  g_g492_p
  (
    .dout(g492_p),
    .din1(g487_n),
    .din2(g490_p)
  );


  orX
  g_g493_n
  (
    .dout(g493_n),
    .din1(g491_p),
    .din2(g492_p)
  );


  andX
  g_g494_p
  (
    .dout(g494_p),
    .din1(ffc_149_p),
    .din2(ffc_153_p_spl_10)
  );


  orX
  g_g494_n
  (
    .dout(g494_n),
    .din1(ffc_149_n),
    .din2(ffc_153_n_spl_10)
  );


  andX
  g_g495_p
  (
    .dout(g495_p),
    .din1(ffc_154_n_spl_0),
    .din2(ffc_155_p_spl_0)
  );


  orX
  g_g495_n
  (
    .dout(g495_n),
    .din1(ffc_154_p_spl_0),
    .din2(ffc_155_n_spl_0)
  );


  andX
  g_g496_p
  (
    .dout(g496_p),
    .din1(ffc_154_p_spl_0),
    .din2(ffc_155_n_spl_0)
  );


  orX
  g_g496_n
  (
    .dout(g496_n),
    .din1(ffc_154_n_spl_0),
    .din2(ffc_155_p_spl_0)
  );


  andX
  g_g497_p
  (
    .dout(g497_p),
    .din1(g495_n),
    .din2(g496_n)
  );


  orX
  g_g497_n
  (
    .dout(g497_n),
    .din1(g495_p),
    .din2(g496_p)
  );


  orX
  g_g498_n
  (
    .dout(g498_n),
    .din1(g494_p),
    .din2(g497_p)
  );


  orX
  g_g499_n
  (
    .dout(g499_n),
    .din1(g494_n),
    .din2(g497_n)
  );


  andX
  g_g500_p
  (
    .dout(g500_p),
    .din1(g498_n),
    .din2(g499_n)
  );


  orX
  g_g501_n
  (
    .dout(g501_n),
    .din1(g493_n_spl_),
    .din2(g500_p_spl_)
  );


  andX
  g_g502_p
  (
    .dout(g502_p),
    .din1(g493_n_spl_),
    .din2(g500_p_spl_)
  );


  andX
  g_g503_p
  (
    .dout(g503_p),
    .din1(ffc_107_p_spl_0),
    .din2(ffc_111_n_spl_)
  );


  orX
  g_g503_n
  (
    .dout(g503_n),
    .din1(ffc_107_n_spl_),
    .din2(ffc_111_p_spl_0)
  );


  andX
  g_g504_p
  (
    .dout(g504_p),
    .din1(ffc_107_n_spl_),
    .din2(ffc_111_p_spl_0)
  );


  orX
  g_g504_n
  (
    .dout(g504_n),
    .din1(ffc_107_p_spl_0),
    .din2(ffc_111_n_spl_)
  );


  andX
  g_g505_p
  (
    .dout(g505_p),
    .din1(g503_n),
    .din2(g504_n)
  );


  orX
  g_g505_n
  (
    .dout(g505_n),
    .din1(g503_p),
    .din2(g504_p)
  );


  andX
  g_g506_p
  (
    .dout(g506_p),
    .din1(ffc_115_p_spl_0),
    .din2(ffc_119_n_spl_)
  );


  orX
  g_g506_n
  (
    .dout(g506_n),
    .din1(ffc_115_n_spl_),
    .din2(ffc_119_p_spl_0)
  );


  andX
  g_g507_p
  (
    .dout(g507_p),
    .din1(ffc_115_n_spl_),
    .din2(ffc_119_p_spl_0)
  );


  orX
  g_g507_n
  (
    .dout(g507_n),
    .din1(ffc_115_p_spl_0),
    .din2(ffc_119_n_spl_)
  );


  andX
  g_g508_p
  (
    .dout(g508_p),
    .din1(g506_n),
    .din2(g507_n)
  );


  orX
  g_g508_n
  (
    .dout(g508_n),
    .din1(g506_p),
    .din2(g507_p)
  );


  andX
  g_g509_p
  (
    .dout(g509_p),
    .din1(g505_p),
    .din2(g508_n)
  );


  andX
  g_g510_p
  (
    .dout(g510_p),
    .din1(g505_n),
    .din2(g508_p)
  );


  orX
  g_g511_n
  (
    .dout(g511_n),
    .din1(g509_p),
    .din2(g510_p)
  );


  andX
  g_g512_p
  (
    .dout(g512_p),
    .din1(ffc_150_p),
    .din2(ffc_153_p_spl_10)
  );


  orX
  g_g512_n
  (
    .dout(g512_n),
    .din1(ffc_150_n),
    .din2(ffc_153_n_spl_10)
  );


  andX
  g_g513_p
  (
    .dout(g513_p),
    .din1(ffc_156_n_spl_0),
    .din2(ffc_157_p_spl_0)
  );


  orX
  g_g513_n
  (
    .dout(g513_n),
    .din1(ffc_156_p_spl_0),
    .din2(ffc_157_n_spl_0)
  );


  andX
  g_g514_p
  (
    .dout(g514_p),
    .din1(ffc_156_p_spl_0),
    .din2(ffc_157_n_spl_0)
  );


  orX
  g_g514_n
  (
    .dout(g514_n),
    .din1(ffc_156_n_spl_0),
    .din2(ffc_157_p_spl_0)
  );


  andX
  g_g515_p
  (
    .dout(g515_p),
    .din1(g513_n),
    .din2(g514_n)
  );


  orX
  g_g515_n
  (
    .dout(g515_n),
    .din1(g513_p),
    .din2(g514_p)
  );


  orX
  g_g516_n
  (
    .dout(g516_n),
    .din1(g512_p),
    .din2(g515_p)
  );


  orX
  g_g517_n
  (
    .dout(g517_n),
    .din1(g512_n),
    .din2(g515_n)
  );


  andX
  g_g518_p
  (
    .dout(g518_p),
    .din1(g516_n),
    .din2(g517_n)
  );


  orX
  g_g519_n
  (
    .dout(g519_n),
    .din1(g511_n_spl_),
    .din2(g518_p_spl_)
  );


  andX
  g_g520_p
  (
    .dout(g520_p),
    .din1(g511_n_spl_),
    .din2(g518_p_spl_)
  );


  andX
  g_g521_p
  (
    .dout(g521_p),
    .din1(ffc_108_p_spl_0),
    .din2(ffc_112_n_spl_)
  );


  orX
  g_g521_n
  (
    .dout(g521_n),
    .din1(ffc_108_n_spl_),
    .din2(ffc_112_p_spl_0)
  );


  andX
  g_g522_p
  (
    .dout(g522_p),
    .din1(ffc_108_n_spl_),
    .din2(ffc_112_p_spl_0)
  );


  orX
  g_g522_n
  (
    .dout(g522_n),
    .din1(ffc_108_p_spl_0),
    .din2(ffc_112_n_spl_)
  );


  andX
  g_g523_p
  (
    .dout(g523_p),
    .din1(g521_n),
    .din2(g522_n)
  );


  orX
  g_g523_n
  (
    .dout(g523_n),
    .din1(g521_p),
    .din2(g522_p)
  );


  andX
  g_g524_p
  (
    .dout(g524_p),
    .din1(ffc_116_p_spl_0),
    .din2(ffc_120_n_spl_)
  );


  orX
  g_g524_n
  (
    .dout(g524_n),
    .din1(ffc_116_n_spl_),
    .din2(ffc_120_p_spl_0)
  );


  andX
  g_g525_p
  (
    .dout(g525_p),
    .din1(ffc_116_n_spl_),
    .din2(ffc_120_p_spl_0)
  );


  orX
  g_g525_n
  (
    .dout(g525_n),
    .din1(ffc_116_p_spl_0),
    .din2(ffc_120_n_spl_)
  );


  andX
  g_g526_p
  (
    .dout(g526_p),
    .din1(g524_n),
    .din2(g525_n)
  );


  orX
  g_g526_n
  (
    .dout(g526_n),
    .din1(g524_p),
    .din2(g525_p)
  );


  andX
  g_g527_p
  (
    .dout(g527_p),
    .din1(g523_p),
    .din2(g526_n)
  );


  andX
  g_g528_p
  (
    .dout(g528_p),
    .din1(g523_n),
    .din2(g526_p)
  );


  orX
  g_g529_n
  (
    .dout(g529_n),
    .din1(g527_p),
    .din2(g528_p)
  );


  andX
  g_g530_p
  (
    .dout(g530_p),
    .din1(ffc_151_p),
    .din2(ffc_153_p_spl_11)
  );


  orX
  g_g530_n
  (
    .dout(g530_n),
    .din1(ffc_151_n),
    .din2(ffc_153_n_spl_11)
  );


  andX
  g_g531_p
  (
    .dout(g531_p),
    .din1(ffc_154_n_spl_1),
    .din2(ffc_156_p_spl_1)
  );


  orX
  g_g531_n
  (
    .dout(g531_n),
    .din1(ffc_154_p_spl_1),
    .din2(ffc_156_n_spl_1)
  );


  andX
  g_g532_p
  (
    .dout(g532_p),
    .din1(ffc_154_p_spl_1),
    .din2(ffc_156_n_spl_1)
  );


  orX
  g_g532_n
  (
    .dout(g532_n),
    .din1(ffc_154_n_spl_1),
    .din2(ffc_156_p_spl_1)
  );


  andX
  g_g533_p
  (
    .dout(g533_p),
    .din1(g531_n),
    .din2(g532_n)
  );


  orX
  g_g533_n
  (
    .dout(g533_n),
    .din1(g531_p),
    .din2(g532_p)
  );


  orX
  g_g534_n
  (
    .dout(g534_n),
    .din1(g530_p),
    .din2(g533_p)
  );


  orX
  g_g535_n
  (
    .dout(g535_n),
    .din1(g530_n),
    .din2(g533_n)
  );


  andX
  g_g536_p
  (
    .dout(g536_p),
    .din1(g534_n),
    .din2(g535_n)
  );


  orX
  g_g537_n
  (
    .dout(g537_n),
    .din1(g529_n_spl_),
    .din2(g536_p_spl_)
  );


  andX
  g_g538_p
  (
    .dout(g538_p),
    .din1(g529_n_spl_),
    .din2(g536_p_spl_)
  );


  andX
  g_g539_p
  (
    .dout(g539_p),
    .din1(ffc_109_p_spl_0),
    .din2(ffc_113_n_spl_)
  );


  orX
  g_g539_n
  (
    .dout(g539_n),
    .din1(ffc_109_n_spl_),
    .din2(ffc_113_p_spl_0)
  );


  andX
  g_g540_p
  (
    .dout(g540_p),
    .din1(ffc_109_n_spl_),
    .din2(ffc_113_p_spl_0)
  );


  orX
  g_g540_n
  (
    .dout(g540_n),
    .din1(ffc_109_p_spl_0),
    .din2(ffc_113_n_spl_)
  );


  andX
  g_g541_p
  (
    .dout(g541_p),
    .din1(g539_n),
    .din2(g540_n)
  );


  orX
  g_g541_n
  (
    .dout(g541_n),
    .din1(g539_p),
    .din2(g540_p)
  );


  andX
  g_g542_p
  (
    .dout(g542_p),
    .din1(ffc_117_p_spl_0),
    .din2(ffc_121_n_spl_)
  );


  orX
  g_g542_n
  (
    .dout(g542_n),
    .din1(ffc_117_n_spl_),
    .din2(ffc_121_p_spl_0)
  );


  andX
  g_g543_p
  (
    .dout(g543_p),
    .din1(ffc_117_n_spl_),
    .din2(ffc_121_p_spl_0)
  );


  orX
  g_g543_n
  (
    .dout(g543_n),
    .din1(ffc_117_p_spl_0),
    .din2(ffc_121_n_spl_)
  );


  andX
  g_g544_p
  (
    .dout(g544_p),
    .din1(g542_n),
    .din2(g543_n)
  );


  orX
  g_g544_n
  (
    .dout(g544_n),
    .din1(g542_p),
    .din2(g543_p)
  );


  andX
  g_g545_p
  (
    .dout(g545_p),
    .din1(g541_p),
    .din2(g544_n)
  );


  andX
  g_g546_p
  (
    .dout(g546_p),
    .din1(g541_n),
    .din2(g544_p)
  );


  orX
  g_g547_n
  (
    .dout(g547_n),
    .din1(g545_p),
    .din2(g546_p)
  );


  andX
  g_g548_p
  (
    .dout(g548_p),
    .din1(ffc_152_p),
    .din2(ffc_153_p_spl_11)
  );


  orX
  g_g548_n
  (
    .dout(g548_n),
    .din1(ffc_152_n),
    .din2(ffc_153_n_spl_11)
  );


  andX
  g_g549_p
  (
    .dout(g549_p),
    .din1(ffc_155_n_spl_1),
    .din2(ffc_157_p_spl_1)
  );


  orX
  g_g549_n
  (
    .dout(g549_n),
    .din1(ffc_155_p_spl_1),
    .din2(ffc_157_n_spl_1)
  );


  andX
  g_g550_p
  (
    .dout(g550_p),
    .din1(ffc_155_p_spl_1),
    .din2(ffc_157_n_spl_1)
  );


  orX
  g_g550_n
  (
    .dout(g550_n),
    .din1(ffc_155_n_spl_1),
    .din2(ffc_157_p_spl_1)
  );


  andX
  g_g551_p
  (
    .dout(g551_p),
    .din1(g549_n),
    .din2(g550_n)
  );


  orX
  g_g551_n
  (
    .dout(g551_n),
    .din1(g549_p),
    .din2(g550_p)
  );


  orX
  g_g552_n
  (
    .dout(g552_n),
    .din1(g548_p),
    .din2(g551_p)
  );


  orX
  g_g553_n
  (
    .dout(g553_n),
    .din1(g548_n),
    .din2(g551_n)
  );


  andX
  g_g554_p
  (
    .dout(g554_p),
    .din1(g552_n),
    .din2(g553_n)
  );


  orX
  g_g555_n
  (
    .dout(g555_n),
    .din1(g547_n_spl_),
    .din2(g554_p_spl_)
  );


  andX
  g_g556_p
  (
    .dout(g556_p),
    .din1(g547_n_spl_),
    .din2(g554_p_spl_)
  );


  andX
  g_g557_p
  (
    .dout(g557_p),
    .din1(ffc_162_p_spl_0),
    .din2(ffc_163_n_spl_)
  );


  orX
  g_g557_n
  (
    .dout(g557_n),
    .din1(ffc_162_n_spl_),
    .din2(ffc_163_p_spl_0)
  );


  andX
  g_g558_p
  (
    .dout(g558_p),
    .din1(ffc_162_n_spl_),
    .din2(ffc_163_p_spl_0)
  );


  orX
  g_g558_n
  (
    .dout(g558_n),
    .din1(ffc_162_p_spl_0),
    .din2(ffc_163_n_spl_)
  );


  andX
  g_g559_p
  (
    .dout(g559_p),
    .din1(g557_n),
    .din2(g558_n)
  );


  orX
  g_g559_n
  (
    .dout(g559_n),
    .din1(g557_p),
    .din2(g558_p)
  );


  andX
  g_g560_p
  (
    .dout(g560_p),
    .din1(ffc_164_p_spl_0),
    .din2(ffc_165_n_spl_)
  );


  orX
  g_g560_n
  (
    .dout(g560_n),
    .din1(ffc_164_n_spl_),
    .din2(ffc_165_p_spl_0)
  );


  andX
  g_g561_p
  (
    .dout(g561_p),
    .din1(ffc_164_n_spl_),
    .din2(ffc_165_p_spl_0)
  );


  orX
  g_g561_n
  (
    .dout(g561_n),
    .din1(ffc_164_p_spl_0),
    .din2(ffc_165_n_spl_)
  );


  andX
  g_g562_p
  (
    .dout(g562_p),
    .din1(g560_n),
    .din2(g561_n)
  );


  orX
  g_g562_n
  (
    .dout(g562_n),
    .din1(g560_p),
    .din2(g561_p)
  );


  andX
  g_g563_p
  (
    .dout(g563_p),
    .din1(g559_p),
    .din2(g562_n)
  );


  andX
  g_g564_p
  (
    .dout(g564_p),
    .din1(g559_n),
    .din2(g562_p)
  );


  orX
  g_g565_n
  (
    .dout(g565_n),
    .din1(g563_p),
    .din2(g564_p)
  );


  andX
  g_g566_p
  (
    .dout(g566_p),
    .din1(ffc_166_p_spl_0),
    .din2(ffc_167_n_spl_)
  );


  orX
  g_g566_n
  (
    .dout(g566_n),
    .din1(ffc_166_n_spl_),
    .din2(ffc_167_p_spl_0)
  );


  andX
  g_g567_p
  (
    .dout(g567_p),
    .din1(ffc_166_n_spl_),
    .din2(ffc_167_p_spl_0)
  );


  orX
  g_g567_n
  (
    .dout(g567_n),
    .din1(ffc_166_p_spl_0),
    .din2(ffc_167_n_spl_)
  );


  andX
  g_g568_p
  (
    .dout(g568_p),
    .din1(g566_n),
    .din2(g567_n)
  );


  orX
  g_g568_n
  (
    .dout(g568_n),
    .din1(g566_p),
    .din2(g567_p)
  );


  andX
  g_g569_p
  (
    .dout(g569_p),
    .din1(ffc_168_p_spl_0),
    .din2(ffc_169_n_spl_)
  );


  orX
  g_g569_n
  (
    .dout(g569_n),
    .din1(ffc_168_n_spl_),
    .din2(ffc_169_p_spl_0)
  );


  andX
  g_g570_p
  (
    .dout(g570_p),
    .din1(ffc_168_n_spl_),
    .din2(ffc_169_p_spl_0)
  );


  orX
  g_g570_n
  (
    .dout(g570_n),
    .din1(ffc_168_p_spl_0),
    .din2(ffc_169_n_spl_)
  );


  andX
  g_g571_p
  (
    .dout(g571_p),
    .din1(g569_n),
    .din2(g570_n)
  );


  orX
  g_g571_n
  (
    .dout(g571_n),
    .din1(g569_p),
    .din2(g570_p)
  );


  andX
  g_g572_p
  (
    .dout(g572_p),
    .din1(g568_p),
    .din2(g571_n)
  );


  andX
  g_g573_p
  (
    .dout(g573_p),
    .din1(g568_n),
    .din2(g571_p)
  );


  orX
  g_g574_n
  (
    .dout(g574_n),
    .din1(g572_p),
    .din2(g573_p)
  );


  andX
  g_g575_p
  (
    .dout(g575_p),
    .din1(ffc_170_p_spl_0),
    .din2(ffc_171_n_spl_)
  );


  orX
  g_g575_n
  (
    .dout(g575_n),
    .din1(ffc_170_n_spl_),
    .din2(ffc_171_p_spl_0)
  );


  andX
  g_g576_p
  (
    .dout(g576_p),
    .din1(ffc_170_n_spl_),
    .din2(ffc_171_p_spl_0)
  );


  orX
  g_g576_n
  (
    .dout(g576_n),
    .din1(ffc_170_p_spl_0),
    .din2(ffc_171_n_spl_)
  );


  andX
  g_g577_p
  (
    .dout(g577_p),
    .din1(g575_n),
    .din2(g576_n)
  );


  orX
  g_g577_n
  (
    .dout(g577_n),
    .din1(g575_p),
    .din2(g576_p)
  );


  andX
  g_g578_p
  (
    .dout(g578_p),
    .din1(ffc_172_p_spl_0),
    .din2(ffc_173_n_spl_)
  );


  orX
  g_g578_n
  (
    .dout(g578_n),
    .din1(ffc_172_n_spl_),
    .din2(ffc_173_p_spl_0)
  );


  andX
  g_g579_p
  (
    .dout(g579_p),
    .din1(ffc_172_n_spl_),
    .din2(ffc_173_p_spl_0)
  );


  orX
  g_g579_n
  (
    .dout(g579_n),
    .din1(ffc_172_p_spl_0),
    .din2(ffc_173_n_spl_)
  );


  andX
  g_g580_p
  (
    .dout(g580_p),
    .din1(g578_n),
    .din2(g579_n)
  );


  orX
  g_g580_n
  (
    .dout(g580_n),
    .din1(g578_p),
    .din2(g579_p)
  );


  andX
  g_g581_p
  (
    .dout(g581_p),
    .din1(g577_p),
    .din2(g580_n)
  );


  andX
  g_g582_p
  (
    .dout(g582_p),
    .din1(g577_n),
    .din2(g580_p)
  );


  orX
  g_g583_n
  (
    .dout(g583_n),
    .din1(g581_p),
    .din2(g582_p)
  );


  andX
  g_g584_p
  (
    .dout(g584_p),
    .din1(ffc_174_p_spl_0),
    .din2(ffc_175_n_spl_)
  );


  orX
  g_g584_n
  (
    .dout(g584_n),
    .din1(ffc_174_n_spl_),
    .din2(ffc_175_p_spl_0)
  );


  andX
  g_g585_p
  (
    .dout(g585_p),
    .din1(ffc_174_n_spl_),
    .din2(ffc_175_p_spl_0)
  );


  orX
  g_g585_n
  (
    .dout(g585_n),
    .din1(ffc_174_p_spl_0),
    .din2(ffc_175_n_spl_)
  );


  andX
  g_g586_p
  (
    .dout(g586_p),
    .din1(g584_n),
    .din2(g585_n)
  );


  orX
  g_g586_n
  (
    .dout(g586_n),
    .din1(g584_p),
    .din2(g585_p)
  );


  andX
  g_g587_p
  (
    .dout(g587_p),
    .din1(ffc_176_p_spl_0),
    .din2(ffc_177_n_spl_)
  );


  orX
  g_g587_n
  (
    .dout(g587_n),
    .din1(ffc_176_n_spl_),
    .din2(ffc_177_p_spl_0)
  );


  andX
  g_g588_p
  (
    .dout(g588_p),
    .din1(ffc_176_n_spl_),
    .din2(ffc_177_p_spl_0)
  );


  orX
  g_g588_n
  (
    .dout(g588_n),
    .din1(ffc_176_p_spl_0),
    .din2(ffc_177_n_spl_)
  );


  andX
  g_g589_p
  (
    .dout(g589_p),
    .din1(g587_n),
    .din2(g588_n)
  );


  orX
  g_g589_n
  (
    .dout(g589_n),
    .din1(g587_p),
    .din2(g588_p)
  );


  andX
  g_g590_p
  (
    .dout(g590_p),
    .din1(g586_p),
    .din2(g589_n)
  );


  andX
  g_g591_p
  (
    .dout(g591_p),
    .din1(g586_n),
    .din2(g589_p)
  );


  orX
  g_g592_n
  (
    .dout(g592_n),
    .din1(g590_p),
    .din2(g591_p)
  );


  andX
  g_g593_p
  (
    .dout(g593_p),
    .din1(ffc_178_p_spl_0),
    .din2(ffc_179_n_spl_)
  );


  orX
  g_g593_n
  (
    .dout(g593_n),
    .din1(ffc_178_n_spl_),
    .din2(ffc_179_p_spl_0)
  );


  andX
  g_g594_p
  (
    .dout(g594_p),
    .din1(ffc_178_n_spl_),
    .din2(ffc_179_p_spl_0)
  );


  orX
  g_g594_n
  (
    .dout(g594_n),
    .din1(ffc_178_p_spl_0),
    .din2(ffc_179_n_spl_)
  );


  andX
  g_g595_p
  (
    .dout(g595_p),
    .din1(g593_n),
    .din2(g594_n)
  );


  orX
  g_g595_n
  (
    .dout(g595_n),
    .din1(g593_p),
    .din2(g594_p)
  );


  andX
  g_g596_p
  (
    .dout(g596_p),
    .din1(ffc_180_p_spl_0),
    .din2(ffc_181_n_spl_)
  );


  orX
  g_g596_n
  (
    .dout(g596_n),
    .din1(ffc_180_n_spl_),
    .din2(ffc_181_p_spl_0)
  );


  andX
  g_g597_p
  (
    .dout(g597_p),
    .din1(ffc_180_n_spl_),
    .din2(ffc_181_p_spl_0)
  );


  orX
  g_g597_n
  (
    .dout(g597_n),
    .din1(ffc_180_p_spl_0),
    .din2(ffc_181_n_spl_)
  );


  andX
  g_g598_p
  (
    .dout(g598_p),
    .din1(g596_n),
    .din2(g597_n)
  );


  orX
  g_g598_n
  (
    .dout(g598_n),
    .din1(g596_p),
    .din2(g597_p)
  );


  andX
  g_g599_p
  (
    .dout(g599_p),
    .din1(g595_p),
    .din2(g598_n)
  );


  andX
  g_g600_p
  (
    .dout(g600_p),
    .din1(g595_n),
    .din2(g598_p)
  );


  orX
  g_g601_n
  (
    .dout(g601_n),
    .din1(g599_p),
    .din2(g600_p)
  );


  andX
  g_g602_p
  (
    .dout(g602_p),
    .din1(ffc_182_p_spl_0),
    .din2(ffc_183_n_spl_)
  );


  orX
  g_g602_n
  (
    .dout(g602_n),
    .din1(ffc_182_n_spl_),
    .din2(ffc_183_p_spl_0)
  );


  andX
  g_g603_p
  (
    .dout(g603_p),
    .din1(ffc_182_n_spl_),
    .din2(ffc_183_p_spl_0)
  );


  orX
  g_g603_n
  (
    .dout(g603_n),
    .din1(ffc_182_p_spl_0),
    .din2(ffc_183_n_spl_)
  );


  andX
  g_g604_p
  (
    .dout(g604_p),
    .din1(g602_n),
    .din2(g603_n)
  );


  orX
  g_g604_n
  (
    .dout(g604_n),
    .din1(g602_p),
    .din2(g603_p)
  );


  andX
  g_g605_p
  (
    .dout(g605_p),
    .din1(ffc_184_p_spl_0),
    .din2(ffc_185_n_spl_)
  );


  orX
  g_g605_n
  (
    .dout(g605_n),
    .din1(ffc_184_n_spl_),
    .din2(ffc_185_p_spl_0)
  );


  andX
  g_g606_p
  (
    .dout(g606_p),
    .din1(ffc_184_n_spl_),
    .din2(ffc_185_p_spl_0)
  );


  orX
  g_g606_n
  (
    .dout(g606_n),
    .din1(ffc_184_p_spl_0),
    .din2(ffc_185_n_spl_)
  );


  andX
  g_g607_p
  (
    .dout(g607_p),
    .din1(g605_n),
    .din2(g606_n)
  );


  orX
  g_g607_n
  (
    .dout(g607_n),
    .din1(g605_p),
    .din2(g606_p)
  );


  andX
  g_g608_p
  (
    .dout(g608_p),
    .din1(g604_p),
    .din2(g607_n)
  );


  andX
  g_g609_p
  (
    .dout(g609_p),
    .din1(g604_n),
    .din2(g607_p)
  );


  orX
  g_g610_n
  (
    .dout(g610_n),
    .din1(g608_p),
    .din2(g609_p)
  );


  andX
  g_g611_p
  (
    .dout(g611_p),
    .din1(ffc_186_p_spl_0),
    .din2(ffc_187_n_spl_)
  );


  orX
  g_g611_n
  (
    .dout(g611_n),
    .din1(ffc_186_n_spl_),
    .din2(ffc_187_p_spl_0)
  );


  andX
  g_g612_p
  (
    .dout(g612_p),
    .din1(ffc_186_n_spl_),
    .din2(ffc_187_p_spl_0)
  );


  orX
  g_g612_n
  (
    .dout(g612_n),
    .din1(ffc_186_p_spl_0),
    .din2(ffc_187_n_spl_)
  );


  andX
  g_g613_p
  (
    .dout(g613_p),
    .din1(g611_n),
    .din2(g612_n)
  );


  orX
  g_g613_n
  (
    .dout(g613_n),
    .din1(g611_p),
    .din2(g612_p)
  );


  andX
  g_g614_p
  (
    .dout(g614_p),
    .din1(ffc_188_p_spl_0),
    .din2(ffc_189_n_spl_)
  );


  orX
  g_g614_n
  (
    .dout(g614_n),
    .din1(ffc_188_n_spl_),
    .din2(ffc_189_p_spl_0)
  );


  andX
  g_g615_p
  (
    .dout(g615_p),
    .din1(ffc_188_n_spl_),
    .din2(ffc_189_p_spl_0)
  );


  orX
  g_g615_n
  (
    .dout(g615_n),
    .din1(ffc_188_p_spl_0),
    .din2(ffc_189_n_spl_)
  );


  andX
  g_g616_p
  (
    .dout(g616_p),
    .din1(g614_n),
    .din2(g615_n)
  );


  orX
  g_g616_n
  (
    .dout(g616_n),
    .din1(g614_p),
    .din2(g615_p)
  );


  andX
  g_g617_p
  (
    .dout(g617_p),
    .din1(g613_p),
    .din2(g616_n)
  );


  andX
  g_g618_p
  (
    .dout(g618_p),
    .din1(g613_n),
    .din2(g616_p)
  );


  orX
  g_g619_n
  (
    .dout(g619_n),
    .din1(g617_p),
    .din2(g618_p)
  );


  andX
  g_g620_p
  (
    .dout(g620_p),
    .din1(ffc_190_p_spl_0),
    .din2(ffc_191_n_spl_)
  );


  orX
  g_g620_n
  (
    .dout(g620_n),
    .din1(ffc_190_n_spl_),
    .din2(ffc_191_p_spl_0)
  );


  andX
  g_g621_p
  (
    .dout(g621_p),
    .din1(ffc_190_n_spl_),
    .din2(ffc_191_p_spl_0)
  );


  orX
  g_g621_n
  (
    .dout(g621_n),
    .din1(ffc_190_p_spl_0),
    .din2(ffc_191_n_spl_)
  );


  andX
  g_g622_p
  (
    .dout(g622_p),
    .din1(g620_n),
    .din2(g621_n)
  );


  orX
  g_g622_n
  (
    .dout(g622_n),
    .din1(g620_p),
    .din2(g621_p)
  );


  andX
  g_g623_p
  (
    .dout(g623_p),
    .din1(ffc_192_p_spl_0),
    .din2(ffc_193_n_spl_)
  );


  orX
  g_g623_n
  (
    .dout(g623_n),
    .din1(ffc_192_n_spl_),
    .din2(ffc_193_p_spl_0)
  );


  andX
  g_g624_p
  (
    .dout(g624_p),
    .din1(ffc_192_n_spl_),
    .din2(ffc_193_p_spl_0)
  );


  orX
  g_g624_n
  (
    .dout(g624_n),
    .din1(ffc_192_p_spl_0),
    .din2(ffc_193_n_spl_)
  );


  andX
  g_g625_p
  (
    .dout(g625_p),
    .din1(g623_n),
    .din2(g624_n)
  );


  orX
  g_g625_n
  (
    .dout(g625_n),
    .din1(g623_p),
    .din2(g624_p)
  );


  andX
  g_g626_p
  (
    .dout(g626_p),
    .din1(g622_p),
    .din2(g625_n)
  );


  andX
  g_g627_p
  (
    .dout(g627_p),
    .din1(g622_n),
    .din2(g625_p)
  );


  orX
  g_g628_n
  (
    .dout(g628_n),
    .din1(g626_p),
    .din2(g627_p)
  );


  buf

  (
    G468_p,
    g242_n
  );


  buf

  (
    G469_p,
    g246_n
  );


  buf

  (
    G470_p,
    g250_n
  );


  buf

  (
    G471_p,
    g254_n
  );


  buf

  (
    G472_p,
    g260_n
  );


  buf

  (
    G473_p,
    g264_n
  );


  buf

  (
    G474_p,
    g268_n
  );


  buf

  (
    G475_p,
    g272_n
  );


  buf

  (
    G476_p,
    g278_n
  );


  buf

  (
    G477_p,
    g282_n
  );


  buf

  (
    G478_p,
    g286_n
  );


  buf

  (
    G479_p,
    g290_n
  );


  buf

  (
    G480_p,
    g296_n
  );


  buf

  (
    G481_p,
    g300_n
  );


  buf

  (
    G482_p,
    g304_n
  );


  buf

  (
    G483_p,
    g308_n
  );


  buf

  (
    G484_p,
    g314_n
  );


  buf

  (
    G485_p,
    g318_n
  );


  buf

  (
    G486_p,
    g322_n
  );


  buf

  (
    G487_p,
    g326_n
  );


  buf

  (
    G488_p,
    g332_n
  );


  buf

  (
    G489_p,
    g336_n
  );


  buf

  (
    G490_p,
    g340_n
  );


  buf

  (
    G491_p,
    g344_n
  );


  buf

  (
    G492_p,
    g350_n
  );


  buf

  (
    G493_p,
    g354_n
  );


  buf

  (
    G494_p,
    g358_n
  );


  buf

  (
    G495_p,
    g362_n
  );


  buf

  (
    G496_p,
    g368_n
  );


  buf

  (
    G497_p,
    g372_n
  );


  buf

  (
    G498_p,
    g376_n
  );


  buf

  (
    G499_p,
    g380_n
  );


  DROC
  ffc_0
  (
    .doutp(ffc_0_p),
    .doutn(ffc_0_n),
    .din(ffc_41_p)
  );


  DROC
  ffc_1
  (
    .doutp(ffc_1_p),
    .doutn(ffc_1_n),
    .din(ffc_42_p)
  );


  DROC
  ffc_2
  (
    .doutp(ffc_2_p),
    .doutn(ffc_2_n),
    .din(ffc_43_p)
  );


  DROC
  ffc_3
  (
    .doutp(ffc_3_p),
    .doutn(ffc_3_n),
    .din(ffc_44_p)
  );


  DROC
  ffc_4
  (
    .doutp(ffc_4_p),
    .doutn(ffc_4_n),
    .din(ffc_45_p)
  );


  DROC
  ffc_5
  (
    .doutp(ffc_5_p),
    .doutn(ffc_5_n),
    .din(ffc_46_p)
  );


  DROC
  ffc_6
  (
    .doutp(ffc_6_p),
    .doutn(ffc_6_n),
    .din(ffc_47_p)
  );


  DROC
  ffc_7
  (
    .doutp(ffc_7_p),
    .doutn(ffc_7_n),
    .din(ffc_48_p)
  );


  DROC
  ffc_8
  (
    .doutp(ffc_8_p),
    .doutn(ffc_8_n),
    .din(ffc_49_p)
  );


  DROC
  ffc_9
  (
    .doutp(ffc_9_p),
    .doutn(ffc_9_n),
    .din(ffc_50_p)
  );


  DROC
  ffc_10
  (
    .doutp(ffc_10_p),
    .doutn(ffc_10_n),
    .din(ffc_51_p)
  );


  DROC
  ffc_11
  (
    .doutp(ffc_11_p),
    .doutn(ffc_11_n),
    .din(ffc_52_p)
  );


  DROC
  ffc_12
  (
    .doutp(ffc_12_p),
    .doutn(ffc_12_n),
    .din(ffc_53_p)
  );


  DROC
  ffc_13
  (
    .doutp(ffc_13_p),
    .doutn(ffc_13_n),
    .din(ffc_54_p)
  );


  DROC
  ffc_14
  (
    .doutp(ffc_14_p),
    .doutn(ffc_14_n),
    .din(ffc_55_p)
  );


  DROC
  ffc_15
  (
    .doutp(ffc_15_p),
    .doutn(ffc_15_n),
    .din(ffc_56_p)
  );


  DROC
  ffc_16
  (
    .doutp(ffc_16_p),
    .doutn(ffc_16_n),
    .din(ffc_57_p)
  );


  DROC
  ffc_17
  (
    .doutp(ffc_17_p),
    .doutn(ffc_17_n),
    .din(ffc_58_p)
  );


  DROC
  ffc_18
  (
    .doutp(ffc_18_p),
    .doutn(ffc_18_n),
    .din(ffc_59_p)
  );


  DROC
  ffc_19
  (
    .doutp(ffc_19_p),
    .doutn(ffc_19_n),
    .din(ffc_60_p)
  );


  DROC
  ffc_20
  (
    .doutp(ffc_20_p),
    .doutn(ffc_20_n),
    .din(ffc_61_p)
  );


  DROC
  ffc_21
  (
    .doutp(ffc_21_p),
    .doutn(ffc_21_n),
    .din(ffc_62_p)
  );


  DROC
  ffc_22
  (
    .doutp(ffc_22_p),
    .doutn(ffc_22_n),
    .din(ffc_63_p)
  );


  DROC
  ffc_23
  (
    .doutp(ffc_23_p),
    .doutn(ffc_23_n),
    .din(ffc_64_p)
  );


  DROC
  ffc_24
  (
    .doutp(ffc_24_p),
    .doutn(ffc_24_n),
    .din(ffc_65_p)
  );


  DROC
  ffc_25
  (
    .doutp(ffc_25_p),
    .doutn(ffc_25_n),
    .din(ffc_66_p)
  );


  DROC
  ffc_26
  (
    .doutp(ffc_26_p),
    .doutn(ffc_26_n),
    .din(ffc_67_p)
  );


  DROC
  ffc_27
  (
    .doutp(ffc_27_p),
    .doutn(ffc_27_n),
    .din(ffc_68_p)
  );


  DROC
  ffc_28
  (
    .doutp(ffc_28_p),
    .doutn(ffc_28_n),
    .din(ffc_69_p)
  );


  DROC
  ffc_29
  (
    .doutp(ffc_29_p),
    .doutn(ffc_29_n),
    .din(ffc_70_p)
  );


  DROC
  ffc_30
  (
    .doutp(ffc_30_p),
    .doutn(ffc_30_n),
    .din(ffc_71_p)
  );


  DROC
  ffc_31
  (
    .doutp(ffc_31_p),
    .doutn(ffc_31_n),
    .din(ffc_72_p)
  );


  DROC
  ffc_32
  (
    .doutp(ffc_32_p),
    .doutn(ffc_32_n),
    .din(G33_p)
  );


  DROC
  ffc_33
  (
    .doutp(ffc_33_p),
    .doutn(ffc_33_n),
    .din(G34_p)
  );


  DROC
  ffc_34
  (
    .doutp(ffc_34_p),
    .doutn(ffc_34_n),
    .din(G35_p)
  );


  DROC
  ffc_35
  (
    .doutp(ffc_35_p),
    .doutn(ffc_35_n),
    .din(G36_p)
  );


  DROC
  ffc_36
  (
    .doutp(ffc_36_p),
    .doutn(ffc_36_n),
    .din(G37_p)
  );


  DROC
  ffc_37
  (
    .doutp(ffc_37_p),
    .doutn(ffc_37_n),
    .din(G38_p)
  );


  DROC
  ffc_38
  (
    .doutp(ffc_38_p),
    .doutn(ffc_38_n),
    .din(G39_p)
  );


  DROC
  ffc_39
  (
    .doutp(ffc_39_p),
    .doutn(ffc_39_n),
    .din(G40_p)
  );


  DROC
  ffc_40
  (
    .doutp(ffc_40_p),
    .doutn(ffc_40_n),
    .din(G41_p)
  );


  DROC
  ffc_41
  (
    .doutp(ffc_41_p),
    .doutn(ffc_41_n),
    .din(ffc_90_p_spl_)
  );


  DROC
  ffc_42
  (
    .doutp(ffc_42_p),
    .doutn(ffc_42_n),
    .din(ffc_91_p_spl_)
  );


  DROC
  ffc_43
  (
    .doutp(ffc_43_p),
    .doutn(ffc_43_n),
    .din(ffc_92_p_spl_)
  );


  DROC
  ffc_44
  (
    .doutp(ffc_44_p),
    .doutn(ffc_44_n),
    .din(ffc_93_p_spl_)
  );


  DROC
  ffc_45
  (
    .doutp(ffc_45_p),
    .doutn(ffc_45_n),
    .din(ffc_94_p_spl_)
  );


  DROC
  ffc_46
  (
    .doutp(ffc_46_p),
    .doutn(ffc_46_n),
    .din(ffc_95_p_spl_)
  );


  DROC
  ffc_47
  (
    .doutp(ffc_47_p),
    .doutn(ffc_47_n),
    .din(ffc_96_p_spl_)
  );


  DROC
  ffc_48
  (
    .doutp(ffc_48_p),
    .doutn(ffc_48_n),
    .din(ffc_97_p_spl_)
  );


  DROC
  ffc_49
  (
    .doutp(ffc_49_p),
    .doutn(ffc_49_n),
    .din(ffc_98_p_spl_)
  );


  DROC
  ffc_50
  (
    .doutp(ffc_50_p),
    .doutn(ffc_50_n),
    .din(ffc_99_p_spl_)
  );


  DROC
  ffc_51
  (
    .doutp(ffc_51_p),
    .doutn(ffc_51_n),
    .din(ffc_100_p_spl_)
  );


  DROC
  ffc_52
  (
    .doutp(ffc_52_p),
    .doutn(ffc_52_n),
    .din(ffc_101_p_spl_)
  );


  DROC
  ffc_53
  (
    .doutp(ffc_53_p),
    .doutn(ffc_53_n),
    .din(ffc_102_p_spl_)
  );


  DROC
  ffc_54
  (
    .doutp(ffc_54_p),
    .doutn(ffc_54_n),
    .din(ffc_103_p_spl_)
  );


  DROC
  ffc_55
  (
    .doutp(ffc_55_p),
    .doutn(ffc_55_n),
    .din(ffc_104_p_spl_)
  );


  DROC
  ffc_56
  (
    .doutp(ffc_56_p),
    .doutn(ffc_56_n),
    .din(ffc_105_p_spl_)
  );


  DROC
  ffc_57
  (
    .doutp(ffc_57_p),
    .doutn(ffc_57_n),
    .din(ffc_106_p_spl_)
  );


  DROC
  ffc_58
  (
    .doutp(ffc_58_p),
    .doutn(ffc_58_n),
    .din(ffc_107_p_spl_)
  );


  DROC
  ffc_59
  (
    .doutp(ffc_59_p),
    .doutn(ffc_59_n),
    .din(ffc_108_p_spl_)
  );


  DROC
  ffc_60
  (
    .doutp(ffc_60_p),
    .doutn(ffc_60_n),
    .din(ffc_109_p_spl_)
  );


  DROC
  ffc_61
  (
    .doutp(ffc_61_p),
    .doutn(ffc_61_n),
    .din(ffc_110_p_spl_)
  );


  DROC
  ffc_62
  (
    .doutp(ffc_62_p),
    .doutn(ffc_62_n),
    .din(ffc_111_p_spl_)
  );


  DROC
  ffc_63
  (
    .doutp(ffc_63_p),
    .doutn(ffc_63_n),
    .din(ffc_112_p_spl_)
  );


  DROC
  ffc_64
  (
    .doutp(ffc_64_p),
    .doutn(ffc_64_n),
    .din(ffc_113_p_spl_)
  );


  DROC
  ffc_65
  (
    .doutp(ffc_65_p),
    .doutn(ffc_65_n),
    .din(ffc_114_p_spl_)
  );


  DROC
  ffc_66
  (
    .doutp(ffc_66_p),
    .doutn(ffc_66_n),
    .din(ffc_115_p_spl_)
  );


  DROC
  ffc_67
  (
    .doutp(ffc_67_p),
    .doutn(ffc_67_n),
    .din(ffc_116_p_spl_)
  );


  DROC
  ffc_68
  (
    .doutp(ffc_68_p),
    .doutn(ffc_68_n),
    .din(ffc_117_p_spl_)
  );


  DROC
  ffc_69
  (
    .doutp(ffc_69_p),
    .doutn(ffc_69_n),
    .din(ffc_118_p_spl_)
  );


  DROC
  ffc_70
  (
    .doutp(ffc_70_p),
    .doutn(ffc_70_n),
    .din(ffc_119_p_spl_)
  );


  DROC
  ffc_71
  (
    .doutp(ffc_71_p),
    .doutn(ffc_71_n),
    .din(ffc_120_p_spl_)
  );


  DROC
  ffc_72
  (
    .doutp(ffc_72_p),
    .doutn(ffc_72_n),
    .din(ffc_121_p_spl_)
  );


  DROC
  ffc_73
  (
    .doutp(ffc_73_p),
    .doutn(ffc_73_n),
    .din(g381_n_spl_)
  );


  DROC
  ffc_74
  (
    .doutp(ffc_74_p),
    .doutn(ffc_74_n),
    .din(g382_n_spl_)
  );


  DROC
  ffc_75
  (
    .doutp(ffc_75_p),
    .doutn(ffc_75_n),
    .din(g383_n_spl_)
  );


  DROC
  ffc_76
  (
    .doutp(ffc_76_p),
    .doutn(ffc_76_n),
    .din(g384_n_spl_)
  );


  DROC
  ffc_77
  (
    .doutp(ffc_77_p),
    .doutn(ffc_77_n),
    .din(g385_n_spl_)
  );


  DROC
  ffc_78
  (
    .doutp(ffc_78_p),
    .doutn(ffc_78_n),
    .din(g386_n_spl_)
  );


  DROC
  ffc_79
  (
    .doutp(ffc_79_p),
    .doutn(ffc_79_n),
    .din(g387_n_spl_)
  );


  DROC
  ffc_80
  (
    .doutp(ffc_80_p),
    .doutn(ffc_80_n),
    .din(g388_n_spl_)
  );


  DROC
  ffc_81
  (
    .doutp(ffc_81_n),
    .doutn(ffc_81_p),
    .din(g389_n_spl_)
  );


  DROC
  ffc_82
  (
    .doutp(ffc_82_n),
    .doutn(ffc_82_p),
    .din(g390_n_spl_)
  );


  DROC
  ffc_83
  (
    .doutp(ffc_83_n),
    .doutn(ffc_83_p),
    .din(g391_n_spl_)
  );


  DROC
  ffc_84
  (
    .doutp(ffc_84_p),
    .doutn(ffc_84_n),
    .din(g392_n_spl_)
  );


  DROC
  ffc_85
  (
    .doutp(ffc_85_n),
    .doutn(ffc_85_p),
    .din(g393_n_spl_)
  );


  DROC
  ffc_86
  (
    .doutp(ffc_86_n),
    .doutn(ffc_86_p),
    .din(g394_n_spl_)
  );


  DROC
  ffc_87
  (
    .doutp(ffc_87_n),
    .doutn(ffc_87_p),
    .din(g396_n_spl_)
  );


  DROC
  ffc_88
  (
    .doutp(ffc_88_n),
    .doutn(ffc_88_p),
    .din(g397_n_spl_)
  );


  DROC
  ffc_89
  (
    .doutp(ffc_89_p),
    .doutn(ffc_89_n),
    .din(g398_n_spl_)
  );


  DROC
  ffc_90
  (
    .doutp(ffc_90_p),
    .doutn(ffc_90_n),
    .din(ffc_162_p_spl_)
  );


  DROC
  ffc_91
  (
    .doutp(ffc_91_p),
    .doutn(ffc_91_n),
    .din(ffc_163_p_spl_)
  );


  DROC
  ffc_92
  (
    .doutp(ffc_92_p),
    .doutn(ffc_92_n),
    .din(ffc_164_p_spl_)
  );


  DROC
  ffc_93
  (
    .doutp(ffc_93_p),
    .doutn(ffc_93_n),
    .din(ffc_165_p_spl_)
  );


  DROC
  ffc_94
  (
    .doutp(ffc_94_p),
    .doutn(ffc_94_n),
    .din(ffc_166_p_spl_)
  );


  DROC
  ffc_95
  (
    .doutp(ffc_95_p),
    .doutn(ffc_95_n),
    .din(ffc_167_p_spl_)
  );


  DROC
  ffc_96
  (
    .doutp(ffc_96_p),
    .doutn(ffc_96_n),
    .din(ffc_168_p_spl_)
  );


  DROC
  ffc_97
  (
    .doutp(ffc_97_p),
    .doutn(ffc_97_n),
    .din(ffc_169_p_spl_)
  );


  DROC
  ffc_98
  (
    .doutp(ffc_98_p),
    .doutn(ffc_98_n),
    .din(ffc_170_p_spl_)
  );


  DROC
  ffc_99
  (
    .doutp(ffc_99_p),
    .doutn(ffc_99_n),
    .din(ffc_171_p_spl_)
  );


  DROC
  ffc_100
  (
    .doutp(ffc_100_p),
    .doutn(ffc_100_n),
    .din(ffc_172_p_spl_)
  );


  DROC
  ffc_101
  (
    .doutp(ffc_101_p),
    .doutn(ffc_101_n),
    .din(ffc_173_p_spl_)
  );


  DROC
  ffc_102
  (
    .doutp(ffc_102_p),
    .doutn(ffc_102_n),
    .din(ffc_174_p_spl_)
  );


  DROC
  ffc_103
  (
    .doutp(ffc_103_p),
    .doutn(ffc_103_n),
    .din(ffc_175_p_spl_)
  );


  DROC
  ffc_104
  (
    .doutp(ffc_104_p),
    .doutn(ffc_104_n),
    .din(ffc_176_p_spl_)
  );


  DROC
  ffc_105
  (
    .doutp(ffc_105_p),
    .doutn(ffc_105_n),
    .din(ffc_177_p_spl_)
  );


  DROC
  ffc_106
  (
    .doutp(ffc_106_p),
    .doutn(ffc_106_n),
    .din(ffc_178_p_spl_)
  );


  DROC
  ffc_107
  (
    .doutp(ffc_107_p),
    .doutn(ffc_107_n),
    .din(ffc_179_p_spl_)
  );


  DROC
  ffc_108
  (
    .doutp(ffc_108_p),
    .doutn(ffc_108_n),
    .din(ffc_180_p_spl_)
  );


  DROC
  ffc_109
  (
    .doutp(ffc_109_p),
    .doutn(ffc_109_n),
    .din(ffc_181_p_spl_)
  );


  DROC
  ffc_110
  (
    .doutp(ffc_110_p),
    .doutn(ffc_110_n),
    .din(ffc_182_p_spl_)
  );


  DROC
  ffc_111
  (
    .doutp(ffc_111_p),
    .doutn(ffc_111_n),
    .din(ffc_183_p_spl_)
  );


  DROC
  ffc_112
  (
    .doutp(ffc_112_p),
    .doutn(ffc_112_n),
    .din(ffc_184_p_spl_)
  );


  DROC
  ffc_113
  (
    .doutp(ffc_113_p),
    .doutn(ffc_113_n),
    .din(ffc_185_p_spl_)
  );


  DROC
  ffc_114
  (
    .doutp(ffc_114_p),
    .doutn(ffc_114_n),
    .din(ffc_186_p_spl_)
  );


  DROC
  ffc_115
  (
    .doutp(ffc_115_p),
    .doutn(ffc_115_n),
    .din(ffc_187_p_spl_)
  );


  DROC
  ffc_116
  (
    .doutp(ffc_116_p),
    .doutn(ffc_116_n),
    .din(ffc_188_p_spl_)
  );


  DROC
  ffc_117
  (
    .doutp(ffc_117_p),
    .doutn(ffc_117_n),
    .din(ffc_189_p_spl_)
  );


  DROC
  ffc_118
  (
    .doutp(ffc_118_p),
    .doutn(ffc_118_n),
    .din(ffc_190_p_spl_)
  );


  DROC
  ffc_119
  (
    .doutp(ffc_119_p),
    .doutn(ffc_119_n),
    .din(ffc_191_p_spl_)
  );


  DROC
  ffc_120
  (
    .doutp(ffc_120_p),
    .doutn(ffc_120_n),
    .din(ffc_192_p_spl_)
  );


  DROC
  ffc_121
  (
    .doutp(ffc_121_p),
    .doutn(ffc_121_n),
    .din(ffc_193_p_spl_)
  );


  DROC
  ffc_122
  (
    .doutp(ffc_122_n),
    .doutn(ffc_122_p),
    .din(g401_n)
  );


  DROC
  ffc_123
  (
    .doutp(ffc_123_n),
    .doutn(ffc_123_p),
    .din(g403_n)
  );


  DROC
  ffc_124
  (
    .doutp(ffc_124_p),
    .doutn(ffc_124_n),
    .din(g404_p)
  );


  DROC
  ffc_125
  (
    .doutp(ffc_125_p),
    .doutn(ffc_125_n),
    .din(g405_p)
  );


  DROC
  ffc_126
  (
    .doutp(ffc_126_p),
    .doutn(ffc_126_n),
    .din(g406_p)
  );


  DROC
  ffc_127
  (
    .doutp(ffc_127_p),
    .doutn(ffc_127_n),
    .din(g407_p)
  );


  DROC
  ffc_128
  (
    .doutp(ffc_128_p),
    .doutn(ffc_128_n),
    .din(g412_p)
  );


  DROC
  ffc_129
  (
    .doutp(ffc_129_n),
    .doutn(ffc_129_p),
    .din(g429_n)
  );


  DROC
  ffc_130
  (
    .doutp(ffc_130_p),
    .doutn(ffc_130_n),
    .din(g430_p)
  );


  DROC
  ffc_131
  (
    .doutp(ffc_131_n),
    .doutn(ffc_131_p),
    .din(g447_n)
  );


  DROC
  ffc_132
  (
    .doutp(ffc_132_p),
    .doutn(ffc_132_n),
    .din(g448_p)
  );


  DROC
  ffc_133
  (
    .doutp(ffc_133_n),
    .doutn(ffc_133_p),
    .din(g465_n)
  );


  DROC
  ffc_134
  (
    .doutp(ffc_134_p),
    .doutn(ffc_134_n),
    .din(g466_p)
  );


  DROC
  ffc_135
  (
    .doutp(ffc_135_n),
    .doutn(ffc_135_p),
    .din(g483_n)
  );


  DROC
  ffc_136
  (
    .doutp(ffc_136_p),
    .doutn(ffc_136_n),
    .din(g484_p)
  );


  DROC
  ffc_137
  (
    .doutp(ffc_137_n),
    .doutn(ffc_137_p),
    .din(g501_n)
  );


  DROC
  ffc_138
  (
    .doutp(ffc_138_p),
    .doutn(ffc_138_n),
    .din(g502_p)
  );


  DROC
  ffc_139
  (
    .doutp(ffc_139_n),
    .doutn(ffc_139_p),
    .din(g519_n)
  );


  DROC
  ffc_140
  (
    .doutp(ffc_140_p),
    .doutn(ffc_140_n),
    .din(g520_p)
  );


  DROC
  ffc_141
  (
    .doutp(ffc_141_n),
    .doutn(ffc_141_p),
    .din(g537_n)
  );


  DROC
  ffc_142
  (
    .doutp(ffc_142_p),
    .doutn(ffc_142_n),
    .din(g538_p)
  );


  DROC
  ffc_143
  (
    .doutp(ffc_143_n),
    .doutn(ffc_143_p),
    .din(g555_n)
  );


  DROC
  ffc_144
  (
    .doutp(ffc_144_p),
    .doutn(ffc_144_n),
    .din(g556_p)
  );


  DROC
  ffc_145
  (
    .doutp(ffc_145_p),
    .doutn(ffc_145_n),
    .din(ffc_32_p)
  );


  DROC
  ffc_146
  (
    .doutp(ffc_146_p),
    .doutn(ffc_146_n),
    .din(ffc_33_p)
  );


  DROC
  ffc_147
  (
    .doutp(ffc_147_p),
    .doutn(ffc_147_n),
    .din(ffc_34_p)
  );


  DROC
  ffc_148
  (
    .doutp(ffc_148_p),
    .doutn(ffc_148_n),
    .din(ffc_35_p)
  );


  DROC
  ffc_149
  (
    .doutp(ffc_149_p),
    .doutn(ffc_149_n),
    .din(ffc_36_p)
  );


  DROC
  ffc_150
  (
    .doutp(ffc_150_p),
    .doutn(ffc_150_n),
    .din(ffc_37_p)
  );


  DROC
  ffc_151
  (
    .doutp(ffc_151_p),
    .doutn(ffc_151_n),
    .din(ffc_38_p)
  );


  DROC
  ffc_152
  (
    .doutp(ffc_152_p),
    .doutn(ffc_152_n),
    .din(ffc_39_p)
  );


  DROC
  ffc_153
  (
    .doutp(ffc_153_p),
    .doutn(ffc_153_n),
    .din(ffc_40_p)
  );


  DROC
  ffc_154
  (
    .doutp(ffc_154_p),
    .doutn(ffc_154_n),
    .din(g565_n)
  );


  DROC
  ffc_155
  (
    .doutp(ffc_155_p),
    .doutn(ffc_155_n),
    .din(g574_n)
  );


  DROC
  ffc_156
  (
    .doutp(ffc_156_p),
    .doutn(ffc_156_n),
    .din(g583_n)
  );


  DROC
  ffc_157
  (
    .doutp(ffc_157_p),
    .doutn(ffc_157_n),
    .din(g592_n)
  );


  DROC
  ffc_158
  (
    .doutp(ffc_158_p),
    .doutn(ffc_158_n),
    .din(g601_n)
  );


  DROC
  ffc_159
  (
    .doutp(ffc_159_p),
    .doutn(ffc_159_n),
    .din(g610_n)
  );


  DROC
  ffc_160
  (
    .doutp(ffc_160_p),
    .doutn(ffc_160_n),
    .din(g619_n)
  );


  DROC
  ffc_161
  (
    .doutp(ffc_161_p),
    .doutn(ffc_161_n),
    .din(g628_n)
  );


  DROC
  ffc_162
  (
    .doutp(ffc_162_p),
    .doutn(ffc_162_n),
    .din(G1_p)
  );


  DROC
  ffc_163
  (
    .doutp(ffc_163_p),
    .doutn(ffc_163_n),
    .din(G2_p)
  );


  DROC
  ffc_164
  (
    .doutp(ffc_164_p),
    .doutn(ffc_164_n),
    .din(G3_p)
  );


  DROC
  ffc_165
  (
    .doutp(ffc_165_p),
    .doutn(ffc_165_n),
    .din(G4_p)
  );


  DROC
  ffc_166
  (
    .doutp(ffc_166_p),
    .doutn(ffc_166_n),
    .din(G5_p)
  );


  DROC
  ffc_167
  (
    .doutp(ffc_167_p),
    .doutn(ffc_167_n),
    .din(G6_p)
  );


  DROC
  ffc_168
  (
    .doutp(ffc_168_p),
    .doutn(ffc_168_n),
    .din(G7_p)
  );


  DROC
  ffc_169
  (
    .doutp(ffc_169_p),
    .doutn(ffc_169_n),
    .din(G8_p)
  );


  DROC
  ffc_170
  (
    .doutp(ffc_170_p),
    .doutn(ffc_170_n),
    .din(G9_p)
  );


  DROC
  ffc_171
  (
    .doutp(ffc_171_p),
    .doutn(ffc_171_n),
    .din(G10_p)
  );


  DROC
  ffc_172
  (
    .doutp(ffc_172_p),
    .doutn(ffc_172_n),
    .din(G11_p)
  );


  DROC
  ffc_173
  (
    .doutp(ffc_173_p),
    .doutn(ffc_173_n),
    .din(G12_p)
  );


  DROC
  ffc_174
  (
    .doutp(ffc_174_p),
    .doutn(ffc_174_n),
    .din(G13_p)
  );


  DROC
  ffc_175
  (
    .doutp(ffc_175_p),
    .doutn(ffc_175_n),
    .din(G14_p)
  );


  DROC
  ffc_176
  (
    .doutp(ffc_176_p),
    .doutn(ffc_176_n),
    .din(G15_p)
  );


  DROC
  ffc_177
  (
    .doutp(ffc_177_p),
    .doutn(ffc_177_n),
    .din(G16_p)
  );


  DROC
  ffc_178
  (
    .doutp(ffc_178_p),
    .doutn(ffc_178_n),
    .din(G17_p)
  );


  DROC
  ffc_179
  (
    .doutp(ffc_179_p),
    .doutn(ffc_179_n),
    .din(G18_p)
  );


  DROC
  ffc_180
  (
    .doutp(ffc_180_p),
    .doutn(ffc_180_n),
    .din(G19_p)
  );


  DROC
  ffc_181
  (
    .doutp(ffc_181_p),
    .doutn(ffc_181_n),
    .din(G20_p)
  );


  DROC
  ffc_182
  (
    .doutp(ffc_182_p),
    .doutn(ffc_182_n),
    .din(G21_p)
  );


  DROC
  ffc_183
  (
    .doutp(ffc_183_p),
    .doutn(ffc_183_n),
    .din(G22_p)
  );


  DROC
  ffc_184
  (
    .doutp(ffc_184_p),
    .doutn(ffc_184_n),
    .din(G23_p)
  );


  DROC
  ffc_185
  (
    .doutp(ffc_185_p),
    .doutn(ffc_185_n),
    .din(G24_p)
  );


  DROC
  ffc_186
  (
    .doutp(ffc_186_p),
    .doutn(ffc_186_n),
    .din(G25_p)
  );


  DROC
  ffc_187
  (
    .doutp(ffc_187_p),
    .doutn(ffc_187_n),
    .din(G26_p)
  );


  DROC
  ffc_188
  (
    .doutp(ffc_188_p),
    .doutn(ffc_188_n),
    .din(G27_p)
  );


  DROC
  ffc_189
  (
    .doutp(ffc_189_p),
    .doutn(ffc_189_n),
    .din(G28_p)
  );


  DROC
  ffc_190
  (
    .doutp(ffc_190_p),
    .doutn(ffc_190_n),
    .din(G29_p)
  );


  DROC
  ffc_191
  (
    .doutp(ffc_191_p),
    .doutn(ffc_191_n),
    .din(G30_p)
  );


  DROC
  ffc_192
  (
    .doutp(ffc_192_p),
    .doutn(ffc_192_n),
    .din(G31_p)
  );


  DROC
  ffc_193
  (
    .doutp(ffc_193_p),
    .doutn(ffc_193_n),
    .din(G32_p)
  );


  buf

  (
    g236_n_spl_,
    g236_n
  );


  buf

  (
    g236_n_spl_0,
    g236_n_spl_
  );


  buf

  (
    g236_n_spl_1,
    g236_n_spl_
  );


  buf

  (
    g236_p_spl_,
    g236_p
  );


  buf

  (
    g236_p_spl_0,
    g236_p_spl_
  );


  buf

  (
    g236_p_spl_1,
    g236_p_spl_
  );


  buf

  (
    ffc_73_p_spl_,
    ffc_73_p
  );


  buf

  (
    ffc_73_p_spl_0,
    ffc_73_p_spl_
  );


  buf

  (
    ffc_73_p_spl_1,
    ffc_73_p_spl_
  );


  buf

  (
    g238_p_spl_,
    g238_p
  );


  buf

  (
    g238_p_spl_0,
    g238_p_spl_
  );


  buf

  (
    g238_p_spl_1,
    g238_p_spl_
  );


  buf

  (
    ffc_73_n_spl_,
    ffc_73_n
  );


  buf

  (
    ffc_73_n_spl_0,
    ffc_73_n_spl_
  );


  buf

  (
    ffc_73_n_spl_1,
    ffc_73_n_spl_
  );


  buf

  (
    g238_n_spl_,
    g238_n
  );


  buf

  (
    g238_n_spl_0,
    g238_n_spl_
  );


  buf

  (
    g238_n_spl_1,
    g238_n_spl_
  );


  buf

  (
    ffc_74_p_spl_,
    ffc_74_p
  );


  buf

  (
    ffc_74_p_spl_0,
    ffc_74_p_spl_
  );


  buf

  (
    ffc_74_p_spl_00,
    ffc_74_p_spl_0
  );


  buf

  (
    ffc_74_p_spl_1,
    ffc_74_p_spl_
  );


  buf

  (
    ffc_74_n_spl_,
    ffc_74_n
  );


  buf

  (
    ffc_74_n_spl_0,
    ffc_74_n_spl_
  );


  buf

  (
    ffc_74_n_spl_00,
    ffc_74_n_spl_0
  );


  buf

  (
    ffc_74_n_spl_1,
    ffc_74_n_spl_
  );


  buf

  (
    ffc_75_p_spl_,
    ffc_75_p
  );


  buf

  (
    ffc_75_p_spl_0,
    ffc_75_p_spl_
  );


  buf

  (
    ffc_75_p_spl_00,
    ffc_75_p_spl_0
  );


  buf

  (
    ffc_75_p_spl_01,
    ffc_75_p_spl_0
  );


  buf

  (
    ffc_75_p_spl_1,
    ffc_75_p_spl_
  );


  buf

  (
    ffc_75_n_spl_,
    ffc_75_n
  );


  buf

  (
    ffc_75_n_spl_0,
    ffc_75_n_spl_
  );


  buf

  (
    ffc_75_n_spl_00,
    ffc_75_n_spl_0
  );


  buf

  (
    ffc_75_n_spl_01,
    ffc_75_n_spl_0
  );


  buf

  (
    ffc_75_n_spl_1,
    ffc_75_n_spl_
  );


  buf

  (
    ffc_76_p_spl_,
    ffc_76_p
  );


  buf

  (
    ffc_76_p_spl_0,
    ffc_76_p_spl_
  );


  buf

  (
    ffc_76_p_spl_1,
    ffc_76_p_spl_
  );


  buf

  (
    ffc_76_n_spl_,
    ffc_76_n
  );


  buf

  (
    ffc_76_n_spl_0,
    ffc_76_n_spl_
  );


  buf

  (
    ffc_76_n_spl_1,
    ffc_76_n_spl_
  );


  buf

  (
    g256_p_spl_,
    g256_p
  );


  buf

  (
    g256_p_spl_0,
    g256_p_spl_
  );


  buf

  (
    g256_p_spl_1,
    g256_p_spl_
  );


  buf

  (
    g256_n_spl_,
    g256_n
  );


  buf

  (
    g256_n_spl_0,
    g256_n_spl_
  );


  buf

  (
    g256_n_spl_1,
    g256_n_spl_
  );


  buf

  (
    g274_p_spl_,
    g274_p
  );


  buf

  (
    g274_p_spl_0,
    g274_p_spl_
  );


  buf

  (
    g274_p_spl_1,
    g274_p_spl_
  );


  buf

  (
    g274_n_spl_,
    g274_n
  );


  buf

  (
    g274_n_spl_0,
    g274_n_spl_
  );


  buf

  (
    g274_n_spl_1,
    g274_n_spl_
  );


  buf

  (
    g292_p_spl_,
    g292_p
  );


  buf

  (
    g292_p_spl_0,
    g292_p_spl_
  );


  buf

  (
    g292_p_spl_1,
    g292_p_spl_
  );


  buf

  (
    g292_n_spl_,
    g292_n
  );


  buf

  (
    g292_n_spl_0,
    g292_n_spl_
  );


  buf

  (
    g292_n_spl_1,
    g292_n_spl_
  );


  buf

  (
    ffc_128_p_spl_,
    ffc_128_p
  );


  buf

  (
    ffc_128_p_spl_0,
    ffc_128_p_spl_
  );


  buf

  (
    ffc_128_p_spl_1,
    ffc_128_p_spl_
  );


  buf

  (
    ffc_128_n_spl_,
    ffc_128_n
  );


  buf

  (
    ffc_128_n_spl_0,
    ffc_128_n_spl_
  );


  buf

  (
    ffc_128_n_spl_1,
    ffc_128_n_spl_
  );


  buf

  (
    ffc_77_p_spl_,
    ffc_77_p
  );


  buf

  (
    ffc_77_p_spl_0,
    ffc_77_p_spl_
  );


  buf

  (
    ffc_77_p_spl_1,
    ffc_77_p_spl_
  );


  buf

  (
    g310_p_spl_,
    g310_p
  );


  buf

  (
    g310_p_spl_0,
    g310_p_spl_
  );


  buf

  (
    g310_p_spl_1,
    g310_p_spl_
  );


  buf

  (
    ffc_77_n_spl_,
    ffc_77_n
  );


  buf

  (
    ffc_77_n_spl_0,
    ffc_77_n_spl_
  );


  buf

  (
    ffc_77_n_spl_1,
    ffc_77_n_spl_
  );


  buf

  (
    g310_n_spl_,
    g310_n
  );


  buf

  (
    g310_n_spl_0,
    g310_n_spl_
  );


  buf

  (
    g310_n_spl_1,
    g310_n_spl_
  );


  buf

  (
    ffc_78_p_spl_,
    ffc_78_p
  );


  buf

  (
    ffc_78_p_spl_0,
    ffc_78_p_spl_
  );


  buf

  (
    ffc_78_p_spl_1,
    ffc_78_p_spl_
  );


  buf

  (
    ffc_78_n_spl_,
    ffc_78_n
  );


  buf

  (
    ffc_78_n_spl_0,
    ffc_78_n_spl_
  );


  buf

  (
    ffc_78_n_spl_1,
    ffc_78_n_spl_
  );


  buf

  (
    ffc_79_p_spl_,
    ffc_79_p
  );


  buf

  (
    ffc_79_p_spl_0,
    ffc_79_p_spl_
  );


  buf

  (
    ffc_79_p_spl_1,
    ffc_79_p_spl_
  );


  buf

  (
    ffc_79_n_spl_,
    ffc_79_n
  );


  buf

  (
    ffc_79_n_spl_0,
    ffc_79_n_spl_
  );


  buf

  (
    ffc_79_n_spl_1,
    ffc_79_n_spl_
  );


  buf

  (
    ffc_80_p_spl_,
    ffc_80_p
  );


  buf

  (
    ffc_80_p_spl_0,
    ffc_80_p_spl_
  );


  buf

  (
    ffc_80_p_spl_1,
    ffc_80_p_spl_
  );


  buf

  (
    ffc_80_n_spl_,
    ffc_80_n
  );


  buf

  (
    ffc_80_n_spl_0,
    ffc_80_n_spl_
  );


  buf

  (
    ffc_80_n_spl_1,
    ffc_80_n_spl_
  );


  buf

  (
    g328_p_spl_,
    g328_p
  );


  buf

  (
    g328_p_spl_0,
    g328_p_spl_
  );


  buf

  (
    g328_p_spl_1,
    g328_p_spl_
  );


  buf

  (
    g328_n_spl_,
    g328_n
  );


  buf

  (
    g328_n_spl_0,
    g328_n_spl_
  );


  buf

  (
    g328_n_spl_1,
    g328_n_spl_
  );


  buf

  (
    g346_p_spl_,
    g346_p
  );


  buf

  (
    g346_p_spl_0,
    g346_p_spl_
  );


  buf

  (
    g346_p_spl_1,
    g346_p_spl_
  );


  buf

  (
    g346_n_spl_,
    g346_n
  );


  buf

  (
    g346_n_spl_0,
    g346_n_spl_
  );


  buf

  (
    g346_n_spl_1,
    g346_n_spl_
  );


  buf

  (
    g364_p_spl_,
    g364_p
  );


  buf

  (
    g364_p_spl_0,
    g364_p_spl_
  );


  buf

  (
    g364_p_spl_1,
    g364_p_spl_
  );


  buf

  (
    g364_n_spl_,
    g364_n
  );


  buf

  (
    g364_n_spl_0,
    g364_n_spl_
  );


  buf

  (
    g364_n_spl_1,
    g364_n_spl_
  );


  buf

  (
    g382_n_spl_,
    g382_n
  );


  buf

  (
    g382_n_spl_0,
    g382_n_spl_
  );


  buf

  (
    g383_n_spl_,
    g383_n
  );


  buf

  (
    g383_n_spl_0,
    g383_n_spl_
  );


  buf

  (
    g385_p_spl_,
    g385_p
  );


  buf

  (
    g385_p_spl_0,
    g385_p_spl_
  );


  buf

  (
    g388_p_spl_,
    g388_p
  );


  buf

  (
    g388_p_spl_0,
    g388_p_spl_
  );


  buf

  (
    g385_n_spl_,
    g385_n
  );


  buf

  (
    g385_n_spl_0,
    g385_n_spl_
  );


  buf

  (
    g388_n_spl_,
    g388_n
  );


  buf

  (
    g388_n_spl_0,
    g388_n_spl_
  );


  buf

  (
    g386_p_spl_,
    g386_p
  );


  buf

  (
    g386_p_spl_0,
    g386_p_spl_
  );


  buf

  (
    g387_p_spl_,
    g387_p
  );


  buf

  (
    g387_p_spl_0,
    g387_p_spl_
  );


  buf

  (
    g381_n_spl_,
    g381_n
  );


  buf

  (
    g381_n_spl_0,
    g381_n_spl_
  );


  buf

  (
    g390_n_spl_,
    g390_n
  );


  buf

  (
    g384_n_spl_,
    g384_n
  );


  buf

  (
    g384_n_spl_0,
    g384_n_spl_
  );


  buf

  (
    g395_n_spl_,
    g395_n
  );


  buf

  (
    g389_n_spl_,
    g389_n
  );


  buf

  (
    g386_n_spl_,
    g386_n
  );


  buf

  (
    g386_n_spl_0,
    g386_n_spl_
  );


  buf

  (
    g387_n_spl_,
    g387_n
  );


  buf

  (
    g387_n_spl_0,
    g387_n_spl_
  );


  buf

  (
    g394_n_spl_,
    g394_n
  );


  buf

  (
    g396_n_spl_,
    g396_n
  );


  buf

  (
    g397_n_spl_,
    g397_n
  );


  buf

  (
    g391_n_spl_,
    g391_n
  );


  buf

  (
    g392_n_spl_,
    g392_n
  );


  buf

  (
    g398_n_spl_,
    g398_n
  );


  buf

  (
    g393_n_spl_,
    g393_n
  );


  buf

  (
    ffc_90_p_spl_,
    ffc_90_p
  );


  buf

  (
    ffc_90_p_spl_0,
    ffc_90_p_spl_
  );


  buf

  (
    ffc_94_n_spl_,
    ffc_94_n
  );


  buf

  (
    ffc_90_n_spl_,
    ffc_90_n
  );


  buf

  (
    ffc_94_p_spl_,
    ffc_94_p
  );


  buf

  (
    ffc_94_p_spl_0,
    ffc_94_p_spl_
  );


  buf

  (
    ffc_98_p_spl_,
    ffc_98_p
  );


  buf

  (
    ffc_98_p_spl_0,
    ffc_98_p_spl_
  );


  buf

  (
    ffc_102_n_spl_,
    ffc_102_n
  );


  buf

  (
    ffc_98_n_spl_,
    ffc_98_n
  );


  buf

  (
    ffc_102_p_spl_,
    ffc_102_p
  );


  buf

  (
    ffc_102_p_spl_0,
    ffc_102_p_spl_
  );


  buf

  (
    ffc_153_p_spl_,
    ffc_153_p
  );


  buf

  (
    ffc_153_p_spl_0,
    ffc_153_p_spl_
  );


  buf

  (
    ffc_153_p_spl_00,
    ffc_153_p_spl_0
  );


  buf

  (
    ffc_153_p_spl_01,
    ffc_153_p_spl_0
  );


  buf

  (
    ffc_153_p_spl_1,
    ffc_153_p_spl_
  );


  buf

  (
    ffc_153_p_spl_10,
    ffc_153_p_spl_1
  );


  buf

  (
    ffc_153_p_spl_11,
    ffc_153_p_spl_1
  );


  buf

  (
    ffc_153_n_spl_,
    ffc_153_n
  );


  buf

  (
    ffc_153_n_spl_0,
    ffc_153_n_spl_
  );


  buf

  (
    ffc_153_n_spl_00,
    ffc_153_n_spl_0
  );


  buf

  (
    ffc_153_n_spl_01,
    ffc_153_n_spl_0
  );


  buf

  (
    ffc_153_n_spl_1,
    ffc_153_n_spl_
  );


  buf

  (
    ffc_153_n_spl_10,
    ffc_153_n_spl_1
  );


  buf

  (
    ffc_153_n_spl_11,
    ffc_153_n_spl_1
  );


  buf

  (
    ffc_158_n_spl_,
    ffc_158_n
  );


  buf

  (
    ffc_158_n_spl_0,
    ffc_158_n_spl_
  );


  buf

  (
    ffc_158_n_spl_1,
    ffc_158_n_spl_
  );


  buf

  (
    ffc_159_p_spl_,
    ffc_159_p
  );


  buf

  (
    ffc_159_p_spl_0,
    ffc_159_p_spl_
  );


  buf

  (
    ffc_159_p_spl_1,
    ffc_159_p_spl_
  );


  buf

  (
    ffc_158_p_spl_,
    ffc_158_p
  );


  buf

  (
    ffc_158_p_spl_0,
    ffc_158_p_spl_
  );


  buf

  (
    ffc_158_p_spl_1,
    ffc_158_p_spl_
  );


  buf

  (
    ffc_159_n_spl_,
    ffc_159_n
  );


  buf

  (
    ffc_159_n_spl_0,
    ffc_159_n_spl_
  );


  buf

  (
    ffc_159_n_spl_1,
    ffc_159_n_spl_
  );


  buf

  (
    g421_n_spl_,
    g421_n
  );


  buf

  (
    g428_p_spl_,
    g428_p
  );


  buf

  (
    ffc_91_p_spl_,
    ffc_91_p
  );


  buf

  (
    ffc_91_p_spl_0,
    ffc_91_p_spl_
  );


  buf

  (
    ffc_95_n_spl_,
    ffc_95_n
  );


  buf

  (
    ffc_91_n_spl_,
    ffc_91_n
  );


  buf

  (
    ffc_95_p_spl_,
    ffc_95_p
  );


  buf

  (
    ffc_95_p_spl_0,
    ffc_95_p_spl_
  );


  buf

  (
    ffc_99_p_spl_,
    ffc_99_p
  );


  buf

  (
    ffc_99_p_spl_0,
    ffc_99_p_spl_
  );


  buf

  (
    ffc_103_n_spl_,
    ffc_103_n
  );


  buf

  (
    ffc_99_n_spl_,
    ffc_99_n
  );


  buf

  (
    ffc_103_p_spl_,
    ffc_103_p
  );


  buf

  (
    ffc_103_p_spl_0,
    ffc_103_p_spl_
  );


  buf

  (
    ffc_160_p_spl_,
    ffc_160_p
  );


  buf

  (
    ffc_160_p_spl_0,
    ffc_160_p_spl_
  );


  buf

  (
    ffc_160_p_spl_1,
    ffc_160_p_spl_
  );


  buf

  (
    ffc_161_n_spl_,
    ffc_161_n
  );


  buf

  (
    ffc_161_n_spl_0,
    ffc_161_n_spl_
  );


  buf

  (
    ffc_161_n_spl_1,
    ffc_161_n_spl_
  );


  buf

  (
    ffc_160_n_spl_,
    ffc_160_n
  );


  buf

  (
    ffc_160_n_spl_0,
    ffc_160_n_spl_
  );


  buf

  (
    ffc_160_n_spl_1,
    ffc_160_n_spl_
  );


  buf

  (
    ffc_161_p_spl_,
    ffc_161_p
  );


  buf

  (
    ffc_161_p_spl_0,
    ffc_161_p_spl_
  );


  buf

  (
    ffc_161_p_spl_1,
    ffc_161_p_spl_
  );


  buf

  (
    g439_n_spl_,
    g439_n
  );


  buf

  (
    g446_p_spl_,
    g446_p
  );


  buf

  (
    ffc_92_p_spl_,
    ffc_92_p
  );


  buf

  (
    ffc_92_p_spl_0,
    ffc_92_p_spl_
  );


  buf

  (
    ffc_96_n_spl_,
    ffc_96_n
  );


  buf

  (
    ffc_92_n_spl_,
    ffc_92_n
  );


  buf

  (
    ffc_96_p_spl_,
    ffc_96_p
  );


  buf

  (
    ffc_96_p_spl_0,
    ffc_96_p_spl_
  );


  buf

  (
    ffc_100_p_spl_,
    ffc_100_p
  );


  buf

  (
    ffc_100_p_spl_0,
    ffc_100_p_spl_
  );


  buf

  (
    ffc_104_n_spl_,
    ffc_104_n
  );


  buf

  (
    ffc_100_n_spl_,
    ffc_100_n
  );


  buf

  (
    ffc_104_p_spl_,
    ffc_104_p
  );


  buf

  (
    ffc_104_p_spl_0,
    ffc_104_p_spl_
  );


  buf

  (
    g457_n_spl_,
    g457_n
  );


  buf

  (
    g464_p_spl_,
    g464_p
  );


  buf

  (
    ffc_93_p_spl_,
    ffc_93_p
  );


  buf

  (
    ffc_93_p_spl_0,
    ffc_93_p_spl_
  );


  buf

  (
    ffc_97_n_spl_,
    ffc_97_n
  );


  buf

  (
    ffc_93_n_spl_,
    ffc_93_n
  );


  buf

  (
    ffc_97_p_spl_,
    ffc_97_p
  );


  buf

  (
    ffc_97_p_spl_0,
    ffc_97_p_spl_
  );


  buf

  (
    ffc_101_p_spl_,
    ffc_101_p
  );


  buf

  (
    ffc_101_p_spl_0,
    ffc_101_p_spl_
  );


  buf

  (
    ffc_105_n_spl_,
    ffc_105_n
  );


  buf

  (
    ffc_101_n_spl_,
    ffc_101_n
  );


  buf

  (
    ffc_105_p_spl_,
    ffc_105_p
  );


  buf

  (
    ffc_105_p_spl_0,
    ffc_105_p_spl_
  );


  buf

  (
    g475_n_spl_,
    g475_n
  );


  buf

  (
    g482_p_spl_,
    g482_p
  );


  buf

  (
    ffc_106_p_spl_,
    ffc_106_p
  );


  buf

  (
    ffc_106_p_spl_0,
    ffc_106_p_spl_
  );


  buf

  (
    ffc_110_n_spl_,
    ffc_110_n
  );


  buf

  (
    ffc_106_n_spl_,
    ffc_106_n
  );


  buf

  (
    ffc_110_p_spl_,
    ffc_110_p
  );


  buf

  (
    ffc_110_p_spl_0,
    ffc_110_p_spl_
  );


  buf

  (
    ffc_114_p_spl_,
    ffc_114_p
  );


  buf

  (
    ffc_114_p_spl_0,
    ffc_114_p_spl_
  );


  buf

  (
    ffc_118_n_spl_,
    ffc_118_n
  );


  buf

  (
    ffc_114_n_spl_,
    ffc_114_n
  );


  buf

  (
    ffc_118_p_spl_,
    ffc_118_p
  );


  buf

  (
    ffc_118_p_spl_0,
    ffc_118_p_spl_
  );


  buf

  (
    ffc_154_n_spl_,
    ffc_154_n
  );


  buf

  (
    ffc_154_n_spl_0,
    ffc_154_n_spl_
  );


  buf

  (
    ffc_154_n_spl_1,
    ffc_154_n_spl_
  );


  buf

  (
    ffc_155_p_spl_,
    ffc_155_p
  );


  buf

  (
    ffc_155_p_spl_0,
    ffc_155_p_spl_
  );


  buf

  (
    ffc_155_p_spl_1,
    ffc_155_p_spl_
  );


  buf

  (
    ffc_154_p_spl_,
    ffc_154_p
  );


  buf

  (
    ffc_154_p_spl_0,
    ffc_154_p_spl_
  );


  buf

  (
    ffc_154_p_spl_1,
    ffc_154_p_spl_
  );


  buf

  (
    ffc_155_n_spl_,
    ffc_155_n
  );


  buf

  (
    ffc_155_n_spl_0,
    ffc_155_n_spl_
  );


  buf

  (
    ffc_155_n_spl_1,
    ffc_155_n_spl_
  );


  buf

  (
    g493_n_spl_,
    g493_n
  );


  buf

  (
    g500_p_spl_,
    g500_p
  );


  buf

  (
    ffc_107_p_spl_,
    ffc_107_p
  );


  buf

  (
    ffc_107_p_spl_0,
    ffc_107_p_spl_
  );


  buf

  (
    ffc_111_n_spl_,
    ffc_111_n
  );


  buf

  (
    ffc_107_n_spl_,
    ffc_107_n
  );


  buf

  (
    ffc_111_p_spl_,
    ffc_111_p
  );


  buf

  (
    ffc_111_p_spl_0,
    ffc_111_p_spl_
  );


  buf

  (
    ffc_115_p_spl_,
    ffc_115_p
  );


  buf

  (
    ffc_115_p_spl_0,
    ffc_115_p_spl_
  );


  buf

  (
    ffc_119_n_spl_,
    ffc_119_n
  );


  buf

  (
    ffc_115_n_spl_,
    ffc_115_n
  );


  buf

  (
    ffc_119_p_spl_,
    ffc_119_p
  );


  buf

  (
    ffc_119_p_spl_0,
    ffc_119_p_spl_
  );


  buf

  (
    ffc_156_n_spl_,
    ffc_156_n
  );


  buf

  (
    ffc_156_n_spl_0,
    ffc_156_n_spl_
  );


  buf

  (
    ffc_156_n_spl_1,
    ffc_156_n_spl_
  );


  buf

  (
    ffc_157_p_spl_,
    ffc_157_p
  );


  buf

  (
    ffc_157_p_spl_0,
    ffc_157_p_spl_
  );


  buf

  (
    ffc_157_p_spl_1,
    ffc_157_p_spl_
  );


  buf

  (
    ffc_156_p_spl_,
    ffc_156_p
  );


  buf

  (
    ffc_156_p_spl_0,
    ffc_156_p_spl_
  );


  buf

  (
    ffc_156_p_spl_1,
    ffc_156_p_spl_
  );


  buf

  (
    ffc_157_n_spl_,
    ffc_157_n
  );


  buf

  (
    ffc_157_n_spl_0,
    ffc_157_n_spl_
  );


  buf

  (
    ffc_157_n_spl_1,
    ffc_157_n_spl_
  );


  buf

  (
    g511_n_spl_,
    g511_n
  );


  buf

  (
    g518_p_spl_,
    g518_p
  );


  buf

  (
    ffc_108_p_spl_,
    ffc_108_p
  );


  buf

  (
    ffc_108_p_spl_0,
    ffc_108_p_spl_
  );


  buf

  (
    ffc_112_n_spl_,
    ffc_112_n
  );


  buf

  (
    ffc_108_n_spl_,
    ffc_108_n
  );


  buf

  (
    ffc_112_p_spl_,
    ffc_112_p
  );


  buf

  (
    ffc_112_p_spl_0,
    ffc_112_p_spl_
  );


  buf

  (
    ffc_116_p_spl_,
    ffc_116_p
  );


  buf

  (
    ffc_116_p_spl_0,
    ffc_116_p_spl_
  );


  buf

  (
    ffc_120_n_spl_,
    ffc_120_n
  );


  buf

  (
    ffc_116_n_spl_,
    ffc_116_n
  );


  buf

  (
    ffc_120_p_spl_,
    ffc_120_p
  );


  buf

  (
    ffc_120_p_spl_0,
    ffc_120_p_spl_
  );


  buf

  (
    g529_n_spl_,
    g529_n
  );


  buf

  (
    g536_p_spl_,
    g536_p
  );


  buf

  (
    ffc_109_p_spl_,
    ffc_109_p
  );


  buf

  (
    ffc_109_p_spl_0,
    ffc_109_p_spl_
  );


  buf

  (
    ffc_113_n_spl_,
    ffc_113_n
  );


  buf

  (
    ffc_109_n_spl_,
    ffc_109_n
  );


  buf

  (
    ffc_113_p_spl_,
    ffc_113_p
  );


  buf

  (
    ffc_113_p_spl_0,
    ffc_113_p_spl_
  );


  buf

  (
    ffc_117_p_spl_,
    ffc_117_p
  );


  buf

  (
    ffc_117_p_spl_0,
    ffc_117_p_spl_
  );


  buf

  (
    ffc_121_n_spl_,
    ffc_121_n
  );


  buf

  (
    ffc_117_n_spl_,
    ffc_117_n
  );


  buf

  (
    ffc_121_p_spl_,
    ffc_121_p
  );


  buf

  (
    ffc_121_p_spl_0,
    ffc_121_p_spl_
  );


  buf

  (
    g547_n_spl_,
    g547_n
  );


  buf

  (
    g554_p_spl_,
    g554_p
  );


  buf

  (
    ffc_162_p_spl_,
    ffc_162_p
  );


  buf

  (
    ffc_162_p_spl_0,
    ffc_162_p_spl_
  );


  buf

  (
    ffc_163_n_spl_,
    ffc_163_n
  );


  buf

  (
    ffc_162_n_spl_,
    ffc_162_n
  );


  buf

  (
    ffc_163_p_spl_,
    ffc_163_p
  );


  buf

  (
    ffc_163_p_spl_0,
    ffc_163_p_spl_
  );


  buf

  (
    ffc_164_p_spl_,
    ffc_164_p
  );


  buf

  (
    ffc_164_p_spl_0,
    ffc_164_p_spl_
  );


  buf

  (
    ffc_165_n_spl_,
    ffc_165_n
  );


  buf

  (
    ffc_164_n_spl_,
    ffc_164_n
  );


  buf

  (
    ffc_165_p_spl_,
    ffc_165_p
  );


  buf

  (
    ffc_165_p_spl_0,
    ffc_165_p_spl_
  );


  buf

  (
    ffc_166_p_spl_,
    ffc_166_p
  );


  buf

  (
    ffc_166_p_spl_0,
    ffc_166_p_spl_
  );


  buf

  (
    ffc_167_n_spl_,
    ffc_167_n
  );


  buf

  (
    ffc_166_n_spl_,
    ffc_166_n
  );


  buf

  (
    ffc_167_p_spl_,
    ffc_167_p
  );


  buf

  (
    ffc_167_p_spl_0,
    ffc_167_p_spl_
  );


  buf

  (
    ffc_168_p_spl_,
    ffc_168_p
  );


  buf

  (
    ffc_168_p_spl_0,
    ffc_168_p_spl_
  );


  buf

  (
    ffc_169_n_spl_,
    ffc_169_n
  );


  buf

  (
    ffc_168_n_spl_,
    ffc_168_n
  );


  buf

  (
    ffc_169_p_spl_,
    ffc_169_p
  );


  buf

  (
    ffc_169_p_spl_0,
    ffc_169_p_spl_
  );


  buf

  (
    ffc_170_p_spl_,
    ffc_170_p
  );


  buf

  (
    ffc_170_p_spl_0,
    ffc_170_p_spl_
  );


  buf

  (
    ffc_171_n_spl_,
    ffc_171_n
  );


  buf

  (
    ffc_170_n_spl_,
    ffc_170_n
  );


  buf

  (
    ffc_171_p_spl_,
    ffc_171_p
  );


  buf

  (
    ffc_171_p_spl_0,
    ffc_171_p_spl_
  );


  buf

  (
    ffc_172_p_spl_,
    ffc_172_p
  );


  buf

  (
    ffc_172_p_spl_0,
    ffc_172_p_spl_
  );


  buf

  (
    ffc_173_n_spl_,
    ffc_173_n
  );


  buf

  (
    ffc_172_n_spl_,
    ffc_172_n
  );


  buf

  (
    ffc_173_p_spl_,
    ffc_173_p
  );


  buf

  (
    ffc_173_p_spl_0,
    ffc_173_p_spl_
  );


  buf

  (
    ffc_174_p_spl_,
    ffc_174_p
  );


  buf

  (
    ffc_174_p_spl_0,
    ffc_174_p_spl_
  );


  buf

  (
    ffc_175_n_spl_,
    ffc_175_n
  );


  buf

  (
    ffc_174_n_spl_,
    ffc_174_n
  );


  buf

  (
    ffc_175_p_spl_,
    ffc_175_p
  );


  buf

  (
    ffc_175_p_spl_0,
    ffc_175_p_spl_
  );


  buf

  (
    ffc_176_p_spl_,
    ffc_176_p
  );


  buf

  (
    ffc_176_p_spl_0,
    ffc_176_p_spl_
  );


  buf

  (
    ffc_177_n_spl_,
    ffc_177_n
  );


  buf

  (
    ffc_176_n_spl_,
    ffc_176_n
  );


  buf

  (
    ffc_177_p_spl_,
    ffc_177_p
  );


  buf

  (
    ffc_177_p_spl_0,
    ffc_177_p_spl_
  );


  buf

  (
    ffc_178_p_spl_,
    ffc_178_p
  );


  buf

  (
    ffc_178_p_spl_0,
    ffc_178_p_spl_
  );


  buf

  (
    ffc_179_n_spl_,
    ffc_179_n
  );


  buf

  (
    ffc_178_n_spl_,
    ffc_178_n
  );


  buf

  (
    ffc_179_p_spl_,
    ffc_179_p
  );


  buf

  (
    ffc_179_p_spl_0,
    ffc_179_p_spl_
  );


  buf

  (
    ffc_180_p_spl_,
    ffc_180_p
  );


  buf

  (
    ffc_180_p_spl_0,
    ffc_180_p_spl_
  );


  buf

  (
    ffc_181_n_spl_,
    ffc_181_n
  );


  buf

  (
    ffc_180_n_spl_,
    ffc_180_n
  );


  buf

  (
    ffc_181_p_spl_,
    ffc_181_p
  );


  buf

  (
    ffc_181_p_spl_0,
    ffc_181_p_spl_
  );


  buf

  (
    ffc_182_p_spl_,
    ffc_182_p
  );


  buf

  (
    ffc_182_p_spl_0,
    ffc_182_p_spl_
  );


  buf

  (
    ffc_183_n_spl_,
    ffc_183_n
  );


  buf

  (
    ffc_182_n_spl_,
    ffc_182_n
  );


  buf

  (
    ffc_183_p_spl_,
    ffc_183_p
  );


  buf

  (
    ffc_183_p_spl_0,
    ffc_183_p_spl_
  );


  buf

  (
    ffc_184_p_spl_,
    ffc_184_p
  );


  buf

  (
    ffc_184_p_spl_0,
    ffc_184_p_spl_
  );


  buf

  (
    ffc_185_n_spl_,
    ffc_185_n
  );


  buf

  (
    ffc_184_n_spl_,
    ffc_184_n
  );


  buf

  (
    ffc_185_p_spl_,
    ffc_185_p
  );


  buf

  (
    ffc_185_p_spl_0,
    ffc_185_p_spl_
  );


  buf

  (
    ffc_186_p_spl_,
    ffc_186_p
  );


  buf

  (
    ffc_186_p_spl_0,
    ffc_186_p_spl_
  );


  buf

  (
    ffc_187_n_spl_,
    ffc_187_n
  );


  buf

  (
    ffc_186_n_spl_,
    ffc_186_n
  );


  buf

  (
    ffc_187_p_spl_,
    ffc_187_p
  );


  buf

  (
    ffc_187_p_spl_0,
    ffc_187_p_spl_
  );


  buf

  (
    ffc_188_p_spl_,
    ffc_188_p
  );


  buf

  (
    ffc_188_p_spl_0,
    ffc_188_p_spl_
  );


  buf

  (
    ffc_189_n_spl_,
    ffc_189_n
  );


  buf

  (
    ffc_188_n_spl_,
    ffc_188_n
  );


  buf

  (
    ffc_189_p_spl_,
    ffc_189_p
  );


  buf

  (
    ffc_189_p_spl_0,
    ffc_189_p_spl_
  );


  buf

  (
    ffc_190_p_spl_,
    ffc_190_p
  );


  buf

  (
    ffc_190_p_spl_0,
    ffc_190_p_spl_
  );


  buf

  (
    ffc_191_n_spl_,
    ffc_191_n
  );


  buf

  (
    ffc_190_n_spl_,
    ffc_190_n
  );


  buf

  (
    ffc_191_p_spl_,
    ffc_191_p
  );


  buf

  (
    ffc_191_p_spl_0,
    ffc_191_p_spl_
  );


  buf

  (
    ffc_192_p_spl_,
    ffc_192_p
  );


  buf

  (
    ffc_192_p_spl_0,
    ffc_192_p_spl_
  );


  buf

  (
    ffc_193_n_spl_,
    ffc_193_n
  );


  buf

  (
    ffc_192_n_spl_,
    ffc_192_n
  );


  buf

  (
    ffc_193_p_spl_,
    ffc_193_p
  );


  buf

  (
    ffc_193_p_spl_0,
    ffc_193_p_spl_
  );


endmodule
