// Benchmark "mymod" written by ABC on Wed Nov  1 23:37:39 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41,
    G468, G469, G470, G471, G472, G473, G474, G475, G476, G477, G478, G479,
    G480, G481, G482, G483, G484, G485, G486, G487, G488, G489, G490, G491,
    G492, G493, G494, G495, G496, G497, G498, G499  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41;
  output G468, G469, G470, G471, G472, G473, G474, G475, G476, G477, G478,
    G479, G480, G481, G482, G483, G484, G485, G486, G487, G488, G489, G490,
    G491, G492, G493, G494, G495, G496, G497, G498, G499;
  reg n286_lo, n298_lo, n310_lo, n322_lo, n334_lo, n346_lo, n358_lo,
    n370_lo, n382_lo, n394_lo, n406_lo, n418_lo, n430_lo, n442_lo, n454_lo,
    n466_lo, n478_lo, n490_lo, n502_lo, n514_lo, n526_lo, n538_lo, n550_lo,
    n562_lo, n574_lo, n586_lo, n598_lo, n610_lo, n622_lo, n634_lo, n646_lo,
    n658_lo, n661_lo, n673_lo, n685_lo, n697_lo, n709_lo, n721_lo, n733_lo,
    n745_lo, n757_lo, n1589_o2, n1590_o2, n1591_o2, n1592_o2, n1593_o2,
    n1594_o2, n1595_o2, n1596_o2, n1597_o2, n1598_o2, n1599_o2, n1600_o2,
    n1601_o2, n1602_o2, n1603_o2, n1604_o2, n1605_o2, n1606_o2, n1607_o2,
    n1608_o2, n1609_o2, n1610_o2, n1611_o2, n1612_o2, n1613_o2, n1614_o2,
    n1615_o2, n1616_o2, n1617_o2, n1618_o2, n1619_o2, n1620_o2, n602_o2,
    n639_o2, n678_o2, n658_o2, n783_o2, n802_o2, n726_o2, n763_o2, n685_o2,
    n680_o2, n822_o2, n843_o2, n842_o2, n681_o2, n684_o2, n686_o2, n823_o2,
    lo002_buf_o2, lo006_buf_o2, lo010_buf_o2, lo014_buf_o2, lo018_buf_o2,
    lo022_buf_o2, lo026_buf_o2, lo030_buf_o2, lo034_buf_o2, lo038_buf_o2,
    lo042_buf_o2, lo046_buf_o2, lo050_buf_o2, lo054_buf_o2, lo058_buf_o2,
    lo062_buf_o2, lo066_buf_o2, lo070_buf_o2, lo074_buf_o2, lo078_buf_o2,
    lo082_buf_o2, lo086_buf_o2, lo090_buf_o2, lo094_buf_o2, lo098_buf_o2,
    lo102_buf_o2, lo106_buf_o2, lo110_buf_o2, lo114_buf_o2, lo118_buf_o2,
    lo122_buf_o2, lo126_buf_o2, n683_o2, n688_o2, n803_o2, n862_o2,
    n764_o2, n863_o2, n886_o2, n600_o2, n601_o2, n637_o2, n638_o2, n676_o2,
    n677_o2, n656_o2, n657_o2, n781_o2, n782_o2, n800_o2, n801_o2, n724_o2,
    n725_o2, n761_o2, n762_o2, lo129_buf_o2, lo133_buf_o2, lo137_buf_o2,
    lo141_buf_o2, lo145_buf_o2, lo149_buf_o2, lo153_buf_o2, lo157_buf_o2,
    lo161_buf_o2, n708_o2, n745_o2, n717_o2, n754_o2, n584_o2, n593_o2,
    n630_o2, n621_o2, lo001_buf_o2, lo005_buf_o2, lo009_buf_o2,
    lo013_buf_o2, lo017_buf_o2, lo021_buf_o2, lo025_buf_o2, lo029_buf_o2,
    lo033_buf_o2, lo037_buf_o2, lo041_buf_o2, lo045_buf_o2, lo049_buf_o2,
    lo053_buf_o2, lo057_buf_o2, lo061_buf_o2, lo065_buf_o2, lo069_buf_o2,
    lo073_buf_o2, lo077_buf_o2, lo081_buf_o2, lo085_buf_o2, lo089_buf_o2,
    lo093_buf_o2, lo097_buf_o2, lo101_buf_o2, lo105_buf_o2, lo109_buf_o2,
    lo113_buf_o2, lo117_buf_o2, lo121_buf_o2, lo125_buf_o2;
  wire new_new_n462__, new_new_n464__, new_new_n466__, new_new_n468__,
    new_new_n470__, new_new_n472__, new_new_n474__, new_new_n476__,
    new_new_n478__, new_new_n480__, new_new_n482__, new_new_n484__,
    new_new_n486__, new_new_n488__, new_new_n490__, new_new_n492__,
    new_new_n494__, new_new_n496__, new_new_n498__, new_new_n500__,
    new_new_n502__, new_new_n504__, new_new_n506__, new_new_n508__,
    new_new_n510__, new_new_n512__, new_new_n514__, new_new_n516__,
    new_new_n518__, new_new_n520__, new_new_n522__, new_new_n524__,
    new_new_n526__, new_new_n528__, new_new_n530__, new_new_n532__,
    new_new_n534__, new_new_n536__, new_new_n538__, new_new_n540__,
    new_new_n542__, new_new_n544__, new_new_n545__, new_new_n546__,
    new_new_n547__, new_new_n548__, new_new_n549__, new_new_n550__,
    new_new_n551__, new_new_n552__, new_new_n553__, new_new_n554__,
    new_new_n555__, new_new_n556__, new_new_n557__, new_new_n558__,
    new_new_n559__, new_new_n560__, new_new_n561__, new_new_n562__,
    new_new_n563__, new_new_n564__, new_new_n565__, new_new_n566__,
    new_new_n567__, new_new_n568__, new_new_n569__, new_new_n570__,
    new_new_n571__, new_new_n572__, new_new_n573__, new_new_n574__,
    new_new_n575__, new_new_n576__, new_new_n577__, new_new_n578__,
    new_new_n579__, new_new_n580__, new_new_n581__, new_new_n582__,
    new_new_n583__, new_new_n584__, new_new_n585__, new_new_n586__,
    new_new_n587__, new_new_n588__, new_new_n589__, new_new_n590__,
    new_new_n591__, new_new_n592__, new_new_n593__, new_new_n594__,
    new_new_n595__, new_new_n596__, new_new_n597__, new_new_n598__,
    new_new_n599__, new_new_n600__, new_new_n601__, new_new_n602__,
    new_new_n603__, new_new_n604__, new_new_n605__, new_new_n606__,
    new_new_n607__, new_new_n608__, new_new_n610__, new_new_n612__,
    new_new_n614__, new_new_n616__, new_new_n618__, new_new_n620__,
    new_new_n622__, new_new_n624__, new_new_n626__, new_new_n628__,
    new_new_n630__, new_new_n632__, new_new_n634__, new_new_n636__,
    new_new_n638__, new_new_n640__, new_new_n642__, new_new_n644__,
    new_new_n646__, new_new_n648__, new_new_n650__, new_new_n652__,
    new_new_n654__, new_new_n656__, new_new_n658__, new_new_n660__,
    new_new_n662__, new_new_n664__, new_new_n666__, new_new_n668__,
    new_new_n670__, new_new_n672__, new_new_n674__, new_new_n676__,
    new_new_n678__, new_new_n680__, new_new_n682__, new_new_n684__,
    new_new_n686__, new_new_n688__, new_new_n690__, new_new_n691__,
    new_new_n692__, new_new_n693__, new_new_n694__, new_new_n695__,
    new_new_n696__, new_new_n697__, new_new_n698__, new_new_n699__,
    new_new_n700__, new_new_n701__, new_new_n702__, new_new_n703__,
    new_new_n704__, new_new_n705__, new_new_n706__, new_new_n707__,
    new_new_n708__, new_new_n709__, new_new_n710__, new_new_n711__,
    new_new_n712__, new_new_n713__, new_new_n714__, new_new_n715__,
    new_new_n716__, new_new_n717__, new_new_n718__, new_new_n719__,
    new_new_n720__, new_new_n721__, new_new_n722__, new_new_n723__,
    new_new_n724__, new_new_n725__, new_new_n726__, new_new_n727__,
    new_new_n728__, new_new_n729__, new_new_n730__, new_new_n731__,
    new_new_n732__, new_new_n733__, new_new_n734__, new_new_n735__,
    new_new_n736__, new_new_n737__, new_new_n738__, new_new_n739__,
    new_new_n740__, new_new_n741__, new_new_n742__, new_new_n743__,
    new_new_n744__, new_new_n745__, new_new_n746__, new_new_n747__,
    new_new_n748__, new_new_n749__, new_new_n750__, new_new_n751__,
    new_new_n752__, new_new_n753__, new_new_n754__, new_new_n755__,
    new_new_n756__, new_new_n757__, new_new_n758__, new_new_n759__,
    new_new_n760__, new_new_n761__, new_new_n762__, new_new_n763__,
    new_new_n764__, new_new_n765__, new_new_n766__, new_new_n767__,
    new_new_n768__, new_new_n769__, new_new_n770__, new_new_n771__,
    new_new_n772__, new_new_n773__, new_new_n774__, new_new_n775__,
    new_new_n776__, new_new_n777__, new_new_n778__, new_new_n779__,
    new_new_n780__, new_new_n781__, new_new_n782__, new_new_n783__,
    new_new_n784__, new_new_n785__, new_new_n786__, new_new_n787__,
    new_new_n788__, new_new_n789__, new_new_n790__, new_new_n791__,
    new_new_n792__, new_new_n793__, new_new_n794__, new_new_n795__,
    new_new_n796__, new_new_n797__, new_new_n798__, new_new_n799__,
    new_new_n800__, new_new_n801__, new_new_n802__, new_new_n803__,
    new_new_n804__, new_new_n805__, new_new_n806__, new_new_n807__,
    new_new_n808__, new_new_n809__, new_new_n810__, new_new_n811__,
    new_new_n812__, new_new_n813__, new_new_n814__, new_new_n815__,
    new_new_n816__, new_new_n817__, new_new_n818__, new_new_n819__,
    new_new_n820__, new_new_n821__, new_new_n822__, new_new_n823__,
    new_new_n824__, new_new_n825__, new_new_n826__, new_new_n827__,
    new_new_n828__, new_new_n829__, new_new_n830__, new_new_n831__,
    new_new_n832__, new_new_n833__, new_new_n834__, new_new_n835__,
    new_new_n836__, new_new_n837__, new_new_n838__, new_new_n839__,
    new_new_n840__, new_new_n841__, new_new_n842__, new_new_n843__,
    new_new_n844__, new_new_n845__, new_new_n846__, new_new_n847__,
    new_new_n848__, new_new_n849__, new_new_n850__, new_new_n851__,
    new_new_n852__, new_new_n853__, new_new_n854__, new_new_n855__,
    new_new_n856__, new_new_n857__, new_new_n858__, new_new_n859__,
    new_new_n860__, new_new_n861__, new_new_n862__, new_new_n863__,
    new_new_n864__, new_new_n865__, new_new_n866__, new_new_n867__,
    new_new_n868__, new_new_n869__, new_new_n870__, new_new_n871__,
    new_new_n872__, new_new_n873__, new_new_n874__, new_new_n875__,
    new_new_n876__, new_new_n877__, new_new_n878__, new_new_n879__,
    new_new_n880__, new_new_n881__, new_new_n882__, new_new_n883__,
    new_new_n884__, new_new_n885__, new_new_n886__, new_new_n887__,
    new_new_n888__, new_new_n889__, new_new_n890__, new_new_n891__,
    new_new_n892__, new_new_n893__, new_new_n894__, new_new_n895__,
    new_new_n896__, new_new_n897__, new_new_n898__, new_new_n899__,
    new_new_n900__, new_new_n901__, new_new_n902__, new_new_n903__,
    new_new_n904__, new_new_n905__, new_new_n906__, new_new_n907__,
    new_new_n908__, new_new_n909__, new_new_n910__, new_new_n911__,
    new_new_n912__, new_new_n913__, new_new_n914__, new_new_n915__,
    new_new_n916__, new_new_n917__, new_new_n918__, new_new_n919__,
    new_new_n920__, new_new_n921__, new_new_n922__, new_new_n923__,
    new_new_n924__, new_new_n925__, new_new_n926__, new_new_n927__,
    new_new_n928__, new_new_n929__, new_new_n930__, new_new_n931__,
    new_new_n932__, new_new_n933__, new_new_n934__, new_new_n935__,
    new_new_n936__, new_new_n937__, new_new_n938__, new_new_n939__,
    new_new_n940__, new_new_n941__, new_new_n942__, new_new_n943__,
    new_new_n944__, new_new_n945__, new_new_n946__, new_new_n947__,
    new_new_n948__, new_new_n949__, new_new_n950__, new_new_n951__,
    new_new_n952__, new_new_n953__, new_new_n954__, new_new_n955__,
    new_new_n956__, new_new_n957__, new_new_n958__, new_new_n959__,
    new_new_n960__, new_new_n961__, new_new_n962__, new_new_n963__,
    new_new_n964__, new_new_n965__, new_new_n966__, new_new_n967__,
    new_new_n968__, new_new_n969__, new_new_n970__, new_new_n971__,
    new_new_n972__, new_new_n973__, new_new_n974__, new_new_n975__,
    new_new_n976__, new_new_n977__, new_new_n978__, new_new_n979__,
    new_new_n980__, new_new_n981__, new_new_n982__, new_new_n983__,
    new_new_n984__, new_new_n985__, new_new_n986__, new_new_n987__,
    new_new_n988__, new_new_n989__, new_new_n990__, new_new_n991__,
    new_new_n992__, new_new_n993__, new_new_n994__, new_new_n995__,
    new_new_n996__, new_new_n997__, new_new_n998__, new_new_n999__,
    new_new_n1000__, new_new_n1001__, new_new_n1002__, new_new_n1003__,
    new_new_n1004__, new_new_n1005__, new_new_n1006__, new_new_n1007__,
    new_new_n1008__, new_new_n1009__, new_new_n1010__, new_new_n1011__,
    new_new_n1012__, new_new_n1013__, new_new_n1014__, new_new_n1015__,
    new_new_n1016__, new_new_n1017__, new_new_n1018__, new_new_n1019__,
    new_new_n1020__, new_new_n1021__, new_new_n1022__, new_new_n1023__,
    new_new_n1024__, new_new_n1025__, new_new_n1026__, new_new_n1027__,
    new_new_n1028__, new_new_n1029__, new_new_n1030__, new_new_n1031__,
    new_new_n1032__, new_new_n1033__, new_new_n1034__, new_new_n1035__,
    new_new_n1036__, new_new_n1037__, new_new_n1038__, new_new_n1039__,
    new_new_n1040__, new_new_n1041__, new_new_n1042__, new_new_n1043__,
    new_new_n1044__, new_new_n1045__, new_new_n1046__, new_new_n1047__,
    new_new_n1048__, new_new_n1049__, new_new_n1050__, new_new_n1051__,
    new_new_n1052__, new_new_n1053__, new_new_n1054__, new_new_n1055__,
    new_new_n1056__, new_new_n1057__, new_new_n1058__, new_new_n1059__,
    new_new_n1060__, new_new_n1061__, new_new_n1062__, new_new_n1063__,
    new_new_n1064__, new_new_n1065__, new_new_n1066__, new_new_n1067__,
    new_new_n1068__, new_new_n1069__, new_new_n1070__, new_new_n1071__,
    new_new_n1072__, new_new_n1073__, new_new_n1074__, new_new_n1075__,
    new_new_n1076__, new_new_n1077__, new_new_n1078__, new_new_n1079__,
    new_new_n1080__, new_new_n1081__, new_new_n1082__, new_new_n1083__,
    new_new_n1084__, new_new_n1085__, new_new_n1086__, new_new_n1087__,
    new_new_n1088__, new_new_n1089__, new_new_n1090__, new_new_n1091__,
    new_new_n1092__, new_new_n1093__, new_new_n1094__, new_new_n1095__,
    new_new_n1096__, new_new_n1097__, new_new_n1098__, new_new_n1099__,
    new_new_n1100__, new_new_n1101__, new_new_n1102__, new_new_n1103__,
    new_new_n1104__, new_new_n1105__, new_new_n1106__, new_new_n1107__,
    new_new_n1108__, new_new_n1109__, new_new_n1110__, new_new_n1111__,
    new_new_n1112__, new_new_n1113__, new_new_n1114__, new_new_n1115__,
    new_new_n1116__, new_new_n1117__, new_new_n1118__, new_new_n1119__,
    new_new_n1120__, new_new_n1121__, new_new_n1122__, new_new_n1123__,
    new_new_n1124__, new_new_n1125__, new_new_n1126__, new_new_n1127__,
    new_new_n1128__, new_new_n1129__, new_new_n1130__, new_new_n1131__,
    new_new_n1132__, new_new_n1133__, new_new_n1134__, new_new_n1135__,
    new_new_n1136__, new_new_n1137__, new_new_n1138__, new_new_n1139__,
    new_new_n1140__, new_new_n1141__, new_new_n1142__, new_new_n1143__,
    new_new_n1144__, new_new_n1145__, new_new_n1146__, new_new_n1147__,
    new_new_n1148__, new_new_n1149__, new_new_n1150__, new_new_n1151__,
    new_new_n1152__, new_new_n1153__, new_new_n1154__, new_new_n1155__,
    new_new_n1156__, new_new_n1157__, new_new_n1158__, new_new_n1159__,
    new_new_n1160__, new_new_n1161__, new_new_n1162__, new_new_n1163__,
    new_new_n1164__, new_new_n1165__, new_new_n1166__, new_new_n1167__,
    new_new_n1168__, new_new_n1169__, new_new_n1170__, new_new_n1171__,
    new_new_n1172__, new_new_n1173__, new_new_n1174__, new_new_n1175__,
    new_new_n1176__, new_new_n1177__, new_new_n1178__, new_new_n1179__,
    new_new_n1180__, new_new_n1181__, new_new_n1182__, new_new_n1183__,
    new_new_n1184__, new_new_n1185__, new_new_n1186__, new_new_n1187__,
    new_new_n1188__, new_new_n1189__, new_new_n1190__, new_new_n1191__,
    new_new_n1192__, new_new_n1193__, new_new_n1194__, new_new_n1195__,
    new_new_n1196__, new_new_n1197__, new_new_n1198__, new_new_n1199__,
    new_new_n1200__, new_new_n1201__, new_new_n1202__, new_new_n1203__,
    new_new_n1204__, new_new_n1205__, new_new_n1206__, new_new_n1207__,
    new_new_n1208__, new_new_n1209__, new_new_n1210__, new_new_n1211__,
    new_new_n1212__, new_new_n1213__, new_new_n1214__, new_new_n1215__,
    new_new_n1216__, new_new_n1217__, new_new_n1218__, new_new_n1219__,
    new_new_n1220__, new_new_n1221__, new_new_n1222__, new_new_n1223__,
    new_new_n1224__, new_new_n1225__, new_new_n1226__, new_new_n1227__,
    new_new_n1228__, new_new_n1229__, new_new_n1230__, new_new_n1231__,
    new_new_n1232__, new_new_n1233__, new_new_n1234__, new_new_n1235__,
    new_new_n1236__, new_new_n1237__, new_new_n1238__, new_new_n1239__,
    new_new_n1240__, new_new_n1241__, new_new_n1242__, new_new_n1243__,
    new_new_n1244__, new_new_n1245__, new_new_n1246__, new_new_n1247__,
    new_new_n1248__, new_new_n1249__, new_new_n1250__, new_new_n1251__,
    new_new_n1252__, new_new_n1253__, new_new_n1254__, new_new_n1255__,
    new_new_n1256__, new_new_n1257__, new_new_n1258__, new_new_n1259__,
    new_new_n1260__, new_new_n1261__, new_new_n1262__, new_new_n1263__,
    new_new_n1264__, new_new_n1265__, new_new_n1266__, new_new_n1267__,
    new_new_n1268__, new_new_n1269__, new_new_n1270__, new_new_n1271__,
    new_new_n1272__, new_new_n1273__, new_new_n1274__, new_new_n1275__,
    new_new_n1276__, new_new_n1277__, new_new_n1278__, new_new_n1279__,
    new_new_n1280__, new_new_n1281__, new_new_n1282__, new_new_n1283__,
    new_new_n1284__, new_new_n1285__, new_new_n1286__, new_new_n1287__,
    new_new_n1288__, new_new_n1289__, new_new_n1290__, new_new_n1291__,
    new_new_n1292__, new_new_n1293__, new_new_n1294__, new_new_n1295__,
    new_new_n1296__, new_new_n1297__, new_new_n1298__, new_new_n1299__,
    new_new_n1300__, new_new_n1301__, new_new_n1302__, new_new_n1303__,
    new_new_n1304__, new_new_n1305__, new_new_n1306__, new_new_n1307__,
    new_new_n1308__, new_new_n1309__, new_new_n1310__, new_new_n1311__,
    new_new_n1312__, new_new_n1313__, new_new_n1314__, new_new_n1315__,
    new_new_n1316__, new_new_n1317__, new_new_n1318__, new_new_n1319__,
    new_new_n1320__, new_new_n1321__, new_new_n1322__, new_new_n1323__,
    new_new_n1324__, new_new_n1325__, new_new_n1326__, new_new_n1327__,
    new_new_n1328__, new_new_n1329__, new_new_n1330__, new_new_n1331__,
    new_new_n1332__, new_new_n1333__, new_new_n1334__, new_new_n1335__,
    new_new_n1336__, new_new_n1337__, new_new_n1338__, new_new_n1339__,
    new_new_n1340__, new_new_n1341__, new_new_n1342__, new_new_n1343__,
    new_new_n1344__, new_new_n1345__, new_new_n1346__, new_new_n1347__,
    new_new_n1348__, new_new_n1349__, new_new_n1350__, new_new_n1351__,
    new_new_n1352__, new_new_n1353__, new_new_n1354__, new_new_n1355__,
    new_new_n1356__, new_new_n1357__, new_new_n1358__, new_new_n1359__,
    new_new_n1360__, new_new_n1361__, new_new_n1362__, new_new_n1363__,
    new_new_n1364__, new_new_n1365__, new_new_n1366__, new_new_n1367__,
    new_new_n1368__, new_new_n1369__, new_new_n1370__, new_new_n1371__,
    new_new_n1372__, new_new_n1373__, new_new_n1374__, new_new_n1375__,
    new_new_n1376__, new_new_n1377__, new_new_n1378__, new_new_n1379__,
    new_new_n1380__, new_new_n1381__, new_new_n1382__, new_new_n1383__,
    new_new_n1384__, new_new_n1385__, new_new_n1386__, new_new_n1387__,
    new_new_n1388__, new_new_n1389__, new_new_n1390__, new_new_n1391__,
    new_new_n1392__, new_new_n1393__, new_new_n1394__, new_new_n1395__,
    new_new_n1396__, new_new_n1397__, new_new_n1398__, new_new_n1399__,
    new_new_n1400__, new_new_n1401__, new_new_n1402__, new_new_n1403__,
    new_new_n1404__, new_new_n1405__, new_new_n1406__, new_new_n1407__,
    new_new_n1408__, new_new_n1409__, new_new_n1410__, new_new_n1411__,
    new_new_n1412__, new_new_n1413__, new_new_n1414__, new_new_n1415__,
    new_new_n1416__, new_new_n1417__, new_new_n1418__, new_new_n1419__,
    new_new_n1420__, new_new_n1421__, new_new_n1422__, new_new_n1423__,
    new_new_n1424__, new_new_n1425__, new_new_n1426__, new_new_n1427__,
    new_new_n1428__, new_new_n1429__, new_new_n1430__, new_new_n1431__,
    new_new_n1432__, new_new_n1433__, new_new_n1434__, new_new_n1435__,
    new_new_n1436__, new_new_n1437__, new_new_n1438__, new_new_n1439__,
    new_new_n1440__, new_new_n1441__, new_new_n1442__, new_new_n1443__,
    new_new_n1444__, new_new_n1445__, new_new_n1446__, new_new_n1447__,
    new_new_n1448__, new_new_n1449__, new_new_n1450__, new_new_n1451__,
    new_new_n1452__, new_new_n1453__, new_new_n1454__, new_new_n1455__,
    new_new_n1456__, new_new_n1457__, new_new_n1458__, new_new_n1459__,
    new_new_n1460__, new_new_n1461__, new_new_n1462__, new_new_n1463__,
    new_new_n1464__, new_new_n1465__, new_new_n1466__, new_new_n1467__,
    new_new_n1468__, new_new_n1469__, new_new_n1470__, new_new_n1471__,
    new_new_n1472__, new_new_n1473__, new_new_n1474__, new_new_n1475__,
    new_new_n1476__, new_new_n1477__, new_new_n1478__, new_new_n1479__,
    new_new_n1480__, new_new_n1481__, new_new_n1482__, new_new_n1483__,
    new_new_n1484__, new_new_n1485__, new_new_n1486__, new_new_n1487__,
    new_new_n1488__, new_new_n1489__, new_new_n1490__, new_new_n1491__,
    new_new_n1492__, new_new_n1493__, new_new_n1494__, new_new_n1495__,
    new_new_n1496__, new_new_n1497__, new_new_n1498__, new_new_n1499__,
    new_new_n1500__, new_new_n1501__, new_new_n1502__, new_new_n1503__,
    new_new_n1504__, new_new_n1505__, new_new_n1506__, new_new_n1507__,
    new_new_n1508__, new_new_n1509__, new_new_n1510__, new_new_n1511__,
    new_new_n1738__, new_new_n1739__, new_new_n1740__, new_new_n1741__,
    new_new_n1742__, new_new_n1743__, new_new_n1744__, new_new_n1745__,
    new_new_n1746__, new_new_n1747__, new_new_n1748__, new_new_n1749__,
    new_new_n1750__, new_new_n1751__, new_new_n1752__, new_new_n1753__,
    new_new_n1754__, new_new_n1755__, new_new_n1756__, new_new_n1757__,
    new_new_n1758__, new_new_n1759__, new_new_n1760__, new_new_n1761__,
    new_new_n1762__, new_new_n1763__, new_new_n1764__, new_new_n1765__,
    new_new_n1766__, new_new_n1767__, new_new_n1768__, new_new_n1769__,
    new_new_n1770__, new_new_n1771__, new_new_n1772__, new_new_n1773__,
    new_new_n1774__, new_new_n1775__, new_new_n1776__, new_new_n1777__,
    new_new_n1778__, new_new_n1779__, new_new_n1780__, new_new_n1781__,
    new_new_n1782__, new_new_n1783__, new_new_n1784__, new_new_n1785__,
    new_new_n1786__, new_new_n1787__, new_new_n1788__, new_new_n1789__,
    new_new_n1790__, new_new_n1791__, new_new_n1792__, new_new_n1793__,
    new_new_n1794__, new_new_n1795__, new_new_n1796__, new_new_n1797__,
    new_new_n1798__, new_new_n1799__, new_new_n1800__, new_new_n1801__,
    new_new_n1802__, new_new_n1803__, new_new_n1804__, new_new_n1805__,
    new_new_n1806__, new_new_n1807__, new_new_n1808__, new_new_n1809__,
    new_new_n1810__, new_new_n1811__, new_new_n1812__, new_new_n1813__,
    new_new_n1814__, new_new_n1815__, new_new_n1816__, new_new_n1817__,
    new_new_n1818__, new_new_n1819__, new_new_n1820__, new_new_n1821__,
    new_new_n1822__, new_new_n1823__, new_new_n1824__, new_new_n1825__,
    new_new_n1826__, new_new_n1827__, new_new_n1828__, new_new_n1829__,
    new_new_n1830__, new_new_n1831__, new_new_n1832__, new_new_n1833__,
    new_new_n1834__, new_new_n1835__, new_new_n1836__, new_new_n1837__,
    new_new_n1838__, new_new_n1839__, new_new_n1840__, new_new_n1841__,
    new_new_n1842__, new_new_n1843__, new_new_n1844__, new_new_n1845__,
    new_new_n1846__, new_new_n1847__, new_new_n1848__, new_new_n1849__,
    new_new_n1850__, new_new_n1851__, new_new_n1852__, new_new_n1853__,
    new_new_n1854__, new_new_n1855__, new_new_n1856__, new_new_n1857__,
    new_new_n1858__, new_new_n1859__, new_new_n1860__, new_new_n1861__,
    new_new_n1862__, new_new_n1863__, new_new_n1864__, new_new_n1865__,
    new_new_n1866__, new_new_n1867__, new_new_n1868__, new_new_n1869__,
    new_new_n1870__, new_new_n1871__, new_new_n1872__, new_new_n1873__,
    new_new_n1874__, new_new_n1875__, new_new_n1876__, new_new_n1877__,
    new_new_n1878__, new_new_n1879__, new_new_n1880__, new_new_n1881__,
    new_new_n1882__, new_new_n1883__, new_new_n1884__, new_new_n1885__,
    new_new_n1886__, new_new_n1887__, new_new_n1888__, new_new_n1889__,
    new_new_n1890__, new_new_n1891__, new_new_n1892__, new_new_n1893__,
    new_new_n1894__, new_new_n1895__, new_new_n1896__, new_new_n1897__,
    new_new_n1898__, new_new_n1899__, new_new_n1900__, new_new_n1901__,
    new_new_n1902__, new_new_n1903__, new_new_n1904__, new_new_n1905__,
    new_new_n1906__, new_new_n1907__, new_new_n1908__, new_new_n1909__,
    new_new_n1910__, new_new_n1911__, new_new_n1912__, new_new_n1913__,
    new_new_n1914__, new_new_n1915__, new_new_n1916__, new_new_n1917__,
    new_new_n1918__, new_new_n1919__, new_new_n1920__, new_new_n1921__,
    new_new_n1922__, new_new_n1923__, new_new_n1924__, new_new_n1925__,
    new_new_n1926__, new_new_n1927__, new_new_n1928__, new_new_n1929__,
    new_new_n1930__, new_new_n1931__, new_new_n1932__, new_new_n1933__,
    new_new_n1934__, new_new_n1935__, new_new_n1936__, new_new_n1937__,
    new_new_n1938__, new_new_n1939__, new_new_n1940__, new_new_n1941__,
    new_new_n1942__, new_new_n1943__, new_new_n1944__, new_new_n1945__,
    new_new_n1946__, new_new_n1947__, new_new_n1948__, new_new_n1949__,
    new_new_n1950__, new_new_n1951__, new_new_n1952__, new_new_n1953__,
    new_new_n1954__, new_new_n1955__, new_new_n1956__, new_new_n1957__,
    new_new_n1958__, new_new_n1959__, new_new_n1960__, new_new_n1961__,
    new_new_n1962__, new_new_n1963__, new_new_n1964__, new_new_n1965__,
    new_new_n1966__, new_new_n1967__, new_new_n1968__, new_new_n1969__,
    new_new_n1970__, new_new_n1971__, new_new_n1972__, new_new_n1973__,
    new_new_n1974__, new_new_n1975__, new_new_n1976__, new_new_n1977__,
    new_new_n1978__, new_new_n1979__, new_new_n1980__, new_new_n1981__,
    new_new_n1982__, new_new_n1983__, new_new_n1984__, new_new_n1985__,
    new_new_n1986__, new_new_n1987__, new_new_n1988__, new_new_n1989__,
    new_new_n1990__, new_new_n1991__, new_new_n1992__, new_new_n1993__,
    new_new_n1994__, new_new_n1995__, new_new_n1996__, new_new_n1997__,
    new_new_n1998__, new_new_n1999__, new_new_n2000__, new_new_n2001__,
    new_new_n2002__, new_new_n2003__, new_new_n2004__, new_new_n2005__,
    new_new_n2006__, new_new_n2007__, new_new_n2008__, new_new_n2009__,
    new_new_n2010__, new_new_n2011__, new_new_n2012__, new_new_n2013__,
    new_new_n2014__, new_new_n2015__, new_new_n2016__, new_new_n2017__,
    new_new_n2018__, new_new_n2019__, new_new_n2020__, new_new_n2021__,
    new_new_n2022__, new_new_n2023__, new_new_n2024__, new_new_n2025__,
    new_new_n2026__, new_new_n2027__, new_new_n2028__, new_new_n2029__,
    new_new_n2030__, new_new_n2031__, new_new_n2032__, new_new_n2033__,
    new_new_n2034__, new_new_n2035__, new_new_n2036__, new_new_n2037__,
    new_new_n2038__, new_new_n2039__, new_new_n2040__, new_new_n2041__,
    new_new_n2042__, new_new_n2043__, new_new_n2044__, new_new_n2045__,
    new_new_n2046__, new_new_n2047__, new_new_n2048__, new_new_n2049__,
    new_new_n2050__, new_new_n2051__, new_new_n2052__, new_new_n2053__,
    new_new_n2054__, new_new_n2055__, new_new_n2056__, new_new_n2057__,
    new_new_n2058__, new_new_n2059__, new_new_n2060__, new_new_n2061__,
    new_new_n2062__, new_new_n2063__, new_new_n2064__, new_new_n2065__,
    new_new_n2066__, new_new_n2067__, new_new_n2068__, new_new_n2069__,
    new_new_n2070__, new_new_n2071__, new_new_n2072__, new_new_n2073__,
    new_new_n2074__, new_new_n2075__, new_new_n2076__, new_new_n2077__,
    new_new_n2078__, new_new_n2079__, new_new_n2080__, new_new_n2081__,
    new_new_n2082__, new_new_n2083__, new_new_n2084__, new_new_n2085__,
    new_new_n2086__, new_new_n2087__, new_new_n2088__, new_new_n2089__,
    new_new_n2090__, new_new_n2091__, new_new_n2092__, new_new_n2093__,
    new_new_n2094__, new_new_n2095__, new_new_n2096__, new_new_n2097__,
    new_new_n2098__, new_new_n2099__, new_new_n2100__, new_new_n2101__,
    new_new_n2102__, new_new_n2103__, new_new_n2104__, new_new_n2105__,
    new_new_n2106__, new_new_n2107__, new_new_n2108__, new_new_n2109__,
    new_new_n2110__, new_new_n2111__, new_new_n2112__, new_new_n2113__,
    new_new_n2114__, new_new_n2115__, new_new_n2116__, new_new_n2117__,
    new_new_n2118__, new_new_n2119__, new_new_n2120__, new_new_n2121__,
    new_new_n2122__, new_new_n2123__, new_new_n2124__, new_new_n2125__,
    new_new_n2126__, new_new_n2127__, new_new_n2128__, new_new_n2129__,
    new_new_n2130__, new_new_n2131__, new_new_n2132__, new_new_n2133__,
    new_new_n2134__, new_new_n2135__, new_new_n2136__, new_new_n2137__,
    new_new_n2138__, new_new_n2139__, new_new_n2140__, new_new_n2141__,
    new_new_n2142__, new_new_n2143__, new_new_n2144__, new_new_n2145__,
    new_new_n2146__, new_new_n2147__, new_new_n2148__, new_new_n2149__,
    new_new_n2150__, new_new_n2151__, new_new_n2152__, new_new_n2153__,
    new_new_n2154__, new_new_n2155__, n3533, n3536, n3539, n3542, n3545,
    n3548, n3551, n3554, n3557, n3560, n3563, n3566, n3569, n3572, n3575,
    n3578, n3581, n3584, n3587, n3590, n3593, n3596, n3599, n3602, n3605,
    n3608, n3611, n3614, n3617, n3620, n3623, n3626, n3629, n3632, n3635,
    n3638, n3641, n3644, n3647, n3650, n3653, n3656, n3659, n3662, n3665,
    n3668, n3671, n3674, n3677, n3680, n3683, n3686, n3689, n3692, n3695,
    n3698, n3701, n3704, n3707, n3710, n3713, n3716, n3719, n3722, n3725,
    n3728, n3731, n3734, n3737, n3740, n3743, n3746, n3749, n3752, n3755,
    n3758, n3761, n3764, n3767, n3770, n3773, n3776, n3779, n3782, n3785,
    n3788, n3791, n3794, n3797, n3800, n3803, n3806, n3809, n3812, n3815,
    n3818, n3821, n3824, n3827, n3830, n3833, n3836, n3839, n3842, n3845,
    n3848, n3851, n3854, n3857, n3860, n3863, n3866, n3869, n3872, n3875,
    n3878, n3881, n3884, n3887, n3890, n3893, n3896, n3899, n3902, n3905,
    n3908, n3911, n3914, n3917, n3920, n3923, n3926, n3929, n3932, n3935,
    n3938, n3941, n3944, n3947, n3950, n3953, n3956, n3959, n3962, n3965,
    n3968, n3971, n3974, n3977, n3980, n3983, n3986, n3989, n3992, n3995,
    n3998, n4001, n4004, n4007, n4010, n4013, n4016, n4019, n4022, n4025,
    n4028, n4031, n4034, n4037, n4040, n4043, n4046, n4049, n4052, n4055,
    n4058, n4061, n4064, n4067, n4070, n4073, n4076, n4079, n4082, n4085,
    n4088, n4091, n4094, n4097, n4100, n4103, n4106, n4109, n4112;
  buf1  g0000(.din(G1), .dout(new_new_n462__));
  buf1  g0001(.din(G2), .dout(new_new_n464__));
  buf1  g0002(.din(G3), .dout(new_new_n466__));
  buf1  g0003(.din(G4), .dout(new_new_n468__));
  buf1  g0004(.din(G5), .dout(new_new_n470__));
  buf1  g0005(.din(G6), .dout(new_new_n472__));
  buf1  g0006(.din(G7), .dout(new_new_n474__));
  buf1  g0007(.din(G8), .dout(new_new_n476__));
  buf1  g0008(.din(G9), .dout(new_new_n478__));
  buf1  g0009(.din(G10), .dout(new_new_n480__));
  buf1  g0010(.din(G11), .dout(new_new_n482__));
  buf1  g0011(.din(G12), .dout(new_new_n484__));
  buf1  g0012(.din(G13), .dout(new_new_n486__));
  buf1  g0013(.din(G14), .dout(new_new_n488__));
  buf1  g0014(.din(G15), .dout(new_new_n490__));
  buf1  g0015(.din(G16), .dout(new_new_n492__));
  buf1  g0016(.din(G17), .dout(new_new_n494__));
  buf1  g0017(.din(G18), .dout(new_new_n496__));
  buf1  g0018(.din(G19), .dout(new_new_n498__));
  buf1  g0019(.din(G20), .dout(new_new_n500__));
  buf1  g0020(.din(G21), .dout(new_new_n502__));
  buf1  g0021(.din(G22), .dout(new_new_n504__));
  buf1  g0022(.din(G23), .dout(new_new_n506__));
  buf1  g0023(.din(G24), .dout(new_new_n508__));
  buf1  g0024(.din(G25), .dout(new_new_n510__));
  buf1  g0025(.din(G26), .dout(new_new_n512__));
  buf1  g0026(.din(G27), .dout(new_new_n514__));
  buf1  g0027(.din(G28), .dout(new_new_n516__));
  buf1  g0028(.din(G29), .dout(new_new_n518__));
  buf1  g0029(.din(G30), .dout(new_new_n520__));
  buf1  g0030(.din(G31), .dout(new_new_n522__));
  buf1  g0031(.din(G32), .dout(new_new_n524__));
  buf1  g0032(.din(G33), .dout(new_new_n526__));
  buf1  g0033(.din(G34), .dout(new_new_n528__));
  buf1  g0034(.din(G35), .dout(new_new_n530__));
  buf1  g0035(.din(G36), .dout(new_new_n532__));
  buf1  g0036(.din(G37), .dout(new_new_n534__));
  buf1  g0037(.din(G38), .dout(new_new_n536__));
  buf1  g0038(.din(G39), .dout(new_new_n538__));
  buf1  g0039(.din(G40), .dout(new_new_n540__));
  buf1  g0040(.din(G41), .dout(new_new_n542__));
  buf1  g0041(.din(n286_lo), .dout(new_new_n544__));
  not1  g0042(.din(n286_lo), .dout(new_new_n545__));
  buf1  g0043(.din(n298_lo), .dout(new_new_n546__));
  not1  g0044(.din(n298_lo), .dout(new_new_n547__));
  buf1  g0045(.din(n310_lo), .dout(new_new_n548__));
  not1  g0046(.din(n310_lo), .dout(new_new_n549__));
  buf1  g0047(.din(n322_lo), .dout(new_new_n550__));
  not1  g0048(.din(n322_lo), .dout(new_new_n551__));
  buf1  g0049(.din(n334_lo), .dout(new_new_n552__));
  not1  g0050(.din(n334_lo), .dout(new_new_n553__));
  buf1  g0051(.din(n346_lo), .dout(new_new_n554__));
  not1  g0052(.din(n346_lo), .dout(new_new_n555__));
  buf1  g0053(.din(n358_lo), .dout(new_new_n556__));
  not1  g0054(.din(n358_lo), .dout(new_new_n557__));
  buf1  g0055(.din(n370_lo), .dout(new_new_n558__));
  not1  g0056(.din(n370_lo), .dout(new_new_n559__));
  buf1  g0057(.din(n382_lo), .dout(new_new_n560__));
  not1  g0058(.din(n382_lo), .dout(new_new_n561__));
  buf1  g0059(.din(n394_lo), .dout(new_new_n562__));
  not1  g0060(.din(n394_lo), .dout(new_new_n563__));
  buf1  g0061(.din(n406_lo), .dout(new_new_n564__));
  not1  g0062(.din(n406_lo), .dout(new_new_n565__));
  buf1  g0063(.din(n418_lo), .dout(new_new_n566__));
  not1  g0064(.din(n418_lo), .dout(new_new_n567__));
  buf1  g0065(.din(n430_lo), .dout(new_new_n568__));
  not1  g0066(.din(n430_lo), .dout(new_new_n569__));
  buf1  g0067(.din(n442_lo), .dout(new_new_n570__));
  not1  g0068(.din(n442_lo), .dout(new_new_n571__));
  buf1  g0069(.din(n454_lo), .dout(new_new_n572__));
  not1  g0070(.din(n454_lo), .dout(new_new_n573__));
  buf1  g0071(.din(n466_lo), .dout(new_new_n574__));
  not1  g0072(.din(n466_lo), .dout(new_new_n575__));
  buf1  g0073(.din(n478_lo), .dout(new_new_n576__));
  not1  g0074(.din(n478_lo), .dout(new_new_n577__));
  buf1  g0075(.din(n490_lo), .dout(new_new_n578__));
  not1  g0076(.din(n490_lo), .dout(new_new_n579__));
  buf1  g0077(.din(n502_lo), .dout(new_new_n580__));
  not1  g0078(.din(n502_lo), .dout(new_new_n581__));
  buf1  g0079(.din(n514_lo), .dout(new_new_n582__));
  not1  g0080(.din(n514_lo), .dout(new_new_n583__));
  buf1  g0081(.din(n526_lo), .dout(new_new_n584__));
  not1  g0082(.din(n526_lo), .dout(new_new_n585__));
  buf1  g0083(.din(n538_lo), .dout(new_new_n586__));
  not1  g0084(.din(n538_lo), .dout(new_new_n587__));
  buf1  g0085(.din(n550_lo), .dout(new_new_n588__));
  not1  g0086(.din(n550_lo), .dout(new_new_n589__));
  buf1  g0087(.din(n562_lo), .dout(new_new_n590__));
  not1  g0088(.din(n562_lo), .dout(new_new_n591__));
  buf1  g0089(.din(n574_lo), .dout(new_new_n592__));
  not1  g0090(.din(n574_lo), .dout(new_new_n593__));
  buf1  g0091(.din(n586_lo), .dout(new_new_n594__));
  not1  g0092(.din(n586_lo), .dout(new_new_n595__));
  buf1  g0093(.din(n598_lo), .dout(new_new_n596__));
  not1  g0094(.din(n598_lo), .dout(new_new_n597__));
  buf1  g0095(.din(n610_lo), .dout(new_new_n598__));
  not1  g0096(.din(n610_lo), .dout(new_new_n599__));
  buf1  g0097(.din(n622_lo), .dout(new_new_n600__));
  not1  g0098(.din(n622_lo), .dout(new_new_n601__));
  buf1  g0099(.din(n634_lo), .dout(new_new_n602__));
  not1  g0100(.din(n634_lo), .dout(new_new_n603__));
  buf1  g0101(.din(n646_lo), .dout(new_new_n604__));
  not1  g0102(.din(n646_lo), .dout(new_new_n605__));
  buf1  g0103(.din(n658_lo), .dout(new_new_n606__));
  not1  g0104(.din(n658_lo), .dout(new_new_n607__));
  buf1  g0105(.din(n661_lo), .dout(new_new_n608__));
  buf1  g0106(.din(n673_lo), .dout(new_new_n610__));
  buf1  g0107(.din(n685_lo), .dout(new_new_n612__));
  buf1  g0108(.din(n697_lo), .dout(new_new_n614__));
  buf1  g0109(.din(n709_lo), .dout(new_new_n616__));
  buf1  g0110(.din(n721_lo), .dout(new_new_n618__));
  buf1  g0111(.din(n733_lo), .dout(new_new_n620__));
  buf1  g0112(.din(n745_lo), .dout(new_new_n622__));
  buf1  g0113(.din(n757_lo), .dout(new_new_n624__));
  buf1  g0114(.din(n1589_o2), .dout(new_new_n626__));
  buf1  g0115(.din(n1590_o2), .dout(new_new_n628__));
  buf1  g0116(.din(n1591_o2), .dout(new_new_n630__));
  buf1  g0117(.din(n1592_o2), .dout(new_new_n632__));
  buf1  g0118(.din(n1593_o2), .dout(new_new_n634__));
  buf1  g0119(.din(n1594_o2), .dout(new_new_n636__));
  buf1  g0120(.din(n1595_o2), .dout(new_new_n638__));
  buf1  g0121(.din(n1596_o2), .dout(new_new_n640__));
  buf1  g0122(.din(n1597_o2), .dout(new_new_n642__));
  buf1  g0123(.din(n1598_o2), .dout(new_new_n644__));
  buf1  g0124(.din(n1599_o2), .dout(new_new_n646__));
  buf1  g0125(.din(n1600_o2), .dout(new_new_n648__));
  buf1  g0126(.din(n1601_o2), .dout(new_new_n650__));
  buf1  g0127(.din(n1602_o2), .dout(new_new_n652__));
  buf1  g0128(.din(n1603_o2), .dout(new_new_n654__));
  buf1  g0129(.din(n1604_o2), .dout(new_new_n656__));
  buf1  g0130(.din(n1605_o2), .dout(new_new_n658__));
  buf1  g0131(.din(n1606_o2), .dout(new_new_n660__));
  buf1  g0132(.din(n1607_o2), .dout(new_new_n662__));
  buf1  g0133(.din(n1608_o2), .dout(new_new_n664__));
  buf1  g0134(.din(n1609_o2), .dout(new_new_n666__));
  buf1  g0135(.din(n1610_o2), .dout(new_new_n668__));
  buf1  g0136(.din(n1611_o2), .dout(new_new_n670__));
  buf1  g0137(.din(n1612_o2), .dout(new_new_n672__));
  buf1  g0138(.din(n1613_o2), .dout(new_new_n674__));
  buf1  g0139(.din(n1614_o2), .dout(new_new_n676__));
  buf1  g0140(.din(n1615_o2), .dout(new_new_n678__));
  buf1  g0141(.din(n1616_o2), .dout(new_new_n680__));
  buf1  g0142(.din(n1617_o2), .dout(new_new_n682__));
  buf1  g0143(.din(n1618_o2), .dout(new_new_n684__));
  buf1  g0144(.din(n1619_o2), .dout(new_new_n686__));
  buf1  g0145(.din(n1620_o2), .dout(new_new_n688__));
  buf1  g0146(.din(n602_o2), .dout(new_new_n690__));
  not1  g0147(.din(n602_o2), .dout(new_new_n691__));
  buf1  g0148(.din(n639_o2), .dout(new_new_n692__));
  not1  g0149(.din(n639_o2), .dout(new_new_n693__));
  buf1  g0150(.din(n678_o2), .dout(new_new_n694__));
  not1  g0151(.din(n678_o2), .dout(new_new_n695__));
  buf1  g0152(.din(n658_o2), .dout(new_new_n696__));
  not1  g0153(.din(n658_o2), .dout(new_new_n697__));
  buf1  g0154(.din(n783_o2), .dout(new_new_n698__));
  not1  g0155(.din(n783_o2), .dout(new_new_n699__));
  buf1  g0156(.din(n802_o2), .dout(new_new_n700__));
  not1  g0157(.din(n802_o2), .dout(new_new_n701__));
  buf1  g0158(.din(n726_o2), .dout(new_new_n702__));
  not1  g0159(.din(n726_o2), .dout(new_new_n703__));
  buf1  g0160(.din(n763_o2), .dout(new_new_n704__));
  not1  g0161(.din(n763_o2), .dout(new_new_n705__));
  buf1  g0162(.din(n685_o2), .dout(new_new_n706__));
  not1  g0163(.din(n685_o2), .dout(new_new_n707__));
  buf1  g0164(.din(n680_o2), .dout(new_new_n708__));
  not1  g0165(.din(n680_o2), .dout(new_new_n709__));
  buf1  g0166(.din(n822_o2), .dout(new_new_n710__));
  not1  g0167(.din(n822_o2), .dout(new_new_n711__));
  buf1  g0168(.din(n843_o2), .dout(new_new_n712__));
  not1  g0169(.din(n843_o2), .dout(new_new_n713__));
  buf1  g0170(.din(n842_o2), .dout(new_new_n714__));
  not1  g0171(.din(n842_o2), .dout(new_new_n715__));
  buf1  g0172(.din(n681_o2), .dout(new_new_n716__));
  not1  g0173(.din(n681_o2), .dout(new_new_n717__));
  buf1  g0174(.din(n684_o2), .dout(new_new_n718__));
  not1  g0175(.din(n684_o2), .dout(new_new_n719__));
  buf1  g0176(.din(n686_o2), .dout(new_new_n720__));
  not1  g0177(.din(n686_o2), .dout(new_new_n721__));
  buf1  g0178(.din(n823_o2), .dout(new_new_n722__));
  not1  g0179(.din(n823_o2), .dout(new_new_n723__));
  buf1  g0180(.din(lo002_buf_o2), .dout(new_new_n724__));
  not1  g0181(.din(lo002_buf_o2), .dout(new_new_n725__));
  buf1  g0182(.din(lo006_buf_o2), .dout(new_new_n726__));
  not1  g0183(.din(lo006_buf_o2), .dout(new_new_n727__));
  buf1  g0184(.din(lo010_buf_o2), .dout(new_new_n728__));
  not1  g0185(.din(lo010_buf_o2), .dout(new_new_n729__));
  buf1  g0186(.din(lo014_buf_o2), .dout(new_new_n730__));
  not1  g0187(.din(lo014_buf_o2), .dout(new_new_n731__));
  buf1  g0188(.din(lo018_buf_o2), .dout(new_new_n732__));
  not1  g0189(.din(lo018_buf_o2), .dout(new_new_n733__));
  buf1  g0190(.din(lo022_buf_o2), .dout(new_new_n734__));
  not1  g0191(.din(lo022_buf_o2), .dout(new_new_n735__));
  buf1  g0192(.din(lo026_buf_o2), .dout(new_new_n736__));
  not1  g0193(.din(lo026_buf_o2), .dout(new_new_n737__));
  buf1  g0194(.din(lo030_buf_o2), .dout(new_new_n738__));
  not1  g0195(.din(lo030_buf_o2), .dout(new_new_n739__));
  buf1  g0196(.din(lo034_buf_o2), .dout(new_new_n740__));
  not1  g0197(.din(lo034_buf_o2), .dout(new_new_n741__));
  buf1  g0198(.din(lo038_buf_o2), .dout(new_new_n742__));
  not1  g0199(.din(lo038_buf_o2), .dout(new_new_n743__));
  buf1  g0200(.din(lo042_buf_o2), .dout(new_new_n744__));
  not1  g0201(.din(lo042_buf_o2), .dout(new_new_n745__));
  buf1  g0202(.din(lo046_buf_o2), .dout(new_new_n746__));
  not1  g0203(.din(lo046_buf_o2), .dout(new_new_n747__));
  buf1  g0204(.din(lo050_buf_o2), .dout(new_new_n748__));
  not1  g0205(.din(lo050_buf_o2), .dout(new_new_n749__));
  buf1  g0206(.din(lo054_buf_o2), .dout(new_new_n750__));
  not1  g0207(.din(lo054_buf_o2), .dout(new_new_n751__));
  buf1  g0208(.din(lo058_buf_o2), .dout(new_new_n752__));
  not1  g0209(.din(lo058_buf_o2), .dout(new_new_n753__));
  buf1  g0210(.din(lo062_buf_o2), .dout(new_new_n754__));
  not1  g0211(.din(lo062_buf_o2), .dout(new_new_n755__));
  buf1  g0212(.din(lo066_buf_o2), .dout(new_new_n756__));
  not1  g0213(.din(lo066_buf_o2), .dout(new_new_n757__));
  buf1  g0214(.din(lo070_buf_o2), .dout(new_new_n758__));
  not1  g0215(.din(lo070_buf_o2), .dout(new_new_n759__));
  buf1  g0216(.din(lo074_buf_o2), .dout(new_new_n760__));
  not1  g0217(.din(lo074_buf_o2), .dout(new_new_n761__));
  buf1  g0218(.din(lo078_buf_o2), .dout(new_new_n762__));
  not1  g0219(.din(lo078_buf_o2), .dout(new_new_n763__));
  buf1  g0220(.din(lo082_buf_o2), .dout(new_new_n764__));
  not1  g0221(.din(lo082_buf_o2), .dout(new_new_n765__));
  buf1  g0222(.din(lo086_buf_o2), .dout(new_new_n766__));
  not1  g0223(.din(lo086_buf_o2), .dout(new_new_n767__));
  buf1  g0224(.din(lo090_buf_o2), .dout(new_new_n768__));
  not1  g0225(.din(lo090_buf_o2), .dout(new_new_n769__));
  buf1  g0226(.din(lo094_buf_o2), .dout(new_new_n770__));
  not1  g0227(.din(lo094_buf_o2), .dout(new_new_n771__));
  buf1  g0228(.din(lo098_buf_o2), .dout(new_new_n772__));
  not1  g0229(.din(lo098_buf_o2), .dout(new_new_n773__));
  buf1  g0230(.din(lo102_buf_o2), .dout(new_new_n774__));
  not1  g0231(.din(lo102_buf_o2), .dout(new_new_n775__));
  buf1  g0232(.din(lo106_buf_o2), .dout(new_new_n776__));
  not1  g0233(.din(lo106_buf_o2), .dout(new_new_n777__));
  buf1  g0234(.din(lo110_buf_o2), .dout(new_new_n778__));
  not1  g0235(.din(lo110_buf_o2), .dout(new_new_n779__));
  buf1  g0236(.din(lo114_buf_o2), .dout(new_new_n780__));
  not1  g0237(.din(lo114_buf_o2), .dout(new_new_n781__));
  buf1  g0238(.din(lo118_buf_o2), .dout(new_new_n782__));
  not1  g0239(.din(lo118_buf_o2), .dout(new_new_n783__));
  buf1  g0240(.din(lo122_buf_o2), .dout(new_new_n784__));
  not1  g0241(.din(lo122_buf_o2), .dout(new_new_n785__));
  buf1  g0242(.din(lo126_buf_o2), .dout(new_new_n786__));
  not1  g0243(.din(lo126_buf_o2), .dout(new_new_n787__));
  buf1  g0244(.din(n683_o2), .dout(new_new_n788__));
  not1  g0245(.din(n683_o2), .dout(new_new_n789__));
  buf1  g0246(.din(n688_o2), .dout(new_new_n790__));
  not1  g0247(.din(n688_o2), .dout(new_new_n791__));
  buf1  g0248(.din(n803_o2), .dout(new_new_n792__));
  not1  g0249(.din(n803_o2), .dout(new_new_n793__));
  buf1  g0250(.din(n862_o2), .dout(new_new_n794__));
  not1  g0251(.din(n862_o2), .dout(new_new_n795__));
  buf1  g0252(.din(n764_o2), .dout(new_new_n796__));
  not1  g0253(.din(n764_o2), .dout(new_new_n797__));
  buf1  g0254(.din(n863_o2), .dout(new_new_n798__));
  not1  g0255(.din(n863_o2), .dout(new_new_n799__));
  buf1  g0256(.din(n886_o2), .dout(new_new_n800__));
  not1  g0257(.din(n886_o2), .dout(new_new_n801__));
  buf1  g0258(.din(n600_o2), .dout(new_new_n802__));
  not1  g0259(.din(n600_o2), .dout(new_new_n803__));
  buf1  g0260(.din(n601_o2), .dout(new_new_n804__));
  not1  g0261(.din(n601_o2), .dout(new_new_n805__));
  buf1  g0262(.din(n637_o2), .dout(new_new_n806__));
  not1  g0263(.din(n637_o2), .dout(new_new_n807__));
  buf1  g0264(.din(n638_o2), .dout(new_new_n808__));
  not1  g0265(.din(n638_o2), .dout(new_new_n809__));
  buf1  g0266(.din(n676_o2), .dout(new_new_n810__));
  not1  g0267(.din(n676_o2), .dout(new_new_n811__));
  buf1  g0268(.din(n677_o2), .dout(new_new_n812__));
  not1  g0269(.din(n677_o2), .dout(new_new_n813__));
  buf1  g0270(.din(n656_o2), .dout(new_new_n814__));
  not1  g0271(.din(n656_o2), .dout(new_new_n815__));
  buf1  g0272(.din(n657_o2), .dout(new_new_n816__));
  not1  g0273(.din(n657_o2), .dout(new_new_n817__));
  buf1  g0274(.din(n781_o2), .dout(new_new_n818__));
  not1  g0275(.din(n781_o2), .dout(new_new_n819__));
  buf1  g0276(.din(n782_o2), .dout(new_new_n820__));
  not1  g0277(.din(n782_o2), .dout(new_new_n821__));
  buf1  g0278(.din(n800_o2), .dout(new_new_n822__));
  not1  g0279(.din(n800_o2), .dout(new_new_n823__));
  buf1  g0280(.din(n801_o2), .dout(new_new_n824__));
  not1  g0281(.din(n801_o2), .dout(new_new_n825__));
  buf1  g0282(.din(n724_o2), .dout(new_new_n826__));
  not1  g0283(.din(n724_o2), .dout(new_new_n827__));
  buf1  g0284(.din(n725_o2), .dout(new_new_n828__));
  not1  g0285(.din(n725_o2), .dout(new_new_n829__));
  buf1  g0286(.din(n761_o2), .dout(new_new_n830__));
  not1  g0287(.din(n761_o2), .dout(new_new_n831__));
  buf1  g0288(.din(n762_o2), .dout(new_new_n832__));
  not1  g0289(.din(n762_o2), .dout(new_new_n833__));
  buf1  g0290(.din(lo129_buf_o2), .dout(new_new_n834__));
  not1  g0291(.din(lo129_buf_o2), .dout(new_new_n835__));
  buf1  g0292(.din(lo133_buf_o2), .dout(new_new_n836__));
  not1  g0293(.din(lo133_buf_o2), .dout(new_new_n837__));
  buf1  g0294(.din(lo137_buf_o2), .dout(new_new_n838__));
  not1  g0295(.din(lo137_buf_o2), .dout(new_new_n839__));
  buf1  g0296(.din(lo141_buf_o2), .dout(new_new_n840__));
  not1  g0297(.din(lo141_buf_o2), .dout(new_new_n841__));
  buf1  g0298(.din(lo145_buf_o2), .dout(new_new_n842__));
  not1  g0299(.din(lo145_buf_o2), .dout(new_new_n843__));
  buf1  g0300(.din(lo149_buf_o2), .dout(new_new_n844__));
  not1  g0301(.din(lo149_buf_o2), .dout(new_new_n845__));
  buf1  g0302(.din(lo153_buf_o2), .dout(new_new_n846__));
  not1  g0303(.din(lo153_buf_o2), .dout(new_new_n847__));
  buf1  g0304(.din(lo157_buf_o2), .dout(new_new_n848__));
  not1  g0305(.din(lo157_buf_o2), .dout(new_new_n849__));
  buf1  g0306(.din(lo161_buf_o2), .dout(new_new_n850__));
  not1  g0307(.din(lo161_buf_o2), .dout(new_new_n851__));
  buf1  g0308(.din(n708_o2), .dout(new_new_n852__));
  not1  g0309(.din(n708_o2), .dout(new_new_n853__));
  buf1  g0310(.din(n745_o2), .dout(new_new_n854__));
  not1  g0311(.din(n745_o2), .dout(new_new_n855__));
  buf1  g0312(.din(n717_o2), .dout(new_new_n856__));
  not1  g0313(.din(n717_o2), .dout(new_new_n857__));
  buf1  g0314(.din(n754_o2), .dout(new_new_n858__));
  not1  g0315(.din(n754_o2), .dout(new_new_n859__));
  buf1  g0316(.din(n584_o2), .dout(new_new_n860__));
  not1  g0317(.din(n584_o2), .dout(new_new_n861__));
  buf1  g0318(.din(n593_o2), .dout(new_new_n862__));
  not1  g0319(.din(n593_o2), .dout(new_new_n863__));
  buf1  g0320(.din(n630_o2), .dout(new_new_n864__));
  not1  g0321(.din(n630_o2), .dout(new_new_n865__));
  buf1  g0322(.din(n621_o2), .dout(new_new_n866__));
  not1  g0323(.din(n621_o2), .dout(new_new_n867__));
  buf1  g0324(.din(lo001_buf_o2), .dout(new_new_n868__));
  not1  g0325(.din(lo001_buf_o2), .dout(new_new_n869__));
  buf1  g0326(.din(lo005_buf_o2), .dout(new_new_n870__));
  not1  g0327(.din(lo005_buf_o2), .dout(new_new_n871__));
  buf1  g0328(.din(lo009_buf_o2), .dout(new_new_n872__));
  not1  g0329(.din(lo009_buf_o2), .dout(new_new_n873__));
  buf1  g0330(.din(lo013_buf_o2), .dout(new_new_n874__));
  not1  g0331(.din(lo013_buf_o2), .dout(new_new_n875__));
  buf1  g0332(.din(lo017_buf_o2), .dout(new_new_n876__));
  not1  g0333(.din(lo017_buf_o2), .dout(new_new_n877__));
  buf1  g0334(.din(lo021_buf_o2), .dout(new_new_n878__));
  not1  g0335(.din(lo021_buf_o2), .dout(new_new_n879__));
  buf1  g0336(.din(lo025_buf_o2), .dout(new_new_n880__));
  not1  g0337(.din(lo025_buf_o2), .dout(new_new_n881__));
  buf1  g0338(.din(lo029_buf_o2), .dout(new_new_n882__));
  not1  g0339(.din(lo029_buf_o2), .dout(new_new_n883__));
  buf1  g0340(.din(lo033_buf_o2), .dout(new_new_n884__));
  not1  g0341(.din(lo033_buf_o2), .dout(new_new_n885__));
  buf1  g0342(.din(lo037_buf_o2), .dout(new_new_n886__));
  not1  g0343(.din(lo037_buf_o2), .dout(new_new_n887__));
  buf1  g0344(.din(lo041_buf_o2), .dout(new_new_n888__));
  not1  g0345(.din(lo041_buf_o2), .dout(new_new_n889__));
  buf1  g0346(.din(lo045_buf_o2), .dout(new_new_n890__));
  not1  g0347(.din(lo045_buf_o2), .dout(new_new_n891__));
  buf1  g0348(.din(lo049_buf_o2), .dout(new_new_n892__));
  not1  g0349(.din(lo049_buf_o2), .dout(new_new_n893__));
  buf1  g0350(.din(lo053_buf_o2), .dout(new_new_n894__));
  not1  g0351(.din(lo053_buf_o2), .dout(new_new_n895__));
  buf1  g0352(.din(lo057_buf_o2), .dout(new_new_n896__));
  not1  g0353(.din(lo057_buf_o2), .dout(new_new_n897__));
  buf1  g0354(.din(lo061_buf_o2), .dout(new_new_n898__));
  not1  g0355(.din(lo061_buf_o2), .dout(new_new_n899__));
  buf1  g0356(.din(lo065_buf_o2), .dout(new_new_n900__));
  not1  g0357(.din(lo065_buf_o2), .dout(new_new_n901__));
  buf1  g0358(.din(lo069_buf_o2), .dout(new_new_n902__));
  not1  g0359(.din(lo069_buf_o2), .dout(new_new_n903__));
  buf1  g0360(.din(lo073_buf_o2), .dout(new_new_n904__));
  not1  g0361(.din(lo073_buf_o2), .dout(new_new_n905__));
  buf1  g0362(.din(lo077_buf_o2), .dout(new_new_n906__));
  not1  g0363(.din(lo077_buf_o2), .dout(new_new_n907__));
  buf1  g0364(.din(lo081_buf_o2), .dout(new_new_n908__));
  not1  g0365(.din(lo081_buf_o2), .dout(new_new_n909__));
  buf1  g0366(.din(lo085_buf_o2), .dout(new_new_n910__));
  not1  g0367(.din(lo085_buf_o2), .dout(new_new_n911__));
  buf1  g0368(.din(lo089_buf_o2), .dout(new_new_n912__));
  not1  g0369(.din(lo089_buf_o2), .dout(new_new_n913__));
  buf1  g0370(.din(lo093_buf_o2), .dout(new_new_n914__));
  not1  g0371(.din(lo093_buf_o2), .dout(new_new_n915__));
  buf1  g0372(.din(lo097_buf_o2), .dout(new_new_n916__));
  not1  g0373(.din(lo097_buf_o2), .dout(new_new_n917__));
  buf1  g0374(.din(lo101_buf_o2), .dout(new_new_n918__));
  not1  g0375(.din(lo101_buf_o2), .dout(new_new_n919__));
  buf1  g0376(.din(lo105_buf_o2), .dout(new_new_n920__));
  not1  g0377(.din(lo105_buf_o2), .dout(new_new_n921__));
  buf1  g0378(.din(lo109_buf_o2), .dout(new_new_n922__));
  not1  g0379(.din(lo109_buf_o2), .dout(new_new_n923__));
  buf1  g0380(.din(lo113_buf_o2), .dout(new_new_n924__));
  not1  g0381(.din(lo113_buf_o2), .dout(new_new_n925__));
  buf1  g0382(.din(lo117_buf_o2), .dout(new_new_n926__));
  not1  g0383(.din(lo117_buf_o2), .dout(new_new_n927__));
  buf1  g0384(.din(lo121_buf_o2), .dout(new_new_n928__));
  not1  g0385(.din(lo121_buf_o2), .dout(new_new_n929__));
  buf1  g0386(.din(lo125_buf_o2), .dout(new_new_n930__));
  not1  g0387(.din(lo125_buf_o2), .dout(new_new_n931__));
  and1  g0388(.dina(new_new_n789__), .dinb(new_new_n791__), .dout(new_new_n932__));
  or1   g0389(.dina(new_new_n788__), .dinb(new_new_n790__), .dout(new_new_n933__));
  and1  g0390(.dina(new_new_n792__), .dinb(new_new_n796__), .dout(new_new_n934__));
  or1   g0391(.dina(new_new_n793__), .dinb(new_new_n797__), .dout(new_new_n935__));
  and1  g0392(.dina(new_new_n1739__), .dinb(new_new_n934__), .dout(new_new_n936__));
  or1   g0393(.dina(new_new_n1742__), .dinb(new_new_n935__), .dout(new_new_n937__));
  and1  g0394(.dina(new_new_n1745__), .dinb(new_new_n1748__), .dout(new_new_n938__));
  or1   g0395(.dina(new_new_n1751__), .dinb(new_new_n1754__), .dout(new_new_n939__));
  and1  g0396(.dina(new_new_n545__), .dinb(new_new_n938__), .dout(new_new_n940__));
  and1  g0397(.dina(new_new_n544__), .dinb(new_new_n939__), .dout(new_new_n941__));
  or1   g0398(.dina(new_new_n940__), .dinb(new_new_n941__), .dout(new_new_n942__));
  and1  g0399(.dina(new_new_n1758__), .dinb(new_new_n1748__), .dout(new_new_n943__));
  or1   g0400(.dina(new_new_n1762__), .dinb(new_new_n1754__), .dout(new_new_n944__));
  and1  g0401(.dina(new_new_n547__), .dinb(new_new_n943__), .dout(new_new_n945__));
  and1  g0402(.dina(new_new_n546__), .dinb(new_new_n944__), .dout(new_new_n946__));
  or1   g0403(.dina(new_new_n945__), .dinb(new_new_n946__), .dout(new_new_n947__));
  and1  g0404(.dina(new_new_n1766__), .dinb(new_new_n1749__), .dout(new_new_n948__));
  or1   g0405(.dina(new_new_n1771__), .dinb(new_new_n1755__), .dout(new_new_n949__));
  and1  g0406(.dina(new_new_n549__), .dinb(new_new_n948__), .dout(new_new_n950__));
  and1  g0407(.dina(new_new_n548__), .dinb(new_new_n949__), .dout(new_new_n951__));
  or1   g0408(.dina(new_new_n950__), .dinb(new_new_n951__), .dout(new_new_n952__));
  and1  g0409(.dina(new_new_n1775__), .dinb(new_new_n1749__), .dout(new_new_n953__));
  or1   g0410(.dina(new_new_n1778__), .dinb(new_new_n1755__), .dout(new_new_n954__));
  and1  g0411(.dina(new_new_n551__), .dinb(new_new_n953__), .dout(new_new_n955__));
  and1  g0412(.dina(new_new_n550__), .dinb(new_new_n954__), .dout(new_new_n956__));
  or1   g0413(.dina(new_new_n955__), .dinb(new_new_n956__), .dout(new_new_n957__));
  and1  g0414(.dina(new_new_n710__), .dinb(new_new_n723__), .dout(new_new_n958__));
  or1   g0415(.dina(new_new_n711__), .dinb(new_new_n722__), .dout(new_new_n959__));
  and1  g0416(.dina(new_new_n1739__), .dinb(new_new_n958__), .dout(new_new_n960__));
  or1   g0417(.dina(new_new_n1742__), .dinb(new_new_n959__), .dout(new_new_n961__));
  and1  g0418(.dina(new_new_n1745__), .dinb(new_new_n1781__), .dout(new_new_n962__));
  or1   g0419(.dina(new_new_n1751__), .dinb(new_new_n1784__), .dout(new_new_n963__));
  and1  g0420(.dina(new_new_n553__), .dinb(new_new_n962__), .dout(new_new_n964__));
  and1  g0421(.dina(new_new_n552__), .dinb(new_new_n963__), .dout(new_new_n965__));
  or1   g0422(.dina(new_new_n964__), .dinb(new_new_n965__), .dout(new_new_n966__));
  and1  g0423(.dina(new_new_n1758__), .dinb(new_new_n1781__), .dout(new_new_n967__));
  or1   g0424(.dina(new_new_n1762__), .dinb(new_new_n1784__), .dout(new_new_n968__));
  and1  g0425(.dina(new_new_n555__), .dinb(new_new_n967__), .dout(new_new_n969__));
  and1  g0426(.dina(new_new_n554__), .dinb(new_new_n968__), .dout(new_new_n970__));
  or1   g0427(.dina(new_new_n969__), .dinb(new_new_n970__), .dout(new_new_n971__));
  and1  g0428(.dina(new_new_n1766__), .dinb(new_new_n1782__), .dout(new_new_n972__));
  or1   g0429(.dina(new_new_n1771__), .dinb(new_new_n1785__), .dout(new_new_n973__));
  and1  g0430(.dina(new_new_n557__), .dinb(new_new_n972__), .dout(new_new_n974__));
  and1  g0431(.dina(new_new_n556__), .dinb(new_new_n973__), .dout(new_new_n975__));
  or1   g0432(.dina(new_new_n974__), .dinb(new_new_n975__), .dout(new_new_n976__));
  and1  g0433(.dina(new_new_n1775__), .dinb(new_new_n1782__), .dout(new_new_n977__));
  or1   g0434(.dina(new_new_n1778__), .dinb(new_new_n1785__), .dout(new_new_n978__));
  and1  g0435(.dina(new_new_n559__), .dinb(new_new_n977__), .dout(new_new_n979__));
  and1  g0436(.dina(new_new_n558__), .dinb(new_new_n978__), .dout(new_new_n980__));
  or1   g0437(.dina(new_new_n979__), .dinb(new_new_n980__), .dout(new_new_n981__));
  and1  g0438(.dina(new_new_n713__), .dinb(new_new_n714__), .dout(new_new_n982__));
  or1   g0439(.dina(new_new_n712__), .dinb(new_new_n715__), .dout(new_new_n983__));
  and1  g0440(.dina(new_new_n1740__), .dinb(new_new_n982__), .dout(new_new_n984__));
  or1   g0441(.dina(new_new_n1743__), .dinb(new_new_n983__), .dout(new_new_n985__));
  and1  g0442(.dina(new_new_n1746__), .dinb(new_new_n1787__), .dout(new_new_n986__));
  or1   g0443(.dina(new_new_n1752__), .dinb(new_new_n1790__), .dout(new_new_n987__));
  and1  g0444(.dina(new_new_n561__), .dinb(new_new_n986__), .dout(new_new_n988__));
  and1  g0445(.dina(new_new_n560__), .dinb(new_new_n987__), .dout(new_new_n989__));
  or1   g0446(.dina(new_new_n988__), .dinb(new_new_n989__), .dout(new_new_n990__));
  and1  g0447(.dina(new_new_n1757__), .dinb(new_new_n1787__), .dout(new_new_n991__));
  or1   g0448(.dina(new_new_n1761__), .dinb(new_new_n1790__), .dout(new_new_n992__));
  and1  g0449(.dina(new_new_n563__), .dinb(new_new_n991__), .dout(new_new_n993__));
  and1  g0450(.dina(new_new_n562__), .dinb(new_new_n992__), .dout(new_new_n994__));
  or1   g0451(.dina(new_new_n993__), .dinb(new_new_n994__), .dout(new_new_n995__));
  and1  g0452(.dina(new_new_n1767__), .dinb(new_new_n1788__), .dout(new_new_n996__));
  or1   g0453(.dina(new_new_n1772__), .dinb(new_new_n1791__), .dout(new_new_n997__));
  and1  g0454(.dina(new_new_n565__), .dinb(new_new_n996__), .dout(new_new_n998__));
  and1  g0455(.dina(new_new_n564__), .dinb(new_new_n997__), .dout(new_new_n999__));
  or1   g0456(.dina(new_new_n998__), .dinb(new_new_n999__), .dout(new_new_n1000__));
  and1  g0457(.dina(new_new_n1776__), .dinb(new_new_n1788__), .dout(new_new_n1001__));
  or1   g0458(.dina(new_new_n1779__), .dinb(new_new_n1791__), .dout(new_new_n1002__));
  and1  g0459(.dina(new_new_n567__), .dinb(new_new_n1001__), .dout(new_new_n1003__));
  and1  g0460(.dina(new_new_n566__), .dinb(new_new_n1002__), .dout(new_new_n1004__));
  or1   g0461(.dina(new_new_n1003__), .dinb(new_new_n1004__), .dout(new_new_n1005__));
  and1  g0462(.dina(new_new_n794__), .dinb(new_new_n798__), .dout(new_new_n1006__));
  or1   g0463(.dina(new_new_n795__), .dinb(new_new_n799__), .dout(new_new_n1007__));
  and1  g0464(.dina(new_new_n1740__), .dinb(new_new_n1006__), .dout(new_new_n1008__));
  or1   g0465(.dina(new_new_n1743__), .dinb(new_new_n1007__), .dout(new_new_n1009__));
  and1  g0466(.dina(new_new_n1746__), .dinb(new_new_n1793__), .dout(new_new_n1010__));
  or1   g0467(.dina(new_new_n1752__), .dinb(new_new_n1796__), .dout(new_new_n1011__));
  and1  g0468(.dina(new_new_n569__), .dinb(new_new_n1010__), .dout(new_new_n1012__));
  and1  g0469(.dina(new_new_n568__), .dinb(new_new_n1011__), .dout(new_new_n1013__));
  or1   g0470(.dina(new_new_n1012__), .dinb(new_new_n1013__), .dout(new_new_n1014__));
  and1  g0471(.dina(new_new_n1759__), .dinb(new_new_n1793__), .dout(new_new_n1015__));
  or1   g0472(.dina(new_new_n1763__), .dinb(new_new_n1796__), .dout(new_new_n1016__));
  and1  g0473(.dina(new_new_n571__), .dinb(new_new_n1015__), .dout(new_new_n1017__));
  and1  g0474(.dina(new_new_n570__), .dinb(new_new_n1016__), .dout(new_new_n1018__));
  or1   g0475(.dina(new_new_n1017__), .dinb(new_new_n1018__), .dout(new_new_n1019__));
  and1  g0476(.dina(new_new_n1767__), .dinb(new_new_n1794__), .dout(new_new_n1020__));
  or1   g0477(.dina(new_new_n1772__), .dinb(new_new_n1797__), .dout(new_new_n1021__));
  and1  g0478(.dina(new_new_n573__), .dinb(new_new_n1020__), .dout(new_new_n1022__));
  and1  g0479(.dina(new_new_n572__), .dinb(new_new_n1021__), .dout(new_new_n1023__));
  or1   g0480(.dina(new_new_n1022__), .dinb(new_new_n1023__), .dout(new_new_n1024__));
  and1  g0481(.dina(new_new_n1776__), .dinb(new_new_n1794__), .dout(new_new_n1025__));
  or1   g0482(.dina(new_new_n1779__), .dinb(new_new_n1797__), .dout(new_new_n1026__));
  and1  g0483(.dina(new_new_n575__), .dinb(new_new_n1025__), .dout(new_new_n1027__));
  and1  g0484(.dina(new_new_n574__), .dinb(new_new_n1026__), .dout(new_new_n1028__));
  or1   g0485(.dina(new_new_n1027__), .dinb(new_new_n1028__), .dout(new_new_n1029__));
  and1  g0486(.dina(new_new_n720__), .dinb(new_new_n1799__), .dout(new_new_n1030__));
  or1   g0487(.dina(new_new_n721__), .dinb(new_new_n1802__), .dout(new_new_n1031__));
  and1  g0488(.dina(new_new_n1768__), .dinb(new_new_n1030__), .dout(new_new_n1032__));
  or1   g0489(.dina(new_new_n1773__), .dinb(new_new_n1031__), .dout(new_new_n1033__));
  and1  g0490(.dina(new_new_n1805__), .dinb(new_new_n1808__), .dout(new_new_n1034__));
  or1   g0491(.dina(new_new_n1811__), .dinb(new_new_n1814__), .dout(new_new_n1035__));
  and1  g0492(.dina(new_new_n577__), .dinb(new_new_n1034__), .dout(new_new_n1036__));
  and1  g0493(.dina(new_new_n576__), .dinb(new_new_n1035__), .dout(new_new_n1037__));
  or1   g0494(.dina(new_new_n1036__), .dinb(new_new_n1037__), .dout(new_new_n1038__));
  and1  g0495(.dina(new_new_n1817__), .dinb(new_new_n1808__), .dout(new_new_n1039__));
  or1   g0496(.dina(new_new_n1820__), .dinb(new_new_n1814__), .dout(new_new_n1040__));
  and1  g0497(.dina(new_new_n579__), .dinb(new_new_n1039__), .dout(new_new_n1041__));
  and1  g0498(.dina(new_new_n578__), .dinb(new_new_n1040__), .dout(new_new_n1042__));
  or1   g0499(.dina(new_new_n1041__), .dinb(new_new_n1042__), .dout(new_new_n1043__));
  and1  g0500(.dina(new_new_n1823__), .dinb(new_new_n1809__), .dout(new_new_n1044__));
  or1   g0501(.dina(new_new_n1826__), .dinb(new_new_n1815__), .dout(new_new_n1045__));
  and1  g0502(.dina(new_new_n581__), .dinb(new_new_n1044__), .dout(new_new_n1046__));
  and1  g0503(.dina(new_new_n580__), .dinb(new_new_n1045__), .dout(new_new_n1047__));
  or1   g0504(.dina(new_new_n1046__), .dinb(new_new_n1047__), .dout(new_new_n1048__));
  and1  g0505(.dina(new_new_n1829__), .dinb(new_new_n1809__), .dout(new_new_n1049__));
  or1   g0506(.dina(new_new_n1832__), .dinb(new_new_n1815__), .dout(new_new_n1050__));
  and1  g0507(.dina(new_new_n583__), .dinb(new_new_n1049__), .dout(new_new_n1051__));
  and1  g0508(.dina(new_new_n582__), .dinb(new_new_n1050__), .dout(new_new_n1052__));
  or1   g0509(.dina(new_new_n1051__), .dinb(new_new_n1052__), .dout(new_new_n1053__));
  and1  g0510(.dina(new_new_n706__), .dinb(new_new_n708__), .dout(new_new_n1054__));
  or1   g0511(.dina(new_new_n707__), .dinb(new_new_n709__), .dout(new_new_n1055__));
  and1  g0512(.dina(new_new_n1799__), .dinb(new_new_n1054__), .dout(new_new_n1056__));
  or1   g0513(.dina(new_new_n1802__), .dinb(new_new_n1055__), .dout(new_new_n1057__));
  and1  g0514(.dina(new_new_n1805__), .dinb(new_new_n1835__), .dout(new_new_n1058__));
  or1   g0515(.dina(new_new_n1811__), .dinb(new_new_n1838__), .dout(new_new_n1059__));
  and1  g0516(.dina(new_new_n585__), .dinb(new_new_n1058__), .dout(new_new_n1060__));
  and1  g0517(.dina(new_new_n584__), .dinb(new_new_n1059__), .dout(new_new_n1061__));
  or1   g0518(.dina(new_new_n1060__), .dinb(new_new_n1061__), .dout(new_new_n1062__));
  and1  g0519(.dina(new_new_n1817__), .dinb(new_new_n1835__), .dout(new_new_n1063__));
  or1   g0520(.dina(new_new_n1820__), .dinb(new_new_n1838__), .dout(new_new_n1064__));
  and1  g0521(.dina(new_new_n587__), .dinb(new_new_n1063__), .dout(new_new_n1065__));
  and1  g0522(.dina(new_new_n586__), .dinb(new_new_n1064__), .dout(new_new_n1066__));
  or1   g0523(.dina(new_new_n1065__), .dinb(new_new_n1066__), .dout(new_new_n1067__));
  and1  g0524(.dina(new_new_n1823__), .dinb(new_new_n1836__), .dout(new_new_n1068__));
  or1   g0525(.dina(new_new_n1826__), .dinb(new_new_n1839__), .dout(new_new_n1069__));
  and1  g0526(.dina(new_new_n589__), .dinb(new_new_n1068__), .dout(new_new_n1070__));
  and1  g0527(.dina(new_new_n588__), .dinb(new_new_n1069__), .dout(new_new_n1071__));
  or1   g0528(.dina(new_new_n1070__), .dinb(new_new_n1071__), .dout(new_new_n1072__));
  and1  g0529(.dina(new_new_n1829__), .dinb(new_new_n1836__), .dout(new_new_n1073__));
  or1   g0530(.dina(new_new_n1832__), .dinb(new_new_n1839__), .dout(new_new_n1074__));
  and1  g0531(.dina(new_new_n591__), .dinb(new_new_n1073__), .dout(new_new_n1075__));
  and1  g0532(.dina(new_new_n590__), .dinb(new_new_n1074__), .dout(new_new_n1076__));
  or1   g0533(.dina(new_new_n1075__), .dinb(new_new_n1076__), .dout(new_new_n1077__));
  and1  g0534(.dina(new_new_n1768__), .dinb(new_new_n718__), .dout(new_new_n1078__));
  or1   g0535(.dina(new_new_n1773__), .dinb(new_new_n719__), .dout(new_new_n1079__));
  and1  g0536(.dina(new_new_n1800__), .dinb(new_new_n1078__), .dout(new_new_n1080__));
  or1   g0537(.dina(new_new_n1803__), .dinb(new_new_n1079__), .dout(new_new_n1081__));
  and1  g0538(.dina(new_new_n1806__), .dinb(new_new_n1841__), .dout(new_new_n1082__));
  or1   g0539(.dina(new_new_n1812__), .dinb(new_new_n1844__), .dout(new_new_n1083__));
  and1  g0540(.dina(new_new_n593__), .dinb(new_new_n1082__), .dout(new_new_n1084__));
  and1  g0541(.dina(new_new_n592__), .dinb(new_new_n1083__), .dout(new_new_n1085__));
  or1   g0542(.dina(new_new_n1084__), .dinb(new_new_n1085__), .dout(new_new_n1086__));
  and1  g0543(.dina(new_new_n1818__), .dinb(new_new_n1841__), .dout(new_new_n1087__));
  or1   g0544(.dina(new_new_n1821__), .dinb(new_new_n1844__), .dout(new_new_n1088__));
  and1  g0545(.dina(new_new_n595__), .dinb(new_new_n1087__), .dout(new_new_n1089__));
  and1  g0546(.dina(new_new_n594__), .dinb(new_new_n1088__), .dout(new_new_n1090__));
  or1   g0547(.dina(new_new_n1089__), .dinb(new_new_n1090__), .dout(new_new_n1091__));
  and1  g0548(.dina(new_new_n1824__), .dinb(new_new_n1842__), .dout(new_new_n1092__));
  or1   g0549(.dina(new_new_n1827__), .dinb(new_new_n1845__), .dout(new_new_n1093__));
  and1  g0550(.dina(new_new_n597__), .dinb(new_new_n1092__), .dout(new_new_n1094__));
  and1  g0551(.dina(new_new_n596__), .dinb(new_new_n1093__), .dout(new_new_n1095__));
  or1   g0552(.dina(new_new_n1094__), .dinb(new_new_n1095__), .dout(new_new_n1096__));
  and1  g0553(.dina(new_new_n1830__), .dinb(new_new_n1842__), .dout(new_new_n1097__));
  or1   g0554(.dina(new_new_n1833__), .dinb(new_new_n1845__), .dout(new_new_n1098__));
  and1  g0555(.dina(new_new_n599__), .dinb(new_new_n1097__), .dout(new_new_n1099__));
  and1  g0556(.dina(new_new_n598__), .dinb(new_new_n1098__), .dout(new_new_n1100__));
  or1   g0557(.dina(new_new_n1099__), .dinb(new_new_n1100__), .dout(new_new_n1101__));
  and1  g0558(.dina(new_new_n1759__), .dinb(new_new_n716__), .dout(new_new_n1102__));
  or1   g0559(.dina(new_new_n1763__), .dinb(new_new_n717__), .dout(new_new_n1103__));
  and1  g0560(.dina(new_new_n1800__), .dinb(new_new_n1102__), .dout(new_new_n1104__));
  or1   g0561(.dina(new_new_n1803__), .dinb(new_new_n1103__), .dout(new_new_n1105__));
  and1  g0562(.dina(new_new_n1806__), .dinb(new_new_n1847__), .dout(new_new_n1106__));
  or1   g0563(.dina(new_new_n1812__), .dinb(new_new_n1850__), .dout(new_new_n1107__));
  and1  g0564(.dina(new_new_n601__), .dinb(new_new_n1106__), .dout(new_new_n1108__));
  and1  g0565(.dina(new_new_n600__), .dinb(new_new_n1107__), .dout(new_new_n1109__));
  or1   g0566(.dina(new_new_n1108__), .dinb(new_new_n1109__), .dout(new_new_n1110__));
  and1  g0567(.dina(new_new_n1818__), .dinb(new_new_n1847__), .dout(new_new_n1111__));
  or1   g0568(.dina(new_new_n1821__), .dinb(new_new_n1850__), .dout(new_new_n1112__));
  and1  g0569(.dina(new_new_n603__), .dinb(new_new_n1111__), .dout(new_new_n1113__));
  and1  g0570(.dina(new_new_n602__), .dinb(new_new_n1112__), .dout(new_new_n1114__));
  or1   g0571(.dina(new_new_n1113__), .dinb(new_new_n1114__), .dout(new_new_n1115__));
  and1  g0572(.dina(new_new_n1824__), .dinb(new_new_n1848__), .dout(new_new_n1116__));
  or1   g0573(.dina(new_new_n1827__), .dinb(new_new_n1851__), .dout(new_new_n1117__));
  and1  g0574(.dina(new_new_n605__), .dinb(new_new_n1116__), .dout(new_new_n1118__));
  and1  g0575(.dina(new_new_n604__), .dinb(new_new_n1117__), .dout(new_new_n1119__));
  or1   g0576(.dina(new_new_n1118__), .dinb(new_new_n1119__), .dout(new_new_n1120__));
  and1  g0577(.dina(new_new_n1830__), .dinb(new_new_n1848__), .dout(new_new_n1121__));
  or1   g0578(.dina(new_new_n1833__), .dinb(new_new_n1851__), .dout(new_new_n1122__));
  and1  g0579(.dina(new_new_n607__), .dinb(new_new_n1121__), .dout(new_new_n1123__));
  and1  g0580(.dina(new_new_n606__), .dinb(new_new_n1122__), .dout(new_new_n1124__));
  or1   g0581(.dina(new_new_n1123__), .dinb(new_new_n1124__), .dout(new_new_n1125__));
  and1  g0582(.dina(new_new_n803__), .dinb(new_new_n805__), .dout(new_new_n1126__));
  or1   g0583(.dina(new_new_n802__), .dinb(new_new_n804__), .dout(new_new_n1127__));
  and1  g0584(.dina(new_new_n807__), .dinb(new_new_n809__), .dout(new_new_n1128__));
  or1   g0585(.dina(new_new_n806__), .dinb(new_new_n808__), .dout(new_new_n1129__));
  and1  g0586(.dina(new_new_n811__), .dinb(new_new_n813__), .dout(new_new_n1130__));
  or1   g0587(.dina(new_new_n810__), .dinb(new_new_n812__), .dout(new_new_n1131__));
  and1  g0588(.dina(new_new_n815__), .dinb(new_new_n817__), .dout(new_new_n1132__));
  or1   g0589(.dina(new_new_n814__), .dinb(new_new_n816__), .dout(new_new_n1133__));
  and1  g0590(.dina(new_new_n819__), .dinb(new_new_n821__), .dout(new_new_n1134__));
  or1   g0591(.dina(new_new_n818__), .dinb(new_new_n820__), .dout(new_new_n1135__));
  and1  g0592(.dina(new_new_n823__), .dinb(new_new_n825__), .dout(new_new_n1136__));
  or1   g0593(.dina(new_new_n822__), .dinb(new_new_n824__), .dout(new_new_n1137__));
  and1  g0594(.dina(new_new_n827__), .dinb(new_new_n829__), .dout(new_new_n1138__));
  or1   g0595(.dina(new_new_n826__), .dinb(new_new_n828__), .dout(new_new_n1139__));
  and1  g0596(.dina(new_new_n831__), .dinb(new_new_n833__), .dout(new_new_n1140__));
  or1   g0597(.dina(new_new_n830__), .dinb(new_new_n832__), .dout(new_new_n1141__));
  or1   g0598(.dina(new_new_n1126__), .dinb(new_new_n1853__), .dout(new_new_n1142__));
  or1   g0599(.dina(new_new_n1855__), .dinb(new_new_n1132__), .dout(new_new_n1143__));
  or1   g0600(.dina(new_new_n1857__), .dinb(new_new_n1859__), .dout(new_new_n1144__));
  and1  g0601(.dina(new_new_n1857__), .dinb(new_new_n1859__), .dout(new_new_n1145__));
  or1   g0602(.dina(new_new_n1861__), .dinb(new_new_n1863__), .dout(new_new_n1146__));
  or1   g0603(.dina(new_new_n1865__), .dinb(new_new_n1867__), .dout(new_new_n1147__));
  or1   g0604(.dina(new_new_n1869__), .dinb(new_new_n1870__), .dout(new_new_n1148__));
  or1   g0605(.dina(new_new_n1869__), .dinb(new_new_n1872__), .dout(new_new_n1149__));
  or1   g0606(.dina(new_new_n1128__), .dinb(new_new_n1873__), .dout(new_new_n1150__));
  or1   g0607(.dina(new_new_n1872__), .dinb(new_new_n1874__), .dout(new_new_n1151__));
  and1  g0608(.dina(new_new_n1865__), .dinb(new_new_n1867__), .dout(new_new_n1152__));
  or1   g0609(.dina(new_new_n1876__), .dinb(new_new_n1878__), .dout(new_new_n1153__));
  or1   g0610(.dina(new_new_n1130__), .dinb(new_new_n1873__), .dout(new_new_n1154__));
  and1  g0611(.dina(new_new_n1879__), .dinb(new_new_n1154__), .dout(new_new_n1155__));
  or1   g0612(.dina(new_new_n1853__), .dinb(new_new_n1155__), .dout(new_new_n1156__));
  and1  g0613(.dina(new_new_n1880__), .dinb(new_new_n1881__), .dout(new_new_n1157__));
  or1   g0614(.dina(new_new_n1855__), .dinb(new_new_n1157__), .dout(new_new_n1158__));
  and1  g0615(.dina(new_new_n1861__), .dinb(new_new_n1864__), .dout(new_new_n1159__));
  and1  g0616(.dina(new_new_n1856__), .dinb(new_new_n1876__), .dout(new_new_n1160__));
  and1  g0617(.dina(new_new_n1878__), .dinb(new_new_n1858__), .dout(new_new_n1161__));
  and1  g0618(.dina(new_new_n1866__), .dinb(new_new_n1863__), .dout(new_new_n1162__));
  and1  g0619(.dina(new_new_n1882__), .dinb(new_new_n1883__), .dout(new_new_n1163__));
  or1   g0620(.dina(new_new_n1884__), .dinb(new_new_n1163__), .dout(new_new_n1164__));
  and1  g0621(.dina(new_new_n1145__), .dinb(new_new_n1885__), .dout(new_new_n1165__));
  or1   g0622(.dina(new_new_n1152__), .dinb(new_new_n1165__), .dout(new_new_n1166__));
  and1  g0623(.dina(new_new_n1164__), .dinb(new_new_n1166__), .dout(new_new_n1167__));
  and1  g0624(.dina(new_new_n1887__), .dinb(new_new_n1888__), .dout(new_new_n1168__));
  or1   g0625(.dina(new_new_n1889__), .dinb(new_new_n1891__), .dout(new_new_n1169__));
  and1  g0626(.dina(new_new_n1889__), .dinb(new_new_n1891__), .dout(new_new_n1170__));
  or1   g0627(.dina(new_new_n1887__), .dinb(new_new_n1888__), .dout(new_new_n1171__));
  and1  g0628(.dina(new_new_n1169__), .dinb(new_new_n1171__), .dout(new_new_n1172__));
  or1   g0629(.dina(new_new_n1168__), .dinb(new_new_n1170__), .dout(new_new_n1173__));
  and1  g0630(.dina(new_new_n1893__), .dinb(new_new_n1894__), .dout(new_new_n1174__));
  or1   g0631(.dina(new_new_n1895__), .dinb(new_new_n1897__), .dout(new_new_n1175__));
  and1  g0632(.dina(new_new_n1895__), .dinb(new_new_n1897__), .dout(new_new_n1176__));
  or1   g0633(.dina(new_new_n1893__), .dinb(new_new_n1894__), .dout(new_new_n1177__));
  and1  g0634(.dina(new_new_n1175__), .dinb(new_new_n1177__), .dout(new_new_n1178__));
  or1   g0635(.dina(new_new_n1174__), .dinb(new_new_n1176__), .dout(new_new_n1179__));
  and1  g0636(.dina(new_new_n1172__), .dinb(new_new_n1179__), .dout(new_new_n1180__));
  and1  g0637(.dina(new_new_n1173__), .dinb(new_new_n1178__), .dout(new_new_n1181__));
  or1   g0638(.dina(new_new_n1180__), .dinb(new_new_n1181__), .dout(new_new_n1182__));
  and1  g0639(.dina(new_new_n834__), .dinb(new_new_n1900__), .dout(new_new_n1183__));
  or1   g0640(.dina(new_new_n835__), .dinb(new_new_n1907__), .dout(new_new_n1184__));
  and1  g0641(.dina(new_new_n1913__), .dinb(new_new_n1916__), .dout(new_new_n1185__));
  or1   g0642(.dina(new_new_n1919__), .dinb(new_new_n1922__), .dout(new_new_n1186__));
  and1  g0643(.dina(new_new_n1919__), .dinb(new_new_n1922__), .dout(new_new_n1187__));
  or1   g0644(.dina(new_new_n1913__), .dinb(new_new_n1916__), .dout(new_new_n1188__));
  and1  g0645(.dina(new_new_n1186__), .dinb(new_new_n1188__), .dout(new_new_n1189__));
  or1   g0646(.dina(new_new_n1185__), .dinb(new_new_n1187__), .dout(new_new_n1190__));
  or1   g0647(.dina(new_new_n1183__), .dinb(new_new_n1189__), .dout(new_new_n1191__));
  or1   g0648(.dina(new_new_n1184__), .dinb(new_new_n1190__), .dout(new_new_n1192__));
  and1  g0649(.dina(new_new_n1191__), .dinb(new_new_n1192__), .dout(new_new_n1193__));
  or1   g0650(.dina(new_new_n1924__), .dinb(new_new_n1925__), .dout(new_new_n1194__));
  and1  g0651(.dina(new_new_n1924__), .dinb(new_new_n1925__), .dout(new_new_n1195__));
  and1  g0652(.dina(new_new_n1927__), .dinb(new_new_n1928__), .dout(new_new_n1196__));
  or1   g0653(.dina(new_new_n1929__), .dinb(new_new_n1931__), .dout(new_new_n1197__));
  and1  g0654(.dina(new_new_n1929__), .dinb(new_new_n1931__), .dout(new_new_n1198__));
  or1   g0655(.dina(new_new_n1927__), .dinb(new_new_n1928__), .dout(new_new_n1199__));
  and1  g0656(.dina(new_new_n1197__), .dinb(new_new_n1199__), .dout(new_new_n1200__));
  or1   g0657(.dina(new_new_n1196__), .dinb(new_new_n1198__), .dout(new_new_n1201__));
  and1  g0658(.dina(new_new_n1933__), .dinb(new_new_n1934__), .dout(new_new_n1202__));
  or1   g0659(.dina(new_new_n1935__), .dinb(new_new_n1937__), .dout(new_new_n1203__));
  and1  g0660(.dina(new_new_n1935__), .dinb(new_new_n1937__), .dout(new_new_n1204__));
  or1   g0661(.dina(new_new_n1933__), .dinb(new_new_n1934__), .dout(new_new_n1205__));
  and1  g0662(.dina(new_new_n1203__), .dinb(new_new_n1205__), .dout(new_new_n1206__));
  or1   g0663(.dina(new_new_n1202__), .dinb(new_new_n1204__), .dout(new_new_n1207__));
  and1  g0664(.dina(new_new_n1200__), .dinb(new_new_n1207__), .dout(new_new_n1208__));
  and1  g0665(.dina(new_new_n1201__), .dinb(new_new_n1206__), .dout(new_new_n1209__));
  or1   g0666(.dina(new_new_n1208__), .dinb(new_new_n1209__), .dout(new_new_n1210__));
  and1  g0667(.dina(new_new_n836__), .dinb(new_new_n1900__), .dout(new_new_n1211__));
  or1   g0668(.dina(new_new_n837__), .dinb(new_new_n1907__), .dout(new_new_n1212__));
  and1  g0669(.dina(new_new_n1939__), .dinb(new_new_n1942__), .dout(new_new_n1213__));
  or1   g0670(.dina(new_new_n1945__), .dinb(new_new_n1948__), .dout(new_new_n1214__));
  and1  g0671(.dina(new_new_n1945__), .dinb(new_new_n1948__), .dout(new_new_n1215__));
  or1   g0672(.dina(new_new_n1939__), .dinb(new_new_n1942__), .dout(new_new_n1216__));
  and1  g0673(.dina(new_new_n1214__), .dinb(new_new_n1216__), .dout(new_new_n1217__));
  or1   g0674(.dina(new_new_n1213__), .dinb(new_new_n1215__), .dout(new_new_n1218__));
  or1   g0675(.dina(new_new_n1211__), .dinb(new_new_n1217__), .dout(new_new_n1219__));
  or1   g0676(.dina(new_new_n1212__), .dinb(new_new_n1218__), .dout(new_new_n1220__));
  and1  g0677(.dina(new_new_n1219__), .dinb(new_new_n1220__), .dout(new_new_n1221__));
  or1   g0678(.dina(new_new_n1950__), .dinb(new_new_n1951__), .dout(new_new_n1222__));
  and1  g0679(.dina(new_new_n1950__), .dinb(new_new_n1951__), .dout(new_new_n1223__));
  and1  g0680(.dina(new_new_n1953__), .dinb(new_new_n1954__), .dout(new_new_n1224__));
  or1   g0681(.dina(new_new_n1955__), .dinb(new_new_n1957__), .dout(new_new_n1225__));
  and1  g0682(.dina(new_new_n1955__), .dinb(new_new_n1957__), .dout(new_new_n1226__));
  or1   g0683(.dina(new_new_n1953__), .dinb(new_new_n1954__), .dout(new_new_n1227__));
  and1  g0684(.dina(new_new_n1225__), .dinb(new_new_n1227__), .dout(new_new_n1228__));
  or1   g0685(.dina(new_new_n1224__), .dinb(new_new_n1226__), .dout(new_new_n1229__));
  and1  g0686(.dina(new_new_n1959__), .dinb(new_new_n1960__), .dout(new_new_n1230__));
  or1   g0687(.dina(new_new_n1961__), .dinb(new_new_n1963__), .dout(new_new_n1231__));
  and1  g0688(.dina(new_new_n1961__), .dinb(new_new_n1963__), .dout(new_new_n1232__));
  or1   g0689(.dina(new_new_n1959__), .dinb(new_new_n1960__), .dout(new_new_n1233__));
  and1  g0690(.dina(new_new_n1231__), .dinb(new_new_n1233__), .dout(new_new_n1234__));
  or1   g0691(.dina(new_new_n1230__), .dinb(new_new_n1232__), .dout(new_new_n1235__));
  and1  g0692(.dina(new_new_n1228__), .dinb(new_new_n1235__), .dout(new_new_n1236__));
  and1  g0693(.dina(new_new_n1229__), .dinb(new_new_n1234__), .dout(new_new_n1237__));
  or1   g0694(.dina(new_new_n1236__), .dinb(new_new_n1237__), .dout(new_new_n1238__));
  and1  g0695(.dina(new_new_n838__), .dinb(new_new_n1901__), .dout(new_new_n1239__));
  or1   g0696(.dina(new_new_n839__), .dinb(new_new_n1908__), .dout(new_new_n1240__));
  and1  g0697(.dina(new_new_n1914__), .dinb(new_new_n1940__), .dout(new_new_n1241__));
  or1   g0698(.dina(new_new_n1920__), .dinb(new_new_n1946__), .dout(new_new_n1242__));
  and1  g0699(.dina(new_new_n1920__), .dinb(new_new_n1946__), .dout(new_new_n1243__));
  or1   g0700(.dina(new_new_n1914__), .dinb(new_new_n1940__), .dout(new_new_n1244__));
  and1  g0701(.dina(new_new_n1242__), .dinb(new_new_n1244__), .dout(new_new_n1245__));
  or1   g0702(.dina(new_new_n1241__), .dinb(new_new_n1243__), .dout(new_new_n1246__));
  or1   g0703(.dina(new_new_n1239__), .dinb(new_new_n1245__), .dout(new_new_n1247__));
  or1   g0704(.dina(new_new_n1240__), .dinb(new_new_n1246__), .dout(new_new_n1248__));
  and1  g0705(.dina(new_new_n1247__), .dinb(new_new_n1248__), .dout(new_new_n1249__));
  or1   g0706(.dina(new_new_n1964__), .dinb(new_new_n1965__), .dout(new_new_n1250__));
  and1  g0707(.dina(new_new_n1964__), .dinb(new_new_n1965__), .dout(new_new_n1251__));
  and1  g0708(.dina(new_new_n1967__), .dinb(new_new_n1968__), .dout(new_new_n1252__));
  or1   g0709(.dina(new_new_n1969__), .dinb(new_new_n1971__), .dout(new_new_n1253__));
  and1  g0710(.dina(new_new_n1969__), .dinb(new_new_n1971__), .dout(new_new_n1254__));
  or1   g0711(.dina(new_new_n1967__), .dinb(new_new_n1968__), .dout(new_new_n1255__));
  and1  g0712(.dina(new_new_n1253__), .dinb(new_new_n1255__), .dout(new_new_n1256__));
  or1   g0713(.dina(new_new_n1252__), .dinb(new_new_n1254__), .dout(new_new_n1257__));
  and1  g0714(.dina(new_new_n1973__), .dinb(new_new_n1974__), .dout(new_new_n1258__));
  or1   g0715(.dina(new_new_n1975__), .dinb(new_new_n1977__), .dout(new_new_n1259__));
  and1  g0716(.dina(new_new_n1975__), .dinb(new_new_n1977__), .dout(new_new_n1260__));
  or1   g0717(.dina(new_new_n1973__), .dinb(new_new_n1974__), .dout(new_new_n1261__));
  and1  g0718(.dina(new_new_n1259__), .dinb(new_new_n1261__), .dout(new_new_n1262__));
  or1   g0719(.dina(new_new_n1258__), .dinb(new_new_n1260__), .dout(new_new_n1263__));
  and1  g0720(.dina(new_new_n1256__), .dinb(new_new_n1263__), .dout(new_new_n1264__));
  and1  g0721(.dina(new_new_n1257__), .dinb(new_new_n1262__), .dout(new_new_n1265__));
  or1   g0722(.dina(new_new_n1264__), .dinb(new_new_n1265__), .dout(new_new_n1266__));
  and1  g0723(.dina(new_new_n840__), .dinb(new_new_n1901__), .dout(new_new_n1267__));
  or1   g0724(.dina(new_new_n841__), .dinb(new_new_n1908__), .dout(new_new_n1268__));
  and1  g0725(.dina(new_new_n1923__), .dinb(new_new_n1949__), .dout(new_new_n1269__));
  or1   g0726(.dina(new_new_n1917__), .dinb(new_new_n1943__), .dout(new_new_n1270__));
  and1  g0727(.dina(new_new_n1917__), .dinb(new_new_n1943__), .dout(new_new_n1271__));
  or1   g0728(.dina(new_new_n1923__), .dinb(new_new_n1949__), .dout(new_new_n1272__));
  and1  g0729(.dina(new_new_n1270__), .dinb(new_new_n1272__), .dout(new_new_n1273__));
  or1   g0730(.dina(new_new_n1269__), .dinb(new_new_n1271__), .dout(new_new_n1274__));
  or1   g0731(.dina(new_new_n1267__), .dinb(new_new_n1273__), .dout(new_new_n1275__));
  or1   g0732(.dina(new_new_n1268__), .dinb(new_new_n1274__), .dout(new_new_n1276__));
  and1  g0733(.dina(new_new_n1275__), .dinb(new_new_n1276__), .dout(new_new_n1277__));
  or1   g0734(.dina(new_new_n1978__), .dinb(new_new_n1979__), .dout(new_new_n1278__));
  and1  g0735(.dina(new_new_n1978__), .dinb(new_new_n1979__), .dout(new_new_n1279__));
  and1  g0736(.dina(new_new_n1981__), .dinb(new_new_n1982__), .dout(new_new_n1280__));
  or1   g0737(.dina(new_new_n1983__), .dinb(new_new_n1985__), .dout(new_new_n1281__));
  and1  g0738(.dina(new_new_n1983__), .dinb(new_new_n1985__), .dout(new_new_n1282__));
  or1   g0739(.dina(new_new_n1981__), .dinb(new_new_n1982__), .dout(new_new_n1283__));
  and1  g0740(.dina(new_new_n1281__), .dinb(new_new_n1283__), .dout(new_new_n1284__));
  or1   g0741(.dina(new_new_n1280__), .dinb(new_new_n1282__), .dout(new_new_n1285__));
  and1  g0742(.dina(new_new_n1987__), .dinb(new_new_n1988__), .dout(new_new_n1286__));
  or1   g0743(.dina(new_new_n1989__), .dinb(new_new_n1991__), .dout(new_new_n1287__));
  and1  g0744(.dina(new_new_n1989__), .dinb(new_new_n1991__), .dout(new_new_n1288__));
  or1   g0745(.dina(new_new_n1987__), .dinb(new_new_n1988__), .dout(new_new_n1289__));
  and1  g0746(.dina(new_new_n1287__), .dinb(new_new_n1289__), .dout(new_new_n1290__));
  or1   g0747(.dina(new_new_n1286__), .dinb(new_new_n1288__), .dout(new_new_n1291__));
  and1  g0748(.dina(new_new_n1284__), .dinb(new_new_n1291__), .dout(new_new_n1292__));
  and1  g0749(.dina(new_new_n1285__), .dinb(new_new_n1290__), .dout(new_new_n1293__));
  or1   g0750(.dina(new_new_n1292__), .dinb(new_new_n1293__), .dout(new_new_n1294__));
  and1  g0751(.dina(new_new_n842__), .dinb(new_new_n1903__), .dout(new_new_n1295__));
  or1   g0752(.dina(new_new_n843__), .dinb(new_new_n1910__), .dout(new_new_n1296__));
  and1  g0753(.dina(new_new_n1993__), .dinb(new_new_n1996__), .dout(new_new_n1297__));
  or1   g0754(.dina(new_new_n1999__), .dinb(new_new_n2002__), .dout(new_new_n1298__));
  and1  g0755(.dina(new_new_n1999__), .dinb(new_new_n2002__), .dout(new_new_n1299__));
  or1   g0756(.dina(new_new_n1993__), .dinb(new_new_n1996__), .dout(new_new_n1300__));
  and1  g0757(.dina(new_new_n1298__), .dinb(new_new_n1300__), .dout(new_new_n1301__));
  or1   g0758(.dina(new_new_n1297__), .dinb(new_new_n1299__), .dout(new_new_n1302__));
  or1   g0759(.dina(new_new_n1295__), .dinb(new_new_n1301__), .dout(new_new_n1303__));
  or1   g0760(.dina(new_new_n1296__), .dinb(new_new_n1302__), .dout(new_new_n1304__));
  and1  g0761(.dina(new_new_n1303__), .dinb(new_new_n1304__), .dout(new_new_n1305__));
  or1   g0762(.dina(new_new_n2004__), .dinb(new_new_n2005__), .dout(new_new_n1306__));
  and1  g0763(.dina(new_new_n2004__), .dinb(new_new_n2005__), .dout(new_new_n1307__));
  and1  g0764(.dina(new_new_n2007__), .dinb(new_new_n2008__), .dout(new_new_n1308__));
  or1   g0765(.dina(new_new_n2009__), .dinb(new_new_n2011__), .dout(new_new_n1309__));
  and1  g0766(.dina(new_new_n2009__), .dinb(new_new_n2011__), .dout(new_new_n1310__));
  or1   g0767(.dina(new_new_n2007__), .dinb(new_new_n2008__), .dout(new_new_n1311__));
  and1  g0768(.dina(new_new_n1309__), .dinb(new_new_n1311__), .dout(new_new_n1312__));
  or1   g0769(.dina(new_new_n1308__), .dinb(new_new_n1310__), .dout(new_new_n1313__));
  and1  g0770(.dina(new_new_n2013__), .dinb(new_new_n2014__), .dout(new_new_n1314__));
  or1   g0771(.dina(new_new_n2015__), .dinb(new_new_n2017__), .dout(new_new_n1315__));
  and1  g0772(.dina(new_new_n2015__), .dinb(new_new_n2017__), .dout(new_new_n1316__));
  or1   g0773(.dina(new_new_n2013__), .dinb(new_new_n2014__), .dout(new_new_n1317__));
  and1  g0774(.dina(new_new_n1315__), .dinb(new_new_n1317__), .dout(new_new_n1318__));
  or1   g0775(.dina(new_new_n1314__), .dinb(new_new_n1316__), .dout(new_new_n1319__));
  and1  g0776(.dina(new_new_n1312__), .dinb(new_new_n1319__), .dout(new_new_n1320__));
  and1  g0777(.dina(new_new_n1313__), .dinb(new_new_n1318__), .dout(new_new_n1321__));
  or1   g0778(.dina(new_new_n1320__), .dinb(new_new_n1321__), .dout(new_new_n1322__));
  and1  g0779(.dina(new_new_n844__), .dinb(new_new_n1903__), .dout(new_new_n1323__));
  or1   g0780(.dina(new_new_n845__), .dinb(new_new_n1910__), .dout(new_new_n1324__));
  and1  g0781(.dina(new_new_n2019__), .dinb(new_new_n2022__), .dout(new_new_n1325__));
  or1   g0782(.dina(new_new_n2025__), .dinb(new_new_n2028__), .dout(new_new_n1326__));
  and1  g0783(.dina(new_new_n2025__), .dinb(new_new_n2028__), .dout(new_new_n1327__));
  or1   g0784(.dina(new_new_n2019__), .dinb(new_new_n2022__), .dout(new_new_n1328__));
  and1  g0785(.dina(new_new_n1326__), .dinb(new_new_n1328__), .dout(new_new_n1329__));
  or1   g0786(.dina(new_new_n1325__), .dinb(new_new_n1327__), .dout(new_new_n1330__));
  or1   g0787(.dina(new_new_n1323__), .dinb(new_new_n1329__), .dout(new_new_n1331__));
  or1   g0788(.dina(new_new_n1324__), .dinb(new_new_n1330__), .dout(new_new_n1332__));
  and1  g0789(.dina(new_new_n1331__), .dinb(new_new_n1332__), .dout(new_new_n1333__));
  or1   g0790(.dina(new_new_n2030__), .dinb(new_new_n2031__), .dout(new_new_n1334__));
  and1  g0791(.dina(new_new_n2030__), .dinb(new_new_n2031__), .dout(new_new_n1335__));
  and1  g0792(.dina(new_new_n2033__), .dinb(new_new_n2034__), .dout(new_new_n1336__));
  or1   g0793(.dina(new_new_n2035__), .dinb(new_new_n2037__), .dout(new_new_n1337__));
  and1  g0794(.dina(new_new_n2035__), .dinb(new_new_n2037__), .dout(new_new_n1338__));
  or1   g0795(.dina(new_new_n2033__), .dinb(new_new_n2034__), .dout(new_new_n1339__));
  and1  g0796(.dina(new_new_n1337__), .dinb(new_new_n1339__), .dout(new_new_n1340__));
  or1   g0797(.dina(new_new_n1336__), .dinb(new_new_n1338__), .dout(new_new_n1341__));
  and1  g0798(.dina(new_new_n2039__), .dinb(new_new_n2040__), .dout(new_new_n1342__));
  or1   g0799(.dina(new_new_n2041__), .dinb(new_new_n2043__), .dout(new_new_n1343__));
  and1  g0800(.dina(new_new_n2041__), .dinb(new_new_n2043__), .dout(new_new_n1344__));
  or1   g0801(.dina(new_new_n2039__), .dinb(new_new_n2040__), .dout(new_new_n1345__));
  and1  g0802(.dina(new_new_n1343__), .dinb(new_new_n1345__), .dout(new_new_n1346__));
  or1   g0803(.dina(new_new_n1342__), .dinb(new_new_n1344__), .dout(new_new_n1347__));
  and1  g0804(.dina(new_new_n1340__), .dinb(new_new_n1347__), .dout(new_new_n1348__));
  and1  g0805(.dina(new_new_n1341__), .dinb(new_new_n1346__), .dout(new_new_n1349__));
  or1   g0806(.dina(new_new_n1348__), .dinb(new_new_n1349__), .dout(new_new_n1350__));
  and1  g0807(.dina(new_new_n846__), .dinb(new_new_n1904__), .dout(new_new_n1351__));
  or1   g0808(.dina(new_new_n847__), .dinb(new_new_n1911__), .dout(new_new_n1352__));
  and1  g0809(.dina(new_new_n1994__), .dinb(new_new_n2026__), .dout(new_new_n1353__));
  or1   g0810(.dina(new_new_n2000__), .dinb(new_new_n2020__), .dout(new_new_n1354__));
  and1  g0811(.dina(new_new_n2000__), .dinb(new_new_n2020__), .dout(new_new_n1355__));
  or1   g0812(.dina(new_new_n1994__), .dinb(new_new_n2026__), .dout(new_new_n1356__));
  and1  g0813(.dina(new_new_n1354__), .dinb(new_new_n1356__), .dout(new_new_n1357__));
  or1   g0814(.dina(new_new_n1353__), .dinb(new_new_n1355__), .dout(new_new_n1358__));
  or1   g0815(.dina(new_new_n1351__), .dinb(new_new_n1357__), .dout(new_new_n1359__));
  or1   g0816(.dina(new_new_n1352__), .dinb(new_new_n1358__), .dout(new_new_n1360__));
  and1  g0817(.dina(new_new_n1359__), .dinb(new_new_n1360__), .dout(new_new_n1361__));
  or1   g0818(.dina(new_new_n2044__), .dinb(new_new_n2045__), .dout(new_new_n1362__));
  and1  g0819(.dina(new_new_n2044__), .dinb(new_new_n2045__), .dout(new_new_n1363__));
  and1  g0820(.dina(new_new_n2047__), .dinb(new_new_n2048__), .dout(new_new_n1364__));
  or1   g0821(.dina(new_new_n2049__), .dinb(new_new_n2051__), .dout(new_new_n1365__));
  and1  g0822(.dina(new_new_n2049__), .dinb(new_new_n2051__), .dout(new_new_n1366__));
  or1   g0823(.dina(new_new_n2047__), .dinb(new_new_n2048__), .dout(new_new_n1367__));
  and1  g0824(.dina(new_new_n1365__), .dinb(new_new_n1367__), .dout(new_new_n1368__));
  or1   g0825(.dina(new_new_n1364__), .dinb(new_new_n1366__), .dout(new_new_n1369__));
  and1  g0826(.dina(new_new_n2053__), .dinb(new_new_n2054__), .dout(new_new_n1370__));
  or1   g0827(.dina(new_new_n2055__), .dinb(new_new_n2057__), .dout(new_new_n1371__));
  and1  g0828(.dina(new_new_n2055__), .dinb(new_new_n2057__), .dout(new_new_n1372__));
  or1   g0829(.dina(new_new_n2053__), .dinb(new_new_n2054__), .dout(new_new_n1373__));
  and1  g0830(.dina(new_new_n1371__), .dinb(new_new_n1373__), .dout(new_new_n1374__));
  or1   g0831(.dina(new_new_n1370__), .dinb(new_new_n1372__), .dout(new_new_n1375__));
  and1  g0832(.dina(new_new_n1368__), .dinb(new_new_n1375__), .dout(new_new_n1376__));
  and1  g0833(.dina(new_new_n1369__), .dinb(new_new_n1374__), .dout(new_new_n1377__));
  or1   g0834(.dina(new_new_n1376__), .dinb(new_new_n1377__), .dout(new_new_n1378__));
  and1  g0835(.dina(new_new_n848__), .dinb(new_new_n1904__), .dout(new_new_n1379__));
  or1   g0836(.dina(new_new_n849__), .dinb(new_new_n1911__), .dout(new_new_n1380__));
  and1  g0837(.dina(new_new_n2003__), .dinb(new_new_n2023__), .dout(new_new_n1381__));
  or1   g0838(.dina(new_new_n1997__), .dinb(new_new_n2029__), .dout(new_new_n1382__));
  and1  g0839(.dina(new_new_n1997__), .dinb(new_new_n2029__), .dout(new_new_n1383__));
  or1   g0840(.dina(new_new_n2003__), .dinb(new_new_n2023__), .dout(new_new_n1384__));
  and1  g0841(.dina(new_new_n1382__), .dinb(new_new_n1384__), .dout(new_new_n1385__));
  or1   g0842(.dina(new_new_n1381__), .dinb(new_new_n1383__), .dout(new_new_n1386__));
  or1   g0843(.dina(new_new_n1379__), .dinb(new_new_n1385__), .dout(new_new_n1387__));
  or1   g0844(.dina(new_new_n1380__), .dinb(new_new_n1386__), .dout(new_new_n1388__));
  and1  g0845(.dina(new_new_n1387__), .dinb(new_new_n1388__), .dout(new_new_n1389__));
  or1   g0846(.dina(new_new_n2058__), .dinb(new_new_n2059__), .dout(new_new_n1390__));
  and1  g0847(.dina(new_new_n2058__), .dinb(new_new_n2059__), .dout(new_new_n1391__));
  and1  g0848(.dina(new_new_n2061__), .dinb(new_new_n2062__), .dout(new_new_n1392__));
  or1   g0849(.dina(new_new_n2063__), .dinb(new_new_n2065__), .dout(new_new_n1393__));
  and1  g0850(.dina(new_new_n2063__), .dinb(new_new_n2065__), .dout(new_new_n1394__));
  or1   g0851(.dina(new_new_n2061__), .dinb(new_new_n2062__), .dout(new_new_n1395__));
  and1  g0852(.dina(new_new_n1393__), .dinb(new_new_n1395__), .dout(new_new_n1396__));
  or1   g0853(.dina(new_new_n1392__), .dinb(new_new_n1394__), .dout(new_new_n1397__));
  and1  g0854(.dina(new_new_n2067__), .dinb(new_new_n2068__), .dout(new_new_n1398__));
  or1   g0855(.dina(new_new_n2069__), .dinb(new_new_n2071__), .dout(new_new_n1399__));
  and1  g0856(.dina(new_new_n2069__), .dinb(new_new_n2071__), .dout(new_new_n1400__));
  or1   g0857(.dina(new_new_n2067__), .dinb(new_new_n2068__), .dout(new_new_n1401__));
  and1  g0858(.dina(new_new_n1399__), .dinb(new_new_n1401__), .dout(new_new_n1402__));
  or1   g0859(.dina(new_new_n1398__), .dinb(new_new_n1400__), .dout(new_new_n1403__));
  and1  g0860(.dina(new_new_n1396__), .dinb(new_new_n1403__), .dout(new_new_n1404__));
  and1  g0861(.dina(new_new_n1397__), .dinb(new_new_n1402__), .dout(new_new_n1405__));
  or1   g0862(.dina(new_new_n1404__), .dinb(new_new_n1405__), .dout(new_new_n1406__));
  and1  g0863(.dina(new_new_n2073__), .dinb(new_new_n2074__), .dout(new_new_n1407__));
  or1   g0864(.dina(new_new_n2075__), .dinb(new_new_n2077__), .dout(new_new_n1408__));
  and1  g0865(.dina(new_new_n2075__), .dinb(new_new_n2077__), .dout(new_new_n1409__));
  or1   g0866(.dina(new_new_n2073__), .dinb(new_new_n2074__), .dout(new_new_n1410__));
  and1  g0867(.dina(new_new_n1408__), .dinb(new_new_n1410__), .dout(new_new_n1411__));
  or1   g0868(.dina(new_new_n1407__), .dinb(new_new_n1409__), .dout(new_new_n1412__));
  and1  g0869(.dina(new_new_n2079__), .dinb(new_new_n2080__), .dout(new_new_n1413__));
  or1   g0870(.dina(new_new_n2081__), .dinb(new_new_n2083__), .dout(new_new_n1414__));
  and1  g0871(.dina(new_new_n2081__), .dinb(new_new_n2083__), .dout(new_new_n1415__));
  or1   g0872(.dina(new_new_n2079__), .dinb(new_new_n2080__), .dout(new_new_n1416__));
  and1  g0873(.dina(new_new_n1414__), .dinb(new_new_n1416__), .dout(new_new_n1417__));
  or1   g0874(.dina(new_new_n1413__), .dinb(new_new_n1415__), .dout(new_new_n1418__));
  and1  g0875(.dina(new_new_n1411__), .dinb(new_new_n1418__), .dout(new_new_n1419__));
  and1  g0876(.dina(new_new_n1412__), .dinb(new_new_n1417__), .dout(new_new_n1420__));
  or1   g0877(.dina(new_new_n1419__), .dinb(new_new_n1420__), .dout(new_new_n1421__));
  and1  g0878(.dina(new_new_n2085__), .dinb(new_new_n2086__), .dout(new_new_n1422__));
  or1   g0879(.dina(new_new_n2087__), .dinb(new_new_n2089__), .dout(new_new_n1423__));
  and1  g0880(.dina(new_new_n2087__), .dinb(new_new_n2089__), .dout(new_new_n1424__));
  or1   g0881(.dina(new_new_n2085__), .dinb(new_new_n2086__), .dout(new_new_n1425__));
  and1  g0882(.dina(new_new_n1423__), .dinb(new_new_n1425__), .dout(new_new_n1426__));
  or1   g0883(.dina(new_new_n1422__), .dinb(new_new_n1424__), .dout(new_new_n1427__));
  and1  g0884(.dina(new_new_n2091__), .dinb(new_new_n2092__), .dout(new_new_n1428__));
  or1   g0885(.dina(new_new_n2093__), .dinb(new_new_n2095__), .dout(new_new_n1429__));
  and1  g0886(.dina(new_new_n2093__), .dinb(new_new_n2095__), .dout(new_new_n1430__));
  or1   g0887(.dina(new_new_n2091__), .dinb(new_new_n2092__), .dout(new_new_n1431__));
  and1  g0888(.dina(new_new_n1429__), .dinb(new_new_n1431__), .dout(new_new_n1432__));
  or1   g0889(.dina(new_new_n1428__), .dinb(new_new_n1430__), .dout(new_new_n1433__));
  and1  g0890(.dina(new_new_n1426__), .dinb(new_new_n1433__), .dout(new_new_n1434__));
  and1  g0891(.dina(new_new_n1427__), .dinb(new_new_n1432__), .dout(new_new_n1435__));
  or1   g0892(.dina(new_new_n1434__), .dinb(new_new_n1435__), .dout(new_new_n1436__));
  and1  g0893(.dina(new_new_n2097__), .dinb(new_new_n2098__), .dout(new_new_n1437__));
  or1   g0894(.dina(new_new_n2099__), .dinb(new_new_n2101__), .dout(new_new_n1438__));
  and1  g0895(.dina(new_new_n2099__), .dinb(new_new_n2101__), .dout(new_new_n1439__));
  or1   g0896(.dina(new_new_n2097__), .dinb(new_new_n2098__), .dout(new_new_n1440__));
  and1  g0897(.dina(new_new_n1438__), .dinb(new_new_n1440__), .dout(new_new_n1441__));
  or1   g0898(.dina(new_new_n1437__), .dinb(new_new_n1439__), .dout(new_new_n1442__));
  and1  g0899(.dina(new_new_n2103__), .dinb(new_new_n2104__), .dout(new_new_n1443__));
  or1   g0900(.dina(new_new_n2105__), .dinb(new_new_n2107__), .dout(new_new_n1444__));
  and1  g0901(.dina(new_new_n2105__), .dinb(new_new_n2107__), .dout(new_new_n1445__));
  or1   g0902(.dina(new_new_n2103__), .dinb(new_new_n2104__), .dout(new_new_n1446__));
  and1  g0903(.dina(new_new_n1444__), .dinb(new_new_n1446__), .dout(new_new_n1447__));
  or1   g0904(.dina(new_new_n1443__), .dinb(new_new_n1445__), .dout(new_new_n1448__));
  and1  g0905(.dina(new_new_n1441__), .dinb(new_new_n1448__), .dout(new_new_n1449__));
  and1  g0906(.dina(new_new_n1442__), .dinb(new_new_n1447__), .dout(new_new_n1450__));
  or1   g0907(.dina(new_new_n1449__), .dinb(new_new_n1450__), .dout(new_new_n1451__));
  and1  g0908(.dina(new_new_n2109__), .dinb(new_new_n2110__), .dout(new_new_n1452__));
  or1   g0909(.dina(new_new_n2111__), .dinb(new_new_n2113__), .dout(new_new_n1453__));
  and1  g0910(.dina(new_new_n2111__), .dinb(new_new_n2113__), .dout(new_new_n1454__));
  or1   g0911(.dina(new_new_n2109__), .dinb(new_new_n2110__), .dout(new_new_n1455__));
  and1  g0912(.dina(new_new_n1453__), .dinb(new_new_n1455__), .dout(new_new_n1456__));
  or1   g0913(.dina(new_new_n1452__), .dinb(new_new_n1454__), .dout(new_new_n1457__));
  and1  g0914(.dina(new_new_n2115__), .dinb(new_new_n2116__), .dout(new_new_n1458__));
  or1   g0915(.dina(new_new_n2117__), .dinb(new_new_n2119__), .dout(new_new_n1459__));
  and1  g0916(.dina(new_new_n2117__), .dinb(new_new_n2119__), .dout(new_new_n1460__));
  or1   g0917(.dina(new_new_n2115__), .dinb(new_new_n2116__), .dout(new_new_n1461__));
  and1  g0918(.dina(new_new_n1459__), .dinb(new_new_n1461__), .dout(new_new_n1462__));
  or1   g0919(.dina(new_new_n1458__), .dinb(new_new_n1460__), .dout(new_new_n1463__));
  and1  g0920(.dina(new_new_n1456__), .dinb(new_new_n1463__), .dout(new_new_n1464__));
  and1  g0921(.dina(new_new_n1457__), .dinb(new_new_n1462__), .dout(new_new_n1465__));
  or1   g0922(.dina(new_new_n1464__), .dinb(new_new_n1465__), .dout(new_new_n1466__));
  and1  g0923(.dina(new_new_n2121__), .dinb(new_new_n2122__), .dout(new_new_n1467__));
  or1   g0924(.dina(new_new_n2123__), .dinb(new_new_n2125__), .dout(new_new_n1468__));
  and1  g0925(.dina(new_new_n2123__), .dinb(new_new_n2125__), .dout(new_new_n1469__));
  or1   g0926(.dina(new_new_n2121__), .dinb(new_new_n2122__), .dout(new_new_n1470__));
  and1  g0927(.dina(new_new_n1468__), .dinb(new_new_n1470__), .dout(new_new_n1471__));
  or1   g0928(.dina(new_new_n1467__), .dinb(new_new_n1469__), .dout(new_new_n1472__));
  and1  g0929(.dina(new_new_n2127__), .dinb(new_new_n2128__), .dout(new_new_n1473__));
  or1   g0930(.dina(new_new_n2129__), .dinb(new_new_n2131__), .dout(new_new_n1474__));
  and1  g0931(.dina(new_new_n2129__), .dinb(new_new_n2131__), .dout(new_new_n1475__));
  or1   g0932(.dina(new_new_n2127__), .dinb(new_new_n2128__), .dout(new_new_n1476__));
  and1  g0933(.dina(new_new_n1474__), .dinb(new_new_n1476__), .dout(new_new_n1477__));
  or1   g0934(.dina(new_new_n1473__), .dinb(new_new_n1475__), .dout(new_new_n1478__));
  and1  g0935(.dina(new_new_n1471__), .dinb(new_new_n1478__), .dout(new_new_n1479__));
  and1  g0936(.dina(new_new_n1472__), .dinb(new_new_n1477__), .dout(new_new_n1480__));
  or1   g0937(.dina(new_new_n1479__), .dinb(new_new_n1480__), .dout(new_new_n1481__));
  and1  g0938(.dina(new_new_n2133__), .dinb(new_new_n2134__), .dout(new_new_n1482__));
  or1   g0939(.dina(new_new_n2135__), .dinb(new_new_n2137__), .dout(new_new_n1483__));
  and1  g0940(.dina(new_new_n2135__), .dinb(new_new_n2137__), .dout(new_new_n1484__));
  or1   g0941(.dina(new_new_n2133__), .dinb(new_new_n2134__), .dout(new_new_n1485__));
  and1  g0942(.dina(new_new_n1483__), .dinb(new_new_n1485__), .dout(new_new_n1486__));
  or1   g0943(.dina(new_new_n1482__), .dinb(new_new_n1484__), .dout(new_new_n1487__));
  and1  g0944(.dina(new_new_n2139__), .dinb(new_new_n2140__), .dout(new_new_n1488__));
  or1   g0945(.dina(new_new_n2141__), .dinb(new_new_n2143__), .dout(new_new_n1489__));
  and1  g0946(.dina(new_new_n2141__), .dinb(new_new_n2143__), .dout(new_new_n1490__));
  or1   g0947(.dina(new_new_n2139__), .dinb(new_new_n2140__), .dout(new_new_n1491__));
  and1  g0948(.dina(new_new_n1489__), .dinb(new_new_n1491__), .dout(new_new_n1492__));
  or1   g0949(.dina(new_new_n1488__), .dinb(new_new_n1490__), .dout(new_new_n1493__));
  and1  g0950(.dina(new_new_n1486__), .dinb(new_new_n1493__), .dout(new_new_n1494__));
  and1  g0951(.dina(new_new_n1487__), .dinb(new_new_n1492__), .dout(new_new_n1495__));
  or1   g0952(.dina(new_new_n1494__), .dinb(new_new_n1495__), .dout(new_new_n1496__));
  and1  g0953(.dina(new_new_n2145__), .dinb(new_new_n2146__), .dout(new_new_n1497__));
  or1   g0954(.dina(new_new_n2147__), .dinb(new_new_n2149__), .dout(new_new_n1498__));
  and1  g0955(.dina(new_new_n2147__), .dinb(new_new_n2149__), .dout(new_new_n1499__));
  or1   g0956(.dina(new_new_n2145__), .dinb(new_new_n2146__), .dout(new_new_n1500__));
  and1  g0957(.dina(new_new_n1498__), .dinb(new_new_n1500__), .dout(new_new_n1501__));
  or1   g0958(.dina(new_new_n1497__), .dinb(new_new_n1499__), .dout(new_new_n1502__));
  and1  g0959(.dina(new_new_n2151__), .dinb(new_new_n2152__), .dout(new_new_n1503__));
  or1   g0960(.dina(new_new_n2153__), .dinb(new_new_n2155__), .dout(new_new_n1504__));
  and1  g0961(.dina(new_new_n2153__), .dinb(new_new_n2155__), .dout(new_new_n1505__));
  or1   g0962(.dina(new_new_n2151__), .dinb(new_new_n2152__), .dout(new_new_n1506__));
  and1  g0963(.dina(new_new_n1504__), .dinb(new_new_n1506__), .dout(new_new_n1507__));
  or1   g0964(.dina(new_new_n1503__), .dinb(new_new_n1505__), .dout(new_new_n1508__));
  and1  g0965(.dina(new_new_n1501__), .dinb(new_new_n1508__), .dout(new_new_n1509__));
  and1  g0966(.dina(new_new_n1502__), .dinb(new_new_n1507__), .dout(new_new_n1510__));
  or1   g0967(.dina(new_new_n1509__), .dinb(new_new_n1510__), .dout(new_new_n1511__));
  buf1  g0968(.din(new_new_n942__), .dout(G468));
  buf1  g0969(.din(new_new_n947__), .dout(G469));
  buf1  g0970(.din(new_new_n952__), .dout(G470));
  buf1  g0971(.din(new_new_n957__), .dout(G471));
  buf1  g0972(.din(new_new_n966__), .dout(G472));
  buf1  g0973(.din(new_new_n971__), .dout(G473));
  buf1  g0974(.din(new_new_n976__), .dout(G474));
  buf1  g0975(.din(new_new_n981__), .dout(G475));
  buf1  g0976(.din(new_new_n990__), .dout(G476));
  buf1  g0977(.din(new_new_n995__), .dout(G477));
  buf1  g0978(.din(new_new_n1000__), .dout(G478));
  buf1  g0979(.din(new_new_n1005__), .dout(G479));
  buf1  g0980(.din(new_new_n1014__), .dout(G480));
  buf1  g0981(.din(new_new_n1019__), .dout(G481));
  buf1  g0982(.din(new_new_n1024__), .dout(G482));
  buf1  g0983(.din(new_new_n1029__), .dout(G483));
  buf1  g0984(.din(new_new_n1038__), .dout(G484));
  buf1  g0985(.din(new_new_n1043__), .dout(G485));
  buf1  g0986(.din(new_new_n1048__), .dout(G486));
  buf1  g0987(.din(new_new_n1053__), .dout(G487));
  buf1  g0988(.din(new_new_n1062__), .dout(G488));
  buf1  g0989(.din(new_new_n1067__), .dout(G489));
  buf1  g0990(.din(new_new_n1072__), .dout(G490));
  buf1  g0991(.din(new_new_n1077__), .dout(G491));
  buf1  g0992(.din(new_new_n1086__), .dout(G492));
  buf1  g0993(.din(new_new_n1091__), .dout(G493));
  buf1  g0994(.din(new_new_n1096__), .dout(G494));
  buf1  g0995(.din(new_new_n1101__), .dout(G495));
  buf1  g0996(.din(new_new_n1110__), .dout(G496));
  buf1  g0997(.din(new_new_n1115__), .dout(G497));
  buf1  g0998(.din(new_new_n1120__), .dout(G498));
  buf1  g0999(.din(new_new_n1125__), .dout(G499));
  buf1  g1000(.din(new_new_n626__), .dout(n3533));
  buf1  g1001(.din(new_new_n628__), .dout(n3536));
  buf1  g1002(.din(new_new_n630__), .dout(n3539));
  buf1  g1003(.din(new_new_n632__), .dout(n3542));
  buf1  g1004(.din(new_new_n634__), .dout(n3545));
  buf1  g1005(.din(new_new_n636__), .dout(n3548));
  buf1  g1006(.din(new_new_n638__), .dout(n3551));
  buf1  g1007(.din(new_new_n640__), .dout(n3554));
  buf1  g1008(.din(new_new_n642__), .dout(n3557));
  buf1  g1009(.din(new_new_n644__), .dout(n3560));
  buf1  g1010(.din(new_new_n646__), .dout(n3563));
  buf1  g1011(.din(new_new_n648__), .dout(n3566));
  buf1  g1012(.din(new_new_n650__), .dout(n3569));
  buf1  g1013(.din(new_new_n652__), .dout(n3572));
  buf1  g1014(.din(new_new_n654__), .dout(n3575));
  buf1  g1015(.din(new_new_n656__), .dout(n3578));
  buf1  g1016(.din(new_new_n658__), .dout(n3581));
  buf1  g1017(.din(new_new_n660__), .dout(n3584));
  buf1  g1018(.din(new_new_n662__), .dout(n3587));
  buf1  g1019(.din(new_new_n664__), .dout(n3590));
  buf1  g1020(.din(new_new_n666__), .dout(n3593));
  buf1  g1021(.din(new_new_n668__), .dout(n3596));
  buf1  g1022(.din(new_new_n670__), .dout(n3599));
  buf1  g1023(.din(new_new_n672__), .dout(n3602));
  buf1  g1024(.din(new_new_n674__), .dout(n3605));
  buf1  g1025(.din(new_new_n676__), .dout(n3608));
  buf1  g1026(.din(new_new_n678__), .dout(n3611));
  buf1  g1027(.din(new_new_n680__), .dout(n3614));
  buf1  g1028(.din(new_new_n682__), .dout(n3617));
  buf1  g1029(.din(new_new_n684__), .dout(n3620));
  buf1  g1030(.din(new_new_n686__), .dout(n3623));
  buf1  g1031(.din(new_new_n688__), .dout(n3626));
  buf1  g1032(.din(new_new_n526__), .dout(n3629));
  buf1  g1033(.din(new_new_n528__), .dout(n3632));
  buf1  g1034(.din(new_new_n530__), .dout(n3635));
  buf1  g1035(.din(new_new_n532__), .dout(n3638));
  buf1  g1036(.din(new_new_n534__), .dout(n3641));
  buf1  g1037(.din(new_new_n536__), .dout(n3644));
  buf1  g1038(.din(new_new_n538__), .dout(n3647));
  buf1  g1039(.din(new_new_n540__), .dout(n3650));
  buf1  g1040(.din(new_new_n542__), .dout(n3653));
  buf1  g1041(.din(new_new_n1886__), .dout(n3656));
  buf1  g1042(.din(new_new_n1926__), .dout(n3659));
  buf1  g1043(.din(new_new_n1952__), .dout(n3662));
  buf1  g1044(.din(new_new_n1966__), .dout(n3665));
  buf1  g1045(.din(new_new_n1890__), .dout(n3668));
  buf1  g1046(.din(new_new_n1930__), .dout(n3671));
  buf1  g1047(.din(new_new_n1956__), .dout(n3674));
  buf1  g1048(.din(new_new_n1970__), .dout(n3677));
  buf1  g1049(.din(new_new_n1892__), .dout(n3680));
  buf1  g1050(.din(new_new_n1932__), .dout(n3683));
  buf1  g1051(.din(new_new_n1958__), .dout(n3686));
  buf1  g1052(.din(new_new_n1972__), .dout(n3689));
  buf1  g1053(.din(new_new_n1896__), .dout(n3692));
  buf1  g1054(.din(new_new_n1936__), .dout(n3695));
  buf1  g1055(.din(new_new_n1962__), .dout(n3698));
  buf1  g1056(.din(new_new_n1976__), .dout(n3701));
  buf1  g1057(.din(new_new_n1980__), .dout(n3704));
  buf1  g1058(.din(new_new_n2006__), .dout(n3707));
  buf1  g1059(.din(new_new_n2032__), .dout(n3710));
  buf1  g1060(.din(new_new_n2046__), .dout(n3713));
  buf1  g1061(.din(new_new_n1984__), .dout(n3716));
  buf1  g1062(.din(new_new_n2010__), .dout(n3719));
  buf1  g1063(.din(new_new_n2036__), .dout(n3722));
  buf1  g1064(.din(new_new_n2050__), .dout(n3725));
  buf1  g1065(.din(new_new_n1986__), .dout(n3728));
  buf1  g1066(.din(new_new_n2012__), .dout(n3731));
  buf1  g1067(.din(new_new_n2038__), .dout(n3734));
  buf1  g1068(.din(new_new_n2052__), .dout(n3737));
  buf1  g1069(.din(new_new_n1990__), .dout(n3740));
  buf1  g1070(.din(new_new_n2016__), .dout(n3743));
  buf1  g1071(.din(new_new_n2042__), .dout(n3746));
  buf1  g1072(.din(new_new_n2056__), .dout(n3749));
  buf1  g1073(.din(new_new_n1868__), .dout(n3752));
  buf1  g1074(.din(new_new_n1852__), .dout(n3755));
  buf1  g1075(.din(new_new_n1854__), .dout(n3758));
  buf1  g1076(.din(new_new_n1871__), .dout(n3761));
  buf1  g1077(.din(new_new_n1860__), .dout(n3764));
  buf1  g1078(.din(new_new_n1875__), .dout(n3767));
  buf1  g1079(.din(new_new_n1877__), .dout(n3770));
  buf1  g1080(.din(new_new_n1862__), .dout(n3773));
  not1  g1081(.din(new_new_n1874__), .dout(n3776));
  not1  g1082(.din(new_new_n1870__), .dout(n3779));
  not1  g1083(.din(new_new_n1882__), .dout(n3782));
  buf1  g1084(.din(new_new_n1883__), .dout(n3785));
  not1  g1085(.din(new_new_n1885__), .dout(n3788));
  not1  g1086(.din(new_new_n1879__), .dout(n3791));
  not1  g1087(.din(new_new_n1880__), .dout(n3794));
  not1  g1088(.din(new_new_n1881__), .dout(n3797));
  buf1  g1089(.din(new_new_n1884__), .dout(n3800));
  buf1  g1090(.din(new_new_n2060__), .dout(n3803));
  buf1  g1091(.din(new_new_n2064__), .dout(n3806));
  buf1  g1092(.din(new_new_n2066__), .dout(n3809));
  buf1  g1093(.din(new_new_n2070__), .dout(n3812));
  buf1  g1094(.din(new_new_n2072__), .dout(n3815));
  buf1  g1095(.din(new_new_n2076__), .dout(n3818));
  buf1  g1096(.din(new_new_n2078__), .dout(n3821));
  buf1  g1097(.din(new_new_n2082__), .dout(n3824));
  buf1  g1098(.din(new_new_n2084__), .dout(n3827));
  buf1  g1099(.din(new_new_n2088__), .dout(n3830));
  buf1  g1100(.din(new_new_n2090__), .dout(n3833));
  buf1  g1101(.din(new_new_n2094__), .dout(n3836));
  buf1  g1102(.din(new_new_n2096__), .dout(n3839));
  buf1  g1103(.din(new_new_n2100__), .dout(n3842));
  buf1  g1104(.din(new_new_n2102__), .dout(n3845));
  buf1  g1105(.din(new_new_n2106__), .dout(n3848));
  buf1  g1106(.din(new_new_n2108__), .dout(n3851));
  buf1  g1107(.din(new_new_n2112__), .dout(n3854));
  buf1  g1108(.din(new_new_n2114__), .dout(n3857));
  buf1  g1109(.din(new_new_n2118__), .dout(n3860));
  buf1  g1110(.din(new_new_n2120__), .dout(n3863));
  buf1  g1111(.din(new_new_n2124__), .dout(n3866));
  buf1  g1112(.din(new_new_n2126__), .dout(n3869));
  buf1  g1113(.din(new_new_n2130__), .dout(n3872));
  buf1  g1114(.din(new_new_n2132__), .dout(n3875));
  buf1  g1115(.din(new_new_n2136__), .dout(n3878));
  buf1  g1116(.din(new_new_n2138__), .dout(n3881));
  buf1  g1117(.din(new_new_n2142__), .dout(n3884));
  buf1  g1118(.din(new_new_n2144__), .dout(n3887));
  buf1  g1119(.din(new_new_n2148__), .dout(n3890));
  buf1  g1120(.din(new_new_n2150__), .dout(n3893));
  buf1  g1121(.din(new_new_n2154__), .dout(n3896));
  not1  g1122(.din(new_new_n1156__), .dout(n3899));
  not1  g1123(.din(new_new_n1158__), .dout(n3902));
  buf1  g1124(.din(new_new_n1159__), .dout(n3905));
  buf1  g1125(.din(new_new_n1160__), .dout(n3908));
  buf1  g1126(.din(new_new_n1161__), .dout(n3911));
  buf1  g1127(.din(new_new_n1162__), .dout(n3914));
  buf1  g1128(.din(new_new_n1167__), .dout(n3917));
  not1  g1129(.din(new_new_n1194__), .dout(n3920));
  buf1  g1130(.din(new_new_n1195__), .dout(n3923));
  not1  g1131(.din(new_new_n1222__), .dout(n3926));
  buf1  g1132(.din(new_new_n1223__), .dout(n3929));
  not1  g1133(.din(new_new_n1250__), .dout(n3932));
  buf1  g1134(.din(new_new_n1251__), .dout(n3935));
  not1  g1135(.din(new_new_n1278__), .dout(n3938));
  buf1  g1136(.din(new_new_n1279__), .dout(n3941));
  not1  g1137(.din(new_new_n1306__), .dout(n3944));
  buf1  g1138(.din(new_new_n1307__), .dout(n3947));
  not1  g1139(.din(new_new_n1334__), .dout(n3950));
  buf1  g1140(.din(new_new_n1335__), .dout(n3953));
  not1  g1141(.din(new_new_n1362__), .dout(n3956));
  buf1  g1142(.din(new_new_n1363__), .dout(n3959));
  not1  g1143(.din(new_new_n1390__), .dout(n3962));
  buf1  g1144(.din(new_new_n1391__), .dout(n3965));
  buf1  g1145(.din(new_new_n608__), .dout(n3968));
  buf1  g1146(.din(new_new_n610__), .dout(n3971));
  buf1  g1147(.din(new_new_n612__), .dout(n3974));
  buf1  g1148(.din(new_new_n614__), .dout(n3977));
  buf1  g1149(.din(new_new_n616__), .dout(n3980));
  buf1  g1150(.din(new_new_n618__), .dout(n3983));
  buf1  g1151(.din(new_new_n620__), .dout(n3986));
  buf1  g1152(.din(new_new_n622__), .dout(n3989));
  buf1  g1153(.din(new_new_n624__), .dout(n3992));
  buf1  g1154(.din(new_new_n1406__), .dout(n3995));
  buf1  g1155(.din(new_new_n1421__), .dout(n3998));
  buf1  g1156(.din(new_new_n1436__), .dout(n4001));
  buf1  g1157(.din(new_new_n1451__), .dout(n4004));
  buf1  g1158(.din(new_new_n1466__), .dout(n4007));
  buf1  g1159(.din(new_new_n1481__), .dout(n4010));
  buf1  g1160(.din(new_new_n1496__), .dout(n4013));
  buf1  g1161(.din(new_new_n1511__), .dout(n4016));
  buf1  g1162(.din(new_new_n462__), .dout(n4019));
  buf1  g1163(.din(new_new_n464__), .dout(n4022));
  buf1  g1164(.din(new_new_n466__), .dout(n4025));
  buf1  g1165(.din(new_new_n468__), .dout(n4028));
  buf1  g1166(.din(new_new_n470__), .dout(n4031));
  buf1  g1167(.din(new_new_n472__), .dout(n4034));
  buf1  g1168(.din(new_new_n474__), .dout(n4037));
  buf1  g1169(.din(new_new_n476__), .dout(n4040));
  buf1  g1170(.din(new_new_n478__), .dout(n4043));
  buf1  g1171(.din(new_new_n480__), .dout(n4046));
  buf1  g1172(.din(new_new_n482__), .dout(n4049));
  buf1  g1173(.din(new_new_n484__), .dout(n4052));
  buf1  g1174(.din(new_new_n486__), .dout(n4055));
  buf1  g1175(.din(new_new_n488__), .dout(n4058));
  buf1  g1176(.din(new_new_n490__), .dout(n4061));
  buf1  g1177(.din(new_new_n492__), .dout(n4064));
  buf1  g1178(.din(new_new_n494__), .dout(n4067));
  buf1  g1179(.din(new_new_n496__), .dout(n4070));
  buf1  g1180(.din(new_new_n498__), .dout(n4073));
  buf1  g1181(.din(new_new_n500__), .dout(n4076));
  buf1  g1182(.din(new_new_n502__), .dout(n4079));
  buf1  g1183(.din(new_new_n504__), .dout(n4082));
  buf1  g1184(.din(new_new_n506__), .dout(n4085));
  buf1  g1185(.din(new_new_n508__), .dout(n4088));
  buf1  g1186(.din(new_new_n510__), .dout(n4091));
  buf1  g1187(.din(new_new_n512__), .dout(n4094));
  buf1  g1188(.din(new_new_n514__), .dout(n4097));
  buf1  g1189(.din(new_new_n516__), .dout(n4100));
  buf1  g1190(.din(new_new_n518__), .dout(n4103));
  buf1  g1191(.din(new_new_n520__), .dout(n4106));
  buf1  g1192(.din(new_new_n522__), .dout(n4109));
  buf1  g1193(.din(new_new_n524__), .dout(n4112));
  buf1  g1194(.din(new_new_n933__), .dout(new_new_n1738__));
  buf1  g1195(.din(new_new_n1738__), .dout(new_new_n1739__));
  buf1  g1196(.din(new_new_n1738__), .dout(new_new_n1740__));
  buf1  g1197(.din(new_new_n932__), .dout(new_new_n1741__));
  buf1  g1198(.din(new_new_n1741__), .dout(new_new_n1742__));
  buf1  g1199(.din(new_new_n1741__), .dout(new_new_n1743__));
  buf1  g1200(.din(new_new_n690__), .dout(new_new_n1744__));
  buf1  g1201(.din(new_new_n1744__), .dout(new_new_n1745__));
  buf1  g1202(.din(new_new_n1744__), .dout(new_new_n1746__));
  buf1  g1203(.din(new_new_n936__), .dout(new_new_n1747__));
  buf1  g1204(.din(new_new_n1747__), .dout(new_new_n1748__));
  buf1  g1205(.din(new_new_n1747__), .dout(new_new_n1749__));
  buf1  g1206(.din(new_new_n691__), .dout(new_new_n1750__));
  buf1  g1207(.din(new_new_n1750__), .dout(new_new_n1751__));
  buf1  g1208(.din(new_new_n1750__), .dout(new_new_n1752__));
  buf1  g1209(.din(new_new_n937__), .dout(new_new_n1753__));
  buf1  g1210(.din(new_new_n1753__), .dout(new_new_n1754__));
  buf1  g1211(.din(new_new_n1753__), .dout(new_new_n1755__));
  buf1  g1212(.din(new_new_n692__), .dout(new_new_n1756__));
  buf1  g1213(.din(new_new_n1756__), .dout(new_new_n1757__));
  buf1  g1214(.din(new_new_n1757__), .dout(new_new_n1758__));
  buf1  g1215(.din(new_new_n1756__), .dout(new_new_n1759__));
  buf1  g1216(.din(new_new_n693__), .dout(new_new_n1760__));
  buf1  g1217(.din(new_new_n1760__), .dout(new_new_n1761__));
  buf1  g1218(.din(new_new_n1761__), .dout(new_new_n1762__));
  buf1  g1219(.din(new_new_n1760__), .dout(new_new_n1763__));
  buf1  g1220(.din(new_new_n694__), .dout(new_new_n1764__));
  buf1  g1221(.din(new_new_n1764__), .dout(new_new_n1765__));
  buf1  g1222(.din(new_new_n1765__), .dout(new_new_n1766__));
  buf1  g1223(.din(new_new_n1765__), .dout(new_new_n1767__));
  buf1  g1224(.din(new_new_n1764__), .dout(new_new_n1768__));
  buf1  g1225(.din(new_new_n695__), .dout(new_new_n1769__));
  buf1  g1226(.din(new_new_n1769__), .dout(new_new_n1770__));
  buf1  g1227(.din(new_new_n1770__), .dout(new_new_n1771__));
  buf1  g1228(.din(new_new_n1770__), .dout(new_new_n1772__));
  buf1  g1229(.din(new_new_n1769__), .dout(new_new_n1773__));
  buf1  g1230(.din(new_new_n696__), .dout(new_new_n1774__));
  buf1  g1231(.din(new_new_n1774__), .dout(new_new_n1775__));
  buf1  g1232(.din(new_new_n1774__), .dout(new_new_n1776__));
  buf1  g1233(.din(new_new_n697__), .dout(new_new_n1777__));
  buf1  g1234(.din(new_new_n1777__), .dout(new_new_n1778__));
  buf1  g1235(.din(new_new_n1777__), .dout(new_new_n1779__));
  buf1  g1236(.din(new_new_n960__), .dout(new_new_n1780__));
  buf1  g1237(.din(new_new_n1780__), .dout(new_new_n1781__));
  buf1  g1238(.din(new_new_n1780__), .dout(new_new_n1782__));
  buf1  g1239(.din(new_new_n961__), .dout(new_new_n1783__));
  buf1  g1240(.din(new_new_n1783__), .dout(new_new_n1784__));
  buf1  g1241(.din(new_new_n1783__), .dout(new_new_n1785__));
  buf1  g1242(.din(new_new_n984__), .dout(new_new_n1786__));
  buf1  g1243(.din(new_new_n1786__), .dout(new_new_n1787__));
  buf1  g1244(.din(new_new_n1786__), .dout(new_new_n1788__));
  buf1  g1245(.din(new_new_n985__), .dout(new_new_n1789__));
  buf1  g1246(.din(new_new_n1789__), .dout(new_new_n1790__));
  buf1  g1247(.din(new_new_n1789__), .dout(new_new_n1791__));
  buf1  g1248(.din(new_new_n1008__), .dout(new_new_n1792__));
  buf1  g1249(.din(new_new_n1792__), .dout(new_new_n1793__));
  buf1  g1250(.din(new_new_n1792__), .dout(new_new_n1794__));
  buf1  g1251(.din(new_new_n1009__), .dout(new_new_n1795__));
  buf1  g1252(.din(new_new_n1795__), .dout(new_new_n1796__));
  buf1  g1253(.din(new_new_n1795__), .dout(new_new_n1797__));
  buf1  g1254(.din(new_new_n800__), .dout(new_new_n1798__));
  buf1  g1255(.din(new_new_n1798__), .dout(new_new_n1799__));
  buf1  g1256(.din(new_new_n1798__), .dout(new_new_n1800__));
  buf1  g1257(.din(new_new_n801__), .dout(new_new_n1801__));
  buf1  g1258(.din(new_new_n1801__), .dout(new_new_n1802__));
  buf1  g1259(.din(new_new_n1801__), .dout(new_new_n1803__));
  buf1  g1260(.din(new_new_n698__), .dout(new_new_n1804__));
  buf1  g1261(.din(new_new_n1804__), .dout(new_new_n1805__));
  buf1  g1262(.din(new_new_n1804__), .dout(new_new_n1806__));
  buf1  g1263(.din(new_new_n1032__), .dout(new_new_n1807__));
  buf1  g1264(.din(new_new_n1807__), .dout(new_new_n1808__));
  buf1  g1265(.din(new_new_n1807__), .dout(new_new_n1809__));
  buf1  g1266(.din(new_new_n699__), .dout(new_new_n1810__));
  buf1  g1267(.din(new_new_n1810__), .dout(new_new_n1811__));
  buf1  g1268(.din(new_new_n1810__), .dout(new_new_n1812__));
  buf1  g1269(.din(new_new_n1033__), .dout(new_new_n1813__));
  buf1  g1270(.din(new_new_n1813__), .dout(new_new_n1814__));
  buf1  g1271(.din(new_new_n1813__), .dout(new_new_n1815__));
  buf1  g1272(.din(new_new_n700__), .dout(new_new_n1816__));
  buf1  g1273(.din(new_new_n1816__), .dout(new_new_n1817__));
  buf1  g1274(.din(new_new_n1816__), .dout(new_new_n1818__));
  buf1  g1275(.din(new_new_n701__), .dout(new_new_n1819__));
  buf1  g1276(.din(new_new_n1819__), .dout(new_new_n1820__));
  buf1  g1277(.din(new_new_n1819__), .dout(new_new_n1821__));
  buf1  g1278(.din(new_new_n702__), .dout(new_new_n1822__));
  buf1  g1279(.din(new_new_n1822__), .dout(new_new_n1823__));
  buf1  g1280(.din(new_new_n1822__), .dout(new_new_n1824__));
  buf1  g1281(.din(new_new_n703__), .dout(new_new_n1825__));
  buf1  g1282(.din(new_new_n1825__), .dout(new_new_n1826__));
  buf1  g1283(.din(new_new_n1825__), .dout(new_new_n1827__));
  buf1  g1284(.din(new_new_n704__), .dout(new_new_n1828__));
  buf1  g1285(.din(new_new_n1828__), .dout(new_new_n1829__));
  buf1  g1286(.din(new_new_n1828__), .dout(new_new_n1830__));
  buf1  g1287(.din(new_new_n705__), .dout(new_new_n1831__));
  buf1  g1288(.din(new_new_n1831__), .dout(new_new_n1832__));
  buf1  g1289(.din(new_new_n1831__), .dout(new_new_n1833__));
  buf1  g1290(.din(new_new_n1056__), .dout(new_new_n1834__));
  buf1  g1291(.din(new_new_n1834__), .dout(new_new_n1835__));
  buf1  g1292(.din(new_new_n1834__), .dout(new_new_n1836__));
  buf1  g1293(.din(new_new_n1057__), .dout(new_new_n1837__));
  buf1  g1294(.din(new_new_n1837__), .dout(new_new_n1838__));
  buf1  g1295(.din(new_new_n1837__), .dout(new_new_n1839__));
  buf1  g1296(.din(new_new_n1080__), .dout(new_new_n1840__));
  buf1  g1297(.din(new_new_n1840__), .dout(new_new_n1841__));
  buf1  g1298(.din(new_new_n1840__), .dout(new_new_n1842__));
  buf1  g1299(.din(new_new_n1081__), .dout(new_new_n1843__));
  buf1  g1300(.din(new_new_n1843__), .dout(new_new_n1844__));
  buf1  g1301(.din(new_new_n1843__), .dout(new_new_n1845__));
  buf1  g1302(.din(new_new_n1104__), .dout(new_new_n1846__));
  buf1  g1303(.din(new_new_n1846__), .dout(new_new_n1847__));
  buf1  g1304(.din(new_new_n1846__), .dout(new_new_n1848__));
  buf1  g1305(.din(new_new_n1105__), .dout(new_new_n1849__));
  buf1  g1306(.din(new_new_n1849__), .dout(new_new_n1850__));
  buf1  g1307(.din(new_new_n1849__), .dout(new_new_n1851__));
  buf1  g1308(.din(new_new_n1129__), .dout(new_new_n1852__));
  buf1  g1309(.din(new_new_n1852__), .dout(new_new_n1853__));
  buf1  g1310(.din(new_new_n1131__), .dout(new_new_n1854__));
  buf1  g1311(.din(new_new_n1854__), .dout(new_new_n1855__));
  buf1  g1312(.din(new_new_n1134__), .dout(new_new_n1856__));
  buf1  g1313(.din(new_new_n1856__), .dout(new_new_n1857__));
  buf1  g1314(.din(new_new_n1140__), .dout(new_new_n1858__));
  buf1  g1315(.din(new_new_n1858__), .dout(new_new_n1859__));
  buf1  g1316(.din(new_new_n1135__), .dout(new_new_n1860__));
  buf1  g1317(.din(new_new_n1860__), .dout(new_new_n1861__));
  buf1  g1318(.din(new_new_n1141__), .dout(new_new_n1862__));
  buf1  g1319(.din(new_new_n1862__), .dout(new_new_n1863__));
  buf1  g1320(.din(new_new_n1136__), .dout(new_new_n1864__));
  buf1  g1321(.din(new_new_n1864__), .dout(new_new_n1865__));
  buf1  g1322(.din(new_new_n1138__), .dout(new_new_n1866__));
  buf1  g1323(.din(new_new_n1866__), .dout(new_new_n1867__));
  buf1  g1324(.din(new_new_n1127__), .dout(new_new_n1868__));
  buf1  g1325(.din(new_new_n1868__), .dout(new_new_n1869__));
  buf1  g1326(.din(new_new_n1143__), .dout(new_new_n1870__));
  buf1  g1327(.din(new_new_n1133__), .dout(new_new_n1871__));
  buf1  g1328(.din(new_new_n1871__), .dout(new_new_n1872__));
  buf1  g1329(.din(new_new_n1149__), .dout(new_new_n1873__));
  buf1  g1330(.din(new_new_n1142__), .dout(new_new_n1874__));
  buf1  g1331(.din(new_new_n1137__), .dout(new_new_n1875__));
  buf1  g1332(.din(new_new_n1875__), .dout(new_new_n1876__));
  buf1  g1333(.din(new_new_n1139__), .dout(new_new_n1877__));
  buf1  g1334(.din(new_new_n1877__), .dout(new_new_n1878__));
  buf1  g1335(.din(new_new_n1148__), .dout(new_new_n1879__));
  buf1  g1336(.din(new_new_n1150__), .dout(new_new_n1880__));
  buf1  g1337(.din(new_new_n1151__), .dout(new_new_n1881__));
  buf1  g1338(.din(new_new_n1144__), .dout(new_new_n1882__));
  buf1  g1339(.din(new_new_n1146__), .dout(new_new_n1883__));
  buf1  g1340(.din(new_new_n1153__), .dout(new_new_n1884__));
  buf1  g1341(.din(new_new_n1147__), .dout(new_new_n1885__));
  buf1  g1342(.din(new_new_n724__), .dout(new_new_n1886__));
  buf1  g1343(.din(new_new_n1886__), .dout(new_new_n1887__));
  buf1  g1344(.din(new_new_n733__), .dout(new_new_n1888__));
  buf1  g1345(.din(new_new_n725__), .dout(new_new_n1889__));
  buf1  g1346(.din(new_new_n732__), .dout(new_new_n1890__));
  buf1  g1347(.din(new_new_n1890__), .dout(new_new_n1891__));
  buf1  g1348(.din(new_new_n740__), .dout(new_new_n1892__));
  buf1  g1349(.din(new_new_n1892__), .dout(new_new_n1893__));
  buf1  g1350(.din(new_new_n749__), .dout(new_new_n1894__));
  buf1  g1351(.din(new_new_n741__), .dout(new_new_n1895__));
  buf1  g1352(.din(new_new_n748__), .dout(new_new_n1896__));
  buf1  g1353(.din(new_new_n1896__), .dout(new_new_n1897__));
  buf1  g1354(.din(new_new_n850__), .dout(new_new_n1898__));
  buf1  g1355(.din(new_new_n1898__), .dout(new_new_n1899__));
  buf1  g1356(.din(new_new_n1899__), .dout(new_new_n1900__));
  buf1  g1357(.din(new_new_n1899__), .dout(new_new_n1901__));
  buf1  g1358(.din(new_new_n1898__), .dout(new_new_n1902__));
  buf1  g1359(.din(new_new_n1902__), .dout(new_new_n1903__));
  buf1  g1360(.din(new_new_n1902__), .dout(new_new_n1904__));
  buf1  g1361(.din(new_new_n851__), .dout(new_new_n1905__));
  buf1  g1362(.din(new_new_n1905__), .dout(new_new_n1906__));
  buf1  g1363(.din(new_new_n1906__), .dout(new_new_n1907__));
  buf1  g1364(.din(new_new_n1906__), .dout(new_new_n1908__));
  buf1  g1365(.din(new_new_n1905__), .dout(new_new_n1909__));
  buf1  g1366(.din(new_new_n1909__), .dout(new_new_n1910__));
  buf1  g1367(.din(new_new_n1909__), .dout(new_new_n1911__));
  buf1  g1368(.din(new_new_n861__), .dout(new_new_n1912__));
  buf1  g1369(.din(new_new_n1912__), .dout(new_new_n1913__));
  buf1  g1370(.din(new_new_n1912__), .dout(new_new_n1914__));
  buf1  g1371(.din(new_new_n862__), .dout(new_new_n1915__));
  buf1  g1372(.din(new_new_n1915__), .dout(new_new_n1916__));
  buf1  g1373(.din(new_new_n1915__), .dout(new_new_n1917__));
  buf1  g1374(.din(new_new_n860__), .dout(new_new_n1918__));
  buf1  g1375(.din(new_new_n1918__), .dout(new_new_n1919__));
  buf1  g1376(.din(new_new_n1918__), .dout(new_new_n1920__));
  buf1  g1377(.din(new_new_n863__), .dout(new_new_n1921__));
  buf1  g1378(.din(new_new_n1921__), .dout(new_new_n1922__));
  buf1  g1379(.din(new_new_n1921__), .dout(new_new_n1923__));
  buf1  g1380(.din(new_new_n1182__), .dout(new_new_n1924__));
  buf1  g1381(.din(new_new_n1193__), .dout(new_new_n1925__));
  buf1  g1382(.din(new_new_n726__), .dout(new_new_n1926__));
  buf1  g1383(.din(new_new_n1926__), .dout(new_new_n1927__));
  buf1  g1384(.din(new_new_n735__), .dout(new_new_n1928__));
  buf1  g1385(.din(new_new_n727__), .dout(new_new_n1929__));
  buf1  g1386(.din(new_new_n734__), .dout(new_new_n1930__));
  buf1  g1387(.din(new_new_n1930__), .dout(new_new_n1931__));
  buf1  g1388(.din(new_new_n742__), .dout(new_new_n1932__));
  buf1  g1389(.din(new_new_n1932__), .dout(new_new_n1933__));
  buf1  g1390(.din(new_new_n751__), .dout(new_new_n1934__));
  buf1  g1391(.din(new_new_n743__), .dout(new_new_n1935__));
  buf1  g1392(.din(new_new_n750__), .dout(new_new_n1936__));
  buf1  g1393(.din(new_new_n1936__), .dout(new_new_n1937__));
  buf1  g1394(.din(new_new_n864__), .dout(new_new_n1938__));
  buf1  g1395(.din(new_new_n1938__), .dout(new_new_n1939__));
  buf1  g1396(.din(new_new_n1938__), .dout(new_new_n1940__));
  buf1  g1397(.din(new_new_n867__), .dout(new_new_n1941__));
  buf1  g1398(.din(new_new_n1941__), .dout(new_new_n1942__));
  buf1  g1399(.din(new_new_n1941__), .dout(new_new_n1943__));
  buf1  g1400(.din(new_new_n865__), .dout(new_new_n1944__));
  buf1  g1401(.din(new_new_n1944__), .dout(new_new_n1945__));
  buf1  g1402(.din(new_new_n1944__), .dout(new_new_n1946__));
  buf1  g1403(.din(new_new_n866__), .dout(new_new_n1947__));
  buf1  g1404(.din(new_new_n1947__), .dout(new_new_n1948__));
  buf1  g1405(.din(new_new_n1947__), .dout(new_new_n1949__));
  buf1  g1406(.din(new_new_n1210__), .dout(new_new_n1950__));
  buf1  g1407(.din(new_new_n1221__), .dout(new_new_n1951__));
  buf1  g1408(.din(new_new_n728__), .dout(new_new_n1952__));
  buf1  g1409(.din(new_new_n1952__), .dout(new_new_n1953__));
  buf1  g1410(.din(new_new_n737__), .dout(new_new_n1954__));
  buf1  g1411(.din(new_new_n729__), .dout(new_new_n1955__));
  buf1  g1412(.din(new_new_n736__), .dout(new_new_n1956__));
  buf1  g1413(.din(new_new_n1956__), .dout(new_new_n1957__));
  buf1  g1414(.din(new_new_n744__), .dout(new_new_n1958__));
  buf1  g1415(.din(new_new_n1958__), .dout(new_new_n1959__));
  buf1  g1416(.din(new_new_n753__), .dout(new_new_n1960__));
  buf1  g1417(.din(new_new_n745__), .dout(new_new_n1961__));
  buf1  g1418(.din(new_new_n752__), .dout(new_new_n1962__));
  buf1  g1419(.din(new_new_n1962__), .dout(new_new_n1963__));
  buf1  g1420(.din(new_new_n1238__), .dout(new_new_n1964__));
  buf1  g1421(.din(new_new_n1249__), .dout(new_new_n1965__));
  buf1  g1422(.din(new_new_n730__), .dout(new_new_n1966__));
  buf1  g1423(.din(new_new_n1966__), .dout(new_new_n1967__));
  buf1  g1424(.din(new_new_n739__), .dout(new_new_n1968__));
  buf1  g1425(.din(new_new_n731__), .dout(new_new_n1969__));
  buf1  g1426(.din(new_new_n738__), .dout(new_new_n1970__));
  buf1  g1427(.din(new_new_n1970__), .dout(new_new_n1971__));
  buf1  g1428(.din(new_new_n746__), .dout(new_new_n1972__));
  buf1  g1429(.din(new_new_n1972__), .dout(new_new_n1973__));
  buf1  g1430(.din(new_new_n755__), .dout(new_new_n1974__));
  buf1  g1431(.din(new_new_n747__), .dout(new_new_n1975__));
  buf1  g1432(.din(new_new_n754__), .dout(new_new_n1976__));
  buf1  g1433(.din(new_new_n1976__), .dout(new_new_n1977__));
  buf1  g1434(.din(new_new_n1266__), .dout(new_new_n1978__));
  buf1  g1435(.din(new_new_n1277__), .dout(new_new_n1979__));
  buf1  g1436(.din(new_new_n756__), .dout(new_new_n1980__));
  buf1  g1437(.din(new_new_n1980__), .dout(new_new_n1981__));
  buf1  g1438(.din(new_new_n765__), .dout(new_new_n1982__));
  buf1  g1439(.din(new_new_n757__), .dout(new_new_n1983__));
  buf1  g1440(.din(new_new_n764__), .dout(new_new_n1984__));
  buf1  g1441(.din(new_new_n1984__), .dout(new_new_n1985__));
  buf1  g1442(.din(new_new_n772__), .dout(new_new_n1986__));
  buf1  g1443(.din(new_new_n1986__), .dout(new_new_n1987__));
  buf1  g1444(.din(new_new_n781__), .dout(new_new_n1988__));
  buf1  g1445(.din(new_new_n773__), .dout(new_new_n1989__));
  buf1  g1446(.din(new_new_n780__), .dout(new_new_n1990__));
  buf1  g1447(.din(new_new_n1990__), .dout(new_new_n1991__));
  buf1  g1448(.din(new_new_n853__), .dout(new_new_n1992__));
  buf1  g1449(.din(new_new_n1992__), .dout(new_new_n1993__));
  buf1  g1450(.din(new_new_n1992__), .dout(new_new_n1994__));
  buf1  g1451(.din(new_new_n854__), .dout(new_new_n1995__));
  buf1  g1452(.din(new_new_n1995__), .dout(new_new_n1996__));
  buf1  g1453(.din(new_new_n1995__), .dout(new_new_n1997__));
  buf1  g1454(.din(new_new_n852__), .dout(new_new_n1998__));
  buf1  g1455(.din(new_new_n1998__), .dout(new_new_n1999__));
  buf1  g1456(.din(new_new_n1998__), .dout(new_new_n2000__));
  buf1  g1457(.din(new_new_n855__), .dout(new_new_n2001__));
  buf1  g1458(.din(new_new_n2001__), .dout(new_new_n2002__));
  buf1  g1459(.din(new_new_n2001__), .dout(new_new_n2003__));
  buf1  g1460(.din(new_new_n1294__), .dout(new_new_n2004__));
  buf1  g1461(.din(new_new_n1305__), .dout(new_new_n2005__));
  buf1  g1462(.din(new_new_n758__), .dout(new_new_n2006__));
  buf1  g1463(.din(new_new_n2006__), .dout(new_new_n2007__));
  buf1  g1464(.din(new_new_n767__), .dout(new_new_n2008__));
  buf1  g1465(.din(new_new_n759__), .dout(new_new_n2009__));
  buf1  g1466(.din(new_new_n766__), .dout(new_new_n2010__));
  buf1  g1467(.din(new_new_n2010__), .dout(new_new_n2011__));
  buf1  g1468(.din(new_new_n774__), .dout(new_new_n2012__));
  buf1  g1469(.din(new_new_n2012__), .dout(new_new_n2013__));
  buf1  g1470(.din(new_new_n783__), .dout(new_new_n2014__));
  buf1  g1471(.din(new_new_n775__), .dout(new_new_n2015__));
  buf1  g1472(.din(new_new_n782__), .dout(new_new_n2016__));
  buf1  g1473(.din(new_new_n2016__), .dout(new_new_n2017__));
  buf1  g1474(.din(new_new_n857__), .dout(new_new_n2018__));
  buf1  g1475(.din(new_new_n2018__), .dout(new_new_n2019__));
  buf1  g1476(.din(new_new_n2018__), .dout(new_new_n2020__));
  buf1  g1477(.din(new_new_n858__), .dout(new_new_n2021__));
  buf1  g1478(.din(new_new_n2021__), .dout(new_new_n2022__));
  buf1  g1479(.din(new_new_n2021__), .dout(new_new_n2023__));
  buf1  g1480(.din(new_new_n856__), .dout(new_new_n2024__));
  buf1  g1481(.din(new_new_n2024__), .dout(new_new_n2025__));
  buf1  g1482(.din(new_new_n2024__), .dout(new_new_n2026__));
  buf1  g1483(.din(new_new_n859__), .dout(new_new_n2027__));
  buf1  g1484(.din(new_new_n2027__), .dout(new_new_n2028__));
  buf1  g1485(.din(new_new_n2027__), .dout(new_new_n2029__));
  buf1  g1486(.din(new_new_n1322__), .dout(new_new_n2030__));
  buf1  g1487(.din(new_new_n1333__), .dout(new_new_n2031__));
  buf1  g1488(.din(new_new_n760__), .dout(new_new_n2032__));
  buf1  g1489(.din(new_new_n2032__), .dout(new_new_n2033__));
  buf1  g1490(.din(new_new_n769__), .dout(new_new_n2034__));
  buf1  g1491(.din(new_new_n761__), .dout(new_new_n2035__));
  buf1  g1492(.din(new_new_n768__), .dout(new_new_n2036__));
  buf1  g1493(.din(new_new_n2036__), .dout(new_new_n2037__));
  buf1  g1494(.din(new_new_n776__), .dout(new_new_n2038__));
  buf1  g1495(.din(new_new_n2038__), .dout(new_new_n2039__));
  buf1  g1496(.din(new_new_n785__), .dout(new_new_n2040__));
  buf1  g1497(.din(new_new_n777__), .dout(new_new_n2041__));
  buf1  g1498(.din(new_new_n784__), .dout(new_new_n2042__));
  buf1  g1499(.din(new_new_n2042__), .dout(new_new_n2043__));
  buf1  g1500(.din(new_new_n1350__), .dout(new_new_n2044__));
  buf1  g1501(.din(new_new_n1361__), .dout(new_new_n2045__));
  buf1  g1502(.din(new_new_n762__), .dout(new_new_n2046__));
  buf1  g1503(.din(new_new_n2046__), .dout(new_new_n2047__));
  buf1  g1504(.din(new_new_n771__), .dout(new_new_n2048__));
  buf1  g1505(.din(new_new_n763__), .dout(new_new_n2049__));
  buf1  g1506(.din(new_new_n770__), .dout(new_new_n2050__));
  buf1  g1507(.din(new_new_n2050__), .dout(new_new_n2051__));
  buf1  g1508(.din(new_new_n778__), .dout(new_new_n2052__));
  buf1  g1509(.din(new_new_n2052__), .dout(new_new_n2053__));
  buf1  g1510(.din(new_new_n787__), .dout(new_new_n2054__));
  buf1  g1511(.din(new_new_n779__), .dout(new_new_n2055__));
  buf1  g1512(.din(new_new_n786__), .dout(new_new_n2056__));
  buf1  g1513(.din(new_new_n2056__), .dout(new_new_n2057__));
  buf1  g1514(.din(new_new_n1378__), .dout(new_new_n2058__));
  buf1  g1515(.din(new_new_n1389__), .dout(new_new_n2059__));
  buf1  g1516(.din(new_new_n868__), .dout(new_new_n2060__));
  buf1  g1517(.din(new_new_n2060__), .dout(new_new_n2061__));
  buf1  g1518(.din(new_new_n871__), .dout(new_new_n2062__));
  buf1  g1519(.din(new_new_n869__), .dout(new_new_n2063__));
  buf1  g1520(.din(new_new_n870__), .dout(new_new_n2064__));
  buf1  g1521(.din(new_new_n2064__), .dout(new_new_n2065__));
  buf1  g1522(.din(new_new_n872__), .dout(new_new_n2066__));
  buf1  g1523(.din(new_new_n2066__), .dout(new_new_n2067__));
  buf1  g1524(.din(new_new_n875__), .dout(new_new_n2068__));
  buf1  g1525(.din(new_new_n873__), .dout(new_new_n2069__));
  buf1  g1526(.din(new_new_n874__), .dout(new_new_n2070__));
  buf1  g1527(.din(new_new_n2070__), .dout(new_new_n2071__));
  buf1  g1528(.din(new_new_n876__), .dout(new_new_n2072__));
  buf1  g1529(.din(new_new_n2072__), .dout(new_new_n2073__));
  buf1  g1530(.din(new_new_n879__), .dout(new_new_n2074__));
  buf1  g1531(.din(new_new_n877__), .dout(new_new_n2075__));
  buf1  g1532(.din(new_new_n878__), .dout(new_new_n2076__));
  buf1  g1533(.din(new_new_n2076__), .dout(new_new_n2077__));
  buf1  g1534(.din(new_new_n880__), .dout(new_new_n2078__));
  buf1  g1535(.din(new_new_n2078__), .dout(new_new_n2079__));
  buf1  g1536(.din(new_new_n883__), .dout(new_new_n2080__));
  buf1  g1537(.din(new_new_n881__), .dout(new_new_n2081__));
  buf1  g1538(.din(new_new_n882__), .dout(new_new_n2082__));
  buf1  g1539(.din(new_new_n2082__), .dout(new_new_n2083__));
  buf1  g1540(.din(new_new_n884__), .dout(new_new_n2084__));
  buf1  g1541(.din(new_new_n2084__), .dout(new_new_n2085__));
  buf1  g1542(.din(new_new_n887__), .dout(new_new_n2086__));
  buf1  g1543(.din(new_new_n885__), .dout(new_new_n2087__));
  buf1  g1544(.din(new_new_n886__), .dout(new_new_n2088__));
  buf1  g1545(.din(new_new_n2088__), .dout(new_new_n2089__));
  buf1  g1546(.din(new_new_n888__), .dout(new_new_n2090__));
  buf1  g1547(.din(new_new_n2090__), .dout(new_new_n2091__));
  buf1  g1548(.din(new_new_n891__), .dout(new_new_n2092__));
  buf1  g1549(.din(new_new_n889__), .dout(new_new_n2093__));
  buf1  g1550(.din(new_new_n890__), .dout(new_new_n2094__));
  buf1  g1551(.din(new_new_n2094__), .dout(new_new_n2095__));
  buf1  g1552(.din(new_new_n892__), .dout(new_new_n2096__));
  buf1  g1553(.din(new_new_n2096__), .dout(new_new_n2097__));
  buf1  g1554(.din(new_new_n895__), .dout(new_new_n2098__));
  buf1  g1555(.din(new_new_n893__), .dout(new_new_n2099__));
  buf1  g1556(.din(new_new_n894__), .dout(new_new_n2100__));
  buf1  g1557(.din(new_new_n2100__), .dout(new_new_n2101__));
  buf1  g1558(.din(new_new_n896__), .dout(new_new_n2102__));
  buf1  g1559(.din(new_new_n2102__), .dout(new_new_n2103__));
  buf1  g1560(.din(new_new_n899__), .dout(new_new_n2104__));
  buf1  g1561(.din(new_new_n897__), .dout(new_new_n2105__));
  buf1  g1562(.din(new_new_n898__), .dout(new_new_n2106__));
  buf1  g1563(.din(new_new_n2106__), .dout(new_new_n2107__));
  buf1  g1564(.din(new_new_n900__), .dout(new_new_n2108__));
  buf1  g1565(.din(new_new_n2108__), .dout(new_new_n2109__));
  buf1  g1566(.din(new_new_n903__), .dout(new_new_n2110__));
  buf1  g1567(.din(new_new_n901__), .dout(new_new_n2111__));
  buf1  g1568(.din(new_new_n902__), .dout(new_new_n2112__));
  buf1  g1569(.din(new_new_n2112__), .dout(new_new_n2113__));
  buf1  g1570(.din(new_new_n904__), .dout(new_new_n2114__));
  buf1  g1571(.din(new_new_n2114__), .dout(new_new_n2115__));
  buf1  g1572(.din(new_new_n907__), .dout(new_new_n2116__));
  buf1  g1573(.din(new_new_n905__), .dout(new_new_n2117__));
  buf1  g1574(.din(new_new_n906__), .dout(new_new_n2118__));
  buf1  g1575(.din(new_new_n2118__), .dout(new_new_n2119__));
  buf1  g1576(.din(new_new_n908__), .dout(new_new_n2120__));
  buf1  g1577(.din(new_new_n2120__), .dout(new_new_n2121__));
  buf1  g1578(.din(new_new_n911__), .dout(new_new_n2122__));
  buf1  g1579(.din(new_new_n909__), .dout(new_new_n2123__));
  buf1  g1580(.din(new_new_n910__), .dout(new_new_n2124__));
  buf1  g1581(.din(new_new_n2124__), .dout(new_new_n2125__));
  buf1  g1582(.din(new_new_n912__), .dout(new_new_n2126__));
  buf1  g1583(.din(new_new_n2126__), .dout(new_new_n2127__));
  buf1  g1584(.din(new_new_n915__), .dout(new_new_n2128__));
  buf1  g1585(.din(new_new_n913__), .dout(new_new_n2129__));
  buf1  g1586(.din(new_new_n914__), .dout(new_new_n2130__));
  buf1  g1587(.din(new_new_n2130__), .dout(new_new_n2131__));
  buf1  g1588(.din(new_new_n916__), .dout(new_new_n2132__));
  buf1  g1589(.din(new_new_n2132__), .dout(new_new_n2133__));
  buf1  g1590(.din(new_new_n919__), .dout(new_new_n2134__));
  buf1  g1591(.din(new_new_n917__), .dout(new_new_n2135__));
  buf1  g1592(.din(new_new_n918__), .dout(new_new_n2136__));
  buf1  g1593(.din(new_new_n2136__), .dout(new_new_n2137__));
  buf1  g1594(.din(new_new_n920__), .dout(new_new_n2138__));
  buf1  g1595(.din(new_new_n2138__), .dout(new_new_n2139__));
  buf1  g1596(.din(new_new_n923__), .dout(new_new_n2140__));
  buf1  g1597(.din(new_new_n921__), .dout(new_new_n2141__));
  buf1  g1598(.din(new_new_n922__), .dout(new_new_n2142__));
  buf1  g1599(.din(new_new_n2142__), .dout(new_new_n2143__));
  buf1  g1600(.din(new_new_n924__), .dout(new_new_n2144__));
  buf1  g1601(.din(new_new_n2144__), .dout(new_new_n2145__));
  buf1  g1602(.din(new_new_n927__), .dout(new_new_n2146__));
  buf1  g1603(.din(new_new_n925__), .dout(new_new_n2147__));
  buf1  g1604(.din(new_new_n926__), .dout(new_new_n2148__));
  buf1  g1605(.din(new_new_n2148__), .dout(new_new_n2149__));
  buf1  g1606(.din(new_new_n928__), .dout(new_new_n2150__));
  buf1  g1607(.din(new_new_n2150__), .dout(new_new_n2151__));
  buf1  g1608(.din(new_new_n931__), .dout(new_new_n2152__));
  buf1  g1609(.din(new_new_n929__), .dout(new_new_n2153__));
  buf1  g1610(.din(new_new_n930__), .dout(new_new_n2154__));
  buf1  g1611(.din(new_new_n2154__), .dout(new_new_n2155__));
  always @ (posedge clock) begin
    n286_lo <= n3533;
    n298_lo <= n3536;
    n310_lo <= n3539;
    n322_lo <= n3542;
    n334_lo <= n3545;
    n346_lo <= n3548;
    n358_lo <= n3551;
    n370_lo <= n3554;
    n382_lo <= n3557;
    n394_lo <= n3560;
    n406_lo <= n3563;
    n418_lo <= n3566;
    n430_lo <= n3569;
    n442_lo <= n3572;
    n454_lo <= n3575;
    n466_lo <= n3578;
    n478_lo <= n3581;
    n490_lo <= n3584;
    n502_lo <= n3587;
    n514_lo <= n3590;
    n526_lo <= n3593;
    n538_lo <= n3596;
    n550_lo <= n3599;
    n562_lo <= n3602;
    n574_lo <= n3605;
    n586_lo <= n3608;
    n598_lo <= n3611;
    n610_lo <= n3614;
    n622_lo <= n3617;
    n634_lo <= n3620;
    n646_lo <= n3623;
    n658_lo <= n3626;
    n661_lo <= n3629;
    n673_lo <= n3632;
    n685_lo <= n3635;
    n697_lo <= n3638;
    n709_lo <= n3641;
    n721_lo <= n3644;
    n733_lo <= n3647;
    n745_lo <= n3650;
    n757_lo <= n3653;
    n1589_o2 <= n3656;
    n1590_o2 <= n3659;
    n1591_o2 <= n3662;
    n1592_o2 <= n3665;
    n1593_o2 <= n3668;
    n1594_o2 <= n3671;
    n1595_o2 <= n3674;
    n1596_o2 <= n3677;
    n1597_o2 <= n3680;
    n1598_o2 <= n3683;
    n1599_o2 <= n3686;
    n1600_o2 <= n3689;
    n1601_o2 <= n3692;
    n1602_o2 <= n3695;
    n1603_o2 <= n3698;
    n1604_o2 <= n3701;
    n1605_o2 <= n3704;
    n1606_o2 <= n3707;
    n1607_o2 <= n3710;
    n1608_o2 <= n3713;
    n1609_o2 <= n3716;
    n1610_o2 <= n3719;
    n1611_o2 <= n3722;
    n1612_o2 <= n3725;
    n1613_o2 <= n3728;
    n1614_o2 <= n3731;
    n1615_o2 <= n3734;
    n1616_o2 <= n3737;
    n1617_o2 <= n3740;
    n1618_o2 <= n3743;
    n1619_o2 <= n3746;
    n1620_o2 <= n3749;
    n602_o2 <= n3752;
    n639_o2 <= n3755;
    n678_o2 <= n3758;
    n658_o2 <= n3761;
    n783_o2 <= n3764;
    n802_o2 <= n3767;
    n726_o2 <= n3770;
    n763_o2 <= n3773;
    n685_o2 <= n3776;
    n680_o2 <= n3779;
    n822_o2 <= n3782;
    n843_o2 <= n3785;
    n842_o2 <= n3788;
    n681_o2 <= n3791;
    n684_o2 <= n3794;
    n686_o2 <= n3797;
    n823_o2 <= n3800;
    lo002_buf_o2 <= n3803;
    lo006_buf_o2 <= n3806;
    lo010_buf_o2 <= n3809;
    lo014_buf_o2 <= n3812;
    lo018_buf_o2 <= n3815;
    lo022_buf_o2 <= n3818;
    lo026_buf_o2 <= n3821;
    lo030_buf_o2 <= n3824;
    lo034_buf_o2 <= n3827;
    lo038_buf_o2 <= n3830;
    lo042_buf_o2 <= n3833;
    lo046_buf_o2 <= n3836;
    lo050_buf_o2 <= n3839;
    lo054_buf_o2 <= n3842;
    lo058_buf_o2 <= n3845;
    lo062_buf_o2 <= n3848;
    lo066_buf_o2 <= n3851;
    lo070_buf_o2 <= n3854;
    lo074_buf_o2 <= n3857;
    lo078_buf_o2 <= n3860;
    lo082_buf_o2 <= n3863;
    lo086_buf_o2 <= n3866;
    lo090_buf_o2 <= n3869;
    lo094_buf_o2 <= n3872;
    lo098_buf_o2 <= n3875;
    lo102_buf_o2 <= n3878;
    lo106_buf_o2 <= n3881;
    lo110_buf_o2 <= n3884;
    lo114_buf_o2 <= n3887;
    lo118_buf_o2 <= n3890;
    lo122_buf_o2 <= n3893;
    lo126_buf_o2 <= n3896;
    n683_o2 <= n3899;
    n688_o2 <= n3902;
    n803_o2 <= n3905;
    n862_o2 <= n3908;
    n764_o2 <= n3911;
    n863_o2 <= n3914;
    n886_o2 <= n3917;
    n600_o2 <= n3920;
    n601_o2 <= n3923;
    n637_o2 <= n3926;
    n638_o2 <= n3929;
    n676_o2 <= n3932;
    n677_o2 <= n3935;
    n656_o2 <= n3938;
    n657_o2 <= n3941;
    n781_o2 <= n3944;
    n782_o2 <= n3947;
    n800_o2 <= n3950;
    n801_o2 <= n3953;
    n724_o2 <= n3956;
    n725_o2 <= n3959;
    n761_o2 <= n3962;
    n762_o2 <= n3965;
    lo129_buf_o2 <= n3968;
    lo133_buf_o2 <= n3971;
    lo137_buf_o2 <= n3974;
    lo141_buf_o2 <= n3977;
    lo145_buf_o2 <= n3980;
    lo149_buf_o2 <= n3983;
    lo153_buf_o2 <= n3986;
    lo157_buf_o2 <= n3989;
    lo161_buf_o2 <= n3992;
    n708_o2 <= n3995;
    n745_o2 <= n3998;
    n717_o2 <= n4001;
    n754_o2 <= n4004;
    n584_o2 <= n4007;
    n593_o2 <= n4010;
    n630_o2 <= n4013;
    n621_o2 <= n4016;
    lo001_buf_o2 <= n4019;
    lo005_buf_o2 <= n4022;
    lo009_buf_o2 <= n4025;
    lo013_buf_o2 <= n4028;
    lo017_buf_o2 <= n4031;
    lo021_buf_o2 <= n4034;
    lo025_buf_o2 <= n4037;
    lo029_buf_o2 <= n4040;
    lo033_buf_o2 <= n4043;
    lo037_buf_o2 <= n4046;
    lo041_buf_o2 <= n4049;
    lo045_buf_o2 <= n4052;
    lo049_buf_o2 <= n4055;
    lo053_buf_o2 <= n4058;
    lo057_buf_o2 <= n4061;
    lo061_buf_o2 <= n4064;
    lo065_buf_o2 <= n4067;
    lo069_buf_o2 <= n4070;
    lo073_buf_o2 <= n4073;
    lo077_buf_o2 <= n4076;
    lo081_buf_o2 <= n4079;
    lo085_buf_o2 <= n4082;
    lo089_buf_o2 <= n4085;
    lo093_buf_o2 <= n4088;
    lo097_buf_o2 <= n4091;
    lo101_buf_o2 <= n4094;
    lo105_buf_o2 <= n4097;
    lo109_buf_o2 <= n4100;
    lo113_buf_o2 <= n4103;
    lo117_buf_o2 <= n4106;
    lo121_buf_o2 <= n4109;
    lo125_buf_o2 <= n4112;
  end
  initial begin
    n286_lo <= 1'b0;
    n298_lo <= 1'b0;
    n310_lo <= 1'b0;
    n322_lo <= 1'b0;
    n334_lo <= 1'b0;
    n346_lo <= 1'b0;
    n358_lo <= 1'b0;
    n370_lo <= 1'b0;
    n382_lo <= 1'b0;
    n394_lo <= 1'b0;
    n406_lo <= 1'b0;
    n418_lo <= 1'b0;
    n430_lo <= 1'b0;
    n442_lo <= 1'b0;
    n454_lo <= 1'b0;
    n466_lo <= 1'b0;
    n478_lo <= 1'b0;
    n490_lo <= 1'b0;
    n502_lo <= 1'b0;
    n514_lo <= 1'b0;
    n526_lo <= 1'b0;
    n538_lo <= 1'b0;
    n550_lo <= 1'b0;
    n562_lo <= 1'b0;
    n574_lo <= 1'b0;
    n586_lo <= 1'b0;
    n598_lo <= 1'b0;
    n610_lo <= 1'b0;
    n622_lo <= 1'b0;
    n634_lo <= 1'b0;
    n646_lo <= 1'b0;
    n658_lo <= 1'b0;
    n661_lo <= 1'b0;
    n673_lo <= 1'b0;
    n685_lo <= 1'b0;
    n697_lo <= 1'b0;
    n709_lo <= 1'b0;
    n721_lo <= 1'b0;
    n733_lo <= 1'b0;
    n745_lo <= 1'b0;
    n757_lo <= 1'b0;
    n1589_o2 <= 1'b0;
    n1590_o2 <= 1'b0;
    n1591_o2 <= 1'b0;
    n1592_o2 <= 1'b0;
    n1593_o2 <= 1'b0;
    n1594_o2 <= 1'b0;
    n1595_o2 <= 1'b0;
    n1596_o2 <= 1'b0;
    n1597_o2 <= 1'b0;
    n1598_o2 <= 1'b0;
    n1599_o2 <= 1'b0;
    n1600_o2 <= 1'b0;
    n1601_o2 <= 1'b0;
    n1602_o2 <= 1'b0;
    n1603_o2 <= 1'b0;
    n1604_o2 <= 1'b0;
    n1605_o2 <= 1'b0;
    n1606_o2 <= 1'b0;
    n1607_o2 <= 1'b0;
    n1608_o2 <= 1'b0;
    n1609_o2 <= 1'b0;
    n1610_o2 <= 1'b0;
    n1611_o2 <= 1'b0;
    n1612_o2 <= 1'b0;
    n1613_o2 <= 1'b0;
    n1614_o2 <= 1'b0;
    n1615_o2 <= 1'b0;
    n1616_o2 <= 1'b0;
    n1617_o2 <= 1'b0;
    n1618_o2 <= 1'b0;
    n1619_o2 <= 1'b0;
    n1620_o2 <= 1'b0;
    n602_o2 <= 1'b0;
    n639_o2 <= 1'b0;
    n678_o2 <= 1'b0;
    n658_o2 <= 1'b0;
    n783_o2 <= 1'b0;
    n802_o2 <= 1'b0;
    n726_o2 <= 1'b0;
    n763_o2 <= 1'b0;
    n685_o2 <= 1'b0;
    n680_o2 <= 1'b0;
    n822_o2 <= 1'b0;
    n843_o2 <= 1'b0;
    n842_o2 <= 1'b0;
    n681_o2 <= 1'b0;
    n684_o2 <= 1'b0;
    n686_o2 <= 1'b0;
    n823_o2 <= 1'b0;
    lo002_buf_o2 <= 1'b0;
    lo006_buf_o2 <= 1'b0;
    lo010_buf_o2 <= 1'b0;
    lo014_buf_o2 <= 1'b0;
    lo018_buf_o2 <= 1'b0;
    lo022_buf_o2 <= 1'b0;
    lo026_buf_o2 <= 1'b0;
    lo030_buf_o2 <= 1'b0;
    lo034_buf_o2 <= 1'b0;
    lo038_buf_o2 <= 1'b0;
    lo042_buf_o2 <= 1'b0;
    lo046_buf_o2 <= 1'b0;
    lo050_buf_o2 <= 1'b0;
    lo054_buf_o2 <= 1'b0;
    lo058_buf_o2 <= 1'b0;
    lo062_buf_o2 <= 1'b0;
    lo066_buf_o2 <= 1'b0;
    lo070_buf_o2 <= 1'b0;
    lo074_buf_o2 <= 1'b0;
    lo078_buf_o2 <= 1'b0;
    lo082_buf_o2 <= 1'b0;
    lo086_buf_o2 <= 1'b0;
    lo090_buf_o2 <= 1'b0;
    lo094_buf_o2 <= 1'b0;
    lo098_buf_o2 <= 1'b0;
    lo102_buf_o2 <= 1'b0;
    lo106_buf_o2 <= 1'b0;
    lo110_buf_o2 <= 1'b0;
    lo114_buf_o2 <= 1'b0;
    lo118_buf_o2 <= 1'b0;
    lo122_buf_o2 <= 1'b0;
    lo126_buf_o2 <= 1'b0;
    n683_o2 <= 1'b0;
    n688_o2 <= 1'b0;
    n803_o2 <= 1'b0;
    n862_o2 <= 1'b0;
    n764_o2 <= 1'b0;
    n863_o2 <= 1'b0;
    n886_o2 <= 1'b0;
    n600_o2 <= 1'b0;
    n601_o2 <= 1'b0;
    n637_o2 <= 1'b0;
    n638_o2 <= 1'b0;
    n676_o2 <= 1'b0;
    n677_o2 <= 1'b0;
    n656_o2 <= 1'b0;
    n657_o2 <= 1'b0;
    n781_o2 <= 1'b0;
    n782_o2 <= 1'b0;
    n800_o2 <= 1'b0;
    n801_o2 <= 1'b0;
    n724_o2 <= 1'b0;
    n725_o2 <= 1'b0;
    n761_o2 <= 1'b0;
    n762_o2 <= 1'b0;
    lo129_buf_o2 <= 1'b0;
    lo133_buf_o2 <= 1'b0;
    lo137_buf_o2 <= 1'b0;
    lo141_buf_o2 <= 1'b0;
    lo145_buf_o2 <= 1'b0;
    lo149_buf_o2 <= 1'b0;
    lo153_buf_o2 <= 1'b0;
    lo157_buf_o2 <= 1'b0;
    lo161_buf_o2 <= 1'b0;
    n708_o2 <= 1'b0;
    n745_o2 <= 1'b0;
    n717_o2 <= 1'b0;
    n754_o2 <= 1'b0;
    n584_o2 <= 1'b0;
    n593_o2 <= 1'b0;
    n630_o2 <= 1'b0;
    n621_o2 <= 1'b0;
    lo001_buf_o2 <= 1'b0;
    lo005_buf_o2 <= 1'b0;
    lo009_buf_o2 <= 1'b0;
    lo013_buf_o2 <= 1'b0;
    lo017_buf_o2 <= 1'b0;
    lo021_buf_o2 <= 1'b0;
    lo025_buf_o2 <= 1'b0;
    lo029_buf_o2 <= 1'b0;
    lo033_buf_o2 <= 1'b0;
    lo037_buf_o2 <= 1'b0;
    lo041_buf_o2 <= 1'b0;
    lo045_buf_o2 <= 1'b0;
    lo049_buf_o2 <= 1'b0;
    lo053_buf_o2 <= 1'b0;
    lo057_buf_o2 <= 1'b0;
    lo061_buf_o2 <= 1'b0;
    lo065_buf_o2 <= 1'b0;
    lo069_buf_o2 <= 1'b0;
    lo073_buf_o2 <= 1'b0;
    lo077_buf_o2 <= 1'b0;
    lo081_buf_o2 <= 1'b0;
    lo085_buf_o2 <= 1'b0;
    lo089_buf_o2 <= 1'b0;
    lo093_buf_o2 <= 1'b0;
    lo097_buf_o2 <= 1'b0;
    lo101_buf_o2 <= 1'b0;
    lo105_buf_o2 <= 1'b0;
    lo109_buf_o2 <= 1'b0;
    lo113_buf_o2 <= 1'b0;
    lo117_buf_o2 <= 1'b0;
    lo121_buf_o2 <= 1'b0;
    lo125_buf_o2 <= 1'b0;
  end
endmodule


