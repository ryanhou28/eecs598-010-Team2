module c3540(G1,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,
  G24,G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G34,G35,G3519,G3520,G3521,G3522,
  G3523,G3524,G3525,G3526,G3527,G3528,G3529,G3530,G3531,G3532,G3533,G3534,
  G3535,G3536,G3537,G3538,G3539,G3540,G36,G37,G38,G39,G4,G40,G41,G42,G43,G44,
  G45,G46,G47,G48,G49,G5,G50,G6,G7,G8,G9);
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
  G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,
  G40,G41,G42,G43,G44,G45,G46,G47,G48,G49,G50;
output G3519,G3520,G3521,G3522,G3523,G3524,G3525,G3526,G3527,G3528,G3529,G3530,
  G3531,G3532,G3533,G3534,G3535,G3536,G3537,G3538,G3539,G3540;

  wire G353,G363,G368,G377,G381,G384,G388,G397,G400,G404,G413,G422,G425,G434,
    G438,G447,G451,G461,G466,G467,G470,G477,G480,G484,G491,G492,G496,G501,G518,
    G519,G523,G527,G530,G533,G534,G537,G540,G543,G546,G549,G552,G556,G559,G562,
    G565,G568,G572,G575,G578,G581,G584,G587,G588,G589,G590,G593,G594,G611,G612,
    G613,G614,G615,G618,G621,G624,G627,G630,G633,G636,G639,G642,G645,G648,G651,
    G654,G657,G660,G663,G666,G667,G684,G685,G686,G691,G708,G713,G714,G715,G716,
    G717,G718,G719,G720,G721,G722,G723,G724,G725,G726,G727,G730,G731,G734,G735,
    G736,G739,G742,G745,G749,G753,G762,G769,G772,G775,G778,G781,G784,G785,G786,
    G787,G790,G791,G792,G793,G794,G795,G796,G797,G798,G799,G800,G805,G810,G813,
    G816,G831,G848,G849,G850,G851,G852,G853,G854,G855,G856,G873,G874,G875,G882,
    G883,G884,G887,G890,G891,G892,G893,G894,G897,G898,G901,G904,G907,G910,G913,
    G916,G919,G922,G925,G928,G929,G930,G931,G932,G933,G934,G935,G939,G956,G957,
    G958,G959,G960,G961,G962,G963,G964,G965,G966,G967,G968,G969,G970,G971,G972,
    G973,G974,G975,G976,G977,G978,G979,G980,G981,G982,G983,G984,G985,G986,G989,
    G992,G993,G994,G995,G996,G997,G998,G999,G1000,G1001,G1002,G1003,G1004,
    G1005,G1008,G1011,G1012,G1015,G1016,G1017,G1018,G1019,G1020,G1021,G1022,
    G1023,G1024,G1025,G1034,G1043,G1048,G1051,G1052,G1053,G1054,G1055,G1056,
    G1057,G1058,G1059,G1060,G1061,G1062,G1063,G1064,G1065,G1066,G1067,G1068,
    G1069,G1070,G1071,G1072,G1073,G1074,G1077,G1080,G1083,G1086,G1089,G1092,
    G1095,G1104,G1113,G1114,G1115,G1116,G1117,G1118,G1119,G1120,G1121,G1122,
    G1123,G1124,G1125,G1126,G1127,G1128,G1129,G1130,G1131,G1132,G1133,G1134,
    G1135,G1136,G1137,G1140,G1141,G1142,G1145,G1146,G1147,G1150,G1151,G1152,
    G1155,G1156,G1157,G1160,G1161,G1162,G1165,G1166,G1167,G1170,G1171,G1172,
    G1175,G1176,G1179,G1180,G1184,G1189,G1193,G1197,G1200,G1203,G1206,G1207,
    G1208,G1209,G1210,G1211,G1212,G1213,G1214,G1215,G1216,G1217,G1218,G1219,
    G1222,G1223,G1224,G1225,G1226,G1227,G1228,G1229,G1230,G1231,G1232,G1233,
    G1234,G1235,G1236,G1237,G1238,G1239,G1240,G1241,G1242,G1243,G1244,G1249,
    G1258,G1263,G1272,G1275,G1278,G1281,G1284,G1287,G1290,G1293,G1296,G1297,
    G1298,G1299,G1300,G1301,G1302,G1303,G1304,G1305,G1306,G1307,G1308,G1309,
    G1310,G1311,G1312,G1313,G1314,G1315,G1316,G1317,G1318,G1319,G1320,G1321,
    G1322,G1323,G1324,G1325,G1326,G1327,G1328,G1345,G1348,G1349,G1350,G1351,
    G1352,G1353,G1354,G1357,G1360,G1363,G1366,G1369,G1372,G1375,G1378,G1379,
    G1380,G1381,G1390,G1399,G1400,G1401,G1402,G1403,G1404,G1405,G1406,G1407,
    G1408,G1409,G1410,G1411,G1412,G1413,G1414,G1415,G1418,G1421,G1424,G1427,
    G1430,G1433,G1436,G1439,G1442,G1445,G1448,G1451,G1454,G1457,G1460,G1463,
    G1466,G1467,G1468,G1469,G1470,G1471,G1472,G1473,G1474,G1475,G1476,G1477,
    G1478,G1479,G1482,G1485,G1486,G1487,G1488,G1489,G1490,G1491,G1492,G1493,
    G1494,G1495,G1496,G1497,G1498,G1499,G1500,G1501,G1502,G1503,G1504,G1505,
    G1506,G1507,G1508,G1509,G1510,G1511,G1512,G1513,G1514,G1517,G1518,G1519,
    G1520,G1521,G1522,G1523,G1524,G1527,G1528,G1529,G1538,G1547,G1556,G1565,
    G1574,G1583,G1592,G1601,G1610,G1619,G1628,G1637,G1646,G1655,G1664,G1673,
    G1674,G1675,G1676,G1677,G1678,G1679,G1680,G1681,G1682,G1683,G1684,G1685,
    G1686,G1687,G1688,G1689,G1693,G1697,G1700,G1703,G1707,G1711,G1714,G1718,
    G1722,G1725,G1729,G1733,G1738,G1743,G1747,G1751,G1756,G1760,G1764,G1769,
    G1770,G1771,G1772,G1773,G1774,G1775,G1776,G1777,G1778,G1779,G1780,G1781,
    G1782,G1783,G1784,G1785,G1786,G1787,G1788,G1789,G1790,G1791,G1792,G1793,
    G1794,G1795,G1796,G1799,G1802,G1805,G1806,G1807,G1808,G1809,G1810,G1811,
    G1812,G1813,G1816,G1819,G1823,G1826,G1827,G1828,G1829,G1830,G1831,G1832,
    G1833,G1834,G1835,G1836,G1837,G1838,G1839,G1840,G1841,G1842,G1843,G1844,
    G1845,G1846,G1847,G1848,G1849,G1850,G1851,G1852,G1853,G1854,G1855,G1856,
    G1857,G1858,G1859,G1860,G1861,G1862,G1863,G1864,G1865,G1866,G1867,G1868,
    G1869,G1870,G1871,G1872,G1873,G1874,G1875,G1876,G1877,G1878,G1879,G1880,
    G1881,G1882,G1883,G1884,G1885,G1886,G1887,G1888,G1889,G1890,G1891,G1892,
    G1893,G1894,G1895,G1896,G1897,G1898,G1899,G1900,G1901,G1902,G1903,G1904,
    G1905,G1906,G1907,G1908,G1909,G1910,G1911,G1912,G1913,G1914,G1915,G1916,
    G1917,G1918,G1919,G1920,G1921,G1922,G1923,G1924,G1925,G1926,G1927,G1928,
    G1929,G1930,G1931,G1932,G1933,G1934,G1935,G1936,G1937,G1938,G1939,G1940,
    G1941,G1942,G1943,G1944,G1945,G1946,G1947,G1948,G1949,G1950,G1951,G1952,
    G1953,G1954,G1955,G1958,G1961,G1962,G1965,G1968,G1971,G1974,G1977,G1978,
    G1981,G1984,G1985,G1988,G1991,G1992,G1995,G1998,G2001,G2004,G2007,G2008,
    G2011,G2014,G2015,G2018,G2021,G2024,G2027,G2030,G2033,G2034,G2035,G2036,
    G2037,G2038,G2039,G2040,G2041,G2042,G2043,G2044,G2045,G2046,G2047,G2048,
    G2049,G2050,G2051,G2052,G2053,G2054,G2055,G2056,G2057,G2058,G2059,G2060,
    G2061,G2062,G2063,G2064,G2065,G2066,G2067,G2068,G2069,G2070,G2071,G2072,
    G2073,G2074,G2075,G2076,G2077,G2078,G2079,G2080,G2081,G2082,G2083,G2084,
    G2085,G2086,G2087,G2088,G2089,G2090,G2091,G2092,G2093,G2094,G2095,G2096,
    G2097,G2098,G2099,G2100,G2101,G2102,G2103,G2104,G2105,G2106,G2107,G2108,
    G2109,G2110,G2111,G2112,G2113,G2114,G2115,G2116,G2117,G2118,G2119,G2120,
    G2121,G2122,G2123,G2124,G2125,G2126,G2127,G2128,G2129,G2130,G2131,G2132,
    G2133,G2134,G2135,G2136,G2137,G2138,G2139,G2140,G2141,G2142,G2143,G2144,
    G2145,G2146,G2147,G2148,G2149,G2150,G2151,G2152,G2153,G2154,G2155,G2156,
    G2157,G2158,G2159,G2160,G2161,G2162,G2163,G2164,G2165,G2166,G2167,G2168,
    G2169,G2172,G2173,G2174,G2175,G2176,G2177,G2178,G2179,G2180,G2181,G2182,
    G2183,G2184,G2185,G2186,G2187,G2188,G2189,G2190,G2191,G2192,G2195,G2198,
    G2199,G2200,G2204,G2208,G2211,G2214,G2215,G2216,G2219,G2222,G2223,G2224,
    G2227,G2230,G2231,G2232,G2236,G2240,G2243,G2246,G2247,G2248,G2251,G2254,
    G2255,G2256,G2257,G2260,G2263,G2266,G2269,G2272,G2275,G2278,G2281,G2284,
    G2287,G2290,G2293,G2296,G2299,G2302,G2305,G2308,G2311,G2312,G2313,G2314,
    G2315,G2316,G2317,G2318,G2319,G2320,G2321,G2322,G2323,G2324,G2325,G2326,
    G2327,G2328,G2329,G2330,G2331,G2332,G2333,G2334,G2335,G2336,G2337,G2338,
    G2339,G2340,G2341,G2342,G2343,G2344,G2345,G2346,G2347,G2348,G2349,G2350,
    G2351,G2352,G2353,G2354,G2355,G2356,G2359,G2362,G2363,G2364,G2365,G2368,
    G2369,G2372,G2373,G2374,G2375,G2378,G2381,G2382,G2383,G2384,G2387,G2388,
    G2391,G2392,G2393,G2396,G2397,G2398,G2399,G2400,G2401,G2404,G2405,G2406,
    G2407,G2408,G2411,G2414,G2415,G2416,G2417,G2418,G2419,G2420,G2421,G2422,
    G2423,G2424,G2425,G2426,G2427,G2428,G2429,G2430,G2436,G2437,G2441,G2444,
    G2450,G2451,G2455,G2458,G2459,G2460,G2461,G2462,G2463,G2464,G2465,G2466,
    G2467,G2468,G2471,G2472,G2475,G2476,G2479,G2482,G2485,G2488,G2491,G2494,
    G2497,G2500,G2501,G2502,G2507,G2512,G2515,G2518,G2521,G2524,G2527,G2530,
    G2531,G2532,G2533,G2534,G2535,G2536,G2537,G2538,G2539,G2542,G2543,G2546,
    G2547,G2550,G2551,G2552,G2556,G2557,G2558,G2561,G2562,G2563,G2566,G2569,
    G2570,G2571,G2574,G2577,G2580,G2583,G2586,G2589,G2592,G2595,G2598,G2601,
    G2604,G2607,G2610,G2613,G2614,G2615,G2616,G2617,G2618,G2619,G2620,G2623,
    G2624,G2625,G2626,G2627,G2628,G2629,G2630,G2631,G2632,G2633,G2634,G2635,
    G2636,G2637,G2638,G2639,G2640,G2643,G2646,G2647,G2648,G2651,G2654,G2655,
    G2656,G2657,G2658,G2659,G2660,G2661,G2662,G2663,G2664,G2665,G2666,G2669,
    G2673,G2674,G2675,G2676,G2677,G2678,G2679,G2680,G2681,G2682,G2683,G2684,
    G2685,G2686,G2687,G2690,G2693,G2694,G2697,G2698,G2699,G2705,G2708,G2711,
    G2712,G2713,G2714,G2715,G2716,G2717,G2718,G2719,G2720,G2721,G2728,G2733,
    G2736,G2739,G2740,G2741,G2742,G2743,G2744,G2745,G2746,G2747,G2750,G2753,
    G2759,G2763,G2768,G2773,G2778,G2779,G2780,G2781,G2784,G2787,G2788,G2789,
    G2790,G2791,G2792,G2793,G2794,G2795,G2796,G2799,G2803,G2804,G2805,G2808,
    G2809,G2810,G2811,G2816,G2820,G2821,G2822,G2823,G2826,G2827,G2828,G2829,
    G2830,G2831,G2832,G2833,G2836,G2839,G2842,G2845,G2848,G2851,G2854,G2857,
    G2860,G2863,G2866,G2869,G2872,G2875,G2876,G2877,G2880,G2883,G2884,G2887,
    G2890,G2893,G2896,G2899,G2902,G2905,G2906,G2909,G2910,G2911,G2912,G2913,
    G2916,G2917,G2918,G2919,G2920,G2923,G2926,G2929,G2932,G2935,G2936,G2937,
    G2938,G2939,G2942,G2943,G2944,G2947,G2950,G2951,G2952,G2953,G2954,G2955,
    G2956,G2957,G2958,G2959,G2960,G2961,G2962,G2965,G2968,G2971,G2974,G2975,
    G2978,G2979,G2980,G2981,G2984,G2985,G2986,G2990,G2991,G2994,G2995,G2996,
    G2999,G3002,G3005,G3006,G3007,G3010,G3011,G3012,G3015,G3016,G3017,G3018,
    G3021,G3024,G3027,G3030,G3031,G3032,G3033,G3034,G3035,G3036,G3037,G3038,
    G3039,G3042,G3045,G3048,G3051,G3054,G3057,G3058,G3059,G3060,G3061,G3062,
    G3063,G3064,G3065,G3066,G3067,G3068,G3069,G3072,G3075,G3078,G3081,G3082,
    G3083,G3084,G3085,G3086,G3089,G3090,G3094,G3095,G3099,G3100,G3103,G3106,
    G3107,G3110,G3114,G3115,G3116,G3117,G3118,G3119,G3120,G3121,G3122,G3126,
    G3129,G3132,G3135,G3136,G3137,G3138,G3139,G3140,G3143,G3146,G3149,G3152,
    G3155,G3158,G3159,G3160,G3164,G3165,G3168,G3169,G3170,G3171,G3174,G3177,
    G3180,G3183,G3186,G3189,G3190,G3191,G3192,G3193,G3194,G3195,G3199,G3202,
    G3203,G3206,G3207,G3208,G3209,G3210,G3211,G3212,G3213,G3214,G3215,G3216,
    G3217,G3220,G3223,G3226,G3227,G3230,G3231,G3232,G3233,G3234,G3235,G3236,
    G3237,G3240,G3243,G3246,G3247,G3248,G3249,G3250,G3251,G3254,G3257,G3258,
    G3259,G3260,G3261,G3262,G3265,G3266,G3267,G3268,G3269,G3270,G3271,G3272,
    G3275,G3278,G3281,G3284,G3287,G3288,G3291,G3294,G3297,G3300,G3301,G3302,
    G3305,G3308,G3311,G3312,G3317,G3320,G3323,G3326,G3329,G3332,G3337,G3340,
    G3341,G3342,G3343,G3344,G3345,G3346,G3347,G3350,G3353,G3356,G3359,G3360,
    G3363,G3366,G3367,G3370,G3373,G3376,G3379,G3380,G3383,G3386,G3387,G3388,
    G3391,G3394,G3395,G3396,G3399,G3402,G3403,G3404,G3405,G3406,G3407,G3408,
    G3409,G3412,G3415,G3416,G3417,G3418,G3419,G3420,G3421,G3422,G3423,G3424,
    G3425,G3428,G3429,G3430,G3431,G3432,G3436,G3437,G3438,G3439,G3440,G3441,
    G3444,G3445,G3448,G3449,G3452,G3453,G3456,G3459,G3460,G3461,G3464,G3465,
    G3466,G3467,G3468,G3471,G3474,G3475,G3478,G3481,G3484,G3487,G3488,G3489,
    G3490,G3491,G3494,G3497,G3500,G3503,G3504,G3505,G3506,G3507,G3508,G3509,
    G3510,G3511,G3512,G3513,G3514,G3515,G3516,G3517,G3518;

  not (G353,G7);
  not (G363,G7);
  not (G368,G8);
  not (G377,G8);
  not (G381,G9);
  not (G384,G9);
  not (G388,G9);
  not (G397,G10);
  not (G400,G10);
  not (G404,G10);
  not (G413,G11);
  not (G422,G11);
  not (G425,G12);
  not (G434,G12);
  not (G438,G13);
  not (G447,G13);
  not (G451,G14);
  not (G461,G14);
  or (G466,G35,G36);
  not (G467,G1);
  not (G470,G1);
  not (G477,G1);
  not (G480,G2);
  not (G484,G2);
  and (G491,G2,G3);
  not (G492,G3);
  not (G496,G3);
  not (G501,G3);
  not (G518,G4);
  not (G519,G4);
  not (G523,G4);
  and (G527,G4,G5);
  not (G530,G5);
  or (G533,G5,G6);
  not (G534,G6);
  not (G537,G6);
  not (G540,G7);
  not (G543,G8);
  not (G546,G8);
  not (G549,G9);
  not (G552,G9);
  not (G556,G11);
  not (G559,G11);
  not (G562,G12);
  not (G565,G12);
  not (G568,G13);
  not (G572,G1);
  not (G575,G9);
  not (G578,G13);
  not (G581,G3);
  not (G584,G25);
  not (G587,G26);
  and (G588,G3,G26);
  nand (G589,G3,G26);
  and (G590,G3,G24);
  not (G593,G3);
  or (G594,G49,G4);
  nand (G611,G1,G2);
  nand (G612,G1,G3,G4);
  not (G613,G3);
  not (G614,G4);
  not (G615,G24);
  not (G618,G27);
  not (G621,G48);
  not (G624,G30);
  not (G627,G31);
  not (G630,G32);
  not (G633,G33);
  not (G636,G34);
  not (G639,G35);
  not (G642,G36);
  not (G645,G37);
  not (G648,G7);
  not (G651,G8);
  not (G654,G8);
  not (G657,G12);
  not (G660,G12);
  not (G663,G47);
  and (G666,G34,G466);
  or (G667,G518,G3);
  or (G684,G593,G23);
  not (G685,G491);
  or (G686,G613,G1);
  and (G691,G611,G612);
  or (G708,G614,G1);
  and (G713,G540,G546,G552);
  nand (G714,G30,G353);
  nand (G715,G31,G368);
  nand (G716,G32,G388);
  nand (G717,G33,G404);
  nand (G718,G34,G413);
  nand (G719,G35,G425);
  nand (G720,G36,G438);
  nand (G721,G37,G451);
  not (G722,G624);
  not (G723,G627);
  not (G724,G630);
  not (G725,G633);
  nand (G726,G377,G384);
  nand (G727,G434,G447);
  nand (G730,G381,G397);
  not (G731,G363);
  not (G734,G651);
  not (G735,G657);
  not (G736,G537);
  not (G739,G537);
  not (G742,G480);
  not (G745,G523);
  not (G749,G530);
  and (G753,G477,G533);
  and (G762,G477,G534,G530);
  and (G769,G467,G534);
  and (G772,G470,G484,G496);
  nand (G775,G470,G484,G496);
  nand (G778,G470,G484);
  not (G781,G572);
  nand (G784,G480,G492,G6);
  nand (G785,G540,G546,G552);
  not (G786,G654);
  and (G787,G559,G565,G568);
  nand (G790,G559,G565,G568);
  not (G791,G660);
  not (G792,G501);
  not (G793,G501);
  not (G794,G501);
  not (G795,G501);
  not (G796,G501);
  not (G797,G501);
  not (G798,G501);
  not (G799,G501);
  or (G800,G581,G584);
  nor (G805,G581,G584);
  not (G810,G590);
  not (G813,G590);
  not (G816,G519);
  not (G831,G523);
  not (G848,G594);
  not (G849,G594);
  not (G850,G594);
  not (G851,G594);
  not (G852,G594);
  not (G853,G594);
  not (G854,G594);
  not (G855,G594);
  or (G856,G1,G685);
  not (G873,G527);
  not (G874,G527);
  and (G875,G467,G480,G492);
  not (G882,G615);
  not (G883,G663);
  or (G884,G618,G621);
  nor (G887,G618,G621);
  not (G890,G636);
  not (G891,G639);
  not (G892,G642);
  not (G893,G645);
  not (G894,G377);
  not (G897,G648);
  not (G898,G384);
  not (G901,G400);
  not (G904,G422);
  not (G907,G434);
  not (G910,G447);
  not (G913,G461);
  not (G916,G575);
  not (G919,G575);
  not (G922,G578);
  not (G925,G578);
  nand (G928,G400,G713);
  and (G929,G714,G715,G716,G717);
  and (G930,G718,G719,G720,G721);
  nand (G931,G627,G722);
  nand (G932,G624,G723);
  nand (G933,G633,G724);
  nand (G934,G630,G725);
  and (G935,G353,G726);
  and (G939,G572,G784);
  not (G956,G667);
  and (G957,G501,G667);
  and (G958,G785,G792);
  not (G959,G667);
  and (G960,G501,G667);
  not (G961,G667);
  and (G962,G501,G667);
  and (G963,G552,G794);
  not (G964,G667);
  and (G965,G501,G667);
  and (G966,G10,G795);
  not (G967,G667);
  and (G968,G501,G667);
  and (G969,G790,G796);
  not (G970,G667);
  and (G971,G501,G667);
  not (G972,G667);
  and (G973,G501,G667);
  and (G974,G568,G798);
  not (G975,G667);
  and (G976,G501,G667);
  and (G977,G14,G799);
  and (G978,G28,G848);
  and (G979,G29,G849);
  and (G980,G30,G850);
  and (G981,G31,G851);
  and (G982,G32,G852);
  and (G983,G33,G853);
  and (G984,G34,G854);
  and (G985,G35,G855);
  and (G986,G1,G2,G873);
  and (G989,G1,G2,G874);
  not (G992,G691);
  not (G993,G691);
  not (G994,G691);
  not (G995,G691);
  not (G996,G691);
  not (G997,G691);
  not (G998,G691);
  not (G999,G691);
  nand (G1000,G639,G890);
  nand (G1001,G636,G891);
  nand (G1002,G645,G892);
  nand (G1003,G642,G893);
  and (G1004,G11,G727);
  nand (G1005,G931,G932);
  nand (G1008,G933,G934);
  nand (G1011,G929,G930);
  and (G1012,G461,G787);
  nand (G1015,G461,G787);
  not (G1016,G731);
  nand (G1017,G916,G734);
  not (G1018,G916);
  and (G1019,G381,G731);
  nand (G1020,G922,G735);
  not (G1021,G922);
  nand (G1022,G11,G727);
  not (G1023,G736);
  not (G1024,G739);
  nand (G1025,G772,G519);
  nand (G1034,G772,G523);
  nand (G1043,G470,G742,G496);
  nand (G1048,G470,G484,G496,G749);
  nand (G1051,G919,G786);
  not (G1052,G919);
  nand (G1053,G925,G791);
  not (G1054,G925);
  not (G1055,G775);
  not (G1056,G781);
  not (G1057,G778);
  and (G1058,G543,G956);
  and (G1059,G21,G957);
  and (G1060,G549,G959);
  and (G1061,G22,G960);
  and (G1062,G10,G961);
  and (G1063,G7,G962);
  and (G1064,G556,G964);
  and (G1065,G543,G965);
  and (G1066,G562,G967);
  and (G1067,G549,G968);
  and (G1068,G13,G970);
  and (G1069,G10,G971);
  and (G1070,G14,G972);
  and (G1071,G556,G973);
  and (G1072,G39,G975);
  and (G1073,G562,G976);
  and (G1074,G26,G810);
  and (G1077,G587,G810);
  and (G1080,G588,G813);
  and (G1083,G589,G813);
  nand (G1086,G745,G749);
  nand (G1089,G519,G749);
  nand (G1092,G470,G742,G684);
  nand (G1095,G484,G492,G745);
  nand (G1104,G484,G745);
  not (G1113,G816);
  not (G1114,G816);
  not (G1115,G816);
  not (G1116,G816);
  not (G1117,G816);
  not (G1118,G816);
  not (G1119,G816);
  not (G1120,G831);
  and (G1121,G831,G594);
  not (G1122,G831);
  and (G1123,G831,G594);
  not (G1124,G831);
  and (G1125,G831,G594);
  not (G1126,G831);
  and (G1127,G831,G594);
  not (G1128,G831);
  and (G1129,G831,G594);
  not (G1130,G831);
  and (G1131,G831,G594);
  not (G1132,G831);
  and (G1133,G831,G594);
  not (G1134,G831);
  and (G1135,G831,G594);
  and (G1136,G691,G856);
  nor (G1137,G7,G856);
  not (G1140,G753);
  and (G1141,G691,G856);
  nor (G1142,G8,G856);
  not (G1145,G753);
  and (G1146,G691,G856);
  nor (G1147,G9,G856);
  not (G1150,G753);
  and (G1151,G691,G856);
  nor (G1152,G10,G856);
  not (G1155,G753);
  and (G1156,G691,G856);
  nor (G1157,G11,G856);
  not (G1160,G769);
  and (G1161,G691,G856);
  nor (G1162,G12,G856);
  not (G1165,G762);
  and (G1166,G691,G856);
  nor (G1167,G13,G856);
  not (G1170,G762);
  and (G1171,G691,G856);
  nor (G1172,G14,G856);
  not (G1175,G762);
  and (G1176,G875,G27);
  nand (G1179,G875,G27);
  and (G1180,G875,G27,G48);
  nand (G1184,G875,G27,G48);
  and (G1189,G875,G27,G48);
  nand (G1193,G875,G27,G48);
  not (G1197,G887);
  nand (G1200,G1000,G1001);
  nand (G1203,G1002,G1003);
  not (G1206,G894);
  nand (G1207,G894,G897);
  not (G1208,G898);
  not (G1209,G901);
  not (G1210,G904);
  not (G1211,G907);
  not (G1212,G910);
  not (G1213,G913);
  nand (G1214,G651,G1018);
  nand (G1215,G657,G1021);
  and (G1216,G935,G739);
  nand (G1217,G654,G1052);
  nand (G1218,G660,G1054);
  and (G1219,G666,G1055);
  or (G1222,G958,G1058,G1059);
  or (G1223,G963,G1062,G1063);
  or (G1224,G966,G1064,G1065);
  or (G1225,G969,G1066,G1067);
  or (G1226,G974,G1070,G1071);
  or (G1227,G977,G1072,G1073);
  and (G1228,G10,G1120);
  and (G1229,G29,G1121);
  and (G1230,G11,G1122);
  and (G1231,G30,G1123);
  and (G1232,G12,G1124);
  and (G1233,G31,G1125);
  and (G1234,G13,G1126);
  and (G1235,G32,G1127);
  and (G1236,G14,G1128);
  and (G1237,G33,G1129);
  and (G1238,G39,G1130);
  and (G1239,G34,G1131);
  and (G1240,G40,G1132);
  and (G1241,G35,G1133);
  and (G1242,G41,G1134);
  and (G1243,G36,G1135);
  not (G1244,G986);
  not (G1249,G986);
  not (G1258,G989);
  not (G1263,G989);
  and (G1272,G7,G686,G1136);
  and (G1275,G8,G686,G1141);
  and (G1278,G9,G686,G1146);
  and (G1281,G10,G686,G1151);
  and (G1284,G11,G708,G1156);
  and (G1287,G12,G708,G1161);
  and (G1290,G13,G708,G1166);
  and (G1293,G14,G708,G1171);
  not (G1296,G939);
  not (G1297,G939);
  not (G1298,G939);
  not (G1299,G939);
  not (G1300,G939);
  not (G1301,G939);
  not (G1302,G939);
  not (G1303,G939);
  nand (G1304,G648,G1206);
  nand (G1305,G901,G1208);
  nand (G1306,G898,G1209);
  nand (G1307,G907,G1210);
  nand (G1308,G904,G1211);
  nand (G1309,G913,G1212);
  nand (G1310,G910,G1213);
  not (G1311,G1200);
  not (G1312,G1203);
  not (G1313,G1025);
  and (G1314,G1025,G1034);
  not (G1315,G1034);
  nand (G1316,G1017,G1214);
  nand (G1317,G1020,G1215);
  and (G1318,G1012,G730,G363,G8);
  not (G1319,G1025);
  and (G1320,G1025,G1034);
  not (G1321,G1034);
  not (G1322,G1025);
  not (G1323,G1034);
  and (G1324,G1025,G1034);
  not (G1325,G1025);
  not (G1326,G1034);
  and (G1327,G1025,G1034);
  not (G1328,G1048);
  not (G1345,G1048);
  nand (G1348,G1051,G1217);
  nand (G1349,G1053,G1218);
  not (G1350,G1043);
  and (G1351,G1043,G775);
  not (G1352,G1043);
  and (G1353,G778,G1043);
  nand (G1354,G805,G1083);
  nand (G1357,G805,G1080);
  nand (G1360,G800,G1083);
  nand (G1363,G800,G1080);
  nand (G1366,G805,G1077);
  nand (G1369,G805,G1074);
  nand (G1372,G800,G1077);
  nand (G1375,G800,G1074);
  not (G1378,G1086);
  not (G1379,G1089);
  and (G1380,G1086,G1089);
  not (G1381,G1092);
  not (G1390,G1092);
  not (G1399,G1104);
  not (G1400,G1104);
  not (G1401,G1104);
  not (G1402,G1104);
  not (G1403,G1095);
  not (G1404,G1095);
  not (G1405,G1095);
  not (G1406,G1095);
  or (G1407,G1228,G978,G1229);
  or (G1408,G1230,G979,G1231);
  or (G1409,G1232,G980,G1233);
  or (G1410,G1234,G981,G1235);
  or (G1411,G1236,G982,G1237);
  or (G1412,G1238,G983,G1239);
  or (G1413,G1240,G984,G1241);
  or (G1414,G1242,G985,G1243);
  and (G1415,G1222,G992);
  and (G1418,G1223,G994);
  and (G1421,G1224,G995);
  and (G1424,G1225,G996);
  and (G1427,G1226,G998);
  and (G1430,G1227,G999);
  not (G1433,G1184);
  and (G1436,G1197,G50);
  nand (G1439,G1197,G50);
  not (G1442,G1005);
  not (G1445,G1008);
  not (G1448,G1005);
  not (G1451,G1008);
  nand (G1454,G1207,G1304);
  nand (G1457,G1305,G1306);
  nand (G1460,G1307,G1308);
  nand (G1463,G1309,G1310);
  nand (G1466,G1203,G1311);
  nand (G1467,G1200,G1312);
  and (G1468,G422,G1314);
  and (G1469,G1316,G397,G1016);
  and (G1470,G451,G1317);
  and (G1471,G1318,G736);
  and (G1472,G434,G1320);
  and (G1473,G1022,G1323);
  and (G1474,G461,G1324);
  and (G1475,G1015,G1326);
  and (G1476,G447,G1327);
  not (G1477,G1348);
  not (G1478,G1349);
  and (G1479,G935,G1350);
  and (G1482,G1011,G1351);
  and (G1485,G363,G1380);
  and (G1486,G1263,G30,G1140);
  and (G1487,G1263,G38,G753);
  and (G1488,G1258,G1407);
  and (G1489,G1263,G31,G1145);
  and (G1490,G1263,G38,G753);
  and (G1491,G1258,G1408);
  and (G1492,G1263,G32,G1150);
  and (G1493,G1263,G38,G753);
  and (G1494,G1258,G1409);
  and (G1495,G1263,G33,G1155);
  and (G1496,G1263,G38,G753);
  and (G1497,G1258,G1410);
  and (G1498,G1249,G34,G1160);
  and (G1499,G1249,G38,G769);
  and (G1500,G1244,G1411);
  and (G1501,G1249,G35,G1165);
  and (G1502,G1249,G38,G762);
  and (G1503,G1244,G1412);
  and (G1504,G1249,G36,G1170);
  and (G1505,G1249,G38,G762);
  and (G1506,G1244,G1413);
  and (G1507,G1249,G37,G1175);
  and (G1508,G1249,G38,G762);
  and (G1509,G1244,G1414);
  not (G1510,G1442);
  not (G1511,G1445);
  not (G1512,G1448);
  not (G1513,G1451);
  nand (G1514,G1466,G1467);
  not (G1517,G1454);
  not (G1518,G1457);
  not (G1519,G1460);
  not (G1520,G1463);
  or (G1521,G1469,G1019);
  not (G1522,G1345);
  and (G1523,G1345,G781);
  and (G1524,G1470,G1352);
  and (G1527,G1477,G793);
  and (G1528,G1478,G797);
  not (G1529,G1354);
  not (G1538,G1357);
  not (G1547,G1360);
  not (G1556,G1363);
  not (G1565,G1366);
  not (G1574,G1369);
  not (G1583,G1372);
  not (G1592,G1375);
  not (G1601,G1354);
  not (G1610,G1357);
  not (G1619,G1360);
  not (G1628,G1363);
  not (G1637,G1366);
  not (G1646,G1369);
  not (G1655,G1372);
  not (G1664,G1375);
  not (G1673,G1381);
  and (G1674,G1381,G1104);
  not (G1675,G1381);
  and (G1676,G1381,G1104);
  not (G1677,G1381);
  and (G1678,G1381,G1104);
  not (G1679,G1381);
  and (G1680,G1381,G1104);
  not (G1681,G1390);
  and (G1682,G1390,G1095);
  not (G1683,G1390);
  and (G1684,G1390,G1095);
  not (G1685,G1390);
  and (G1686,G1390,G1095);
  not (G1687,G1390);
  and (G1688,G1390,G1095);
  or (G1689,G1415,G1137,G1272);
  nor (G1693,G1415,G1137,G1272);
  or (G1697,G1486,G1487,G1488);
  or (G1700,G1489,G1490,G1491);
  or (G1703,G1418,G1147,G1278);
  nor (G1707,G1418,G1147,G1278);
  or (G1711,G1492,G1493,G1494);
  or (G1714,G1421,G1152,G1281);
  nor (G1718,G1421,G1152,G1281);
  or (G1722,G1495,G1496,G1497);
  or (G1725,G1424,G1157,G1284);
  nor (G1729,G1424,G1157,G1284);
  or (G1733,G1498,G1499,G1500);
  or (G1738,G1501,G1502,G1503);
  or (G1743,G1427,G1167,G1290);
  nor (G1747,G1427,G1167,G1290);
  or (G1751,G1504,G1505,G1506);
  or (G1756,G1430,G1172,G1293);
  nor (G1760,G1430,G1172,G1293);
  or (G1764,G1507,G1508,G1509);
  not (G1769,G1433);
  not (G1770,G1328);
  and (G1771,G939,G1328);
  not (G1772,G1328);
  and (G1773,G939,G1328);
  not (G1774,G1328);
  and (G1775,G939,G1328);
  not (G1776,G1328);
  and (G1777,G939,G1328);
  not (G1778,G1328);
  and (G1779,G939,G1328);
  not (G1780,G1328);
  and (G1781,G939,G1328);
  not (G1782,G1328);
  and (G1783,G939,G1328);
  not (G1784,G1328);
  and (G1785,G939,G1328);
  or (G1786,G1479,G1219,G1482);
  nor (G1787,G1479,G1219,G1482);
  nand (G1788,G1445,G1510);
  nand (G1789,G1442,G1511);
  nand (G1790,G1451,G1512);
  nand (G1791,G1448,G1513);
  nand (G1792,G1457,G1517);
  nand (G1793,G1454,G1518);
  nand (G1794,G1463,G1519);
  nand (G1795,G1460,G1520);
  and (G1796,G935,G1522);
  and (G1799,G1012,G1523);
  and (G1802,G1521,G1057);
  or (G1805,G1527,G1060,G1061);
  or (G1806,G1528,G1068,G1069);
  and (G1807,G363,G1674);
  and (G1808,G377,G1676);
  and (G1809,G384,G1678);
  and (G1810,G400,G1680);
  not (G1811,G1787);
  nand (G1812,G1788,G1789);
  nand (G1813,G1790,G1791);
  not (G1816,G1514);
  nand (G1819,G1792,G1793);
  nand (G1823,G1794,G1795);
  and (G1826,G1514,G1313);
  not (G1827,G1529);
  not (G1828,G1538);
  not (G1829,G1547);
  not (G1830,G1556);
  not (G1831,G1565);
  not (G1832,G1574);
  not (G1833,G1583);
  not (G1834,G1592);
  not (G1835,G1529);
  not (G1836,G1538);
  not (G1837,G1547);
  not (G1838,G1556);
  not (G1839,G1565);
  not (G1840,G1574);
  not (G1841,G1583);
  not (G1842,G1592);
  not (G1843,G1529);
  not (G1844,G1538);
  not (G1845,G1547);
  not (G1846,G1556);
  not (G1847,G1565);
  not (G1848,G1574);
  not (G1849,G1583);
  not (G1850,G1592);
  not (G1851,G1529);
  not (G1852,G1538);
  not (G1853,G1547);
  not (G1854,G1556);
  not (G1855,G1565);
  not (G1856,G1574);
  not (G1857,G1583);
  not (G1858,G1592);
  not (G1859,G1529);
  not (G1860,G1538);
  not (G1861,G1547);
  not (G1862,G1556);
  not (G1863,G1565);
  not (G1864,G1574);
  not (G1865,G1583);
  not (G1866,G1592);
  not (G1867,G1529);
  not (G1868,G1538);
  not (G1869,G1547);
  not (G1870,G1556);
  not (G1871,G1565);
  not (G1872,G1574);
  not (G1873,G1583);
  not (G1874,G1592);
  not (G1875,G1529);
  not (G1876,G1538);
  not (G1877,G1547);
  not (G1878,G1556);
  not (G1879,G1565);
  not (G1880,G1574);
  not (G1881,G1583);
  not (G1882,G1592);
  not (G1883,G1529);
  not (G1884,G1538);
  not (G1885,G1547);
  not (G1886,G1556);
  not (G1887,G1565);
  not (G1888,G1574);
  not (G1889,G1583);
  not (G1890,G1592);
  not (G1891,G1601);
  not (G1892,G1610);
  not (G1893,G1619);
  not (G1894,G1628);
  not (G1895,G1637);
  not (G1896,G1646);
  not (G1897,G1655);
  not (G1898,G1664);
  not (G1899,G1601);
  not (G1900,G1610);
  not (G1901,G1619);
  not (G1902,G1628);
  not (G1903,G1637);
  not (G1904,G1646);
  not (G1905,G1655);
  not (G1906,G1664);
  not (G1907,G1601);
  not (G1908,G1610);
  not (G1909,G1619);
  not (G1910,G1628);
  not (G1911,G1637);
  not (G1912,G1646);
  not (G1913,G1655);
  not (G1914,G1664);
  not (G1915,G1601);
  not (G1916,G1610);
  not (G1917,G1619);
  not (G1918,G1628);
  not (G1919,G1637);
  not (G1920,G1646);
  not (G1921,G1655);
  not (G1922,G1664);
  not (G1923,G1601);
  not (G1924,G1610);
  not (G1925,G1619);
  not (G1926,G1628);
  not (G1927,G1637);
  not (G1928,G1646);
  not (G1929,G1655);
  not (G1930,G1664);
  not (G1931,G1601);
  not (G1932,G1610);
  not (G1933,G1619);
  not (G1934,G1628);
  not (G1935,G1637);
  not (G1936,G1646);
  not (G1937,G1655);
  not (G1938,G1664);
  not (G1939,G1601);
  not (G1940,G1610);
  not (G1941,G1619);
  not (G1942,G1628);
  not (G1943,G1637);
  not (G1944,G1646);
  not (G1945,G1655);
  not (G1946,G1664);
  not (G1947,G1601);
  not (G1948,G1610);
  not (G1949,G1619);
  not (G1950,G1628);
  not (G1951,G1637);
  not (G1952,G1646);
  not (G1953,G1655);
  not (G1954,G1664);
  not (G1955,G1697);
  not (G1958,G1697);
  not (G1961,G1693);
  and (G1962,G1805,G993);
  not (G1965,G1700);
  not (G1968,G1700);
  not (G1971,G1711);
  not (G1974,G1711);
  not (G1977,G1707);
  not (G1978,G1722);
  not (G1981,G1722);
  not (G1984,G1718);
  not (G1985,G1733);
  not (G1988,G1733);
  not (G1991,G1729);
  and (G1992,G1806,G997);
  not (G1995,G1738);
  not (G1998,G1738);
  not (G2001,G1751);
  not (G2004,G1751);
  not (G2007,G1747);
  not (G2008,G1764);
  not (G2011,G1764);
  not (G2014,G1760);
  and (G2015,G1176,G1689);
  and (G2018,G1180,G1703);
  and (G2021,G1180,G1714);
  and (G2024,G1180,G1725);
  and (G2027,G1189,G1743);
  and (G2030,G1189,G1756);
  not (G2033,G1733);
  not (G2034,G1738);
  not (G2035,G1751);
  not (G2036,G1764);
  and (G2037,G1733,G1738,G1751,G1764,G882);
  not (G2038,G1812);
  or (G2039,G1826,G1315,G1468);
  and (G2040,G15,G1827);
  and (G2041,G22,G1828);
  and (G2042,G21,G1829);
  and (G2043,G20,G1830);
  and (G2044,G19,G1831);
  and (G2045,G18,G1832);
  and (G2046,G17,G1833);
  and (G2047,G16,G1834);
  and (G2048,G16,G1835);
  and (G2049,G353,G1836);
  and (G2050,G22,G1837);
  and (G2051,G21,G1838);
  and (G2052,G20,G1839);
  and (G2053,G19,G1840);
  and (G2054,G18,G1841);
  and (G2055,G17,G1842);
  and (G2056,G17,G1843);
  and (G2057,G368,G1844);
  and (G2058,G353,G1845);
  and (G2059,G22,G1846);
  and (G2060,G21,G1847);
  and (G2061,G20,G1848);
  and (G2062,G19,G1849);
  and (G2063,G18,G1850);
  and (G2064,G18,G1851);
  and (G2065,G388,G1852);
  and (G2066,G368,G1853);
  and (G2067,G353,G1854);
  and (G2068,G22,G1855);
  and (G2069,G21,G1856);
  and (G2070,G20,G1857);
  and (G2071,G19,G1858);
  and (G2072,G19,G1859);
  and (G2073,G404,G1860);
  and (G2074,G388,G1861);
  and (G2075,G368,G1862);
  and (G2076,G353,G1863);
  and (G2077,G22,G1864);
  and (G2078,G21,G1865);
  and (G2079,G20,G1866);
  and (G2080,G20,G1867);
  and (G2081,G413,G1868);
  and (G2082,G404,G1869);
  and (G2083,G388,G1870);
  and (G2084,G368,G1871);
  and (G2085,G353,G1872);
  and (G2086,G22,G1873);
  and (G2087,G21,G1874);
  and (G2088,G21,G1875);
  and (G2089,G425,G1876);
  and (G2090,G413,G1877);
  and (G2091,G404,G1878);
  and (G2092,G388,G1879);
  and (G2093,G368,G1880);
  and (G2094,G353,G1881);
  and (G2095,G22,G1882);
  and (G2096,G22,G1883);
  and (G2097,G438,G1884);
  and (G2098,G425,G1885);
  and (G2099,G413,G1886);
  and (G2100,G404,G1887);
  and (G2101,G388,G1888);
  and (G2102,G368,G1889);
  and (G2103,G353,G1890);
  and (G2104,G39,G1891);
  and (G2105,G368,G1892);
  and (G2106,G388,G1893);
  and (G2107,G404,G1894);
  and (G2108,G413,G1895);
  and (G2109,G425,G1896);
  and (G2110,G438,G1897);
  and (G2111,G451,G1898);
  and (G2112,G40,G1899);
  and (G2113,G388,G1900);
  and (G2114,G404,G1901);
  and (G2115,G413,G1902);
  and (G2116,G425,G1903);
  and (G2117,G438,G1904);
  and (G2118,G451,G1905);
  and (G2119,G39,G1906);
  and (G2120,G41,G1907);
  and (G2121,G404,G1908);
  and (G2122,G413,G1909);
  and (G2123,G425,G1910);
  and (G2124,G438,G1911);
  and (G2125,G451,G1912);
  and (G2126,G39,G1913);
  and (G2127,G40,G1914);
  and (G2128,G42,G1915);
  and (G2129,G413,G1916);
  and (G2130,G425,G1917);
  and (G2131,G438,G1918);
  and (G2132,G451,G1919);
  and (G2133,G39,G1920);
  and (G2134,G40,G1921);
  and (G2135,G41,G1922);
  and (G2136,G43,G1923);
  and (G2137,G425,G1924);
  and (G2138,G438,G1925);
  and (G2139,G451,G1926);
  and (G2140,G39,G1927);
  and (G2141,G40,G1928);
  and (G2142,G41,G1929);
  and (G2143,G42,G1930);
  and (G2144,G44,G1931);
  and (G2145,G438,G1932);
  and (G2146,G451,G1933);
  and (G2147,G39,G1934);
  and (G2148,G40,G1935);
  and (G2149,G41,G1936);
  and (G2150,G42,G1937);
  and (G2151,G43,G1938);
  and (G2152,G45,G1939);
  and (G2153,G451,G1940);
  and (G2154,G39,G1941);
  and (G2155,G40,G1942);
  and (G2156,G41,G1943);
  and (G2157,G42,G1944);
  and (G2158,G43,G1945);
  and (G2159,G44,G1946);
  and (G2160,G46,G1947);
  and (G2161,G39,G1948);
  and (G2162,G40,G1949);
  and (G2163,G41,G1950);
  and (G2164,G42,G1951);
  and (G2165,G43,G1952);
  and (G2166,G44,G1953);
  and (G2167,G45,G1954);
  and (G2168,G2033,G2034,G2035,G2036,G615);
  not (G2169,G1823);
  and (G2172,G2038,G1023);
  and (G2173,G1823,G1319);
  and (G2174,G1819,G1024);
  nor (G2175,G2040,G2041,G2042,G2043,G2044,G2045,G2046,G2047);
  nor (G2176,G2048,G2049,G2050,G2051,G2052,G2053,G2054,G2055);
  nor (G2177,G2056,G2057,G2058,G2059,G2060,G2061,G2062,G2063);
  nor (G2178,G2064,G2065,G2066,G2067,G2068,G2069,G2070,G2071);
  nor (G2179,G2072,G2073,G2074,G2075,G2076,G2077,G2078,G2079);
  nor (G2180,G2080,G2081,G2082,G2083,G2084,G2085,G2086,G2087);
  nor (G2181,G2088,G2089,G2090,G2091,G2092,G2093,G2094,G2095);
  nor (G2182,G2096,G2097,G2098,G2099,G2100,G2101,G2102,G2103);
  nor (G2183,G2104,G2105,G2106,G2107,G2108,G2109,G2110,G2111);
  nor (G2184,G2112,G2113,G2114,G2115,G2116,G2117,G2118,G2119);
  nor (G2185,G2120,G2121,G2122,G2123,G2124,G2125,G2126,G2127);
  nor (G2186,G2128,G2129,G2130,G2131,G2132,G2133,G2134,G2135);
  nor (G2187,G2136,G2137,G2138,G2139,G2140,G2141,G2142,G2143);
  nor (G2188,G2144,G2145,G2146,G2147,G2148,G2149,G2150,G2151);
  nor (G2189,G2152,G2153,G2154,G2155,G2156,G2157,G2158,G2159);
  nor (G2190,G2160,G2161,G2162,G2163,G2164,G2165,G2166,G2167);
  and (G2191,G2039,G1682);
  and (G2192,G23,G1689,G1955);
  and (G2195,G24,G1689,G1958);
  and (G2198,G25,G1693,G1958);
  and (G2199,G26,G1693,G1955);
  or (G2200,G1962,G1142,G1275);
  nor (G2204,G1962,G1142,G1275);
  and (G2208,G23,G1703,G1971);
  and (G2211,G24,G1703,G1974);
  and (G2214,G25,G1707,G1974);
  and (G2215,G26,G1707,G1971);
  and (G2216,G23,G1714,G1978);
  and (G2219,G24,G1714,G1981);
  and (G2222,G25,G1718,G1981);
  and (G2223,G26,G1718,G1978);
  and (G2224,G23,G1725,G1985);
  and (G2227,G24,G1725,G1988);
  and (G2230,G25,G1729,G1988);
  and (G2231,G26,G1729,G1985);
  or (G2232,G1992,G1162,G1287);
  nor (G2236,G1992,G1162,G1287);
  and (G2240,G23,G1743,G2001);
  and (G2243,G24,G1743,G2004);
  and (G2246,G25,G1747,G2004);
  and (G2247,G26,G1747,G2001);
  and (G2248,G23,G1756,G2008);
  and (G2251,G24,G1756,G2011);
  and (G2254,G25,G1760,G2011);
  and (G2255,G26,G1760,G2008);
  or (G2256,G2037,G2168);
  not (G2257,G1813);
  not (G2260,G1816);
  not (G2263,G1813);
  not (G2266,G1816);
  not (G2269,G1819);
  not (G2272,G1819);
  not (G2275,G2015);
  not (G2278,G2015);
  not (G2281,G2018);
  not (G2284,G2018);
  not (G2287,G2021);
  not (G2290,G2021);
  not (G2293,G2024);
  not (G2296,G2024);
  not (G2299,G2027);
  not (G2302,G2027);
  not (G2305,G2030);
  not (G2308,G2030);
  nor (G2311,G2172,G1471);
  or (G2312,G2173,G1321,G1472);
  nor (G2313,G2174,G1216);
  and (G2314,G2175,G1378);
  and (G2315,G2183,G1379);
  and (G2316,G2176,G1113);
  and (G2317,G2184,G816);
  and (G2318,G2177,G1114);
  and (G2319,G2185,G816);
  and (G2320,G2178,G1115);
  and (G2321,G2186,G816);
  and (G2322,G2179,G1116);
  and (G2323,G2187,G816);
  and (G2324,G2180,G1117);
  and (G2325,G2188,G816);
  and (G2326,G2181,G1118);
  and (G2327,G2189,G816);
  and (G2328,G2182,G1119);
  and (G2329,G2190,G816);
  or (G2330,G2198,G2199,G1961);
  or (G2331,G2214,G2215,G1977);
  or (G2332,G2222,G2223,G1984);
  or (G2333,G2230,G2231,G1991);
  or (G2334,G2246,G2247,G2007);
  or (G2335,G2254,G2255,G2014);
  and (G2336,G2256,G1769);
  not (G2337,G2263);
  not (G2338,G2266);
  not (G2339,G2272);
  not (G2340,G2269);
  not (G2341,G2257);
  not (G2342,G2260);
  and (G2343,G2313,G1322);
  and (G2344,G2311,G1325);
  or (G2345,G2314,G2315,G1485);
  or (G2346,G2316,G2317);
  or (G2347,G2318,G2319);
  or (G2348,G2320,G2321);
  or (G2349,G2322,G2323);
  or (G2350,G2324,G2325);
  or (G2351,G2326,G2327);
  or (G2352,G2328,G2329);
  and (G2353,G2312,G1684);
  or (G2354,G2192,G2195);
  nor (G2355,G2192,G2195);
  and (G2356,G23,G2200,G1965);
  and (G2359,G24,G2200,G1968);
  and (G2362,G25,G2204,G1968);
  and (G2363,G26,G2204,G1965);
  not (G2364,G2204);
  or (G2365,G2208,G2211);
  nor (G2368,G2208,G2211);
  or (G2369,G2216,G2219);
  nor (G2372,G2216,G2219);
  or (G2373,G2224,G2227);
  nor (G2374,G2224,G2227);
  and (G2375,G23,G2232,G1995);
  and (G2378,G24,G2232,G1998);
  and (G2381,G25,G2236,G1998);
  and (G2382,G26,G2236,G1995);
  not (G2383,G2236);
  or (G2384,G2240,G2243);
  nor (G2387,G2240,G2243);
  or (G2388,G2248,G2251);
  nor (G2391,G2248,G2251);
  not (G2392,G2278);
  and (G2393,G1176,G2200);
  not (G2396,G2281);
  not (G2397,G2284);
  not (G2398,G2287);
  not (G2399,G2290);
  not (G2400,G2296);
  and (G2401,G1189,G2232);
  not (G2404,G2302);
  not (G2405,G2305);
  not (G2406,G2308);
  not (G2407,G2299);
  not (G2408,G2169);
  not (G2411,G2169);
  not (G2414,G2275);
  not (G2415,G2293);
  nand (G2416,G2260,G2341);
  nand (G2417,G2257,G2342);
  nand (G2418,G2266,G2337);
  nand (G2419,G2263,G2338);
  or (G2420,G2343,G1473,G1474);
  or (G2421,G2344,G1475,G1476);
  and (G2422,G2345,G1673);
  and (G2423,G2346,G1675);
  and (G2424,G2347,G1677);
  and (G2425,G2348,G1679);
  and (G2426,G2349,G1681);
  and (G2427,G2350,G1683);
  and (G2428,G2351,G1685);
  and (G2429,G2352,G1687);
  and (G2430,G2355,G2330);
  or (G2436,G2362,G2363,G2364);
  and (G2437,G2368,G2331);
  and (G2441,G2372,G2332);
  and (G2444,G2374,G2333);
  or (G2450,G2381,G2382,G2383);
  and (G2451,G2387,G2334);
  and (G2455,G2391,G2335);
  not (G2458,G2354);
  not (G2459,G2373);
  nand (G2460,G2416,G2417);
  nand (G2461,G2418,G2419);
  nand (G2462,G2411,G2339);
  not (G2463,G2411);
  nand (G2464,G2408,G2340);
  not (G2465,G2408);
  and (G2466,G2421,G1686);
  and (G2467,G2420,G1688);
  or (G2468,G2356,G2359);
  nor (G2471,G2356,G2359);
  or (G2472,G2375,G2378);
  nor (G2475,G2375,G2378);
  and (G2476,G2365,G1184);
  and (G2479,G2369,G1184);
  and (G2482,G2384,G1193);
  and (G2485,G2388,G1193);
  not (G2488,G2393);
  not (G2491,G2393);
  not (G2494,G2401);
  not (G2497,G2401);
  nand (G2500,G2272,G2463);
  nand (G2501,G2269,G2465);
  and (G2502,G2471,G2436);
  and (G2507,G2475,G2450);
  not (G2512,G2430);
  not (G2515,G2437);
  not (G2518,G2441);
  not (G2521,G2444);
  not (G2524,G2451);
  not (G2527,G2455);
  nand (G2530,G2462,G2500);
  nand (G2531,G2464,G2501);
  nand (G2532,G2430,G2468);
  nand (G2533,G2444,G2472);
  not (G2534,G2488);
  not (G2535,G2491);
  not (G2536,G2497);
  not (G2537,G2494);
  and (G2538,G2468,G1179);
  not (G2539,G2479);
  and (G2542,G2472,G1184);
  not (G2543,G2485);
  not (G2546,G2476);
  not (G2547,G2485);
  not (G2550,G2530);
  not (G2551,G2531);
  and (G2552,G2430,G2502,G2437,G2441);
  nand (G2556,G2430,G2502,G2365);
  nand (G2557,G2369,G2502,G2437,G2430);
  and (G2558,G2444,G2507,G2451,G2455);
  nand (G2561,G2444,G2507,G2384);
  nand (G2562,G2388,G2507,G2451,G2444);
  not (G2563,G2502);
  not (G2566,G2507);
  not (G2569,G2538);
  not (G2570,G2542);
  not (G2571,G2512);
  not (G2574,G2512);
  not (G2577,G2515);
  not (G2580,G2515);
  not (G2583,G2518);
  not (G2586,G2518);
  not (G2589,G2521);
  not (G2592,G2521);
  not (G2595,G2524);
  not (G2598,G2524);
  not (G2601,G2527);
  not (G2604,G2527);
  nand (G2607,G2458,G2532,G2556,G2557);
  nand (G2610,G2459,G2533,G2561,G2562);
  not (G2613,G2547);
  nand (G2614,G2574,G2392);
  nand (G2615,G2580,G2397);
  nand (G2616,G2586,G2399);
  nand (G2617,G2592,G2400);
  nand (G2618,G2598,G2404);
  nand (G2619,G2604,G2406);
  not (G2620,G2552);
  not (G2623,G2574);
  not (G2624,G2577);
  nand (G2625,G2577,G2396);
  not (G2626,G2580);
  not (G2627,G2583);
  nand (G2628,G2583,G2398);
  not (G2629,G2586);
  not (G2630,G2592);
  not (G2631,G2598);
  not (G2632,G2601);
  nand (G2633,G2601,G2405);
  not (G2634,G2604);
  not (G2635,G2595);
  nand (G2636,G2595,G2407);
  and (G2637,G2558,G1433);
  not (G2638,G2571);
  nand (G2639,G2571,G2414);
  not (G2640,G2563);
  not (G2643,G2563);
  not (G2646,G2589);
  nand (G2647,G2589,G2415);
  not (G2648,G2566);
  not (G2651,G2566);
  nand (G2654,G2552,G2610);
  not (G2655,G2607);
  nand (G2656,G2278,G2623);
  nand (G2657,G2284,G2626);
  nand (G2658,G2290,G2629);
  nand (G2659,G2296,G2630);
  nand (G2660,G2302,G2631);
  nand (G2661,G2308,G2634);
  nand (G2662,G2281,G2624);
  nand (G2663,G2287,G2627);
  nand (G2664,G2305,G2632);
  nand (G2665,G2299,G2635);
  and (G2666,G2610,G1193);
  or (G2669,G2336,G2637);
  nand (G2673,G2275,G2638);
  nand (G2674,G2293,G2646);
  and (G2675,G2654,G2655);
  nand (G2676,G2656,G2614);
  nand (G2677,G2643,G2535);
  nand (G2678,G2657,G2615);
  nand (G2679,G2658,G2616);
  nand (G2680,G2659,G2617);
  nand (G2681,G2651,G2536);
  nand (G2682,G2660,G2618);
  nand (G2683,G2661,G2619);
  not (G2684,G2640);
  nand (G2685,G2640,G2534);
  not (G2686,G2643);
  nand (G2687,G2662,G2625);
  nand (G2690,G2663,G2628);
  not (G2693,G2651);
  nand (G2694,G2664,G2633);
  not (G2697,G2648);
  nand (G2698,G2648,G2537);
  nand (G2699,G2665,G2636);
  nand (G2705,G2673,G2639);
  nand (G2708,G2674,G2647);
  not (G2711,G2676);
  nand (G2712,G2491,G2686);
  not (G2713,G2678);
  not (G2714,G2679);
  not (G2715,G2680);
  nand (G2716,G2497,G2693);
  not (G2717,G2682);
  not (G2718,G2683);
  nand (G2719,G2488,G2684);
  nand (G2720,G2494,G2697);
  not (G2721,G2666);
  not (G2728,G2669);
  not (G2733,G2666);
  and (G2736,G47,G2669);
  and (G2739,G2711,G1399);
  nand (G2740,G2712,G2677);
  and (G2741,G2713,G1401);
  and (G2742,G2714,G1402);
  and (G2743,G2715,G1403);
  nand (G2744,G2716,G2681);
  and (G2745,G2717,G1405);
  and (G2746,G2718,G1406);
  nand (G2747,G2719,G2685);
  not (G2750,G2687);
  not (G2753,G2687);
  not (G2759,G2690);
  not (G2763,G2690);
  nand (G2768,G2720,G2698);
  not (G2773,G2694);
  and (G2778,G2699,G2543);
  not (G2779,G2705);
  not (G2780,G2708);
  and (G2781,G47,G2694);
  not (G2784,G2699);
  nor (G2787,G2422,G2739,G1807);
  not (G2788,G2740);
  nor (G2789,G2424,G2741,G1809);
  nor (G2790,G2425,G2742,G1810);
  nor (G2791,G2426,G2743,G2191);
  not (G2792,G2744);
  nor (G2793,G2428,G2745,G2466);
  nor (G2794,G2429,G2746,G2467);
  and (G2795,G2721,G2620);
  and (G2796,G2728,G2620);
  or (G2799,G2482,G2778);
  not (G2803,G2736);
  not (G2804,G2721);
  not (G2805,G2721);
  not (G2808,G2733);
  and (G2809,G2788,G1400);
  and (G2810,G2792,G1404);
  not (G2811,G2747);
  or (G2816,G2607,G2795);
  and (G2820,G2728,G2763,G2753);
  and (G2821,G2728,G2759);
  and (G2822,G2773,G2699,G2768);
  and (G2823,G2773,G2699);
  and (G2826,G2721,G2759);
  nand (G2827,G2753,G2539);
  nand (G2828,G2753,G2763,G2721);
  nand (G2829,G2768,G2482);
  nand (G2830,G2768,G2699,G2543);
  nand (G2831,G2784,G2613);
  not (G2832,G2784);
  and (G2833,G47,G2669,G2804);
  and (G2836,G2787,G1771);
  and (G2839,G2789,G1775);
  and (G2842,G2790,G1777);
  and (G2845,G2791,G1779);
  and (G2848,G2793,G1783);
  and (G2851,G2794,G1785);
  not (G2854,G2747);
  not (G2857,G2753);
  not (G2860,G2759);
  not (G2863,G2768);
  not (G2866,G2781);
  not (G2869,G2781);
  and (G2872,G2773,G2773);
  nor (G2875,G2423,G2809,G1808);
  nor (G2876,G2427,G2810,G2353);
  and (G2877,G47,G2821);
  and (G2880,G47,G2822);
  nand (G2883,G2547,G2832);
  not (G2884,G2799);
  not (G2887,G2796);
  nand (G2890,G2546,G2827,G2828);
  or (G2893,G2479,G2826);
  nand (G2896,G2570,G2829,G2830);
  not (G2899,G2799);
  and (G2902,G47,G2820);
  or (G2905,G2833,G2805);
  and (G2906,G2728,G2811,G2753,G2763);
  nand (G2909,G2811,G2476);
  nand (G2910,G2811,G2750,G2539);
  nand (G2911,G2811,G2750,G2763,G2721);
  not (G2912,G2857);
  nand (G2913,G2831,G2883);
  not (G2916,G2866);
  not (G2917,G2869);
  nand (G2918,G2872,G883);
  not (G2919,G2872);
  not (G2920,G2816);
  nor (G2923,G2833,G2805);
  and (G2926,G2875,G1773);
  and (G2929,G2876,G1781);
  not (G2932,G2816);
  not (G2935,G2854);
  not (G2936,G2860);
  nand (G2937,G2860,G2808);
  not (G2938,G2863);
  and (G2939,G47,G2823);
  not (G2942,G2884);
  and (G2943,G2799,G2884);
  and (G2944,G2905,G1056);
  nand (G2947,G2569,G2909,G2910,G2911);
  not (G2950,G2887);
  not (G2951,G2902);
  not (G2952,G2893);
  nand (G2953,G2893,G2912);
  not (G2954,G2896);
  nand (G2955,G2896,G2780);
  nand (G2956,G663,G2919);
  not (G2957,G2890);
  nand (G2958,G2890,G2935);
  nand (G2959,G2733,G2936);
  not (G2960,G2899);
  nand (G2961,G2899,G2938);
  not (G2962,G2877);
  not (G2965,G2877);
  not (G2968,G2880);
  not (G2971,G2880);
  and (G2974,G47,G2823,G2942);
  and (G2975,G47,G2906);
  nand (G2978,G2857,G2952);
  nand (G2979,G2708,G2954);
  not (G2980,G2939);
  nand (G2981,G2918,G2956);
  not (G2984,G2920);
  and (G2985,G2816,G2920);
  not (G2986,G2923);
  not (G2990,G2932);
  not (G2991,G2906);
  nand (G2994,G2854,G2957);
  nand (G2995,G2863,G2960);
  nand (G2996,G2937,G2959);
  not (G2999,G2913);
  not (G3002,G2913);
  or (G3005,G1796,G2944,G1799);
  nor (G3006,G1796,G2944,G1799);
  nand (G3007,G2978,G2953);
  not (G3010,G2962);
  not (G3011,G2965);
  nand (G3012,G2979,G2955);
  not (G3015,G2968);
  not (G3016,G2971);
  and (G3017,G47,G2796,G2984);
  not (G3018,G2947);
  not (G3021,G2947);
  nand (G3024,G2994,G2958);
  nand (G3027,G2995,G2961);
  not (G3030,G3006);
  nand (G3031,G2991,G2950);
  not (G3032,G2991);
  not (G3033,G2996);
  nand (G3034,G2996,G2803);
  not (G3035,G2999);
  nand (G3036,G2999,G2916);
  not (G3037,G3002);
  nand (G3038,G3002,G2917);
  nor (G3039,G3017,G2985);
  and (G3042,G2981,G1303);
  and (G3045,G2981,G1784);
  not (G3048,G2975);
  not (G3051,G2975);
  not (G3054,G2986);
  nand (G3057,G2887,G3032);
  not (G3058,G3021);
  nand (G3059,G3021,G2779);
  not (G3060,G3024);
  nand (G3061,G3024,G2951);
  nand (G3062,G2736,G3033);
  not (G3063,G3027);
  nand (G3064,G3027,G2980);
  nand (G3065,G2866,G3035);
  nand (G3066,G2869,G3037);
  not (G3067,G3018);
  nand (G3068,G3018,G2990);
  not (G3069,G3007);
  not (G3072,G3007);
  not (G3075,G3012);
  not (G3078,G3012);
  nand (G3081,G3031,G3057);
  nand (G3082,G2705,G3058);
  not (G3083,G3048);
  not (G3084,G3051);
  nand (G3085,G2902,G3060);
  nand (G3086,G3062,G3034);
  nand (G3089,G2939,G3063);
  nand (G3090,G3065,G3036);
  nand (G3094,G3066,G3038);
  not (G3095,G3039);
  not (G3099,G3054);
  or (G3100,G3042,G3045,G2851);
  nor (G3103,G3042,G3045,G2851);
  nand (G3106,G2932,G3067);
  nand (G3107,G3082,G3059);
  nand (G3110,G3085,G3061);
  not (G3114,G3069);
  nand (G3115,G3069,G3010);
  not (G3116,G3072);
  nand (G3117,G3072,G3011);
  not (G3118,G3075);
  nand (G3119,G3075,G3015);
  not (G3120,G3078);
  nand (G3121,G3078,G3016);
  nand (G3122,G3089,G3064);
  nand (G3126,G3106,G3068);
  and (G3129,G47,G3081);
  not (G3132,G3094);
  not (G3135,G3103);
  nand (G3136,G2962,G3114);
  nand (G3137,G2965,G3116);
  nand (G3138,G2968,G3118);
  nand (G3139,G2971,G3120);
  and (G3140,G3086,G1299);
  and (G3143,G3086,G1776);
  and (G3146,G3090,G1302);
  not (G3149,G3095);
  and (G3152,G3090,G2923);
  not (G3155,G3100);
  not (G3158,G3126);
  not (G3159,G3129);
  nand (G3160,G3136,G3115);
  nand (G3164,G3137,G3117);
  nand (G3165,G3138,G3119);
  nand (G3168,G3139,G3121);
  nand (G3169,G3132,G3099);
  not (G3170,G3132);
  and (G3171,G3110,G1297);
  and (G3174,G3122,G1301);
  not (G3177,G3107);
  not (G3180,G3107);
  not (G3183,G3110);
  not (G3186,G3122);
  nand (G3189,G3129,G3158);
  nand (G3190,G3126,G3159);
  not (G3191,G3168);
  not (G3192,G3149);
  not (G3193,G3152);
  nand (G3194,G3054,G3170);
  or (G3195,G3140,G3143,G2842);
  nor (G3199,G3140,G3143,G2842);
  not (G3202,G3155);
  not (G3203,G3164);
  nand (G3206,G3189,G3190);
  not (G3207,G3177);
  nand (G3208,G3177,G3083);
  not (G3209,G3180);
  nand (G3210,G3180,G3084);
  nor (G3211,G3191,G2986);
  and (G3212,G3090,G3122,G3165,G2986);
  not (G3213,G3183);
  not (G3214,G3186);
  nand (G3215,G3186,G3193);
  nand (G3216,G3194,G3169);
  and (G3217,G3160,G1298);
  and (G3220,G3165,G1300);
  and (G3223,G3160,G3039);
  not (G3226,G3199);
  and (G3227,G3206,G1353);
  nand (G3230,G3048,G3207);
  nand (G3231,G3051,G3209);
  or (G3232,G3211,G3212);
  nand (G3233,G3203,G3192);
  not (G3234,G3203);
  nand (G3235,G3152,G3214);
  not (G3236,G3216);
  not (G3237,G3195);
  not (G3240,G3195);
  nand (G3243,G3230,G3208);
  nand (G3246,G3231,G3210);
  nand (G3247,G3223,G3213);
  not (G3248,G3223);
  nand (G3249,G3149,G3234);
  nand (G3250,G3235,G3215);
  and (G3251,G3232,G1778);
  and (G3254,G3236,G1782);
  or (G3257,G1802,G1524,G3227);
  nor (G3258,G1802,G1524,G3227);
  not (G3259,G3246);
  nand (G3260,G3183,G3248);
  nand (G3261,G3249,G3233);
  and (G3262,G3250,G1780);
  not (G3265,G3237);
  not (G3266,G3240);
  not (G3267,G3258);
  nor (G3268,G3259,G3095);
  and (G3269,G3160,G3110,G3243,G3095);
  nand (G3270,G3247,G3260);
  not (G3271,G3261);
  and (G3272,G3243,G1296);
  or (G3275,G3220,G3251,G2845);
  nor (G3278,G3220,G3251,G2845);
  or (G3281,G3146,G3254,G2848);
  nor (G3284,G3146,G3254,G2848);
  or (G3287,G3268,G3269);
  and (G3288,G3270,G1772);
  and (G3291,G3271,G1774);
  or (G3294,G3174,G3262,G2929);
  nor (G3297,G3174,G3262,G2929);
  not (G3300,G3278);
  not (G3301,G3284);
  and (G3302,G3287,G1770);
  not (G3305,G3281);
  not (G3308,G3275);
  not (G3311,G3297);
  or (G3312,G3171,G3288,G2926);
  nor (G3317,G3171,G3288,G2926);
  or (G3320,G3217,G3291,G2839);
  nor (G3323,G3217,G3291,G2839);
  and (G3326,G3103,G3284,G3297,G3278);
  not (G3329,G3294);
  or (G3332,G3272,G3302,G2836);
  nor (G3337,G3272,G3302,G2836);
  nand (G3340,G3305,G3202);
  not (G3341,G3305);
  not (G3342,G3308);
  not (G3343,G3323);
  nand (G3344,G3155,G3341);
  not (G3345,G3329);
  nand (G3346,G3329,G3342);
  not (G3347,G3320);
  and (G3350,G3312,G884);
  not (G3353,G3312);
  nand (G3356,G3340,G3344);
  nand (G3359,G3308,G3345);
  and (G3360,G884,G3332);
  and (G3363,G3199,G3323,G3317,G3337);
  and (G3366,G3317,G3337,G887);
  not (G3367,G3332);
  nand (G3370,G3359,G3346);
  not (G3373,G3347);
  not (G3376,G3347);
  not (G3379,G3353);
  not (G3380,G3350);
  not (G3383,G3350);
  and (G3386,G3326,G3363);
  and (G3387,G3326,G3363);
  not (G3388,G3356);
  not (G3391,G3356);
  not (G3394,G3367);
  nand (G3395,G3367,G3379);
  not (G3396,G3360);
  not (G3399,G3360);
  nor (G3402,G3366,G3387);
  nand (G3403,G3373,G3265);
  not (G3404,G3373);
  nand (G3405,G3376,G3266);
  not (G3406,G3376);
  not (G3407,G3380);
  not (G3408,G3383);
  not (G3409,G3370);
  not (G3412,G3370);
  nand (G3415,G3353,G3394);
  and (G3416,G27,G3402);
  not (G3417,G3388);
  not (G3418,G3391);
  nand (G3419,G3237,G3404);
  nand (G3420,G3240,G3406);
  not (G3421,G3396);
  nand (G3422,G3396,G3407);
  nand (G3423,G3399,G3408);
  not (G3424,G3399);
  nand (G3425,G3395,G3415);
  nand (G3428,G3409,G3417);
  not (G3429,G3409);
  nand (G3430,G3412,G3418);
  not (G3431,G3412);
  nand (G3432,G3403,G3419);
  nand (G3436,G3405,G3420);
  nand (G3437,G3380,G3421);
  nand (G3438,G3383,G3424);
  nand (G3439,G3388,G3429);
  nand (G3440,G3391,G3431);
  not (G3441,G3436);
  not (G3444,G3425);
  nand (G3445,G3437,G3422);
  nand (G3448,G3438,G3423);
  nand (G3449,G3428,G3439);
  nand (G3452,G3430,G3440);
  not (G3453,G3448);
  not (G3456,G3432);
  and (G3459,G3432,G3445,G1436);
  and (G3460,G3441,G3445,G1439);
  not (G3461,G3452);
  not (G3464,G3456);
  nand (G3465,G3456,G3444);
  and (G3466,G3432,G3453,G1439);
  and (G3467,G3441,G3453,G1436);
  not (G3468,G3449);
  not (G3471,G3449);
  nand (G3474,G3425,G3464);
  or (G3475,G3459,G3466,G3460,G3467);
  not (G3478,G3461);
  not (G3481,G3461);
  nand (G3484,G3474,G3465);
  not (G3487,G3471);
  not (G3488,G3468);
  not (G3489,G3481);
  not (G3490,G3478);
  not (G3491,G3475);
  not (G3494,G3475);
  not (G3497,G3484);
  not (G3500,G3484);
  nand (G3503,G3491,G3490);
  nand (G3504,G3494,G3489);
  not (G3505,G3494);
  not (G3506,G3491);
  nand (G3507,G3497,G3488);
  nand (G3508,G3500,G3487);
  nand (G3509,G3478,G3506);
  nand (G3510,G3481,G3505);
  not (G3511,G3500);
  not (G3512,G3497);
  nand (G3513,G3468,G3512);
  nand (G3514,G3471,G3511);
  nand (G3515,G3509,G3503);
  nand (G3516,G3510,G3504);
  nand (G3517,G3507,G3513);
  nand (G3518,G3508,G3514);
  not (G3519,G928);
  not (G3520,G1004);
  nand (G3521,G1786,G1811);
  nand (G3522,G2460,G2461);
  nand (G3523,G2550,G2551);
  and (G3524,G2558,G2552);
  not (G3525,G2675);
  or (G3526,G2974,G2943);
  and (G3527,G3005,G3030);
  and (G3528,G3100,G3135);
  and (G3529,G3195,G3226);
  and (G3530,G3257,G3267);
  and (G3531,G3275,G3300);
  and (G3532,G3281,G3301);
  and (G3533,G3294,G3311);
  and (G3534,G3312,G3312);
  and (G3535,G3332,G3332);
  and (G3536,G3320,G3343);
  not (G3537,G3386);
  not (G3538,G3416);
  and (G3539,G3515,G3516);
  nand (G3540,G3517,G3518);

endmodule
