
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  n940_lo,
  n949_lo,
  n961_lo,
  n973_lo,
  n976_lo,
  n985_lo,
  n988_lo,
  n997_lo,
  n1009_lo,
  n1021_lo,
  n1033_lo,
  n1045_lo,
  n1057_lo,
  n1060_lo,
  n1069_lo,
  n1081_lo,
  n1093_lo,
  n1105_lo,
  n1117_lo,
  n1120_lo,
  n1129_lo,
  n1132_lo,
  n1156_lo,
  n1168_lo,
  n1180_lo,
  n1189_lo,
  n1192_lo,
  n1195_lo,
  n1201_lo,
  n1204_lo,
  n1228_lo,
  n1231_lo,
  n1234_lo,
  n1237_lo,
  n1240_lo,
  n1243_lo,
  n1249_lo,
  n1252_lo,
  n1255_lo,
  n1261_lo,
  n1264_lo,
  n1267_lo,
  n1273_lo,
  n1276_lo,
  n1279_lo,
  n1282_lo,
  n1285_lo,
  n1288_lo,
  n1291_lo,
  n1294_lo,
  n1297_lo,
  n1300_lo,
  n1303_lo,
  n1309_lo,
  n1312_lo,
  n1315_lo,
  n1318_lo,
  n1321_lo,
  n1333_lo,
  n1225_o2,
  n1229_o2,
  n1228_o2,
  n1259_o2,
  n1272_o2,
  n1269_o2,
  n1307_o2,
  n1201_o2,
  n1202_o2,
  n1203_o2,
  n1204_o2,
  n622_o2,
  n1205_o2,
  n1206_o2,
  n497_o2,
  n1212_o2,
  n1213_o2,
  n1214_o2,
  n1215_o2,
  n1216_o2,
  n1217_o2,
  n1218_o2,
  n1219_o2,
  n1242_o2,
  n1243_o2,
  n1273_o2,
  n1274_o2,
  n1275_o2,
  n1276_o2,
  n1277_o2,
  n1286_o2,
  n1299_o2,
  n601_o2,
  n625_o2,
  n463_o2,
  lo082_buf_o2,
  n455_o2,
  n642_o2,
  n459_o2,
  n501_o2,
  n599_o2,
  n485_o2,
  lo086_buf_o2,
  lo122_buf_o2,
  n502_o2,
  n627_o2,
  lo038_buf_o2,
  lo046_buf_o2,
  lo050_buf_o2,
  lo058_buf_o2,
  lo070_buf_o2,
  lo094_buf_o2,
  n462_o2,
  lo006_buf_o2,
  lo010_buf_o2,
  lo022_buf_o2,
  lo026_buf_o2,
  lo030_buf_o2,
  lo034_buf_o2,
  lo054_buf_o2,
  lo130_buf_o2,
  n547_o2,
  n424_inv,
  n617_o2,
  lo042_buf_o2,
  lo062_buf_o2,
  lo110_buf_o2,
  n733_o2,
  n734_o2,
  n570_o2,
  n461_o2,
  n644_o2,
  n628_o2,
  n528_o2,
  n460_inv,
  lo002_buf_o2,
  lo014_buf_o2,
  lo018_buf_o2,
  lo078_buf_o2,
  lo090_buf_o2,
  n513_o2,
  lo102_buf_o2,
  lo106_buf_o2,
  n600_o2,
  n529_o2,
  n593_o2,
  lo066_buf_o2,
  n549_o2,
  n550_o2,
  n571_o2,
  n572_o2,
  n495_o2,
  n496_o2,
  n620_o2,
  n482_o2,
  lo081_buf_o2,
  n576_o2,
  n520_o2,
  n521_o2,
  n562_o2,
  n508_o2,
  n509_o2,
  lo074_buf_o2,
  n539_o2,
  n536_o2,
  n516_o2,
  n491_o2,
  n557_o2,
  n586_o2,
  n483_o2,
  n484_o2,
  lo004_buf_o2,
  lo008_buf_o2,
  lo020_buf_o2,
  lo024_buf_o2,
  lo028_buf_o2,
  lo032_buf_o2,
  lo052_buf_o2,
  lo128_buf_o2,
  lo037_buf_o2,
  lo045_buf_o2,
  lo049_buf_o2,
  lo057_buf_o2,
  lo069_buf_o2,
  lo093_buf_o2,
  G1884,
  G1885,
  G1886,
  G1887,
  G1888,
  G1889,
  G1890,
  G1891,
  G1892,
  G1893,
  G1894,
  G1895,
  G1896,
  G1897,
  G1898,
  G1899,
  G1900,
  G1901,
  G1902,
  G1903,
  G1904,
  G1905,
  G1906,
  G1907,
  G1908,
  n2248_li000_li000,
  n2257_li003_li003,
  n2269_li007_li007,
  n2281_li011_li011,
  n2284_li012_li012,
  n2293_li015_li015,
  n2296_li016_li016,
  n2305_li019_li019,
  n2317_li023_li023,
  n2329_li027_li027,
  n2341_li031_li031,
  n2353_li035_li035,
  n2365_li039_li039,
  n2368_li040_li040,
  n2377_li043_li043,
  n2389_li047_li047,
  n2401_li051_li051,
  n2413_li055_li055,
  n2425_li059_li059,
  n2428_li060_li060,
  n2437_li063_li063,
  n2440_li064_li064,
  n2464_li072_li072,
  n2476_li076_li076,
  n2488_li080_li080,
  n2497_li083_li083,
  n2500_li084_li084,
  n2503_li085_li085,
  n2509_li087_li087,
  n2512_li088_li088,
  n2536_li096_li096,
  n2539_li097_li097,
  n2542_li098_li098,
  n2545_li099_li099,
  n2548_li100_li100,
  n2551_li101_li101,
  n2557_li103_li103,
  n2560_li104_li104,
  n2563_li105_li105,
  n2569_li107_li107,
  n2572_li108_li108,
  n2575_li109_li109,
  n2581_li111_li111,
  n2584_li112_li112,
  n2587_li113_li113,
  n2590_li114_li114,
  n2593_li115_li115,
  n2596_li116_li116,
  n2599_li117_li117,
  n2602_li118_li118,
  n2605_li119_li119,
  n2608_li120_li120,
  n2611_li121_li121,
  n2617_li123_li123,
  n2620_li124_li124,
  n2623_li125_li125,
  n2626_li126_li126,
  n2629_li127_li127,
  n2641_li131_li131,
  n1225_i2,
  n1229_i2,
  n1228_i2,
  n1259_i2,
  n1272_i2,
  n1269_i2,
  n1307_i2,
  n1201_i2,
  n1202_i2,
  n1203_i2,
  n1204_i2,
  n622_i2,
  n1205_i2,
  n1206_i2,
  n497_i2,
  n1212_i2,
  n1213_i2,
  n1214_i2,
  n1215_i2,
  n1216_i2,
  n1217_i2,
  n1218_i2,
  n1219_i2,
  n1242_i2,
  n1243_i2,
  n1273_i2,
  n1274_i2,
  n1275_i2,
  n1276_i2,
  n1277_i2,
  n1286_i2,
  n1299_i2,
  n601_i2,
  n625_i2,
  n463_i2,
  lo082_buf_i2,
  n455_i2,
  n642_i2,
  n459_i2,
  n501_i2,
  n599_i2,
  n485_i2,
  lo086_buf_i2,
  lo122_buf_i2,
  n502_i2,
  n627_i2,
  lo038_buf_i2,
  lo046_buf_i2,
  lo050_buf_i2,
  lo058_buf_i2,
  lo070_buf_i2,
  lo094_buf_i2,
  n462_i2,
  lo006_buf_i2,
  lo010_buf_i2,
  lo022_buf_i2,
  lo026_buf_i2,
  lo030_buf_i2,
  lo034_buf_i2,
  lo054_buf_i2,
  lo130_buf_i2,
  n547_i2,
  n568_i2,
  n617_i2,
  lo042_buf_i2,
  lo062_buf_i2,
  lo110_buf_i2,
  n733_i2,
  n734_i2,
  n570_i2,
  n461_i2,
  n644_i2,
  n628_i2,
  n528_i2,
  n592_i2,
  lo002_buf_i2,
  lo014_buf_i2,
  lo018_buf_i2,
  lo078_buf_i2,
  lo090_buf_i2,
  n513_i2,
  lo102_buf_i2,
  lo106_buf_i2,
  n600_i2,
  n529_i2,
  n593_i2,
  lo066_buf_i2,
  n549_i2,
  n550_i2,
  n571_i2,
  n572_i2,
  n495_i2,
  n496_i2,
  n620_i2,
  n482_i2,
  lo081_buf_i2,
  n576_i2,
  n520_i2,
  n521_i2,
  n562_i2,
  n508_i2,
  n509_i2,
  lo074_buf_i2,
  n539_i2,
  n536_i2,
  n516_i2,
  n491_i2,
  n557_i2,
  n586_i2,
  n483_i2,
  n484_i2,
  lo004_buf_i2,
  lo008_buf_i2,
  lo020_buf_i2,
  lo024_buf_i2,
  lo028_buf_i2,
  lo032_buf_i2,
  lo052_buf_i2,
  lo128_buf_i2,
  lo037_buf_i2,
  lo045_buf_i2,
  lo049_buf_i2,
  lo057_buf_i2,
  lo069_buf_i2,
  lo093_buf_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input n940_lo;input n949_lo;input n961_lo;input n973_lo;input n976_lo;input n985_lo;input n988_lo;input n997_lo;input n1009_lo;input n1021_lo;input n1033_lo;input n1045_lo;input n1057_lo;input n1060_lo;input n1069_lo;input n1081_lo;input n1093_lo;input n1105_lo;input n1117_lo;input n1120_lo;input n1129_lo;input n1132_lo;input n1156_lo;input n1168_lo;input n1180_lo;input n1189_lo;input n1192_lo;input n1195_lo;input n1201_lo;input n1204_lo;input n1228_lo;input n1231_lo;input n1234_lo;input n1237_lo;input n1240_lo;input n1243_lo;input n1249_lo;input n1252_lo;input n1255_lo;input n1261_lo;input n1264_lo;input n1267_lo;input n1273_lo;input n1276_lo;input n1279_lo;input n1282_lo;input n1285_lo;input n1288_lo;input n1291_lo;input n1294_lo;input n1297_lo;input n1300_lo;input n1303_lo;input n1309_lo;input n1312_lo;input n1315_lo;input n1318_lo;input n1321_lo;input n1333_lo;input n1225_o2;input n1229_o2;input n1228_o2;input n1259_o2;input n1272_o2;input n1269_o2;input n1307_o2;input n1201_o2;input n1202_o2;input n1203_o2;input n1204_o2;input n622_o2;input n1205_o2;input n1206_o2;input n497_o2;input n1212_o2;input n1213_o2;input n1214_o2;input n1215_o2;input n1216_o2;input n1217_o2;input n1218_o2;input n1219_o2;input n1242_o2;input n1243_o2;input n1273_o2;input n1274_o2;input n1275_o2;input n1276_o2;input n1277_o2;input n1286_o2;input n1299_o2;input n601_o2;input n625_o2;input n463_o2;input lo082_buf_o2;input n455_o2;input n642_o2;input n459_o2;input n501_o2;input n599_o2;input n485_o2;input lo086_buf_o2;input lo122_buf_o2;input n502_o2;input n627_o2;input lo038_buf_o2;input lo046_buf_o2;input lo050_buf_o2;input lo058_buf_o2;input lo070_buf_o2;input lo094_buf_o2;input n462_o2;input lo006_buf_o2;input lo010_buf_o2;input lo022_buf_o2;input lo026_buf_o2;input lo030_buf_o2;input lo034_buf_o2;input lo054_buf_o2;input lo130_buf_o2;input n547_o2;input n424_inv;input n617_o2;input lo042_buf_o2;input lo062_buf_o2;input lo110_buf_o2;input n733_o2;input n734_o2;input n570_o2;input n461_o2;input n644_o2;input n628_o2;input n528_o2;input n460_inv;input lo002_buf_o2;input lo014_buf_o2;input lo018_buf_o2;input lo078_buf_o2;input lo090_buf_o2;input n513_o2;input lo102_buf_o2;input lo106_buf_o2;input n600_o2;input n529_o2;input n593_o2;input lo066_buf_o2;input n549_o2;input n550_o2;input n571_o2;input n572_o2;input n495_o2;input n496_o2;input n620_o2;input n482_o2;input lo081_buf_o2;input n576_o2;input n520_o2;input n521_o2;input n562_o2;input n508_o2;input n509_o2;input lo074_buf_o2;input n539_o2;input n536_o2;input n516_o2;input n491_o2;input n557_o2;input n586_o2;input n483_o2;input n484_o2;input lo004_buf_o2;input lo008_buf_o2;input lo020_buf_o2;input lo024_buf_o2;input lo028_buf_o2;input lo032_buf_o2;input lo052_buf_o2;input lo128_buf_o2;input lo037_buf_o2;input lo045_buf_o2;input lo049_buf_o2;input lo057_buf_o2;input lo069_buf_o2;input lo093_buf_o2;
  output G1884;output G1885;output G1886;output G1887;output G1888;output G1889;output G1890;output G1891;output G1892;output G1893;output G1894;output G1895;output G1896;output G1897;output G1898;output G1899;output G1900;output G1901;output G1902;output G1903;output G1904;output G1905;output G1906;output G1907;output G1908;output n2248_li000_li000;output n2257_li003_li003;output n2269_li007_li007;output n2281_li011_li011;output n2284_li012_li012;output n2293_li015_li015;output n2296_li016_li016;output n2305_li019_li019;output n2317_li023_li023;output n2329_li027_li027;output n2341_li031_li031;output n2353_li035_li035;output n2365_li039_li039;output n2368_li040_li040;output n2377_li043_li043;output n2389_li047_li047;output n2401_li051_li051;output n2413_li055_li055;output n2425_li059_li059;output n2428_li060_li060;output n2437_li063_li063;output n2440_li064_li064;output n2464_li072_li072;output n2476_li076_li076;output n2488_li080_li080;output n2497_li083_li083;output n2500_li084_li084;output n2503_li085_li085;output n2509_li087_li087;output n2512_li088_li088;output n2536_li096_li096;output n2539_li097_li097;output n2542_li098_li098;output n2545_li099_li099;output n2548_li100_li100;output n2551_li101_li101;output n2557_li103_li103;output n2560_li104_li104;output n2563_li105_li105;output n2569_li107_li107;output n2572_li108_li108;output n2575_li109_li109;output n2581_li111_li111;output n2584_li112_li112;output n2587_li113_li113;output n2590_li114_li114;output n2593_li115_li115;output n2596_li116_li116;output n2599_li117_li117;output n2602_li118_li118;output n2605_li119_li119;output n2608_li120_li120;output n2611_li121_li121;output n2617_li123_li123;output n2620_li124_li124;output n2623_li125_li125;output n2626_li126_li126;output n2629_li127_li127;output n2641_li131_li131;output n1225_i2;output n1229_i2;output n1228_i2;output n1259_i2;output n1272_i2;output n1269_i2;output n1307_i2;output n1201_i2;output n1202_i2;output n1203_i2;output n1204_i2;output n622_i2;output n1205_i2;output n1206_i2;output n497_i2;output n1212_i2;output n1213_i2;output n1214_i2;output n1215_i2;output n1216_i2;output n1217_i2;output n1218_i2;output n1219_i2;output n1242_i2;output n1243_i2;output n1273_i2;output n1274_i2;output n1275_i2;output n1276_i2;output n1277_i2;output n1286_i2;output n1299_i2;output n601_i2;output n625_i2;output n463_i2;output lo082_buf_i2;output n455_i2;output n642_i2;output n459_i2;output n501_i2;output n599_i2;output n485_i2;output lo086_buf_i2;output lo122_buf_i2;output n502_i2;output n627_i2;output lo038_buf_i2;output lo046_buf_i2;output lo050_buf_i2;output lo058_buf_i2;output lo070_buf_i2;output lo094_buf_i2;output n462_i2;output lo006_buf_i2;output lo010_buf_i2;output lo022_buf_i2;output lo026_buf_i2;output lo030_buf_i2;output lo034_buf_i2;output lo054_buf_i2;output lo130_buf_i2;output n547_i2;output n568_i2;output n617_i2;output lo042_buf_i2;output lo062_buf_i2;output lo110_buf_i2;output n733_i2;output n734_i2;output n570_i2;output n461_i2;output n644_i2;output n628_i2;output n528_i2;output n592_i2;output lo002_buf_i2;output lo014_buf_i2;output lo018_buf_i2;output lo078_buf_i2;output lo090_buf_i2;output n513_i2;output lo102_buf_i2;output lo106_buf_i2;output n600_i2;output n529_i2;output n593_i2;output lo066_buf_i2;output n549_i2;output n550_i2;output n571_i2;output n572_i2;output n495_i2;output n496_i2;output n620_i2;output n482_i2;output lo081_buf_i2;output n576_i2;output n520_i2;output n521_i2;output n562_i2;output n508_i2;output n509_i2;output lo074_buf_i2;output n539_i2;output n536_i2;output n516_i2;output n491_i2;output n557_i2;output n586_i2;output n483_i2;output n484_i2;output lo004_buf_i2;output lo008_buf_i2;output lo020_buf_i2;output lo024_buf_i2;output lo028_buf_i2;output lo032_buf_i2;output lo052_buf_i2;output lo128_buf_i2;output lo037_buf_i2;output lo045_buf_i2;output lo049_buf_i2;output lo057_buf_i2;output lo069_buf_i2;output lo093_buf_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire n940_lo_p;
  wire n940_lo_n;
  wire n949_lo_p;
  wire n949_lo_n;
  wire n961_lo_p;
  wire n961_lo_n;
  wire n973_lo_p;
  wire n973_lo_n;
  wire n976_lo_p;
  wire n976_lo_n;
  wire n985_lo_p;
  wire n985_lo_n;
  wire n988_lo_p;
  wire n988_lo_n;
  wire n997_lo_p;
  wire n997_lo_n;
  wire n1009_lo_p;
  wire n1009_lo_n;
  wire n1021_lo_p;
  wire n1021_lo_n;
  wire n1033_lo_p;
  wire n1033_lo_n;
  wire n1045_lo_p;
  wire n1045_lo_n;
  wire n1057_lo_p;
  wire n1057_lo_n;
  wire n1060_lo_p;
  wire n1060_lo_n;
  wire n1069_lo_p;
  wire n1069_lo_n;
  wire n1081_lo_p;
  wire n1081_lo_n;
  wire n1093_lo_p;
  wire n1093_lo_n;
  wire n1105_lo_p;
  wire n1105_lo_n;
  wire n1117_lo_p;
  wire n1117_lo_n;
  wire n1120_lo_p;
  wire n1120_lo_n;
  wire n1129_lo_p;
  wire n1129_lo_n;
  wire n1132_lo_p;
  wire n1132_lo_n;
  wire n1156_lo_p;
  wire n1156_lo_n;
  wire n1168_lo_p;
  wire n1168_lo_n;
  wire n1180_lo_p;
  wire n1180_lo_n;
  wire n1189_lo_p;
  wire n1189_lo_n;
  wire n1192_lo_p;
  wire n1192_lo_n;
  wire n1195_lo_p;
  wire n1195_lo_n;
  wire n1201_lo_p;
  wire n1201_lo_n;
  wire n1204_lo_p;
  wire n1204_lo_n;
  wire n1228_lo_p;
  wire n1228_lo_n;
  wire n1231_lo_p;
  wire n1231_lo_n;
  wire n1234_lo_p;
  wire n1234_lo_n;
  wire n1237_lo_p;
  wire n1237_lo_n;
  wire n1240_lo_p;
  wire n1240_lo_n;
  wire n1243_lo_p;
  wire n1243_lo_n;
  wire n1249_lo_p;
  wire n1249_lo_n;
  wire n1252_lo_p;
  wire n1252_lo_n;
  wire n1255_lo_p;
  wire n1255_lo_n;
  wire n1261_lo_p;
  wire n1261_lo_n;
  wire n1264_lo_p;
  wire n1264_lo_n;
  wire n1267_lo_p;
  wire n1267_lo_n;
  wire n1273_lo_p;
  wire n1273_lo_n;
  wire n1276_lo_p;
  wire n1276_lo_n;
  wire n1279_lo_p;
  wire n1279_lo_n;
  wire n1282_lo_p;
  wire n1282_lo_n;
  wire n1285_lo_p;
  wire n1285_lo_n;
  wire n1288_lo_p;
  wire n1288_lo_n;
  wire n1291_lo_p;
  wire n1291_lo_n;
  wire n1294_lo_p;
  wire n1294_lo_n;
  wire n1297_lo_p;
  wire n1297_lo_n;
  wire n1300_lo_p;
  wire n1300_lo_n;
  wire n1303_lo_p;
  wire n1303_lo_n;
  wire n1309_lo_p;
  wire n1309_lo_n;
  wire n1312_lo_p;
  wire n1312_lo_n;
  wire n1315_lo_p;
  wire n1315_lo_n;
  wire n1318_lo_p;
  wire n1318_lo_n;
  wire n1321_lo_p;
  wire n1321_lo_n;
  wire n1333_lo_p;
  wire n1333_lo_n;
  wire n1225_o2_p;
  wire n1225_o2_n;
  wire n1229_o2_p;
  wire n1229_o2_n;
  wire n1228_o2_p;
  wire n1228_o2_n;
  wire n1259_o2_p;
  wire n1259_o2_n;
  wire n1272_o2_p;
  wire n1272_o2_n;
  wire n1269_o2_p;
  wire n1269_o2_n;
  wire n1307_o2_p;
  wire n1307_o2_n;
  wire n1201_o2_p;
  wire n1201_o2_n;
  wire n1202_o2_p;
  wire n1202_o2_n;
  wire n1203_o2_p;
  wire n1203_o2_n;
  wire n1204_o2_p;
  wire n1204_o2_n;
  wire n622_o2_p;
  wire n622_o2_n;
  wire n1205_o2_p;
  wire n1205_o2_n;
  wire n1206_o2_p;
  wire n1206_o2_n;
  wire n497_o2_p;
  wire n497_o2_n;
  wire n1212_o2_p;
  wire n1212_o2_n;
  wire n1213_o2_p;
  wire n1213_o2_n;
  wire n1214_o2_p;
  wire n1214_o2_n;
  wire n1215_o2_p;
  wire n1215_o2_n;
  wire n1216_o2_p;
  wire n1216_o2_n;
  wire n1217_o2_p;
  wire n1217_o2_n;
  wire n1218_o2_p;
  wire n1218_o2_n;
  wire n1219_o2_p;
  wire n1219_o2_n;
  wire n1242_o2_p;
  wire n1242_o2_n;
  wire n1243_o2_p;
  wire n1243_o2_n;
  wire n1273_o2_p;
  wire n1273_o2_n;
  wire n1274_o2_p;
  wire n1274_o2_n;
  wire n1275_o2_p;
  wire n1275_o2_n;
  wire n1276_o2_p;
  wire n1276_o2_n;
  wire n1277_o2_p;
  wire n1277_o2_n;
  wire n1286_o2_p;
  wire n1286_o2_n;
  wire n1299_o2_p;
  wire n1299_o2_n;
  wire n601_o2_p;
  wire n601_o2_n;
  wire n625_o2_p;
  wire n625_o2_n;
  wire n463_o2_p;
  wire n463_o2_n;
  wire lo082_buf_o2_p;
  wire lo082_buf_o2_n;
  wire n455_o2_p;
  wire n455_o2_n;
  wire n642_o2_p;
  wire n642_o2_n;
  wire n459_o2_p;
  wire n459_o2_n;
  wire n501_o2_p;
  wire n501_o2_n;
  wire n599_o2_p;
  wire n599_o2_n;
  wire n485_o2_p;
  wire n485_o2_n;
  wire lo086_buf_o2_p;
  wire lo086_buf_o2_n;
  wire lo122_buf_o2_p;
  wire lo122_buf_o2_n;
  wire n502_o2_p;
  wire n502_o2_n;
  wire n627_o2_p;
  wire n627_o2_n;
  wire lo038_buf_o2_p;
  wire lo038_buf_o2_n;
  wire lo046_buf_o2_p;
  wire lo046_buf_o2_n;
  wire lo050_buf_o2_p;
  wire lo050_buf_o2_n;
  wire lo058_buf_o2_p;
  wire lo058_buf_o2_n;
  wire lo070_buf_o2_p;
  wire lo070_buf_o2_n;
  wire lo094_buf_o2_p;
  wire lo094_buf_o2_n;
  wire n462_o2_p;
  wire n462_o2_n;
  wire lo006_buf_o2_p;
  wire lo006_buf_o2_n;
  wire lo010_buf_o2_p;
  wire lo010_buf_o2_n;
  wire lo022_buf_o2_p;
  wire lo022_buf_o2_n;
  wire lo026_buf_o2_p;
  wire lo026_buf_o2_n;
  wire lo030_buf_o2_p;
  wire lo030_buf_o2_n;
  wire lo034_buf_o2_p;
  wire lo034_buf_o2_n;
  wire lo054_buf_o2_p;
  wire lo054_buf_o2_n;
  wire lo130_buf_o2_p;
  wire lo130_buf_o2_n;
  wire n547_o2_p;
  wire n547_o2_n;
  wire n424_inv_p;
  wire n424_inv_n;
  wire n617_o2_p;
  wire n617_o2_n;
  wire lo042_buf_o2_p;
  wire lo042_buf_o2_n;
  wire lo062_buf_o2_p;
  wire lo062_buf_o2_n;
  wire lo110_buf_o2_p;
  wire lo110_buf_o2_n;
  wire n733_o2_p;
  wire n733_o2_n;
  wire n734_o2_p;
  wire n734_o2_n;
  wire n570_o2_p;
  wire n570_o2_n;
  wire n461_o2_p;
  wire n461_o2_n;
  wire n644_o2_p;
  wire n644_o2_n;
  wire n628_o2_p;
  wire n628_o2_n;
  wire n528_o2_p;
  wire n528_o2_n;
  wire n460_inv_p;
  wire n460_inv_n;
  wire lo002_buf_o2_p;
  wire lo002_buf_o2_n;
  wire lo014_buf_o2_p;
  wire lo014_buf_o2_n;
  wire lo018_buf_o2_p;
  wire lo018_buf_o2_n;
  wire lo078_buf_o2_p;
  wire lo078_buf_o2_n;
  wire lo090_buf_o2_p;
  wire lo090_buf_o2_n;
  wire n513_o2_p;
  wire n513_o2_n;
  wire lo102_buf_o2_p;
  wire lo102_buf_o2_n;
  wire lo106_buf_o2_p;
  wire lo106_buf_o2_n;
  wire n600_o2_p;
  wire n600_o2_n;
  wire n529_o2_p;
  wire n529_o2_n;
  wire n593_o2_p;
  wire n593_o2_n;
  wire lo066_buf_o2_p;
  wire lo066_buf_o2_n;
  wire n549_o2_p;
  wire n549_o2_n;
  wire n550_o2_p;
  wire n550_o2_n;
  wire n571_o2_p;
  wire n571_o2_n;
  wire n572_o2_p;
  wire n572_o2_n;
  wire n495_o2_p;
  wire n495_o2_n;
  wire n496_o2_p;
  wire n496_o2_n;
  wire n620_o2_p;
  wire n620_o2_n;
  wire n482_o2_p;
  wire n482_o2_n;
  wire lo081_buf_o2_p;
  wire lo081_buf_o2_n;
  wire n576_o2_p;
  wire n576_o2_n;
  wire n520_o2_p;
  wire n520_o2_n;
  wire n521_o2_p;
  wire n521_o2_n;
  wire n562_o2_p;
  wire n562_o2_n;
  wire n508_o2_p;
  wire n508_o2_n;
  wire n509_o2_p;
  wire n509_o2_n;
  wire lo074_buf_o2_p;
  wire lo074_buf_o2_n;
  wire n539_o2_p;
  wire n539_o2_n;
  wire n536_o2_p;
  wire n536_o2_n;
  wire n516_o2_p;
  wire n516_o2_n;
  wire n491_o2_p;
  wire n491_o2_n;
  wire n557_o2_p;
  wire n557_o2_n;
  wire n586_o2_p;
  wire n586_o2_n;
  wire n483_o2_p;
  wire n483_o2_n;
  wire n484_o2_p;
  wire n484_o2_n;
  wire lo004_buf_o2_p;
  wire lo004_buf_o2_n;
  wire lo008_buf_o2_p;
  wire lo008_buf_o2_n;
  wire lo020_buf_o2_p;
  wire lo020_buf_o2_n;
  wire lo024_buf_o2_p;
  wire lo024_buf_o2_n;
  wire lo028_buf_o2_p;
  wire lo028_buf_o2_n;
  wire lo032_buf_o2_p;
  wire lo032_buf_o2_n;
  wire lo052_buf_o2_p;
  wire lo052_buf_o2_n;
  wire lo128_buf_o2_p;
  wire lo128_buf_o2_n;
  wire lo037_buf_o2_p;
  wire lo037_buf_o2_n;
  wire lo045_buf_o2_p;
  wire lo045_buf_o2_n;
  wire lo049_buf_o2_p;
  wire lo049_buf_o2_n;
  wire lo057_buf_o2_p;
  wire lo057_buf_o2_n;
  wire lo069_buf_o2_p;
  wire lo069_buf_o2_n;
  wire lo093_buf_o2_p;
  wire lo093_buf_o2_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire n461_o2_n_spl_;
  wire n628_o2_p_spl_;
  wire n461_o2_p_spl_;
  wire n628_o2_n_spl_;
  wire g218_n_spl_;
  wire g218_n_spl_0;
  wire g218_n_spl_00;
  wire g218_n_spl_01;
  wire g218_n_spl_1;
  wire g218_n_spl_10;
  wire g218_p_spl_;
  wire g218_p_spl_0;
  wire g218_p_spl_00;
  wire g218_p_spl_01;
  wire g218_p_spl_1;
  wire g218_p_spl_10;
  wire n644_o2_n_spl_;
  wire n644_o2_n_spl_0;
  wire n644_o2_p_spl_;
  wire n644_o2_p_spl_0;
  wire g231_n_spl_;
  wire g231_n_spl_0;
  wire g231_n_spl_00;
  wire g231_n_spl_01;
  wire g231_n_spl_1;
  wire g231_p_spl_;
  wire g231_p_spl_0;
  wire g231_p_spl_00;
  wire g231_p_spl_01;
  wire g231_p_spl_1;
  wire n501_o2_n_spl_;
  wire n463_o2_n_spl_;
  wire g242_p_spl_;
  wire g242_n_spl_;
  wire g243_n_spl_;
  wire g243_n_spl_0;
  wire g243_n_spl_1;
  wire g243_p_spl_;
  wire g243_p_spl_0;
  wire g243_p_spl_1;
  wire n601_o2_n_spl_;
  wire n625_o2_p_spl_;
  wire n599_o2_p_spl_;
  wire g263_n_spl_;
  wire g263_n_spl_0;
  wire g263_n_spl_1;
  wire g263_p_spl_;
  wire g263_p_spl_0;
  wire g263_p_spl_1;
  wire g276_n_spl_;
  wire g276_n_spl_0;
  wire g276_n_spl_00;
  wire g276_n_spl_01;
  wire g276_n_spl_1;
  wire n1333_lo_p_spl_;
  wire n1333_lo_p_spl_0;
  wire n1309_lo_n_spl_;
  wire n1309_lo_n_spl_0;
  wire n1309_lo_n_spl_00;
  wire n1309_lo_n_spl_1;
  wire n1309_lo_p_spl_;
  wire n1309_lo_p_spl_0;
  wire g276_p_spl_;
  wire g276_p_spl_0;
  wire n459_o2_p_spl_;
  wire n459_o2_p_spl_0;
  wire n459_o2_p_spl_00;
  wire n459_o2_p_spl_01;
  wire n459_o2_p_spl_1;
  wire n1333_lo_n_spl_;
  wire g310_n_spl_;
  wire g310_p_spl_;
  wire g320_n_spl_;
  wire g320_p_spl_;
  wire n600_o2_n_spl_;
  wire lo122_buf_o2_n_spl_;
  wire lo122_buf_o2_p_spl_;
  wire lo122_buf_o2_p_spl_0;
  wire lo122_buf_o2_p_spl_1;
  wire n620_o2_p_spl_;
  wire g331_p_spl_;
  wire n1282_lo_p_spl_;
  wire n1219_o2_p_spl_;
  wire n1219_o2_p_spl_0;
  wire n1219_o2_p_spl_1;
  wire n1294_lo_p_spl_;
  wire n1318_lo_p_spl_;
  wire g332_n_spl_;
  wire n1234_lo_p_spl_;
  wire lo106_buf_o2_p_spl_;
  wire lo102_buf_o2_p_spl_;
  wire g338_n_spl_;
  wire g345_p_spl_;
  wire g333_n_spl_;
  wire g337_p_spl_;
  wire g356_p_spl_;
  wire n1303_lo_p_spl_;
  wire n1303_lo_p_spl_0;
  wire n1303_lo_p_spl_1;
  wire lo090_buf_o2_p_spl_;
  wire lo090_buf_o2_p_spl_0;
  wire n539_o2_n_spl_;
  wire n536_o2_p_spl_;
  wire n539_o2_p_spl_;
  wire n536_o2_n_spl_;
  wire lo074_buf_o2_p_spl_;
  wire lo130_buf_o2_n_spl_;
  wire lo130_buf_o2_n_spl_0;
  wire lo130_buf_o2_n_spl_1;
  wire lo130_buf_o2_p_spl_;
  wire lo130_buf_o2_p_spl_0;
  wire lo130_buf_o2_p_spl_00;
  wire lo130_buf_o2_p_spl_1;
  wire n516_o2_n_spl_;
  wire n516_o2_n_spl_0;
  wire n516_o2_n_spl_1;
  wire n557_o2_p_spl_;
  wire n516_o2_p_spl_;
  wire n516_o2_p_spl_0;
  wire n516_o2_p_spl_1;
  wire n557_o2_n_spl_;
  wire lo050_buf_o2_n_spl_;
  wire n562_o2_p_spl_;
  wire lo050_buf_o2_p_spl_;
  wire lo050_buf_o2_p_spl_0;
  wire n562_o2_n_spl_;
  wire n491_o2_p_spl_;
  wire n491_o2_p_spl_0;
  wire n586_o2_p_spl_;
  wire n586_o2_p_spl_0;
  wire n586_o2_p_spl_1;
  wire n491_o2_n_spl_;
  wire n491_o2_n_spl_0;
  wire n586_o2_n_spl_;
  wire n586_o2_n_spl_0;
  wire n586_o2_n_spl_1;
  wire lo030_buf_o2_n_spl_;
  wire lo014_buf_o2_p_spl_;
  wire lo014_buf_o2_p_spl_0;
  wire lo014_buf_o2_p_spl_00;
  wire lo014_buf_o2_p_spl_1;
  wire lo030_buf_o2_p_spl_;
  wire lo030_buf_o2_p_spl_0;
  wire lo014_buf_o2_n_spl_;
  wire lo014_buf_o2_n_spl_0;
  wire lo014_buf_o2_n_spl_1;
  wire g381_n_spl_;
  wire g384_p_spl_;
  wire g381_p_spl_;
  wire g384_n_spl_;
  wire g361_n_spl_;
  wire g391_p_spl_;
  wire g339_n_spl_;
  wire g392_n_spl_;
  wire g341_n_spl_;
  wire g394_n_spl_;
  wire g340_n_spl_;
  wire g358_n_spl_;
  wire g360_p_spl_;
  wire g399_p_spl_;
  wire g399_n_spl_;
  wire lo006_buf_o2_n_spl_;
  wire g403_n_spl_;
  wire lo006_buf_o2_p_spl_;
  wire lo006_buf_o2_p_spl_0;
  wire g403_p_spl_;
  wire lo002_buf_o2_p_spl_;
  wire lo002_buf_o2_p_spl_0;
  wire g410_p_spl_;
  wire lo002_buf_o2_n_spl_;
  wire g410_n_spl_;
  wire g357_p_spl_;
  wire g357_p_spl_0;
  wire g357_n_spl_;
  wire g357_n_spl_0;
  wire g357_n_spl_1;
  wire lo032_buf_o2_n_spl_;
  wire lo052_buf_o2_n_spl_;
  wire lo032_buf_o2_p_spl_;
  wire lo032_buf_o2_p_spl_0;
  wire lo052_buf_o2_p_spl_;
  wire lo052_buf_o2_p_spl_0;
  wire lo094_buf_o2_p_spl_;
  wire n1303_lo_n_spl_;
  wire n1303_lo_n_spl_0;
  wire g409_n_spl_;
  wire g419_n_spl_;
  wire g369_n_spl_;
  wire n1267_lo_n_spl_;
  wire g426_p_spl_;
  wire g378_p_spl_;
  wire g390_p_spl_;
  wire g390_p_spl_0;
  wire g429_n_spl_;
  wire n1195_lo_p_spl_;
  wire lo054_buf_o2_n_spl_;
  wire lo054_buf_o2_p_spl_;
  wire lo054_buf_o2_p_spl_0;
  wire g438_n_spl_;
  wire g441_p_spl_;
  wire lo081_buf_o2_p_spl_;
  wire lo034_buf_o2_p_spl_;
  wire lo034_buf_o2_p_spl_0;
  wire n482_o2_n_spl_;
  wire lo034_buf_o2_n_spl_;
  wire n482_o2_p_spl_;
  wire g444_p_spl_;
  wire g447_n_spl_;
  wire g444_n_spl_;
  wire g447_p_spl_;
  wire g387_p_spl_;
  wire lo037_buf_o2_p_spl_;
  wire lo037_buf_o2_p_spl_0;
  wire lo037_buf_o2_p_spl_00;
  wire lo037_buf_o2_p_spl_1;
  wire lo057_buf_o2_n_spl_;
  wire lo057_buf_o2_n_spl_0;
  wire lo037_buf_o2_n_spl_;
  wire lo037_buf_o2_n_spl_0;
  wire lo037_buf_o2_n_spl_1;
  wire lo057_buf_o2_p_spl_;
  wire lo057_buf_o2_p_spl_0;
  wire lo057_buf_o2_p_spl_1;
  wire n1120_lo_p_spl_;
  wire n1120_lo_p_spl_0;
  wire g456_n_spl_;
  wire n1120_lo_n_spl_;
  wire g456_p_spl_;
  wire n1132_lo_p_spl_;
  wire lo093_buf_o2_n_spl_;
  wire n988_lo_p_spl_;
  wire n988_lo_p_spl_0;
  wire lo028_buf_o2_n_spl_;
  wire lo028_buf_o2_n_spl_0;
  wire n988_lo_n_spl_;
  wire lo028_buf_o2_p_spl_;
  wire lo028_buf_o2_p_spl_0;
  wire lo028_buf_o2_p_spl_1;
  wire n1168_lo_p_spl_;
  wire lo128_buf_o2_n_spl_;
  wire lo069_buf_o2_p_spl_;
  wire lo093_buf_o2_p_spl_;
  wire lo128_buf_o2_p_spl_;
  wire n1060_lo_n_spl_;
  wire n1060_lo_n_spl_0;
  wire g469_n_spl_;
  wire lo045_buf_o2_n_spl_;
  wire lo045_buf_o2_n_spl_0;
  wire lo045_buf_o2_p_spl_;
  wire lo045_buf_o2_p_spl_0;
  wire lo045_buf_o2_p_spl_1;
  wire lo020_buf_o2_p_spl_;
  wire lo020_buf_o2_p_spl_0;
  wire lo020_buf_o2_p_spl_00;
  wire lo020_buf_o2_p_spl_1;
  wire lo020_buf_o2_n_spl_;
  wire lo020_buf_o2_n_spl_0;
  wire lo020_buf_o2_n_spl_1;
  wire lo008_buf_o2_n_spl_;
  wire lo008_buf_o2_n_spl_0;
  wire lo008_buf_o2_p_spl_;
  wire lo008_buf_o2_p_spl_0;
  wire lo008_buf_o2_p_spl_1;
  wire g422_p_spl_;
  wire lo004_buf_o2_n_spl_;
  wire lo004_buf_o2_p_spl_;
  wire lo004_buf_o2_p_spl_0;
  wire n940_lo_p_spl_;
  wire lo024_buf_o2_p_spl_;
  wire lo024_buf_o2_p_spl_0;
  wire lo024_buf_o2_p_spl_00;
  wire lo024_buf_o2_p_spl_1;
  wire lo024_buf_o2_n_spl_;
  wire lo024_buf_o2_n_spl_0;
  wire lo024_buf_o2_n_spl_1;
  wire n976_lo_p_spl_;
  wire lo049_buf_o2_n_spl_;
  wire lo049_buf_o2_p_spl_;
  wire lo049_buf_o2_p_spl_0;
  wire n1060_lo_p_spl_;
  wire g459_n_spl_;
  wire g459_n_spl_0;
  wire g507_n_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    n940_lo_p,
    n940_lo
  );


  not

  (
    n940_lo_n,
    n940_lo
  );


  buf

  (
    n949_lo_p,
    n949_lo
  );


  not

  (
    n949_lo_n,
    n949_lo
  );


  buf

  (
    n961_lo_p,
    n961_lo
  );


  not

  (
    n961_lo_n,
    n961_lo
  );


  buf

  (
    n973_lo_p,
    n973_lo
  );


  not

  (
    n973_lo_n,
    n973_lo
  );


  buf

  (
    n976_lo_p,
    n976_lo
  );


  not

  (
    n976_lo_n,
    n976_lo
  );


  buf

  (
    n985_lo_p,
    n985_lo
  );


  not

  (
    n985_lo_n,
    n985_lo
  );


  buf

  (
    n988_lo_p,
    n988_lo
  );


  not

  (
    n988_lo_n,
    n988_lo
  );


  buf

  (
    n997_lo_p,
    n997_lo
  );


  not

  (
    n997_lo_n,
    n997_lo
  );


  buf

  (
    n1009_lo_p,
    n1009_lo
  );


  not

  (
    n1009_lo_n,
    n1009_lo
  );


  buf

  (
    n1021_lo_p,
    n1021_lo
  );


  not

  (
    n1021_lo_n,
    n1021_lo
  );


  buf

  (
    n1033_lo_p,
    n1033_lo
  );


  not

  (
    n1033_lo_n,
    n1033_lo
  );


  buf

  (
    n1045_lo_p,
    n1045_lo
  );


  not

  (
    n1045_lo_n,
    n1045_lo
  );


  buf

  (
    n1057_lo_p,
    n1057_lo
  );


  not

  (
    n1057_lo_n,
    n1057_lo
  );


  buf

  (
    n1060_lo_p,
    n1060_lo
  );


  not

  (
    n1060_lo_n,
    n1060_lo
  );


  buf

  (
    n1069_lo_p,
    n1069_lo
  );


  not

  (
    n1069_lo_n,
    n1069_lo
  );


  buf

  (
    n1081_lo_p,
    n1081_lo
  );


  not

  (
    n1081_lo_n,
    n1081_lo
  );


  buf

  (
    n1093_lo_p,
    n1093_lo
  );


  not

  (
    n1093_lo_n,
    n1093_lo
  );


  buf

  (
    n1105_lo_p,
    n1105_lo
  );


  not

  (
    n1105_lo_n,
    n1105_lo
  );


  buf

  (
    n1117_lo_p,
    n1117_lo
  );


  not

  (
    n1117_lo_n,
    n1117_lo
  );


  buf

  (
    n1120_lo_p,
    n1120_lo
  );


  not

  (
    n1120_lo_n,
    n1120_lo
  );


  buf

  (
    n1129_lo_p,
    n1129_lo
  );


  not

  (
    n1129_lo_n,
    n1129_lo
  );


  buf

  (
    n1132_lo_p,
    n1132_lo
  );


  not

  (
    n1132_lo_n,
    n1132_lo
  );


  buf

  (
    n1156_lo_p,
    n1156_lo
  );


  not

  (
    n1156_lo_n,
    n1156_lo
  );


  buf

  (
    n1168_lo_p,
    n1168_lo
  );


  not

  (
    n1168_lo_n,
    n1168_lo
  );


  buf

  (
    n1180_lo_p,
    n1180_lo
  );


  not

  (
    n1180_lo_n,
    n1180_lo
  );


  buf

  (
    n1189_lo_p,
    n1189_lo
  );


  not

  (
    n1189_lo_n,
    n1189_lo
  );


  buf

  (
    n1192_lo_p,
    n1192_lo
  );


  not

  (
    n1192_lo_n,
    n1192_lo
  );


  buf

  (
    n1195_lo_p,
    n1195_lo
  );


  not

  (
    n1195_lo_n,
    n1195_lo
  );


  buf

  (
    n1201_lo_p,
    n1201_lo
  );


  not

  (
    n1201_lo_n,
    n1201_lo
  );


  buf

  (
    n1204_lo_p,
    n1204_lo
  );


  not

  (
    n1204_lo_n,
    n1204_lo
  );


  buf

  (
    n1228_lo_p,
    n1228_lo
  );


  not

  (
    n1228_lo_n,
    n1228_lo
  );


  buf

  (
    n1231_lo_p,
    n1231_lo
  );


  not

  (
    n1231_lo_n,
    n1231_lo
  );


  buf

  (
    n1234_lo_p,
    n1234_lo
  );


  not

  (
    n1234_lo_n,
    n1234_lo
  );


  buf

  (
    n1237_lo_p,
    n1237_lo
  );


  not

  (
    n1237_lo_n,
    n1237_lo
  );


  buf

  (
    n1240_lo_p,
    n1240_lo
  );


  not

  (
    n1240_lo_n,
    n1240_lo
  );


  buf

  (
    n1243_lo_p,
    n1243_lo
  );


  not

  (
    n1243_lo_n,
    n1243_lo
  );


  buf

  (
    n1249_lo_p,
    n1249_lo
  );


  not

  (
    n1249_lo_n,
    n1249_lo
  );


  buf

  (
    n1252_lo_p,
    n1252_lo
  );


  not

  (
    n1252_lo_n,
    n1252_lo
  );


  buf

  (
    n1255_lo_p,
    n1255_lo
  );


  not

  (
    n1255_lo_n,
    n1255_lo
  );


  buf

  (
    n1261_lo_p,
    n1261_lo
  );


  not

  (
    n1261_lo_n,
    n1261_lo
  );


  buf

  (
    n1264_lo_p,
    n1264_lo
  );


  not

  (
    n1264_lo_n,
    n1264_lo
  );


  buf

  (
    n1267_lo_p,
    n1267_lo
  );


  not

  (
    n1267_lo_n,
    n1267_lo
  );


  buf

  (
    n1273_lo_p,
    n1273_lo
  );


  not

  (
    n1273_lo_n,
    n1273_lo
  );


  buf

  (
    n1276_lo_p,
    n1276_lo
  );


  not

  (
    n1276_lo_n,
    n1276_lo
  );


  buf

  (
    n1279_lo_p,
    n1279_lo
  );


  not

  (
    n1279_lo_n,
    n1279_lo
  );


  buf

  (
    n1282_lo_p,
    n1282_lo
  );


  not

  (
    n1282_lo_n,
    n1282_lo
  );


  buf

  (
    n1285_lo_p,
    n1285_lo
  );


  not

  (
    n1285_lo_n,
    n1285_lo
  );


  buf

  (
    n1288_lo_p,
    n1288_lo
  );


  not

  (
    n1288_lo_n,
    n1288_lo
  );


  buf

  (
    n1291_lo_p,
    n1291_lo
  );


  not

  (
    n1291_lo_n,
    n1291_lo
  );


  buf

  (
    n1294_lo_p,
    n1294_lo
  );


  not

  (
    n1294_lo_n,
    n1294_lo
  );


  buf

  (
    n1297_lo_p,
    n1297_lo
  );


  not

  (
    n1297_lo_n,
    n1297_lo
  );


  buf

  (
    n1300_lo_p,
    n1300_lo
  );


  not

  (
    n1300_lo_n,
    n1300_lo
  );


  buf

  (
    n1303_lo_p,
    n1303_lo
  );


  not

  (
    n1303_lo_n,
    n1303_lo
  );


  buf

  (
    n1309_lo_p,
    n1309_lo
  );


  not

  (
    n1309_lo_n,
    n1309_lo
  );


  buf

  (
    n1312_lo_p,
    n1312_lo
  );


  not

  (
    n1312_lo_n,
    n1312_lo
  );


  buf

  (
    n1315_lo_p,
    n1315_lo
  );


  not

  (
    n1315_lo_n,
    n1315_lo
  );


  buf

  (
    n1318_lo_p,
    n1318_lo
  );


  not

  (
    n1318_lo_n,
    n1318_lo
  );


  buf

  (
    n1321_lo_p,
    n1321_lo
  );


  not

  (
    n1321_lo_n,
    n1321_lo
  );


  buf

  (
    n1333_lo_p,
    n1333_lo
  );


  not

  (
    n1333_lo_n,
    n1333_lo
  );


  buf

  (
    n1225_o2_p,
    n1225_o2
  );


  not

  (
    n1225_o2_n,
    n1225_o2
  );


  buf

  (
    n1229_o2_p,
    n1229_o2
  );


  not

  (
    n1229_o2_n,
    n1229_o2
  );


  buf

  (
    n1228_o2_p,
    n1228_o2
  );


  not

  (
    n1228_o2_n,
    n1228_o2
  );


  buf

  (
    n1259_o2_p,
    n1259_o2
  );


  not

  (
    n1259_o2_n,
    n1259_o2
  );


  buf

  (
    n1272_o2_p,
    n1272_o2
  );


  not

  (
    n1272_o2_n,
    n1272_o2
  );


  buf

  (
    n1269_o2_p,
    n1269_o2
  );


  not

  (
    n1269_o2_n,
    n1269_o2
  );


  buf

  (
    n1307_o2_p,
    n1307_o2
  );


  not

  (
    n1307_o2_n,
    n1307_o2
  );


  buf

  (
    n1201_o2_p,
    n1201_o2
  );


  not

  (
    n1201_o2_n,
    n1201_o2
  );


  buf

  (
    n1202_o2_p,
    n1202_o2
  );


  not

  (
    n1202_o2_n,
    n1202_o2
  );


  buf

  (
    n1203_o2_p,
    n1203_o2
  );


  not

  (
    n1203_o2_n,
    n1203_o2
  );


  buf

  (
    n1204_o2_p,
    n1204_o2
  );


  not

  (
    n1204_o2_n,
    n1204_o2
  );


  buf

  (
    n622_o2_p,
    n622_o2
  );


  not

  (
    n622_o2_n,
    n622_o2
  );


  buf

  (
    n1205_o2_p,
    n1205_o2
  );


  not

  (
    n1205_o2_n,
    n1205_o2
  );


  buf

  (
    n1206_o2_p,
    n1206_o2
  );


  not

  (
    n1206_o2_n,
    n1206_o2
  );


  buf

  (
    n497_o2_p,
    n497_o2
  );


  not

  (
    n497_o2_n,
    n497_o2
  );


  buf

  (
    n1212_o2_p,
    n1212_o2
  );


  not

  (
    n1212_o2_n,
    n1212_o2
  );


  buf

  (
    n1213_o2_p,
    n1213_o2
  );


  not

  (
    n1213_o2_n,
    n1213_o2
  );


  buf

  (
    n1214_o2_p,
    n1214_o2
  );


  not

  (
    n1214_o2_n,
    n1214_o2
  );


  buf

  (
    n1215_o2_p,
    n1215_o2
  );


  not

  (
    n1215_o2_n,
    n1215_o2
  );


  buf

  (
    n1216_o2_p,
    n1216_o2
  );


  not

  (
    n1216_o2_n,
    n1216_o2
  );


  buf

  (
    n1217_o2_p,
    n1217_o2
  );


  not

  (
    n1217_o2_n,
    n1217_o2
  );


  buf

  (
    n1218_o2_p,
    n1218_o2
  );


  not

  (
    n1218_o2_n,
    n1218_o2
  );


  buf

  (
    n1219_o2_p,
    n1219_o2
  );


  not

  (
    n1219_o2_n,
    n1219_o2
  );


  buf

  (
    n1242_o2_p,
    n1242_o2
  );


  not

  (
    n1242_o2_n,
    n1242_o2
  );


  buf

  (
    n1243_o2_p,
    n1243_o2
  );


  not

  (
    n1243_o2_n,
    n1243_o2
  );


  buf

  (
    n1273_o2_p,
    n1273_o2
  );


  not

  (
    n1273_o2_n,
    n1273_o2
  );


  buf

  (
    n1274_o2_p,
    n1274_o2
  );


  not

  (
    n1274_o2_n,
    n1274_o2
  );


  buf

  (
    n1275_o2_p,
    n1275_o2
  );


  not

  (
    n1275_o2_n,
    n1275_o2
  );


  buf

  (
    n1276_o2_p,
    n1276_o2
  );


  not

  (
    n1276_o2_n,
    n1276_o2
  );


  buf

  (
    n1277_o2_p,
    n1277_o2
  );


  not

  (
    n1277_o2_n,
    n1277_o2
  );


  buf

  (
    n1286_o2_p,
    n1286_o2
  );


  not

  (
    n1286_o2_n,
    n1286_o2
  );


  buf

  (
    n1299_o2_p,
    n1299_o2
  );


  not

  (
    n1299_o2_n,
    n1299_o2
  );


  buf

  (
    n601_o2_p,
    n601_o2
  );


  not

  (
    n601_o2_n,
    n601_o2
  );


  buf

  (
    n625_o2_p,
    n625_o2
  );


  not

  (
    n625_o2_n,
    n625_o2
  );


  buf

  (
    n463_o2_p,
    n463_o2
  );


  not

  (
    n463_o2_n,
    n463_o2
  );


  buf

  (
    lo082_buf_o2_p,
    lo082_buf_o2
  );


  not

  (
    lo082_buf_o2_n,
    lo082_buf_o2
  );


  buf

  (
    n455_o2_p,
    n455_o2
  );


  not

  (
    n455_o2_n,
    n455_o2
  );


  buf

  (
    n642_o2_p,
    n642_o2
  );


  not

  (
    n642_o2_n,
    n642_o2
  );


  buf

  (
    n459_o2_p,
    n459_o2
  );


  not

  (
    n459_o2_n,
    n459_o2
  );


  buf

  (
    n501_o2_p,
    n501_o2
  );


  not

  (
    n501_o2_n,
    n501_o2
  );


  buf

  (
    n599_o2_p,
    n599_o2
  );


  not

  (
    n599_o2_n,
    n599_o2
  );


  buf

  (
    n485_o2_p,
    n485_o2
  );


  not

  (
    n485_o2_n,
    n485_o2
  );


  buf

  (
    lo086_buf_o2_p,
    lo086_buf_o2
  );


  not

  (
    lo086_buf_o2_n,
    lo086_buf_o2
  );


  buf

  (
    lo122_buf_o2_p,
    lo122_buf_o2
  );


  not

  (
    lo122_buf_o2_n,
    lo122_buf_o2
  );


  buf

  (
    n502_o2_p,
    n502_o2
  );


  not

  (
    n502_o2_n,
    n502_o2
  );


  buf

  (
    n627_o2_p,
    n627_o2
  );


  not

  (
    n627_o2_n,
    n627_o2
  );


  buf

  (
    lo038_buf_o2_p,
    lo038_buf_o2
  );


  not

  (
    lo038_buf_o2_n,
    lo038_buf_o2
  );


  buf

  (
    lo046_buf_o2_p,
    lo046_buf_o2
  );


  not

  (
    lo046_buf_o2_n,
    lo046_buf_o2
  );


  buf

  (
    lo050_buf_o2_p,
    lo050_buf_o2
  );


  not

  (
    lo050_buf_o2_n,
    lo050_buf_o2
  );


  buf

  (
    lo058_buf_o2_p,
    lo058_buf_o2
  );


  not

  (
    lo058_buf_o2_n,
    lo058_buf_o2
  );


  buf

  (
    lo070_buf_o2_p,
    lo070_buf_o2
  );


  not

  (
    lo070_buf_o2_n,
    lo070_buf_o2
  );


  buf

  (
    lo094_buf_o2_p,
    lo094_buf_o2
  );


  not

  (
    lo094_buf_o2_n,
    lo094_buf_o2
  );


  buf

  (
    n462_o2_p,
    n462_o2
  );


  not

  (
    n462_o2_n,
    n462_o2
  );


  buf

  (
    lo006_buf_o2_p,
    lo006_buf_o2
  );


  not

  (
    lo006_buf_o2_n,
    lo006_buf_o2
  );


  buf

  (
    lo010_buf_o2_p,
    lo010_buf_o2
  );


  not

  (
    lo010_buf_o2_n,
    lo010_buf_o2
  );


  buf

  (
    lo022_buf_o2_p,
    lo022_buf_o2
  );


  not

  (
    lo022_buf_o2_n,
    lo022_buf_o2
  );


  buf

  (
    lo026_buf_o2_p,
    lo026_buf_o2
  );


  not

  (
    lo026_buf_o2_n,
    lo026_buf_o2
  );


  buf

  (
    lo030_buf_o2_p,
    lo030_buf_o2
  );


  not

  (
    lo030_buf_o2_n,
    lo030_buf_o2
  );


  buf

  (
    lo034_buf_o2_p,
    lo034_buf_o2
  );


  not

  (
    lo034_buf_o2_n,
    lo034_buf_o2
  );


  buf

  (
    lo054_buf_o2_p,
    lo054_buf_o2
  );


  not

  (
    lo054_buf_o2_n,
    lo054_buf_o2
  );


  buf

  (
    lo130_buf_o2_p,
    lo130_buf_o2
  );


  not

  (
    lo130_buf_o2_n,
    lo130_buf_o2
  );


  buf

  (
    n547_o2_p,
    n547_o2
  );


  not

  (
    n547_o2_n,
    n547_o2
  );


  buf

  (
    n424_inv_p,
    n424_inv
  );


  not

  (
    n424_inv_n,
    n424_inv
  );


  buf

  (
    n617_o2_p,
    n617_o2
  );


  not

  (
    n617_o2_n,
    n617_o2
  );


  buf

  (
    lo042_buf_o2_p,
    lo042_buf_o2
  );


  not

  (
    lo042_buf_o2_n,
    lo042_buf_o2
  );


  buf

  (
    lo062_buf_o2_p,
    lo062_buf_o2
  );


  not

  (
    lo062_buf_o2_n,
    lo062_buf_o2
  );


  buf

  (
    lo110_buf_o2_p,
    lo110_buf_o2
  );


  not

  (
    lo110_buf_o2_n,
    lo110_buf_o2
  );


  buf

  (
    n733_o2_p,
    n733_o2
  );


  not

  (
    n733_o2_n,
    n733_o2
  );


  buf

  (
    n734_o2_p,
    n734_o2
  );


  not

  (
    n734_o2_n,
    n734_o2
  );


  buf

  (
    n570_o2_p,
    n570_o2
  );


  not

  (
    n570_o2_n,
    n570_o2
  );


  buf

  (
    n461_o2_p,
    n461_o2
  );


  not

  (
    n461_o2_n,
    n461_o2
  );


  buf

  (
    n644_o2_p,
    n644_o2
  );


  not

  (
    n644_o2_n,
    n644_o2
  );


  buf

  (
    n628_o2_p,
    n628_o2
  );


  not

  (
    n628_o2_n,
    n628_o2
  );


  buf

  (
    n528_o2_p,
    n528_o2
  );


  not

  (
    n528_o2_n,
    n528_o2
  );


  buf

  (
    n460_inv_p,
    n460_inv
  );


  not

  (
    n460_inv_n,
    n460_inv
  );


  buf

  (
    lo002_buf_o2_p,
    lo002_buf_o2
  );


  not

  (
    lo002_buf_o2_n,
    lo002_buf_o2
  );


  buf

  (
    lo014_buf_o2_p,
    lo014_buf_o2
  );


  not

  (
    lo014_buf_o2_n,
    lo014_buf_o2
  );


  buf

  (
    lo018_buf_o2_p,
    lo018_buf_o2
  );


  not

  (
    lo018_buf_o2_n,
    lo018_buf_o2
  );


  buf

  (
    lo078_buf_o2_p,
    lo078_buf_o2
  );


  not

  (
    lo078_buf_o2_n,
    lo078_buf_o2
  );


  buf

  (
    lo090_buf_o2_p,
    lo090_buf_o2
  );


  not

  (
    lo090_buf_o2_n,
    lo090_buf_o2
  );


  buf

  (
    n513_o2_p,
    n513_o2
  );


  not

  (
    n513_o2_n,
    n513_o2
  );


  buf

  (
    lo102_buf_o2_p,
    lo102_buf_o2
  );


  not

  (
    lo102_buf_o2_n,
    lo102_buf_o2
  );


  buf

  (
    lo106_buf_o2_p,
    lo106_buf_o2
  );


  not

  (
    lo106_buf_o2_n,
    lo106_buf_o2
  );


  buf

  (
    n600_o2_p,
    n600_o2
  );


  not

  (
    n600_o2_n,
    n600_o2
  );


  buf

  (
    n529_o2_p,
    n529_o2
  );


  not

  (
    n529_o2_n,
    n529_o2
  );


  buf

  (
    n593_o2_p,
    n593_o2
  );


  not

  (
    n593_o2_n,
    n593_o2
  );


  buf

  (
    lo066_buf_o2_p,
    lo066_buf_o2
  );


  not

  (
    lo066_buf_o2_n,
    lo066_buf_o2
  );


  buf

  (
    n549_o2_p,
    n549_o2
  );


  not

  (
    n549_o2_n,
    n549_o2
  );


  buf

  (
    n550_o2_p,
    n550_o2
  );


  not

  (
    n550_o2_n,
    n550_o2
  );


  buf

  (
    n571_o2_p,
    n571_o2
  );


  not

  (
    n571_o2_n,
    n571_o2
  );


  buf

  (
    n572_o2_p,
    n572_o2
  );


  not

  (
    n572_o2_n,
    n572_o2
  );


  buf

  (
    n495_o2_p,
    n495_o2
  );


  not

  (
    n495_o2_n,
    n495_o2
  );


  buf

  (
    n496_o2_p,
    n496_o2
  );


  not

  (
    n496_o2_n,
    n496_o2
  );


  buf

  (
    n620_o2_p,
    n620_o2
  );


  not

  (
    n620_o2_n,
    n620_o2
  );


  buf

  (
    n482_o2_p,
    n482_o2
  );


  not

  (
    n482_o2_n,
    n482_o2
  );


  buf

  (
    lo081_buf_o2_p,
    lo081_buf_o2
  );


  not

  (
    lo081_buf_o2_n,
    lo081_buf_o2
  );


  buf

  (
    n576_o2_p,
    n576_o2
  );


  not

  (
    n576_o2_n,
    n576_o2
  );


  buf

  (
    n520_o2_p,
    n520_o2
  );


  not

  (
    n520_o2_n,
    n520_o2
  );


  buf

  (
    n521_o2_p,
    n521_o2
  );


  not

  (
    n521_o2_n,
    n521_o2
  );


  buf

  (
    n562_o2_p,
    n562_o2
  );


  not

  (
    n562_o2_n,
    n562_o2
  );


  buf

  (
    n508_o2_p,
    n508_o2
  );


  not

  (
    n508_o2_n,
    n508_o2
  );


  buf

  (
    n509_o2_p,
    n509_o2
  );


  not

  (
    n509_o2_n,
    n509_o2
  );


  buf

  (
    lo074_buf_o2_p,
    lo074_buf_o2
  );


  not

  (
    lo074_buf_o2_n,
    lo074_buf_o2
  );


  buf

  (
    n539_o2_p,
    n539_o2
  );


  not

  (
    n539_o2_n,
    n539_o2
  );


  buf

  (
    n536_o2_p,
    n536_o2
  );


  not

  (
    n536_o2_n,
    n536_o2
  );


  buf

  (
    n516_o2_p,
    n516_o2
  );


  not

  (
    n516_o2_n,
    n516_o2
  );


  buf

  (
    n491_o2_p,
    n491_o2
  );


  not

  (
    n491_o2_n,
    n491_o2
  );


  buf

  (
    n557_o2_p,
    n557_o2
  );


  not

  (
    n557_o2_n,
    n557_o2
  );


  buf

  (
    n586_o2_p,
    n586_o2
  );


  not

  (
    n586_o2_n,
    n586_o2
  );


  buf

  (
    n483_o2_p,
    n483_o2
  );


  not

  (
    n483_o2_n,
    n483_o2
  );


  buf

  (
    n484_o2_p,
    n484_o2
  );


  not

  (
    n484_o2_n,
    n484_o2
  );


  buf

  (
    lo004_buf_o2_p,
    lo004_buf_o2
  );


  not

  (
    lo004_buf_o2_n,
    lo004_buf_o2
  );


  buf

  (
    lo008_buf_o2_p,
    lo008_buf_o2
  );


  not

  (
    lo008_buf_o2_n,
    lo008_buf_o2
  );


  buf

  (
    lo020_buf_o2_p,
    lo020_buf_o2
  );


  not

  (
    lo020_buf_o2_n,
    lo020_buf_o2
  );


  buf

  (
    lo024_buf_o2_p,
    lo024_buf_o2
  );


  not

  (
    lo024_buf_o2_n,
    lo024_buf_o2
  );


  buf

  (
    lo028_buf_o2_p,
    lo028_buf_o2
  );


  not

  (
    lo028_buf_o2_n,
    lo028_buf_o2
  );


  buf

  (
    lo032_buf_o2_p,
    lo032_buf_o2
  );


  not

  (
    lo032_buf_o2_n,
    lo032_buf_o2
  );


  buf

  (
    lo052_buf_o2_p,
    lo052_buf_o2
  );


  not

  (
    lo052_buf_o2_n,
    lo052_buf_o2
  );


  buf

  (
    lo128_buf_o2_p,
    lo128_buf_o2
  );


  not

  (
    lo128_buf_o2_n,
    lo128_buf_o2
  );


  buf

  (
    lo037_buf_o2_p,
    lo037_buf_o2
  );


  not

  (
    lo037_buf_o2_n,
    lo037_buf_o2
  );


  buf

  (
    lo045_buf_o2_p,
    lo045_buf_o2
  );


  not

  (
    lo045_buf_o2_n,
    lo045_buf_o2
  );


  buf

  (
    lo049_buf_o2_p,
    lo049_buf_o2
  );


  not

  (
    lo049_buf_o2_n,
    lo049_buf_o2
  );


  buf

  (
    lo057_buf_o2_p,
    lo057_buf_o2
  );


  not

  (
    lo057_buf_o2_n,
    lo057_buf_o2
  );


  buf

  (
    lo069_buf_o2_p,
    lo069_buf_o2
  );


  not

  (
    lo069_buf_o2_n,
    lo069_buf_o2
  );


  buf

  (
    lo093_buf_o2_p,
    lo093_buf_o2
  );


  not

  (
    lo093_buf_o2_n,
    lo093_buf_o2
  );


  and

  (
    g218_p,
    n461_o2_n_spl_,
    n628_o2_p_spl_
  );


  or

  (
    g218_n,
    n461_o2_p_spl_,
    n628_o2_n_spl_
  );


  and

  (
    g219_p,
    n949_lo_n,
    g218_n_spl_00
  );


  and

  (
    g220_p,
    n949_lo_p,
    g218_p_spl_00
  );


  or

  (
    g221_n,
    g219_p,
    g220_p
  );


  and

  (
    g222_p,
    n961_lo_n,
    g218_n_spl_00
  );


  and

  (
    g223_p,
    n961_lo_p,
    g218_p_spl_00
  );


  or

  (
    g224_n,
    g222_p,
    g223_p
  );


  and

  (
    g225_p,
    n973_lo_n,
    g218_n_spl_01
  );


  and

  (
    g226_p,
    n973_lo_p,
    g218_p_spl_01
  );


  or

  (
    g227_n,
    g225_p,
    g226_p
  );


  and

  (
    g228_p,
    n985_lo_n,
    g218_n_spl_01
  );


  and

  (
    g229_p,
    n985_lo_p,
    g218_p_spl_01
  );


  or

  (
    g230_n,
    g228_p,
    g229_p
  );


  and

  (
    g231_p,
    n644_o2_n_spl_0,
    n628_o2_p_spl_
  );


  or

  (
    g231_n,
    n644_o2_p_spl_0,
    n628_o2_n_spl_
  );


  and

  (
    g232_p,
    n1057_lo_n,
    g231_n_spl_00
  );


  and

  (
    g233_p,
    n1057_lo_p,
    g231_p_spl_00
  );


  or

  (
    g234_n,
    g232_p,
    g233_p
  );


  and

  (
    g235_p,
    n1117_lo_n,
    g231_n_spl_00
  );


  and

  (
    g236_p,
    n1117_lo_p,
    g231_p_spl_00
  );


  or

  (
    g237_n,
    g235_p,
    g236_p
  );


  and

  (
    g238_p,
    n1129_lo_n,
    g231_n_spl_01
  );


  and

  (
    g239_p,
    n1129_lo_p,
    g231_p_spl_01
  );


  or

  (
    g240_n,
    g238_p,
    g239_p
  );


  and

  (
    g241_p,
    n463_o2_p,
    n501_o2_n_spl_
  );


  or

  (
    g241_n,
    n463_o2_n_spl_,
    n501_o2_p
  );


  and

  (
    g242_p,
    n627_o2_p,
    g241_p
  );


  or

  (
    g242_n,
    n627_o2_n,
    g241_n
  );


  and

  (
    g243_p,
    n461_o2_n_spl_,
    g242_p_spl_
  );


  or

  (
    g243_n,
    n461_o2_p_spl_,
    g242_n_spl_
  );


  and

  (
    g244_p,
    n997_lo_n,
    g243_n_spl_0
  );


  and

  (
    g245_p,
    n997_lo_p,
    g243_p_spl_0
  );


  or

  (
    g246_n,
    g244_p,
    g245_p
  );


  and

  (
    g247_p,
    n1009_lo_n,
    g243_n_spl_0
  );


  and

  (
    g248_p,
    n1009_lo_p,
    g243_p_spl_0
  );


  or

  (
    g249_n,
    g247_p,
    g248_p
  );


  and

  (
    g250_p,
    n1021_lo_n,
    g243_n_spl_1
  );


  and

  (
    g251_p,
    n1021_lo_p,
    g243_p_spl_1
  );


  or

  (
    g252_n,
    g250_p,
    g251_p
  );


  and

  (
    g253_p,
    n1033_lo_n,
    g243_n_spl_1
  );


  and

  (
    g254_p,
    n1033_lo_p,
    g243_p_spl_1
  );


  or

  (
    g255_n,
    g253_p,
    g254_p
  );


  and

  (
    g256_p,
    n644_o2_n_spl_0,
    g242_p_spl_
  );


  or

  (
    g256_n,
    n644_o2_p_spl_0,
    g242_n_spl_
  );


  and

  (
    g257_p,
    n1045_lo_p,
    g256_p
  );


  and

  (
    g258_p,
    n1045_lo_n,
    g256_n
  );


  or

  (
    g259_n,
    g257_p,
    g258_p
  );


  and

  (
    g260_p,
    n601_o2_p,
    n644_o2_n_spl_
  );


  or

  (
    g260_n,
    n601_o2_n_spl_,
    n644_o2_p_spl_
  );


  and

  (
    g261_p,
    n625_o2_p_spl_,
    g260_p
  );


  or

  (
    g261_n,
    n625_o2_n,
    g260_n
  );


  and

  (
    g262_p,
    n502_o2_n,
    g261_p
  );


  or

  (
    g262_n,
    n502_o2_p,
    g261_n
  );


  and

  (
    g263_p,
    n599_o2_p_spl_,
    g262_p
  );


  or

  (
    g263_n,
    n599_o2_n,
    g262_n
  );


  and

  (
    g264_p,
    n1069_lo_n,
    g263_n_spl_0
  );


  and

  (
    g265_p,
    n1069_lo_p,
    g263_p_spl_0
  );


  or

  (
    g266_n,
    g264_p,
    g265_p
  );


  and

  (
    g267_p,
    n1081_lo_n,
    g263_n_spl_0
  );


  and

  (
    g268_p,
    n1081_lo_p,
    g263_p_spl_0
  );


  or

  (
    g269_n,
    g267_p,
    g268_p
  );


  and

  (
    g270_p,
    n1093_lo_n,
    g263_n_spl_1
  );


  and

  (
    g271_p,
    n1093_lo_p,
    g263_p_spl_1
  );


  or

  (
    g272_n,
    g270_p,
    g271_p
  );


  and

  (
    g273_p,
    n1105_lo_n,
    g263_n_spl_1
  );


  and

  (
    g274_p,
    n1105_lo_p,
    g263_p_spl_1
  );


  or

  (
    g275_n,
    g273_p,
    g274_p
  );


  and

  (
    g276_p,
    g218_n_spl_10,
    g231_n_spl_01
  );


  or

  (
    g276_n,
    g218_p_spl_10,
    g231_p_spl_01
  );


  and

  (
    g277_p,
    n1321_lo_p,
    g276_n_spl_00
  );


  and

  (
    g278_p,
    n601_o2_n_spl_,
    n463_o2_n_spl_
  );


  and

  (
    g279_p,
    n501_o2_n_spl_,
    g278_p
  );


  and

  (
    g280_p,
    n625_o2_p_spl_,
    g279_p
  );


  and

  (
    g281_p,
    n599_o2_p_spl_,
    g280_p
  );


  or

  (
    g282_n,
    n1333_lo_p_spl_0,
    g281_p
  );


  or

  (
    g283_n,
    g277_p,
    g282_n
  );


  and

  (
    g284_p,
    n1309_lo_n_spl_00,
    n622_o2_p
  );


  or

  (
    g284_n,
    n1309_lo_p_spl_0,
    n622_o2_n
  );


  and

  (
    g285_p,
    g276_n_spl_00,
    g284_p
  );


  or

  (
    g285_n,
    g276_p_spl_0,
    g284_n
  );


  and

  (
    g286_p,
    n1307_o2_n,
    g285_n
  );


  and

  (
    g287_p,
    n1307_o2_p,
    g285_p
  );


  or

  (
    g288_n,
    g286_p,
    g287_p
  );


  and

  (
    g289_p,
    n459_o2_p_spl_00,
    g288_n
  );


  and

  (
    g290_p,
    n1237_lo_p,
    n1309_lo_n_spl_00
  );


  or

  (
    g290_n,
    n1237_lo_n,
    n1309_lo_p_spl_0
  );


  and

  (
    g291_p,
    g276_n_spl_01,
    g290_p
  );


  or

  (
    g291_n,
    g276_p_spl_0,
    g290_n
  );


  and

  (
    g292_p,
    n497_o2_p,
    g291_n
  );


  and

  (
    g293_p,
    n497_o2_n,
    g291_p
  );


  or

  (
    g294_n,
    g292_p,
    g293_p
  );


  and

  (
    g295_p,
    n459_o2_p_spl_00,
    g294_n
  );


  and

  (
    g296_p,
    n1261_lo_p,
    n1309_lo_n_spl_0
  );


  and

  (
    g297_p,
    g276_n_spl_01,
    g296_p
  );


  or

  (
    g298_n,
    n1269_o2_n,
    g297_p
  );


  and

  (
    g299_p,
    n459_o2_p_spl_01,
    g298_n
  );


  and

  (
    g300_p,
    n1273_lo_p,
    n1309_lo_n_spl_1
  );


  and

  (
    g301_p,
    g276_n_spl_1,
    g300_p
  );


  or

  (
    g302_n,
    n1225_o2_n,
    g301_p
  );


  and

  (
    g303_p,
    n459_o2_p_spl_01,
    g302_n
  );


  and

  (
    g304_p,
    n1309_lo_n_spl_1,
    n1259_o2_p
  );


  and

  (
    g305_p,
    g276_n_spl_1,
    g304_p
  );


  or

  (
    g306_n,
    n1228_o2_p,
    g305_p
  );


  and

  (
    g307_p,
    n459_o2_p_spl_1,
    g306_n
  );


  and

  (
    g308_p,
    n1189_lo_p,
    n1285_lo_p
  );


  or

  (
    g308_n,
    n1189_lo_n,
    n1285_lo_n
  );


  and

  (
    g309_p,
    n1333_lo_n_spl_,
    g308_n
  );


  or

  (
    g309_n,
    n1333_lo_p_spl_0,
    g308_p
  );


  and

  (
    g310_p,
    n1229_o2_p,
    n455_o2_p
  );


  or

  (
    g310_n,
    n1229_o2_n,
    n455_o2_n
  );


  and

  (
    g311_p,
    g218_p_spl_10,
    g310_n_spl_
  );


  or

  (
    g311_n,
    g218_n_spl_10,
    g310_p_spl_
  );


  and

  (
    g312_p,
    g218_n_spl_1,
    g310_p_spl_
  );


  or

  (
    g312_n,
    g218_p_spl_1,
    g310_n_spl_
  );


  and

  (
    g313_p,
    g311_n,
    g312_n
  );


  or

  (
    g313_n,
    g311_p,
    g312_p
  );


  and

  (
    g314_p,
    g309_n,
    g313_n
  );


  and

  (
    g315_p,
    g309_p,
    g313_p
  );


  or

  (
    g316_n,
    g314_p,
    g315_p
  );


  and

  (
    g317_p,
    n1201_lo_p,
    n1297_lo_p
  );


  or

  (
    g317_n,
    n1201_lo_n,
    n1297_lo_n
  );


  and

  (
    g318_p,
    n1333_lo_n_spl_,
    g317_n
  );


  or

  (
    g318_n,
    n1333_lo_p_spl_,
    g317_p
  );


  and

  (
    g319_p,
    n733_o2_n,
    n734_o2_n
  );


  or

  (
    g319_n,
    n733_o2_p,
    n734_o2_p
  );


  and

  (
    g320_p,
    n642_o2_p,
    g319_n
  );


  or

  (
    g320_n,
    n642_o2_n,
    g319_p
  );


  and

  (
    g321_p,
    g231_p_spl_1,
    g320_n_spl_
  );


  or

  (
    g321_n,
    g231_n_spl_1,
    g320_p_spl_
  );


  and

  (
    g322_p,
    g231_n_spl_1,
    g320_p_spl_
  );


  or

  (
    g322_n,
    g231_p_spl_1,
    g320_n_spl_
  );


  and

  (
    g323_p,
    g321_n,
    g322_n
  );


  or

  (
    g323_n,
    g321_p,
    g322_p
  );


  and

  (
    g324_p,
    g318_n,
    g323_n
  );


  and

  (
    g325_p,
    g318_p,
    g323_p
  );


  or

  (
    g326_n,
    g324_p,
    g325_p
  );


  or

  (
    g327_n,
    n1249_lo_n,
    n1309_lo_p_spl_
  );


  or

  (
    g328_n,
    g276_p_spl_,
    g327_n
  );


  and

  (
    g329_p,
    n1272_o2_n,
    g328_n
  );


  and

  (
    g330_p,
    n459_o2_p_spl_1,
    g329_p
  );


  and

  (
    g331_p,
    n1299_o2_p,
    n600_o2_p
  );


  or

  (
    g331_n,
    n1299_o2_n,
    n600_o2_n_spl_
  );


  and

  (
    g332_p,
    n495_o2_n,
    n496_o2_n
  );


  or

  (
    g332_n,
    n495_o2_p,
    n496_o2_p
  );


  or

  (
    g333_n,
    n1205_o2_n,
    n600_o2_n_spl_
  );


  and

  (
    g334_p,
    lo122_buf_o2_n_spl_,
    n620_o2_n
  );


  or

  (
    g334_n,
    lo122_buf_o2_p_spl_0,
    n620_o2_p_spl_
  );


  or

  (
    g335_n,
    g331_p_spl_,
    g334_n
  );


  or

  (
    g336_n,
    g331_n,
    g334_p
  );


  and

  (
    g337_p,
    g335_n,
    g336_n
  );


  or

  (
    g338_n,
    n1276_o2_n,
    n462_o2_n
  );


  or

  (
    g339_n,
    n1282_lo_p_spl_,
    n1219_o2_p_spl_0
  );


  or

  (
    g340_n,
    n1294_lo_p_spl_,
    n1219_o2_p_spl_0
  );


  or

  (
    g341_n,
    n1318_lo_p_spl_,
    n1219_o2_p_spl_1
  );


  and

  (
    g342_p,
    lo122_buf_o2_n_spl_,
    g332_n_spl_
  );


  or

  (
    g342_n,
    lo122_buf_o2_p_spl_0,
    g332_p
  );


  or

  (
    g343_n,
    n1234_lo_p_spl_,
    g342_n
  );


  or

  (
    g344_n,
    n1234_lo_n,
    g342_p
  );


  and

  (
    g345_p,
    g343_n,
    g344_n
  );


  or

  (
    g346_n,
    lo106_buf_o2_p_spl_,
    n529_o2_n
  );


  and

  (
    g347_p,
    n549_o2_n,
    n550_o2_n
  );


  and

  (
    g348_p,
    n571_o2_p,
    n572_o2_n
  );


  and

  (
    g349_p,
    g347_p,
    g348_p
  );


  and

  (
    g350_p,
    g346_n,
    g349_p
  );


  or

  (
    g351_n,
    lo102_buf_o2_n,
    n593_o2_n
  );


  or

  (
    g352_n,
    lo102_buf_o2_p_spl_,
    n593_o2_p
  );


  or

  (
    g353_n,
    lo106_buf_o2_n,
    n529_o2_p
  );


  and

  (
    g354_p,
    g352_n,
    g353_n
  );


  and

  (
    g355_p,
    g351_n,
    g354_p
  );


  and

  (
    g356_p,
    g350_p,
    g355_p
  );


  and

  (
    g357_p,
    n483_o2_n,
    n484_o2_n
  );


  or

  (
    g357_n,
    n483_o2_p,
    n484_o2_p
  );


  or

  (
    g358_n,
    g338_n_spl_,
    g345_p_spl_
  );


  or

  (
    g359_n,
    g333_n_spl_,
    g337_p_spl_
  );


  and

  (
    g360_p,
    g356_p_spl_,
    g359_n
  );


  or

  (
    g361_n,
    n1303_lo_p_spl_0,
    lo090_buf_o2_p_spl_0
  );


  and

  (
    g362_p,
    n539_o2_n_spl_,
    n536_o2_p_spl_
  );


  or

  (
    g362_n,
    n539_o2_p_spl_,
    n536_o2_n_spl_
  );


  and

  (
    g363_p,
    n539_o2_p_spl_,
    n536_o2_n_spl_
  );


  or

  (
    g363_n,
    n539_o2_n_spl_,
    n536_o2_p_spl_
  );


  and

  (
    g364_p,
    g362_n,
    g363_n
  );


  or

  (
    g364_n,
    g362_p,
    g363_p
  );


  and

  (
    g365_p,
    lo090_buf_o2_n,
    lo074_buf_o2_p_spl_
  );


  or

  (
    g365_n,
    lo090_buf_o2_p_spl_0,
    lo074_buf_o2_n
  );


  and

  (
    g366_p,
    lo130_buf_o2_n_spl_0,
    g365_p
  );


  or

  (
    g366_n,
    lo130_buf_o2_p_spl_00,
    g365_n
  );


  and

  (
    g367_p,
    g364_n,
    g366_n
  );


  and

  (
    g368_p,
    g364_p,
    g366_p
  );


  or

  (
    g369_n,
    g367_p,
    g368_p
  );


  and

  (
    g370_p,
    n516_o2_n_spl_0,
    n557_o2_p_spl_
  );


  or

  (
    g370_n,
    n516_o2_p_spl_0,
    n557_o2_n_spl_
  );


  and

  (
    g371_p,
    n516_o2_p_spl_0,
    n557_o2_n_spl_
  );


  or

  (
    g371_n,
    n516_o2_n_spl_0,
    n557_o2_p_spl_
  );


  and

  (
    g372_p,
    g370_n,
    g371_n
  );


  or

  (
    g372_n,
    g370_p,
    g371_p
  );


  and

  (
    g373_p,
    lo050_buf_o2_n_spl_,
    n562_o2_p_spl_
  );


  or

  (
    g373_n,
    lo050_buf_o2_p_spl_0,
    n562_o2_n_spl_
  );


  and

  (
    g374_p,
    lo050_buf_o2_p_spl_0,
    n562_o2_n_spl_
  );


  or

  (
    g374_n,
    lo050_buf_o2_n_spl_,
    n562_o2_p_spl_
  );


  and

  (
    g375_p,
    g373_n,
    g374_n
  );


  or

  (
    g375_n,
    g373_p,
    g374_p
  );


  or

  (
    g376_n,
    g372_p,
    g375_p
  );


  or

  (
    g377_n,
    g372_n,
    g375_n
  );


  and

  (
    g378_p,
    g376_n,
    g377_n
  );


  and

  (
    g379_p,
    n491_o2_p_spl_0,
    n586_o2_p_spl_0
  );


  or

  (
    g379_n,
    n491_o2_n_spl_0,
    n586_o2_n_spl_0
  );


  and

  (
    g380_p,
    n491_o2_n_spl_0,
    n586_o2_n_spl_0
  );


  or

  (
    g380_n,
    n491_o2_p_spl_0,
    n586_o2_p_spl_0
  );


  and

  (
    g381_p,
    g379_n,
    g380_n
  );


  or

  (
    g381_n,
    g379_p,
    g380_p
  );


  and

  (
    g382_p,
    lo030_buf_o2_n_spl_,
    lo014_buf_o2_p_spl_00
  );


  or

  (
    g382_n,
    lo030_buf_o2_p_spl_0,
    lo014_buf_o2_n_spl_0
  );


  and

  (
    g383_p,
    lo030_buf_o2_p_spl_0,
    lo014_buf_o2_n_spl_0
  );


  or

  (
    g383_n,
    lo030_buf_o2_n_spl_,
    lo014_buf_o2_p_spl_00
  );


  and

  (
    g384_p,
    g382_n,
    g383_n
  );


  or

  (
    g384_n,
    g382_p,
    g383_p
  );


  and

  (
    g385_p,
    g381_n_spl_,
    g384_p_spl_
  );


  or

  (
    g385_n,
    g381_p_spl_,
    g384_n_spl_
  );


  and

  (
    g386_p,
    g381_p_spl_,
    g384_n_spl_
  );


  or

  (
    g386_n,
    g381_n_spl_,
    g384_p_spl_
  );


  and

  (
    g387_p,
    g385_n,
    g386_n
  );


  or

  (
    g387_n,
    g385_p,
    g386_p
  );


  and

  (
    g388_p,
    n1286_o2_n,
    n485_o2_p
  );


  and

  (
    g389_p,
    n1286_o2_p,
    n485_o2_n
  );


  and

  (
    g390_p,
    lo074_buf_o2_p_spl_,
    g361_n_spl_
  );


  and

  (
    g391_p,
    n1206_o2_p,
    n1277_o2_n
  );


  or

  (
    g392_n,
    lo122_buf_o2_p_spl_1,
    g391_p_spl_
  );


  or

  (
    g393_n,
    g339_n_spl_,
    g392_n_spl_
  );


  or

  (
    g394_n,
    g341_n_spl_,
    g391_p_spl_
  );


  and

  (
    g395_p,
    g393_n,
    g394_n_spl_
  );


  or

  (
    g396_n,
    g340_n_spl_,
    g392_n_spl_
  );


  and

  (
    g397_p,
    g394_n_spl_,
    g396_n
  );


  and

  (
    g398_p,
    g358_n_spl_,
    g360_p_spl_
  );


  and

  (
    g399_p,
    n508_o2_n,
    n509_o2_n
  );


  or

  (
    g399_n,
    n508_o2_p,
    n509_o2_p
  );


  and

  (
    g400_p,
    n516_o2_p_spl_1,
    g399_p_spl_
  );


  or

  (
    g400_n,
    n516_o2_n_spl_1,
    g399_n_spl_
  );


  and

  (
    g401_p,
    n516_o2_n_spl_1,
    g399_n_spl_
  );


  or

  (
    g401_n,
    n516_o2_p_spl_1,
    g399_p_spl_
  );


  and

  (
    g402_p,
    g400_n,
    g401_n
  );


  or

  (
    g402_n,
    g400_p,
    g401_p
  );


  and

  (
    g403_p,
    n520_o2_n,
    n521_o2_n
  );


  or

  (
    g403_n,
    n520_o2_p,
    n521_o2_p
  );


  and

  (
    g404_p,
    lo006_buf_o2_n_spl_,
    g403_n_spl_
  );


  or

  (
    g404_n,
    lo006_buf_o2_p_spl_0,
    g403_p_spl_
  );


  and

  (
    g405_p,
    lo006_buf_o2_p_spl_0,
    g403_p_spl_
  );


  or

  (
    g405_n,
    lo006_buf_o2_n_spl_,
    g403_n_spl_
  );


  and

  (
    g406_p,
    g404_n,
    g405_n
  );


  or

  (
    g406_n,
    g404_p,
    g405_p
  );


  and

  (
    g407_p,
    g402_n,
    g406_p
  );


  and

  (
    g408_p,
    g402_p,
    g406_n
  );


  or

  (
    g409_n,
    g407_p,
    g408_p
  );


  and

  (
    g410_p,
    lo130_buf_o2_n_spl_0,
    n576_o2_p
  );


  or

  (
    g410_n,
    lo130_buf_o2_p_spl_00,
    n576_o2_n
  );


  and

  (
    g411_p,
    lo002_buf_o2_p_spl_0,
    g410_p_spl_
  );


  or

  (
    g411_n,
    lo002_buf_o2_n_spl_,
    g410_n_spl_
  );


  and

  (
    g412_p,
    lo002_buf_o2_n_spl_,
    g410_n_spl_
  );


  or

  (
    g412_n,
    lo002_buf_o2_p_spl_0,
    g410_p_spl_
  );


  and

  (
    g413_p,
    g411_n,
    g412_n
  );


  or

  (
    g413_n,
    g411_p,
    g412_p
  );


  and

  (
    g414_p,
    n586_o2_p_spl_1,
    g357_p_spl_0
  );


  or

  (
    g414_n,
    n586_o2_n_spl_1,
    g357_n_spl_0
  );


  and

  (
    g415_p,
    n586_o2_n_spl_1,
    g357_n_spl_0
  );


  or

  (
    g415_n,
    n586_o2_p_spl_1,
    g357_p_spl_0
  );


  and

  (
    g416_p,
    g414_n,
    g415_n
  );


  or

  (
    g416_n,
    g414_p,
    g415_p
  );


  and

  (
    g417_p,
    g413_p,
    g416_n
  );


  and

  (
    g418_p,
    g413_n,
    g416_p
  );


  or

  (
    g419_n,
    g417_p,
    g418_p
  );


  and

  (
    g420_p,
    lo032_buf_o2_n_spl_,
    lo052_buf_o2_n_spl_
  );


  or

  (
    g420_n,
    lo032_buf_o2_p_spl_0,
    lo052_buf_o2_p_spl_0
  );


  and

  (
    g421_p,
    lo032_buf_o2_p_spl_0,
    lo052_buf_o2_p_spl_0
  );


  or

  (
    g421_n,
    lo032_buf_o2_n_spl_,
    lo052_buf_o2_n_spl_
  );


  and

  (
    g422_p,
    g420_n,
    g421_n
  );


  or

  (
    g422_n,
    g420_p,
    g421_p
  );


  or

  (
    g423_n,
    n1303_lo_p_spl_0,
    lo094_buf_o2_p_spl_
  );


  and

  (
    g424_p,
    n1303_lo_n_spl_0,
    g409_n_spl_
  );


  and

  (
    g425_p,
    n1303_lo_n_spl_0,
    g419_n_spl_
  );


  and

  (
    g426_p,
    n1303_lo_n_spl_,
    g369_n_spl_
  );


  and

  (
    g427_p,
    n1267_lo_n_spl_,
    g426_p_spl_
  );


  or

  (
    g428_n,
    n1267_lo_n_spl_,
    g426_p_spl_
  );


  or

  (
    g429_n,
    n1303_lo_p_spl_1,
    g378_p_spl_
  );


  or

  (
    g430_n,
    g390_p_spl_0,
    g429_n_spl_
  );


  and

  (
    g431_p,
    g390_p_spl_0,
    g429_n_spl_
  );


  and

  (
    g432_p,
    n1195_lo_p_spl_,
    lo130_buf_o2_n_spl_1
  );


  or

  (
    g432_n,
    n1195_lo_n,
    lo130_buf_o2_p_spl_0
  );


  and

  (
    g433_p,
    lo054_buf_o2_n_spl_,
    lo014_buf_o2_n_spl_1
  );


  or

  (
    g433_n,
    lo054_buf_o2_p_spl_0,
    lo014_buf_o2_p_spl_0
  );


  and

  (
    g434_p,
    lo054_buf_o2_p_spl_0,
    lo014_buf_o2_p_spl_1
  );


  or

  (
    g434_n,
    lo054_buf_o2_n_spl_,
    lo014_buf_o2_n_spl_1
  );


  and

  (
    g435_p,
    g433_n,
    g434_n
  );


  or

  (
    g435_n,
    g433_p,
    g434_p
  );


  and

  (
    g436_p,
    g432_p,
    g435_n
  );


  and

  (
    g437_p,
    g432_n,
    g435_p
  );


  or

  (
    g438_n,
    g436_p,
    g437_p
  );


  or

  (
    g439_n,
    n491_o2_n_spl_,
    g357_n_spl_1
  );


  or

  (
    g440_n,
    n491_o2_p_spl_,
    g357_p_spl_
  );


  and

  (
    g441_p,
    g439_n,
    g440_n
  );


  and

  (
    g442_p,
    g438_n_spl_,
    g441_p_spl_
  );


  or

  (
    g443_n,
    g438_n_spl_,
    g441_p_spl_
  );


  and

  (
    g444_p,
    lo130_buf_o2_n_spl_1,
    lo081_buf_o2_p_spl_
  );


  or

  (
    g444_n,
    lo130_buf_o2_p_spl_1,
    lo081_buf_o2_n
  );


  and

  (
    g445_p,
    lo034_buf_o2_p_spl_0,
    n482_o2_n_spl_
  );


  or

  (
    g445_n,
    lo034_buf_o2_n_spl_,
    n482_o2_p_spl_
  );


  and

  (
    g446_p,
    lo034_buf_o2_n_spl_,
    n482_o2_p_spl_
  );


  or

  (
    g446_n,
    lo034_buf_o2_p_spl_0,
    n482_o2_n_spl_
  );


  and

  (
    g447_p,
    g445_n,
    g446_n
  );


  or

  (
    g447_n,
    g445_p,
    g446_p
  );


  and

  (
    g448_p,
    g444_p_spl_,
    g447_n_spl_
  );


  or

  (
    g448_n,
    g444_n_spl_,
    g447_p_spl_
  );


  and

  (
    g449_p,
    g444_n_spl_,
    g447_p_spl_
  );


  or

  (
    g449_n,
    g444_p_spl_,
    g447_n_spl_
  );


  and

  (
    g450_p,
    g448_n,
    g449_n
  );


  or

  (
    g450_n,
    g448_p,
    g449_p
  );


  and

  (
    g451_p,
    g387_n,
    g450_p
  );


  and

  (
    g452_p,
    g387_p_spl_,
    g450_n
  );


  or

  (
    g453_n,
    g451_p,
    g452_p
  );


  and

  (
    g454_p,
    lo037_buf_o2_p_spl_00,
    lo057_buf_o2_n_spl_0
  );


  or

  (
    g454_n,
    lo037_buf_o2_n_spl_0,
    lo057_buf_o2_p_spl_0
  );


  and

  (
    g455_p,
    lo037_buf_o2_n_spl_0,
    lo057_buf_o2_p_spl_0
  );


  or

  (
    g455_n,
    lo037_buf_o2_p_spl_00,
    lo057_buf_o2_n_spl_0
  );


  and

  (
    g456_p,
    g454_n,
    g455_n
  );


  or

  (
    g456_n,
    g454_p,
    g455_p
  );


  and

  (
    g457_p,
    n1120_lo_p_spl_0,
    g456_n_spl_
  );


  and

  (
    g458_p,
    n1120_lo_n_spl_,
    g456_p_spl_
  );


  or

  (
    g459_n,
    g457_p,
    g458_p
  );


  and

  (
    g460_p,
    n1132_lo_p_spl_,
    lo093_buf_o2_n_spl_
  );


  and

  (
    g461_p,
    n988_lo_p_spl_0,
    lo028_buf_o2_n_spl_0
  );


  and

  (
    g462_p,
    n988_lo_n_spl_,
    lo028_buf_o2_p_spl_0
  );


  and

  (
    g463_p,
    n1168_lo_p_spl_,
    n1204_lo_n
  );


  and

  (
    g464_p,
    lo128_buf_o2_n_spl_,
    g463_p
  );


  and

  (
    g465_p,
    lo069_buf_o2_p_spl_,
    lo093_buf_o2_n_spl_
  );


  or

  (
    g465_n,
    lo069_buf_o2_n,
    lo093_buf_o2_p_spl_
  );


  and

  (
    g466_p,
    lo128_buf_o2_n_spl_,
    g465_p
  );


  or

  (
    g466_n,
    lo128_buf_o2_p_spl_,
    g465_n
  );


  and

  (
    g467_p,
    lo057_buf_o2_p_spl_1,
    g466_n
  );


  and

  (
    g468_p,
    lo057_buf_o2_n_spl_,
    g466_p
  );


  or

  (
    g469_n,
    g467_p,
    g468_p
  );


  and

  (
    g470_p,
    n1060_lo_n_spl_0,
    g469_n_spl_
  );


  or

  (
    g471_n,
    n1060_lo_n_spl_0,
    g469_n_spl_
  );


  and

  (
    g472_p,
    lo045_buf_o2_n_spl_0,
    g456_n_spl_
  );


  and

  (
    g473_p,
    lo045_buf_o2_p_spl_0,
    g456_p_spl_
  );


  or

  (
    g474_n,
    g472_p,
    g473_p
  );


  and

  (
    g475_p,
    lo020_buf_o2_p_spl_00,
    lo028_buf_o2_n_spl_0
  );


  or

  (
    g475_n,
    lo020_buf_o2_n_spl_0,
    lo028_buf_o2_p_spl_0
  );


  and

  (
    g476_p,
    lo020_buf_o2_n_spl_0,
    lo028_buf_o2_p_spl_1
  );


  or

  (
    g476_n,
    lo020_buf_o2_p_spl_00,
    lo028_buf_o2_n_spl_
  );


  and

  (
    g477_p,
    g475_n,
    g476_n
  );


  or

  (
    g477_n,
    g475_p,
    g476_p
  );


  and

  (
    g478_p,
    lo008_buf_o2_n_spl_0,
    g477_n
  );


  and

  (
    g479_p,
    lo008_buf_o2_p_spl_0,
    g477_p
  );


  or

  (
    g480_n,
    g478_p,
    g479_p
  );


  and

  (
    g481_p,
    n1120_lo_p_spl_0,
    g422_n
  );


  and

  (
    g482_p,
    n1120_lo_n_spl_,
    g422_p_spl_
  );


  or

  (
    g483_n,
    g481_p,
    g482_p
  );


  and

  (
    g484_p,
    lo004_buf_o2_n_spl_,
    lo008_buf_o2_n_spl_0
  );


  or

  (
    g484_n,
    lo004_buf_o2_p_spl_0,
    lo008_buf_o2_p_spl_0
  );


  and

  (
    g485_p,
    lo004_buf_o2_p_spl_0,
    lo008_buf_o2_p_spl_1
  );


  or

  (
    g485_n,
    lo004_buf_o2_n_spl_,
    lo008_buf_o2_n_spl_
  );


  and

  (
    g486_p,
    g484_n,
    g485_n
  );


  or

  (
    g486_n,
    g484_p,
    g485_p
  );


  and

  (
    g487_p,
    n940_lo_p_spl_,
    g486_n
  );


  and

  (
    g488_p,
    n940_lo_n,
    g486_p
  );


  or

  (
    g489_n,
    g487_p,
    g488_p
  );


  and

  (
    g490_p,
    lo024_buf_o2_p_spl_00,
    lo037_buf_o2_n_spl_1
  );


  or

  (
    g490_n,
    lo024_buf_o2_n_spl_0,
    lo037_buf_o2_p_spl_0
  );


  and

  (
    g491_p,
    lo024_buf_o2_n_spl_0,
    lo037_buf_o2_p_spl_1
  );


  or

  (
    g491_n,
    lo024_buf_o2_p_spl_00,
    lo037_buf_o2_n_spl_1
  );


  and

  (
    g492_p,
    g490_n,
    g491_n
  );


  or

  (
    g492_n,
    g490_p,
    g491_p
  );


  and

  (
    g493_p,
    n976_lo_n,
    g492_n
  );


  and

  (
    g494_p,
    n976_lo_p_spl_,
    g492_p
  );


  or

  (
    g495_n,
    g493_p,
    g494_p
  );


  and

  (
    g496_p,
    lo020_buf_o2_n_spl_1,
    lo024_buf_o2_n_spl_1
  );


  or

  (
    g496_n,
    lo020_buf_o2_p_spl_0,
    lo024_buf_o2_p_spl_0
  );


  and

  (
    g497_p,
    lo020_buf_o2_p_spl_1,
    lo024_buf_o2_p_spl_1
  );


  or

  (
    g497_n,
    lo020_buf_o2_n_spl_1,
    lo024_buf_o2_n_spl_1
  );


  and

  (
    g498_p,
    g496_n,
    g497_n
  );


  or

  (
    g498_n,
    g496_p,
    g497_p
  );


  and

  (
    g499_p,
    n988_lo_p_spl_0,
    g498_n
  );


  and

  (
    g500_p,
    n988_lo_n_spl_,
    g498_p
  );


  or

  (
    g501_n,
    g499_p,
    g500_p
  );


  and

  (
    g502_p,
    lo045_buf_o2_n_spl_0,
    lo049_buf_o2_n_spl_
  );


  or

  (
    g502_n,
    lo045_buf_o2_p_spl_0,
    lo049_buf_o2_p_spl_0
  );


  and

  (
    g503_p,
    lo045_buf_o2_p_spl_1,
    lo049_buf_o2_p_spl_0
  );


  or

  (
    g503_n,
    lo045_buf_o2_n_spl_,
    lo049_buf_o2_n_spl_
  );


  and

  (
    g504_p,
    g502_n,
    g503_n
  );


  or

  (
    g504_n,
    g502_p,
    g503_p
  );


  and

  (
    g505_p,
    n1060_lo_p_spl_,
    g504_n
  );


  and

  (
    g506_p,
    n1060_lo_n_spl_,
    g504_p
  );


  or

  (
    g507_n,
    g505_p,
    g506_p
  );


  and

  (
    g508_p,
    g459_n_spl_0,
    g507_n_spl_
  );


  or

  (
    g509_n,
    g459_n_spl_0,
    g507_n_spl_
  );


  buf

  (
    G1884,
    g221_n
  );


  buf

  (
    G1885,
    g224_n
  );


  buf

  (
    G1886,
    g227_n
  );


  buf

  (
    G1887,
    g230_n
  );


  buf

  (
    G1888,
    g234_n
  );


  buf

  (
    G1889,
    g237_n
  );


  buf

  (
    G1890,
    g240_n
  );


  buf

  (
    G1891,
    g246_n
  );


  buf

  (
    G1892,
    g249_n
  );


  buf

  (
    G1893,
    g252_n
  );


  buf

  (
    G1894,
    g255_n
  );


  buf

  (
    G1895,
    g259_n
  );


  buf

  (
    G1896,
    g266_n
  );


  buf

  (
    G1897,
    g269_n
  );


  buf

  (
    G1898,
    g272_n
  );


  buf

  (
    G1899,
    g275_n
  );


  buf

  (
    G1900,
    g283_n
  );


  buf

  (
    G1901,
    g289_p
  );


  buf

  (
    G1902,
    g295_p
  );


  buf

  (
    G1903,
    g299_p
  );


  buf

  (
    G1904,
    g303_p
  );


  buf

  (
    G1905,
    g307_p
  );


  buf

  (
    G1906,
    g316_n
  );


  buf

  (
    G1907,
    g326_n
  );


  buf

  (
    G1908,
    g330_p
  );


  buf

  (
    n2248_li000_li000,
    G1_p
  );


  buf

  (
    n2257_li003_li003,
    n1273_o2_p
  );


  buf

  (
    n2269_li007_li007,
    n1212_o2_p
  );


  buf

  (
    n2281_li011_li011,
    n1213_o2_p
  );


  buf

  (
    n2284_li012_li012,
    G4_p
  );


  buf

  (
    n2293_li015_li015,
    n1274_o2_p
  );


  buf

  (
    n2296_li016_li016,
    G5_p
  );


  buf

  (
    n2305_li019_li019,
    n1275_o2_p
  );


  buf

  (
    n2317_li023_li023,
    n1214_o2_p
  );


  buf

  (
    n2329_li027_li027,
    n1215_o2_p
  );


  buf

  (
    n2341_li031_li031,
    n1216_o2_p
  );


  buf

  (
    n2353_li035_li035,
    n1217_o2_p
  );


  buf

  (
    n2365_li039_li039,
    n1201_o2_p
  );


  buf

  (
    n2368_li040_li040,
    G11_p
  );


  buf

  (
    n2377_li043_li043,
    n1242_o2_p
  );


  buf

  (
    n2389_li047_li047,
    n1202_o2_p
  );


  buf

  (
    n2401_li051_li051,
    n1203_o2_p
  );


  buf

  (
    n2413_li055_li055,
    n1218_o2_p
  );


  buf

  (
    n2425_li059_li059,
    n1204_o2_p
  );


  buf

  (
    n2428_li060_li060,
    G16_p
  );


  buf

  (
    n2437_li063_li063,
    n1243_o2_p
  );


  buf

  (
    n2440_li064_li064,
    G17_p
  );


  buf

  (
    n2464_li072_li072,
    G19_p
  );


  buf

  (
    n2476_li076_li076,
    G20_p
  );


  buf

  (
    n2488_li080_li080,
    G21_p
  );


  buf

  (
    n2497_li083_li083,
    lo082_buf_o2_p
  );


  buf

  (
    n2500_li084_li084,
    G22_p
  );


  buf

  (
    n2503_li085_li085,
    n1192_lo_p
  );


  buf

  (
    n2509_li087_li087,
    lo086_buf_o2_p
  );


  buf

  (
    n2512_li088_li088,
    G23_p
  );


  buf

  (
    n2536_li096_li096,
    G25_p
  );


  buf

  (
    n2539_li097_li097,
    n1228_lo_p
  );


  buf

  (
    n2542_li098_li098,
    n1231_lo_p
  );


  buf

  (
    n2545_li099_li099,
    n1234_lo_p_spl_
  );


  buf

  (
    n2548_li100_li100,
    G26_p
  );


  buf

  (
    n2551_li101_li101,
    n1240_lo_p
  );


  buf

  (
    n2557_li103_li103,
    lo102_buf_o2_p_spl_
  );


  buf

  (
    n2560_li104_li104,
    G27_p
  );


  buf

  (
    n2563_li105_li105,
    n1252_lo_p
  );


  buf

  (
    n2569_li107_li107,
    lo106_buf_o2_p_spl_
  );


  buf

  (
    n2572_li108_li108,
    G28_p
  );


  buf

  (
    n2575_li109_li109,
    n1264_lo_p
  );


  buf

  (
    n2581_li111_li111,
    lo110_buf_o2_p
  );


  buf

  (
    n2584_li112_li112,
    G29_p
  );


  buf

  (
    n2587_li113_li113,
    n1276_lo_p
  );


  buf

  (
    n2590_li114_li114,
    n1279_lo_p
  );


  buf

  (
    n2593_li115_li115,
    n1282_lo_p_spl_
  );


  buf

  (
    n2596_li116_li116,
    G30_p
  );


  buf

  (
    n2599_li117_li117,
    n1288_lo_p
  );


  buf

  (
    n2602_li118_li118,
    n1291_lo_p
  );


  buf

  (
    n2605_li119_li119,
    n1294_lo_p_spl_
  );


  buf

  (
    n2608_li120_li120,
    G31_p
  );


  buf

  (
    n2611_li121_li121,
    n1300_lo_p
  );


  buf

  (
    n2617_li123_li123,
    lo122_buf_o2_p_spl_1
  );


  buf

  (
    n2620_li124_li124,
    G32_p
  );


  buf

  (
    n2623_li125_li125,
    n1312_lo_p
  );


  buf

  (
    n2626_li126_li126,
    n1315_lo_p
  );


  buf

  (
    n2629_li127_li127,
    n1318_lo_p_spl_
  );


  buf

  (
    n2641_li131_li131,
    n1219_o2_p_spl_1
  );


  buf

  (
    n1225_i2,
    n547_o2_p
  );


  buf

  (
    n1229_i2,
    n617_o2_p
  );


  buf

  (
    n1228_i2,
    n424_inv_p
  );


  buf

  (
    n1259_i2,
    n570_o2_p
  );


  buf

  (
    n1272_i2,
    n460_inv_p
  );


  buf

  (
    n1269_i2,
    n528_o2_p
  );


  buf

  (
    n1307_i2,
    n620_o2_p_spl_
  );


  buf

  (
    n1201_i2,
    lo038_buf_o2_p
  );


  buf

  (
    n1202_i2,
    lo046_buf_o2_p
  );


  buf

  (
    n1203_i2,
    lo050_buf_o2_p_spl_
  );


  buf

  (
    n1204_i2,
    lo058_buf_o2_p
  );


  buf

  (
    n622_i2,
    g331_p_spl_
  );


  buf

  (
    n1205_i2,
    lo070_buf_o2_p
  );


  buf

  (
    n1206_i2,
    lo094_buf_o2_p_spl_
  );


  buf

  (
    n497_i2,
    g332_n_spl_
  );


  buf

  (
    n1212_i2,
    lo006_buf_o2_p_spl_
  );


  buf

  (
    n1213_i2,
    lo010_buf_o2_p
  );


  buf

  (
    n1214_i2,
    lo022_buf_o2_p
  );


  buf

  (
    n1215_i2,
    lo026_buf_o2_p
  );


  buf

  (
    n1216_i2,
    lo030_buf_o2_p_spl_
  );


  buf

  (
    n1217_i2,
    lo034_buf_o2_p_spl_
  );


  buf

  (
    n1218_i2,
    lo054_buf_o2_p_spl_
  );


  buf

  (
    n1219_i2,
    lo130_buf_o2_p_spl_1
  );


  buf

  (
    n1242_i2,
    lo042_buf_o2_p
  );


  buf

  (
    n1243_i2,
    lo062_buf_o2_p
  );


  buf

  (
    n1273_i2,
    lo002_buf_o2_p_spl_
  );


  buf

  (
    n1274_i2,
    lo014_buf_o2_p_spl_1
  );


  buf

  (
    n1275_i2,
    lo018_buf_o2_p
  );


  buf

  (
    n1276_i2,
    lo078_buf_o2_p
  );


  buf

  (
    n1277_i2,
    lo090_buf_o2_p_spl_
  );


  buf

  (
    n1286_i2,
    n513_o2_p
  );


  buf

  (
    n1299_i2,
    lo066_buf_o2_p
  );


  not

  (
    n601_i2,
    g333_n_spl_
  );


  buf

  (
    n625_i2,
    g337_p_spl_
  );


  not

  (
    n463_i2,
    g338_n_spl_
  );


  buf

  (
    lo082_buf_i2,
    lo081_buf_o2_p_spl_
  );


  buf

  (
    n455_i2,
    g339_n_spl_
  );


  buf

  (
    n642_i2,
    g340_n_spl_
  );


  buf

  (
    n459_i2,
    g341_n_spl_
  );


  not

  (
    n501_i2,
    g345_p_spl_
  );


  buf

  (
    n599_i2,
    g356_p_spl_
  );


  buf

  (
    n485_i2,
    g357_n_spl_1
  );


  buf

  (
    lo086_buf_i2,
    n1195_lo_p_spl_
  );


  buf

  (
    lo122_buf_i2,
    n1303_lo_p_spl_1
  );


  not

  (
    n502_i2,
    g358_n_spl_
  );


  buf

  (
    n627_i2,
    g360_p_spl_
  );


  buf

  (
    lo038_buf_i2,
    lo037_buf_o2_p_spl_1
  );


  buf

  (
    lo046_buf_i2,
    lo045_buf_o2_p_spl_1
  );


  buf

  (
    lo050_buf_i2,
    lo049_buf_o2_p_spl_
  );


  buf

  (
    lo058_buf_i2,
    lo057_buf_o2_p_spl_1
  );


  buf

  (
    lo070_buf_i2,
    lo069_buf_o2_p_spl_
  );


  buf

  (
    lo094_buf_i2,
    lo093_buf_o2_p_spl_
  );


  buf

  (
    n462_i2,
    g361_n_spl_
  );


  buf

  (
    lo006_buf_i2,
    lo004_buf_o2_p_spl_
  );


  buf

  (
    lo010_buf_i2,
    lo008_buf_o2_p_spl_1
  );


  buf

  (
    lo022_buf_i2,
    lo020_buf_o2_p_spl_1
  );


  buf

  (
    lo026_buf_i2,
    lo024_buf_o2_p_spl_1
  );


  buf

  (
    lo030_buf_i2,
    lo028_buf_o2_p_spl_1
  );


  buf

  (
    lo034_buf_i2,
    lo032_buf_o2_p_spl_
  );


  buf

  (
    lo054_buf_i2,
    lo052_buf_o2_p_spl_
  );


  buf

  (
    lo130_buf_i2,
    lo128_buf_o2_p_spl_
  );


  buf

  (
    n547_i2,
    g369_n_spl_
  );


  buf

  (
    n568_i2,
    g378_p_spl_
  );


  buf

  (
    n617_i2,
    g387_p_spl_
  );


  buf

  (
    lo042_buf_i2,
    n1060_lo_p_spl_
  );


  buf

  (
    lo062_buf_i2,
    n1120_lo_p_spl_
  );


  buf

  (
    lo110_buf_i2,
    n1267_lo_p
  );


  buf

  (
    n733_i2,
    g388_p
  );


  buf

  (
    n734_i2,
    g389_p
  );


  buf

  (
    n570_i2,
    g390_p_spl_
  );


  buf

  (
    n461_i2,
    g395_p
  );


  buf

  (
    n644_i2,
    g397_p
  );


  buf

  (
    n628_i2,
    g398_p
  );


  buf

  (
    n528_i2,
    g409_n_spl_
  );


  not

  (
    n592_i2,
    g419_n_spl_
  );


  buf

  (
    lo002_buf_i2,
    n940_lo_p_spl_
  );


  buf

  (
    lo014_buf_i2,
    n976_lo_p_spl_
  );


  buf

  (
    lo018_buf_i2,
    n988_lo_p_spl_
  );


  buf

  (
    lo078_buf_i2,
    n1168_lo_p_spl_
  );


  buf

  (
    lo090_buf_i2,
    n1204_lo_p
  );


  buf

  (
    n513_i2,
    g422_p_spl_
  );


  buf

  (
    lo102_buf_i2,
    n1243_lo_p
  );


  buf

  (
    lo106_buf_i2,
    n1255_lo_p
  );


  buf

  (
    n600_i2,
    g423_n
  );


  buf

  (
    n529_i2,
    g424_p
  );


  not

  (
    n593_i2,
    g425_p
  );


  buf

  (
    lo066_buf_i2,
    n1132_lo_p_spl_
  );


  buf

  (
    n549_i2,
    g427_p
  );


  not

  (
    n550_i2,
    g428_n
  );


  buf

  (
    n571_i2,
    g430_n
  );


  buf

  (
    n572_i2,
    g431_p
  );


  buf

  (
    n495_i2,
    g442_p
  );


  not

  (
    n496_i2,
    g443_n
  );


  buf

  (
    n620_i2,
    g453_n
  );


  not

  (
    n482_i2,
    g459_n_spl_
  );


  buf

  (
    lo081_buf_i2,
    n1180_lo_p
  );


  buf

  (
    n576_i2,
    g460_p
  );


  buf

  (
    n520_i2,
    g461_p
  );


  buf

  (
    n521_i2,
    g462_p
  );


  buf

  (
    n562_i2,
    g464_p
  );


  buf

  (
    n508_i2,
    g470_p
  );


  not

  (
    n509_i2,
    g471_n
  );


  buf

  (
    lo074_buf_i2,
    n1156_lo_p
  );


  buf

  (
    n539_i2,
    g474_n
  );


  buf

  (
    n536_i2,
    g480_n
  );


  buf

  (
    n516_i2,
    g483_n
  );


  buf

  (
    n491_i2,
    g489_n
  );


  buf

  (
    n557_i2,
    g495_n
  );


  buf

  (
    n586_i2,
    g501_n
  );


  buf

  (
    n483_i2,
    g508_p
  );


  not

  (
    n484_i2,
    g509_n
  );


  buf

  (
    lo004_buf_i2,
    G2_p
  );


  buf

  (
    lo008_buf_i2,
    G3_p
  );


  buf

  (
    lo020_buf_i2,
    G6_p
  );


  buf

  (
    lo024_buf_i2,
    G7_p
  );


  buf

  (
    lo028_buf_i2,
    G8_p
  );


  buf

  (
    lo032_buf_i2,
    G9_p
  );


  buf

  (
    lo052_buf_i2,
    G14_p
  );


  buf

  (
    lo128_buf_i2,
    G33_p
  );


  buf

  (
    lo037_buf_i2,
    G10_p
  );


  buf

  (
    lo045_buf_i2,
    G12_p
  );


  buf

  (
    lo049_buf_i2,
    G13_p
  );


  buf

  (
    lo057_buf_i2,
    G15_p
  );


  buf

  (
    lo069_buf_i2,
    G18_p
  );


  buf

  (
    lo093_buf_i2,
    G24_p
  );


  buf

  (
    n461_o2_n_spl_,
    n461_o2_n
  );


  buf

  (
    n628_o2_p_spl_,
    n628_o2_p
  );


  buf

  (
    n461_o2_p_spl_,
    n461_o2_p
  );


  buf

  (
    n628_o2_n_spl_,
    n628_o2_n
  );


  buf

  (
    g218_n_spl_,
    g218_n
  );


  buf

  (
    g218_n_spl_0,
    g218_n_spl_
  );


  buf

  (
    g218_n_spl_00,
    g218_n_spl_0
  );


  buf

  (
    g218_n_spl_01,
    g218_n_spl_0
  );


  buf

  (
    g218_n_spl_1,
    g218_n_spl_
  );


  buf

  (
    g218_n_spl_10,
    g218_n_spl_1
  );


  buf

  (
    g218_p_spl_,
    g218_p
  );


  buf

  (
    g218_p_spl_0,
    g218_p_spl_
  );


  buf

  (
    g218_p_spl_00,
    g218_p_spl_0
  );


  buf

  (
    g218_p_spl_01,
    g218_p_spl_0
  );


  buf

  (
    g218_p_spl_1,
    g218_p_spl_
  );


  buf

  (
    g218_p_spl_10,
    g218_p_spl_1
  );


  buf

  (
    n644_o2_n_spl_,
    n644_o2_n
  );


  buf

  (
    n644_o2_n_spl_0,
    n644_o2_n_spl_
  );


  buf

  (
    n644_o2_p_spl_,
    n644_o2_p
  );


  buf

  (
    n644_o2_p_spl_0,
    n644_o2_p_spl_
  );


  buf

  (
    g231_n_spl_,
    g231_n
  );


  buf

  (
    g231_n_spl_0,
    g231_n_spl_
  );


  buf

  (
    g231_n_spl_00,
    g231_n_spl_0
  );


  buf

  (
    g231_n_spl_01,
    g231_n_spl_0
  );


  buf

  (
    g231_n_spl_1,
    g231_n_spl_
  );


  buf

  (
    g231_p_spl_,
    g231_p
  );


  buf

  (
    g231_p_spl_0,
    g231_p_spl_
  );


  buf

  (
    g231_p_spl_00,
    g231_p_spl_0
  );


  buf

  (
    g231_p_spl_01,
    g231_p_spl_0
  );


  buf

  (
    g231_p_spl_1,
    g231_p_spl_
  );


  buf

  (
    n501_o2_n_spl_,
    n501_o2_n
  );


  buf

  (
    n463_o2_n_spl_,
    n463_o2_n
  );


  buf

  (
    g242_p_spl_,
    g242_p
  );


  buf

  (
    g242_n_spl_,
    g242_n
  );


  buf

  (
    g243_n_spl_,
    g243_n
  );


  buf

  (
    g243_n_spl_0,
    g243_n_spl_
  );


  buf

  (
    g243_n_spl_1,
    g243_n_spl_
  );


  buf

  (
    g243_p_spl_,
    g243_p
  );


  buf

  (
    g243_p_spl_0,
    g243_p_spl_
  );


  buf

  (
    g243_p_spl_1,
    g243_p_spl_
  );


  buf

  (
    n601_o2_n_spl_,
    n601_o2_n
  );


  buf

  (
    n625_o2_p_spl_,
    n625_o2_p
  );


  buf

  (
    n599_o2_p_spl_,
    n599_o2_p
  );


  buf

  (
    g263_n_spl_,
    g263_n
  );


  buf

  (
    g263_n_spl_0,
    g263_n_spl_
  );


  buf

  (
    g263_n_spl_1,
    g263_n_spl_
  );


  buf

  (
    g263_p_spl_,
    g263_p
  );


  buf

  (
    g263_p_spl_0,
    g263_p_spl_
  );


  buf

  (
    g263_p_spl_1,
    g263_p_spl_
  );


  buf

  (
    g276_n_spl_,
    g276_n
  );


  buf

  (
    g276_n_spl_0,
    g276_n_spl_
  );


  buf

  (
    g276_n_spl_00,
    g276_n_spl_0
  );


  buf

  (
    g276_n_spl_01,
    g276_n_spl_0
  );


  buf

  (
    g276_n_spl_1,
    g276_n_spl_
  );


  buf

  (
    n1333_lo_p_spl_,
    n1333_lo_p
  );


  buf

  (
    n1333_lo_p_spl_0,
    n1333_lo_p_spl_
  );


  buf

  (
    n1309_lo_n_spl_,
    n1309_lo_n
  );


  buf

  (
    n1309_lo_n_spl_0,
    n1309_lo_n_spl_
  );


  buf

  (
    n1309_lo_n_spl_00,
    n1309_lo_n_spl_0
  );


  buf

  (
    n1309_lo_n_spl_1,
    n1309_lo_n_spl_
  );


  buf

  (
    n1309_lo_p_spl_,
    n1309_lo_p
  );


  buf

  (
    n1309_lo_p_spl_0,
    n1309_lo_p_spl_
  );


  buf

  (
    g276_p_spl_,
    g276_p
  );


  buf

  (
    g276_p_spl_0,
    g276_p_spl_
  );


  buf

  (
    n459_o2_p_spl_,
    n459_o2_p
  );


  buf

  (
    n459_o2_p_spl_0,
    n459_o2_p_spl_
  );


  buf

  (
    n459_o2_p_spl_00,
    n459_o2_p_spl_0
  );


  buf

  (
    n459_o2_p_spl_01,
    n459_o2_p_spl_0
  );


  buf

  (
    n459_o2_p_spl_1,
    n459_o2_p_spl_
  );


  buf

  (
    n1333_lo_n_spl_,
    n1333_lo_n
  );


  buf

  (
    g310_n_spl_,
    g310_n
  );


  buf

  (
    g310_p_spl_,
    g310_p
  );


  buf

  (
    g320_n_spl_,
    g320_n
  );


  buf

  (
    g320_p_spl_,
    g320_p
  );


  buf

  (
    n600_o2_n_spl_,
    n600_o2_n
  );


  buf

  (
    lo122_buf_o2_n_spl_,
    lo122_buf_o2_n
  );


  buf

  (
    lo122_buf_o2_p_spl_,
    lo122_buf_o2_p
  );


  buf

  (
    lo122_buf_o2_p_spl_0,
    lo122_buf_o2_p_spl_
  );


  buf

  (
    lo122_buf_o2_p_spl_1,
    lo122_buf_o2_p_spl_
  );


  buf

  (
    n620_o2_p_spl_,
    n620_o2_p
  );


  buf

  (
    g331_p_spl_,
    g331_p
  );


  buf

  (
    n1282_lo_p_spl_,
    n1282_lo_p
  );


  buf

  (
    n1219_o2_p_spl_,
    n1219_o2_p
  );


  buf

  (
    n1219_o2_p_spl_0,
    n1219_o2_p_spl_
  );


  buf

  (
    n1219_o2_p_spl_1,
    n1219_o2_p_spl_
  );


  buf

  (
    n1294_lo_p_spl_,
    n1294_lo_p
  );


  buf

  (
    n1318_lo_p_spl_,
    n1318_lo_p
  );


  buf

  (
    g332_n_spl_,
    g332_n
  );


  buf

  (
    n1234_lo_p_spl_,
    n1234_lo_p
  );


  buf

  (
    lo106_buf_o2_p_spl_,
    lo106_buf_o2_p
  );


  buf

  (
    lo102_buf_o2_p_spl_,
    lo102_buf_o2_p
  );


  buf

  (
    g338_n_spl_,
    g338_n
  );


  buf

  (
    g345_p_spl_,
    g345_p
  );


  buf

  (
    g333_n_spl_,
    g333_n
  );


  buf

  (
    g337_p_spl_,
    g337_p
  );


  buf

  (
    g356_p_spl_,
    g356_p
  );


  buf

  (
    n1303_lo_p_spl_,
    n1303_lo_p
  );


  buf

  (
    n1303_lo_p_spl_0,
    n1303_lo_p_spl_
  );


  buf

  (
    n1303_lo_p_spl_1,
    n1303_lo_p_spl_
  );


  buf

  (
    lo090_buf_o2_p_spl_,
    lo090_buf_o2_p
  );


  buf

  (
    lo090_buf_o2_p_spl_0,
    lo090_buf_o2_p_spl_
  );


  buf

  (
    n539_o2_n_spl_,
    n539_o2_n
  );


  buf

  (
    n536_o2_p_spl_,
    n536_o2_p
  );


  buf

  (
    n539_o2_p_spl_,
    n539_o2_p
  );


  buf

  (
    n536_o2_n_spl_,
    n536_o2_n
  );


  buf

  (
    lo074_buf_o2_p_spl_,
    lo074_buf_o2_p
  );


  buf

  (
    lo130_buf_o2_n_spl_,
    lo130_buf_o2_n
  );


  buf

  (
    lo130_buf_o2_n_spl_0,
    lo130_buf_o2_n_spl_
  );


  buf

  (
    lo130_buf_o2_n_spl_1,
    lo130_buf_o2_n_spl_
  );


  buf

  (
    lo130_buf_o2_p_spl_,
    lo130_buf_o2_p
  );


  buf

  (
    lo130_buf_o2_p_spl_0,
    lo130_buf_o2_p_spl_
  );


  buf

  (
    lo130_buf_o2_p_spl_00,
    lo130_buf_o2_p_spl_0
  );


  buf

  (
    lo130_buf_o2_p_spl_1,
    lo130_buf_o2_p_spl_
  );


  buf

  (
    n516_o2_n_spl_,
    n516_o2_n
  );


  buf

  (
    n516_o2_n_spl_0,
    n516_o2_n_spl_
  );


  buf

  (
    n516_o2_n_spl_1,
    n516_o2_n_spl_
  );


  buf

  (
    n557_o2_p_spl_,
    n557_o2_p
  );


  buf

  (
    n516_o2_p_spl_,
    n516_o2_p
  );


  buf

  (
    n516_o2_p_spl_0,
    n516_o2_p_spl_
  );


  buf

  (
    n516_o2_p_spl_1,
    n516_o2_p_spl_
  );


  buf

  (
    n557_o2_n_spl_,
    n557_o2_n
  );


  buf

  (
    lo050_buf_o2_n_spl_,
    lo050_buf_o2_n
  );


  buf

  (
    n562_o2_p_spl_,
    n562_o2_p
  );


  buf

  (
    lo050_buf_o2_p_spl_,
    lo050_buf_o2_p
  );


  buf

  (
    lo050_buf_o2_p_spl_0,
    lo050_buf_o2_p_spl_
  );


  buf

  (
    n562_o2_n_spl_,
    n562_o2_n
  );


  buf

  (
    n491_o2_p_spl_,
    n491_o2_p
  );


  buf

  (
    n491_o2_p_spl_0,
    n491_o2_p_spl_
  );


  buf

  (
    n586_o2_p_spl_,
    n586_o2_p
  );


  buf

  (
    n586_o2_p_spl_0,
    n586_o2_p_spl_
  );


  buf

  (
    n586_o2_p_spl_1,
    n586_o2_p_spl_
  );


  buf

  (
    n491_o2_n_spl_,
    n491_o2_n
  );


  buf

  (
    n491_o2_n_spl_0,
    n491_o2_n_spl_
  );


  buf

  (
    n586_o2_n_spl_,
    n586_o2_n
  );


  buf

  (
    n586_o2_n_spl_0,
    n586_o2_n_spl_
  );


  buf

  (
    n586_o2_n_spl_1,
    n586_o2_n_spl_
  );


  buf

  (
    lo030_buf_o2_n_spl_,
    lo030_buf_o2_n
  );


  buf

  (
    lo014_buf_o2_p_spl_,
    lo014_buf_o2_p
  );


  buf

  (
    lo014_buf_o2_p_spl_0,
    lo014_buf_o2_p_spl_
  );


  buf

  (
    lo014_buf_o2_p_spl_00,
    lo014_buf_o2_p_spl_0
  );


  buf

  (
    lo014_buf_o2_p_spl_1,
    lo014_buf_o2_p_spl_
  );


  buf

  (
    lo030_buf_o2_p_spl_,
    lo030_buf_o2_p
  );


  buf

  (
    lo030_buf_o2_p_spl_0,
    lo030_buf_o2_p_spl_
  );


  buf

  (
    lo014_buf_o2_n_spl_,
    lo014_buf_o2_n
  );


  buf

  (
    lo014_buf_o2_n_spl_0,
    lo014_buf_o2_n_spl_
  );


  buf

  (
    lo014_buf_o2_n_spl_1,
    lo014_buf_o2_n_spl_
  );


  buf

  (
    g381_n_spl_,
    g381_n
  );


  buf

  (
    g384_p_spl_,
    g384_p
  );


  buf

  (
    g381_p_spl_,
    g381_p
  );


  buf

  (
    g384_n_spl_,
    g384_n
  );


  buf

  (
    g361_n_spl_,
    g361_n
  );


  buf

  (
    g391_p_spl_,
    g391_p
  );


  buf

  (
    g339_n_spl_,
    g339_n
  );


  buf

  (
    g392_n_spl_,
    g392_n
  );


  buf

  (
    g341_n_spl_,
    g341_n
  );


  buf

  (
    g394_n_spl_,
    g394_n
  );


  buf

  (
    g340_n_spl_,
    g340_n
  );


  buf

  (
    g358_n_spl_,
    g358_n
  );


  buf

  (
    g360_p_spl_,
    g360_p
  );


  buf

  (
    g399_p_spl_,
    g399_p
  );


  buf

  (
    g399_n_spl_,
    g399_n
  );


  buf

  (
    lo006_buf_o2_n_spl_,
    lo006_buf_o2_n
  );


  buf

  (
    g403_n_spl_,
    g403_n
  );


  buf

  (
    lo006_buf_o2_p_spl_,
    lo006_buf_o2_p
  );


  buf

  (
    lo006_buf_o2_p_spl_0,
    lo006_buf_o2_p_spl_
  );


  buf

  (
    g403_p_spl_,
    g403_p
  );


  buf

  (
    lo002_buf_o2_p_spl_,
    lo002_buf_o2_p
  );


  buf

  (
    lo002_buf_o2_p_spl_0,
    lo002_buf_o2_p_spl_
  );


  buf

  (
    g410_p_spl_,
    g410_p
  );


  buf

  (
    lo002_buf_o2_n_spl_,
    lo002_buf_o2_n
  );


  buf

  (
    g410_n_spl_,
    g410_n
  );


  buf

  (
    g357_p_spl_,
    g357_p
  );


  buf

  (
    g357_p_spl_0,
    g357_p_spl_
  );


  buf

  (
    g357_n_spl_,
    g357_n
  );


  buf

  (
    g357_n_spl_0,
    g357_n_spl_
  );


  buf

  (
    g357_n_spl_1,
    g357_n_spl_
  );


  buf

  (
    lo032_buf_o2_n_spl_,
    lo032_buf_o2_n
  );


  buf

  (
    lo052_buf_o2_n_spl_,
    lo052_buf_o2_n
  );


  buf

  (
    lo032_buf_o2_p_spl_,
    lo032_buf_o2_p
  );


  buf

  (
    lo032_buf_o2_p_spl_0,
    lo032_buf_o2_p_spl_
  );


  buf

  (
    lo052_buf_o2_p_spl_,
    lo052_buf_o2_p
  );


  buf

  (
    lo052_buf_o2_p_spl_0,
    lo052_buf_o2_p_spl_
  );


  buf

  (
    lo094_buf_o2_p_spl_,
    lo094_buf_o2_p
  );


  buf

  (
    n1303_lo_n_spl_,
    n1303_lo_n
  );


  buf

  (
    n1303_lo_n_spl_0,
    n1303_lo_n_spl_
  );


  buf

  (
    g409_n_spl_,
    g409_n
  );


  buf

  (
    g419_n_spl_,
    g419_n
  );


  buf

  (
    g369_n_spl_,
    g369_n
  );


  buf

  (
    n1267_lo_n_spl_,
    n1267_lo_n
  );


  buf

  (
    g426_p_spl_,
    g426_p
  );


  buf

  (
    g378_p_spl_,
    g378_p
  );


  buf

  (
    g390_p_spl_,
    g390_p
  );


  buf

  (
    g390_p_spl_0,
    g390_p_spl_
  );


  buf

  (
    g429_n_spl_,
    g429_n
  );


  buf

  (
    n1195_lo_p_spl_,
    n1195_lo_p
  );


  buf

  (
    lo054_buf_o2_n_spl_,
    lo054_buf_o2_n
  );


  buf

  (
    lo054_buf_o2_p_spl_,
    lo054_buf_o2_p
  );


  buf

  (
    lo054_buf_o2_p_spl_0,
    lo054_buf_o2_p_spl_
  );


  buf

  (
    g438_n_spl_,
    g438_n
  );


  buf

  (
    g441_p_spl_,
    g441_p
  );


  buf

  (
    lo081_buf_o2_p_spl_,
    lo081_buf_o2_p
  );


  buf

  (
    lo034_buf_o2_p_spl_,
    lo034_buf_o2_p
  );


  buf

  (
    lo034_buf_o2_p_spl_0,
    lo034_buf_o2_p_spl_
  );


  buf

  (
    n482_o2_n_spl_,
    n482_o2_n
  );


  buf

  (
    lo034_buf_o2_n_spl_,
    lo034_buf_o2_n
  );


  buf

  (
    n482_o2_p_spl_,
    n482_o2_p
  );


  buf

  (
    g444_p_spl_,
    g444_p
  );


  buf

  (
    g447_n_spl_,
    g447_n
  );


  buf

  (
    g444_n_spl_,
    g444_n
  );


  buf

  (
    g447_p_spl_,
    g447_p
  );


  buf

  (
    g387_p_spl_,
    g387_p
  );


  buf

  (
    lo037_buf_o2_p_spl_,
    lo037_buf_o2_p
  );


  buf

  (
    lo037_buf_o2_p_spl_0,
    lo037_buf_o2_p_spl_
  );


  buf

  (
    lo037_buf_o2_p_spl_00,
    lo037_buf_o2_p_spl_0
  );


  buf

  (
    lo037_buf_o2_p_spl_1,
    lo037_buf_o2_p_spl_
  );


  buf

  (
    lo057_buf_o2_n_spl_,
    lo057_buf_o2_n
  );


  buf

  (
    lo057_buf_o2_n_spl_0,
    lo057_buf_o2_n_spl_
  );


  buf

  (
    lo037_buf_o2_n_spl_,
    lo037_buf_o2_n
  );


  buf

  (
    lo037_buf_o2_n_spl_0,
    lo037_buf_o2_n_spl_
  );


  buf

  (
    lo037_buf_o2_n_spl_1,
    lo037_buf_o2_n_spl_
  );


  buf

  (
    lo057_buf_o2_p_spl_,
    lo057_buf_o2_p
  );


  buf

  (
    lo057_buf_o2_p_spl_0,
    lo057_buf_o2_p_spl_
  );


  buf

  (
    lo057_buf_o2_p_spl_1,
    lo057_buf_o2_p_spl_
  );


  buf

  (
    n1120_lo_p_spl_,
    n1120_lo_p
  );


  buf

  (
    n1120_lo_p_spl_0,
    n1120_lo_p_spl_
  );


  buf

  (
    g456_n_spl_,
    g456_n
  );


  buf

  (
    n1120_lo_n_spl_,
    n1120_lo_n
  );


  buf

  (
    g456_p_spl_,
    g456_p
  );


  buf

  (
    n1132_lo_p_spl_,
    n1132_lo_p
  );


  buf

  (
    lo093_buf_o2_n_spl_,
    lo093_buf_o2_n
  );


  buf

  (
    n988_lo_p_spl_,
    n988_lo_p
  );


  buf

  (
    n988_lo_p_spl_0,
    n988_lo_p_spl_
  );


  buf

  (
    lo028_buf_o2_n_spl_,
    lo028_buf_o2_n
  );


  buf

  (
    lo028_buf_o2_n_spl_0,
    lo028_buf_o2_n_spl_
  );


  buf

  (
    n988_lo_n_spl_,
    n988_lo_n
  );


  buf

  (
    lo028_buf_o2_p_spl_,
    lo028_buf_o2_p
  );


  buf

  (
    lo028_buf_o2_p_spl_0,
    lo028_buf_o2_p_spl_
  );


  buf

  (
    lo028_buf_o2_p_spl_1,
    lo028_buf_o2_p_spl_
  );


  buf

  (
    n1168_lo_p_spl_,
    n1168_lo_p
  );


  buf

  (
    lo128_buf_o2_n_spl_,
    lo128_buf_o2_n
  );


  buf

  (
    lo069_buf_o2_p_spl_,
    lo069_buf_o2_p
  );


  buf

  (
    lo093_buf_o2_p_spl_,
    lo093_buf_o2_p
  );


  buf

  (
    lo128_buf_o2_p_spl_,
    lo128_buf_o2_p
  );


  buf

  (
    n1060_lo_n_spl_,
    n1060_lo_n
  );


  buf

  (
    n1060_lo_n_spl_0,
    n1060_lo_n_spl_
  );


  buf

  (
    g469_n_spl_,
    g469_n
  );


  buf

  (
    lo045_buf_o2_n_spl_,
    lo045_buf_o2_n
  );


  buf

  (
    lo045_buf_o2_n_spl_0,
    lo045_buf_o2_n_spl_
  );


  buf

  (
    lo045_buf_o2_p_spl_,
    lo045_buf_o2_p
  );


  buf

  (
    lo045_buf_o2_p_spl_0,
    lo045_buf_o2_p_spl_
  );


  buf

  (
    lo045_buf_o2_p_spl_1,
    lo045_buf_o2_p_spl_
  );


  buf

  (
    lo020_buf_o2_p_spl_,
    lo020_buf_o2_p
  );


  buf

  (
    lo020_buf_o2_p_spl_0,
    lo020_buf_o2_p_spl_
  );


  buf

  (
    lo020_buf_o2_p_spl_00,
    lo020_buf_o2_p_spl_0
  );


  buf

  (
    lo020_buf_o2_p_spl_1,
    lo020_buf_o2_p_spl_
  );


  buf

  (
    lo020_buf_o2_n_spl_,
    lo020_buf_o2_n
  );


  buf

  (
    lo020_buf_o2_n_spl_0,
    lo020_buf_o2_n_spl_
  );


  buf

  (
    lo020_buf_o2_n_spl_1,
    lo020_buf_o2_n_spl_
  );


  buf

  (
    lo008_buf_o2_n_spl_,
    lo008_buf_o2_n
  );


  buf

  (
    lo008_buf_o2_n_spl_0,
    lo008_buf_o2_n_spl_
  );


  buf

  (
    lo008_buf_o2_p_spl_,
    lo008_buf_o2_p
  );


  buf

  (
    lo008_buf_o2_p_spl_0,
    lo008_buf_o2_p_spl_
  );


  buf

  (
    lo008_buf_o2_p_spl_1,
    lo008_buf_o2_p_spl_
  );


  buf

  (
    g422_p_spl_,
    g422_p
  );


  buf

  (
    lo004_buf_o2_n_spl_,
    lo004_buf_o2_n
  );


  buf

  (
    lo004_buf_o2_p_spl_,
    lo004_buf_o2_p
  );


  buf

  (
    lo004_buf_o2_p_spl_0,
    lo004_buf_o2_p_spl_
  );


  buf

  (
    n940_lo_p_spl_,
    n940_lo_p
  );


  buf

  (
    lo024_buf_o2_p_spl_,
    lo024_buf_o2_p
  );


  buf

  (
    lo024_buf_o2_p_spl_0,
    lo024_buf_o2_p_spl_
  );


  buf

  (
    lo024_buf_o2_p_spl_00,
    lo024_buf_o2_p_spl_0
  );


  buf

  (
    lo024_buf_o2_p_spl_1,
    lo024_buf_o2_p_spl_
  );


  buf

  (
    lo024_buf_o2_n_spl_,
    lo024_buf_o2_n
  );


  buf

  (
    lo024_buf_o2_n_spl_0,
    lo024_buf_o2_n_spl_
  );


  buf

  (
    lo024_buf_o2_n_spl_1,
    lo024_buf_o2_n_spl_
  );


  buf

  (
    n976_lo_p_spl_,
    n976_lo_p
  );


  buf

  (
    lo049_buf_o2_n_spl_,
    lo049_buf_o2_n
  );


  buf

  (
    lo049_buf_o2_p_spl_,
    lo049_buf_o2_p
  );


  buf

  (
    lo049_buf_o2_p_spl_0,
    lo049_buf_o2_p_spl_
  );


  buf

  (
    n1060_lo_p_spl_,
    n1060_lo_p
  );


  buf

  (
    g459_n_spl_,
    g459_n
  );


  buf

  (
    g459_n_spl_0,
    g459_n_spl_
  );


  buf

  (
    g507_n_spl_,
    g507_n
  );


endmodule
