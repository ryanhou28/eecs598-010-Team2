
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  G42,
  G43,
  G44,
  G45,
  G46,
  G47,
  G48,
  G49,
  G50,
  G3519,
  G3520,
  G3521,
  G3522,
  G3523,
  G3524,
  G3525,
  G3526,
  G3527,
  G3528,
  G3529,
  G3530,
  G3531,
  G3532,
  G3533,
  G3534,
  G3535,
  G3536,
  G3537,
  G3538,
  G3539,
  G3540
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input G42;input G43;input G44;input G45;input G46;input G47;input G48;input G49;input G50;
  output G3519;output G3520;output G3521;output G3522;output G3523;output G3524;output G3525;output G3526;output G3527;output G3528;output G3529;output G3530;output G3531;output G3532;output G3533;output G3534;output G3535;output G3536;output G3537;output G3538;output G3539;output G3540;
  wire new_n73_;wire new_n74_;wire new_n76_;wire new_n78_;wire new_n79_;wire new_n80_;wire new_n81_;wire new_n82_;wire new_n83_;wire new_n84_;wire new_n85_;wire new_n86_;wire new_n87_;wire new_n88_;wire new_n89_;wire new_n90_;wire new_n91_;wire new_n92_;wire new_n93_;wire new_n94_;wire new_n95_;wire new_n96_;wire new_n97_;wire new_n98_;wire new_n99_;wire new_n100_;wire new_n101_;wire new_n102_;wire new_n103_;wire new_n104_;wire new_n105_;wire new_n107_;wire new_n108_;wire new_n109_;wire new_n110_;wire new_n111_;wire new_n112_;wire new_n113_;wire new_n114_;wire new_n115_;wire new_n116_;wire new_n117_;wire new_n118_;wire new_n119_;wire new_n120_;wire new_n121_;wire new_n122_;wire new_n123_;wire new_n124_;wire new_n125_;wire new_n126_;wire new_n128_;wire new_n129_;wire new_n130_;wire new_n131_;wire new_n132_;wire new_n133_;wire new_n134_;wire new_n135_;wire new_n136_;wire new_n137_;wire new_n138_;wire new_n139_;wire new_n140_;wire new_n141_;wire new_n142_;wire new_n143_;wire new_n144_;wire new_n145_;wire new_n146_;wire new_n148_;wire new_n149_;wire new_n150_;wire new_n151_;wire new_n152_;wire new_n153_;wire new_n154_;wire new_n155_;wire new_n156_;wire new_n157_;wire new_n158_;wire new_n159_;wire new_n160_;wire new_n161_;wire new_n162_;wire new_n163_;wire new_n164_;wire new_n165_;wire new_n166_;wire new_n167_;wire new_n168_;wire new_n169_;wire new_n170_;wire new_n171_;wire new_n172_;wire new_n173_;wire new_n174_;wire new_n175_;wire new_n176_;wire new_n177_;wire new_n178_;wire new_n179_;wire new_n180_;wire new_n181_;wire new_n182_;wire new_n183_;wire new_n184_;wire new_n185_;wire new_n186_;wire new_n187_;wire new_n188_;wire new_n189_;wire new_n190_;wire new_n191_;wire new_n192_;wire new_n193_;wire new_n194_;wire new_n195_;wire new_n196_;wire new_n197_;wire new_n198_;wire new_n199_;wire new_n200_;wire new_n201_;wire new_n202_;wire new_n203_;wire new_n204_;wire new_n205_;wire new_n206_;wire new_n207_;wire new_n208_;wire new_n209_;wire new_n210_;wire new_n211_;wire new_n212_;wire new_n213_;wire new_n214_;wire new_n215_;wire new_n216_;wire new_n217_;wire new_n218_;wire new_n219_;wire new_n220_;wire new_n221_;wire new_n222_;wire new_n223_;wire new_n224_;wire new_n225_;wire new_n226_;wire new_n227_;wire new_n228_;wire new_n229_;wire new_n230_;wire new_n231_;wire new_n232_;wire new_n233_;wire new_n234_;wire new_n235_;wire new_n236_;wire new_n237_;wire new_n238_;wire new_n239_;wire new_n240_;wire new_n241_;wire new_n242_;wire new_n243_;wire new_n244_;wire new_n245_;wire new_n246_;wire new_n247_;wire new_n248_;wire new_n249_;wire new_n250_;wire new_n251_;wire new_n252_;wire new_n253_;wire new_n254_;wire new_n255_;wire new_n256_;wire new_n257_;wire new_n258_;wire new_n259_;wire new_n260_;wire new_n261_;wire new_n262_;wire new_n263_;wire new_n264_;wire new_n265_;wire new_n266_;wire new_n267_;wire new_n268_;wire new_n269_;wire new_n270_;wire new_n271_;wire new_n272_;wire new_n273_;wire new_n274_;wire new_n275_;wire new_n276_;wire new_n277_;wire new_n278_;wire new_n279_;wire new_n280_;wire new_n281_;wire new_n282_;wire new_n283_;wire new_n284_;wire new_n285_;wire new_n286_;wire new_n287_;wire new_n288_;wire new_n289_;wire new_n290_;wire new_n291_;wire new_n292_;wire new_n293_;wire new_n294_;wire new_n295_;wire new_n296_;wire new_n297_;wire new_n298_;wire new_n299_;wire new_n300_;wire new_n301_;wire new_n302_;wire new_n303_;wire new_n304_;wire new_n305_;wire new_n306_;wire new_n307_;wire new_n308_;wire new_n309_;wire new_n310_;wire new_n311_;wire new_n312_;wire new_n313_;wire new_n314_;wire new_n315_;wire new_n316_;wire new_n317_;wire new_n318_;wire new_n319_;wire new_n320_;wire new_n321_;wire new_n322_;wire new_n323_;wire new_n324_;wire new_n325_;wire new_n326_;wire new_n327_;wire new_n328_;wire new_n329_;wire new_n330_;wire new_n331_;wire new_n332_;wire new_n333_;wire new_n334_;wire new_n335_;wire new_n336_;wire new_n337_;wire new_n338_;wire new_n339_;wire new_n340_;wire new_n341_;wire new_n342_;wire new_n343_;wire new_n344_;wire new_n345_;wire new_n346_;wire new_n347_;wire new_n348_;wire new_n349_;wire new_n350_;wire new_n351_;wire new_n352_;wire new_n353_;wire new_n354_;wire new_n355_;wire new_n356_;wire new_n357_;wire new_n358_;wire new_n359_;wire new_n360_;wire new_n361_;wire new_n362_;wire new_n363_;wire new_n364_;wire new_n365_;wire new_n366_;wire new_n367_;wire new_n368_;wire new_n369_;wire new_n370_;wire new_n371_;wire new_n372_;wire new_n373_;wire new_n375_;wire new_n376_;wire new_n377_;wire new_n378_;wire new_n379_;wire new_n380_;wire new_n381_;wire new_n382_;wire new_n383_;wire new_n384_;wire new_n385_;wire new_n386_;wire new_n387_;wire new_n389_;wire new_n390_;wire new_n391_;wire new_n392_;wire new_n393_;wire new_n394_;wire new_n395_;wire new_n396_;wire new_n397_;wire new_n398_;wire new_n399_;wire new_n401_;wire new_n402_;wire new_n403_;wire new_n404_;wire new_n406_;wire new_n407_;wire new_n408_;wire new_n409_;wire new_n410_;wire new_n411_;wire new_n412_;wire new_n413_;wire new_n414_;wire new_n415_;wire new_n416_;wire new_n417_;wire new_n418_;wire new_n419_;wire new_n420_;wire new_n421_;wire new_n422_;wire new_n423_;wire new_n424_;wire new_n425_;wire new_n426_;wire new_n427_;wire new_n428_;wire new_n429_;wire new_n430_;wire new_n431_;wire new_n432_;wire new_n433_;wire new_n434_;wire new_n435_;wire new_n436_;wire new_n437_;wire new_n438_;wire new_n439_;wire new_n440_;wire new_n441_;wire new_n442_;wire new_n443_;wire new_n444_;wire new_n445_;wire new_n446_;wire new_n447_;wire new_n448_;wire new_n449_;wire new_n450_;wire new_n451_;wire new_n452_;wire new_n453_;wire new_n454_;wire new_n455_;wire new_n456_;wire new_n457_;wire new_n458_;wire new_n459_;wire new_n460_;wire new_n461_;wire new_n462_;wire new_n463_;wire new_n464_;wire new_n465_;wire new_n466_;wire new_n467_;wire new_n468_;wire new_n469_;wire new_n470_;wire new_n471_;wire new_n472_;wire new_n473_;wire new_n474_;wire new_n476_;wire new_n477_;wire new_n478_;wire new_n479_;wire new_n480_;wire new_n481_;wire new_n482_;wire new_n483_;wire new_n484_;wire new_n485_;wire new_n486_;wire new_n487_;wire new_n488_;wire new_n489_;wire new_n490_;wire new_n491_;wire new_n492_;wire new_n493_;wire new_n494_;wire new_n495_;wire new_n496_;wire new_n497_;wire new_n498_;wire new_n499_;wire new_n500_;wire new_n501_;wire new_n502_;wire new_n503_;wire new_n504_;wire new_n505_;wire new_n506_;wire new_n507_;wire new_n508_;wire new_n509_;wire new_n510_;wire new_n511_;wire new_n512_;wire new_n513_;wire new_n514_;wire new_n515_;wire new_n516_;wire new_n517_;wire new_n518_;wire new_n519_;wire new_n520_;wire new_n521_;wire new_n522_;wire new_n523_;wire new_n524_;wire new_n525_;wire new_n526_;wire new_n527_;wire new_n528_;wire new_n529_;wire new_n530_;wire new_n532_;wire new_n533_;wire new_n534_;wire new_n535_;wire new_n536_;wire new_n537_;wire new_n538_;wire new_n539_;wire new_n540_;wire new_n541_;wire new_n542_;wire new_n543_;wire new_n544_;wire new_n545_;wire new_n546_;wire new_n547_;wire new_n548_;wire new_n549_;wire new_n550_;wire new_n551_;wire new_n552_;wire new_n553_;wire new_n554_;wire new_n555_;wire new_n556_;wire new_n557_;wire new_n558_;wire new_n559_;wire new_n560_;wire new_n561_;wire new_n562_;wire new_n563_;wire new_n564_;wire new_n565_;wire new_n566_;wire new_n567_;wire new_n568_;wire new_n569_;wire new_n570_;wire new_n571_;wire new_n572_;wire new_n574_;wire new_n575_;wire new_n576_;wire new_n577_;wire new_n578_;wire new_n579_;wire new_n580_;wire new_n581_;wire new_n582_;wire new_n583_;wire new_n584_;wire new_n585_;wire new_n586_;wire new_n587_;wire new_n588_;wire new_n589_;wire new_n590_;wire new_n591_;wire new_n592_;wire new_n593_;wire new_n594_;wire new_n595_;wire new_n596_;wire new_n597_;wire new_n598_;wire new_n599_;wire new_n600_;wire new_n601_;wire new_n602_;wire new_n603_;wire new_n604_;wire new_n605_;wire new_n606_;wire new_n607_;wire new_n608_;wire new_n609_;wire new_n610_;wire new_n611_;wire new_n612_;wire new_n613_;wire new_n614_;wire new_n615_;wire new_n616_;wire new_n617_;wire new_n618_;wire new_n619_;wire new_n620_;wire new_n621_;wire new_n622_;wire new_n623_;wire new_n624_;wire new_n625_;wire new_n626_;wire new_n627_;wire new_n628_;wire new_n629_;wire new_n630_;wire new_n631_;wire new_n632_;wire new_n633_;wire new_n634_;wire new_n635_;wire new_n636_;wire new_n637_;wire new_n638_;wire new_n639_;wire new_n640_;wire new_n641_;wire new_n642_;wire new_n644_;wire new_n645_;wire new_n646_;wire new_n647_;wire new_n648_;wire new_n649_;wire new_n650_;wire new_n651_;wire new_n652_;wire new_n653_;wire new_n654_;wire new_n655_;wire new_n656_;wire new_n657_;wire new_n658_;wire new_n659_;wire new_n660_;wire new_n661_;wire new_n662_;wire new_n663_;wire new_n664_;wire new_n665_;wire new_n666_;wire new_n667_;wire new_n668_;wire new_n669_;wire new_n670_;wire new_n671_;wire new_n672_;wire new_n673_;wire new_n674_;wire new_n675_;wire new_n676_;wire new_n677_;wire new_n678_;wire new_n679_;wire new_n680_;wire new_n681_;wire new_n682_;wire new_n683_;wire new_n685_;wire new_n686_;wire new_n687_;wire new_n688_;wire new_n689_;wire new_n690_;wire new_n691_;wire new_n692_;wire new_n693_;wire new_n694_;wire new_n695_;wire new_n696_;wire new_n697_;wire new_n698_;wire new_n699_;wire new_n700_;wire new_n701_;wire new_n702_;wire new_n703_;wire new_n704_;wire new_n705_;wire new_n706_;wire new_n707_;wire new_n708_;wire new_n709_;wire new_n710_;wire new_n711_;wire new_n712_;wire new_n713_;wire new_n714_;wire new_n715_;wire new_n716_;wire new_n717_;wire new_n718_;wire new_n719_;wire new_n720_;wire new_n721_;wire new_n722_;wire new_n723_;wire new_n724_;wire new_n726_;wire new_n727_;wire new_n728_;wire new_n729_;wire new_n730_;wire new_n731_;wire new_n732_;wire new_n733_;wire new_n734_;wire new_n735_;wire new_n736_;wire new_n737_;wire new_n738_;wire new_n739_;wire new_n740_;wire new_n741_;wire new_n742_;wire new_n743_;wire new_n744_;wire new_n745_;wire new_n746_;wire new_n747_;wire new_n748_;wire new_n749_;wire new_n750_;wire new_n751_;wire new_n752_;wire new_n753_;wire new_n754_;wire new_n755_;wire new_n756_;wire new_n757_;wire new_n758_;wire new_n759_;wire new_n760_;wire new_n761_;wire new_n762_;wire new_n763_;wire new_n764_;wire new_n765_;wire new_n766_;wire new_n767_;wire new_n768_;wire new_n769_;wire new_n770_;wire new_n771_;wire new_n772_;wire new_n773_;wire new_n774_;wire new_n775_;wire new_n776_;wire new_n777_;wire new_n778_;wire new_n780_;wire new_n781_;wire new_n782_;wire new_n783_;wire new_n784_;wire new_n785_;wire new_n786_;wire new_n787_;wire new_n788_;wire new_n789_;wire new_n790_;wire new_n791_;wire new_n792_;wire new_n793_;wire new_n794_;wire new_n795_;wire new_n796_;wire new_n797_;wire new_n798_;wire new_n799_;wire new_n800_;wire new_n801_;wire new_n802_;wire new_n803_;wire new_n804_;wire new_n805_;wire new_n806_;wire new_n807_;wire new_n808_;wire new_n809_;wire new_n810_;wire new_n811_;wire new_n812_;wire new_n813_;wire new_n814_;wire new_n815_;wire new_n816_;wire new_n817_;wire new_n818_;wire new_n819_;wire new_n820_;wire new_n821_;wire new_n822_;wire new_n823_;wire new_n824_;wire new_n825_;wire new_n827_;wire new_n828_;wire new_n829_;wire new_n830_;wire new_n831_;wire new_n832_;wire new_n833_;wire new_n834_;wire new_n835_;wire new_n836_;wire new_n837_;wire new_n838_;wire new_n839_;wire new_n840_;wire new_n841_;wire new_n842_;wire new_n843_;wire new_n844_;wire new_n845_;wire new_n846_;wire new_n847_;wire new_n848_;wire new_n849_;wire new_n850_;wire new_n851_;wire new_n852_;wire new_n853_;wire new_n854_;wire new_n855_;wire new_n856_;wire new_n857_;wire new_n858_;wire new_n859_;wire new_n860_;wire new_n861_;wire new_n863_;wire new_n864_;wire new_n865_;wire new_n866_;wire new_n867_;wire new_n868_;wire new_n870_;wire new_n871_;wire new_n872_;wire new_n874_;wire new_n875_;wire new_n876_;wire new_n877_;wire new_n878_;wire new_n879_;wire new_n880_;wire new_n881_;wire new_n882_;wire new_n883_;wire new_n884_;wire new_n885_;wire new_n886_;wire new_n887_;wire new_n888_;wire new_n889_;wire new_n890_;wire new_n891_;wire new_n892_;wire new_n893_;wire new_n895_;wire new_n896_;wire new_n897_;wire new_n898_;wire new_n899_;
  wire G7_spl_;
  wire G7_spl_0;
  wire G7_spl_00;
  wire G7_spl_000;
  wire G7_spl_001;
  wire G7_spl_01;
  wire G7_spl_010;
  wire G7_spl_011;
  wire G7_spl_1;
  wire G7_spl_10;
  wire G7_spl_100;
  wire G7_spl_101;
  wire G7_spl_11;
  wire G7_spl_110;
  wire G7_spl_111;
  wire G8_spl_;
  wire G8_spl_0;
  wire G8_spl_00;
  wire G8_spl_000;
  wire G8_spl_001;
  wire G8_spl_01;
  wire G8_spl_010;
  wire G8_spl_011;
  wire G8_spl_1;
  wire G8_spl_10;
  wire G8_spl_100;
  wire G8_spl_101;
  wire G8_spl_11;
  wire new_n73__spl_;
  wire G9_spl_;
  wire G9_spl_0;
  wire G9_spl_00;
  wire G9_spl_000;
  wire G9_spl_001;
  wire G9_spl_01;
  wire G9_spl_010;
  wire G9_spl_011;
  wire G9_spl_1;
  wire G9_spl_10;
  wire G9_spl_100;
  wire G9_spl_101;
  wire G9_spl_11;
  wire G9_spl_110;
  wire new_n74__spl_;
  wire G10_spl_;
  wire G10_spl_0;
  wire G10_spl_00;
  wire G10_spl_000;
  wire G10_spl_001;
  wire G10_spl_01;
  wire G10_spl_010;
  wire G10_spl_011;
  wire G10_spl_1;
  wire G10_spl_10;
  wire G10_spl_100;
  wire G10_spl_101;
  wire G10_spl_11;
  wire G10_spl_110;
  wire G12_spl_;
  wire G12_spl_0;
  wire G12_spl_00;
  wire G12_spl_000;
  wire G12_spl_001;
  wire G12_spl_01;
  wire G12_spl_010;
  wire G12_spl_011;
  wire G12_spl_1;
  wire G12_spl_10;
  wire G12_spl_100;
  wire G12_spl_101;
  wire G12_spl_11;
  wire G13_spl_;
  wire G13_spl_0;
  wire G13_spl_00;
  wire G13_spl_000;
  wire G13_spl_001;
  wire G13_spl_01;
  wire G13_spl_010;
  wire G13_spl_011;
  wire G13_spl_1;
  wire G13_spl_10;
  wire G13_spl_100;
  wire G13_spl_101;
  wire G13_spl_11;
  wire G13_spl_110;
  wire new_n76__spl_;
  wire G11_spl_;
  wire G11_spl_0;
  wire G11_spl_00;
  wire G11_spl_000;
  wire G11_spl_001;
  wire G11_spl_01;
  wire G11_spl_010;
  wire G11_spl_011;
  wire G11_spl_1;
  wire G11_spl_10;
  wire G11_spl_100;
  wire G11_spl_101;
  wire G11_spl_11;
  wire G1_spl_;
  wire G1_spl_0;
  wire G1_spl_00;
  wire G1_spl_000;
  wire G1_spl_001;
  wire G1_spl_01;
  wire G1_spl_010;
  wire G1_spl_1;
  wire G1_spl_10;
  wire G1_spl_11;
  wire G3_spl_;
  wire G3_spl_0;
  wire G3_spl_00;
  wire G3_spl_000;
  wire G3_spl_0000;
  wire G3_spl_0001;
  wire G3_spl_001;
  wire G3_spl_0010;
  wire G3_spl_0011;
  wire G3_spl_01;
  wire G3_spl_010;
  wire G3_spl_0100;
  wire G3_spl_011;
  wire G3_spl_1;
  wire G3_spl_10;
  wire G3_spl_100;
  wire G3_spl_101;
  wire G3_spl_11;
  wire G3_spl_110;
  wire G3_spl_111;
  wire G34_spl_;
  wire G34_spl_0;
  wire G34_spl_00;
  wire G34_spl_01;
  wire G34_spl_1;
  wire G34_spl_10;
  wire G32_spl_;
  wire G32_spl_0;
  wire G32_spl_00;
  wire G32_spl_01;
  wire G32_spl_1;
  wire G30_spl_;
  wire G30_spl_0;
  wire G30_spl_00;
  wire G30_spl_01;
  wire G30_spl_1;
  wire G33_spl_;
  wire G33_spl_0;
  wire G33_spl_00;
  wire G33_spl_01;
  wire G33_spl_1;
  wire G14_spl_;
  wire G14_spl_0;
  wire G14_spl_00;
  wire G14_spl_000;
  wire G14_spl_001;
  wire G14_spl_01;
  wire G14_spl_010;
  wire G14_spl_011;
  wire G14_spl_1;
  wire G14_spl_10;
  wire G14_spl_100;
  wire G14_spl_101;
  wire G14_spl_11;
  wire G14_spl_110;
  wire G14_spl_111;
  wire G37_spl_;
  wire G37_spl_0;
  wire G37_spl_1;
  wire G31_spl_;
  wire G31_spl_0;
  wire G31_spl_00;
  wire G31_spl_01;
  wire G31_spl_1;
  wire G35_spl_;
  wire G35_spl_0;
  wire G35_spl_00;
  wire G35_spl_01;
  wire G35_spl_1;
  wire G35_spl_10;
  wire G36_spl_;
  wire G36_spl_0;
  wire G36_spl_00;
  wire G36_spl_01;
  wire G36_spl_1;
  wire G2_spl_;
  wire G2_spl_0;
  wire G2_spl_00;
  wire G2_spl_1;
  wire new_n95__spl_;
  wire new_n95__spl_0;
  wire new_n97__spl_;
  wire new_n96__spl_;
  wire new_n96__spl_0;
  wire new_n98__spl_;
  wire new_n98__spl_0;
  wire new_n100__spl_;
  wire new_n100__spl_0;
  wire new_n101__spl_;
  wire new_n101__spl_0;
  wire new_n101__spl_1;
  wire new_n109__spl_;
  wire new_n112__spl_;
  wire new_n118__spl_;
  wire new_n121__spl_;
  wire new_n115__spl_;
  wire new_n124__spl_;
  wire new_n128__spl_;
  wire new_n130__spl_;
  wire new_n133__spl_;
  wire new_n138__spl_;
  wire new_n141__spl_;
  wire new_n136__spl_;
  wire new_n144__spl_;
  wire new_n144__spl_0;
  wire G4_spl_;
  wire G4_spl_0;
  wire G4_spl_00;
  wire G4_spl_000;
  wire G4_spl_0000;
  wire G4_spl_00000;
  wire G4_spl_00001;
  wire G4_spl_0001;
  wire G4_spl_00010;
  wire G4_spl_00011;
  wire G4_spl_001;
  wire G4_spl_0010;
  wire G4_spl_00100;
  wire G4_spl_00101;
  wire G4_spl_0011;
  wire G4_spl_00110;
  wire G4_spl_01;
  wire G4_spl_010;
  wire G4_spl_0100;
  wire G4_spl_0101;
  wire G4_spl_011;
  wire G4_spl_0110;
  wire G4_spl_0111;
  wire G4_spl_1;
  wire G4_spl_10;
  wire G4_spl_100;
  wire G4_spl_1000;
  wire G4_spl_1001;
  wire G4_spl_101;
  wire G4_spl_1010;
  wire G4_spl_1011;
  wire G4_spl_11;
  wire G4_spl_110;
  wire G4_spl_1100;
  wire G4_spl_1101;
  wire G4_spl_111;
  wire G4_spl_1110;
  wire G4_spl_1111;
  wire new_n148__spl_;
  wire new_n154__spl_;
  wire new_n154__spl_0;
  wire new_n154__spl_1;
  wire G39_spl_;
  wire G39_spl_0;
  wire G39_spl_00;
  wire G39_spl_000;
  wire G39_spl_01;
  wire G39_spl_1;
  wire G39_spl_10;
  wire G39_spl_11;
  wire new_n153__spl_;
  wire new_n153__spl_0;
  wire new_n153__spl_1;
  wire new_n151__spl_;
  wire new_n151__spl_0;
  wire new_n151__spl_00;
  wire new_n151__spl_000;
  wire new_n151__spl_001;
  wire new_n151__spl_01;
  wire new_n151__spl_1;
  wire new_n151__spl_10;
  wire new_n151__spl_11;
  wire new_n160__spl_;
  wire new_n160__spl_0;
  wire new_n160__spl_00;
  wire new_n160__spl_01;
  wire new_n160__spl_1;
  wire new_n160__spl_10;
  wire new_n160__spl_11;
  wire new_n162__spl_;
  wire new_n165__spl_;
  wire new_n165__spl_0;
  wire new_n164__spl_;
  wire new_n164__spl_0;
  wire new_n164__spl_1;
  wire G5_spl_;
  wire G5_spl_0;
  wire G5_spl_00;
  wire G5_spl_01;
  wire G5_spl_1;
  wire new_n170__spl_;
  wire new_n171__spl_;
  wire new_n171__spl_0;
  wire new_n171__spl_00;
  wire new_n171__spl_000;
  wire new_n171__spl_01;
  wire new_n171__spl_1;
  wire new_n171__spl_10;
  wire new_n171__spl_11;
  wire G6_spl_;
  wire G6_spl_0;
  wire G6_spl_00;
  wire G6_spl_1;
  wire new_n173__spl_;
  wire new_n173__spl_0;
  wire new_n172__spl_;
  wire new_n172__spl_0;
  wire new_n174__spl_;
  wire new_n174__spl_0;
  wire new_n174__spl_1;
  wire G41_spl_;
  wire G41_spl_0;
  wire G41_spl_00;
  wire G41_spl_01;
  wire G41_spl_1;
  wire G41_spl_10;
  wire new_n180__spl_;
  wire new_n180__spl_0;
  wire new_n180__spl_00;
  wire new_n180__spl_01;
  wire new_n180__spl_1;
  wire new_n180__spl_10;
  wire new_n180__spl_11;
  wire new_n175__spl_;
  wire new_n175__spl_0;
  wire G25_spl_;
  wire G26_spl_;
  wire G26_spl_0;
  wire new_n185__spl_;
  wire new_n185__spl_0;
  wire new_n185__spl_1;
  wire new_n186__spl_;
  wire new_n186__spl_0;
  wire new_n186__spl_00;
  wire new_n186__spl_000;
  wire new_n186__spl_01;
  wire new_n186__spl_1;
  wire new_n186__spl_10;
  wire new_n186__spl_11;
  wire new_n169__spl_;
  wire new_n169__spl_0;
  wire G23_spl_;
  wire G24_spl_;
  wire G24_spl_0;
  wire G24_spl_1;
  wire new_n189__spl_;
  wire new_n189__spl_0;
  wire new_n189__spl_00;
  wire new_n189__spl_01;
  wire new_n189__spl_1;
  wire new_n189__spl_10;
  wire new_n189__spl_11;
  wire new_n191__spl_;
  wire new_n191__spl_0;
  wire new_n197__spl_;
  wire G40_spl_;
  wire G40_spl_0;
  wire G40_spl_00;
  wire G40_spl_01;
  wire G40_spl_1;
  wire G40_spl_10;
  wire new_n210__spl_;
  wire new_n210__spl_0;
  wire new_n210__spl_1;
  wire new_n201__spl_;
  wire new_n201__spl_0;
  wire new_n214__spl_;
  wire new_n214__spl_0;
  wire new_n152__spl_;
  wire new_n152__spl_0;
  wire new_n152__spl_1;
  wire new_n236__spl_;
  wire new_n236__spl_0;
  wire new_n236__spl_1;
  wire new_n226__spl_;
  wire new_n226__spl_0;
  wire new_n240__spl_;
  wire new_n155__spl_;
  wire new_n155__spl_0;
  wire new_n155__spl_1;
  wire new_n248__spl_;
  wire new_n262__spl_;
  wire new_n262__spl_0;
  wire new_n262__spl_1;
  wire new_n253__spl_;
  wire new_n253__spl_0;
  wire new_n266__spl_;
  wire new_n266__spl_0;
  wire new_n241__spl_;
  wire new_n241__spl_0;
  wire new_n241__spl_1;
  wire new_n267__spl_;
  wire new_n267__spl_0;
  wire new_n215__spl_;
  wire new_n215__spl_0;
  wire new_n268__spl_;
  wire new_n192__spl_;
  wire new_n192__spl_0;
  wire new_n269__spl_;
  wire new_n277__spl_;
  wire new_n277__spl_0;
  wire new_n277__spl_1;
  wire new_n283__spl_;
  wire new_n283__spl_0;
  wire new_n283__spl_00;
  wire new_n283__spl_1;
  wire new_n284__spl_;
  wire new_n284__spl_0;
  wire new_n284__spl_1;
  wire new_n293__spl_;
  wire new_n281__spl_;
  wire new_n281__spl_0;
  wire new_n297__spl_;
  wire new_n297__spl_0;
  wire new_n315__spl_;
  wire new_n306__spl_;
  wire new_n306__spl_0;
  wire new_n319__spl_;
  wire new_n319__spl_0;
  wire G21_spl_;
  wire G21_spl_0;
  wire G21_spl_00;
  wire G21_spl_01;
  wire G21_spl_1;
  wire G21_spl_10;
  wire G21_spl_11;
  wire G29_spl_;
  wire new_n339__spl_;
  wire new_n330__spl_;
  wire new_n330__spl_0;
  wire new_n343__spl_;
  wire G22_spl_;
  wire G22_spl_0;
  wire G22_spl_00;
  wire G22_spl_01;
  wire G22_spl_1;
  wire G22_spl_10;
  wire G22_spl_11;
  wire new_n351__spl_;
  wire new_n365__spl_;
  wire new_n356__spl_;
  wire new_n356__spl_0;
  wire new_n369__spl_;
  wire new_n369__spl_0;
  wire new_n344__spl_;
  wire new_n344__spl_0;
  wire new_n344__spl_1;
  wire new_n370__spl_;
  wire new_n370__spl_0;
  wire new_n320__spl_;
  wire new_n320__spl_0;
  wire new_n371__spl_;
  wire new_n298__spl_;
  wire new_n298__spl_0;
  wire new_n372__spl_;
  wire new_n270__spl_;
  wire new_n373__spl_;
  wire new_n373__spl_0;
  wire new_n373__spl_1;
  wire new_n380__spl_;
  wire new_n387__spl_;
  wire G27_spl_;
  wire G27_spl_0;
  wire G48_spl_;
  wire new_n389__spl_;
  wire new_n389__spl_0;
  wire new_n389__spl_1;
  wire new_n390__spl_;
  wire new_n390__spl_0;
  wire new_n390__spl_00;
  wire new_n390__spl_000;
  wire new_n390__spl_001;
  wire new_n390__spl_01;
  wire new_n390__spl_010;
  wire new_n390__spl_011;
  wire new_n390__spl_1;
  wire new_n390__spl_10;
  wire new_n390__spl_100;
  wire new_n390__spl_101;
  wire new_n390__spl_11;
  wire new_n391__spl_;
  wire new_n395__spl_;
  wire G47_spl_;
  wire G47_spl_0;
  wire G47_spl_00;
  wire G47_spl_01;
  wire G47_spl_1;
  wire G47_spl_10;
  wire new_n398__spl_;
  wire new_n398__spl_0;
  wire new_n398__spl_1;
  wire new_n394__spl_;
  wire new_n394__spl_0;
  wire new_n394__spl_1;
  wire new_n401__spl_;
  wire new_n401__spl_0;
  wire new_n401__spl_00;
  wire new_n401__spl_01;
  wire new_n401__spl_1;
  wire new_n401__spl_10;
  wire new_n401__spl_11;
  wire new_n403__spl_;
  wire new_n403__spl_0;
  wire new_n403__spl_00;
  wire new_n403__spl_01;
  wire new_n403__spl_1;
  wire new_n403__spl_10;
  wire new_n407__spl_;
  wire new_n409__spl_;
  wire new_n409__spl_0;
  wire new_n409__spl_00;
  wire new_n409__spl_01;
  wire new_n409__spl_1;
  wire new_n409__spl_10;
  wire new_n411__spl_;
  wire new_n411__spl_0;
  wire new_n410__spl_;
  wire new_n410__spl_0;
  wire new_n410__spl_00;
  wire new_n410__spl_000;
  wire new_n410__spl_001;
  wire new_n410__spl_01;
  wire new_n410__spl_1;
  wire new_n410__spl_10;
  wire new_n410__spl_11;
  wire new_n414__spl_;
  wire new_n414__spl_0;
  wire new_n414__spl_1;
  wire new_n418__spl_;
  wire new_n417__spl_;
  wire new_n417__spl_0;
  wire new_n417__spl_00;
  wire new_n417__spl_000;
  wire new_n417__spl_01;
  wire new_n417__spl_1;
  wire new_n417__spl_10;
  wire new_n417__spl_11;
  wire new_n428__spl_;
  wire new_n428__spl_0;
  wire new_n427__spl_;
  wire new_n427__spl_0;
  wire new_n427__spl_1;
  wire new_n429__spl_;
  wire G45_spl_;
  wire new_n430__spl_;
  wire new_n430__spl_0;
  wire new_n430__spl_00;
  wire new_n430__spl_000;
  wire new_n430__spl_0000;
  wire new_n430__spl_001;
  wire new_n430__spl_01;
  wire new_n430__spl_010;
  wire new_n430__spl_011;
  wire new_n430__spl_1;
  wire new_n430__spl_10;
  wire new_n430__spl_100;
  wire new_n430__spl_101;
  wire new_n430__spl_11;
  wire new_n430__spl_110;
  wire new_n430__spl_111;
  wire new_n432__spl_;
  wire new_n433__spl_;
  wire new_n433__spl_0;
  wire new_n433__spl_00;
  wire new_n433__spl_000;
  wire new_n433__spl_0000;
  wire new_n433__spl_0001;
  wire new_n433__spl_001;
  wire new_n433__spl_01;
  wire new_n433__spl_010;
  wire new_n433__spl_011;
  wire new_n433__spl_1;
  wire new_n433__spl_10;
  wire new_n433__spl_100;
  wire new_n433__spl_101;
  wire new_n433__spl_11;
  wire new_n433__spl_110;
  wire new_n433__spl_111;
  wire new_n435__spl_;
  wire new_n435__spl_0;
  wire new_n435__spl_00;
  wire new_n435__spl_000;
  wire new_n435__spl_001;
  wire new_n435__spl_01;
  wire new_n435__spl_010;
  wire new_n435__spl_011;
  wire new_n435__spl_1;
  wire new_n435__spl_10;
  wire new_n435__spl_100;
  wire new_n435__spl_101;
  wire new_n435__spl_11;
  wire new_n435__spl_110;
  wire new_n435__spl_111;
  wire G44_spl_;
  wire G44_spl_0;
  wire G43_spl_;
  wire G43_spl_0;
  wire G43_spl_1;
  wire new_n437__spl_;
  wire new_n437__spl_0;
  wire new_n437__spl_00;
  wire new_n437__spl_000;
  wire new_n437__spl_0000;
  wire new_n437__spl_001;
  wire new_n437__spl_01;
  wire new_n437__spl_010;
  wire new_n437__spl_011;
  wire new_n437__spl_1;
  wire new_n437__spl_10;
  wire new_n437__spl_100;
  wire new_n437__spl_101;
  wire new_n437__spl_11;
  wire new_n437__spl_110;
  wire new_n437__spl_111;
  wire new_n439__spl_;
  wire new_n439__spl_0;
  wire new_n439__spl_00;
  wire new_n439__spl_000;
  wire new_n439__spl_001;
  wire new_n439__spl_01;
  wire new_n439__spl_010;
  wire new_n439__spl_011;
  wire new_n439__spl_1;
  wire new_n439__spl_10;
  wire new_n439__spl_100;
  wire new_n439__spl_101;
  wire new_n439__spl_11;
  wire G42_spl_;
  wire G42_spl_0;
  wire G42_spl_1;
  wire new_n445__spl_;
  wire new_n445__spl_0;
  wire new_n445__spl_00;
  wire new_n445__spl_000;
  wire new_n445__spl_001;
  wire new_n445__spl_01;
  wire new_n445__spl_010;
  wire new_n445__spl_011;
  wire new_n445__spl_1;
  wire new_n445__spl_10;
  wire new_n445__spl_11;
  wire new_n443__spl_;
  wire new_n458__spl_;
  wire new_n455__spl_;
  wire new_n457__spl_;
  wire new_n456__spl_;
  wire new_n460__spl_;
  wire new_n459__spl_;
  wire new_n477__spl_;
  wire new_n476__spl_;
  wire new_n476__spl_0;
  wire new_n476__spl_1;
  wire new_n480__spl_;
  wire new_n480__spl_0;
  wire new_n480__spl_1;
  wire G18_spl_;
  wire G18_spl_0;
  wire G18_spl_1;
  wire G19_spl_;
  wire G19_spl_0;
  wire G19_spl_1;
  wire G20_spl_;
  wire G20_spl_0;
  wire G20_spl_00;
  wire G20_spl_1;
  wire new_n522__spl_;
  wire new_n522__spl_0;
  wire new_n525__spl_;
  wire new_n523__spl_;
  wire new_n526__spl_;
  wire new_n532__spl_;
  wire new_n536__spl_;
  wire new_n535__spl_;
  wire new_n535__spl_0;
  wire new_n535__spl_00;
  wire new_n535__spl_1;
  wire new_n539__spl_;
  wire new_n539__spl_0;
  wire new_n539__spl_00;
  wire new_n539__spl_1;
  wire new_n540__spl_;
  wire new_n541__spl_;
  wire new_n542__spl_;
  wire new_n543__spl_;
  wire new_n543__spl_0;
  wire new_n550__spl_;
  wire new_n550__spl_0;
  wire new_n552__spl_;
  wire new_n549__spl_;
  wire new_n549__spl_0;
  wire new_n556__spl_;
  wire new_n556__spl_0;
  wire new_n556__spl_1;
  wire new_n547__spl_;
  wire new_n559__spl_;
  wire new_n574__spl_;
  wire new_n577__spl_;
  wire new_n577__spl_0;
  wire new_n583__spl_;
  wire new_n594__spl_;
  wire new_n603__spl_;
  wire new_n611__spl_;
  wire G3526_spl_;
  wire new_n614__spl_;
  wire new_n614__spl_0;
  wire new_n614__spl_00;
  wire new_n614__spl_1;
  wire new_n617__spl_;
  wire new_n618__spl_;
  wire new_n620__spl_;
  wire new_n622__spl_;
  wire new_n615__spl_;
  wire new_n625__spl_;
  wire new_n630__spl_;
  wire new_n634__spl_;
  wire new_n633__spl_;
  wire new_n633__spl_0;
  wire new_n633__spl_1;
  wire new_n637__spl_;
  wire new_n637__spl_0;
  wire new_n637__spl_1;
  wire new_n663__spl_;
  wire new_n664__spl_;
  wire new_n662__spl_;
  wire new_n680__spl_;
  wire new_n680__spl_0;
  wire new_n701__spl_;
  wire new_n712__spl_;
  wire new_n710__spl_;
  wire new_n726__spl_;
  wire new_n729__spl_;
  wire new_n727__spl_;
  wire new_n727__spl_0;
  wire new_n732__spl_;
  wire new_n733__spl_;
  wire new_n733__spl_0;
  wire new_n736__spl_;
  wire new_n738__spl_;
  wire new_n741__spl_;
  wire new_n741__spl_0;
  wire new_n741__spl_1;
  wire new_n743__spl_;
  wire new_n743__spl_0;
  wire new_n735__spl_;
  wire new_n735__spl_0;
  wire new_n735__spl_1;
  wire new_n744__spl_;
  wire new_n744__spl_0;
  wire G16_spl_;
  wire G17_spl_;
  wire G17_spl_0;
  wire new_n777__spl_;
  wire new_n748__spl_;
  wire new_n780__spl_;
  wire new_n783__spl_;
  wire new_n783__spl_0;
  wire new_n817__spl_;
  wire new_n778__spl_;
  wire G3535_spl_;
  wire G3529_spl_;
  wire G3536_spl_;
  wire G3531_spl_;
  wire G3533_spl_;
  wire G3528_spl_;
  wire G3532_spl_;
  wire new_n865__spl_;
  wire new_n866__spl_;
  wire new_n864__spl_;
  wire new_n863__spl_;
  wire new_n863__spl_0;
  wire new_n870__spl_;
  wire new_n875__spl_;
  wire new_n877__spl_;
  wire G50_spl_;
  wire new_n884__spl_;
  wire new_n884__spl_0;
  wire new_n884__spl_1;
  wire new_n882__spl_;
  wire new_n882__spl_0;
  wire new_n882__spl_1;
  wire new_n888__spl_;
  wire new_n880__spl_;
  wire new_n880__spl_0;
  wire new_n880__spl_1;
  wire new_n891__spl_;
  wire new_n897__spl_;

  nor1
  g000
  (
    .dina(G7_spl_000),
    .dinb(G8_spl_000),
    .dout(new_n73_)
  );


  anb1
  g001
  (
    .dina(new_n73__spl_),
    .dinb(G9_spl_000),
    .dout(new_n74_)
  );


  anb1
  g002
  (
    .dina(new_n74__spl_),
    .dinb(G10_spl_000),
    .dout(G3519)
  );


  nor1
  g003
  (
    .dina(G12_spl_000),
    .dinb(G13_spl_000),
    .dout(new_n76_)
  );


  anb2
  g004
  (
    .dina(new_n76__spl_),
    .dinb(G11_spl_000),
    .dout(G3520)
  );


  nor1
  g005
  (
    .dina(G1_spl_000),
    .dinb(G3_spl_0000),
    .dout(new_n78_)
  );


  anb1
  g006
  (
    .dina(G34_spl_00),
    .dinb(G11_spl_000),
    .dout(new_n79_)
  );


  anb2
  g007
  (
    .dina(G9_spl_000),
    .dinb(G32_spl_00),
    .dout(new_n80_)
  );


  anb2
  g008
  (
    .dina(new_n79_),
    .dinb(new_n80_),
    .dout(new_n81_)
  );


  anb2
  g009
  (
    .dina(G7_spl_000),
    .dinb(G30_spl_00),
    .dout(new_n82_)
  );


  anb1
  g010
  (
    .dina(G33_spl_00),
    .dinb(G10_spl_000),
    .dout(new_n83_)
  );


  anb1
  g011
  (
    .dina(new_n82_),
    .dinb(new_n83_),
    .dout(new_n84_)
  );


  anb2
  g012
  (
    .dina(new_n81_),
    .dinb(new_n84_),
    .dout(new_n85_)
  );


  anb2
  g013
  (
    .dina(G14_spl_000),
    .dinb(G37_spl_0),
    .dout(new_n86_)
  );


  anb1
  g014
  (
    .dina(G31_spl_00),
    .dinb(G8_spl_000),
    .dout(new_n87_)
  );


  anb1
  g015
  (
    .dina(new_n86_),
    .dinb(new_n87_),
    .dout(new_n88_)
  );


  anb1
  g016
  (
    .dina(G35_spl_00),
    .dinb(G12_spl_000),
    .dout(new_n89_)
  );


  anb2
  g017
  (
    .dina(G13_spl_000),
    .dinb(G36_spl_00),
    .dout(new_n90_)
  );


  anb2
  g018
  (
    .dina(new_n89_),
    .dinb(new_n90_),
    .dout(new_n91_)
  );


  anb1
  g019
  (
    .dina(new_n88_),
    .dinb(new_n91_),
    .dout(new_n92_)
  );


  anb2
  g020
  (
    .dina(new_n85_),
    .dinb(new_n92_),
    .dout(new_n93_)
  );


  anb2
  g021
  (
    .dina(new_n78_),
    .dinb(new_n93_),
    .dout(new_n94_)
  );


  anb2
  g022
  (
    .dina(G1_spl_000),
    .dinb(G2_spl_00),
    .dout(new_n95_)
  );


  nor1
  g023
  (
    .dina(G3_spl_0000),
    .dinb(new_n95__spl_0),
    .dout(new_n96_)
  );


  and2
  g024
  (
    .dina(G8_spl_001),
    .dinb(G9_spl_001),
    .dout(new_n97_)
  );


  nab1
  g025
  (
    .dina(G7_spl_001),
    .dinb(new_n97__spl_),
    .dout(new_n98_)
  );


  and1
  g026
  (
    .dina(new_n96__spl_0),
    .dinb(new_n98__spl_0),
    .dout(new_n99_)
  );


  and2
  g027
  (
    .dina(G1_spl_001),
    .dinb(G2_spl_00),
    .dout(new_n100_)
  );


  and2
  g028
  (
    .dina(G3_spl_0001),
    .dinb(new_n100__spl_0),
    .dout(new_n101_)
  );


  nor1
  g029
  (
    .dina(G35_spl_00),
    .dinb(G36_spl_00),
    .dout(new_n102_)
  );


  anb1
  g030
  (
    .dina(G34_spl_00),
    .dinb(new_n102_),
    .dout(new_n103_)
  );


  anb2
  g031
  (
    .dina(new_n101__spl_0),
    .dinb(new_n103_),
    .dout(new_n104_)
  );


  anb2
  g032
  (
    .dina(new_n99_),
    .dinb(new_n104_),
    .dout(new_n105_)
  );


  anb1
  g033
  (
    .dina(new_n94_),
    .dinb(new_n105_),
    .dout(G3521)
  );


  anb2
  g034
  (
    .dina(G37_spl_0),
    .dinb(G36_spl_01),
    .dout(new_n107_)
  );


  anb1
  g035
  (
    .dina(G37_spl_1),
    .dinb(G36_spl_01),
    .dout(new_n108_)
  );


  anb1
  g036
  (
    .dina(new_n107_),
    .dinb(new_n108_),
    .dout(new_n109_)
  );


  anb2
  g037
  (
    .dina(G35_spl_01),
    .dinb(G34_spl_01),
    .dout(new_n110_)
  );


  anb1
  g038
  (
    .dina(G35_spl_01),
    .dinb(G34_spl_01),
    .dout(new_n111_)
  );


  anb1
  g039
  (
    .dina(new_n110_),
    .dinb(new_n111_),
    .dout(new_n112_)
  );


  anb2
  g040
  (
    .dina(new_n109__spl_),
    .dinb(new_n112__spl_),
    .dout(new_n113_)
  );


  anb1
  g041
  (
    .dina(new_n109__spl_),
    .dinb(new_n112__spl_),
    .dout(new_n114_)
  );


  anb1
  g042
  (
    .dina(new_n113_),
    .dinb(new_n114_),
    .dout(new_n115_)
  );


  anb2
  g043
  (
    .dina(G33_spl_00),
    .dinb(G32_spl_00),
    .dout(new_n116_)
  );


  anb1
  g044
  (
    .dina(G33_spl_01),
    .dinb(G32_spl_01),
    .dout(new_n117_)
  );


  anb1
  g045
  (
    .dina(new_n116_),
    .dinb(new_n117_),
    .dout(new_n118_)
  );


  anb2
  g046
  (
    .dina(G31_spl_00),
    .dinb(G30_spl_00),
    .dout(new_n119_)
  );


  anb1
  g047
  (
    .dina(G31_spl_01),
    .dinb(G30_spl_01),
    .dout(new_n120_)
  );


  anb1
  g048
  (
    .dina(new_n119_),
    .dinb(new_n120_),
    .dout(new_n121_)
  );


  anb1
  g049
  (
    .dina(new_n118__spl_),
    .dinb(new_n121__spl_),
    .dout(new_n122_)
  );


  anb2
  g050
  (
    .dina(new_n118__spl_),
    .dinb(new_n121__spl_),
    .dout(new_n123_)
  );


  anb2
  g051
  (
    .dina(new_n122_),
    .dinb(new_n123_),
    .dout(new_n124_)
  );


  anb2
  g052
  (
    .dina(new_n115__spl_),
    .dinb(new_n124__spl_),
    .dout(new_n125_)
  );


  anb1
  g053
  (
    .dina(new_n115__spl_),
    .dinb(new_n124__spl_),
    .dout(new_n126_)
  );


  anb1
  g054
  (
    .dina(new_n125_),
    .dinb(new_n126_),
    .dout(G3522)
  );


  and2
  g055
  (
    .dina(G11_spl_001),
    .dinb(G12_spl_001),
    .dout(new_n128_)
  );


  and1
  g056
  (
    .dina(G11_spl_001),
    .dinb(G12_spl_001),
    .dout(new_n129_)
  );


  anb1
  g057
  (
    .dina(new_n128__spl_),
    .dinb(new_n129_),
    .dout(new_n130_)
  );


  anb1
  g058
  (
    .dina(G13_spl_001),
    .dinb(G14_spl_000),
    .dout(new_n131_)
  );


  anb2
  g059
  (
    .dina(G13_spl_001),
    .dinb(G14_spl_001),
    .dout(new_n132_)
  );


  anb2
  g060
  (
    .dina(new_n131_),
    .dinb(new_n132_),
    .dout(new_n133_)
  );


  anb1
  g061
  (
    .dina(new_n130__spl_),
    .dinb(new_n133__spl_),
    .dout(new_n134_)
  );


  anb2
  g062
  (
    .dina(new_n130__spl_),
    .dinb(new_n133__spl_),
    .dout(new_n135_)
  );


  anb2
  g063
  (
    .dina(new_n134_),
    .dinb(new_n135_),
    .dout(new_n136_)
  );


  nor2
  g064
  (
    .dina(G7_spl_001),
    .dinb(G8_spl_001),
    .dout(new_n137_)
  );


  anb2
  g065
  (
    .dina(new_n73__spl_),
    .dinb(new_n137_),
    .dout(new_n138_)
  );


  nor1
  g066
  (
    .dina(G9_spl_001),
    .dinb(G10_spl_001),
    .dout(new_n139_)
  );


  nor2
  g067
  (
    .dina(G9_spl_010),
    .dinb(G10_spl_001),
    .dout(new_n140_)
  );


  anb2
  g068
  (
    .dina(new_n139_),
    .dinb(new_n140_),
    .dout(new_n141_)
  );


  anb2
  g069
  (
    .dina(new_n138__spl_),
    .dinb(new_n141__spl_),
    .dout(new_n142_)
  );


  anb1
  g070
  (
    .dina(new_n138__spl_),
    .dinb(new_n141__spl_),
    .dout(new_n143_)
  );


  nab2
  g071
  (
    .dina(new_n142_),
    .dinb(new_n143_),
    .dout(new_n144_)
  );


  anb1
  g072
  (
    .dina(new_n136__spl_),
    .dinb(new_n144__spl_0),
    .dout(new_n145_)
  );


  anb2
  g073
  (
    .dina(new_n136__spl_),
    .dinb(new_n144__spl_0),
    .dout(new_n146_)
  );


  anb2
  g074
  (
    .dina(new_n145_),
    .dinb(new_n146_),
    .dout(G3523)
  );


  nor2
  g075
  (
    .dina(G1_spl_001),
    .dinb(G2_spl_0),
    .dout(new_n148_)
  );


  nor2
  g076
  (
    .dina(G1_spl_010),
    .dinb(G3_spl_0001),
    .dout(new_n149_)
  );


  anb1
  g077
  (
    .dina(G4_spl_00000),
    .dinb(new_n149_),
    .dout(new_n150_)
  );


  anb1
  g078
  (
    .dina(new_n148__spl_),
    .dinb(new_n150_),
    .dout(new_n151_)
  );


  anb1
  g079
  (
    .dina(G4_spl_00000),
    .dinb(G3_spl_0010),
    .dout(new_n152_)
  );


  anb2
  g080
  (
    .dina(G3_spl_0010),
    .dinb(G4_spl_00001),
    .dout(new_n153_)
  );


  nor1
  g081
  (
    .dina(G3_spl_0011),
    .dinb(G4_spl_00001),
    .dout(new_n154_)
  );


  and2
  g082
  (
    .dina(G3_spl_0011),
    .dinb(G4_spl_00010),
    .dout(new_n155_)
  );


  anb1
  g083
  (
    .dina(new_n154__spl_0),
    .dinb(G12_spl_010),
    .dout(new_n156_)
  );


  nab2
  g084
  (
    .dina(G39_spl_000),
    .dinb(new_n153__spl_0),
    .dout(new_n157_)
  );


  anb2
  g085
  (
    .dina(new_n156_),
    .dinb(new_n157_),
    .dout(new_n158_)
  );


  nab1
  g086
  (
    .dina(new_n151__spl_000),
    .dinb(new_n158_),
    .dout(new_n159_)
  );


  nab2
  g087
  (
    .dina(G3_spl_0100),
    .dinb(new_n95__spl_0),
    .dout(new_n160_)
  );


  nab1
  g088
  (
    .dina(G14_spl_001),
    .dinb(new_n160__spl_00),
    .dout(new_n161_)
  );


  and1
  g089
  (
    .dina(new_n151__spl_000),
    .dinb(new_n160__spl_00),
    .dout(new_n162_)
  );


  anb1
  g090
  (
    .dina(G4_spl_00010),
    .dinb(G1_spl_010),
    .dout(new_n163_)
  );


  anb1
  g091
  (
    .dina(new_n162__spl_),
    .dinb(new_n163_),
    .dout(new_n164_)
  );


  anb1
  g092
  (
    .dina(G3_spl_0100),
    .dinb(new_n151__spl_001),
    .dout(new_n165_)
  );


  anb1
  g093
  (
    .dina(G14_spl_010),
    .dinb(new_n165__spl_0),
    .dout(new_n166_)
  );


  anb2
  g094
  (
    .dina(new_n164__spl_0),
    .dinb(new_n166_),
    .dout(new_n167_)
  );


  anb2
  g095
  (
    .dina(new_n161_),
    .dinb(new_n167_),
    .dout(new_n168_)
  );


  anb2
  g096
  (
    .dina(new_n159_),
    .dinb(new_n168_),
    .dout(new_n169_)
  );


  and1
  g097
  (
    .dina(G4_spl_00011),
    .dinb(G5_spl_00),
    .dout(new_n170_)
  );


  nor1
  g098
  (
    .dina(new_n148__spl_),
    .dinb(new_n170__spl_),
    .dout(new_n171_)
  );


  anb2
  g099
  (
    .dina(new_n171__spl_000),
    .dinb(G38),
    .dout(new_n172_)
  );


  nor1
  g100
  (
    .dina(G1_spl_01),
    .dinb(G6_spl_00),
    .dout(new_n173_)
  );


  anb1
  g101
  (
    .dina(new_n173__spl_0),
    .dinb(G5_spl_00),
    .dout(new_n174_)
  );


  nab1
  g102
  (
    .dina(new_n172__spl_0),
    .dinb(new_n174__spl_0),
    .dout(new_n175_)
  );


  anb1
  g103
  (
    .dina(G37_spl_1),
    .dinb(new_n174__spl_0),
    .dout(new_n176_)
  );


  nor1
  g104
  (
    .dina(G4_spl_00011),
    .dinb(G41_spl_00),
    .dout(new_n177_)
  );


  anb2
  g105
  (
    .dina(G36_spl_1),
    .dinb(G4_spl_00100),
    .dout(new_n178_)
  );


  anb2
  g106
  (
    .dina(new_n177_),
    .dinb(new_n178_),
    .dout(new_n179_)
  );


  and2
  g107
  (
    .dina(G4_spl_00100),
    .dinb(G49),
    .dout(new_n180_)
  );


  anb1
  g108
  (
    .dina(G35_spl_10),
    .dinb(new_n180__spl_00),
    .dout(new_n181_)
  );


  anb1
  g109
  (
    .dina(new_n179_),
    .dinb(new_n181_),
    .dout(new_n182_)
  );


  anb2
  g110
  (
    .dina(new_n176_),
    .dinb(new_n182_),
    .dout(new_n183_)
  );


  anb2
  g111
  (
    .dina(new_n171__spl_000),
    .dinb(new_n183_),
    .dout(new_n184_)
  );


  anb2
  g112
  (
    .dina(new_n175__spl_0),
    .dinb(new_n184_),
    .dout(new_n185_)
  );


  nor1
  g113
  (
    .dina(G25_spl_),
    .dinb(G26_spl_0),
    .dout(new_n186_)
  );


  and2
  g114
  (
    .dina(new_n185__spl_0),
    .dinb(new_n186__spl_000),
    .dout(new_n187_)
  );


  anb2
  g115
  (
    .dina(new_n169__spl_0),
    .dinb(new_n187_),
    .dout(new_n188_)
  );


  and2
  g116
  (
    .dina(G23_spl_),
    .dinb(G24_spl_0),
    .dout(new_n189_)
  );


  anb2
  g117
  (
    .dina(new_n185__spl_0),
    .dinb(new_n189__spl_00),
    .dout(new_n190_)
  );


  anb2
  g118
  (
    .dina(new_n190_),
    .dinb(new_n169__spl_0),
    .dout(new_n191_)
  );


  and1
  g119
  (
    .dina(new_n188_),
    .dinb(new_n191__spl_0),
    .dout(new_n192_)
  );


  anb1
  g120
  (
    .dina(new_n154__spl_0),
    .dinb(G11_spl_010),
    .dout(new_n193_)
  );


  nab2
  g121
  (
    .dina(G14_spl_010),
    .dinb(new_n153__spl_0),
    .dout(new_n194_)
  );


  anb2
  g122
  (
    .dina(new_n193_),
    .dinb(new_n194_),
    .dout(new_n195_)
  );


  anb2
  g123
  (
    .dina(new_n151__spl_001),
    .dinb(new_n195_),
    .dout(new_n196_)
  );


  nab2
  g124
  (
    .dina(new_n160__spl_01),
    .dinb(new_n165__spl_0),
    .dout(new_n197_)
  );


  and1
  g125
  (
    .dina(G13_spl_010),
    .dinb(new_n164__spl_0),
    .dout(new_n198_)
  );


  nab1
  g126
  (
    .dina(G13_spl_010),
    .dinb(new_n197__spl_),
    .dout(new_n199_)
  );


  anb1
  g127
  (
    .dina(new_n196_),
    .dinb(new_n198_),
    .dout(new_n200_)
  );


  anb2
  g128
  (
    .dina(new_n199_),
    .dinb(new_n200_),
    .dout(new_n201_)
  );


  anb1
  g129
  (
    .dina(G36_spl_1),
    .dinb(new_n174__spl_1),
    .dout(new_n202_)
  );


  nor1
  g130
  (
    .dina(G4_spl_00101),
    .dinb(G40_spl_00),
    .dout(new_n203_)
  );


  anb2
  g131
  (
    .dina(G35_spl_10),
    .dinb(G4_spl_00101),
    .dout(new_n204_)
  );


  anb2
  g132
  (
    .dina(new_n203_),
    .dinb(new_n204_),
    .dout(new_n205_)
  );


  anb1
  g133
  (
    .dina(G34_spl_10),
    .dinb(new_n180__spl_00),
    .dout(new_n206_)
  );


  anb1
  g134
  (
    .dina(new_n205_),
    .dinb(new_n206_),
    .dout(new_n207_)
  );


  anb2
  g135
  (
    .dina(new_n202_),
    .dinb(new_n207_),
    .dout(new_n208_)
  );


  anb2
  g136
  (
    .dina(new_n171__spl_00),
    .dinb(new_n208_),
    .dout(new_n209_)
  );


  nab1
  g137
  (
    .dina(new_n175__spl_0),
    .dinb(new_n209_),
    .dout(new_n210_)
  );


  anb2
  g138
  (
    .dina(new_n186__spl_000),
    .dinb(new_n210__spl_0),
    .dout(new_n211_)
  );


  anb1
  g139
  (
    .dina(new_n211_),
    .dinb(new_n201__spl_0),
    .dout(new_n212_)
  );


  nor2
  g140
  (
    .dina(new_n189__spl_00),
    .dinb(new_n210__spl_0),
    .dout(new_n213_)
  );


  anb2
  g141
  (
    .dina(new_n213_),
    .dinb(new_n201__spl_0),
    .dout(new_n214_)
  );


  anb2
  g142
  (
    .dina(new_n212_),
    .dinb(new_n214__spl_0),
    .dout(new_n215_)
  );


  anb2
  g143
  (
    .dina(new_n164__spl_1),
    .dinb(G11_spl_010),
    .dout(new_n216_)
  );


  nab1
  g144
  (
    .dina(G11_spl_011),
    .dinb(new_n160__spl_01),
    .dout(new_n217_)
  );


  anb1
  g145
  (
    .dina(new_n216_),
    .dinb(new_n217_),
    .dout(new_n218_)
  );


  anb1
  g146
  (
    .dina(new_n154__spl_1),
    .dinb(G9_spl_010),
    .dout(new_n219_)
  );


  anb2
  g147
  (
    .dina(G12_spl_010),
    .dinb(new_n152__spl_0),
    .dout(new_n220_)
  );


  nor1
  g148
  (
    .dina(G13_spl_011),
    .dinb(new_n128__spl_),
    .dout(new_n221_)
  );


  anb1
  g149
  (
    .dina(G3_spl_010),
    .dinb(new_n221_),
    .dout(new_n222_)
  );


  anb1
  g150
  (
    .dina(new_n220_),
    .dinb(new_n222_),
    .dout(new_n223_)
  );


  anb2
  g151
  (
    .dina(new_n219_),
    .dinb(new_n223_),
    .dout(new_n224_)
  );


  anb2
  g152
  (
    .dina(new_n151__spl_01),
    .dinb(new_n224_),
    .dout(new_n225_)
  );


  anb2
  g153
  (
    .dina(new_n218_),
    .dinb(new_n225_),
    .dout(new_n226_)
  );


  anb2
  g154
  (
    .dina(new_n172__spl_0),
    .dinb(new_n173__spl_0),
    .dout(new_n227_)
  );


  anb1
  g155
  (
    .dina(G32_spl_01),
    .dinb(new_n180__spl_01),
    .dout(new_n228_)
  );


  nor2
  g156
  (
    .dina(G4_spl_00110),
    .dinb(G33_spl_01),
    .dout(new_n229_)
  );


  anb1
  g157
  (
    .dina(G14_spl_011),
    .dinb(G4_spl_00110),
    .dout(new_n230_)
  );


  anb1
  g158
  (
    .dina(new_n229_),
    .dinb(new_n230_),
    .dout(new_n231_)
  );


  anb1
  g159
  (
    .dina(G34_spl_10),
    .dinb(new_n173__spl_),
    .dout(new_n232_)
  );


  anb1
  g160
  (
    .dina(new_n231_),
    .dinb(new_n232_),
    .dout(new_n233_)
  );


  anb2
  g161
  (
    .dina(new_n228_),
    .dinb(new_n233_),
    .dout(new_n234_)
  );


  nab1
  g162
  (
    .dina(new_n171__spl_01),
    .dinb(new_n234_),
    .dout(new_n235_)
  );


  anb1
  g163
  (
    .dina(new_n227_),
    .dinb(new_n235_),
    .dout(new_n236_)
  );


  anb2
  g164
  (
    .dina(new_n186__spl_00),
    .dinb(new_n236__spl_0),
    .dout(new_n237_)
  );


  anb2
  g165
  (
    .dina(new_n226__spl_0),
    .dinb(new_n237_),
    .dout(new_n238_)
  );


  nor2
  g166
  (
    .dina(new_n189__spl_01),
    .dinb(new_n236__spl_0),
    .dout(new_n239_)
  );


  anb2
  g167
  (
    .dina(new_n239_),
    .dinb(new_n226__spl_0),
    .dout(new_n240_)
  );


  and1
  g168
  (
    .dina(new_n238_),
    .dinb(new_n240__spl_),
    .dout(new_n241_)
  );


  anb1
  g169
  (
    .dina(G12_spl_011),
    .dinb(new_n164__spl_1),
    .dout(new_n242_)
  );


  anb2
  g170
  (
    .dina(G12_spl_011),
    .dinb(new_n160__spl_10),
    .dout(new_n243_)
  );


  anb2
  g171
  (
    .dina(new_n242_),
    .dinb(new_n243_),
    .dout(new_n244_)
  );


  anb1
  g172
  (
    .dina(G10_spl_010),
    .dinb(new_n155__spl_0),
    .dout(new_n245_)
  );


  nab2
  g173
  (
    .dina(G13_spl_011),
    .dinb(new_n153__spl_1),
    .dout(new_n246_)
  );


  nor2
  g174
  (
    .dina(G12_spl_100),
    .dinb(G13_spl_100),
    .dout(new_n247_)
  );


  anb2
  g175
  (
    .dina(new_n76__spl_),
    .dinb(new_n247_),
    .dout(new_n248_)
  );


  anb1
  g176
  (
    .dina(G3_spl_011),
    .dinb(new_n248__spl_),
    .dout(new_n249_)
  );


  anb1
  g177
  (
    .dina(new_n246_),
    .dinb(new_n249_),
    .dout(new_n250_)
  );


  anb2
  g178
  (
    .dina(new_n245_),
    .dinb(new_n250_),
    .dout(new_n251_)
  );


  nab1
  g179
  (
    .dina(new_n151__spl_01),
    .dinb(new_n251_),
    .dout(new_n252_)
  );


  anb1
  g180
  (
    .dina(new_n244_),
    .dinb(new_n252_),
    .dout(new_n253_)
  );


  anb1
  g181
  (
    .dina(G35_spl_1),
    .dinb(new_n174__spl_1),
    .dout(new_n254_)
  );


  nor1
  g182
  (
    .dina(G4_spl_0011),
    .dinb(G39_spl_000),
    .dout(new_n255_)
  );


  anb2
  g183
  (
    .dina(G34_spl_1),
    .dinb(G4_spl_0100),
    .dout(new_n256_)
  );


  anb2
  g184
  (
    .dina(new_n255_),
    .dinb(new_n256_),
    .dout(new_n257_)
  );


  anb1
  g185
  (
    .dina(G33_spl_1),
    .dinb(new_n180__spl_01),
    .dout(new_n258_)
  );


  anb1
  g186
  (
    .dina(new_n257_),
    .dinb(new_n258_),
    .dout(new_n259_)
  );


  anb2
  g187
  (
    .dina(new_n254_),
    .dinb(new_n259_),
    .dout(new_n260_)
  );


  anb2
  g188
  (
    .dina(new_n171__spl_01),
    .dinb(new_n260_),
    .dout(new_n261_)
  );


  anb2
  g189
  (
    .dina(new_n175__spl_),
    .dinb(new_n261_),
    .dout(new_n262_)
  );


  nor1
  g190
  (
    .dina(new_n186__spl_01),
    .dinb(new_n262__spl_0),
    .dout(new_n263_)
  );


  anb2
  g191
  (
    .dina(new_n263_),
    .dinb(new_n253__spl_0),
    .dout(new_n264_)
  );


  anb1
  g192
  (
    .dina(new_n189__spl_01),
    .dinb(new_n262__spl_0),
    .dout(new_n265_)
  );


  anb2
  g193
  (
    .dina(new_n253__spl_0),
    .dinb(new_n265_),
    .dout(new_n266_)
  );


  and1
  g194
  (
    .dina(new_n264_),
    .dinb(new_n266__spl_0),
    .dout(new_n267_)
  );


  nor2
  g195
  (
    .dina(new_n241__spl_0),
    .dinb(new_n267__spl_0),
    .dout(new_n268_)
  );


  and2
  g196
  (
    .dina(new_n215__spl_0),
    .dinb(new_n268__spl_),
    .dout(new_n269_)
  );


  anb1
  g197
  (
    .dina(new_n192__spl_0),
    .dinb(new_n269__spl_),
    .dout(new_n270_)
  );


  anb1
  g198
  (
    .dina(new_n154__spl_1),
    .dinb(G8_spl_010),
    .dout(new_n271_)
  );


  anb2
  g199
  (
    .dina(G11_spl_011),
    .dinb(new_n152__spl_0),
    .dout(new_n272_)
  );


  anb2
  g200
  (
    .dina(new_n271_),
    .dinb(new_n272_),
    .dout(new_n273_)
  );


  anb2
  g201
  (
    .dina(new_n151__spl_10),
    .dinb(new_n273_),
    .dout(new_n274_)
  );


  anb2
  g202
  (
    .dina(G10_spl_010),
    .dinb(new_n160__spl_10),
    .dout(new_n275_)
  );


  anb1
  g203
  (
    .dina(G3_spl_011),
    .dinb(G1_spl_10),
    .dout(new_n276_)
  );


  anb1
  g204
  (
    .dina(new_n162__spl_),
    .dinb(new_n276_),
    .dout(new_n277_)
  );


  anb1
  g205
  (
    .dina(G10_spl_011),
    .dinb(new_n165__spl_),
    .dout(new_n278_)
  );


  anb1
  g206
  (
    .dina(new_n278_),
    .dinb(new_n277__spl_0),
    .dout(new_n279_)
  );


  anb1
  g207
  (
    .dina(new_n275_),
    .dinb(new_n279_),
    .dout(new_n280_)
  );


  anb1
  g208
  (
    .dina(new_n274_),
    .dinb(new_n280_),
    .dout(new_n281_)
  );


  and2
  g209
  (
    .dina(G5_spl_01),
    .dinb(G6_spl_00),
    .dout(new_n282_)
  );


  nab1
  g210
  (
    .dina(G1_spl_10),
    .dinb(new_n282_),
    .dout(new_n283_)
  );


  anb2
  g211
  (
    .dina(new_n172__spl_),
    .dinb(new_n283__spl_00),
    .dout(new_n284_)
  );


  anb1
  g212
  (
    .dina(G33_spl_1),
    .dinb(new_n283__spl_00),
    .dout(new_n285_)
  );


  nor1
  g213
  (
    .dina(G4_spl_0100),
    .dinb(G13_spl_100),
    .dout(new_n286_)
  );


  anb2
  g214
  (
    .dina(G32_spl_1),
    .dinb(G4_spl_0101),
    .dout(new_n287_)
  );


  anb2
  g215
  (
    .dina(new_n286_),
    .dinb(new_n287_),
    .dout(new_n288_)
  );


  anb1
  g216
  (
    .dina(G31_spl_01),
    .dinb(new_n180__spl_10),
    .dout(new_n289_)
  );


  anb1
  g217
  (
    .dina(new_n288_),
    .dinb(new_n289_),
    .dout(new_n290_)
  );


  anb2
  g218
  (
    .dina(new_n285_),
    .dinb(new_n290_),
    .dout(new_n291_)
  );


  nab1
  g219
  (
    .dina(new_n171__spl_10),
    .dinb(new_n291_),
    .dout(new_n292_)
  );


  anb1
  g220
  (
    .dina(new_n284__spl_0),
    .dinb(new_n292_),
    .dout(new_n293_)
  );


  anb1
  g221
  (
    .dina(new_n293__spl_),
    .dinb(new_n186__spl_01),
    .dout(new_n294_)
  );


  anb1
  g222
  (
    .dina(new_n281__spl_0),
    .dinb(new_n294_),
    .dout(new_n295_)
  );


  nab2
  g223
  (
    .dina(new_n189__spl_10),
    .dinb(new_n281__spl_0),
    .dout(new_n296_)
  );


  nab2
  g224
  (
    .dina(new_n293__spl_),
    .dinb(new_n296_),
    .dout(new_n297_)
  );


  anb2
  g225
  (
    .dina(new_n295_),
    .dinb(new_n297__spl_0),
    .dout(new_n298_)
  );


  anb1
  g226
  (
    .dina(G7_spl_010),
    .dinb(new_n155__spl_0),
    .dout(new_n299_)
  );


  nab2
  g227
  (
    .dina(G10_spl_011),
    .dinb(new_n153__spl_1),
    .dout(new_n300_)
  );


  anb2
  g228
  (
    .dina(new_n299_),
    .dinb(new_n300_),
    .dout(new_n301_)
  );


  anb2
  g229
  (
    .dina(new_n151__spl_10),
    .dinb(new_n301_),
    .dout(new_n302_)
  );


  and1
  g230
  (
    .dina(G9_spl_011),
    .dinb(new_n277__spl_0),
    .dout(new_n303_)
  );


  nab1
  g231
  (
    .dina(G9_spl_011),
    .dinb(new_n197__spl_),
    .dout(new_n304_)
  );


  anb1
  g232
  (
    .dina(new_n302_),
    .dinb(new_n303_),
    .dout(new_n305_)
  );


  anb2
  g233
  (
    .dina(new_n304_),
    .dinb(new_n305_),
    .dout(new_n306_)
  );


  anb1
  g234
  (
    .dina(G32_spl_1),
    .dinb(new_n283__spl_0),
    .dout(new_n307_)
  );


  nor1
  g235
  (
    .dina(G4_spl_0101),
    .dinb(G12_spl_100),
    .dout(new_n308_)
  );


  anb2
  g236
  (
    .dina(G31_spl_1),
    .dinb(G4_spl_0110),
    .dout(new_n309_)
  );


  anb2
  g237
  (
    .dina(new_n308_),
    .dinb(new_n309_),
    .dout(new_n310_)
  );


  anb1
  g238
  (
    .dina(G30_spl_01),
    .dinb(new_n180__spl_10),
    .dout(new_n311_)
  );


  anb1
  g239
  (
    .dina(new_n310_),
    .dinb(new_n311_),
    .dout(new_n312_)
  );


  anb2
  g240
  (
    .dina(new_n307_),
    .dinb(new_n312_),
    .dout(new_n313_)
  );


  nab1
  g241
  (
    .dina(new_n171__spl_10),
    .dinb(new_n313_),
    .dout(new_n314_)
  );


  anb1
  g242
  (
    .dina(new_n284__spl_0),
    .dinb(new_n314_),
    .dout(new_n315_)
  );


  anb2
  g243
  (
    .dina(new_n186__spl_10),
    .dinb(new_n315__spl_),
    .dout(new_n316_)
  );


  anb2
  g244
  (
    .dina(new_n306__spl_0),
    .dinb(new_n316_),
    .dout(new_n317_)
  );


  nor2
  g245
  (
    .dina(new_n189__spl_10),
    .dinb(new_n315__spl_),
    .dout(new_n318_)
  );


  anb1
  g246
  (
    .dina(new_n306__spl_0),
    .dinb(new_n318_),
    .dout(new_n319_)
  );


  anb1
  g247
  (
    .dina(new_n317_),
    .dinb(new_n319__spl_0),
    .dout(new_n320_)
  );


  anb2
  g248
  (
    .dina(new_n277__spl_1),
    .dinb(G7_spl_010),
    .dout(new_n321_)
  );


  nab1
  g249
  (
    .dina(G7_spl_011),
    .dinb(new_n160__spl_11),
    .dout(new_n322_)
  );


  anb1
  g250
  (
    .dina(new_n321_),
    .dinb(new_n322_),
    .dout(new_n323_)
  );


  anb1
  g251
  (
    .dina(G21_spl_00),
    .dinb(new_n155__spl_1),
    .dout(new_n324_)
  );


  anb2
  g252
  (
    .dina(G8_spl_010),
    .dinb(new_n152__spl_1),
    .dout(new_n325_)
  );


  anb1
  g253
  (
    .dina(G3_spl_100),
    .dinb(new_n74__spl_),
    .dout(new_n326_)
  );


  anb1
  g254
  (
    .dina(new_n325_),
    .dinb(new_n326_),
    .dout(new_n327_)
  );


  anb2
  g255
  (
    .dina(new_n324_),
    .dinb(new_n327_),
    .dout(new_n328_)
  );


  anb2
  g256
  (
    .dina(new_n151__spl_11),
    .dinb(new_n328_),
    .dout(new_n329_)
  );


  anb2
  g257
  (
    .dina(new_n323_),
    .dinb(new_n329_),
    .dout(new_n330_)
  );


  anb1
  g258
  (
    .dina(G30_spl_1),
    .dinb(new_n283__spl_1),
    .dout(new_n331_)
  );


  nor1
  g259
  (
    .dina(G4_spl_0110),
    .dinb(G10_spl_100),
    .dout(new_n332_)
  );


  anb2
  g260
  (
    .dina(G29_spl_),
    .dinb(G4_spl_0111),
    .dout(new_n333_)
  );


  anb2
  g261
  (
    .dina(new_n332_),
    .dinb(new_n333_),
    .dout(new_n334_)
  );


  anb1
  g262
  (
    .dina(G28),
    .dinb(new_n180__spl_11),
    .dout(new_n335_)
  );


  anb1
  g263
  (
    .dina(new_n334_),
    .dinb(new_n335_),
    .dout(new_n336_)
  );


  anb2
  g264
  (
    .dina(new_n331_),
    .dinb(new_n336_),
    .dout(new_n337_)
  );


  nab1
  g265
  (
    .dina(new_n171__spl_11),
    .dinb(new_n337_),
    .dout(new_n338_)
  );


  anb1
  g266
  (
    .dina(new_n284__spl_1),
    .dinb(new_n338_),
    .dout(new_n339_)
  );


  anb2
  g267
  (
    .dina(new_n186__spl_10),
    .dinb(new_n339__spl_),
    .dout(new_n340_)
  );


  anb2
  g268
  (
    .dina(new_n330__spl_0),
    .dinb(new_n340_),
    .dout(new_n341_)
  );


  nor2
  g269
  (
    .dina(new_n189__spl_11),
    .dinb(new_n330__spl_0),
    .dout(new_n342_)
  );


  nab2
  g270
  (
    .dina(new_n339__spl_),
    .dinb(new_n342_),
    .dout(new_n343_)
  );


  and1
  g271
  (
    .dina(new_n341_),
    .dinb(new_n343__spl_),
    .dout(new_n344_)
  );


  anb2
  g272
  (
    .dina(new_n277__spl_1),
    .dinb(G8_spl_011),
    .dout(new_n345_)
  );


  nab1
  g273
  (
    .dina(G8_spl_011),
    .dinb(new_n160__spl_11),
    .dout(new_n346_)
  );


  anb1
  g274
  (
    .dina(new_n345_),
    .dinb(new_n346_),
    .dout(new_n347_)
  );


  anb1
  g275
  (
    .dina(G22_spl_00),
    .dinb(new_n155__spl_1),
    .dout(new_n348_)
  );


  anb2
  g276
  (
    .dina(G9_spl_100),
    .dinb(new_n152__spl_1),
    .dout(new_n349_)
  );


  and1
  g277
  (
    .dina(G8_spl_100),
    .dinb(G9_spl_100),
    .dout(new_n350_)
  );


  nab2
  g278
  (
    .dina(new_n97__spl_),
    .dinb(new_n350_),
    .dout(new_n351_)
  );


  anb1
  g279
  (
    .dina(G3_spl_100),
    .dinb(new_n351__spl_),
    .dout(new_n352_)
  );


  anb1
  g280
  (
    .dina(new_n349_),
    .dinb(new_n352_),
    .dout(new_n353_)
  );


  anb2
  g281
  (
    .dina(new_n348_),
    .dinb(new_n353_),
    .dout(new_n354_)
  );


  anb2
  g282
  (
    .dina(new_n151__spl_11),
    .dinb(new_n354_),
    .dout(new_n355_)
  );


  anb2
  g283
  (
    .dina(new_n347_),
    .dinb(new_n355_),
    .dout(new_n356_)
  );


  anb1
  g284
  (
    .dina(G31_spl_1),
    .dinb(new_n283__spl_1),
    .dout(new_n357_)
  );


  nor1
  g285
  (
    .dina(G4_spl_0111),
    .dinb(G11_spl_100),
    .dout(new_n358_)
  );


  anb2
  g286
  (
    .dina(G30_spl_1),
    .dinb(G4_spl_1000),
    .dout(new_n359_)
  );


  anb2
  g287
  (
    .dina(new_n358_),
    .dinb(new_n359_),
    .dout(new_n360_)
  );


  anb1
  g288
  (
    .dina(G29_spl_),
    .dinb(new_n180__spl_11),
    .dout(new_n361_)
  );


  anb1
  g289
  (
    .dina(new_n360_),
    .dinb(new_n361_),
    .dout(new_n362_)
  );


  anb2
  g290
  (
    .dina(new_n357_),
    .dinb(new_n362_),
    .dout(new_n363_)
  );


  nab1
  g291
  (
    .dina(new_n171__spl_11),
    .dinb(new_n363_),
    .dout(new_n364_)
  );


  anb1
  g292
  (
    .dina(new_n284__spl_1),
    .dinb(new_n364_),
    .dout(new_n365_)
  );


  anb2
  g293
  (
    .dina(new_n186__spl_11),
    .dinb(new_n365__spl_),
    .dout(new_n366_)
  );


  anb1
  g294
  (
    .dina(new_n366_),
    .dinb(new_n356__spl_0),
    .dout(new_n367_)
  );


  nor2
  g295
  (
    .dina(new_n189__spl_11),
    .dinb(new_n365__spl_),
    .dout(new_n368_)
  );


  anb2
  g296
  (
    .dina(new_n368_),
    .dinb(new_n356__spl_0),
    .dout(new_n369_)
  );


  anb2
  g297
  (
    .dina(new_n367_),
    .dinb(new_n369__spl_0),
    .dout(new_n370_)
  );


  nab2
  g298
  (
    .dina(new_n344__spl_0),
    .dinb(new_n370__spl_0),
    .dout(new_n371_)
  );


  anb1
  g299
  (
    .dina(new_n320__spl_0),
    .dinb(new_n371__spl_),
    .dout(new_n372_)
  );


  anb2
  g300
  (
    .dina(new_n298__spl_0),
    .dinb(new_n372__spl_),
    .dout(new_n373_)
  );


  anb1
  g301
  (
    .dina(new_n270__spl_),
    .dinb(new_n373__spl_0),
    .dout(G3524)
  );


  and2
  g302
  (
    .dina(new_n191__spl_0),
    .dinb(new_n269__spl_),
    .dout(new_n375_)
  );


  nor1
  g303
  (
    .dina(new_n214__spl_0),
    .dinb(new_n268__spl_),
    .dout(new_n376_)
  );


  anb1
  g304
  (
    .dina(new_n241__spl_0),
    .dinb(new_n266__spl_0),
    .dout(new_n377_)
  );


  anb1
  g305
  (
    .dina(new_n240__spl_),
    .dinb(new_n377_),
    .dout(new_n378_)
  );


  anb2
  g306
  (
    .dina(new_n376_),
    .dinb(new_n378_),
    .dout(new_n379_)
  );


  anb1
  g307
  (
    .dina(new_n375_),
    .dinb(new_n379_),
    .dout(new_n380_)
  );


  nor1
  g308
  (
    .dina(new_n373__spl_0),
    .dinb(new_n380__spl_),
    .dout(new_n381_)
  );


  anb2
  g309
  (
    .dina(new_n297__spl_0),
    .dinb(new_n372__spl_),
    .dout(new_n382_)
  );


  anb1
  g310
  (
    .dina(new_n319__spl_0),
    .dinb(new_n371__spl_),
    .dout(new_n383_)
  );


  anb1
  g311
  (
    .dina(new_n344__spl_0),
    .dinb(new_n369__spl_0),
    .dout(new_n384_)
  );


  anb1
  g312
  (
    .dina(new_n343__spl_),
    .dinb(new_n384_),
    .dout(new_n385_)
  );


  anb2
  g313
  (
    .dina(new_n383_),
    .dinb(new_n385_),
    .dout(new_n386_)
  );


  anb1
  g314
  (
    .dina(new_n382_),
    .dinb(new_n386_),
    .dout(new_n387_)
  );


  anb2
  g315
  (
    .dina(new_n381_),
    .dinb(new_n387__spl_),
    .dout(G3525)
  );


  nab2
  g316
  (
    .dina(G27_spl_0),
    .dinb(new_n101__spl_0),
    .dout(new_n389_)
  );


  nab2
  g317
  (
    .dina(G48_spl_),
    .dinb(new_n389__spl_0),
    .dout(new_n390_)
  );


  anb1
  g318
  (
    .dina(new_n201__spl_),
    .dinb(new_n390__spl_000),
    .dout(new_n391_)
  );


  anb1
  g319
  (
    .dina(new_n215__spl_0),
    .dinb(new_n391__spl_),
    .dout(new_n392_)
  );


  anb2
  g320
  (
    .dina(new_n215__spl_),
    .dinb(new_n391__spl_),
    .dout(new_n393_)
  );


  anb2
  g321
  (
    .dina(new_n392_),
    .dinb(new_n393_),
    .dout(new_n394_)
  );


  anb2
  g322
  (
    .dina(new_n390__spl_000),
    .dinb(new_n169__spl_),
    .dout(new_n395_)
  );


  anb2
  g323
  (
    .dina(new_n192__spl_0),
    .dinb(new_n395__spl_),
    .dout(new_n396_)
  );


  anb1
  g324
  (
    .dina(new_n192__spl_),
    .dinb(new_n395__spl_),
    .dout(new_n397_)
  );


  anb1
  g325
  (
    .dina(new_n396_),
    .dinb(new_n397_),
    .dout(new_n398_)
  );


  nor2
  g326
  (
    .dina(G47_spl_00),
    .dinb(new_n398__spl_0),
    .dout(new_n399_)
  );


  anb1
  g327
  (
    .dina(new_n394__spl_0),
    .dinb(new_n399_),
    .dout(G3526)
  );


  anb1
  g328
  (
    .dina(G5_spl_01),
    .dinb(new_n101__spl_1),
    .dout(new_n401_)
  );


  anb1
  g329
  (
    .dina(new_n98__spl_0),
    .dinb(new_n401__spl_00),
    .dout(new_n402_)
  );


  nab1
  g330
  (
    .dina(new_n380__spl_),
    .dinb(new_n390__spl_001),
    .dout(new_n403_)
  );


  anb2
  g331
  (
    .dina(G1_spl_11),
    .dinb(new_n403__spl_00),
    .dout(new_n404_)
  );


  anb2
  g332
  (
    .dina(new_n402_),
    .dinb(new_n404_),
    .dout(G3527)
  );


  anb1
  g333
  (
    .dina(new_n398__spl_0),
    .dinb(G47_spl_00),
    .dout(new_n406_)
  );


  and2
  g334
  (
    .dina(G2_spl_1),
    .dinb(G3_spl_101),
    .dout(new_n407_)
  );


  nab2
  g335
  (
    .dina(G6_spl_0),
    .dinb(new_n407__spl_),
    .dout(new_n408_)
  );


  anb2
  g336
  (
    .dina(G1_spl_11),
    .dinb(new_n408_),
    .dout(new_n409_)
  );


  nab2
  g337
  (
    .dina(new_n401__spl_00),
    .dinb(new_n409__spl_00),
    .dout(new_n410_)
  );


  anb2
  g338
  (
    .dina(new_n398__spl_1),
    .dinb(G47_spl_01),
    .dout(new_n411_)
  );


  anb2
  g339
  (
    .dina(new_n406_),
    .dinb(new_n411__spl_0),
    .dout(new_n412_)
  );


  anb1
  g340
  (
    .dina(new_n410__spl_000),
    .dinb(new_n412_),
    .dout(new_n413_)
  );


  nab2
  g341
  (
    .dina(G4_spl_1000),
    .dinb(new_n407__spl_),
    .dout(new_n414_)
  );


  anb1
  g342
  (
    .dina(new_n398__spl_1),
    .dinb(new_n414__spl_0),
    .dout(new_n415_)
  );


  anb2
  g343
  (
    .dina(G23_spl_),
    .dinb(G3_spl_101),
    .dout(new_n416_)
  );


  anb1
  g344
  (
    .dina(new_n416_),
    .dinb(new_n95__spl_),
    .dout(new_n417_)
  );


  nor1
  g345
  (
    .dina(G4_spl_1001),
    .dinb(new_n101__spl_1),
    .dout(new_n418_)
  );


  anb2
  g346
  (
    .dina(new_n418__spl_),
    .dinb(G14_spl_011),
    .dout(new_n419_)
  );


  anb2
  g347
  (
    .dina(G6_spl_1),
    .dinb(new_n144__spl_),
    .dout(new_n420_)
  );


  anb1
  g348
  (
    .dina(G6_spl_1),
    .dinb(new_n98__spl_),
    .dout(new_n421_)
  );


  nab1
  g349
  (
    .dina(G3520),
    .dinb(new_n418__spl_),
    .dout(new_n422_)
  );


  anb2
  g350
  (
    .dina(new_n421_),
    .dinb(new_n422_),
    .dout(new_n423_)
  );


  anb1
  g351
  (
    .dina(new_n420_),
    .dinb(new_n423_),
    .dout(new_n424_)
  );


  anb1
  g352
  (
    .dina(new_n419_),
    .dinb(new_n424_),
    .dout(new_n425_)
  );


  anb1
  g353
  (
    .dina(new_n417__spl_000),
    .dinb(new_n425_),
    .dout(new_n426_)
  );


  nor2
  g354
  (
    .dina(G3_spl_110),
    .dinb(G25_spl_),
    .dout(new_n427_)
  );


  and1
  g355
  (
    .dina(G3_spl_110),
    .dinb(G24_spl_0),
    .dout(new_n428_)
  );


  anb2
  g356
  (
    .dina(new_n428__spl_0),
    .dinb(G26_spl_0),
    .dout(new_n429_)
  );


  anb1
  g357
  (
    .dina(new_n427__spl_0),
    .dinb(new_n429__spl_),
    .dout(new_n430_)
  );


  anb1
  g358
  (
    .dina(G45_spl_),
    .dinb(new_n430__spl_0000),
    .dout(new_n431_)
  );


  and2
  g359
  (
    .dina(G26_spl_),
    .dinb(new_n428__spl_0),
    .dout(new_n432_)
  );


  nor1
  g360
  (
    .dina(new_n427__spl_0),
    .dinb(new_n432__spl_),
    .dout(new_n433_)
  );


  anb2
  g361
  (
    .dina(new_n433__spl_0000),
    .dinb(G46),
    .dout(new_n434_)
  );


  anb1
  g362
  (
    .dina(new_n427__spl_1),
    .dinb(new_n432__spl_),
    .dout(new_n435_)
  );


  anb2
  g363
  (
    .dina(new_n435__spl_000),
    .dinb(G44_spl_0),
    .dout(new_n436_)
  );


  and2
  g364
  (
    .dina(new_n427__spl_1),
    .dinb(new_n429__spl_),
    .dout(new_n437_)
  );


  and1
  g365
  (
    .dina(G43_spl_0),
    .dinb(new_n437__spl_0000),
    .dout(new_n438_)
  );


  nor2
  g366
  (
    .dina(G3_spl_111),
    .dinb(new_n430__spl_0000),
    .dout(new_n439_)
  );


  and1
  g367
  (
    .dina(G41_spl_00),
    .dinb(new_n439__spl_000),
    .dout(new_n440_)
  );


  anb1
  g368
  (
    .dina(G42_spl_0),
    .dinb(new_n433__spl_0000),
    .dout(new_n441_)
  );


  nor2
  g369
  (
    .dina(G39_spl_00),
    .dinb(new_n437__spl_0000),
    .dout(new_n442_)
  );


  anb2
  g370
  (
    .dina(new_n441_),
    .dinb(new_n442_),
    .dout(new_n443_)
  );


  anb2
  g371
  (
    .dina(new_n186__spl_11),
    .dinb(G3_spl_111),
    .dout(new_n444_)
  );


  anb2
  g372
  (
    .dina(new_n428__spl_),
    .dinb(new_n444_),
    .dout(new_n445_)
  );


  nor2
  g373
  (
    .dina(G40_spl_00),
    .dinb(new_n445__spl_000),
    .dout(new_n446_)
  );


  anb2
  g374
  (
    .dina(new_n431_),
    .dinb(new_n436_),
    .dout(new_n447_)
  );


  anb1
  g375
  (
    .dina(new_n434_),
    .dinb(new_n438_),
    .dout(new_n448_)
  );


  nab1
  g376
  (
    .dina(new_n443__spl_),
    .dinb(new_n448_),
    .dout(new_n449_)
  );


  anb2
  g377
  (
    .dina(new_n447_),
    .dinb(new_n449_),
    .dout(new_n450_)
  );


  anb2
  g378
  (
    .dina(new_n440_),
    .dinb(G4_spl_1001),
    .dout(new_n451_)
  );


  anb1
  g379
  (
    .dina(new_n446_),
    .dinb(new_n451_),
    .dout(new_n452_)
  );


  anb2
  g380
  (
    .dina(new_n450_),
    .dinb(new_n452_),
    .dout(new_n453_)
  );


  nor1
  g381
  (
    .dina(G8_spl_100),
    .dinb(new_n435__spl_000),
    .dout(new_n454_)
  );


  nab1
  g382
  (
    .dina(G12_spl_101),
    .dinb(new_n445__spl_000),
    .dout(new_n455_)
  );


  nab1
  g383
  (
    .dina(G13_spl_101),
    .dinb(new_n437__spl_000),
    .dout(new_n456_)
  );


  anb2
  g384
  (
    .dina(new_n433__spl_0001),
    .dinb(G22_spl_00),
    .dout(new_n457_)
  );


  anb2
  g385
  (
    .dina(G9_spl_101),
    .dinb(new_n437__spl_001),
    .dout(new_n458_)
  );


  nab1
  g386
  (
    .dina(G4_spl_1010),
    .dinb(new_n458__spl_),
    .dout(new_n459_)
  );


  nab1
  g387
  (
    .dina(G11_spl_100),
    .dinb(new_n439__spl_000),
    .dout(new_n460_)
  );


  and2
  g388
  (
    .dina(G10_spl_100),
    .dinb(new_n433__spl_0001),
    .dout(new_n461_)
  );


  and2
  g389
  (
    .dina(G7_spl_011),
    .dinb(new_n430__spl_000),
    .dout(new_n462_)
  );


  anb2
  g390
  (
    .dina(new_n454_),
    .dinb(new_n462_),
    .dout(new_n463_)
  );


  anb2
  g391
  (
    .dina(new_n455__spl_),
    .dinb(new_n457__spl_),
    .dout(new_n464_)
  );


  nab1
  g392
  (
    .dina(new_n456__spl_),
    .dinb(new_n461_),
    .dout(new_n465_)
  );


  anb1
  g393
  (
    .dina(new_n465_),
    .dinb(new_n460__spl_),
    .dout(new_n466_)
  );


  anb1
  g394
  (
    .dina(new_n459__spl_),
    .dinb(new_n464_),
    .dout(new_n467_)
  );


  anb2
  g395
  (
    .dina(new_n463_),
    .dinb(new_n467_),
    .dout(new_n468_)
  );


  anb1
  g396
  (
    .dina(new_n466_),
    .dinb(new_n468_),
    .dout(new_n469_)
  );


  anb1
  g397
  (
    .dina(new_n453_),
    .dinb(new_n469_),
    .dout(new_n470_)
  );


  anb2
  g398
  (
    .dina(new_n417__spl_000),
    .dinb(new_n470_),
    .dout(new_n471_)
  );


  anb2
  g399
  (
    .dina(new_n426_),
    .dinb(new_n471_),
    .dout(new_n472_)
  );


  anb1
  g400
  (
    .dina(new_n472_),
    .dinb(new_n410__spl_000),
    .dout(new_n473_)
  );


  anb2
  g401
  (
    .dina(new_n415_),
    .dinb(new_n473_),
    .dout(new_n474_)
  );


  anb2
  g402
  (
    .dina(new_n413_),
    .dinb(new_n474_),
    .dout(G3528)
  );


  anb2
  g403
  (
    .dina(G2_spl_1),
    .dinb(G4_spl_1010),
    .dout(new_n476_)
  );


  nor1
  g404
  (
    .dina(new_n281__spl_),
    .dinb(new_n390__spl_001),
    .dout(new_n477_)
  );


  anb1
  g405
  (
    .dina(new_n298__spl_0),
    .dinb(new_n477__spl_),
    .dout(new_n478_)
  );


  anb2
  g406
  (
    .dina(new_n298__spl_),
    .dinb(new_n477__spl_),
    .dout(new_n479_)
  );


  anb2
  g407
  (
    .dina(new_n478_),
    .dinb(new_n479_),
    .dout(new_n480_)
  );


  and2
  g408
  (
    .dina(new_n476__spl_0),
    .dinb(new_n480__spl_0),
    .dout(new_n481_)
  );


  anb2
  g409
  (
    .dina(new_n433__spl_001),
    .dinb(G18_spl_0),
    .dout(new_n482_)
  );


  anb1
  g410
  (
    .dina(G19_spl_0),
    .dinb(new_n430__spl_001),
    .dout(new_n483_)
  );


  anb1
  g411
  (
    .dina(new_n482_),
    .dinb(new_n483_),
    .dout(new_n484_)
  );


  nab1
  g412
  (
    .dina(G8_spl_101),
    .dinb(new_n445__spl_001),
    .dout(new_n485_)
  );


  anb1
  g413
  (
    .dina(G20_spl_00),
    .dinb(new_n435__spl_001),
    .dout(new_n486_)
  );


  nab1
  g414
  (
    .dina(G7_spl_100),
    .dinb(new_n439__spl_001),
    .dout(new_n487_)
  );


  nor2
  g415
  (
    .dina(G21_spl_00),
    .dinb(new_n437__spl_001),
    .dout(new_n488_)
  );


  anb2
  g416
  (
    .dina(new_n486_),
    .dinb(new_n488_),
    .dout(new_n489_)
  );


  anb1
  g417
  (
    .dina(new_n484_),
    .dinb(new_n489_),
    .dout(new_n490_)
  );


  anb1
  g418
  (
    .dina(new_n457__spl_),
    .dinb(new_n485_),
    .dout(new_n491_)
  );


  and1
  g419
  (
    .dina(new_n459__spl_),
    .dinb(new_n491_),
    .dout(new_n492_)
  );


  anb2
  g420
  (
    .dina(new_n487_),
    .dinb(new_n492_),
    .dout(new_n493_)
  );


  anb1
  g421
  (
    .dina(new_n490_),
    .dinb(new_n493_),
    .dout(new_n494_)
  );


  nor1
  g422
  (
    .dina(G14_spl_100),
    .dinb(new_n433__spl_001),
    .dout(new_n495_)
  );


  anb2
  g423
  (
    .dina(new_n430__spl_001),
    .dinb(G41_spl_01),
    .dout(new_n496_)
  );


  anb2
  g424
  (
    .dina(new_n495_),
    .dinb(new_n496_),
    .dout(new_n497_)
  );


  anb2
  g425
  (
    .dina(new_n435__spl_001),
    .dinb(G40_spl_01),
    .dout(new_n498_)
  );


  nab1
  g426
  (
    .dina(G11_spl_101),
    .dinb(new_n437__spl_010),
    .dout(new_n499_)
  );


  anb1
  g427
  (
    .dina(new_n498_),
    .dinb(new_n499_),
    .dout(new_n500_)
  );


  anb2
  g428
  (
    .dina(new_n497_),
    .dinb(new_n500_),
    .dout(new_n501_)
  );


  anb2
  g429
  (
    .dina(G13_spl_101),
    .dinb(new_n439__spl_001),
    .dout(new_n502_)
  );


  anb1
  g430
  (
    .dina(G4_spl_1011),
    .dinb(new_n455__spl_),
    .dout(new_n503_)
  );


  anb2
  g431
  (
    .dina(new_n443__spl_),
    .dinb(new_n503_),
    .dout(new_n504_)
  );


  anb1
  g432
  (
    .dina(new_n502_),
    .dinb(new_n504_),
    .dout(new_n505_)
  );


  anb2
  g433
  (
    .dina(new_n501_),
    .dinb(new_n505_),
    .dout(new_n506_)
  );


  anb2
  g434
  (
    .dina(new_n494_),
    .dinb(new_n506_),
    .dout(new_n507_)
  );


  anb2
  g435
  (
    .dina(new_n417__spl_00),
    .dinb(new_n507_),
    .dout(new_n508_)
  );


  anb2
  g436
  (
    .dina(new_n410__spl_001),
    .dinb(new_n508_),
    .dout(new_n509_)
  );


  anb1
  g437
  (
    .dina(new_n481_),
    .dinb(new_n509_),
    .dout(new_n510_)
  );


  anb1
  g438
  (
    .dina(new_n185__spl_1),
    .dinb(new_n210__spl_1),
    .dout(new_n511_)
  );


  anb2
  g439
  (
    .dina(new_n236__spl_1),
    .dinb(new_n262__spl_1),
    .dout(new_n512_)
  );


  anb1
  g440
  (
    .dina(new_n511_),
    .dinb(new_n512_),
    .dout(new_n513_)
  );


  anb1
  g441
  (
    .dina(G24_spl_1),
    .dinb(new_n513_),
    .dout(new_n514_)
  );


  anb2
  g442
  (
    .dina(new_n185__spl_1),
    .dinb(new_n210__spl_1),
    .dout(new_n515_)
  );


  anb1
  g443
  (
    .dina(new_n236__spl_1),
    .dinb(new_n262__spl_1),
    .dout(new_n516_)
  );


  anb2
  g444
  (
    .dina(new_n515_),
    .dinb(new_n516_),
    .dout(new_n517_)
  );


  anb2
  g445
  (
    .dina(G24_spl_1),
    .dinb(new_n517_),
    .dout(new_n518_)
  );


  anb2
  g446
  (
    .dina(new_n514_),
    .dinb(new_n518_),
    .dout(new_n519_)
  );


  nab2
  g447
  (
    .dina(new_n390__spl_010),
    .dinb(new_n519_),
    .dout(new_n520_)
  );


  anb1
  g448
  (
    .dina(new_n270__spl_),
    .dinb(new_n390__spl_010),
    .dout(new_n521_)
  );


  anb1
  g449
  (
    .dina(new_n520_),
    .dinb(new_n521_),
    .dout(new_n522_)
  );


  anb1
  g450
  (
    .dina(G47_spl_01),
    .dinb(new_n522__spl_0),
    .dout(new_n523_)
  );


  and1
  g451
  (
    .dina(new_n403__spl_00),
    .dinb(new_n480__spl_0),
    .dout(new_n524_)
  );


  and2
  g452
  (
    .dina(new_n403__spl_01),
    .dinb(new_n480__spl_1),
    .dout(new_n525_)
  );


  anb2
  g453
  (
    .dina(new_n524_),
    .dinb(new_n525__spl_),
    .dout(new_n526_)
  );


  nab2
  g454
  (
    .dina(new_n523__spl_),
    .dinb(new_n526__spl_),
    .dout(new_n527_)
  );


  nab1
  g455
  (
    .dina(new_n523__spl_),
    .dinb(new_n526__spl_),
    .dout(new_n528_)
  );


  anb1
  g456
  (
    .dina(new_n527_),
    .dinb(new_n528_),
    .dout(new_n529_)
  );


  nab2
  g457
  (
    .dina(new_n410__spl_001),
    .dinb(new_n529_),
    .dout(new_n530_)
  );


  anb2
  g458
  (
    .dina(new_n510_),
    .dinb(new_n530_),
    .dout(G3529)
  );


  anb2
  g459
  (
    .dina(new_n390__spl_011),
    .dinb(new_n306__spl_),
    .dout(new_n532_)
  );


  anb2
  g460
  (
    .dina(new_n320__spl_0),
    .dinb(new_n532__spl_),
    .dout(new_n533_)
  );


  anb1
  g461
  (
    .dina(new_n320__spl_),
    .dinb(new_n532__spl_),
    .dout(new_n534_)
  );


  anb1
  g462
  (
    .dina(new_n533_),
    .dinb(new_n534_),
    .dout(new_n535_)
  );


  anb1
  g463
  (
    .dina(new_n356__spl_),
    .dinb(new_n389__spl_0),
    .dout(new_n536_)
  );


  nab2
  g464
  (
    .dina(new_n370__spl_0),
    .dinb(new_n536__spl_),
    .dout(new_n537_)
  );


  nab1
  g465
  (
    .dina(new_n370__spl_),
    .dinb(new_n536__spl_),
    .dout(new_n538_)
  );


  anb1
  g466
  (
    .dina(new_n537_),
    .dinb(new_n538_),
    .dout(new_n539_)
  );


  and1
  g467
  (
    .dina(new_n535__spl_00),
    .dinb(new_n539__spl_00),
    .dout(new_n540_)
  );


  anb2
  g468
  (
    .dina(new_n480__spl_1),
    .dinb(new_n522__spl_0),
    .dout(new_n541_)
  );


  anb1
  g469
  (
    .dina(new_n540__spl_),
    .dinb(new_n541__spl_),
    .dout(new_n542_)
  );


  and1
  g470
  (
    .dina(new_n373__spl_1),
    .dinb(new_n522__spl_),
    .dout(new_n543_)
  );


  anb2
  g471
  (
    .dina(new_n542__spl_),
    .dinb(new_n543__spl_0),
    .dout(new_n544_)
  );


  anb1
  g472
  (
    .dina(new_n542__spl_),
    .dinb(new_n543__spl_0),
    .dout(new_n545_)
  );


  anb1
  g473
  (
    .dina(new_n544_),
    .dinb(new_n545_),
    .dout(new_n546_)
  );


  anb1
  g474
  (
    .dina(G47_spl_10),
    .dinb(new_n546_),
    .dout(new_n547_)
  );


  anb1
  g475
  (
    .dina(new_n373__spl_1),
    .dinb(new_n403__spl_01),
    .dout(new_n548_)
  );


  anb1
  g476
  (
    .dina(new_n387__spl_),
    .dinb(new_n548_),
    .dout(new_n549_)
  );


  anb1
  g477
  (
    .dina(new_n390__spl_011),
    .dinb(new_n297__spl_),
    .dout(new_n550_)
  );


  anb2
  g478
  (
    .dina(new_n550__spl_0),
    .dinb(new_n540__spl_),
    .dout(new_n551_)
  );


  nor2
  g479
  (
    .dina(new_n319__spl_),
    .dinb(new_n390__spl_100),
    .dout(new_n552_)
  );


  anb1
  g480
  (
    .dina(new_n539__spl_00),
    .dinb(new_n552__spl_),
    .dout(new_n553_)
  );


  anb2
  g481
  (
    .dina(new_n369__spl_),
    .dinb(new_n389__spl_1),
    .dout(new_n554_)
  );


  anb2
  g482
  (
    .dina(new_n553_),
    .dinb(new_n554_),
    .dout(new_n555_)
  );


  anb1
  g483
  (
    .dina(new_n551_),
    .dinb(new_n555_),
    .dout(new_n556_)
  );


  anb1
  g484
  (
    .dina(new_n549__spl_0),
    .dinb(new_n556__spl_0),
    .dout(new_n557_)
  );


  anb2
  g485
  (
    .dina(new_n549__spl_0),
    .dinb(new_n556__spl_0),
    .dout(new_n558_)
  );


  anb2
  g486
  (
    .dina(new_n557_),
    .dinb(new_n558_),
    .dout(new_n559_)
  );


  anb1
  g487
  (
    .dina(new_n547__spl_),
    .dinb(new_n559__spl_),
    .dout(new_n560_)
  );


  anb2
  g488
  (
    .dina(new_n547__spl_),
    .dinb(new_n559__spl_),
    .dout(new_n561_)
  );


  anb2
  g489
  (
    .dina(new_n560_),
    .dinb(new_n561_),
    .dout(new_n562_)
  );


  anb2
  g490
  (
    .dina(new_n96__spl_0),
    .dinb(new_n100__spl_0),
    .dout(new_n563_)
  );


  anb1
  g491
  (
    .dina(new_n562_),
    .dinb(new_n563_),
    .dout(new_n564_)
  );


  anb2
  g492
  (
    .dina(G14_spl_100),
    .dinb(new_n96__spl_),
    .dout(new_n565_)
  );


  anb2
  g493
  (
    .dina(new_n565_),
    .dinb(new_n248__spl_),
    .dout(new_n566_)
  );


  anb2
  g494
  (
    .dina(G10_spl_101),
    .dinb(new_n351__spl_),
    .dout(new_n567_)
  );


  anb2
  g495
  (
    .dina(G7_spl_100),
    .dinb(new_n567_),
    .dout(new_n568_)
  );


  nor2
  g496
  (
    .dina(G7_spl_101),
    .dinb(G9_spl_101),
    .dout(new_n569_)
  );


  anb2
  g497
  (
    .dina(new_n100__spl_),
    .dinb(new_n569_),
    .dout(new_n570_)
  );


  anb1
  g498
  (
    .dina(new_n568_),
    .dinb(new_n570_),
    .dout(new_n571_)
  );


  anb1
  g499
  (
    .dina(new_n566_),
    .dinb(new_n571_),
    .dout(new_n572_)
  );


  anb2
  g500
  (
    .dina(new_n564_),
    .dinb(new_n572_),
    .dout(G3530)
  );


  anb2
  g501
  (
    .dina(new_n390__spl_100),
    .dinb(new_n226__spl_),
    .dout(new_n574_)
  );


  nab1
  g502
  (
    .dina(new_n241__spl_1),
    .dinb(new_n574__spl_),
    .dout(new_n575_)
  );


  nab2
  g503
  (
    .dina(new_n241__spl_1),
    .dinb(new_n574__spl_),
    .dout(new_n576_)
  );


  anb2
  g504
  (
    .dina(new_n575_),
    .dinb(new_n576_),
    .dout(new_n577_)
  );


  and2
  g505
  (
    .dina(new_n414__spl_0),
    .dinb(new_n577__spl_0),
    .dout(new_n578_)
  );


  and2
  g506
  (
    .dina(G39_spl_01),
    .dinb(G43_spl_0),
    .dout(new_n579_)
  );


  anb2
  g507
  (
    .dina(new_n433__spl_010),
    .dinb(new_n579_),
    .dout(new_n580_)
  );


  nab1
  g508
  (
    .dina(G13_spl_110),
    .dinb(new_n445__spl_001),
    .dout(new_n581_)
  );


  anb2
  g509
  (
    .dina(new_n430__spl_010),
    .dinb(G42_spl_0),
    .dout(new_n582_)
  );


  anb2
  g510
  (
    .dina(G40_spl_01),
    .dinb(G12_spl_101),
    .dout(new_n583_)
  );


  and1
  g511
  (
    .dina(new_n437__spl_010),
    .dinb(new_n583__spl_),
    .dout(new_n584_)
  );


  anb1
  g512
  (
    .dina(new_n580_),
    .dinb(new_n584_),
    .dout(new_n585_)
  );


  anb2
  g513
  (
    .dina(new_n581_),
    .dinb(new_n582_),
    .dout(new_n586_)
  );


  anb1
  g514
  (
    .dina(new_n585_),
    .dinb(new_n586_),
    .dout(new_n587_)
  );


  nab1
  g515
  (
    .dina(G14_spl_101),
    .dinb(new_n439__spl_010),
    .dout(new_n588_)
  );


  anb1
  g516
  (
    .dina(G41_spl_01),
    .dinb(new_n435__spl_010),
    .dout(new_n589_)
  );


  anb1
  g517
  (
    .dina(G4_spl_1011),
    .dinb(new_n589_),
    .dout(new_n590_)
  );


  anb2
  g518
  (
    .dina(new_n588_),
    .dinb(new_n590_),
    .dout(new_n591_)
  );


  anb1
  g519
  (
    .dina(new_n587_),
    .dinb(new_n591_),
    .dout(new_n592_)
  );


  anb1
  g520
  (
    .dina(G20_spl_00),
    .dinb(new_n430__spl_010),
    .dout(new_n593_)
  );


  anb1
  g521
  (
    .dina(G7_spl_101),
    .dinb(G19_spl_0),
    .dout(new_n594_)
  );


  and2
  g522
  (
    .dina(new_n433__spl_010),
    .dinb(new_n594__spl_),
    .dout(new_n595_)
  );


  anb2
  g523
  (
    .dina(new_n593_),
    .dinb(new_n595_),
    .dout(new_n596_)
  );


  anb2
  g524
  (
    .dina(new_n435__spl_010),
    .dinb(G21_spl_01),
    .dout(new_n597_)
  );


  anb1
  g525
  (
    .dina(G10_spl_101),
    .dinb(G22_spl_01),
    .dout(new_n598_)
  );


  anb1
  g526
  (
    .dina(new_n437__spl_011),
    .dinb(new_n598_),
    .dout(new_n599_)
  );


  anb1
  g527
  (
    .dina(new_n597_),
    .dinb(new_n599_),
    .dout(new_n600_)
  );


  anb2
  g528
  (
    .dina(new_n596_),
    .dinb(new_n600_),
    .dout(new_n601_)
  );


  anb2
  g529
  (
    .dina(G8_spl_101),
    .dinb(new_n439__spl_010),
    .dout(new_n602_)
  );


  nab1
  g530
  (
    .dina(G9_spl_110),
    .dinb(new_n445__spl_010),
    .dout(new_n603_)
  );


  and2
  g531
  (
    .dina(G4_spl_1100),
    .dinb(new_n603__spl_),
    .dout(new_n604_)
  );


  anb1
  g532
  (
    .dina(new_n602_),
    .dinb(new_n604_),
    .dout(new_n605_)
  );


  anb2
  g533
  (
    .dina(new_n601_),
    .dinb(new_n605_),
    .dout(new_n606_)
  );


  anb2
  g534
  (
    .dina(new_n592_),
    .dinb(new_n606_),
    .dout(new_n607_)
  );


  anb2
  g535
  (
    .dina(new_n417__spl_01),
    .dinb(new_n607_),
    .dout(new_n608_)
  );


  anb2
  g536
  (
    .dina(new_n410__spl_01),
    .dinb(new_n608_),
    .dout(new_n609_)
  );


  anb1
  g537
  (
    .dina(new_n578_),
    .dinb(new_n609_),
    .dout(new_n610_)
  );


  and2
  g538
  (
    .dina(new_n253__spl_),
    .dinb(new_n390__spl_101),
    .dout(new_n611_)
  );


  anb2
  g539
  (
    .dina(new_n267__spl_0),
    .dinb(new_n611__spl_),
    .dout(new_n612_)
  );


  anb1
  g540
  (
    .dina(new_n267__spl_),
    .dinb(new_n611__spl_),
    .dout(new_n613_)
  );


  anb1
  g541
  (
    .dina(new_n612_),
    .dinb(new_n613_),
    .dout(new_n614_)
  );


  anb1
  g542
  (
    .dina(G3526_spl_),
    .dinb(new_n614__spl_00),
    .dout(new_n615_)
  );


  anb1
  g543
  (
    .dina(new_n390__spl_101),
    .dinb(new_n266__spl_),
    .dout(new_n616_)
  );


  anb1
  g544
  (
    .dina(new_n390__spl_11),
    .dinb(new_n191__spl_),
    .dout(new_n617_)
  );


  anb1
  g545
  (
    .dina(new_n394__spl_0),
    .dinb(new_n617__spl_),
    .dout(new_n618_)
  );


  anb2
  g546
  (
    .dina(new_n214__spl_),
    .dinb(new_n390__spl_11),
    .dout(new_n619_)
  );


  anb2
  g547
  (
    .dina(new_n618__spl_),
    .dinb(new_n619_),
    .dout(new_n620_)
  );


  anb2
  g548
  (
    .dina(new_n614__spl_00),
    .dinb(new_n620__spl_),
    .dout(new_n621_)
  );


  anb2
  g549
  (
    .dina(new_n616_),
    .dinb(new_n621_),
    .dout(new_n622_)
  );


  anb1
  g550
  (
    .dina(new_n577__spl_0),
    .dinb(new_n622__spl_),
    .dout(new_n623_)
  );


  anb2
  g551
  (
    .dina(new_n577__spl_),
    .dinb(new_n622__spl_),
    .dout(new_n624_)
  );


  anb2
  g552
  (
    .dina(new_n623_),
    .dinb(new_n624_),
    .dout(new_n625_)
  );


  anb2
  g553
  (
    .dina(new_n615__spl_),
    .dinb(new_n625__spl_),
    .dout(new_n626_)
  );


  anb1
  g554
  (
    .dina(new_n615__spl_),
    .dinb(new_n625__spl_),
    .dout(new_n627_)
  );


  anb1
  g555
  (
    .dina(new_n626_),
    .dinb(new_n627_),
    .dout(new_n628_)
  );


  anb2
  g556
  (
    .dina(new_n394__spl_1),
    .dinb(new_n617__spl_),
    .dout(new_n629_)
  );


  nab1
  g557
  (
    .dina(new_n618__spl_),
    .dinb(new_n629_),
    .dout(new_n630_)
  );


  anb1
  g558
  (
    .dina(new_n411__spl_0),
    .dinb(new_n630__spl_),
    .dout(new_n631_)
  );


  anb2
  g559
  (
    .dina(new_n411__spl_),
    .dinb(new_n630__spl_),
    .dout(new_n632_)
  );


  anb2
  g560
  (
    .dina(new_n631_),
    .dinb(new_n632_),
    .dout(new_n633_)
  );


  anb2
  g561
  (
    .dina(G3526_spl_),
    .dinb(new_n620__spl_),
    .dout(new_n634_)
  );


  nab2
  g562
  (
    .dina(new_n614__spl_0),
    .dinb(new_n634__spl_),
    .dout(new_n635_)
  );


  nab1
  g563
  (
    .dina(new_n614__spl_1),
    .dinb(new_n634__spl_),
    .dout(new_n636_)
  );


  anb1
  g564
  (
    .dina(new_n635_),
    .dinb(new_n636_),
    .dout(new_n637_)
  );


  anb1
  g565
  (
    .dina(new_n633__spl_0),
    .dinb(new_n637__spl_0),
    .dout(new_n638_)
  );


  anb2
  g566
  (
    .dina(new_n638_),
    .dinb(new_n403__spl_10),
    .dout(new_n639_)
  );


  anb2
  g567
  (
    .dina(new_n401__spl_01),
    .dinb(new_n639_),
    .dout(new_n640_)
  );


  anb2
  g568
  (
    .dina(new_n409__spl_00),
    .dinb(new_n640_),
    .dout(new_n641_)
  );


  anb2
  g569
  (
    .dina(new_n628_),
    .dinb(new_n641_),
    .dout(new_n642_)
  );


  anb2
  g570
  (
    .dina(new_n610_),
    .dinb(new_n642_),
    .dout(G3531)
  );


  nor1
  g571
  (
    .dina(new_n394__spl_1),
    .dinb(new_n414__spl_1),
    .dout(new_n644_)
  );


  anb1
  g572
  (
    .dina(G14_spl_101),
    .dinb(G42_spl_1),
    .dout(new_n645_)
  );


  nab2
  g573
  (
    .dina(new_n437__spl_011),
    .dinb(new_n645_),
    .dout(new_n646_)
  );


  anb1
  g574
  (
    .dina(G43_spl_1),
    .dinb(new_n435__spl_011),
    .dout(new_n647_)
  );


  and2
  g575
  (
    .dina(G41_spl_10),
    .dinb(G45_spl_),
    .dout(new_n648_)
  );


  nab1
  g576
  (
    .dina(new_n433__spl_011),
    .dinb(new_n648_),
    .dout(new_n649_)
  );


  and1
  g577
  (
    .dina(G39_spl_01),
    .dinb(new_n445__spl_010),
    .dout(new_n650_)
  );


  and1
  g578
  (
    .dina(G40_spl_10),
    .dinb(new_n439__spl_011),
    .dout(new_n651_)
  );


  anb2
  g579
  (
    .dina(new_n430__spl_011),
    .dinb(G44_spl_0),
    .dout(new_n652_)
  );


  anb1
  g580
  (
    .dina(new_n646_),
    .dinb(new_n649_),
    .dout(new_n653_)
  );


  anb2
  g581
  (
    .dina(new_n647_),
    .dinb(new_n652_),
    .dout(new_n654_)
  );


  anb1
  g582
  (
    .dina(new_n653_),
    .dinb(new_n654_),
    .dout(new_n655_)
  );


  anb1
  g583
  (
    .dina(G4_spl_1100),
    .dinb(new_n650_),
    .dout(new_n656_)
  );


  anb2
  g584
  (
    .dina(new_n651_),
    .dinb(new_n656_),
    .dout(new_n657_)
  );


  anb1
  g585
  (
    .dina(new_n655_),
    .dinb(new_n657_),
    .dout(new_n658_)
  );


  nab1
  g586
  (
    .dina(G10_spl_110),
    .dinb(new_n439__spl_011),
    .dout(new_n659_)
  );


  anb2
  g587
  (
    .dina(G12_spl_11),
    .dinb(new_n437__spl_100),
    .dout(new_n660_)
  );


  nab1
  g588
  (
    .dina(G4_spl_1101),
    .dinb(new_n660_),
    .dout(new_n661_)
  );


  anb2
  g589
  (
    .dina(new_n659_),
    .dinb(new_n661_),
    .dout(new_n662_)
  );


  anb2
  g590
  (
    .dina(G11_spl_101),
    .dinb(new_n445__spl_011),
    .dout(new_n663_)
  );


  nab1
  g591
  (
    .dina(G8_spl_11),
    .dinb(new_n437__spl_100),
    .dout(new_n664_)
  );


  anb1
  g592
  (
    .dina(new_n663__spl_),
    .dinb(new_n664__spl_),
    .dout(new_n665_)
  );


  nor1
  g593
  (
    .dina(G7_spl_110),
    .dinb(new_n435__spl_011),
    .dout(new_n666_)
  );


  anb2
  g594
  (
    .dina(new_n430__spl_011),
    .dinb(G22_spl_01),
    .dout(new_n667_)
  );


  anb2
  g595
  (
    .dina(new_n666_),
    .dinb(new_n667_),
    .dout(new_n668_)
  );


  anb2
  g596
  (
    .dina(G21_spl_01),
    .dinb(G9_spl_110),
    .dout(new_n669_)
  );


  anb2
  g597
  (
    .dina(new_n433__spl_011),
    .dinb(new_n669_),
    .dout(new_n670_)
  );


  anb2
  g598
  (
    .dina(new_n668_),
    .dinb(new_n670_),
    .dout(new_n671_)
  );


  anb1
  g599
  (
    .dina(new_n665_),
    .dinb(new_n671_),
    .dout(new_n672_)
  );


  anb2
  g600
  (
    .dina(new_n662__spl_),
    .dinb(new_n672_),
    .dout(new_n673_)
  );


  anb2
  g601
  (
    .dina(new_n658_),
    .dinb(new_n673_),
    .dout(new_n674_)
  );


  anb2
  g602
  (
    .dina(new_n417__spl_01),
    .dinb(new_n674_),
    .dout(new_n675_)
  );


  anb1
  g603
  (
    .dina(new_n675_),
    .dinb(new_n410__spl_01),
    .dout(new_n676_)
  );


  anb2
  g604
  (
    .dina(new_n644_),
    .dinb(new_n676_),
    .dout(new_n677_)
  );


  nab2
  g605
  (
    .dina(new_n403__spl_10),
    .dinb(new_n633__spl_0),
    .dout(new_n678_)
  );


  and1
  g606
  (
    .dina(new_n409__spl_01),
    .dinb(new_n633__spl_1),
    .dout(new_n679_)
  );


  nab1
  g607
  (
    .dina(new_n403__spl_1),
    .dinb(new_n633__spl_1),
    .dout(new_n680_)
  );


  anb1
  g608
  (
    .dina(new_n678_),
    .dinb(new_n680__spl_0),
    .dout(new_n681_)
  );


  anb1
  g609
  (
    .dina(new_n681_),
    .dinb(new_n401__spl_01),
    .dout(new_n682_)
  );


  anb1
  g610
  (
    .dina(new_n677_),
    .dinb(new_n679_),
    .dout(new_n683_)
  );


  anb2
  g611
  (
    .dina(new_n682_),
    .dinb(new_n683_),
    .dout(G3532)
  );


  anb1
  g612
  (
    .dina(new_n637__spl_0),
    .dinb(new_n680__spl_0),
    .dout(new_n685_)
  );


  anb2
  g613
  (
    .dina(new_n637__spl_1),
    .dinb(new_n680__spl_),
    .dout(new_n686_)
  );


  anb2
  g614
  (
    .dina(new_n685_),
    .dinb(new_n686_),
    .dout(new_n687_)
  );


  nab1
  g615
  (
    .dina(new_n401__spl_10),
    .dinb(new_n687_),
    .dout(new_n688_)
  );


  nab2
  g616
  (
    .dina(new_n409__spl_01),
    .dinb(new_n637__spl_1),
    .dout(new_n689_)
  );


  anb2
  g617
  (
    .dina(new_n414__spl_1),
    .dinb(new_n614__spl_1),
    .dout(new_n690_)
  );


  and2
  g618
  (
    .dina(G40_spl_10),
    .dinb(G44_spl_),
    .dout(new_n691_)
  );


  anb2
  g619
  (
    .dina(new_n433__spl_100),
    .dinb(new_n691_),
    .dout(new_n692_)
  );


  anb2
  g620
  (
    .dina(G41_spl_10),
    .dinb(G13_spl_110),
    .dout(new_n693_)
  );


  nab1
  g621
  (
    .dina(G14_spl_110),
    .dinb(new_n445__spl_011),
    .dout(new_n694_)
  );


  anb1
  g622
  (
    .dina(G42_spl_1),
    .dinb(new_n435__spl_100),
    .dout(new_n695_)
  );


  and1
  g623
  (
    .dina(G39_spl_10),
    .dinb(new_n439__spl_100),
    .dout(new_n696_)
  );


  anb2
  g624
  (
    .dina(new_n430__spl_100),
    .dinb(G43_spl_1),
    .dout(new_n697_)
  );


  nor2
  g625
  (
    .dina(G41_spl_1),
    .dinb(new_n437__spl_101),
    .dout(new_n698_)
  );


  anb2
  g626
  (
    .dina(new_n695_),
    .dinb(new_n698_),
    .dout(new_n699_)
  );


  anb1
  g627
  (
    .dina(new_n692_),
    .dinb(new_n699_),
    .dout(new_n700_)
  );


  anb1
  g628
  (
    .dina(G4_spl_1101),
    .dinb(new_n456__spl_),
    .dout(new_n701_)
  );


  anb2
  g629
  (
    .dina(new_n694_),
    .dinb(new_n697_),
    .dout(new_n702_)
  );


  anb1
  g630
  (
    .dina(new_n701__spl_),
    .dinb(new_n702_),
    .dout(new_n703_)
  );


  anb2
  g631
  (
    .dina(new_n696_),
    .dinb(new_n703_),
    .dout(new_n704_)
  );


  anb1
  g632
  (
    .dina(new_n700_),
    .dinb(new_n704_),
    .dout(new_n705_)
  );


  anb1
  g633
  (
    .dina(G22_spl_10),
    .dinb(new_n435__spl_100),
    .dout(new_n706_)
  );


  and1
  g634
  (
    .dina(G7_spl_110),
    .dinb(G11_spl_11),
    .dout(new_n707_)
  );


  nab2
  g635
  (
    .dina(new_n437__spl_101),
    .dinb(new_n707_),
    .dout(new_n708_)
  );


  anb2
  g636
  (
    .dina(new_n430__spl_100),
    .dinb(G21_spl_10),
    .dout(new_n709_)
  );


  nab1
  g637
  (
    .dina(G10_spl_110),
    .dinb(new_n445__spl_10),
    .dout(new_n710_)
  );


  anb2
  g638
  (
    .dina(G9_spl_11),
    .dinb(new_n439__spl_100),
    .dout(new_n711_)
  );


  anb2
  g639
  (
    .dina(G20_spl_0),
    .dinb(G8_spl_11),
    .dout(new_n712_)
  );


  anb2
  g640
  (
    .dina(new_n433__spl_100),
    .dinb(new_n712__spl_),
    .dout(new_n713_)
  );


  anb2
  g641
  (
    .dina(new_n710__spl_),
    .dinb(new_n713_),
    .dout(new_n714_)
  );


  anb2
  g642
  (
    .dina(new_n706_),
    .dinb(new_n709_),
    .dout(new_n715_)
  );


  nab1
  g643
  (
    .dina(G4_spl_1110),
    .dinb(new_n711_),
    .dout(new_n716_)
  );


  anb2
  g644
  (
    .dina(new_n715_),
    .dinb(new_n716_),
    .dout(new_n717_)
  );


  anb1
  g645
  (
    .dina(new_n708_),
    .dinb(new_n714_),
    .dout(new_n718_)
  );


  anb2
  g646
  (
    .dina(new_n717_),
    .dinb(new_n718_),
    .dout(new_n719_)
  );


  anb2
  g647
  (
    .dina(new_n705_),
    .dinb(new_n719_),
    .dout(new_n720_)
  );


  anb2
  g648
  (
    .dina(new_n417__spl_10),
    .dinb(new_n720_),
    .dout(new_n721_)
  );


  anb2
  g649
  (
    .dina(new_n410__spl_10),
    .dinb(new_n721_),
    .dout(new_n722_)
  );


  anb1
  g650
  (
    .dina(new_n690_),
    .dinb(new_n722_),
    .dout(new_n723_)
  );


  anb1
  g651
  (
    .dina(new_n689_),
    .dinb(new_n723_),
    .dout(new_n724_)
  );


  anb2
  g652
  (
    .dina(new_n688_),
    .dinb(new_n724_),
    .dout(G3533)
  );


  nab2
  g653
  (
    .dina(G47_spl_10),
    .dinb(new_n541__spl_),
    .dout(new_n726_)
  );


  anb1
  g654
  (
    .dina(new_n535__spl_00),
    .dinb(new_n726__spl_),
    .dout(new_n727_)
  );


  anb1
  g655
  (
    .dina(new_n535__spl_0),
    .dinb(new_n550__spl_0),
    .dout(new_n728_)
  );


  nab2
  g656
  (
    .dina(new_n552__spl_),
    .dinb(new_n728_),
    .dout(new_n729_)
  );


  anb1
  g657
  (
    .dina(new_n539__spl_0),
    .dinb(new_n729__spl_),
    .dout(new_n730_)
  );


  anb2
  g658
  (
    .dina(new_n539__spl_1),
    .dinb(new_n729__spl_),
    .dout(new_n731_)
  );


  anb2
  g659
  (
    .dina(new_n730_),
    .dinb(new_n731_),
    .dout(new_n732_)
  );


  anb1
  g660
  (
    .dina(new_n727__spl_0),
    .dinb(new_n732__spl_),
    .dout(new_n733_)
  );


  anb2
  g661
  (
    .dina(new_n727__spl_0),
    .dinb(new_n732__spl_),
    .dout(new_n734_)
  );


  nab1
  g662
  (
    .dina(new_n733__spl_0),
    .dinb(new_n734_),
    .dout(new_n735_)
  );


  nab2
  g663
  (
    .dina(new_n525__spl_),
    .dinb(new_n550__spl_),
    .dout(new_n736_)
  );


  anb2
  g664
  (
    .dina(new_n535__spl_1),
    .dinb(new_n726__spl_),
    .dout(new_n737_)
  );


  anb2
  g665
  (
    .dina(new_n727__spl_),
    .dinb(new_n737_),
    .dout(new_n738_)
  );


  anb2
  g666
  (
    .dina(new_n736__spl_),
    .dinb(new_n738__spl_),
    .dout(new_n739_)
  );


  anb1
  g667
  (
    .dina(new_n736__spl_),
    .dinb(new_n738__spl_),
    .dout(new_n740_)
  );


  anb1
  g668
  (
    .dina(new_n739_),
    .dinb(new_n740_),
    .dout(new_n741_)
  );


  and1
  g669
  (
    .dina(G47_spl_1),
    .dinb(new_n543__spl_),
    .dout(new_n742_)
  );


  anb2
  g670
  (
    .dina(new_n549__spl_),
    .dinb(new_n742_),
    .dout(new_n743_)
  );


  nab1
  g671
  (
    .dina(new_n741__spl_0),
    .dinb(new_n743__spl_0),
    .dout(new_n744_)
  );


  anb1
  g672
  (
    .dina(new_n735__spl_0),
    .dinb(new_n744__spl_0),
    .dout(new_n745_)
  );


  anb2
  g673
  (
    .dina(new_n735__spl_0),
    .dinb(new_n744__spl_0),
    .dout(new_n746_)
  );


  anb2
  g674
  (
    .dina(new_n745_),
    .dinb(new_n746_),
    .dout(new_n747_)
  );


  nab1
  g675
  (
    .dina(new_n401__spl_10),
    .dinb(new_n747_),
    .dout(new_n748_)
  );


  nab1
  g676
  (
    .dina(new_n476__spl_0),
    .dinb(new_n539__spl_1),
    .dout(new_n749_)
  );


  nor1
  g677
  (
    .dina(G14_spl_110),
    .dinb(new_n435__spl_101),
    .dout(new_n750_)
  );


  anb2
  g678
  (
    .dina(new_n430__spl_101),
    .dinb(G39_spl_10),
    .dout(new_n751_)
  );


  anb2
  g679
  (
    .dina(new_n433__spl_101),
    .dinb(new_n583__spl_),
    .dout(new_n752_)
  );


  anb2
  g680
  (
    .dina(new_n750_),
    .dinb(new_n751_),
    .dout(new_n753_)
  );


  anb1
  g681
  (
    .dina(new_n752_),
    .dinb(new_n753_),
    .dout(new_n754_)
  );


  nab2
  g682
  (
    .dina(new_n458__spl_),
    .dinb(new_n710__spl_),
    .dout(new_n755_)
  );


  anb1
  g683
  (
    .dina(new_n701__spl_),
    .dinb(new_n755_),
    .dout(new_n756_)
  );


  anb2
  g684
  (
    .dina(new_n460__spl_),
    .dinb(new_n756_),
    .dout(new_n757_)
  );


  anb1
  g685
  (
    .dina(new_n754_),
    .dinb(new_n757_),
    .dout(new_n758_)
  );


  anb1
  g686
  (
    .dina(G18_spl_0),
    .dinb(new_n435__spl_101),
    .dout(new_n759_)
  );


  and2
  g687
  (
    .dina(G16_spl_),
    .dinb(G20_spl_1),
    .dout(new_n760_)
  );


  anb2
  g688
  (
    .dina(new_n433__spl_101),
    .dinb(new_n760_),
    .dout(new_n761_)
  );


  nor2
  g689
  (
    .dina(G22_spl_10),
    .dinb(new_n445__spl_10),
    .dout(new_n762_)
  );


  anb1
  g690
  (
    .dina(new_n437__spl_110),
    .dinb(new_n594__spl_),
    .dout(new_n763_)
  );


  anb1
  g691
  (
    .dina(new_n761_),
    .dinb(new_n763_),
    .dout(new_n764_)
  );


  and1
  g692
  (
    .dina(G21_spl_10),
    .dinb(new_n439__spl_101),
    .dout(new_n765_)
  );


  anb2
  g693
  (
    .dina(new_n430__spl_101),
    .dinb(G17_spl_0),
    .dout(new_n766_)
  );


  anb2
  g694
  (
    .dina(new_n765_),
    .dinb(new_n766_),
    .dout(new_n767_)
  );


  nab1
  g695
  (
    .dina(G4_spl_1110),
    .dinb(new_n762_),
    .dout(new_n768_)
  );


  anb2
  g696
  (
    .dina(new_n759_),
    .dinb(new_n764_),
    .dout(new_n769_)
  );


  anb1
  g697
  (
    .dina(new_n768_),
    .dinb(new_n769_),
    .dout(new_n770_)
  );


  anb2
  g698
  (
    .dina(new_n767_),
    .dinb(new_n770_),
    .dout(new_n771_)
  );


  anb2
  g699
  (
    .dina(new_n758_),
    .dinb(new_n771_),
    .dout(new_n772_)
  );


  anb2
  g700
  (
    .dina(new_n417__spl_10),
    .dinb(new_n772_),
    .dout(new_n773_)
  );


  anb1
  g701
  (
    .dina(new_n773_),
    .dinb(new_n410__spl_10),
    .dout(new_n774_)
  );


  anb2
  g702
  (
    .dina(new_n749_),
    .dinb(new_n774_),
    .dout(new_n775_)
  );


  anb1
  g703
  (
    .dina(new_n409__spl_10),
    .dinb(new_n735__spl_1),
    .dout(new_n776_)
  );


  anb1
  g704
  (
    .dina(new_n775_),
    .dinb(new_n776_),
    .dout(new_n777_)
  );


  anb1
  g705
  (
    .dina(new_n777__spl_),
    .dinb(new_n748__spl_),
    .dout(new_n778_)
  );


  anb2
  g706
  (
    .dina(new_n748__spl_),
    .dinb(new_n777__spl_),
    .dout(G3534)
  );


  anb2
  g707
  (
    .dina(new_n389__spl_1),
    .dinb(new_n330__spl_),
    .dout(new_n780_)
  );


  nab1
  g708
  (
    .dina(new_n344__spl_1),
    .dinb(new_n780__spl_),
    .dout(new_n781_)
  );


  nab2
  g709
  (
    .dina(new_n344__spl_1),
    .dinb(new_n780__spl_),
    .dout(new_n782_)
  );


  anb2
  g710
  (
    .dina(new_n781_),
    .dinb(new_n782_),
    .dout(new_n783_)
  );


  and2
  g711
  (
    .dina(new_n476__spl_1),
    .dinb(new_n783__spl_0),
    .dout(new_n784_)
  );


  nor1
  g712
  (
    .dina(G5_spl_1),
    .dinb(G7_spl_111),
    .dout(new_n785_)
  );


  anb1
  g713
  (
    .dina(G17_spl_0),
    .dinb(new_n435__spl_110),
    .dout(new_n786_)
  );


  nor1
  g714
  (
    .dina(G18_spl_1),
    .dinb(G22_spl_11),
    .dout(new_n787_)
  );


  anb1
  g715
  (
    .dina(new_n437__spl_110),
    .dinb(new_n787_),
    .dout(new_n788_)
  );


  and2
  g716
  (
    .dina(G15),
    .dinb(G19_spl_1),
    .dout(new_n789_)
  );


  anb2
  g717
  (
    .dina(new_n433__spl_110),
    .dinb(new_n789_),
    .dout(new_n790_)
  );


  nor2
  g718
  (
    .dina(G21_spl_11),
    .dinb(new_n445__spl_11),
    .dout(new_n791_)
  );


  and1
  g719
  (
    .dina(G20_spl_1),
    .dinb(new_n439__spl_101),
    .dout(new_n792_)
  );


  anb1
  g720
  (
    .dina(G16_spl_),
    .dinb(new_n430__spl_110),
    .dout(new_n793_)
  );


  anb2
  g721
  (
    .dina(new_n788_),
    .dinb(new_n790_),
    .dout(new_n794_)
  );


  anb1
  g722
  (
    .dina(new_n791_),
    .dinb(new_n793_),
    .dout(new_n795_)
  );


  anb2
  g723
  (
    .dina(new_n794_),
    .dinb(new_n795_),
    .dout(new_n796_)
  );


  anb1
  g724
  (
    .dina(new_n170__spl_),
    .dinb(new_n786_),
    .dout(new_n797_)
  );


  anb1
  g725
  (
    .dina(new_n797_),
    .dinb(new_n792_),
    .dout(new_n798_)
  );


  anb2
  g726
  (
    .dina(new_n796_),
    .dinb(new_n798_),
    .dout(new_n799_)
  );


  anb2
  g727
  (
    .dina(new_n785_),
    .dinb(new_n799_),
    .dout(new_n800_)
  );


  anb1
  g728
  (
    .dina(G5_spl_1),
    .dinb(new_n603__spl_),
    .dout(new_n801_)
  );


  nor1
  g729
  (
    .dina(G13_spl_11),
    .dinb(new_n435__spl_110),
    .dout(new_n802_)
  );


  anb2
  g730
  (
    .dina(G39_spl_11),
    .dinb(G11_spl_11),
    .dout(new_n803_)
  );


  anb2
  g731
  (
    .dina(new_n433__spl_110),
    .dinb(new_n803_),
    .dout(new_n804_)
  );


  and2
  g732
  (
    .dina(G14_spl_111),
    .dinb(new_n430__spl_110),
    .dout(new_n805_)
  );


  anb2
  g733
  (
    .dina(new_n802_),
    .dinb(new_n805_),
    .dout(new_n806_)
  );


  anb2
  g734
  (
    .dina(new_n664__spl_),
    .dinb(new_n804_),
    .dout(new_n807_)
  );


  and2
  g735
  (
    .dina(new_n806_),
    .dinb(new_n807_),
    .dout(new_n808_)
  );


  anb1
  g736
  (
    .dina(new_n801_),
    .dinb(new_n808_),
    .dout(new_n809_)
  );


  anb2
  g737
  (
    .dina(new_n662__spl_),
    .dinb(new_n809_),
    .dout(new_n810_)
  );


  anb2
  g738
  (
    .dina(new_n800_),
    .dinb(new_n810_),
    .dout(new_n811_)
  );


  anb2
  g739
  (
    .dina(new_n417__spl_11),
    .dinb(new_n811_),
    .dout(new_n812_)
  );


  anb2
  g740
  (
    .dina(new_n410__spl_11),
    .dinb(new_n812_),
    .dout(new_n813_)
  );


  anb1
  g741
  (
    .dina(new_n784_),
    .dinb(new_n813_),
    .dout(new_n814_)
  );


  nab1
  g742
  (
    .dina(new_n556__spl_1),
    .dinb(new_n783__spl_0),
    .dout(new_n815_)
  );


  nab2
  g743
  (
    .dina(new_n556__spl_1),
    .dinb(new_n783__spl_),
    .dout(new_n816_)
  );


  anb2
  g744
  (
    .dina(new_n815_),
    .dinb(new_n816_),
    .dout(new_n817_)
  );


  anb2
  g745
  (
    .dina(new_n733__spl_0),
    .dinb(new_n817__spl_),
    .dout(new_n818_)
  );


  anb1
  g746
  (
    .dina(new_n733__spl_),
    .dinb(new_n817__spl_),
    .dout(new_n819_)
  );


  anb1
  g747
  (
    .dina(new_n818_),
    .dinb(new_n819_),
    .dout(new_n820_)
  );


  and2
  g748
  (
    .dina(new_n735__spl_1),
    .dinb(new_n741__spl_0),
    .dout(new_n821_)
  );


  anb2
  g749
  (
    .dina(new_n743__spl_0),
    .dinb(new_n821_),
    .dout(new_n822_)
  );


  anb2
  g750
  (
    .dina(new_n401__spl_11),
    .dinb(new_n822_),
    .dout(new_n823_)
  );


  anb2
  g751
  (
    .dina(new_n409__spl_10),
    .dinb(new_n823_),
    .dout(new_n824_)
  );


  anb2
  g752
  (
    .dina(new_n820_),
    .dinb(new_n824_),
    .dout(new_n825_)
  );


  anb2
  g753
  (
    .dina(new_n814_),
    .dinb(new_n825_),
    .dout(G3535)
  );


  anb2
  g754
  (
    .dina(new_n476__spl_1),
    .dinb(new_n535__spl_1),
    .dout(new_n827_)
  );


  anb2
  g755
  (
    .dina(new_n435__spl_111),
    .dinb(G19_spl_1),
    .dout(new_n828_)
  );


  nab1
  g756
  (
    .dina(G7_spl_111),
    .dinb(new_n445__spl_11),
    .dout(new_n829_)
  );


  nor2
  g757
  (
    .dina(new_n437__spl_111),
    .dinb(new_n712__spl_),
    .dout(new_n830_)
  );


  anb1
  g758
  (
    .dina(G18_spl_1),
    .dinb(new_n430__spl_111),
    .dout(new_n831_)
  );


  anb1
  g759
  (
    .dina(new_n828_),
    .dinb(new_n831_),
    .dout(new_n832_)
  );


  anb2
  g760
  (
    .dina(new_n829_),
    .dinb(new_n830_),
    .dout(new_n833_)
  );


  anb1
  g761
  (
    .dina(new_n832_),
    .dinb(new_n833_),
    .dout(new_n834_)
  );


  and1
  g762
  (
    .dina(G22_spl_11),
    .dinb(new_n439__spl_11),
    .dout(new_n835_)
  );


  and2
  g763
  (
    .dina(G17_spl_),
    .dinb(G21_spl_11),
    .dout(new_n836_)
  );


  anb2
  g764
  (
    .dina(new_n433__spl_111),
    .dinb(new_n836_),
    .dout(new_n837_)
  );


  nab1
  g765
  (
    .dina(G4_spl_1111),
    .dinb(new_n837_),
    .dout(new_n838_)
  );


  anb2
  g766
  (
    .dina(new_n835_),
    .dinb(new_n838_),
    .dout(new_n839_)
  );


  anb1
  g767
  (
    .dina(new_n834_),
    .dinb(new_n839_),
    .dout(new_n840_)
  );


  and1
  g768
  (
    .dina(G10_spl_11),
    .dinb(G14_spl_111),
    .dout(new_n841_)
  );


  anb1
  g769
  (
    .dina(new_n437__spl_111),
    .dinb(new_n841_),
    .dout(new_n842_)
  );


  anb2
  g770
  (
    .dina(new_n430__spl_111),
    .dinb(G40_spl_1),
    .dout(new_n843_)
  );


  anb2
  g771
  (
    .dina(new_n433__spl_111),
    .dinb(new_n693_),
    .dout(new_n844_)
  );


  anb1
  g772
  (
    .dina(G39_spl_11),
    .dinb(new_n435__spl_111),
    .dout(new_n845_)
  );


  anb2
  g773
  (
    .dina(new_n842_),
    .dinb(new_n844_),
    .dout(new_n846_)
  );


  nab1
  g774
  (
    .dina(G12_spl_11),
    .dinb(new_n439__spl_11),
    .dout(new_n847_)
  );


  anb1
  g775
  (
    .dina(new_n663__spl_),
    .dinb(new_n846_),
    .dout(new_n848_)
  );


  anb2
  g776
  (
    .dina(new_n845_),
    .dinb(G4_spl_1111),
    .dout(new_n849_)
  );


  anb1
  g777
  (
    .dina(new_n843_),
    .dinb(new_n847_),
    .dout(new_n850_)
  );


  anb2
  g778
  (
    .dina(new_n849_),
    .dinb(new_n850_),
    .dout(new_n851_)
  );


  anb1
  g779
  (
    .dina(new_n848_),
    .dinb(new_n851_),
    .dout(new_n852_)
  );


  and2
  g780
  (
    .dina(new_n840_),
    .dinb(new_n852_),
    .dout(new_n853_)
  );


  anb2
  g781
  (
    .dina(new_n417__spl_11),
    .dinb(new_n853_),
    .dout(new_n854_)
  );


  anb2
  g782
  (
    .dina(new_n410__spl_11),
    .dinb(new_n854_),
    .dout(new_n855_)
  );


  anb1
  g783
  (
    .dina(new_n827_),
    .dinb(new_n855_),
    .dout(new_n856_)
  );


  anb1
  g784
  (
    .dina(new_n741__spl_1),
    .dinb(new_n743__spl_),
    .dout(new_n857_)
  );


  anb1
  g785
  (
    .dina(new_n409__spl_1),
    .dinb(new_n741__spl_1),
    .dout(new_n858_)
  );


  and2
  g786
  (
    .dina(new_n401__spl_11),
    .dinb(new_n744__spl_),
    .dout(new_n859_)
  );


  anb2
  g787
  (
    .dina(new_n858_),
    .dinb(new_n859_),
    .dout(new_n860_)
  );


  anb2
  g788
  (
    .dina(new_n857_),
    .dinb(new_n860_),
    .dout(new_n861_)
  );


  anb2
  g789
  (
    .dina(new_n856_),
    .dinb(new_n861_),
    .dout(G3536)
  );


  anb1
  g790
  (
    .dina(new_n778__spl_),
    .dinb(G3535_spl_),
    .dout(new_n863_)
  );


  and2
  g791
  (
    .dina(G3529_spl_),
    .dinb(G3536_spl_),
    .dout(new_n864_)
  );


  nor1
  g792
  (
    .dina(G3531_spl_),
    .dinb(G3533_spl_),
    .dout(new_n865_)
  );


  and2
  g793
  (
    .dina(G3528_spl_),
    .dinb(G3532_spl_),
    .dout(new_n866_)
  );


  anb1
  g794
  (
    .dina(new_n865__spl_),
    .dinb(new_n866__spl_),
    .dout(new_n867_)
  );


  anb2
  g795
  (
    .dina(new_n864__spl_),
    .dinb(new_n867_),
    .dout(new_n868_)
  );


  nab2
  g796
  (
    .dina(new_n863__spl_0),
    .dinb(new_n868_),
    .dout(G3537)
  );


  nor2
  g797
  (
    .dina(G27_spl_0),
    .dinb(G48_spl_),
    .dout(new_n870_)
  );


  anb1
  g798
  (
    .dina(new_n863__spl_0),
    .dinb(new_n870__spl_),
    .dout(new_n871_)
  );


  and1
  g799
  (
    .dina(G27_spl_),
    .dinb(G3537),
    .dout(new_n872_)
  );


  anb2
  g800
  (
    .dina(new_n871_),
    .dinb(new_n872_),
    .dout(G3538)
  );


  and1
  g801
  (
    .dina(G3528_spl_),
    .dinb(G3532_spl_),
    .dout(new_n874_)
  );


  nab2
  g802
  (
    .dina(new_n866__spl_),
    .dinb(new_n874_),
    .dout(new_n875_)
  );


  nor2
  g803
  (
    .dina(G3531_spl_),
    .dinb(G3533_spl_),
    .dout(new_n876_)
  );


  anb2
  g804
  (
    .dina(new_n865__spl_),
    .dinb(new_n876_),
    .dout(new_n877_)
  );


  anb2
  g805
  (
    .dina(new_n875__spl_),
    .dinb(new_n877__spl_),
    .dout(new_n878_)
  );


  anb1
  g806
  (
    .dina(new_n875__spl_),
    .dinb(new_n877__spl_),
    .dout(new_n879_)
  );


  anb1
  g807
  (
    .dina(new_n878_),
    .dinb(new_n879_),
    .dout(new_n880_)
  );


  and1
  g808
  (
    .dina(G3529_spl_),
    .dinb(G3536_spl_),
    .dout(new_n881_)
  );


  nab2
  g809
  (
    .dina(new_n864__spl_),
    .dinb(new_n881_),
    .dout(new_n882_)
  );


  anb2
  g810
  (
    .dina(new_n778__spl_),
    .dinb(G3535_spl_),
    .dout(new_n883_)
  );


  anb2
  g811
  (
    .dina(new_n863__spl_),
    .dinb(new_n883_),
    .dout(new_n884_)
  );


  anb1
  g812
  (
    .dina(G50_spl_),
    .dinb(new_n884__spl_0),
    .dout(new_n885_)
  );


  nab1
  g813
  (
    .dina(G50_spl_),
    .dinb(new_n884__spl_0),
    .dout(new_n886_)
  );


  anb1
  g814
  (
    .dina(new_n870__spl_),
    .dinb(new_n885_),
    .dout(new_n887_)
  );


  anb2
  g815
  (
    .dina(new_n886_),
    .dinb(new_n887_),
    .dout(new_n888_)
  );


  anb2
  g816
  (
    .dina(new_n882__spl_0),
    .dinb(new_n888__spl_),
    .dout(new_n889_)
  );


  anb1
  g817
  (
    .dina(new_n882__spl_0),
    .dinb(new_n888__spl_),
    .dout(new_n890_)
  );


  anb1
  g818
  (
    .dina(new_n889_),
    .dinb(new_n890_),
    .dout(new_n891_)
  );


  anb2
  g819
  (
    .dina(new_n880__spl_0),
    .dinb(new_n891__spl_),
    .dout(new_n892_)
  );


  anb1
  g820
  (
    .dina(new_n880__spl_0),
    .dinb(new_n891__spl_),
    .dout(new_n893_)
  );


  nab2
  g821
  (
    .dina(new_n892_),
    .dinb(new_n893_),
    .dout(G3539)
  );


  anb2
  g822
  (
    .dina(new_n882__spl_1),
    .dinb(new_n884__spl_1),
    .dout(new_n895_)
  );


  anb1
  g823
  (
    .dina(new_n882__spl_1),
    .dinb(new_n884__spl_1),
    .dout(new_n896_)
  );


  anb1
  g824
  (
    .dina(new_n895_),
    .dinb(new_n896_),
    .dout(new_n897_)
  );


  anb2
  g825
  (
    .dina(new_n880__spl_1),
    .dinb(new_n897__spl_),
    .dout(new_n898_)
  );


  anb1
  g826
  (
    .dina(new_n880__spl_1),
    .dinb(new_n897__spl_),
    .dout(new_n899_)
  );


  anb1
  g827
  (
    .dina(new_n898_),
    .dinb(new_n899_),
    .dout(G3540)
  );


  splt
  gG7
  (
    .dout(G7_spl_),
    .din(G7)
  );


  splt
  gG7_spl_
  (
    .dout(G7_spl_0),
    .din(G7_spl_)
  );


  splt
  gG7_spl_0
  (
    .dout(G7_spl_00),
    .din(G7_spl_0)
  );


  splt
  gG7_spl_00
  (
    .dout(G7_spl_000),
    .din(G7_spl_00)
  );


  splt
  gG7_spl_00
  (
    .dout(G7_spl_001),
    .din(G7_spl_00)
  );


  splt
  gG7_spl_0
  (
    .dout(G7_spl_01),
    .din(G7_spl_0)
  );


  splt
  gG7_spl_01
  (
    .dout(G7_spl_010),
    .din(G7_spl_01)
  );


  splt
  gG7_spl_01
  (
    .dout(G7_spl_011),
    .din(G7_spl_01)
  );


  splt
  gG7_spl_
  (
    .dout(G7_spl_1),
    .din(G7_spl_)
  );


  splt
  gG7_spl_1
  (
    .dout(G7_spl_10),
    .din(G7_spl_1)
  );


  splt
  gG7_spl_10
  (
    .dout(G7_spl_100),
    .din(G7_spl_10)
  );


  splt
  gG7_spl_10
  (
    .dout(G7_spl_101),
    .din(G7_spl_10)
  );


  splt
  gG7_spl_1
  (
    .dout(G7_spl_11),
    .din(G7_spl_1)
  );


  splt
  gG7_spl_11
  (
    .dout(G7_spl_110),
    .din(G7_spl_11)
  );


  splt
  gG7_spl_11
  (
    .dout(G7_spl_111),
    .din(G7_spl_11)
  );


  splt
  gG8
  (
    .dout(G8_spl_),
    .din(G8)
  );


  splt
  gG8_spl_
  (
    .dout(G8_spl_0),
    .din(G8_spl_)
  );


  splt
  gG8_spl_0
  (
    .dout(G8_spl_00),
    .din(G8_spl_0)
  );


  splt
  gG8_spl_00
  (
    .dout(G8_spl_000),
    .din(G8_spl_00)
  );


  splt
  gG8_spl_00
  (
    .dout(G8_spl_001),
    .din(G8_spl_00)
  );


  splt
  gG8_spl_0
  (
    .dout(G8_spl_01),
    .din(G8_spl_0)
  );


  splt
  gG8_spl_01
  (
    .dout(G8_spl_010),
    .din(G8_spl_01)
  );


  splt
  gG8_spl_01
  (
    .dout(G8_spl_011),
    .din(G8_spl_01)
  );


  splt
  gG8_spl_
  (
    .dout(G8_spl_1),
    .din(G8_spl_)
  );


  splt
  gG8_spl_1
  (
    .dout(G8_spl_10),
    .din(G8_spl_1)
  );


  splt
  gG8_spl_10
  (
    .dout(G8_spl_100),
    .din(G8_spl_10)
  );


  splt
  gG8_spl_10
  (
    .dout(G8_spl_101),
    .din(G8_spl_10)
  );


  splt
  gG8_spl_1
  (
    .dout(G8_spl_11),
    .din(G8_spl_1)
  );


  splt
  gnew_n73_
  (
    .dout(new_n73__spl_),
    .din(new_n73_)
  );


  splt
  gG9
  (
    .dout(G9_spl_),
    .din(G9)
  );


  splt
  gG9_spl_
  (
    .dout(G9_spl_0),
    .din(G9_spl_)
  );


  splt
  gG9_spl_0
  (
    .dout(G9_spl_00),
    .din(G9_spl_0)
  );


  splt
  gG9_spl_00
  (
    .dout(G9_spl_000),
    .din(G9_spl_00)
  );


  splt
  gG9_spl_00
  (
    .dout(G9_spl_001),
    .din(G9_spl_00)
  );


  splt
  gG9_spl_0
  (
    .dout(G9_spl_01),
    .din(G9_spl_0)
  );


  splt
  gG9_spl_01
  (
    .dout(G9_spl_010),
    .din(G9_spl_01)
  );


  splt
  gG9_spl_01
  (
    .dout(G9_spl_011),
    .din(G9_spl_01)
  );


  splt
  gG9_spl_
  (
    .dout(G9_spl_1),
    .din(G9_spl_)
  );


  splt
  gG9_spl_1
  (
    .dout(G9_spl_10),
    .din(G9_spl_1)
  );


  splt
  gG9_spl_10
  (
    .dout(G9_spl_100),
    .din(G9_spl_10)
  );


  splt
  gG9_spl_10
  (
    .dout(G9_spl_101),
    .din(G9_spl_10)
  );


  splt
  gG9_spl_1
  (
    .dout(G9_spl_11),
    .din(G9_spl_1)
  );


  splt
  gG9_spl_11
  (
    .dout(G9_spl_110),
    .din(G9_spl_11)
  );


  splt
  gnew_n74_
  (
    .dout(new_n74__spl_),
    .din(new_n74_)
  );


  splt
  gG10
  (
    .dout(G10_spl_),
    .din(G10)
  );


  splt
  gG10_spl_
  (
    .dout(G10_spl_0),
    .din(G10_spl_)
  );


  splt
  gG10_spl_0
  (
    .dout(G10_spl_00),
    .din(G10_spl_0)
  );


  splt
  gG10_spl_00
  (
    .dout(G10_spl_000),
    .din(G10_spl_00)
  );


  splt
  gG10_spl_00
  (
    .dout(G10_spl_001),
    .din(G10_spl_00)
  );


  splt
  gG10_spl_0
  (
    .dout(G10_spl_01),
    .din(G10_spl_0)
  );


  splt
  gG10_spl_01
  (
    .dout(G10_spl_010),
    .din(G10_spl_01)
  );


  splt
  gG10_spl_01
  (
    .dout(G10_spl_011),
    .din(G10_spl_01)
  );


  splt
  gG10_spl_
  (
    .dout(G10_spl_1),
    .din(G10_spl_)
  );


  splt
  gG10_spl_1
  (
    .dout(G10_spl_10),
    .din(G10_spl_1)
  );


  splt
  gG10_spl_10
  (
    .dout(G10_spl_100),
    .din(G10_spl_10)
  );


  splt
  gG10_spl_10
  (
    .dout(G10_spl_101),
    .din(G10_spl_10)
  );


  splt
  gG10_spl_1
  (
    .dout(G10_spl_11),
    .din(G10_spl_1)
  );


  splt
  gG10_spl_11
  (
    .dout(G10_spl_110),
    .din(G10_spl_11)
  );


  splt
  gG12
  (
    .dout(G12_spl_),
    .din(G12)
  );


  splt
  gG12_spl_
  (
    .dout(G12_spl_0),
    .din(G12_spl_)
  );


  splt
  gG12_spl_0
  (
    .dout(G12_spl_00),
    .din(G12_spl_0)
  );


  splt
  gG12_spl_00
  (
    .dout(G12_spl_000),
    .din(G12_spl_00)
  );


  splt
  gG12_spl_00
  (
    .dout(G12_spl_001),
    .din(G12_spl_00)
  );


  splt
  gG12_spl_0
  (
    .dout(G12_spl_01),
    .din(G12_spl_0)
  );


  splt
  gG12_spl_01
  (
    .dout(G12_spl_010),
    .din(G12_spl_01)
  );


  splt
  gG12_spl_01
  (
    .dout(G12_spl_011),
    .din(G12_spl_01)
  );


  splt
  gG12_spl_
  (
    .dout(G12_spl_1),
    .din(G12_spl_)
  );


  splt
  gG12_spl_1
  (
    .dout(G12_spl_10),
    .din(G12_spl_1)
  );


  splt
  gG12_spl_10
  (
    .dout(G12_spl_100),
    .din(G12_spl_10)
  );


  splt
  gG12_spl_10
  (
    .dout(G12_spl_101),
    .din(G12_spl_10)
  );


  splt
  gG12_spl_1
  (
    .dout(G12_spl_11),
    .din(G12_spl_1)
  );


  splt
  gG13
  (
    .dout(G13_spl_),
    .din(G13)
  );


  splt
  gG13_spl_
  (
    .dout(G13_spl_0),
    .din(G13_spl_)
  );


  splt
  gG13_spl_0
  (
    .dout(G13_spl_00),
    .din(G13_spl_0)
  );


  splt
  gG13_spl_00
  (
    .dout(G13_spl_000),
    .din(G13_spl_00)
  );


  splt
  gG13_spl_00
  (
    .dout(G13_spl_001),
    .din(G13_spl_00)
  );


  splt
  gG13_spl_0
  (
    .dout(G13_spl_01),
    .din(G13_spl_0)
  );


  splt
  gG13_spl_01
  (
    .dout(G13_spl_010),
    .din(G13_spl_01)
  );


  splt
  gG13_spl_01
  (
    .dout(G13_spl_011),
    .din(G13_spl_01)
  );


  splt
  gG13_spl_
  (
    .dout(G13_spl_1),
    .din(G13_spl_)
  );


  splt
  gG13_spl_1
  (
    .dout(G13_spl_10),
    .din(G13_spl_1)
  );


  splt
  gG13_spl_10
  (
    .dout(G13_spl_100),
    .din(G13_spl_10)
  );


  splt
  gG13_spl_10
  (
    .dout(G13_spl_101),
    .din(G13_spl_10)
  );


  splt
  gG13_spl_1
  (
    .dout(G13_spl_11),
    .din(G13_spl_1)
  );


  splt
  gG13_spl_11
  (
    .dout(G13_spl_110),
    .din(G13_spl_11)
  );


  splt
  gnew_n76_
  (
    .dout(new_n76__spl_),
    .din(new_n76_)
  );


  splt
  gG11
  (
    .dout(G11_spl_),
    .din(G11)
  );


  splt
  gG11_spl_
  (
    .dout(G11_spl_0),
    .din(G11_spl_)
  );


  splt
  gG11_spl_0
  (
    .dout(G11_spl_00),
    .din(G11_spl_0)
  );


  splt
  gG11_spl_00
  (
    .dout(G11_spl_000),
    .din(G11_spl_00)
  );


  splt
  gG11_spl_00
  (
    .dout(G11_spl_001),
    .din(G11_spl_00)
  );


  splt
  gG11_spl_0
  (
    .dout(G11_spl_01),
    .din(G11_spl_0)
  );


  splt
  gG11_spl_01
  (
    .dout(G11_spl_010),
    .din(G11_spl_01)
  );


  splt
  gG11_spl_01
  (
    .dout(G11_spl_011),
    .din(G11_spl_01)
  );


  splt
  gG11_spl_
  (
    .dout(G11_spl_1),
    .din(G11_spl_)
  );


  splt
  gG11_spl_1
  (
    .dout(G11_spl_10),
    .din(G11_spl_1)
  );


  splt
  gG11_spl_10
  (
    .dout(G11_spl_100),
    .din(G11_spl_10)
  );


  splt
  gG11_spl_10
  (
    .dout(G11_spl_101),
    .din(G11_spl_10)
  );


  splt
  gG11_spl_1
  (
    .dout(G11_spl_11),
    .din(G11_spl_1)
  );


  splt
  gG1
  (
    .dout(G1_spl_),
    .din(G1)
  );


  splt
  gG1_spl_
  (
    .dout(G1_spl_0),
    .din(G1_spl_)
  );


  splt
  gG1_spl_0
  (
    .dout(G1_spl_00),
    .din(G1_spl_0)
  );


  splt
  gG1_spl_00
  (
    .dout(G1_spl_000),
    .din(G1_spl_00)
  );


  splt
  gG1_spl_00
  (
    .dout(G1_spl_001),
    .din(G1_spl_00)
  );


  splt
  gG1_spl_0
  (
    .dout(G1_spl_01),
    .din(G1_spl_0)
  );


  splt
  gG1_spl_01
  (
    .dout(G1_spl_010),
    .din(G1_spl_01)
  );


  splt
  gG1_spl_
  (
    .dout(G1_spl_1),
    .din(G1_spl_)
  );


  splt
  gG1_spl_1
  (
    .dout(G1_spl_10),
    .din(G1_spl_1)
  );


  splt
  gG1_spl_1
  (
    .dout(G1_spl_11),
    .din(G1_spl_1)
  );


  splt
  gG3
  (
    .dout(G3_spl_),
    .din(G3)
  );


  splt
  gG3_spl_
  (
    .dout(G3_spl_0),
    .din(G3_spl_)
  );


  splt
  gG3_spl_0
  (
    .dout(G3_spl_00),
    .din(G3_spl_0)
  );


  splt
  gG3_spl_00
  (
    .dout(G3_spl_000),
    .din(G3_spl_00)
  );


  splt
  gG3_spl_000
  (
    .dout(G3_spl_0000),
    .din(G3_spl_000)
  );


  splt
  gG3_spl_000
  (
    .dout(G3_spl_0001),
    .din(G3_spl_000)
  );


  splt
  gG3_spl_00
  (
    .dout(G3_spl_001),
    .din(G3_spl_00)
  );


  splt
  gG3_spl_001
  (
    .dout(G3_spl_0010),
    .din(G3_spl_001)
  );


  splt
  gG3_spl_001
  (
    .dout(G3_spl_0011),
    .din(G3_spl_001)
  );


  splt
  gG3_spl_0
  (
    .dout(G3_spl_01),
    .din(G3_spl_0)
  );


  splt
  gG3_spl_01
  (
    .dout(G3_spl_010),
    .din(G3_spl_01)
  );


  splt
  gG3_spl_010
  (
    .dout(G3_spl_0100),
    .din(G3_spl_010)
  );


  splt
  gG3_spl_01
  (
    .dout(G3_spl_011),
    .din(G3_spl_01)
  );


  splt
  gG3_spl_
  (
    .dout(G3_spl_1),
    .din(G3_spl_)
  );


  splt
  gG3_spl_1
  (
    .dout(G3_spl_10),
    .din(G3_spl_1)
  );


  splt
  gG3_spl_10
  (
    .dout(G3_spl_100),
    .din(G3_spl_10)
  );


  splt
  gG3_spl_10
  (
    .dout(G3_spl_101),
    .din(G3_spl_10)
  );


  splt
  gG3_spl_1
  (
    .dout(G3_spl_11),
    .din(G3_spl_1)
  );


  splt
  gG3_spl_11
  (
    .dout(G3_spl_110),
    .din(G3_spl_11)
  );


  splt
  gG3_spl_11
  (
    .dout(G3_spl_111),
    .din(G3_spl_11)
  );


  splt
  gG34
  (
    .dout(G34_spl_),
    .din(G34)
  );


  splt
  gG34_spl_
  (
    .dout(G34_spl_0),
    .din(G34_spl_)
  );


  splt
  gG34_spl_0
  (
    .dout(G34_spl_00),
    .din(G34_spl_0)
  );


  splt
  gG34_spl_0
  (
    .dout(G34_spl_01),
    .din(G34_spl_0)
  );


  splt
  gG34_spl_
  (
    .dout(G34_spl_1),
    .din(G34_spl_)
  );


  splt
  gG34_spl_1
  (
    .dout(G34_spl_10),
    .din(G34_spl_1)
  );


  splt
  gG32
  (
    .dout(G32_spl_),
    .din(G32)
  );


  splt
  gG32_spl_
  (
    .dout(G32_spl_0),
    .din(G32_spl_)
  );


  splt
  gG32_spl_0
  (
    .dout(G32_spl_00),
    .din(G32_spl_0)
  );


  splt
  gG32_spl_0
  (
    .dout(G32_spl_01),
    .din(G32_spl_0)
  );


  splt
  gG32_spl_
  (
    .dout(G32_spl_1),
    .din(G32_spl_)
  );


  splt
  gG30
  (
    .dout(G30_spl_),
    .din(G30)
  );


  splt
  gG30_spl_
  (
    .dout(G30_spl_0),
    .din(G30_spl_)
  );


  splt
  gG30_spl_0
  (
    .dout(G30_spl_00),
    .din(G30_spl_0)
  );


  splt
  gG30_spl_0
  (
    .dout(G30_spl_01),
    .din(G30_spl_0)
  );


  splt
  gG30_spl_
  (
    .dout(G30_spl_1),
    .din(G30_spl_)
  );


  splt
  gG33
  (
    .dout(G33_spl_),
    .din(G33)
  );


  splt
  gG33_spl_
  (
    .dout(G33_spl_0),
    .din(G33_spl_)
  );


  splt
  gG33_spl_0
  (
    .dout(G33_spl_00),
    .din(G33_spl_0)
  );


  splt
  gG33_spl_0
  (
    .dout(G33_spl_01),
    .din(G33_spl_0)
  );


  splt
  gG33_spl_
  (
    .dout(G33_spl_1),
    .din(G33_spl_)
  );


  splt
  gG14
  (
    .dout(G14_spl_),
    .din(G14)
  );


  splt
  gG14_spl_
  (
    .dout(G14_spl_0),
    .din(G14_spl_)
  );


  splt
  gG14_spl_0
  (
    .dout(G14_spl_00),
    .din(G14_spl_0)
  );


  splt
  gG14_spl_00
  (
    .dout(G14_spl_000),
    .din(G14_spl_00)
  );


  splt
  gG14_spl_00
  (
    .dout(G14_spl_001),
    .din(G14_spl_00)
  );


  splt
  gG14_spl_0
  (
    .dout(G14_spl_01),
    .din(G14_spl_0)
  );


  splt
  gG14_spl_01
  (
    .dout(G14_spl_010),
    .din(G14_spl_01)
  );


  splt
  gG14_spl_01
  (
    .dout(G14_spl_011),
    .din(G14_spl_01)
  );


  splt
  gG14_spl_
  (
    .dout(G14_spl_1),
    .din(G14_spl_)
  );


  splt
  gG14_spl_1
  (
    .dout(G14_spl_10),
    .din(G14_spl_1)
  );


  splt
  gG14_spl_10
  (
    .dout(G14_spl_100),
    .din(G14_spl_10)
  );


  splt
  gG14_spl_10
  (
    .dout(G14_spl_101),
    .din(G14_spl_10)
  );


  splt
  gG14_spl_1
  (
    .dout(G14_spl_11),
    .din(G14_spl_1)
  );


  splt
  gG14_spl_11
  (
    .dout(G14_spl_110),
    .din(G14_spl_11)
  );


  splt
  gG14_spl_11
  (
    .dout(G14_spl_111),
    .din(G14_spl_11)
  );


  splt
  gG37
  (
    .dout(G37_spl_),
    .din(G37)
  );


  splt
  gG37_spl_
  (
    .dout(G37_spl_0),
    .din(G37_spl_)
  );


  splt
  gG37_spl_
  (
    .dout(G37_spl_1),
    .din(G37_spl_)
  );


  splt
  gG31
  (
    .dout(G31_spl_),
    .din(G31)
  );


  splt
  gG31_spl_
  (
    .dout(G31_spl_0),
    .din(G31_spl_)
  );


  splt
  gG31_spl_0
  (
    .dout(G31_spl_00),
    .din(G31_spl_0)
  );


  splt
  gG31_spl_0
  (
    .dout(G31_spl_01),
    .din(G31_spl_0)
  );


  splt
  gG31_spl_
  (
    .dout(G31_spl_1),
    .din(G31_spl_)
  );


  splt
  gG35
  (
    .dout(G35_spl_),
    .din(G35)
  );


  splt
  gG35_spl_
  (
    .dout(G35_spl_0),
    .din(G35_spl_)
  );


  splt
  gG35_spl_0
  (
    .dout(G35_spl_00),
    .din(G35_spl_0)
  );


  splt
  gG35_spl_0
  (
    .dout(G35_spl_01),
    .din(G35_spl_0)
  );


  splt
  gG35_spl_
  (
    .dout(G35_spl_1),
    .din(G35_spl_)
  );


  splt
  gG35_spl_1
  (
    .dout(G35_spl_10),
    .din(G35_spl_1)
  );


  splt
  gG36
  (
    .dout(G36_spl_),
    .din(G36)
  );


  splt
  gG36_spl_
  (
    .dout(G36_spl_0),
    .din(G36_spl_)
  );


  splt
  gG36_spl_0
  (
    .dout(G36_spl_00),
    .din(G36_spl_0)
  );


  splt
  gG36_spl_0
  (
    .dout(G36_spl_01),
    .din(G36_spl_0)
  );


  splt
  gG36_spl_
  (
    .dout(G36_spl_1),
    .din(G36_spl_)
  );


  splt
  gG2
  (
    .dout(G2_spl_),
    .din(G2)
  );


  splt
  gG2_spl_
  (
    .dout(G2_spl_0),
    .din(G2_spl_)
  );


  splt
  gG2_spl_0
  (
    .dout(G2_spl_00),
    .din(G2_spl_0)
  );


  splt
  gG2_spl_
  (
    .dout(G2_spl_1),
    .din(G2_spl_)
  );


  splt
  gnew_n95_
  (
    .dout(new_n95__spl_),
    .din(new_n95_)
  );


  splt
  gnew_n95__spl_
  (
    .dout(new_n95__spl_0),
    .din(new_n95__spl_)
  );


  splt
  gnew_n97_
  (
    .dout(new_n97__spl_),
    .din(new_n97_)
  );


  splt
  gnew_n96_
  (
    .dout(new_n96__spl_),
    .din(new_n96_)
  );


  splt
  gnew_n96__spl_
  (
    .dout(new_n96__spl_0),
    .din(new_n96__spl_)
  );


  splt
  gnew_n98_
  (
    .dout(new_n98__spl_),
    .din(new_n98_)
  );


  splt
  gnew_n98__spl_
  (
    .dout(new_n98__spl_0),
    .din(new_n98__spl_)
  );


  splt
  gnew_n100_
  (
    .dout(new_n100__spl_),
    .din(new_n100_)
  );


  splt
  gnew_n100__spl_
  (
    .dout(new_n100__spl_0),
    .din(new_n100__spl_)
  );


  splt
  gnew_n101_
  (
    .dout(new_n101__spl_),
    .din(new_n101_)
  );


  splt
  gnew_n101__spl_
  (
    .dout(new_n101__spl_0),
    .din(new_n101__spl_)
  );


  splt
  gnew_n101__spl_
  (
    .dout(new_n101__spl_1),
    .din(new_n101__spl_)
  );


  splt
  gnew_n109_
  (
    .dout(new_n109__spl_),
    .din(new_n109_)
  );


  splt
  gnew_n112_
  (
    .dout(new_n112__spl_),
    .din(new_n112_)
  );


  splt
  gnew_n118_
  (
    .dout(new_n118__spl_),
    .din(new_n118_)
  );


  splt
  gnew_n121_
  (
    .dout(new_n121__spl_),
    .din(new_n121_)
  );


  splt
  gnew_n115_
  (
    .dout(new_n115__spl_),
    .din(new_n115_)
  );


  splt
  gnew_n124_
  (
    .dout(new_n124__spl_),
    .din(new_n124_)
  );


  splt
  gnew_n128_
  (
    .dout(new_n128__spl_),
    .din(new_n128_)
  );


  splt
  gnew_n130_
  (
    .dout(new_n130__spl_),
    .din(new_n130_)
  );


  splt
  gnew_n133_
  (
    .dout(new_n133__spl_),
    .din(new_n133_)
  );


  splt
  gnew_n138_
  (
    .dout(new_n138__spl_),
    .din(new_n138_)
  );


  splt
  gnew_n141_
  (
    .dout(new_n141__spl_),
    .din(new_n141_)
  );


  splt
  gnew_n136_
  (
    .dout(new_n136__spl_),
    .din(new_n136_)
  );


  splt
  gnew_n144_
  (
    .dout(new_n144__spl_),
    .din(new_n144_)
  );


  splt
  gnew_n144__spl_
  (
    .dout(new_n144__spl_0),
    .din(new_n144__spl_)
  );


  splt
  gG4
  (
    .dout(G4_spl_),
    .din(G4)
  );


  splt
  gG4_spl_
  (
    .dout(G4_spl_0),
    .din(G4_spl_)
  );


  splt
  gG4_spl_0
  (
    .dout(G4_spl_00),
    .din(G4_spl_0)
  );


  splt
  gG4_spl_00
  (
    .dout(G4_spl_000),
    .din(G4_spl_00)
  );


  splt
  gG4_spl_000
  (
    .dout(G4_spl_0000),
    .din(G4_spl_000)
  );


  splt
  gG4_spl_0000
  (
    .dout(G4_spl_00000),
    .din(G4_spl_0000)
  );


  splt
  gG4_spl_0000
  (
    .dout(G4_spl_00001),
    .din(G4_spl_0000)
  );


  splt
  gG4_spl_000
  (
    .dout(G4_spl_0001),
    .din(G4_spl_000)
  );


  splt
  gG4_spl_0001
  (
    .dout(G4_spl_00010),
    .din(G4_spl_0001)
  );


  splt
  gG4_spl_0001
  (
    .dout(G4_spl_00011),
    .din(G4_spl_0001)
  );


  splt
  gG4_spl_00
  (
    .dout(G4_spl_001),
    .din(G4_spl_00)
  );


  splt
  gG4_spl_001
  (
    .dout(G4_spl_0010),
    .din(G4_spl_001)
  );


  splt
  gG4_spl_0010
  (
    .dout(G4_spl_00100),
    .din(G4_spl_0010)
  );


  splt
  gG4_spl_0010
  (
    .dout(G4_spl_00101),
    .din(G4_spl_0010)
  );


  splt
  gG4_spl_001
  (
    .dout(G4_spl_0011),
    .din(G4_spl_001)
  );


  splt
  gG4_spl_0011
  (
    .dout(G4_spl_00110),
    .din(G4_spl_0011)
  );


  splt
  gG4_spl_0
  (
    .dout(G4_spl_01),
    .din(G4_spl_0)
  );


  splt
  gG4_spl_01
  (
    .dout(G4_spl_010),
    .din(G4_spl_01)
  );


  splt
  gG4_spl_010
  (
    .dout(G4_spl_0100),
    .din(G4_spl_010)
  );


  splt
  gG4_spl_010
  (
    .dout(G4_spl_0101),
    .din(G4_spl_010)
  );


  splt
  gG4_spl_01
  (
    .dout(G4_spl_011),
    .din(G4_spl_01)
  );


  splt
  gG4_spl_011
  (
    .dout(G4_spl_0110),
    .din(G4_spl_011)
  );


  splt
  gG4_spl_011
  (
    .dout(G4_spl_0111),
    .din(G4_spl_011)
  );


  splt
  gG4_spl_
  (
    .dout(G4_spl_1),
    .din(G4_spl_)
  );


  splt
  gG4_spl_1
  (
    .dout(G4_spl_10),
    .din(G4_spl_1)
  );


  splt
  gG4_spl_10
  (
    .dout(G4_spl_100),
    .din(G4_spl_10)
  );


  splt
  gG4_spl_100
  (
    .dout(G4_spl_1000),
    .din(G4_spl_100)
  );


  splt
  gG4_spl_100
  (
    .dout(G4_spl_1001),
    .din(G4_spl_100)
  );


  splt
  gG4_spl_10
  (
    .dout(G4_spl_101),
    .din(G4_spl_10)
  );


  splt
  gG4_spl_101
  (
    .dout(G4_spl_1010),
    .din(G4_spl_101)
  );


  splt
  gG4_spl_101
  (
    .dout(G4_spl_1011),
    .din(G4_spl_101)
  );


  splt
  gG4_spl_1
  (
    .dout(G4_spl_11),
    .din(G4_spl_1)
  );


  splt
  gG4_spl_11
  (
    .dout(G4_spl_110),
    .din(G4_spl_11)
  );


  splt
  gG4_spl_110
  (
    .dout(G4_spl_1100),
    .din(G4_spl_110)
  );


  splt
  gG4_spl_110
  (
    .dout(G4_spl_1101),
    .din(G4_spl_110)
  );


  splt
  gG4_spl_11
  (
    .dout(G4_spl_111),
    .din(G4_spl_11)
  );


  splt
  gG4_spl_111
  (
    .dout(G4_spl_1110),
    .din(G4_spl_111)
  );


  splt
  gG4_spl_111
  (
    .dout(G4_spl_1111),
    .din(G4_spl_111)
  );


  splt
  gnew_n148_
  (
    .dout(new_n148__spl_),
    .din(new_n148_)
  );


  splt
  gnew_n154_
  (
    .dout(new_n154__spl_),
    .din(new_n154_)
  );


  splt
  gnew_n154__spl_
  (
    .dout(new_n154__spl_0),
    .din(new_n154__spl_)
  );


  splt
  gnew_n154__spl_
  (
    .dout(new_n154__spl_1),
    .din(new_n154__spl_)
  );


  splt
  gG39
  (
    .dout(G39_spl_),
    .din(G39)
  );


  splt
  gG39_spl_
  (
    .dout(G39_spl_0),
    .din(G39_spl_)
  );


  splt
  gG39_spl_0
  (
    .dout(G39_spl_00),
    .din(G39_spl_0)
  );


  splt
  gG39_spl_00
  (
    .dout(G39_spl_000),
    .din(G39_spl_00)
  );


  splt
  gG39_spl_0
  (
    .dout(G39_spl_01),
    .din(G39_spl_0)
  );


  splt
  gG39_spl_
  (
    .dout(G39_spl_1),
    .din(G39_spl_)
  );


  splt
  gG39_spl_1
  (
    .dout(G39_spl_10),
    .din(G39_spl_1)
  );


  splt
  gG39_spl_1
  (
    .dout(G39_spl_11),
    .din(G39_spl_1)
  );


  splt
  gnew_n153_
  (
    .dout(new_n153__spl_),
    .din(new_n153_)
  );


  splt
  gnew_n153__spl_
  (
    .dout(new_n153__spl_0),
    .din(new_n153__spl_)
  );


  splt
  gnew_n153__spl_
  (
    .dout(new_n153__spl_1),
    .din(new_n153__spl_)
  );


  splt
  gnew_n151_
  (
    .dout(new_n151__spl_),
    .din(new_n151_)
  );


  splt
  gnew_n151__spl_
  (
    .dout(new_n151__spl_0),
    .din(new_n151__spl_)
  );


  splt
  gnew_n151__spl_0
  (
    .dout(new_n151__spl_00),
    .din(new_n151__spl_0)
  );


  splt
  gnew_n151__spl_00
  (
    .dout(new_n151__spl_000),
    .din(new_n151__spl_00)
  );


  splt
  gnew_n151__spl_00
  (
    .dout(new_n151__spl_001),
    .din(new_n151__spl_00)
  );


  splt
  gnew_n151__spl_0
  (
    .dout(new_n151__spl_01),
    .din(new_n151__spl_0)
  );


  splt
  gnew_n151__spl_
  (
    .dout(new_n151__spl_1),
    .din(new_n151__spl_)
  );


  splt
  gnew_n151__spl_1
  (
    .dout(new_n151__spl_10),
    .din(new_n151__spl_1)
  );


  splt
  gnew_n151__spl_1
  (
    .dout(new_n151__spl_11),
    .din(new_n151__spl_1)
  );


  splt
  gnew_n160_
  (
    .dout(new_n160__spl_),
    .din(new_n160_)
  );


  splt
  gnew_n160__spl_
  (
    .dout(new_n160__spl_0),
    .din(new_n160__spl_)
  );


  splt
  gnew_n160__spl_0
  (
    .dout(new_n160__spl_00),
    .din(new_n160__spl_0)
  );


  splt
  gnew_n160__spl_0
  (
    .dout(new_n160__spl_01),
    .din(new_n160__spl_0)
  );


  splt
  gnew_n160__spl_
  (
    .dout(new_n160__spl_1),
    .din(new_n160__spl_)
  );


  splt
  gnew_n160__spl_1
  (
    .dout(new_n160__spl_10),
    .din(new_n160__spl_1)
  );


  splt
  gnew_n160__spl_1
  (
    .dout(new_n160__spl_11),
    .din(new_n160__spl_1)
  );


  splt
  gnew_n162_
  (
    .dout(new_n162__spl_),
    .din(new_n162_)
  );


  splt
  gnew_n165_
  (
    .dout(new_n165__spl_),
    .din(new_n165_)
  );


  splt
  gnew_n165__spl_
  (
    .dout(new_n165__spl_0),
    .din(new_n165__spl_)
  );


  splt
  gnew_n164_
  (
    .dout(new_n164__spl_),
    .din(new_n164_)
  );


  splt
  gnew_n164__spl_
  (
    .dout(new_n164__spl_0),
    .din(new_n164__spl_)
  );


  splt
  gnew_n164__spl_
  (
    .dout(new_n164__spl_1),
    .din(new_n164__spl_)
  );


  splt
  gG5
  (
    .dout(G5_spl_),
    .din(G5)
  );


  splt
  gG5_spl_
  (
    .dout(G5_spl_0),
    .din(G5_spl_)
  );


  splt
  gG5_spl_0
  (
    .dout(G5_spl_00),
    .din(G5_spl_0)
  );


  splt
  gG5_spl_0
  (
    .dout(G5_spl_01),
    .din(G5_spl_0)
  );


  splt
  gG5_spl_
  (
    .dout(G5_spl_1),
    .din(G5_spl_)
  );


  splt
  gnew_n170_
  (
    .dout(new_n170__spl_),
    .din(new_n170_)
  );


  splt
  gnew_n171_
  (
    .dout(new_n171__spl_),
    .din(new_n171_)
  );


  splt
  gnew_n171__spl_
  (
    .dout(new_n171__spl_0),
    .din(new_n171__spl_)
  );


  splt
  gnew_n171__spl_0
  (
    .dout(new_n171__spl_00),
    .din(new_n171__spl_0)
  );


  splt
  gnew_n171__spl_00
  (
    .dout(new_n171__spl_000),
    .din(new_n171__spl_00)
  );


  splt
  gnew_n171__spl_0
  (
    .dout(new_n171__spl_01),
    .din(new_n171__spl_0)
  );


  splt
  gnew_n171__spl_
  (
    .dout(new_n171__spl_1),
    .din(new_n171__spl_)
  );


  splt
  gnew_n171__spl_1
  (
    .dout(new_n171__spl_10),
    .din(new_n171__spl_1)
  );


  splt
  gnew_n171__spl_1
  (
    .dout(new_n171__spl_11),
    .din(new_n171__spl_1)
  );


  splt
  gG6
  (
    .dout(G6_spl_),
    .din(G6)
  );


  splt
  gG6_spl_
  (
    .dout(G6_spl_0),
    .din(G6_spl_)
  );


  splt
  gG6_spl_0
  (
    .dout(G6_spl_00),
    .din(G6_spl_0)
  );


  splt
  gG6_spl_
  (
    .dout(G6_spl_1),
    .din(G6_spl_)
  );


  splt
  gnew_n173_
  (
    .dout(new_n173__spl_),
    .din(new_n173_)
  );


  splt
  gnew_n173__spl_
  (
    .dout(new_n173__spl_0),
    .din(new_n173__spl_)
  );


  splt
  gnew_n172_
  (
    .dout(new_n172__spl_),
    .din(new_n172_)
  );


  splt
  gnew_n172__spl_
  (
    .dout(new_n172__spl_0),
    .din(new_n172__spl_)
  );


  splt
  gnew_n174_
  (
    .dout(new_n174__spl_),
    .din(new_n174_)
  );


  splt
  gnew_n174__spl_
  (
    .dout(new_n174__spl_0),
    .din(new_n174__spl_)
  );


  splt
  gnew_n174__spl_
  (
    .dout(new_n174__spl_1),
    .din(new_n174__spl_)
  );


  splt
  gG41
  (
    .dout(G41_spl_),
    .din(G41)
  );


  splt
  gG41_spl_
  (
    .dout(G41_spl_0),
    .din(G41_spl_)
  );


  splt
  gG41_spl_0
  (
    .dout(G41_spl_00),
    .din(G41_spl_0)
  );


  splt
  gG41_spl_0
  (
    .dout(G41_spl_01),
    .din(G41_spl_0)
  );


  splt
  gG41_spl_
  (
    .dout(G41_spl_1),
    .din(G41_spl_)
  );


  splt
  gG41_spl_1
  (
    .dout(G41_spl_10),
    .din(G41_spl_1)
  );


  splt
  gnew_n180_
  (
    .dout(new_n180__spl_),
    .din(new_n180_)
  );


  splt
  gnew_n180__spl_
  (
    .dout(new_n180__spl_0),
    .din(new_n180__spl_)
  );


  splt
  gnew_n180__spl_0
  (
    .dout(new_n180__spl_00),
    .din(new_n180__spl_0)
  );


  splt
  gnew_n180__spl_0
  (
    .dout(new_n180__spl_01),
    .din(new_n180__spl_0)
  );


  splt
  gnew_n180__spl_
  (
    .dout(new_n180__spl_1),
    .din(new_n180__spl_)
  );


  splt
  gnew_n180__spl_1
  (
    .dout(new_n180__spl_10),
    .din(new_n180__spl_1)
  );


  splt
  gnew_n180__spl_1
  (
    .dout(new_n180__spl_11),
    .din(new_n180__spl_1)
  );


  splt
  gnew_n175_
  (
    .dout(new_n175__spl_),
    .din(new_n175_)
  );


  splt
  gnew_n175__spl_
  (
    .dout(new_n175__spl_0),
    .din(new_n175__spl_)
  );


  splt
  gG25
  (
    .dout(G25_spl_),
    .din(G25)
  );


  splt
  gG26
  (
    .dout(G26_spl_),
    .din(G26)
  );


  splt
  gG26_spl_
  (
    .dout(G26_spl_0),
    .din(G26_spl_)
  );


  splt
  gnew_n185_
  (
    .dout(new_n185__spl_),
    .din(new_n185_)
  );


  splt
  gnew_n185__spl_
  (
    .dout(new_n185__spl_0),
    .din(new_n185__spl_)
  );


  splt
  gnew_n185__spl_
  (
    .dout(new_n185__spl_1),
    .din(new_n185__spl_)
  );


  splt
  gnew_n186_
  (
    .dout(new_n186__spl_),
    .din(new_n186_)
  );


  splt
  gnew_n186__spl_
  (
    .dout(new_n186__spl_0),
    .din(new_n186__spl_)
  );


  splt
  gnew_n186__spl_0
  (
    .dout(new_n186__spl_00),
    .din(new_n186__spl_0)
  );


  splt
  gnew_n186__spl_00
  (
    .dout(new_n186__spl_000),
    .din(new_n186__spl_00)
  );


  splt
  gnew_n186__spl_0
  (
    .dout(new_n186__spl_01),
    .din(new_n186__spl_0)
  );


  splt
  gnew_n186__spl_
  (
    .dout(new_n186__spl_1),
    .din(new_n186__spl_)
  );


  splt
  gnew_n186__spl_1
  (
    .dout(new_n186__spl_10),
    .din(new_n186__spl_1)
  );


  splt
  gnew_n186__spl_1
  (
    .dout(new_n186__spl_11),
    .din(new_n186__spl_1)
  );


  splt
  gnew_n169_
  (
    .dout(new_n169__spl_),
    .din(new_n169_)
  );


  splt
  gnew_n169__spl_
  (
    .dout(new_n169__spl_0),
    .din(new_n169__spl_)
  );


  splt
  gG23
  (
    .dout(G23_spl_),
    .din(G23)
  );


  splt
  gG24
  (
    .dout(G24_spl_),
    .din(G24)
  );


  splt
  gG24_spl_
  (
    .dout(G24_spl_0),
    .din(G24_spl_)
  );


  splt
  gG24_spl_
  (
    .dout(G24_spl_1),
    .din(G24_spl_)
  );


  splt
  gnew_n189_
  (
    .dout(new_n189__spl_),
    .din(new_n189_)
  );


  splt
  gnew_n189__spl_
  (
    .dout(new_n189__spl_0),
    .din(new_n189__spl_)
  );


  splt
  gnew_n189__spl_0
  (
    .dout(new_n189__spl_00),
    .din(new_n189__spl_0)
  );


  splt
  gnew_n189__spl_0
  (
    .dout(new_n189__spl_01),
    .din(new_n189__spl_0)
  );


  splt
  gnew_n189__spl_
  (
    .dout(new_n189__spl_1),
    .din(new_n189__spl_)
  );


  splt
  gnew_n189__spl_1
  (
    .dout(new_n189__spl_10),
    .din(new_n189__spl_1)
  );


  splt
  gnew_n189__spl_1
  (
    .dout(new_n189__spl_11),
    .din(new_n189__spl_1)
  );


  splt
  gnew_n191_
  (
    .dout(new_n191__spl_),
    .din(new_n191_)
  );


  splt
  gnew_n191__spl_
  (
    .dout(new_n191__spl_0),
    .din(new_n191__spl_)
  );


  splt
  gnew_n197_
  (
    .dout(new_n197__spl_),
    .din(new_n197_)
  );


  splt
  gG40
  (
    .dout(G40_spl_),
    .din(G40)
  );


  splt
  gG40_spl_
  (
    .dout(G40_spl_0),
    .din(G40_spl_)
  );


  splt
  gG40_spl_0
  (
    .dout(G40_spl_00),
    .din(G40_spl_0)
  );


  splt
  gG40_spl_0
  (
    .dout(G40_spl_01),
    .din(G40_spl_0)
  );


  splt
  gG40_spl_
  (
    .dout(G40_spl_1),
    .din(G40_spl_)
  );


  splt
  gG40_spl_1
  (
    .dout(G40_spl_10),
    .din(G40_spl_1)
  );


  splt
  gnew_n210_
  (
    .dout(new_n210__spl_),
    .din(new_n210_)
  );


  splt
  gnew_n210__spl_
  (
    .dout(new_n210__spl_0),
    .din(new_n210__spl_)
  );


  splt
  gnew_n210__spl_
  (
    .dout(new_n210__spl_1),
    .din(new_n210__spl_)
  );


  splt
  gnew_n201_
  (
    .dout(new_n201__spl_),
    .din(new_n201_)
  );


  splt
  gnew_n201__spl_
  (
    .dout(new_n201__spl_0),
    .din(new_n201__spl_)
  );


  splt
  gnew_n214_
  (
    .dout(new_n214__spl_),
    .din(new_n214_)
  );


  splt
  gnew_n214__spl_
  (
    .dout(new_n214__spl_0),
    .din(new_n214__spl_)
  );


  splt
  gnew_n152_
  (
    .dout(new_n152__spl_),
    .din(new_n152_)
  );


  splt
  gnew_n152__spl_
  (
    .dout(new_n152__spl_0),
    .din(new_n152__spl_)
  );


  splt
  gnew_n152__spl_
  (
    .dout(new_n152__spl_1),
    .din(new_n152__spl_)
  );


  splt
  gnew_n236_
  (
    .dout(new_n236__spl_),
    .din(new_n236_)
  );


  splt
  gnew_n236__spl_
  (
    .dout(new_n236__spl_0),
    .din(new_n236__spl_)
  );


  splt
  gnew_n236__spl_
  (
    .dout(new_n236__spl_1),
    .din(new_n236__spl_)
  );


  splt
  gnew_n226_
  (
    .dout(new_n226__spl_),
    .din(new_n226_)
  );


  splt
  gnew_n226__spl_
  (
    .dout(new_n226__spl_0),
    .din(new_n226__spl_)
  );


  splt
  gnew_n240_
  (
    .dout(new_n240__spl_),
    .din(new_n240_)
  );


  splt
  gnew_n155_
  (
    .dout(new_n155__spl_),
    .din(new_n155_)
  );


  splt
  gnew_n155__spl_
  (
    .dout(new_n155__spl_0),
    .din(new_n155__spl_)
  );


  splt
  gnew_n155__spl_
  (
    .dout(new_n155__spl_1),
    .din(new_n155__spl_)
  );


  splt
  gnew_n248_
  (
    .dout(new_n248__spl_),
    .din(new_n248_)
  );


  splt
  gnew_n262_
  (
    .dout(new_n262__spl_),
    .din(new_n262_)
  );


  splt
  gnew_n262__spl_
  (
    .dout(new_n262__spl_0),
    .din(new_n262__spl_)
  );


  splt
  gnew_n262__spl_
  (
    .dout(new_n262__spl_1),
    .din(new_n262__spl_)
  );


  splt
  gnew_n253_
  (
    .dout(new_n253__spl_),
    .din(new_n253_)
  );


  splt
  gnew_n253__spl_
  (
    .dout(new_n253__spl_0),
    .din(new_n253__spl_)
  );


  splt
  gnew_n266_
  (
    .dout(new_n266__spl_),
    .din(new_n266_)
  );


  splt
  gnew_n266__spl_
  (
    .dout(new_n266__spl_0),
    .din(new_n266__spl_)
  );


  splt
  gnew_n241_
  (
    .dout(new_n241__spl_),
    .din(new_n241_)
  );


  splt
  gnew_n241__spl_
  (
    .dout(new_n241__spl_0),
    .din(new_n241__spl_)
  );


  splt
  gnew_n241__spl_
  (
    .dout(new_n241__spl_1),
    .din(new_n241__spl_)
  );


  splt
  gnew_n267_
  (
    .dout(new_n267__spl_),
    .din(new_n267_)
  );


  splt
  gnew_n267__spl_
  (
    .dout(new_n267__spl_0),
    .din(new_n267__spl_)
  );


  splt
  gnew_n215_
  (
    .dout(new_n215__spl_),
    .din(new_n215_)
  );


  splt
  gnew_n215__spl_
  (
    .dout(new_n215__spl_0),
    .din(new_n215__spl_)
  );


  splt
  gnew_n268_
  (
    .dout(new_n268__spl_),
    .din(new_n268_)
  );


  splt
  gnew_n192_
  (
    .dout(new_n192__spl_),
    .din(new_n192_)
  );


  splt
  gnew_n192__spl_
  (
    .dout(new_n192__spl_0),
    .din(new_n192__spl_)
  );


  splt
  gnew_n269_
  (
    .dout(new_n269__spl_),
    .din(new_n269_)
  );


  splt
  gnew_n277_
  (
    .dout(new_n277__spl_),
    .din(new_n277_)
  );


  splt
  gnew_n277__spl_
  (
    .dout(new_n277__spl_0),
    .din(new_n277__spl_)
  );


  splt
  gnew_n277__spl_
  (
    .dout(new_n277__spl_1),
    .din(new_n277__spl_)
  );


  splt
  gnew_n283_
  (
    .dout(new_n283__spl_),
    .din(new_n283_)
  );


  splt
  gnew_n283__spl_
  (
    .dout(new_n283__spl_0),
    .din(new_n283__spl_)
  );


  splt
  gnew_n283__spl_0
  (
    .dout(new_n283__spl_00),
    .din(new_n283__spl_0)
  );


  splt
  gnew_n283__spl_
  (
    .dout(new_n283__spl_1),
    .din(new_n283__spl_)
  );


  splt
  gnew_n284_
  (
    .dout(new_n284__spl_),
    .din(new_n284_)
  );


  splt
  gnew_n284__spl_
  (
    .dout(new_n284__spl_0),
    .din(new_n284__spl_)
  );


  splt
  gnew_n284__spl_
  (
    .dout(new_n284__spl_1),
    .din(new_n284__spl_)
  );


  splt
  gnew_n293_
  (
    .dout(new_n293__spl_),
    .din(new_n293_)
  );


  splt
  gnew_n281_
  (
    .dout(new_n281__spl_),
    .din(new_n281_)
  );


  splt
  gnew_n281__spl_
  (
    .dout(new_n281__spl_0),
    .din(new_n281__spl_)
  );


  splt
  gnew_n297_
  (
    .dout(new_n297__spl_),
    .din(new_n297_)
  );


  splt
  gnew_n297__spl_
  (
    .dout(new_n297__spl_0),
    .din(new_n297__spl_)
  );


  splt
  gnew_n315_
  (
    .dout(new_n315__spl_),
    .din(new_n315_)
  );


  splt
  gnew_n306_
  (
    .dout(new_n306__spl_),
    .din(new_n306_)
  );


  splt
  gnew_n306__spl_
  (
    .dout(new_n306__spl_0),
    .din(new_n306__spl_)
  );


  splt
  gnew_n319_
  (
    .dout(new_n319__spl_),
    .din(new_n319_)
  );


  splt
  gnew_n319__spl_
  (
    .dout(new_n319__spl_0),
    .din(new_n319__spl_)
  );


  splt
  gG21
  (
    .dout(G21_spl_),
    .din(G21)
  );


  splt
  gG21_spl_
  (
    .dout(G21_spl_0),
    .din(G21_spl_)
  );


  splt
  gG21_spl_0
  (
    .dout(G21_spl_00),
    .din(G21_spl_0)
  );


  splt
  gG21_spl_0
  (
    .dout(G21_spl_01),
    .din(G21_spl_0)
  );


  splt
  gG21_spl_
  (
    .dout(G21_spl_1),
    .din(G21_spl_)
  );


  splt
  gG21_spl_1
  (
    .dout(G21_spl_10),
    .din(G21_spl_1)
  );


  splt
  gG21_spl_1
  (
    .dout(G21_spl_11),
    .din(G21_spl_1)
  );


  splt
  gG29
  (
    .dout(G29_spl_),
    .din(G29)
  );


  splt
  gnew_n339_
  (
    .dout(new_n339__spl_),
    .din(new_n339_)
  );


  splt
  gnew_n330_
  (
    .dout(new_n330__spl_),
    .din(new_n330_)
  );


  splt
  gnew_n330__spl_
  (
    .dout(new_n330__spl_0),
    .din(new_n330__spl_)
  );


  splt
  gnew_n343_
  (
    .dout(new_n343__spl_),
    .din(new_n343_)
  );


  splt
  gG22
  (
    .dout(G22_spl_),
    .din(G22)
  );


  splt
  gG22_spl_
  (
    .dout(G22_spl_0),
    .din(G22_spl_)
  );


  splt
  gG22_spl_0
  (
    .dout(G22_spl_00),
    .din(G22_spl_0)
  );


  splt
  gG22_spl_0
  (
    .dout(G22_spl_01),
    .din(G22_spl_0)
  );


  splt
  gG22_spl_
  (
    .dout(G22_spl_1),
    .din(G22_spl_)
  );


  splt
  gG22_spl_1
  (
    .dout(G22_spl_10),
    .din(G22_spl_1)
  );


  splt
  gG22_spl_1
  (
    .dout(G22_spl_11),
    .din(G22_spl_1)
  );


  splt
  gnew_n351_
  (
    .dout(new_n351__spl_),
    .din(new_n351_)
  );


  splt
  gnew_n365_
  (
    .dout(new_n365__spl_),
    .din(new_n365_)
  );


  splt
  gnew_n356_
  (
    .dout(new_n356__spl_),
    .din(new_n356_)
  );


  splt
  gnew_n356__spl_
  (
    .dout(new_n356__spl_0),
    .din(new_n356__spl_)
  );


  splt
  gnew_n369_
  (
    .dout(new_n369__spl_),
    .din(new_n369_)
  );


  splt
  gnew_n369__spl_
  (
    .dout(new_n369__spl_0),
    .din(new_n369__spl_)
  );


  splt
  gnew_n344_
  (
    .dout(new_n344__spl_),
    .din(new_n344_)
  );


  splt
  gnew_n344__spl_
  (
    .dout(new_n344__spl_0),
    .din(new_n344__spl_)
  );


  splt
  gnew_n344__spl_
  (
    .dout(new_n344__spl_1),
    .din(new_n344__spl_)
  );


  splt
  gnew_n370_
  (
    .dout(new_n370__spl_),
    .din(new_n370_)
  );


  splt
  gnew_n370__spl_
  (
    .dout(new_n370__spl_0),
    .din(new_n370__spl_)
  );


  splt
  gnew_n320_
  (
    .dout(new_n320__spl_),
    .din(new_n320_)
  );


  splt
  gnew_n320__spl_
  (
    .dout(new_n320__spl_0),
    .din(new_n320__spl_)
  );


  splt
  gnew_n371_
  (
    .dout(new_n371__spl_),
    .din(new_n371_)
  );


  splt
  gnew_n298_
  (
    .dout(new_n298__spl_),
    .din(new_n298_)
  );


  splt
  gnew_n298__spl_
  (
    .dout(new_n298__spl_0),
    .din(new_n298__spl_)
  );


  splt
  gnew_n372_
  (
    .dout(new_n372__spl_),
    .din(new_n372_)
  );


  splt
  gnew_n270_
  (
    .dout(new_n270__spl_),
    .din(new_n270_)
  );


  splt
  gnew_n373_
  (
    .dout(new_n373__spl_),
    .din(new_n373_)
  );


  splt
  gnew_n373__spl_
  (
    .dout(new_n373__spl_0),
    .din(new_n373__spl_)
  );


  splt
  gnew_n373__spl_
  (
    .dout(new_n373__spl_1),
    .din(new_n373__spl_)
  );


  splt
  gnew_n380_
  (
    .dout(new_n380__spl_),
    .din(new_n380_)
  );


  splt
  gnew_n387_
  (
    .dout(new_n387__spl_),
    .din(new_n387_)
  );


  splt
  gG27
  (
    .dout(G27_spl_),
    .din(G27)
  );


  splt
  gG27_spl_
  (
    .dout(G27_spl_0),
    .din(G27_spl_)
  );


  splt
  gG48
  (
    .dout(G48_spl_),
    .din(G48)
  );


  splt
  gnew_n389_
  (
    .dout(new_n389__spl_),
    .din(new_n389_)
  );


  splt
  gnew_n389__spl_
  (
    .dout(new_n389__spl_0),
    .din(new_n389__spl_)
  );


  splt
  gnew_n389__spl_
  (
    .dout(new_n389__spl_1),
    .din(new_n389__spl_)
  );


  splt
  gnew_n390_
  (
    .dout(new_n390__spl_),
    .din(new_n390_)
  );


  splt
  gnew_n390__spl_
  (
    .dout(new_n390__spl_0),
    .din(new_n390__spl_)
  );


  splt
  gnew_n390__spl_0
  (
    .dout(new_n390__spl_00),
    .din(new_n390__spl_0)
  );


  splt
  gnew_n390__spl_00
  (
    .dout(new_n390__spl_000),
    .din(new_n390__spl_00)
  );


  splt
  gnew_n390__spl_00
  (
    .dout(new_n390__spl_001),
    .din(new_n390__spl_00)
  );


  splt
  gnew_n390__spl_0
  (
    .dout(new_n390__spl_01),
    .din(new_n390__spl_0)
  );


  splt
  gnew_n390__spl_01
  (
    .dout(new_n390__spl_010),
    .din(new_n390__spl_01)
  );


  splt
  gnew_n390__spl_01
  (
    .dout(new_n390__spl_011),
    .din(new_n390__spl_01)
  );


  splt
  gnew_n390__spl_
  (
    .dout(new_n390__spl_1),
    .din(new_n390__spl_)
  );


  splt
  gnew_n390__spl_1
  (
    .dout(new_n390__spl_10),
    .din(new_n390__spl_1)
  );


  splt
  gnew_n390__spl_10
  (
    .dout(new_n390__spl_100),
    .din(new_n390__spl_10)
  );


  splt
  gnew_n390__spl_10
  (
    .dout(new_n390__spl_101),
    .din(new_n390__spl_10)
  );


  splt
  gnew_n390__spl_1
  (
    .dout(new_n390__spl_11),
    .din(new_n390__spl_1)
  );


  splt
  gnew_n391_
  (
    .dout(new_n391__spl_),
    .din(new_n391_)
  );


  splt
  gnew_n395_
  (
    .dout(new_n395__spl_),
    .din(new_n395_)
  );


  splt
  gG47
  (
    .dout(G47_spl_),
    .din(G47)
  );


  splt
  gG47_spl_
  (
    .dout(G47_spl_0),
    .din(G47_spl_)
  );


  splt
  gG47_spl_0
  (
    .dout(G47_spl_00),
    .din(G47_spl_0)
  );


  splt
  gG47_spl_0
  (
    .dout(G47_spl_01),
    .din(G47_spl_0)
  );


  splt
  gG47_spl_
  (
    .dout(G47_spl_1),
    .din(G47_spl_)
  );


  splt
  gG47_spl_1
  (
    .dout(G47_spl_10),
    .din(G47_spl_1)
  );


  splt
  gnew_n398_
  (
    .dout(new_n398__spl_),
    .din(new_n398_)
  );


  splt
  gnew_n398__spl_
  (
    .dout(new_n398__spl_0),
    .din(new_n398__spl_)
  );


  splt
  gnew_n398__spl_
  (
    .dout(new_n398__spl_1),
    .din(new_n398__spl_)
  );


  splt
  gnew_n394_
  (
    .dout(new_n394__spl_),
    .din(new_n394_)
  );


  splt
  gnew_n394__spl_
  (
    .dout(new_n394__spl_0),
    .din(new_n394__spl_)
  );


  splt
  gnew_n394__spl_
  (
    .dout(new_n394__spl_1),
    .din(new_n394__spl_)
  );


  splt
  gnew_n401_
  (
    .dout(new_n401__spl_),
    .din(new_n401_)
  );


  splt
  gnew_n401__spl_
  (
    .dout(new_n401__spl_0),
    .din(new_n401__spl_)
  );


  splt
  gnew_n401__spl_0
  (
    .dout(new_n401__spl_00),
    .din(new_n401__spl_0)
  );


  splt
  gnew_n401__spl_0
  (
    .dout(new_n401__spl_01),
    .din(new_n401__spl_0)
  );


  splt
  gnew_n401__spl_
  (
    .dout(new_n401__spl_1),
    .din(new_n401__spl_)
  );


  splt
  gnew_n401__spl_1
  (
    .dout(new_n401__spl_10),
    .din(new_n401__spl_1)
  );


  splt
  gnew_n401__spl_1
  (
    .dout(new_n401__spl_11),
    .din(new_n401__spl_1)
  );


  splt
  gnew_n403_
  (
    .dout(new_n403__spl_),
    .din(new_n403_)
  );


  splt
  gnew_n403__spl_
  (
    .dout(new_n403__spl_0),
    .din(new_n403__spl_)
  );


  splt
  gnew_n403__spl_0
  (
    .dout(new_n403__spl_00),
    .din(new_n403__spl_0)
  );


  splt
  gnew_n403__spl_0
  (
    .dout(new_n403__spl_01),
    .din(new_n403__spl_0)
  );


  splt
  gnew_n403__spl_
  (
    .dout(new_n403__spl_1),
    .din(new_n403__spl_)
  );


  splt
  gnew_n403__spl_1
  (
    .dout(new_n403__spl_10),
    .din(new_n403__spl_1)
  );


  splt
  gnew_n407_
  (
    .dout(new_n407__spl_),
    .din(new_n407_)
  );


  splt
  gnew_n409_
  (
    .dout(new_n409__spl_),
    .din(new_n409_)
  );


  splt
  gnew_n409__spl_
  (
    .dout(new_n409__spl_0),
    .din(new_n409__spl_)
  );


  splt
  gnew_n409__spl_0
  (
    .dout(new_n409__spl_00),
    .din(new_n409__spl_0)
  );


  splt
  gnew_n409__spl_0
  (
    .dout(new_n409__spl_01),
    .din(new_n409__spl_0)
  );


  splt
  gnew_n409__spl_
  (
    .dout(new_n409__spl_1),
    .din(new_n409__spl_)
  );


  splt
  gnew_n409__spl_1
  (
    .dout(new_n409__spl_10),
    .din(new_n409__spl_1)
  );


  splt
  gnew_n411_
  (
    .dout(new_n411__spl_),
    .din(new_n411_)
  );


  splt
  gnew_n411__spl_
  (
    .dout(new_n411__spl_0),
    .din(new_n411__spl_)
  );


  splt
  gnew_n410_
  (
    .dout(new_n410__spl_),
    .din(new_n410_)
  );


  splt
  gnew_n410__spl_
  (
    .dout(new_n410__spl_0),
    .din(new_n410__spl_)
  );


  splt
  gnew_n410__spl_0
  (
    .dout(new_n410__spl_00),
    .din(new_n410__spl_0)
  );


  splt
  gnew_n410__spl_00
  (
    .dout(new_n410__spl_000),
    .din(new_n410__spl_00)
  );


  splt
  gnew_n410__spl_00
  (
    .dout(new_n410__spl_001),
    .din(new_n410__spl_00)
  );


  splt
  gnew_n410__spl_0
  (
    .dout(new_n410__spl_01),
    .din(new_n410__spl_0)
  );


  splt
  gnew_n410__spl_
  (
    .dout(new_n410__spl_1),
    .din(new_n410__spl_)
  );


  splt
  gnew_n410__spl_1
  (
    .dout(new_n410__spl_10),
    .din(new_n410__spl_1)
  );


  splt
  gnew_n410__spl_1
  (
    .dout(new_n410__spl_11),
    .din(new_n410__spl_1)
  );


  splt
  gnew_n414_
  (
    .dout(new_n414__spl_),
    .din(new_n414_)
  );


  splt
  gnew_n414__spl_
  (
    .dout(new_n414__spl_0),
    .din(new_n414__spl_)
  );


  splt
  gnew_n414__spl_
  (
    .dout(new_n414__spl_1),
    .din(new_n414__spl_)
  );


  splt
  gnew_n418_
  (
    .dout(new_n418__spl_),
    .din(new_n418_)
  );


  splt
  gnew_n417_
  (
    .dout(new_n417__spl_),
    .din(new_n417_)
  );


  splt
  gnew_n417__spl_
  (
    .dout(new_n417__spl_0),
    .din(new_n417__spl_)
  );


  splt
  gnew_n417__spl_0
  (
    .dout(new_n417__spl_00),
    .din(new_n417__spl_0)
  );


  splt
  gnew_n417__spl_00
  (
    .dout(new_n417__spl_000),
    .din(new_n417__spl_00)
  );


  splt
  gnew_n417__spl_0
  (
    .dout(new_n417__spl_01),
    .din(new_n417__spl_0)
  );


  splt
  gnew_n417__spl_
  (
    .dout(new_n417__spl_1),
    .din(new_n417__spl_)
  );


  splt
  gnew_n417__spl_1
  (
    .dout(new_n417__spl_10),
    .din(new_n417__spl_1)
  );


  splt
  gnew_n417__spl_1
  (
    .dout(new_n417__spl_11),
    .din(new_n417__spl_1)
  );


  splt
  gnew_n428_
  (
    .dout(new_n428__spl_),
    .din(new_n428_)
  );


  splt
  gnew_n428__spl_
  (
    .dout(new_n428__spl_0),
    .din(new_n428__spl_)
  );


  splt
  gnew_n427_
  (
    .dout(new_n427__spl_),
    .din(new_n427_)
  );


  splt
  gnew_n427__spl_
  (
    .dout(new_n427__spl_0),
    .din(new_n427__spl_)
  );


  splt
  gnew_n427__spl_
  (
    .dout(new_n427__spl_1),
    .din(new_n427__spl_)
  );


  splt
  gnew_n429_
  (
    .dout(new_n429__spl_),
    .din(new_n429_)
  );


  splt
  gG45
  (
    .dout(G45_spl_),
    .din(G45)
  );


  splt
  gnew_n430_
  (
    .dout(new_n430__spl_),
    .din(new_n430_)
  );


  splt
  gnew_n430__spl_
  (
    .dout(new_n430__spl_0),
    .din(new_n430__spl_)
  );


  splt
  gnew_n430__spl_0
  (
    .dout(new_n430__spl_00),
    .din(new_n430__spl_0)
  );


  splt
  gnew_n430__spl_00
  (
    .dout(new_n430__spl_000),
    .din(new_n430__spl_00)
  );


  splt
  gnew_n430__spl_000
  (
    .dout(new_n430__spl_0000),
    .din(new_n430__spl_000)
  );


  splt
  gnew_n430__spl_00
  (
    .dout(new_n430__spl_001),
    .din(new_n430__spl_00)
  );


  splt
  gnew_n430__spl_0
  (
    .dout(new_n430__spl_01),
    .din(new_n430__spl_0)
  );


  splt
  gnew_n430__spl_01
  (
    .dout(new_n430__spl_010),
    .din(new_n430__spl_01)
  );


  splt
  gnew_n430__spl_01
  (
    .dout(new_n430__spl_011),
    .din(new_n430__spl_01)
  );


  splt
  gnew_n430__spl_
  (
    .dout(new_n430__spl_1),
    .din(new_n430__spl_)
  );


  splt
  gnew_n430__spl_1
  (
    .dout(new_n430__spl_10),
    .din(new_n430__spl_1)
  );


  splt
  gnew_n430__spl_10
  (
    .dout(new_n430__spl_100),
    .din(new_n430__spl_10)
  );


  splt
  gnew_n430__spl_10
  (
    .dout(new_n430__spl_101),
    .din(new_n430__spl_10)
  );


  splt
  gnew_n430__spl_1
  (
    .dout(new_n430__spl_11),
    .din(new_n430__spl_1)
  );


  splt
  gnew_n430__spl_11
  (
    .dout(new_n430__spl_110),
    .din(new_n430__spl_11)
  );


  splt
  gnew_n430__spl_11
  (
    .dout(new_n430__spl_111),
    .din(new_n430__spl_11)
  );


  splt
  gnew_n432_
  (
    .dout(new_n432__spl_),
    .din(new_n432_)
  );


  splt
  gnew_n433_
  (
    .dout(new_n433__spl_),
    .din(new_n433_)
  );


  splt
  gnew_n433__spl_
  (
    .dout(new_n433__spl_0),
    .din(new_n433__spl_)
  );


  splt
  gnew_n433__spl_0
  (
    .dout(new_n433__spl_00),
    .din(new_n433__spl_0)
  );


  splt
  gnew_n433__spl_00
  (
    .dout(new_n433__spl_000),
    .din(new_n433__spl_00)
  );


  splt
  gnew_n433__spl_000
  (
    .dout(new_n433__spl_0000),
    .din(new_n433__spl_000)
  );


  splt
  gnew_n433__spl_000
  (
    .dout(new_n433__spl_0001),
    .din(new_n433__spl_000)
  );


  splt
  gnew_n433__spl_00
  (
    .dout(new_n433__spl_001),
    .din(new_n433__spl_00)
  );


  splt
  gnew_n433__spl_0
  (
    .dout(new_n433__spl_01),
    .din(new_n433__spl_0)
  );


  splt
  gnew_n433__spl_01
  (
    .dout(new_n433__spl_010),
    .din(new_n433__spl_01)
  );


  splt
  gnew_n433__spl_01
  (
    .dout(new_n433__spl_011),
    .din(new_n433__spl_01)
  );


  splt
  gnew_n433__spl_
  (
    .dout(new_n433__spl_1),
    .din(new_n433__spl_)
  );


  splt
  gnew_n433__spl_1
  (
    .dout(new_n433__spl_10),
    .din(new_n433__spl_1)
  );


  splt
  gnew_n433__spl_10
  (
    .dout(new_n433__spl_100),
    .din(new_n433__spl_10)
  );


  splt
  gnew_n433__spl_10
  (
    .dout(new_n433__spl_101),
    .din(new_n433__spl_10)
  );


  splt
  gnew_n433__spl_1
  (
    .dout(new_n433__spl_11),
    .din(new_n433__spl_1)
  );


  splt
  gnew_n433__spl_11
  (
    .dout(new_n433__spl_110),
    .din(new_n433__spl_11)
  );


  splt
  gnew_n433__spl_11
  (
    .dout(new_n433__spl_111),
    .din(new_n433__spl_11)
  );


  splt
  gnew_n435_
  (
    .dout(new_n435__spl_),
    .din(new_n435_)
  );


  splt
  gnew_n435__spl_
  (
    .dout(new_n435__spl_0),
    .din(new_n435__spl_)
  );


  splt
  gnew_n435__spl_0
  (
    .dout(new_n435__spl_00),
    .din(new_n435__spl_0)
  );


  splt
  gnew_n435__spl_00
  (
    .dout(new_n435__spl_000),
    .din(new_n435__spl_00)
  );


  splt
  gnew_n435__spl_00
  (
    .dout(new_n435__spl_001),
    .din(new_n435__spl_00)
  );


  splt
  gnew_n435__spl_0
  (
    .dout(new_n435__spl_01),
    .din(new_n435__spl_0)
  );


  splt
  gnew_n435__spl_01
  (
    .dout(new_n435__spl_010),
    .din(new_n435__spl_01)
  );


  splt
  gnew_n435__spl_01
  (
    .dout(new_n435__spl_011),
    .din(new_n435__spl_01)
  );


  splt
  gnew_n435__spl_
  (
    .dout(new_n435__spl_1),
    .din(new_n435__spl_)
  );


  splt
  gnew_n435__spl_1
  (
    .dout(new_n435__spl_10),
    .din(new_n435__spl_1)
  );


  splt
  gnew_n435__spl_10
  (
    .dout(new_n435__spl_100),
    .din(new_n435__spl_10)
  );


  splt
  gnew_n435__spl_10
  (
    .dout(new_n435__spl_101),
    .din(new_n435__spl_10)
  );


  splt
  gnew_n435__spl_1
  (
    .dout(new_n435__spl_11),
    .din(new_n435__spl_1)
  );


  splt
  gnew_n435__spl_11
  (
    .dout(new_n435__spl_110),
    .din(new_n435__spl_11)
  );


  splt
  gnew_n435__spl_11
  (
    .dout(new_n435__spl_111),
    .din(new_n435__spl_11)
  );


  splt
  gG44
  (
    .dout(G44_spl_),
    .din(G44)
  );


  splt
  gG44_spl_
  (
    .dout(G44_spl_0),
    .din(G44_spl_)
  );


  splt
  gG43
  (
    .dout(G43_spl_),
    .din(G43)
  );


  splt
  gG43_spl_
  (
    .dout(G43_spl_0),
    .din(G43_spl_)
  );


  splt
  gG43_spl_
  (
    .dout(G43_spl_1),
    .din(G43_spl_)
  );


  splt
  gnew_n437_
  (
    .dout(new_n437__spl_),
    .din(new_n437_)
  );


  splt
  gnew_n437__spl_
  (
    .dout(new_n437__spl_0),
    .din(new_n437__spl_)
  );


  splt
  gnew_n437__spl_0
  (
    .dout(new_n437__spl_00),
    .din(new_n437__spl_0)
  );


  splt
  gnew_n437__spl_00
  (
    .dout(new_n437__spl_000),
    .din(new_n437__spl_00)
  );


  splt
  gnew_n437__spl_000
  (
    .dout(new_n437__spl_0000),
    .din(new_n437__spl_000)
  );


  splt
  gnew_n437__spl_00
  (
    .dout(new_n437__spl_001),
    .din(new_n437__spl_00)
  );


  splt
  gnew_n437__spl_0
  (
    .dout(new_n437__spl_01),
    .din(new_n437__spl_0)
  );


  splt
  gnew_n437__spl_01
  (
    .dout(new_n437__spl_010),
    .din(new_n437__spl_01)
  );


  splt
  gnew_n437__spl_01
  (
    .dout(new_n437__spl_011),
    .din(new_n437__spl_01)
  );


  splt
  gnew_n437__spl_
  (
    .dout(new_n437__spl_1),
    .din(new_n437__spl_)
  );


  splt
  gnew_n437__spl_1
  (
    .dout(new_n437__spl_10),
    .din(new_n437__spl_1)
  );


  splt
  gnew_n437__spl_10
  (
    .dout(new_n437__spl_100),
    .din(new_n437__spl_10)
  );


  splt
  gnew_n437__spl_10
  (
    .dout(new_n437__spl_101),
    .din(new_n437__spl_10)
  );


  splt
  gnew_n437__spl_1
  (
    .dout(new_n437__spl_11),
    .din(new_n437__spl_1)
  );


  splt
  gnew_n437__spl_11
  (
    .dout(new_n437__spl_110),
    .din(new_n437__spl_11)
  );


  splt
  gnew_n437__spl_11
  (
    .dout(new_n437__spl_111),
    .din(new_n437__spl_11)
  );


  splt
  gnew_n439_
  (
    .dout(new_n439__spl_),
    .din(new_n439_)
  );


  splt
  gnew_n439__spl_
  (
    .dout(new_n439__spl_0),
    .din(new_n439__spl_)
  );


  splt
  gnew_n439__spl_0
  (
    .dout(new_n439__spl_00),
    .din(new_n439__spl_0)
  );


  splt
  gnew_n439__spl_00
  (
    .dout(new_n439__spl_000),
    .din(new_n439__spl_00)
  );


  splt
  gnew_n439__spl_00
  (
    .dout(new_n439__spl_001),
    .din(new_n439__spl_00)
  );


  splt
  gnew_n439__spl_0
  (
    .dout(new_n439__spl_01),
    .din(new_n439__spl_0)
  );


  splt
  gnew_n439__spl_01
  (
    .dout(new_n439__spl_010),
    .din(new_n439__spl_01)
  );


  splt
  gnew_n439__spl_01
  (
    .dout(new_n439__spl_011),
    .din(new_n439__spl_01)
  );


  splt
  gnew_n439__spl_
  (
    .dout(new_n439__spl_1),
    .din(new_n439__spl_)
  );


  splt
  gnew_n439__spl_1
  (
    .dout(new_n439__spl_10),
    .din(new_n439__spl_1)
  );


  splt
  gnew_n439__spl_10
  (
    .dout(new_n439__spl_100),
    .din(new_n439__spl_10)
  );


  splt
  gnew_n439__spl_10
  (
    .dout(new_n439__spl_101),
    .din(new_n439__spl_10)
  );


  splt
  gnew_n439__spl_1
  (
    .dout(new_n439__spl_11),
    .din(new_n439__spl_1)
  );


  splt
  gG42
  (
    .dout(G42_spl_),
    .din(G42)
  );


  splt
  gG42_spl_
  (
    .dout(G42_spl_0),
    .din(G42_spl_)
  );


  splt
  gG42_spl_
  (
    .dout(G42_spl_1),
    .din(G42_spl_)
  );


  splt
  gnew_n445_
  (
    .dout(new_n445__spl_),
    .din(new_n445_)
  );


  splt
  gnew_n445__spl_
  (
    .dout(new_n445__spl_0),
    .din(new_n445__spl_)
  );


  splt
  gnew_n445__spl_0
  (
    .dout(new_n445__spl_00),
    .din(new_n445__spl_0)
  );


  splt
  gnew_n445__spl_00
  (
    .dout(new_n445__spl_000),
    .din(new_n445__spl_00)
  );


  splt
  gnew_n445__spl_00
  (
    .dout(new_n445__spl_001),
    .din(new_n445__spl_00)
  );


  splt
  gnew_n445__spl_0
  (
    .dout(new_n445__spl_01),
    .din(new_n445__spl_0)
  );


  splt
  gnew_n445__spl_01
  (
    .dout(new_n445__spl_010),
    .din(new_n445__spl_01)
  );


  splt
  gnew_n445__spl_01
  (
    .dout(new_n445__spl_011),
    .din(new_n445__spl_01)
  );


  splt
  gnew_n445__spl_
  (
    .dout(new_n445__spl_1),
    .din(new_n445__spl_)
  );


  splt
  gnew_n445__spl_1
  (
    .dout(new_n445__spl_10),
    .din(new_n445__spl_1)
  );


  splt
  gnew_n445__spl_1
  (
    .dout(new_n445__spl_11),
    .din(new_n445__spl_1)
  );


  splt
  gnew_n443_
  (
    .dout(new_n443__spl_),
    .din(new_n443_)
  );


  splt
  gnew_n458_
  (
    .dout(new_n458__spl_),
    .din(new_n458_)
  );


  splt
  gnew_n455_
  (
    .dout(new_n455__spl_),
    .din(new_n455_)
  );


  splt
  gnew_n457_
  (
    .dout(new_n457__spl_),
    .din(new_n457_)
  );


  splt
  gnew_n456_
  (
    .dout(new_n456__spl_),
    .din(new_n456_)
  );


  splt
  gnew_n460_
  (
    .dout(new_n460__spl_),
    .din(new_n460_)
  );


  splt
  gnew_n459_
  (
    .dout(new_n459__spl_),
    .din(new_n459_)
  );


  splt
  gnew_n477_
  (
    .dout(new_n477__spl_),
    .din(new_n477_)
  );


  splt
  gnew_n476_
  (
    .dout(new_n476__spl_),
    .din(new_n476_)
  );


  splt
  gnew_n476__spl_
  (
    .dout(new_n476__spl_0),
    .din(new_n476__spl_)
  );


  splt
  gnew_n476__spl_
  (
    .dout(new_n476__spl_1),
    .din(new_n476__spl_)
  );


  splt
  gnew_n480_
  (
    .dout(new_n480__spl_),
    .din(new_n480_)
  );


  splt
  gnew_n480__spl_
  (
    .dout(new_n480__spl_0),
    .din(new_n480__spl_)
  );


  splt
  gnew_n480__spl_
  (
    .dout(new_n480__spl_1),
    .din(new_n480__spl_)
  );


  splt
  gG18
  (
    .dout(G18_spl_),
    .din(G18)
  );


  splt
  gG18_spl_
  (
    .dout(G18_spl_0),
    .din(G18_spl_)
  );


  splt
  gG18_spl_
  (
    .dout(G18_spl_1),
    .din(G18_spl_)
  );


  splt
  gG19
  (
    .dout(G19_spl_),
    .din(G19)
  );


  splt
  gG19_spl_
  (
    .dout(G19_spl_0),
    .din(G19_spl_)
  );


  splt
  gG19_spl_
  (
    .dout(G19_spl_1),
    .din(G19_spl_)
  );


  splt
  gG20
  (
    .dout(G20_spl_),
    .din(G20)
  );


  splt
  gG20_spl_
  (
    .dout(G20_spl_0),
    .din(G20_spl_)
  );


  splt
  gG20_spl_0
  (
    .dout(G20_spl_00),
    .din(G20_spl_0)
  );


  splt
  gG20_spl_
  (
    .dout(G20_spl_1),
    .din(G20_spl_)
  );


  splt
  gnew_n522_
  (
    .dout(new_n522__spl_),
    .din(new_n522_)
  );


  splt
  gnew_n522__spl_
  (
    .dout(new_n522__spl_0),
    .din(new_n522__spl_)
  );


  splt
  gnew_n525_
  (
    .dout(new_n525__spl_),
    .din(new_n525_)
  );


  splt
  gnew_n523_
  (
    .dout(new_n523__spl_),
    .din(new_n523_)
  );


  splt
  gnew_n526_
  (
    .dout(new_n526__spl_),
    .din(new_n526_)
  );


  splt
  gnew_n532_
  (
    .dout(new_n532__spl_),
    .din(new_n532_)
  );


  splt
  gnew_n536_
  (
    .dout(new_n536__spl_),
    .din(new_n536_)
  );


  splt
  gnew_n535_
  (
    .dout(new_n535__spl_),
    .din(new_n535_)
  );


  splt
  gnew_n535__spl_
  (
    .dout(new_n535__spl_0),
    .din(new_n535__spl_)
  );


  splt
  gnew_n535__spl_0
  (
    .dout(new_n535__spl_00),
    .din(new_n535__spl_0)
  );


  splt
  gnew_n535__spl_
  (
    .dout(new_n535__spl_1),
    .din(new_n535__spl_)
  );


  splt
  gnew_n539_
  (
    .dout(new_n539__spl_),
    .din(new_n539_)
  );


  splt
  gnew_n539__spl_
  (
    .dout(new_n539__spl_0),
    .din(new_n539__spl_)
  );


  splt
  gnew_n539__spl_0
  (
    .dout(new_n539__spl_00),
    .din(new_n539__spl_0)
  );


  splt
  gnew_n539__spl_
  (
    .dout(new_n539__spl_1),
    .din(new_n539__spl_)
  );


  splt
  gnew_n540_
  (
    .dout(new_n540__spl_),
    .din(new_n540_)
  );


  splt
  gnew_n541_
  (
    .dout(new_n541__spl_),
    .din(new_n541_)
  );


  splt
  gnew_n542_
  (
    .dout(new_n542__spl_),
    .din(new_n542_)
  );


  splt
  gnew_n543_
  (
    .dout(new_n543__spl_),
    .din(new_n543_)
  );


  splt
  gnew_n543__spl_
  (
    .dout(new_n543__spl_0),
    .din(new_n543__spl_)
  );


  splt
  gnew_n550_
  (
    .dout(new_n550__spl_),
    .din(new_n550_)
  );


  splt
  gnew_n550__spl_
  (
    .dout(new_n550__spl_0),
    .din(new_n550__spl_)
  );


  splt
  gnew_n552_
  (
    .dout(new_n552__spl_),
    .din(new_n552_)
  );


  splt
  gnew_n549_
  (
    .dout(new_n549__spl_),
    .din(new_n549_)
  );


  splt
  gnew_n549__spl_
  (
    .dout(new_n549__spl_0),
    .din(new_n549__spl_)
  );


  splt
  gnew_n556_
  (
    .dout(new_n556__spl_),
    .din(new_n556_)
  );


  splt
  gnew_n556__spl_
  (
    .dout(new_n556__spl_0),
    .din(new_n556__spl_)
  );


  splt
  gnew_n556__spl_
  (
    .dout(new_n556__spl_1),
    .din(new_n556__spl_)
  );


  splt
  gnew_n547_
  (
    .dout(new_n547__spl_),
    .din(new_n547_)
  );


  splt
  gnew_n559_
  (
    .dout(new_n559__spl_),
    .din(new_n559_)
  );


  splt
  gnew_n574_
  (
    .dout(new_n574__spl_),
    .din(new_n574_)
  );


  splt
  gnew_n577_
  (
    .dout(new_n577__spl_),
    .din(new_n577_)
  );


  splt
  gnew_n577__spl_
  (
    .dout(new_n577__spl_0),
    .din(new_n577__spl_)
  );


  splt
  gnew_n583_
  (
    .dout(new_n583__spl_),
    .din(new_n583_)
  );


  splt
  gnew_n594_
  (
    .dout(new_n594__spl_),
    .din(new_n594_)
  );


  splt
  gnew_n603_
  (
    .dout(new_n603__spl_),
    .din(new_n603_)
  );


  splt
  gnew_n611_
  (
    .dout(new_n611__spl_),
    .din(new_n611_)
  );


  splt
  gG3526
  (
    .dout(G3526_spl_),
    .din(G3526)
  );


  splt
  gnew_n614_
  (
    .dout(new_n614__spl_),
    .din(new_n614_)
  );


  splt
  gnew_n614__spl_
  (
    .dout(new_n614__spl_0),
    .din(new_n614__spl_)
  );


  splt
  gnew_n614__spl_0
  (
    .dout(new_n614__spl_00),
    .din(new_n614__spl_0)
  );


  splt
  gnew_n614__spl_
  (
    .dout(new_n614__spl_1),
    .din(new_n614__spl_)
  );


  splt
  gnew_n617_
  (
    .dout(new_n617__spl_),
    .din(new_n617_)
  );


  splt
  gnew_n618_
  (
    .dout(new_n618__spl_),
    .din(new_n618_)
  );


  splt
  gnew_n620_
  (
    .dout(new_n620__spl_),
    .din(new_n620_)
  );


  splt
  gnew_n622_
  (
    .dout(new_n622__spl_),
    .din(new_n622_)
  );


  splt
  gnew_n615_
  (
    .dout(new_n615__spl_),
    .din(new_n615_)
  );


  splt
  gnew_n625_
  (
    .dout(new_n625__spl_),
    .din(new_n625_)
  );


  splt
  gnew_n630_
  (
    .dout(new_n630__spl_),
    .din(new_n630_)
  );


  splt
  gnew_n634_
  (
    .dout(new_n634__spl_),
    .din(new_n634_)
  );


  splt
  gnew_n633_
  (
    .dout(new_n633__spl_),
    .din(new_n633_)
  );


  splt
  gnew_n633__spl_
  (
    .dout(new_n633__spl_0),
    .din(new_n633__spl_)
  );


  splt
  gnew_n633__spl_
  (
    .dout(new_n633__spl_1),
    .din(new_n633__spl_)
  );


  splt
  gnew_n637_
  (
    .dout(new_n637__spl_),
    .din(new_n637_)
  );


  splt
  gnew_n637__spl_
  (
    .dout(new_n637__spl_0),
    .din(new_n637__spl_)
  );


  splt
  gnew_n637__spl_
  (
    .dout(new_n637__spl_1),
    .din(new_n637__spl_)
  );


  splt
  gnew_n663_
  (
    .dout(new_n663__spl_),
    .din(new_n663_)
  );


  splt
  gnew_n664_
  (
    .dout(new_n664__spl_),
    .din(new_n664_)
  );


  splt
  gnew_n662_
  (
    .dout(new_n662__spl_),
    .din(new_n662_)
  );


  splt
  gnew_n680_
  (
    .dout(new_n680__spl_),
    .din(new_n680_)
  );


  splt
  gnew_n680__spl_
  (
    .dout(new_n680__spl_0),
    .din(new_n680__spl_)
  );


  splt
  gnew_n701_
  (
    .dout(new_n701__spl_),
    .din(new_n701_)
  );


  splt
  gnew_n712_
  (
    .dout(new_n712__spl_),
    .din(new_n712_)
  );


  splt
  gnew_n710_
  (
    .dout(new_n710__spl_),
    .din(new_n710_)
  );


  splt
  gnew_n726_
  (
    .dout(new_n726__spl_),
    .din(new_n726_)
  );


  splt
  gnew_n729_
  (
    .dout(new_n729__spl_),
    .din(new_n729_)
  );


  splt
  gnew_n727_
  (
    .dout(new_n727__spl_),
    .din(new_n727_)
  );


  splt
  gnew_n727__spl_
  (
    .dout(new_n727__spl_0),
    .din(new_n727__spl_)
  );


  splt
  gnew_n732_
  (
    .dout(new_n732__spl_),
    .din(new_n732_)
  );


  splt
  gnew_n733_
  (
    .dout(new_n733__spl_),
    .din(new_n733_)
  );


  splt
  gnew_n733__spl_
  (
    .dout(new_n733__spl_0),
    .din(new_n733__spl_)
  );


  splt
  gnew_n736_
  (
    .dout(new_n736__spl_),
    .din(new_n736_)
  );


  splt
  gnew_n738_
  (
    .dout(new_n738__spl_),
    .din(new_n738_)
  );


  splt
  gnew_n741_
  (
    .dout(new_n741__spl_),
    .din(new_n741_)
  );


  splt
  gnew_n741__spl_
  (
    .dout(new_n741__spl_0),
    .din(new_n741__spl_)
  );


  splt
  gnew_n741__spl_
  (
    .dout(new_n741__spl_1),
    .din(new_n741__spl_)
  );


  splt
  gnew_n743_
  (
    .dout(new_n743__spl_),
    .din(new_n743_)
  );


  splt
  gnew_n743__spl_
  (
    .dout(new_n743__spl_0),
    .din(new_n743__spl_)
  );


  splt
  gnew_n735_
  (
    .dout(new_n735__spl_),
    .din(new_n735_)
  );


  splt
  gnew_n735__spl_
  (
    .dout(new_n735__spl_0),
    .din(new_n735__spl_)
  );


  splt
  gnew_n735__spl_
  (
    .dout(new_n735__spl_1),
    .din(new_n735__spl_)
  );


  splt
  gnew_n744_
  (
    .dout(new_n744__spl_),
    .din(new_n744_)
  );


  splt
  gnew_n744__spl_
  (
    .dout(new_n744__spl_0),
    .din(new_n744__spl_)
  );


  splt
  gG16
  (
    .dout(G16_spl_),
    .din(G16)
  );


  splt
  gG17
  (
    .dout(G17_spl_),
    .din(G17)
  );


  splt
  gG17_spl_
  (
    .dout(G17_spl_0),
    .din(G17_spl_)
  );


  splt
  gnew_n777_
  (
    .dout(new_n777__spl_),
    .din(new_n777_)
  );


  splt
  gnew_n748_
  (
    .dout(new_n748__spl_),
    .din(new_n748_)
  );


  splt
  gnew_n780_
  (
    .dout(new_n780__spl_),
    .din(new_n780_)
  );


  splt
  gnew_n783_
  (
    .dout(new_n783__spl_),
    .din(new_n783_)
  );


  splt
  gnew_n783__spl_
  (
    .dout(new_n783__spl_0),
    .din(new_n783__spl_)
  );


  splt
  gnew_n817_
  (
    .dout(new_n817__spl_),
    .din(new_n817_)
  );


  splt
  gnew_n778_
  (
    .dout(new_n778__spl_),
    .din(new_n778_)
  );


  splt
  gG3535
  (
    .dout(G3535_spl_),
    .din(G3535)
  );


  splt
  gG3529
  (
    .dout(G3529_spl_),
    .din(G3529)
  );


  splt
  gG3536
  (
    .dout(G3536_spl_),
    .din(G3536)
  );


  splt
  gG3531
  (
    .dout(G3531_spl_),
    .din(G3531)
  );


  splt
  gG3533
  (
    .dout(G3533_spl_),
    .din(G3533)
  );


  splt
  gG3528
  (
    .dout(G3528_spl_),
    .din(G3528)
  );


  splt
  gG3532
  (
    .dout(G3532_spl_),
    .din(G3532)
  );


  splt
  gnew_n865_
  (
    .dout(new_n865__spl_),
    .din(new_n865_)
  );


  splt
  gnew_n866_
  (
    .dout(new_n866__spl_),
    .din(new_n866_)
  );


  splt
  gnew_n864_
  (
    .dout(new_n864__spl_),
    .din(new_n864_)
  );


  splt
  gnew_n863_
  (
    .dout(new_n863__spl_),
    .din(new_n863_)
  );


  splt
  gnew_n863__spl_
  (
    .dout(new_n863__spl_0),
    .din(new_n863__spl_)
  );


  splt
  gnew_n870_
  (
    .dout(new_n870__spl_),
    .din(new_n870_)
  );


  splt
  gnew_n875_
  (
    .dout(new_n875__spl_),
    .din(new_n875_)
  );


  splt
  gnew_n877_
  (
    .dout(new_n877__spl_),
    .din(new_n877_)
  );


  splt
  gG50
  (
    .dout(G50_spl_),
    .din(G50)
  );


  splt
  gnew_n884_
  (
    .dout(new_n884__spl_),
    .din(new_n884_)
  );


  splt
  gnew_n884__spl_
  (
    .dout(new_n884__spl_0),
    .din(new_n884__spl_)
  );


  splt
  gnew_n884__spl_
  (
    .dout(new_n884__spl_1),
    .din(new_n884__spl_)
  );


  splt
  gnew_n882_
  (
    .dout(new_n882__spl_),
    .din(new_n882_)
  );


  splt
  gnew_n882__spl_
  (
    .dout(new_n882__spl_0),
    .din(new_n882__spl_)
  );


  splt
  gnew_n882__spl_
  (
    .dout(new_n882__spl_1),
    .din(new_n882__spl_)
  );


  splt
  gnew_n888_
  (
    .dout(new_n888__spl_),
    .din(new_n888_)
  );


  splt
  gnew_n880_
  (
    .dout(new_n880__spl_),
    .din(new_n880_)
  );


  splt
  gnew_n880__spl_
  (
    .dout(new_n880__spl_0),
    .din(new_n880__spl_)
  );


  splt
  gnew_n880__spl_
  (
    .dout(new_n880__spl_1),
    .din(new_n880__spl_)
  );


  splt
  gnew_n891_
  (
    .dout(new_n891__spl_),
    .din(new_n891_)
  );


  splt
  gnew_n897_
  (
    .dout(new_n897__spl_),
    .din(new_n897_)
  );


endmodule
