
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  n286_lo,
  n298_lo,
  n310_lo,
  n322_lo,
  n334_lo,
  n346_lo,
  n358_lo,
  n370_lo,
  n382_lo,
  n394_lo,
  n406_lo,
  n418_lo,
  n430_lo,
  n442_lo,
  n454_lo,
  n466_lo,
  n478_lo,
  n490_lo,
  n502_lo,
  n514_lo,
  n526_lo,
  n538_lo,
  n550_lo,
  n562_lo,
  n574_lo,
  n586_lo,
  n598_lo,
  n610_lo,
  n622_lo,
  n634_lo,
  n646_lo,
  n658_lo,
  n661_lo,
  n673_lo,
  n685_lo,
  n697_lo,
  n709_lo,
  n721_lo,
  n733_lo,
  n745_lo,
  n757_lo,
  n1589_o2,
  n1590_o2,
  n1591_o2,
  n1592_o2,
  n1593_o2,
  n1594_o2,
  n1595_o2,
  n1596_o2,
  n1597_o2,
  n1598_o2,
  n1599_o2,
  n1600_o2,
  n1601_o2,
  n1602_o2,
  n1603_o2,
  n1604_o2,
  n1605_o2,
  n1606_o2,
  n1607_o2,
  n1608_o2,
  n1609_o2,
  n1610_o2,
  n1611_o2,
  n1612_o2,
  n1613_o2,
  n1614_o2,
  n1615_o2,
  n1616_o2,
  n1617_o2,
  n1618_o2,
  n1619_o2,
  n1620_o2,
  n602_o2,
  n639_o2,
  n678_o2,
  n658_o2,
  n783_o2,
  n802_o2,
  n726_o2,
  n763_o2,
  n685_o2,
  n680_o2,
  n822_o2,
  n843_o2,
  n842_o2,
  n681_o2,
  n684_o2,
  n686_o2,
  n823_o2,
  lo002_buf_o2,
  lo006_buf_o2,
  lo010_buf_o2,
  lo014_buf_o2,
  lo018_buf_o2,
  lo022_buf_o2,
  lo026_buf_o2,
  lo030_buf_o2,
  lo034_buf_o2,
  lo038_buf_o2,
  lo042_buf_o2,
  lo046_buf_o2,
  lo050_buf_o2,
  lo054_buf_o2,
  lo058_buf_o2,
  lo062_buf_o2,
  lo066_buf_o2,
  lo070_buf_o2,
  lo074_buf_o2,
  lo078_buf_o2,
  lo082_buf_o2,
  lo086_buf_o2,
  lo090_buf_o2,
  lo094_buf_o2,
  lo098_buf_o2,
  lo102_buf_o2,
  lo106_buf_o2,
  lo110_buf_o2,
  lo114_buf_o2,
  lo118_buf_o2,
  lo122_buf_o2,
  lo126_buf_o2,
  n683_o2,
  n688_o2,
  n803_o2,
  n862_o2,
  n764_o2,
  n863_o2,
  n886_o2,
  n600_o2,
  n601_o2,
  n637_o2,
  n638_o2,
  n676_o2,
  n677_o2,
  n656_o2,
  n657_o2,
  n781_o2,
  n782_o2,
  n800_o2,
  n801_o2,
  n724_o2,
  n725_o2,
  n761_o2,
  n762_o2,
  lo129_buf_o2,
  lo133_buf_o2,
  lo137_buf_o2,
  lo141_buf_o2,
  lo145_buf_o2,
  lo149_buf_o2,
  lo153_buf_o2,
  lo157_buf_o2,
  lo161_buf_o2,
  n708_o2,
  n745_o2,
  n717_o2,
  n754_o2,
  n584_o2,
  n593_o2,
  n630_o2,
  n621_o2,
  lo001_buf_o2,
  lo005_buf_o2,
  lo009_buf_o2,
  lo013_buf_o2,
  lo017_buf_o2,
  lo021_buf_o2,
  lo025_buf_o2,
  lo029_buf_o2,
  lo033_buf_o2,
  lo037_buf_o2,
  lo041_buf_o2,
  lo045_buf_o2,
  lo049_buf_o2,
  lo053_buf_o2,
  lo057_buf_o2,
  lo061_buf_o2,
  lo065_buf_o2,
  lo069_buf_o2,
  lo073_buf_o2,
  lo077_buf_o2,
  lo081_buf_o2,
  lo085_buf_o2,
  lo089_buf_o2,
  lo093_buf_o2,
  lo097_buf_o2,
  lo101_buf_o2,
  lo105_buf_o2,
  lo109_buf_o2,
  lo113_buf_o2,
  lo117_buf_o2,
  lo121_buf_o2,
  lo125_buf_o2,
  G468,
  G469,
  G470,
  G471,
  G472,
  G473,
  G474,
  G475,
  G476,
  G477,
  G478,
  G479,
  G480,
  G481,
  G482,
  G483,
  G484,
  G485,
  G486,
  G487,
  G488,
  G489,
  G490,
  G491,
  G492,
  G493,
  G494,
  G495,
  G496,
  G497,
  G498,
  G499,
  n1020_li003_li003,
  n1032_li007_li007,
  n1044_li011_li011,
  n1056_li015_li015,
  n1068_li019_li019,
  n1080_li023_li023,
  n1092_li027_li027,
  n1104_li031_li031,
  n1116_li035_li035,
  n1128_li039_li039,
  n1140_li043_li043,
  n1152_li047_li047,
  n1164_li051_li051,
  n1176_li055_li055,
  n1188_li059_li059,
  n1200_li063_li063,
  n1212_li067_li067,
  n1224_li071_li071,
  n1236_li075_li075,
  n1248_li079_li079,
  n1260_li083_li083,
  n1272_li087_li087,
  n1284_li091_li091,
  n1296_li095_li095,
  n1308_li099_li099,
  n1320_li103_li103,
  n1332_li107_li107,
  n1344_li111_li111,
  n1356_li115_li115,
  n1368_li119_li119,
  n1380_li123_li123,
  n1392_li127_li127,
  n1395_li128_li128,
  n1407_li132_li132,
  n1419_li136_li136,
  n1431_li140_li140,
  n1443_li144_li144,
  n1455_li148_li148,
  n1467_li152_li152,
  n1479_li156_li156,
  n1491_li160_li160,
  n1589_i2,
  n1590_i2,
  n1591_i2,
  n1592_i2,
  n1593_i2,
  n1594_i2,
  n1595_i2,
  n1596_i2,
  n1597_i2,
  n1598_i2,
  n1599_i2,
  n1600_i2,
  n1601_i2,
  n1602_i2,
  n1603_i2,
  n1604_i2,
  n1605_i2,
  n1606_i2,
  n1607_i2,
  n1608_i2,
  n1609_i2,
  n1610_i2,
  n1611_i2,
  n1612_i2,
  n1613_i2,
  n1614_i2,
  n1615_i2,
  n1616_i2,
  n1617_i2,
  n1618_i2,
  n1619_i2,
  n1620_i2,
  n602_i2,
  n639_i2,
  n678_i2,
  n658_i2,
  n783_i2,
  n802_i2,
  n726_i2,
  n763_i2,
  n685_i2,
  n680_i2,
  n822_i2,
  n843_i2,
  n842_i2,
  n681_i2,
  n684_i2,
  n686_i2,
  n823_i2,
  lo002_buf_i2,
  lo006_buf_i2,
  lo010_buf_i2,
  lo014_buf_i2,
  lo018_buf_i2,
  lo022_buf_i2,
  lo026_buf_i2,
  lo030_buf_i2,
  lo034_buf_i2,
  lo038_buf_i2,
  lo042_buf_i2,
  lo046_buf_i2,
  lo050_buf_i2,
  lo054_buf_i2,
  lo058_buf_i2,
  lo062_buf_i2,
  lo066_buf_i2,
  lo070_buf_i2,
  lo074_buf_i2,
  lo078_buf_i2,
  lo082_buf_i2,
  lo086_buf_i2,
  lo090_buf_i2,
  lo094_buf_i2,
  lo098_buf_i2,
  lo102_buf_i2,
  lo106_buf_i2,
  lo110_buf_i2,
  lo114_buf_i2,
  lo118_buf_i2,
  lo122_buf_i2,
  lo126_buf_i2,
  n683_i2,
  n688_i2,
  n803_i2,
  n862_i2,
  n764_i2,
  n863_i2,
  n886_i2,
  n600_i2,
  n601_i2,
  n637_i2,
  n638_i2,
  n676_i2,
  n677_i2,
  n656_i2,
  n657_i2,
  n781_i2,
  n782_i2,
  n800_i2,
  n801_i2,
  n724_i2,
  n725_i2,
  n761_i2,
  n762_i2,
  lo129_buf_i2,
  lo133_buf_i2,
  lo137_buf_i2,
  lo141_buf_i2,
  lo145_buf_i2,
  lo149_buf_i2,
  lo153_buf_i2,
  lo157_buf_i2,
  lo161_buf_i2,
  n708_i2,
  n745_i2,
  n717_i2,
  n754_i2,
  n584_i2,
  n593_i2,
  n630_i2,
  n621_i2,
  lo001_buf_i2,
  lo005_buf_i2,
  lo009_buf_i2,
  lo013_buf_i2,
  lo017_buf_i2,
  lo021_buf_i2,
  lo025_buf_i2,
  lo029_buf_i2,
  lo033_buf_i2,
  lo037_buf_i2,
  lo041_buf_i2,
  lo045_buf_i2,
  lo049_buf_i2,
  lo053_buf_i2,
  lo057_buf_i2,
  lo061_buf_i2,
  lo065_buf_i2,
  lo069_buf_i2,
  lo073_buf_i2,
  lo077_buf_i2,
  lo081_buf_i2,
  lo085_buf_i2,
  lo089_buf_i2,
  lo093_buf_i2,
  lo097_buf_i2,
  lo101_buf_i2,
  lo105_buf_i2,
  lo109_buf_i2,
  lo113_buf_i2,
  lo117_buf_i2,
  lo121_buf_i2,
  lo125_buf_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input n286_lo;input n298_lo;input n310_lo;input n322_lo;input n334_lo;input n346_lo;input n358_lo;input n370_lo;input n382_lo;input n394_lo;input n406_lo;input n418_lo;input n430_lo;input n442_lo;input n454_lo;input n466_lo;input n478_lo;input n490_lo;input n502_lo;input n514_lo;input n526_lo;input n538_lo;input n550_lo;input n562_lo;input n574_lo;input n586_lo;input n598_lo;input n610_lo;input n622_lo;input n634_lo;input n646_lo;input n658_lo;input n661_lo;input n673_lo;input n685_lo;input n697_lo;input n709_lo;input n721_lo;input n733_lo;input n745_lo;input n757_lo;input n1589_o2;input n1590_o2;input n1591_o2;input n1592_o2;input n1593_o2;input n1594_o2;input n1595_o2;input n1596_o2;input n1597_o2;input n1598_o2;input n1599_o2;input n1600_o2;input n1601_o2;input n1602_o2;input n1603_o2;input n1604_o2;input n1605_o2;input n1606_o2;input n1607_o2;input n1608_o2;input n1609_o2;input n1610_o2;input n1611_o2;input n1612_o2;input n1613_o2;input n1614_o2;input n1615_o2;input n1616_o2;input n1617_o2;input n1618_o2;input n1619_o2;input n1620_o2;input n602_o2;input n639_o2;input n678_o2;input n658_o2;input n783_o2;input n802_o2;input n726_o2;input n763_o2;input n685_o2;input n680_o2;input n822_o2;input n843_o2;input n842_o2;input n681_o2;input n684_o2;input n686_o2;input n823_o2;input lo002_buf_o2;input lo006_buf_o2;input lo010_buf_o2;input lo014_buf_o2;input lo018_buf_o2;input lo022_buf_o2;input lo026_buf_o2;input lo030_buf_o2;input lo034_buf_o2;input lo038_buf_o2;input lo042_buf_o2;input lo046_buf_o2;input lo050_buf_o2;input lo054_buf_o2;input lo058_buf_o2;input lo062_buf_o2;input lo066_buf_o2;input lo070_buf_o2;input lo074_buf_o2;input lo078_buf_o2;input lo082_buf_o2;input lo086_buf_o2;input lo090_buf_o2;input lo094_buf_o2;input lo098_buf_o2;input lo102_buf_o2;input lo106_buf_o2;input lo110_buf_o2;input lo114_buf_o2;input lo118_buf_o2;input lo122_buf_o2;input lo126_buf_o2;input n683_o2;input n688_o2;input n803_o2;input n862_o2;input n764_o2;input n863_o2;input n886_o2;input n600_o2;input n601_o2;input n637_o2;input n638_o2;input n676_o2;input n677_o2;input n656_o2;input n657_o2;input n781_o2;input n782_o2;input n800_o2;input n801_o2;input n724_o2;input n725_o2;input n761_o2;input n762_o2;input lo129_buf_o2;input lo133_buf_o2;input lo137_buf_o2;input lo141_buf_o2;input lo145_buf_o2;input lo149_buf_o2;input lo153_buf_o2;input lo157_buf_o2;input lo161_buf_o2;input n708_o2;input n745_o2;input n717_o2;input n754_o2;input n584_o2;input n593_o2;input n630_o2;input n621_o2;input lo001_buf_o2;input lo005_buf_o2;input lo009_buf_o2;input lo013_buf_o2;input lo017_buf_o2;input lo021_buf_o2;input lo025_buf_o2;input lo029_buf_o2;input lo033_buf_o2;input lo037_buf_o2;input lo041_buf_o2;input lo045_buf_o2;input lo049_buf_o2;input lo053_buf_o2;input lo057_buf_o2;input lo061_buf_o2;input lo065_buf_o2;input lo069_buf_o2;input lo073_buf_o2;input lo077_buf_o2;input lo081_buf_o2;input lo085_buf_o2;input lo089_buf_o2;input lo093_buf_o2;input lo097_buf_o2;input lo101_buf_o2;input lo105_buf_o2;input lo109_buf_o2;input lo113_buf_o2;input lo117_buf_o2;input lo121_buf_o2;input lo125_buf_o2;
  output G468;output G469;output G470;output G471;output G472;output G473;output G474;output G475;output G476;output G477;output G478;output G479;output G480;output G481;output G482;output G483;output G484;output G485;output G486;output G487;output G488;output G489;output G490;output G491;output G492;output G493;output G494;output G495;output G496;output G497;output G498;output G499;output n1020_li003_li003;output n1032_li007_li007;output n1044_li011_li011;output n1056_li015_li015;output n1068_li019_li019;output n1080_li023_li023;output n1092_li027_li027;output n1104_li031_li031;output n1116_li035_li035;output n1128_li039_li039;output n1140_li043_li043;output n1152_li047_li047;output n1164_li051_li051;output n1176_li055_li055;output n1188_li059_li059;output n1200_li063_li063;output n1212_li067_li067;output n1224_li071_li071;output n1236_li075_li075;output n1248_li079_li079;output n1260_li083_li083;output n1272_li087_li087;output n1284_li091_li091;output n1296_li095_li095;output n1308_li099_li099;output n1320_li103_li103;output n1332_li107_li107;output n1344_li111_li111;output n1356_li115_li115;output n1368_li119_li119;output n1380_li123_li123;output n1392_li127_li127;output n1395_li128_li128;output n1407_li132_li132;output n1419_li136_li136;output n1431_li140_li140;output n1443_li144_li144;output n1455_li148_li148;output n1467_li152_li152;output n1479_li156_li156;output n1491_li160_li160;output n1589_i2;output n1590_i2;output n1591_i2;output n1592_i2;output n1593_i2;output n1594_i2;output n1595_i2;output n1596_i2;output n1597_i2;output n1598_i2;output n1599_i2;output n1600_i2;output n1601_i2;output n1602_i2;output n1603_i2;output n1604_i2;output n1605_i2;output n1606_i2;output n1607_i2;output n1608_i2;output n1609_i2;output n1610_i2;output n1611_i2;output n1612_i2;output n1613_i2;output n1614_i2;output n1615_i2;output n1616_i2;output n1617_i2;output n1618_i2;output n1619_i2;output n1620_i2;output n602_i2;output n639_i2;output n678_i2;output n658_i2;output n783_i2;output n802_i2;output n726_i2;output n763_i2;output n685_i2;output n680_i2;output n822_i2;output n843_i2;output n842_i2;output n681_i2;output n684_i2;output n686_i2;output n823_i2;output lo002_buf_i2;output lo006_buf_i2;output lo010_buf_i2;output lo014_buf_i2;output lo018_buf_i2;output lo022_buf_i2;output lo026_buf_i2;output lo030_buf_i2;output lo034_buf_i2;output lo038_buf_i2;output lo042_buf_i2;output lo046_buf_i2;output lo050_buf_i2;output lo054_buf_i2;output lo058_buf_i2;output lo062_buf_i2;output lo066_buf_i2;output lo070_buf_i2;output lo074_buf_i2;output lo078_buf_i2;output lo082_buf_i2;output lo086_buf_i2;output lo090_buf_i2;output lo094_buf_i2;output lo098_buf_i2;output lo102_buf_i2;output lo106_buf_i2;output lo110_buf_i2;output lo114_buf_i2;output lo118_buf_i2;output lo122_buf_i2;output lo126_buf_i2;output n683_i2;output n688_i2;output n803_i2;output n862_i2;output n764_i2;output n863_i2;output n886_i2;output n600_i2;output n601_i2;output n637_i2;output n638_i2;output n676_i2;output n677_i2;output n656_i2;output n657_i2;output n781_i2;output n782_i2;output n800_i2;output n801_i2;output n724_i2;output n725_i2;output n761_i2;output n762_i2;output lo129_buf_i2;output lo133_buf_i2;output lo137_buf_i2;output lo141_buf_i2;output lo145_buf_i2;output lo149_buf_i2;output lo153_buf_i2;output lo157_buf_i2;output lo161_buf_i2;output n708_i2;output n745_i2;output n717_i2;output n754_i2;output n584_i2;output n593_i2;output n630_i2;output n621_i2;output lo001_buf_i2;output lo005_buf_i2;output lo009_buf_i2;output lo013_buf_i2;output lo017_buf_i2;output lo021_buf_i2;output lo025_buf_i2;output lo029_buf_i2;output lo033_buf_i2;output lo037_buf_i2;output lo041_buf_i2;output lo045_buf_i2;output lo049_buf_i2;output lo053_buf_i2;output lo057_buf_i2;output lo061_buf_i2;output lo065_buf_i2;output lo069_buf_i2;output lo073_buf_i2;output lo077_buf_i2;output lo081_buf_i2;output lo085_buf_i2;output lo089_buf_i2;output lo093_buf_i2;output lo097_buf_i2;output lo101_buf_i2;output lo105_buf_i2;output lo109_buf_i2;output lo113_buf_i2;output lo117_buf_i2;output lo121_buf_i2;output lo125_buf_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire n286_lo_p;
  wire n286_lo_n;
  wire n298_lo_p;
  wire n298_lo_n;
  wire n310_lo_p;
  wire n310_lo_n;
  wire n322_lo_p;
  wire n322_lo_n;
  wire n334_lo_p;
  wire n334_lo_n;
  wire n346_lo_p;
  wire n346_lo_n;
  wire n358_lo_p;
  wire n358_lo_n;
  wire n370_lo_p;
  wire n370_lo_n;
  wire n382_lo_p;
  wire n382_lo_n;
  wire n394_lo_p;
  wire n394_lo_n;
  wire n406_lo_p;
  wire n406_lo_n;
  wire n418_lo_p;
  wire n418_lo_n;
  wire n430_lo_p;
  wire n430_lo_n;
  wire n442_lo_p;
  wire n442_lo_n;
  wire n454_lo_p;
  wire n454_lo_n;
  wire n466_lo_p;
  wire n466_lo_n;
  wire n478_lo_p;
  wire n478_lo_n;
  wire n490_lo_p;
  wire n490_lo_n;
  wire n502_lo_p;
  wire n502_lo_n;
  wire n514_lo_p;
  wire n514_lo_n;
  wire n526_lo_p;
  wire n526_lo_n;
  wire n538_lo_p;
  wire n538_lo_n;
  wire n550_lo_p;
  wire n550_lo_n;
  wire n562_lo_p;
  wire n562_lo_n;
  wire n574_lo_p;
  wire n574_lo_n;
  wire n586_lo_p;
  wire n586_lo_n;
  wire n598_lo_p;
  wire n598_lo_n;
  wire n610_lo_p;
  wire n610_lo_n;
  wire n622_lo_p;
  wire n622_lo_n;
  wire n634_lo_p;
  wire n634_lo_n;
  wire n646_lo_p;
  wire n646_lo_n;
  wire n658_lo_p;
  wire n658_lo_n;
  wire n661_lo_p;
  wire n661_lo_n;
  wire n673_lo_p;
  wire n673_lo_n;
  wire n685_lo_p;
  wire n685_lo_n;
  wire n697_lo_p;
  wire n697_lo_n;
  wire n709_lo_p;
  wire n709_lo_n;
  wire n721_lo_p;
  wire n721_lo_n;
  wire n733_lo_p;
  wire n733_lo_n;
  wire n745_lo_p;
  wire n745_lo_n;
  wire n757_lo_p;
  wire n757_lo_n;
  wire n1589_o2_p;
  wire n1589_o2_n;
  wire n1590_o2_p;
  wire n1590_o2_n;
  wire n1591_o2_p;
  wire n1591_o2_n;
  wire n1592_o2_p;
  wire n1592_o2_n;
  wire n1593_o2_p;
  wire n1593_o2_n;
  wire n1594_o2_p;
  wire n1594_o2_n;
  wire n1595_o2_p;
  wire n1595_o2_n;
  wire n1596_o2_p;
  wire n1596_o2_n;
  wire n1597_o2_p;
  wire n1597_o2_n;
  wire n1598_o2_p;
  wire n1598_o2_n;
  wire n1599_o2_p;
  wire n1599_o2_n;
  wire n1600_o2_p;
  wire n1600_o2_n;
  wire n1601_o2_p;
  wire n1601_o2_n;
  wire n1602_o2_p;
  wire n1602_o2_n;
  wire n1603_o2_p;
  wire n1603_o2_n;
  wire n1604_o2_p;
  wire n1604_o2_n;
  wire n1605_o2_p;
  wire n1605_o2_n;
  wire n1606_o2_p;
  wire n1606_o2_n;
  wire n1607_o2_p;
  wire n1607_o2_n;
  wire n1608_o2_p;
  wire n1608_o2_n;
  wire n1609_o2_p;
  wire n1609_o2_n;
  wire n1610_o2_p;
  wire n1610_o2_n;
  wire n1611_o2_p;
  wire n1611_o2_n;
  wire n1612_o2_p;
  wire n1612_o2_n;
  wire n1613_o2_p;
  wire n1613_o2_n;
  wire n1614_o2_p;
  wire n1614_o2_n;
  wire n1615_o2_p;
  wire n1615_o2_n;
  wire n1616_o2_p;
  wire n1616_o2_n;
  wire n1617_o2_p;
  wire n1617_o2_n;
  wire n1618_o2_p;
  wire n1618_o2_n;
  wire n1619_o2_p;
  wire n1619_o2_n;
  wire n1620_o2_p;
  wire n1620_o2_n;
  wire n602_o2_p;
  wire n602_o2_n;
  wire n639_o2_p;
  wire n639_o2_n;
  wire n678_o2_p;
  wire n678_o2_n;
  wire n658_o2_p;
  wire n658_o2_n;
  wire n783_o2_p;
  wire n783_o2_n;
  wire n802_o2_p;
  wire n802_o2_n;
  wire n726_o2_p;
  wire n726_o2_n;
  wire n763_o2_p;
  wire n763_o2_n;
  wire n685_o2_p;
  wire n685_o2_n;
  wire n680_o2_p;
  wire n680_o2_n;
  wire n822_o2_p;
  wire n822_o2_n;
  wire n843_o2_p;
  wire n843_o2_n;
  wire n842_o2_p;
  wire n842_o2_n;
  wire n681_o2_p;
  wire n681_o2_n;
  wire n684_o2_p;
  wire n684_o2_n;
  wire n686_o2_p;
  wire n686_o2_n;
  wire n823_o2_p;
  wire n823_o2_n;
  wire lo002_buf_o2_p;
  wire lo002_buf_o2_n;
  wire lo006_buf_o2_p;
  wire lo006_buf_o2_n;
  wire lo010_buf_o2_p;
  wire lo010_buf_o2_n;
  wire lo014_buf_o2_p;
  wire lo014_buf_o2_n;
  wire lo018_buf_o2_p;
  wire lo018_buf_o2_n;
  wire lo022_buf_o2_p;
  wire lo022_buf_o2_n;
  wire lo026_buf_o2_p;
  wire lo026_buf_o2_n;
  wire lo030_buf_o2_p;
  wire lo030_buf_o2_n;
  wire lo034_buf_o2_p;
  wire lo034_buf_o2_n;
  wire lo038_buf_o2_p;
  wire lo038_buf_o2_n;
  wire lo042_buf_o2_p;
  wire lo042_buf_o2_n;
  wire lo046_buf_o2_p;
  wire lo046_buf_o2_n;
  wire lo050_buf_o2_p;
  wire lo050_buf_o2_n;
  wire lo054_buf_o2_p;
  wire lo054_buf_o2_n;
  wire lo058_buf_o2_p;
  wire lo058_buf_o2_n;
  wire lo062_buf_o2_p;
  wire lo062_buf_o2_n;
  wire lo066_buf_o2_p;
  wire lo066_buf_o2_n;
  wire lo070_buf_o2_p;
  wire lo070_buf_o2_n;
  wire lo074_buf_o2_p;
  wire lo074_buf_o2_n;
  wire lo078_buf_o2_p;
  wire lo078_buf_o2_n;
  wire lo082_buf_o2_p;
  wire lo082_buf_o2_n;
  wire lo086_buf_o2_p;
  wire lo086_buf_o2_n;
  wire lo090_buf_o2_p;
  wire lo090_buf_o2_n;
  wire lo094_buf_o2_p;
  wire lo094_buf_o2_n;
  wire lo098_buf_o2_p;
  wire lo098_buf_o2_n;
  wire lo102_buf_o2_p;
  wire lo102_buf_o2_n;
  wire lo106_buf_o2_p;
  wire lo106_buf_o2_n;
  wire lo110_buf_o2_p;
  wire lo110_buf_o2_n;
  wire lo114_buf_o2_p;
  wire lo114_buf_o2_n;
  wire lo118_buf_o2_p;
  wire lo118_buf_o2_n;
  wire lo122_buf_o2_p;
  wire lo122_buf_o2_n;
  wire lo126_buf_o2_p;
  wire lo126_buf_o2_n;
  wire n683_o2_p;
  wire n683_o2_n;
  wire n688_o2_p;
  wire n688_o2_n;
  wire n803_o2_p;
  wire n803_o2_n;
  wire n862_o2_p;
  wire n862_o2_n;
  wire n764_o2_p;
  wire n764_o2_n;
  wire n863_o2_p;
  wire n863_o2_n;
  wire n886_o2_p;
  wire n886_o2_n;
  wire n600_o2_p;
  wire n600_o2_n;
  wire n601_o2_p;
  wire n601_o2_n;
  wire n637_o2_p;
  wire n637_o2_n;
  wire n638_o2_p;
  wire n638_o2_n;
  wire n676_o2_p;
  wire n676_o2_n;
  wire n677_o2_p;
  wire n677_o2_n;
  wire n656_o2_p;
  wire n656_o2_n;
  wire n657_o2_p;
  wire n657_o2_n;
  wire n781_o2_p;
  wire n781_o2_n;
  wire n782_o2_p;
  wire n782_o2_n;
  wire n800_o2_p;
  wire n800_o2_n;
  wire n801_o2_p;
  wire n801_o2_n;
  wire n724_o2_p;
  wire n724_o2_n;
  wire n725_o2_p;
  wire n725_o2_n;
  wire n761_o2_p;
  wire n761_o2_n;
  wire n762_o2_p;
  wire n762_o2_n;
  wire lo129_buf_o2_p;
  wire lo129_buf_o2_n;
  wire lo133_buf_o2_p;
  wire lo133_buf_o2_n;
  wire lo137_buf_o2_p;
  wire lo137_buf_o2_n;
  wire lo141_buf_o2_p;
  wire lo141_buf_o2_n;
  wire lo145_buf_o2_p;
  wire lo145_buf_o2_n;
  wire lo149_buf_o2_p;
  wire lo149_buf_o2_n;
  wire lo153_buf_o2_p;
  wire lo153_buf_o2_n;
  wire lo157_buf_o2_p;
  wire lo157_buf_o2_n;
  wire lo161_buf_o2_p;
  wire lo161_buf_o2_n;
  wire n708_o2_p;
  wire n708_o2_n;
  wire n745_o2_p;
  wire n745_o2_n;
  wire n717_o2_p;
  wire n717_o2_n;
  wire n754_o2_p;
  wire n754_o2_n;
  wire n584_o2_p;
  wire n584_o2_n;
  wire n593_o2_p;
  wire n593_o2_n;
  wire n630_o2_p;
  wire n630_o2_n;
  wire n621_o2_p;
  wire n621_o2_n;
  wire lo001_buf_o2_p;
  wire lo001_buf_o2_n;
  wire lo005_buf_o2_p;
  wire lo005_buf_o2_n;
  wire lo009_buf_o2_p;
  wire lo009_buf_o2_n;
  wire lo013_buf_o2_p;
  wire lo013_buf_o2_n;
  wire lo017_buf_o2_p;
  wire lo017_buf_o2_n;
  wire lo021_buf_o2_p;
  wire lo021_buf_o2_n;
  wire lo025_buf_o2_p;
  wire lo025_buf_o2_n;
  wire lo029_buf_o2_p;
  wire lo029_buf_o2_n;
  wire lo033_buf_o2_p;
  wire lo033_buf_o2_n;
  wire lo037_buf_o2_p;
  wire lo037_buf_o2_n;
  wire lo041_buf_o2_p;
  wire lo041_buf_o2_n;
  wire lo045_buf_o2_p;
  wire lo045_buf_o2_n;
  wire lo049_buf_o2_p;
  wire lo049_buf_o2_n;
  wire lo053_buf_o2_p;
  wire lo053_buf_o2_n;
  wire lo057_buf_o2_p;
  wire lo057_buf_o2_n;
  wire lo061_buf_o2_p;
  wire lo061_buf_o2_n;
  wire lo065_buf_o2_p;
  wire lo065_buf_o2_n;
  wire lo069_buf_o2_p;
  wire lo069_buf_o2_n;
  wire lo073_buf_o2_p;
  wire lo073_buf_o2_n;
  wire lo077_buf_o2_p;
  wire lo077_buf_o2_n;
  wire lo081_buf_o2_p;
  wire lo081_buf_o2_n;
  wire lo085_buf_o2_p;
  wire lo085_buf_o2_n;
  wire lo089_buf_o2_p;
  wire lo089_buf_o2_n;
  wire lo093_buf_o2_p;
  wire lo093_buf_o2_n;
  wire lo097_buf_o2_p;
  wire lo097_buf_o2_n;
  wire lo101_buf_o2_p;
  wire lo101_buf_o2_n;
  wire lo105_buf_o2_p;
  wire lo105_buf_o2_n;
  wire lo109_buf_o2_p;
  wire lo109_buf_o2_n;
  wire lo113_buf_o2_p;
  wire lo113_buf_o2_n;
  wire lo117_buf_o2_p;
  wire lo117_buf_o2_n;
  wire lo121_buf_o2_p;
  wire lo121_buf_o2_n;
  wire lo125_buf_o2_p;
  wire lo125_buf_o2_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g236_n_spl_;
  wire g236_n_spl_0;
  wire g236_n_spl_1;
  wire g236_p_spl_;
  wire g236_p_spl_0;
  wire g236_p_spl_1;
  wire n602_o2_p_spl_;
  wire n602_o2_p_spl_0;
  wire n602_o2_p_spl_1;
  wire g238_p_spl_;
  wire g238_p_spl_0;
  wire g238_p_spl_1;
  wire n602_o2_n_spl_;
  wire n602_o2_n_spl_0;
  wire n602_o2_n_spl_1;
  wire g238_n_spl_;
  wire g238_n_spl_0;
  wire g238_n_spl_1;
  wire n639_o2_p_spl_;
  wire n639_o2_p_spl_0;
  wire n639_o2_p_spl_00;
  wire n639_o2_p_spl_1;
  wire n639_o2_n_spl_;
  wire n639_o2_n_spl_0;
  wire n639_o2_n_spl_00;
  wire n639_o2_n_spl_1;
  wire n678_o2_p_spl_;
  wire n678_o2_p_spl_0;
  wire n678_o2_p_spl_00;
  wire n678_o2_p_spl_01;
  wire n678_o2_p_spl_1;
  wire n678_o2_n_spl_;
  wire n678_o2_n_spl_0;
  wire n678_o2_n_spl_00;
  wire n678_o2_n_spl_01;
  wire n678_o2_n_spl_1;
  wire n658_o2_p_spl_;
  wire n658_o2_p_spl_0;
  wire n658_o2_p_spl_1;
  wire n658_o2_n_spl_;
  wire n658_o2_n_spl_0;
  wire n658_o2_n_spl_1;
  wire g256_p_spl_;
  wire g256_p_spl_0;
  wire g256_p_spl_1;
  wire g256_n_spl_;
  wire g256_n_spl_0;
  wire g256_n_spl_1;
  wire g274_p_spl_;
  wire g274_p_spl_0;
  wire g274_p_spl_1;
  wire g274_n_spl_;
  wire g274_n_spl_0;
  wire g274_n_spl_1;
  wire g292_p_spl_;
  wire g292_p_spl_0;
  wire g292_p_spl_1;
  wire g292_n_spl_;
  wire g292_n_spl_0;
  wire g292_n_spl_1;
  wire n886_o2_p_spl_;
  wire n886_o2_p_spl_0;
  wire n886_o2_p_spl_1;
  wire n886_o2_n_spl_;
  wire n886_o2_n_spl_0;
  wire n886_o2_n_spl_1;
  wire n783_o2_p_spl_;
  wire n783_o2_p_spl_0;
  wire n783_o2_p_spl_1;
  wire g310_p_spl_;
  wire g310_p_spl_0;
  wire g310_p_spl_1;
  wire n783_o2_n_spl_;
  wire n783_o2_n_spl_0;
  wire n783_o2_n_spl_1;
  wire g310_n_spl_;
  wire g310_n_spl_0;
  wire g310_n_spl_1;
  wire n802_o2_p_spl_;
  wire n802_o2_p_spl_0;
  wire n802_o2_p_spl_1;
  wire n802_o2_n_spl_;
  wire n802_o2_n_spl_0;
  wire n802_o2_n_spl_1;
  wire n726_o2_p_spl_;
  wire n726_o2_p_spl_0;
  wire n726_o2_p_spl_1;
  wire n726_o2_n_spl_;
  wire n726_o2_n_spl_0;
  wire n726_o2_n_spl_1;
  wire n763_o2_p_spl_;
  wire n763_o2_p_spl_0;
  wire n763_o2_p_spl_1;
  wire n763_o2_n_spl_;
  wire n763_o2_n_spl_0;
  wire n763_o2_n_spl_1;
  wire g328_p_spl_;
  wire g328_p_spl_0;
  wire g328_p_spl_1;
  wire g328_n_spl_;
  wire g328_n_spl_0;
  wire g328_n_spl_1;
  wire g346_p_spl_;
  wire g346_p_spl_0;
  wire g346_p_spl_1;
  wire g346_n_spl_;
  wire g346_n_spl_0;
  wire g346_n_spl_1;
  wire g364_p_spl_;
  wire g364_p_spl_0;
  wire g364_p_spl_1;
  wire g364_n_spl_;
  wire g364_n_spl_0;
  wire g364_n_spl_1;
  wire g382_n_spl_;
  wire g382_n_spl_0;
  wire g383_n_spl_;
  wire g383_n_spl_0;
  wire g385_p_spl_;
  wire g385_p_spl_0;
  wire g388_p_spl_;
  wire g388_p_spl_0;
  wire g385_n_spl_;
  wire g385_n_spl_0;
  wire g388_n_spl_;
  wire g388_n_spl_0;
  wire g386_p_spl_;
  wire g386_p_spl_0;
  wire g387_p_spl_;
  wire g387_p_spl_0;
  wire g381_n_spl_;
  wire g381_n_spl_0;
  wire g390_n_spl_;
  wire g384_n_spl_;
  wire g384_n_spl_0;
  wire g395_n_spl_;
  wire g389_n_spl_;
  wire g386_n_spl_;
  wire g386_n_spl_0;
  wire g387_n_spl_;
  wire g387_n_spl_0;
  wire g394_n_spl_;
  wire g396_n_spl_;
  wire g397_n_spl_;
  wire g391_n_spl_;
  wire g392_n_spl_;
  wire g398_n_spl_;
  wire g393_n_spl_;
  wire lo002_buf_o2_p_spl_;
  wire lo002_buf_o2_p_spl_0;
  wire lo018_buf_o2_n_spl_;
  wire lo002_buf_o2_n_spl_;
  wire lo018_buf_o2_p_spl_;
  wire lo018_buf_o2_p_spl_0;
  wire lo034_buf_o2_p_spl_;
  wire lo034_buf_o2_p_spl_0;
  wire lo050_buf_o2_n_spl_;
  wire lo034_buf_o2_n_spl_;
  wire lo050_buf_o2_p_spl_;
  wire lo050_buf_o2_p_spl_0;
  wire lo161_buf_o2_p_spl_;
  wire lo161_buf_o2_p_spl_0;
  wire lo161_buf_o2_p_spl_00;
  wire lo161_buf_o2_p_spl_01;
  wire lo161_buf_o2_p_spl_1;
  wire lo161_buf_o2_p_spl_10;
  wire lo161_buf_o2_p_spl_11;
  wire lo161_buf_o2_n_spl_;
  wire lo161_buf_o2_n_spl_0;
  wire lo161_buf_o2_n_spl_00;
  wire lo161_buf_o2_n_spl_01;
  wire lo161_buf_o2_n_spl_1;
  wire lo161_buf_o2_n_spl_10;
  wire lo161_buf_o2_n_spl_11;
  wire n584_o2_n_spl_;
  wire n584_o2_n_spl_0;
  wire n584_o2_n_spl_1;
  wire n593_o2_p_spl_;
  wire n593_o2_p_spl_0;
  wire n593_o2_p_spl_1;
  wire n584_o2_p_spl_;
  wire n584_o2_p_spl_0;
  wire n584_o2_p_spl_1;
  wire n593_o2_n_spl_;
  wire n593_o2_n_spl_0;
  wire n593_o2_n_spl_1;
  wire g421_n_spl_;
  wire g428_p_spl_;
  wire lo006_buf_o2_p_spl_;
  wire lo006_buf_o2_p_spl_0;
  wire lo022_buf_o2_n_spl_;
  wire lo006_buf_o2_n_spl_;
  wire lo022_buf_o2_p_spl_;
  wire lo022_buf_o2_p_spl_0;
  wire lo038_buf_o2_p_spl_;
  wire lo038_buf_o2_p_spl_0;
  wire lo054_buf_o2_n_spl_;
  wire lo038_buf_o2_n_spl_;
  wire lo054_buf_o2_p_spl_;
  wire lo054_buf_o2_p_spl_0;
  wire n630_o2_p_spl_;
  wire n630_o2_p_spl_0;
  wire n630_o2_p_spl_1;
  wire n621_o2_n_spl_;
  wire n621_o2_n_spl_0;
  wire n621_o2_n_spl_1;
  wire n630_o2_n_spl_;
  wire n630_o2_n_spl_0;
  wire n630_o2_n_spl_1;
  wire n621_o2_p_spl_;
  wire n621_o2_p_spl_0;
  wire n621_o2_p_spl_1;
  wire g439_n_spl_;
  wire g446_p_spl_;
  wire lo010_buf_o2_p_spl_;
  wire lo010_buf_o2_p_spl_0;
  wire lo026_buf_o2_n_spl_;
  wire lo010_buf_o2_n_spl_;
  wire lo026_buf_o2_p_spl_;
  wire lo026_buf_o2_p_spl_0;
  wire lo042_buf_o2_p_spl_;
  wire lo042_buf_o2_p_spl_0;
  wire lo058_buf_o2_n_spl_;
  wire lo042_buf_o2_n_spl_;
  wire lo058_buf_o2_p_spl_;
  wire lo058_buf_o2_p_spl_0;
  wire g457_n_spl_;
  wire g464_p_spl_;
  wire lo014_buf_o2_p_spl_;
  wire lo014_buf_o2_p_spl_0;
  wire lo030_buf_o2_n_spl_;
  wire lo014_buf_o2_n_spl_;
  wire lo030_buf_o2_p_spl_;
  wire lo030_buf_o2_p_spl_0;
  wire lo046_buf_o2_p_spl_;
  wire lo046_buf_o2_p_spl_0;
  wire lo062_buf_o2_n_spl_;
  wire lo046_buf_o2_n_spl_;
  wire lo062_buf_o2_p_spl_;
  wire lo062_buf_o2_p_spl_0;
  wire g475_n_spl_;
  wire g482_p_spl_;
  wire lo066_buf_o2_p_spl_;
  wire lo066_buf_o2_p_spl_0;
  wire lo082_buf_o2_n_spl_;
  wire lo066_buf_o2_n_spl_;
  wire lo082_buf_o2_p_spl_;
  wire lo082_buf_o2_p_spl_0;
  wire lo098_buf_o2_p_spl_;
  wire lo098_buf_o2_p_spl_0;
  wire lo114_buf_o2_n_spl_;
  wire lo098_buf_o2_n_spl_;
  wire lo114_buf_o2_p_spl_;
  wire lo114_buf_o2_p_spl_0;
  wire n708_o2_n_spl_;
  wire n708_o2_n_spl_0;
  wire n708_o2_n_spl_1;
  wire n745_o2_p_spl_;
  wire n745_o2_p_spl_0;
  wire n745_o2_p_spl_1;
  wire n708_o2_p_spl_;
  wire n708_o2_p_spl_0;
  wire n708_o2_p_spl_1;
  wire n745_o2_n_spl_;
  wire n745_o2_n_spl_0;
  wire n745_o2_n_spl_1;
  wire g493_n_spl_;
  wire g500_p_spl_;
  wire lo070_buf_o2_p_spl_;
  wire lo070_buf_o2_p_spl_0;
  wire lo086_buf_o2_n_spl_;
  wire lo070_buf_o2_n_spl_;
  wire lo086_buf_o2_p_spl_;
  wire lo086_buf_o2_p_spl_0;
  wire lo102_buf_o2_p_spl_;
  wire lo102_buf_o2_p_spl_0;
  wire lo118_buf_o2_n_spl_;
  wire lo102_buf_o2_n_spl_;
  wire lo118_buf_o2_p_spl_;
  wire lo118_buf_o2_p_spl_0;
  wire n717_o2_n_spl_;
  wire n717_o2_n_spl_0;
  wire n717_o2_n_spl_1;
  wire n754_o2_p_spl_;
  wire n754_o2_p_spl_0;
  wire n754_o2_p_spl_1;
  wire n717_o2_p_spl_;
  wire n717_o2_p_spl_0;
  wire n717_o2_p_spl_1;
  wire n754_o2_n_spl_;
  wire n754_o2_n_spl_0;
  wire n754_o2_n_spl_1;
  wire g511_n_spl_;
  wire g518_p_spl_;
  wire lo074_buf_o2_p_spl_;
  wire lo074_buf_o2_p_spl_0;
  wire lo090_buf_o2_n_spl_;
  wire lo074_buf_o2_n_spl_;
  wire lo090_buf_o2_p_spl_;
  wire lo090_buf_o2_p_spl_0;
  wire lo106_buf_o2_p_spl_;
  wire lo106_buf_o2_p_spl_0;
  wire lo122_buf_o2_n_spl_;
  wire lo106_buf_o2_n_spl_;
  wire lo122_buf_o2_p_spl_;
  wire lo122_buf_o2_p_spl_0;
  wire g529_n_spl_;
  wire g536_p_spl_;
  wire lo078_buf_o2_p_spl_;
  wire lo078_buf_o2_p_spl_0;
  wire lo094_buf_o2_n_spl_;
  wire lo078_buf_o2_n_spl_;
  wire lo094_buf_o2_p_spl_;
  wire lo094_buf_o2_p_spl_0;
  wire lo110_buf_o2_p_spl_;
  wire lo110_buf_o2_p_spl_0;
  wire lo126_buf_o2_n_spl_;
  wire lo110_buf_o2_n_spl_;
  wire lo126_buf_o2_p_spl_;
  wire lo126_buf_o2_p_spl_0;
  wire g547_n_spl_;
  wire g554_p_spl_;
  wire lo001_buf_o2_p_spl_;
  wire lo001_buf_o2_p_spl_0;
  wire lo005_buf_o2_n_spl_;
  wire lo001_buf_o2_n_spl_;
  wire lo005_buf_o2_p_spl_;
  wire lo005_buf_o2_p_spl_0;
  wire lo009_buf_o2_p_spl_;
  wire lo009_buf_o2_p_spl_0;
  wire lo013_buf_o2_n_spl_;
  wire lo009_buf_o2_n_spl_;
  wire lo013_buf_o2_p_spl_;
  wire lo013_buf_o2_p_spl_0;
  wire lo017_buf_o2_p_spl_;
  wire lo017_buf_o2_p_spl_0;
  wire lo021_buf_o2_n_spl_;
  wire lo017_buf_o2_n_spl_;
  wire lo021_buf_o2_p_spl_;
  wire lo021_buf_o2_p_spl_0;
  wire lo025_buf_o2_p_spl_;
  wire lo025_buf_o2_p_spl_0;
  wire lo029_buf_o2_n_spl_;
  wire lo025_buf_o2_n_spl_;
  wire lo029_buf_o2_p_spl_;
  wire lo029_buf_o2_p_spl_0;
  wire lo033_buf_o2_p_spl_;
  wire lo033_buf_o2_p_spl_0;
  wire lo037_buf_o2_n_spl_;
  wire lo033_buf_o2_n_spl_;
  wire lo037_buf_o2_p_spl_;
  wire lo037_buf_o2_p_spl_0;
  wire lo041_buf_o2_p_spl_;
  wire lo041_buf_o2_p_spl_0;
  wire lo045_buf_o2_n_spl_;
  wire lo041_buf_o2_n_spl_;
  wire lo045_buf_o2_p_spl_;
  wire lo045_buf_o2_p_spl_0;
  wire lo049_buf_o2_p_spl_;
  wire lo049_buf_o2_p_spl_0;
  wire lo053_buf_o2_n_spl_;
  wire lo049_buf_o2_n_spl_;
  wire lo053_buf_o2_p_spl_;
  wire lo053_buf_o2_p_spl_0;
  wire lo057_buf_o2_p_spl_;
  wire lo057_buf_o2_p_spl_0;
  wire lo061_buf_o2_n_spl_;
  wire lo057_buf_o2_n_spl_;
  wire lo061_buf_o2_p_spl_;
  wire lo061_buf_o2_p_spl_0;
  wire lo065_buf_o2_p_spl_;
  wire lo065_buf_o2_p_spl_0;
  wire lo069_buf_o2_n_spl_;
  wire lo065_buf_o2_n_spl_;
  wire lo069_buf_o2_p_spl_;
  wire lo069_buf_o2_p_spl_0;
  wire lo073_buf_o2_p_spl_;
  wire lo073_buf_o2_p_spl_0;
  wire lo077_buf_o2_n_spl_;
  wire lo073_buf_o2_n_spl_;
  wire lo077_buf_o2_p_spl_;
  wire lo077_buf_o2_p_spl_0;
  wire lo081_buf_o2_p_spl_;
  wire lo081_buf_o2_p_spl_0;
  wire lo085_buf_o2_n_spl_;
  wire lo081_buf_o2_n_spl_;
  wire lo085_buf_o2_p_spl_;
  wire lo085_buf_o2_p_spl_0;
  wire lo089_buf_o2_p_spl_;
  wire lo089_buf_o2_p_spl_0;
  wire lo093_buf_o2_n_spl_;
  wire lo089_buf_o2_n_spl_;
  wire lo093_buf_o2_p_spl_;
  wire lo093_buf_o2_p_spl_0;
  wire lo097_buf_o2_p_spl_;
  wire lo097_buf_o2_p_spl_0;
  wire lo101_buf_o2_n_spl_;
  wire lo097_buf_o2_n_spl_;
  wire lo101_buf_o2_p_spl_;
  wire lo101_buf_o2_p_spl_0;
  wire lo105_buf_o2_p_spl_;
  wire lo105_buf_o2_p_spl_0;
  wire lo109_buf_o2_n_spl_;
  wire lo105_buf_o2_n_spl_;
  wire lo109_buf_o2_p_spl_;
  wire lo109_buf_o2_p_spl_0;
  wire lo113_buf_o2_p_spl_;
  wire lo113_buf_o2_p_spl_0;
  wire lo117_buf_o2_n_spl_;
  wire lo113_buf_o2_n_spl_;
  wire lo117_buf_o2_p_spl_;
  wire lo117_buf_o2_p_spl_0;
  wire lo121_buf_o2_p_spl_;
  wire lo121_buf_o2_p_spl_0;
  wire lo125_buf_o2_n_spl_;
  wire lo121_buf_o2_n_spl_;
  wire lo125_buf_o2_p_spl_;
  wire lo125_buf_o2_p_spl_0;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  buf

  (
    n286_lo_p,
    n286_lo
  );


  not

  (
    n286_lo_n,
    n286_lo
  );


  buf

  (
    n298_lo_p,
    n298_lo
  );


  not

  (
    n298_lo_n,
    n298_lo
  );


  buf

  (
    n310_lo_p,
    n310_lo
  );


  not

  (
    n310_lo_n,
    n310_lo
  );


  buf

  (
    n322_lo_p,
    n322_lo
  );


  not

  (
    n322_lo_n,
    n322_lo
  );


  buf

  (
    n334_lo_p,
    n334_lo
  );


  not

  (
    n334_lo_n,
    n334_lo
  );


  buf

  (
    n346_lo_p,
    n346_lo
  );


  not

  (
    n346_lo_n,
    n346_lo
  );


  buf

  (
    n358_lo_p,
    n358_lo
  );


  not

  (
    n358_lo_n,
    n358_lo
  );


  buf

  (
    n370_lo_p,
    n370_lo
  );


  not

  (
    n370_lo_n,
    n370_lo
  );


  buf

  (
    n382_lo_p,
    n382_lo
  );


  not

  (
    n382_lo_n,
    n382_lo
  );


  buf

  (
    n394_lo_p,
    n394_lo
  );


  not

  (
    n394_lo_n,
    n394_lo
  );


  buf

  (
    n406_lo_p,
    n406_lo
  );


  not

  (
    n406_lo_n,
    n406_lo
  );


  buf

  (
    n418_lo_p,
    n418_lo
  );


  not

  (
    n418_lo_n,
    n418_lo
  );


  buf

  (
    n430_lo_p,
    n430_lo
  );


  not

  (
    n430_lo_n,
    n430_lo
  );


  buf

  (
    n442_lo_p,
    n442_lo
  );


  not

  (
    n442_lo_n,
    n442_lo
  );


  buf

  (
    n454_lo_p,
    n454_lo
  );


  not

  (
    n454_lo_n,
    n454_lo
  );


  buf

  (
    n466_lo_p,
    n466_lo
  );


  not

  (
    n466_lo_n,
    n466_lo
  );


  buf

  (
    n478_lo_p,
    n478_lo
  );


  not

  (
    n478_lo_n,
    n478_lo
  );


  buf

  (
    n490_lo_p,
    n490_lo
  );


  not

  (
    n490_lo_n,
    n490_lo
  );


  buf

  (
    n502_lo_p,
    n502_lo
  );


  not

  (
    n502_lo_n,
    n502_lo
  );


  buf

  (
    n514_lo_p,
    n514_lo
  );


  not

  (
    n514_lo_n,
    n514_lo
  );


  buf

  (
    n526_lo_p,
    n526_lo
  );


  not

  (
    n526_lo_n,
    n526_lo
  );


  buf

  (
    n538_lo_p,
    n538_lo
  );


  not

  (
    n538_lo_n,
    n538_lo
  );


  buf

  (
    n550_lo_p,
    n550_lo
  );


  not

  (
    n550_lo_n,
    n550_lo
  );


  buf

  (
    n562_lo_p,
    n562_lo
  );


  not

  (
    n562_lo_n,
    n562_lo
  );


  buf

  (
    n574_lo_p,
    n574_lo
  );


  not

  (
    n574_lo_n,
    n574_lo
  );


  buf

  (
    n586_lo_p,
    n586_lo
  );


  not

  (
    n586_lo_n,
    n586_lo
  );


  buf

  (
    n598_lo_p,
    n598_lo
  );


  not

  (
    n598_lo_n,
    n598_lo
  );


  buf

  (
    n610_lo_p,
    n610_lo
  );


  not

  (
    n610_lo_n,
    n610_lo
  );


  buf

  (
    n622_lo_p,
    n622_lo
  );


  not

  (
    n622_lo_n,
    n622_lo
  );


  buf

  (
    n634_lo_p,
    n634_lo
  );


  not

  (
    n634_lo_n,
    n634_lo
  );


  buf

  (
    n646_lo_p,
    n646_lo
  );


  not

  (
    n646_lo_n,
    n646_lo
  );


  buf

  (
    n658_lo_p,
    n658_lo
  );


  not

  (
    n658_lo_n,
    n658_lo
  );


  buf

  (
    n661_lo_p,
    n661_lo
  );


  not

  (
    n661_lo_n,
    n661_lo
  );


  buf

  (
    n673_lo_p,
    n673_lo
  );


  not

  (
    n673_lo_n,
    n673_lo
  );


  buf

  (
    n685_lo_p,
    n685_lo
  );


  not

  (
    n685_lo_n,
    n685_lo
  );


  buf

  (
    n697_lo_p,
    n697_lo
  );


  not

  (
    n697_lo_n,
    n697_lo
  );


  buf

  (
    n709_lo_p,
    n709_lo
  );


  not

  (
    n709_lo_n,
    n709_lo
  );


  buf

  (
    n721_lo_p,
    n721_lo
  );


  not

  (
    n721_lo_n,
    n721_lo
  );


  buf

  (
    n733_lo_p,
    n733_lo
  );


  not

  (
    n733_lo_n,
    n733_lo
  );


  buf

  (
    n745_lo_p,
    n745_lo
  );


  not

  (
    n745_lo_n,
    n745_lo
  );


  buf

  (
    n757_lo_p,
    n757_lo
  );


  not

  (
    n757_lo_n,
    n757_lo
  );


  buf

  (
    n1589_o2_p,
    n1589_o2
  );


  not

  (
    n1589_o2_n,
    n1589_o2
  );


  buf

  (
    n1590_o2_p,
    n1590_o2
  );


  not

  (
    n1590_o2_n,
    n1590_o2
  );


  buf

  (
    n1591_o2_p,
    n1591_o2
  );


  not

  (
    n1591_o2_n,
    n1591_o2
  );


  buf

  (
    n1592_o2_p,
    n1592_o2
  );


  not

  (
    n1592_o2_n,
    n1592_o2
  );


  buf

  (
    n1593_o2_p,
    n1593_o2
  );


  not

  (
    n1593_o2_n,
    n1593_o2
  );


  buf

  (
    n1594_o2_p,
    n1594_o2
  );


  not

  (
    n1594_o2_n,
    n1594_o2
  );


  buf

  (
    n1595_o2_p,
    n1595_o2
  );


  not

  (
    n1595_o2_n,
    n1595_o2
  );


  buf

  (
    n1596_o2_p,
    n1596_o2
  );


  not

  (
    n1596_o2_n,
    n1596_o2
  );


  buf

  (
    n1597_o2_p,
    n1597_o2
  );


  not

  (
    n1597_o2_n,
    n1597_o2
  );


  buf

  (
    n1598_o2_p,
    n1598_o2
  );


  not

  (
    n1598_o2_n,
    n1598_o2
  );


  buf

  (
    n1599_o2_p,
    n1599_o2
  );


  not

  (
    n1599_o2_n,
    n1599_o2
  );


  buf

  (
    n1600_o2_p,
    n1600_o2
  );


  not

  (
    n1600_o2_n,
    n1600_o2
  );


  buf

  (
    n1601_o2_p,
    n1601_o2
  );


  not

  (
    n1601_o2_n,
    n1601_o2
  );


  buf

  (
    n1602_o2_p,
    n1602_o2
  );


  not

  (
    n1602_o2_n,
    n1602_o2
  );


  buf

  (
    n1603_o2_p,
    n1603_o2
  );


  not

  (
    n1603_o2_n,
    n1603_o2
  );


  buf

  (
    n1604_o2_p,
    n1604_o2
  );


  not

  (
    n1604_o2_n,
    n1604_o2
  );


  buf

  (
    n1605_o2_p,
    n1605_o2
  );


  not

  (
    n1605_o2_n,
    n1605_o2
  );


  buf

  (
    n1606_o2_p,
    n1606_o2
  );


  not

  (
    n1606_o2_n,
    n1606_o2
  );


  buf

  (
    n1607_o2_p,
    n1607_o2
  );


  not

  (
    n1607_o2_n,
    n1607_o2
  );


  buf

  (
    n1608_o2_p,
    n1608_o2
  );


  not

  (
    n1608_o2_n,
    n1608_o2
  );


  buf

  (
    n1609_o2_p,
    n1609_o2
  );


  not

  (
    n1609_o2_n,
    n1609_o2
  );


  buf

  (
    n1610_o2_p,
    n1610_o2
  );


  not

  (
    n1610_o2_n,
    n1610_o2
  );


  buf

  (
    n1611_o2_p,
    n1611_o2
  );


  not

  (
    n1611_o2_n,
    n1611_o2
  );


  buf

  (
    n1612_o2_p,
    n1612_o2
  );


  not

  (
    n1612_o2_n,
    n1612_o2
  );


  buf

  (
    n1613_o2_p,
    n1613_o2
  );


  not

  (
    n1613_o2_n,
    n1613_o2
  );


  buf

  (
    n1614_o2_p,
    n1614_o2
  );


  not

  (
    n1614_o2_n,
    n1614_o2
  );


  buf

  (
    n1615_o2_p,
    n1615_o2
  );


  not

  (
    n1615_o2_n,
    n1615_o2
  );


  buf

  (
    n1616_o2_p,
    n1616_o2
  );


  not

  (
    n1616_o2_n,
    n1616_o2
  );


  buf

  (
    n1617_o2_p,
    n1617_o2
  );


  not

  (
    n1617_o2_n,
    n1617_o2
  );


  buf

  (
    n1618_o2_p,
    n1618_o2
  );


  not

  (
    n1618_o2_n,
    n1618_o2
  );


  buf

  (
    n1619_o2_p,
    n1619_o2
  );


  not

  (
    n1619_o2_n,
    n1619_o2
  );


  buf

  (
    n1620_o2_p,
    n1620_o2
  );


  not

  (
    n1620_o2_n,
    n1620_o2
  );


  buf

  (
    n602_o2_p,
    n602_o2
  );


  not

  (
    n602_o2_n,
    n602_o2
  );


  buf

  (
    n639_o2_p,
    n639_o2
  );


  not

  (
    n639_o2_n,
    n639_o2
  );


  buf

  (
    n678_o2_p,
    n678_o2
  );


  not

  (
    n678_o2_n,
    n678_o2
  );


  buf

  (
    n658_o2_p,
    n658_o2
  );


  not

  (
    n658_o2_n,
    n658_o2
  );


  buf

  (
    n783_o2_p,
    n783_o2
  );


  not

  (
    n783_o2_n,
    n783_o2
  );


  buf

  (
    n802_o2_p,
    n802_o2
  );


  not

  (
    n802_o2_n,
    n802_o2
  );


  buf

  (
    n726_o2_p,
    n726_o2
  );


  not

  (
    n726_o2_n,
    n726_o2
  );


  buf

  (
    n763_o2_p,
    n763_o2
  );


  not

  (
    n763_o2_n,
    n763_o2
  );


  buf

  (
    n685_o2_p,
    n685_o2
  );


  not

  (
    n685_o2_n,
    n685_o2
  );


  buf

  (
    n680_o2_p,
    n680_o2
  );


  not

  (
    n680_o2_n,
    n680_o2
  );


  buf

  (
    n822_o2_p,
    n822_o2
  );


  not

  (
    n822_o2_n,
    n822_o2
  );


  buf

  (
    n843_o2_p,
    n843_o2
  );


  not

  (
    n843_o2_n,
    n843_o2
  );


  buf

  (
    n842_o2_p,
    n842_o2
  );


  not

  (
    n842_o2_n,
    n842_o2
  );


  buf

  (
    n681_o2_p,
    n681_o2
  );


  not

  (
    n681_o2_n,
    n681_o2
  );


  buf

  (
    n684_o2_p,
    n684_o2
  );


  not

  (
    n684_o2_n,
    n684_o2
  );


  buf

  (
    n686_o2_p,
    n686_o2
  );


  not

  (
    n686_o2_n,
    n686_o2
  );


  buf

  (
    n823_o2_p,
    n823_o2
  );


  not

  (
    n823_o2_n,
    n823_o2
  );


  buf

  (
    lo002_buf_o2_p,
    lo002_buf_o2
  );


  not

  (
    lo002_buf_o2_n,
    lo002_buf_o2
  );


  buf

  (
    lo006_buf_o2_p,
    lo006_buf_o2
  );


  not

  (
    lo006_buf_o2_n,
    lo006_buf_o2
  );


  buf

  (
    lo010_buf_o2_p,
    lo010_buf_o2
  );


  not

  (
    lo010_buf_o2_n,
    lo010_buf_o2
  );


  buf

  (
    lo014_buf_o2_p,
    lo014_buf_o2
  );


  not

  (
    lo014_buf_o2_n,
    lo014_buf_o2
  );


  buf

  (
    lo018_buf_o2_p,
    lo018_buf_o2
  );


  not

  (
    lo018_buf_o2_n,
    lo018_buf_o2
  );


  buf

  (
    lo022_buf_o2_p,
    lo022_buf_o2
  );


  not

  (
    lo022_buf_o2_n,
    lo022_buf_o2
  );


  buf

  (
    lo026_buf_o2_p,
    lo026_buf_o2
  );


  not

  (
    lo026_buf_o2_n,
    lo026_buf_o2
  );


  buf

  (
    lo030_buf_o2_p,
    lo030_buf_o2
  );


  not

  (
    lo030_buf_o2_n,
    lo030_buf_o2
  );


  buf

  (
    lo034_buf_o2_p,
    lo034_buf_o2
  );


  not

  (
    lo034_buf_o2_n,
    lo034_buf_o2
  );


  buf

  (
    lo038_buf_o2_p,
    lo038_buf_o2
  );


  not

  (
    lo038_buf_o2_n,
    lo038_buf_o2
  );


  buf

  (
    lo042_buf_o2_p,
    lo042_buf_o2
  );


  not

  (
    lo042_buf_o2_n,
    lo042_buf_o2
  );


  buf

  (
    lo046_buf_o2_p,
    lo046_buf_o2
  );


  not

  (
    lo046_buf_o2_n,
    lo046_buf_o2
  );


  buf

  (
    lo050_buf_o2_p,
    lo050_buf_o2
  );


  not

  (
    lo050_buf_o2_n,
    lo050_buf_o2
  );


  buf

  (
    lo054_buf_o2_p,
    lo054_buf_o2
  );


  not

  (
    lo054_buf_o2_n,
    lo054_buf_o2
  );


  buf

  (
    lo058_buf_o2_p,
    lo058_buf_o2
  );


  not

  (
    lo058_buf_o2_n,
    lo058_buf_o2
  );


  buf

  (
    lo062_buf_o2_p,
    lo062_buf_o2
  );


  not

  (
    lo062_buf_o2_n,
    lo062_buf_o2
  );


  buf

  (
    lo066_buf_o2_p,
    lo066_buf_o2
  );


  not

  (
    lo066_buf_o2_n,
    lo066_buf_o2
  );


  buf

  (
    lo070_buf_o2_p,
    lo070_buf_o2
  );


  not

  (
    lo070_buf_o2_n,
    lo070_buf_o2
  );


  buf

  (
    lo074_buf_o2_p,
    lo074_buf_o2
  );


  not

  (
    lo074_buf_o2_n,
    lo074_buf_o2
  );


  buf

  (
    lo078_buf_o2_p,
    lo078_buf_o2
  );


  not

  (
    lo078_buf_o2_n,
    lo078_buf_o2
  );


  buf

  (
    lo082_buf_o2_p,
    lo082_buf_o2
  );


  not

  (
    lo082_buf_o2_n,
    lo082_buf_o2
  );


  buf

  (
    lo086_buf_o2_p,
    lo086_buf_o2
  );


  not

  (
    lo086_buf_o2_n,
    lo086_buf_o2
  );


  buf

  (
    lo090_buf_o2_p,
    lo090_buf_o2
  );


  not

  (
    lo090_buf_o2_n,
    lo090_buf_o2
  );


  buf

  (
    lo094_buf_o2_p,
    lo094_buf_o2
  );


  not

  (
    lo094_buf_o2_n,
    lo094_buf_o2
  );


  buf

  (
    lo098_buf_o2_p,
    lo098_buf_o2
  );


  not

  (
    lo098_buf_o2_n,
    lo098_buf_o2
  );


  buf

  (
    lo102_buf_o2_p,
    lo102_buf_o2
  );


  not

  (
    lo102_buf_o2_n,
    lo102_buf_o2
  );


  buf

  (
    lo106_buf_o2_p,
    lo106_buf_o2
  );


  not

  (
    lo106_buf_o2_n,
    lo106_buf_o2
  );


  buf

  (
    lo110_buf_o2_p,
    lo110_buf_o2
  );


  not

  (
    lo110_buf_o2_n,
    lo110_buf_o2
  );


  buf

  (
    lo114_buf_o2_p,
    lo114_buf_o2
  );


  not

  (
    lo114_buf_o2_n,
    lo114_buf_o2
  );


  buf

  (
    lo118_buf_o2_p,
    lo118_buf_o2
  );


  not

  (
    lo118_buf_o2_n,
    lo118_buf_o2
  );


  buf

  (
    lo122_buf_o2_p,
    lo122_buf_o2
  );


  not

  (
    lo122_buf_o2_n,
    lo122_buf_o2
  );


  buf

  (
    lo126_buf_o2_p,
    lo126_buf_o2
  );


  not

  (
    lo126_buf_o2_n,
    lo126_buf_o2
  );


  buf

  (
    n683_o2_p,
    n683_o2
  );


  not

  (
    n683_o2_n,
    n683_o2
  );


  buf

  (
    n688_o2_p,
    n688_o2
  );


  not

  (
    n688_o2_n,
    n688_o2
  );


  buf

  (
    n803_o2_p,
    n803_o2
  );


  not

  (
    n803_o2_n,
    n803_o2
  );


  buf

  (
    n862_o2_p,
    n862_o2
  );


  not

  (
    n862_o2_n,
    n862_o2
  );


  buf

  (
    n764_o2_p,
    n764_o2
  );


  not

  (
    n764_o2_n,
    n764_o2
  );


  buf

  (
    n863_o2_p,
    n863_o2
  );


  not

  (
    n863_o2_n,
    n863_o2
  );


  buf

  (
    n886_o2_p,
    n886_o2
  );


  not

  (
    n886_o2_n,
    n886_o2
  );


  buf

  (
    n600_o2_p,
    n600_o2
  );


  not

  (
    n600_o2_n,
    n600_o2
  );


  buf

  (
    n601_o2_p,
    n601_o2
  );


  not

  (
    n601_o2_n,
    n601_o2
  );


  buf

  (
    n637_o2_p,
    n637_o2
  );


  not

  (
    n637_o2_n,
    n637_o2
  );


  buf

  (
    n638_o2_p,
    n638_o2
  );


  not

  (
    n638_o2_n,
    n638_o2
  );


  buf

  (
    n676_o2_p,
    n676_o2
  );


  not

  (
    n676_o2_n,
    n676_o2
  );


  buf

  (
    n677_o2_p,
    n677_o2
  );


  not

  (
    n677_o2_n,
    n677_o2
  );


  buf

  (
    n656_o2_p,
    n656_o2
  );


  not

  (
    n656_o2_n,
    n656_o2
  );


  buf

  (
    n657_o2_p,
    n657_o2
  );


  not

  (
    n657_o2_n,
    n657_o2
  );


  buf

  (
    n781_o2_p,
    n781_o2
  );


  not

  (
    n781_o2_n,
    n781_o2
  );


  buf

  (
    n782_o2_p,
    n782_o2
  );


  not

  (
    n782_o2_n,
    n782_o2
  );


  buf

  (
    n800_o2_p,
    n800_o2
  );


  not

  (
    n800_o2_n,
    n800_o2
  );


  buf

  (
    n801_o2_p,
    n801_o2
  );


  not

  (
    n801_o2_n,
    n801_o2
  );


  buf

  (
    n724_o2_p,
    n724_o2
  );


  not

  (
    n724_o2_n,
    n724_o2
  );


  buf

  (
    n725_o2_p,
    n725_o2
  );


  not

  (
    n725_o2_n,
    n725_o2
  );


  buf

  (
    n761_o2_p,
    n761_o2
  );


  not

  (
    n761_o2_n,
    n761_o2
  );


  buf

  (
    n762_o2_p,
    n762_o2
  );


  not

  (
    n762_o2_n,
    n762_o2
  );


  buf

  (
    lo129_buf_o2_p,
    lo129_buf_o2
  );


  not

  (
    lo129_buf_o2_n,
    lo129_buf_o2
  );


  buf

  (
    lo133_buf_o2_p,
    lo133_buf_o2
  );


  not

  (
    lo133_buf_o2_n,
    lo133_buf_o2
  );


  buf

  (
    lo137_buf_o2_p,
    lo137_buf_o2
  );


  not

  (
    lo137_buf_o2_n,
    lo137_buf_o2
  );


  buf

  (
    lo141_buf_o2_p,
    lo141_buf_o2
  );


  not

  (
    lo141_buf_o2_n,
    lo141_buf_o2
  );


  buf

  (
    lo145_buf_o2_p,
    lo145_buf_o2
  );


  not

  (
    lo145_buf_o2_n,
    lo145_buf_o2
  );


  buf

  (
    lo149_buf_o2_p,
    lo149_buf_o2
  );


  not

  (
    lo149_buf_o2_n,
    lo149_buf_o2
  );


  buf

  (
    lo153_buf_o2_p,
    lo153_buf_o2
  );


  not

  (
    lo153_buf_o2_n,
    lo153_buf_o2
  );


  buf

  (
    lo157_buf_o2_p,
    lo157_buf_o2
  );


  not

  (
    lo157_buf_o2_n,
    lo157_buf_o2
  );


  buf

  (
    lo161_buf_o2_p,
    lo161_buf_o2
  );


  not

  (
    lo161_buf_o2_n,
    lo161_buf_o2
  );


  buf

  (
    n708_o2_p,
    n708_o2
  );


  not

  (
    n708_o2_n,
    n708_o2
  );


  buf

  (
    n745_o2_p,
    n745_o2
  );


  not

  (
    n745_o2_n,
    n745_o2
  );


  buf

  (
    n717_o2_p,
    n717_o2
  );


  not

  (
    n717_o2_n,
    n717_o2
  );


  buf

  (
    n754_o2_p,
    n754_o2
  );


  not

  (
    n754_o2_n,
    n754_o2
  );


  buf

  (
    n584_o2_p,
    n584_o2
  );


  not

  (
    n584_o2_n,
    n584_o2
  );


  buf

  (
    n593_o2_p,
    n593_o2
  );


  not

  (
    n593_o2_n,
    n593_o2
  );


  buf

  (
    n630_o2_p,
    n630_o2
  );


  not

  (
    n630_o2_n,
    n630_o2
  );


  buf

  (
    n621_o2_p,
    n621_o2
  );


  not

  (
    n621_o2_n,
    n621_o2
  );


  buf

  (
    lo001_buf_o2_p,
    lo001_buf_o2
  );


  not

  (
    lo001_buf_o2_n,
    lo001_buf_o2
  );


  buf

  (
    lo005_buf_o2_p,
    lo005_buf_o2
  );


  not

  (
    lo005_buf_o2_n,
    lo005_buf_o2
  );


  buf

  (
    lo009_buf_o2_p,
    lo009_buf_o2
  );


  not

  (
    lo009_buf_o2_n,
    lo009_buf_o2
  );


  buf

  (
    lo013_buf_o2_p,
    lo013_buf_o2
  );


  not

  (
    lo013_buf_o2_n,
    lo013_buf_o2
  );


  buf

  (
    lo017_buf_o2_p,
    lo017_buf_o2
  );


  not

  (
    lo017_buf_o2_n,
    lo017_buf_o2
  );


  buf

  (
    lo021_buf_o2_p,
    lo021_buf_o2
  );


  not

  (
    lo021_buf_o2_n,
    lo021_buf_o2
  );


  buf

  (
    lo025_buf_o2_p,
    lo025_buf_o2
  );


  not

  (
    lo025_buf_o2_n,
    lo025_buf_o2
  );


  buf

  (
    lo029_buf_o2_p,
    lo029_buf_o2
  );


  not

  (
    lo029_buf_o2_n,
    lo029_buf_o2
  );


  buf

  (
    lo033_buf_o2_p,
    lo033_buf_o2
  );


  not

  (
    lo033_buf_o2_n,
    lo033_buf_o2
  );


  buf

  (
    lo037_buf_o2_p,
    lo037_buf_o2
  );


  not

  (
    lo037_buf_o2_n,
    lo037_buf_o2
  );


  buf

  (
    lo041_buf_o2_p,
    lo041_buf_o2
  );


  not

  (
    lo041_buf_o2_n,
    lo041_buf_o2
  );


  buf

  (
    lo045_buf_o2_p,
    lo045_buf_o2
  );


  not

  (
    lo045_buf_o2_n,
    lo045_buf_o2
  );


  buf

  (
    lo049_buf_o2_p,
    lo049_buf_o2
  );


  not

  (
    lo049_buf_o2_n,
    lo049_buf_o2
  );


  buf

  (
    lo053_buf_o2_p,
    lo053_buf_o2
  );


  not

  (
    lo053_buf_o2_n,
    lo053_buf_o2
  );


  buf

  (
    lo057_buf_o2_p,
    lo057_buf_o2
  );


  not

  (
    lo057_buf_o2_n,
    lo057_buf_o2
  );


  buf

  (
    lo061_buf_o2_p,
    lo061_buf_o2
  );


  not

  (
    lo061_buf_o2_n,
    lo061_buf_o2
  );


  buf

  (
    lo065_buf_o2_p,
    lo065_buf_o2
  );


  not

  (
    lo065_buf_o2_n,
    lo065_buf_o2
  );


  buf

  (
    lo069_buf_o2_p,
    lo069_buf_o2
  );


  not

  (
    lo069_buf_o2_n,
    lo069_buf_o2
  );


  buf

  (
    lo073_buf_o2_p,
    lo073_buf_o2
  );


  not

  (
    lo073_buf_o2_n,
    lo073_buf_o2
  );


  buf

  (
    lo077_buf_o2_p,
    lo077_buf_o2
  );


  not

  (
    lo077_buf_o2_n,
    lo077_buf_o2
  );


  buf

  (
    lo081_buf_o2_p,
    lo081_buf_o2
  );


  not

  (
    lo081_buf_o2_n,
    lo081_buf_o2
  );


  buf

  (
    lo085_buf_o2_p,
    lo085_buf_o2
  );


  not

  (
    lo085_buf_o2_n,
    lo085_buf_o2
  );


  buf

  (
    lo089_buf_o2_p,
    lo089_buf_o2
  );


  not

  (
    lo089_buf_o2_n,
    lo089_buf_o2
  );


  buf

  (
    lo093_buf_o2_p,
    lo093_buf_o2
  );


  not

  (
    lo093_buf_o2_n,
    lo093_buf_o2
  );


  buf

  (
    lo097_buf_o2_p,
    lo097_buf_o2
  );


  not

  (
    lo097_buf_o2_n,
    lo097_buf_o2
  );


  buf

  (
    lo101_buf_o2_p,
    lo101_buf_o2
  );


  not

  (
    lo101_buf_o2_n,
    lo101_buf_o2
  );


  buf

  (
    lo105_buf_o2_p,
    lo105_buf_o2
  );


  not

  (
    lo105_buf_o2_n,
    lo105_buf_o2
  );


  buf

  (
    lo109_buf_o2_p,
    lo109_buf_o2
  );


  not

  (
    lo109_buf_o2_n,
    lo109_buf_o2
  );


  buf

  (
    lo113_buf_o2_p,
    lo113_buf_o2
  );


  not

  (
    lo113_buf_o2_n,
    lo113_buf_o2
  );


  buf

  (
    lo117_buf_o2_p,
    lo117_buf_o2
  );


  not

  (
    lo117_buf_o2_n,
    lo117_buf_o2
  );


  buf

  (
    lo121_buf_o2_p,
    lo121_buf_o2
  );


  not

  (
    lo121_buf_o2_n,
    lo121_buf_o2
  );


  buf

  (
    lo125_buf_o2_p,
    lo125_buf_o2
  );


  not

  (
    lo125_buf_o2_n,
    lo125_buf_o2
  );


  and

  (
    g236_p,
    n683_o2_n,
    n688_o2_n
  );


  or

  (
    g236_n,
    n683_o2_p,
    n688_o2_p
  );


  and

  (
    g237_p,
    n803_o2_p,
    n764_o2_p
  );


  or

  (
    g237_n,
    n803_o2_n,
    n764_o2_n
  );


  and

  (
    g238_p,
    g236_n_spl_0,
    g237_p
  );


  or

  (
    g238_n,
    g236_p_spl_0,
    g237_n
  );


  and

  (
    g239_p,
    n602_o2_p_spl_0,
    g238_p_spl_0
  );


  or

  (
    g239_n,
    n602_o2_n_spl_0,
    g238_n_spl_0
  );


  and

  (
    g240_p,
    n286_lo_n,
    g239_p
  );


  and

  (
    g241_p,
    n286_lo_p,
    g239_n
  );


  or

  (
    g242_n,
    g240_p,
    g241_p
  );


  and

  (
    g243_p,
    n639_o2_p_spl_00,
    g238_p_spl_0
  );


  or

  (
    g243_n,
    n639_o2_n_spl_00,
    g238_n_spl_0
  );


  and

  (
    g244_p,
    n298_lo_n,
    g243_p
  );


  and

  (
    g245_p,
    n298_lo_p,
    g243_n
  );


  or

  (
    g246_n,
    g244_p,
    g245_p
  );


  and

  (
    g247_p,
    n678_o2_p_spl_00,
    g238_p_spl_1
  );


  or

  (
    g247_n,
    n678_o2_n_spl_00,
    g238_n_spl_1
  );


  and

  (
    g248_p,
    n310_lo_n,
    g247_p
  );


  and

  (
    g249_p,
    n310_lo_p,
    g247_n
  );


  or

  (
    g250_n,
    g248_p,
    g249_p
  );


  and

  (
    g251_p,
    n658_o2_p_spl_0,
    g238_p_spl_1
  );


  or

  (
    g251_n,
    n658_o2_n_spl_0,
    g238_n_spl_1
  );


  and

  (
    g252_p,
    n322_lo_n,
    g251_p
  );


  and

  (
    g253_p,
    n322_lo_p,
    g251_n
  );


  or

  (
    g254_n,
    g252_p,
    g253_p
  );


  and

  (
    g255_p,
    n822_o2_p,
    n823_o2_n
  );


  or

  (
    g255_n,
    n822_o2_n,
    n823_o2_p
  );


  and

  (
    g256_p,
    g236_n_spl_0,
    g255_p
  );


  or

  (
    g256_n,
    g236_p_spl_0,
    g255_n
  );


  and

  (
    g257_p,
    n602_o2_p_spl_0,
    g256_p_spl_0
  );


  or

  (
    g257_n,
    n602_o2_n_spl_0,
    g256_n_spl_0
  );


  and

  (
    g258_p,
    n334_lo_n,
    g257_p
  );


  and

  (
    g259_p,
    n334_lo_p,
    g257_n
  );


  or

  (
    g260_n,
    g258_p,
    g259_p
  );


  and

  (
    g261_p,
    n639_o2_p_spl_00,
    g256_p_spl_0
  );


  or

  (
    g261_n,
    n639_o2_n_spl_00,
    g256_n_spl_0
  );


  and

  (
    g262_p,
    n346_lo_n,
    g261_p
  );


  and

  (
    g263_p,
    n346_lo_p,
    g261_n
  );


  or

  (
    g264_n,
    g262_p,
    g263_p
  );


  and

  (
    g265_p,
    n678_o2_p_spl_00,
    g256_p_spl_1
  );


  or

  (
    g265_n,
    n678_o2_n_spl_00,
    g256_n_spl_1
  );


  and

  (
    g266_p,
    n358_lo_n,
    g265_p
  );


  and

  (
    g267_p,
    n358_lo_p,
    g265_n
  );


  or

  (
    g268_n,
    g266_p,
    g267_p
  );


  and

  (
    g269_p,
    n658_o2_p_spl_0,
    g256_p_spl_1
  );


  or

  (
    g269_n,
    n658_o2_n_spl_0,
    g256_n_spl_1
  );


  and

  (
    g270_p,
    n370_lo_n,
    g269_p
  );


  and

  (
    g271_p,
    n370_lo_p,
    g269_n
  );


  or

  (
    g272_n,
    g270_p,
    g271_p
  );


  and

  (
    g273_p,
    n843_o2_n,
    n842_o2_p
  );


  or

  (
    g273_n,
    n843_o2_p,
    n842_o2_n
  );


  and

  (
    g274_p,
    g236_n_spl_1,
    g273_p
  );


  or

  (
    g274_n,
    g236_p_spl_1,
    g273_n
  );


  and

  (
    g275_p,
    n602_o2_p_spl_1,
    g274_p_spl_0
  );


  or

  (
    g275_n,
    n602_o2_n_spl_1,
    g274_n_spl_0
  );


  and

  (
    g276_p,
    n382_lo_n,
    g275_p
  );


  and

  (
    g277_p,
    n382_lo_p,
    g275_n
  );


  or

  (
    g278_n,
    g276_p,
    g277_p
  );


  and

  (
    g279_p,
    n639_o2_p_spl_0,
    g274_p_spl_0
  );


  or

  (
    g279_n,
    n639_o2_n_spl_0,
    g274_n_spl_0
  );


  and

  (
    g280_p,
    n394_lo_n,
    g279_p
  );


  and

  (
    g281_p,
    n394_lo_p,
    g279_n
  );


  or

  (
    g282_n,
    g280_p,
    g281_p
  );


  and

  (
    g283_p,
    n678_o2_p_spl_01,
    g274_p_spl_1
  );


  or

  (
    g283_n,
    n678_o2_n_spl_01,
    g274_n_spl_1
  );


  and

  (
    g284_p,
    n406_lo_n,
    g283_p
  );


  and

  (
    g285_p,
    n406_lo_p,
    g283_n
  );


  or

  (
    g286_n,
    g284_p,
    g285_p
  );


  and

  (
    g287_p,
    n658_o2_p_spl_1,
    g274_p_spl_1
  );


  or

  (
    g287_n,
    n658_o2_n_spl_1,
    g274_n_spl_1
  );


  and

  (
    g288_p,
    n418_lo_n,
    g287_p
  );


  and

  (
    g289_p,
    n418_lo_p,
    g287_n
  );


  or

  (
    g290_n,
    g288_p,
    g289_p
  );


  and

  (
    g291_p,
    n862_o2_p,
    n863_o2_p
  );


  or

  (
    g291_n,
    n862_o2_n,
    n863_o2_n
  );


  and

  (
    g292_p,
    g236_n_spl_1,
    g291_p
  );


  or

  (
    g292_n,
    g236_p_spl_1,
    g291_n
  );


  and

  (
    g293_p,
    n602_o2_p_spl_1,
    g292_p_spl_0
  );


  or

  (
    g293_n,
    n602_o2_n_spl_1,
    g292_n_spl_0
  );


  and

  (
    g294_p,
    n430_lo_n,
    g293_p
  );


  and

  (
    g295_p,
    n430_lo_p,
    g293_n
  );


  or

  (
    g296_n,
    g294_p,
    g295_p
  );


  and

  (
    g297_p,
    n639_o2_p_spl_1,
    g292_p_spl_0
  );


  or

  (
    g297_n,
    n639_o2_n_spl_1,
    g292_n_spl_0
  );


  and

  (
    g298_p,
    n442_lo_n,
    g297_p
  );


  and

  (
    g299_p,
    n442_lo_p,
    g297_n
  );


  or

  (
    g300_n,
    g298_p,
    g299_p
  );


  and

  (
    g301_p,
    n678_o2_p_spl_01,
    g292_p_spl_1
  );


  or

  (
    g301_n,
    n678_o2_n_spl_01,
    g292_n_spl_1
  );


  and

  (
    g302_p,
    n454_lo_n,
    g301_p
  );


  and

  (
    g303_p,
    n454_lo_p,
    g301_n
  );


  or

  (
    g304_n,
    g302_p,
    g303_p
  );


  and

  (
    g305_p,
    n658_o2_p_spl_1,
    g292_p_spl_1
  );


  or

  (
    g305_n,
    n658_o2_n_spl_1,
    g292_n_spl_1
  );


  and

  (
    g306_p,
    n466_lo_n,
    g305_p
  );


  and

  (
    g307_p,
    n466_lo_p,
    g305_n
  );


  or

  (
    g308_n,
    g306_p,
    g307_p
  );


  and

  (
    g309_p,
    n686_o2_p,
    n886_o2_p_spl_0
  );


  or

  (
    g309_n,
    n686_o2_n,
    n886_o2_n_spl_0
  );


  and

  (
    g310_p,
    n678_o2_p_spl_1,
    g309_p
  );


  or

  (
    g310_n,
    n678_o2_n_spl_1,
    g309_n
  );


  and

  (
    g311_p,
    n783_o2_p_spl_0,
    g310_p_spl_0
  );


  or

  (
    g311_n,
    n783_o2_n_spl_0,
    g310_n_spl_0
  );


  and

  (
    g312_p,
    n478_lo_n,
    g311_p
  );


  and

  (
    g313_p,
    n478_lo_p,
    g311_n
  );


  or

  (
    g314_n,
    g312_p,
    g313_p
  );


  and

  (
    g315_p,
    n802_o2_p_spl_0,
    g310_p_spl_0
  );


  or

  (
    g315_n,
    n802_o2_n_spl_0,
    g310_n_spl_0
  );


  and

  (
    g316_p,
    n490_lo_n,
    g315_p
  );


  and

  (
    g317_p,
    n490_lo_p,
    g315_n
  );


  or

  (
    g318_n,
    g316_p,
    g317_p
  );


  and

  (
    g319_p,
    n726_o2_p_spl_0,
    g310_p_spl_1
  );


  or

  (
    g319_n,
    n726_o2_n_spl_0,
    g310_n_spl_1
  );


  and

  (
    g320_p,
    n502_lo_n,
    g319_p
  );


  and

  (
    g321_p,
    n502_lo_p,
    g319_n
  );


  or

  (
    g322_n,
    g320_p,
    g321_p
  );


  and

  (
    g323_p,
    n763_o2_p_spl_0,
    g310_p_spl_1
  );


  or

  (
    g323_n,
    n763_o2_n_spl_0,
    g310_n_spl_1
  );


  and

  (
    g324_p,
    n514_lo_n,
    g323_p
  );


  and

  (
    g325_p,
    n514_lo_p,
    g323_n
  );


  or

  (
    g326_n,
    g324_p,
    g325_p
  );


  and

  (
    g327_p,
    n685_o2_p,
    n680_o2_p
  );


  or

  (
    g327_n,
    n685_o2_n,
    n680_o2_n
  );


  and

  (
    g328_p,
    n886_o2_p_spl_0,
    g327_p
  );


  or

  (
    g328_n,
    n886_o2_n_spl_0,
    g327_n
  );


  and

  (
    g329_p,
    n783_o2_p_spl_0,
    g328_p_spl_0
  );


  or

  (
    g329_n,
    n783_o2_n_spl_0,
    g328_n_spl_0
  );


  and

  (
    g330_p,
    n526_lo_n,
    g329_p
  );


  and

  (
    g331_p,
    n526_lo_p,
    g329_n
  );


  or

  (
    g332_n,
    g330_p,
    g331_p
  );


  and

  (
    g333_p,
    n802_o2_p_spl_0,
    g328_p_spl_0
  );


  or

  (
    g333_n,
    n802_o2_n_spl_0,
    g328_n_spl_0
  );


  and

  (
    g334_p,
    n538_lo_n,
    g333_p
  );


  and

  (
    g335_p,
    n538_lo_p,
    g333_n
  );


  or

  (
    g336_n,
    g334_p,
    g335_p
  );


  and

  (
    g337_p,
    n726_o2_p_spl_0,
    g328_p_spl_1
  );


  or

  (
    g337_n,
    n726_o2_n_spl_0,
    g328_n_spl_1
  );


  and

  (
    g338_p,
    n550_lo_n,
    g337_p
  );


  and

  (
    g339_p,
    n550_lo_p,
    g337_n
  );


  or

  (
    g340_n,
    g338_p,
    g339_p
  );


  and

  (
    g341_p,
    n763_o2_p_spl_0,
    g328_p_spl_1
  );


  or

  (
    g341_n,
    n763_o2_n_spl_0,
    g328_n_spl_1
  );


  and

  (
    g342_p,
    n562_lo_n,
    g341_p
  );


  and

  (
    g343_p,
    n562_lo_p,
    g341_n
  );


  or

  (
    g344_n,
    g342_p,
    g343_p
  );


  and

  (
    g345_p,
    n678_o2_p_spl_1,
    n684_o2_p
  );


  or

  (
    g345_n,
    n678_o2_n_spl_1,
    n684_o2_n
  );


  and

  (
    g346_p,
    n886_o2_p_spl_1,
    g345_p
  );


  or

  (
    g346_n,
    n886_o2_n_spl_1,
    g345_n
  );


  and

  (
    g347_p,
    n783_o2_p_spl_1,
    g346_p_spl_0
  );


  or

  (
    g347_n,
    n783_o2_n_spl_1,
    g346_n_spl_0
  );


  and

  (
    g348_p,
    n574_lo_n,
    g347_p
  );


  and

  (
    g349_p,
    n574_lo_p,
    g347_n
  );


  or

  (
    g350_n,
    g348_p,
    g349_p
  );


  and

  (
    g351_p,
    n802_o2_p_spl_1,
    g346_p_spl_0
  );


  or

  (
    g351_n,
    n802_o2_n_spl_1,
    g346_n_spl_0
  );


  and

  (
    g352_p,
    n586_lo_n,
    g351_p
  );


  and

  (
    g353_p,
    n586_lo_p,
    g351_n
  );


  or

  (
    g354_n,
    g352_p,
    g353_p
  );


  and

  (
    g355_p,
    n726_o2_p_spl_1,
    g346_p_spl_1
  );


  or

  (
    g355_n,
    n726_o2_n_spl_1,
    g346_n_spl_1
  );


  and

  (
    g356_p,
    n598_lo_n,
    g355_p
  );


  and

  (
    g357_p,
    n598_lo_p,
    g355_n
  );


  or

  (
    g358_n,
    g356_p,
    g357_p
  );


  and

  (
    g359_p,
    n763_o2_p_spl_1,
    g346_p_spl_1
  );


  or

  (
    g359_n,
    n763_o2_n_spl_1,
    g346_n_spl_1
  );


  and

  (
    g360_p,
    n610_lo_n,
    g359_p
  );


  and

  (
    g361_p,
    n610_lo_p,
    g359_n
  );


  or

  (
    g362_n,
    g360_p,
    g361_p
  );


  and

  (
    g363_p,
    n639_o2_p_spl_1,
    n681_o2_p
  );


  or

  (
    g363_n,
    n639_o2_n_spl_1,
    n681_o2_n
  );


  and

  (
    g364_p,
    n886_o2_p_spl_1,
    g363_p
  );


  or

  (
    g364_n,
    n886_o2_n_spl_1,
    g363_n
  );


  and

  (
    g365_p,
    n783_o2_p_spl_1,
    g364_p_spl_0
  );


  or

  (
    g365_n,
    n783_o2_n_spl_1,
    g364_n_spl_0
  );


  and

  (
    g366_p,
    n622_lo_n,
    g365_p
  );


  and

  (
    g367_p,
    n622_lo_p,
    g365_n
  );


  or

  (
    g368_n,
    g366_p,
    g367_p
  );


  and

  (
    g369_p,
    n802_o2_p_spl_1,
    g364_p_spl_0
  );


  or

  (
    g369_n,
    n802_o2_n_spl_1,
    g364_n_spl_0
  );


  and

  (
    g370_p,
    n634_lo_n,
    g369_p
  );


  and

  (
    g371_p,
    n634_lo_p,
    g369_n
  );


  or

  (
    g372_n,
    g370_p,
    g371_p
  );


  and

  (
    g373_p,
    n726_o2_p_spl_1,
    g364_p_spl_1
  );


  or

  (
    g373_n,
    n726_o2_n_spl_1,
    g364_n_spl_1
  );


  and

  (
    g374_p,
    n646_lo_n,
    g373_p
  );


  and

  (
    g375_p,
    n646_lo_p,
    g373_n
  );


  or

  (
    g376_n,
    g374_p,
    g375_p
  );


  and

  (
    g377_p,
    n763_o2_p_spl_1,
    g364_p_spl_1
  );


  or

  (
    g377_n,
    n763_o2_n_spl_1,
    g364_n_spl_1
  );


  and

  (
    g378_p,
    n658_lo_n,
    g377_p
  );


  and

  (
    g379_p,
    n658_lo_p,
    g377_n
  );


  or

  (
    g380_n,
    g378_p,
    g379_p
  );


  and

  (
    g381_p,
    n600_o2_n,
    n601_o2_n
  );


  or

  (
    g381_n,
    n600_o2_p,
    n601_o2_p
  );


  and

  (
    g382_p,
    n637_o2_n,
    n638_o2_n
  );


  or

  (
    g382_n,
    n637_o2_p,
    n638_o2_p
  );


  and

  (
    g383_p,
    n676_o2_n,
    n677_o2_n
  );


  or

  (
    g383_n,
    n676_o2_p,
    n677_o2_p
  );


  and

  (
    g384_p,
    n656_o2_n,
    n657_o2_n
  );


  or

  (
    g384_n,
    n656_o2_p,
    n657_o2_p
  );


  and

  (
    g385_p,
    n781_o2_n,
    n782_o2_n
  );


  or

  (
    g385_n,
    n781_o2_p,
    n782_o2_p
  );


  and

  (
    g386_p,
    n800_o2_n,
    n801_o2_n
  );


  or

  (
    g386_n,
    n800_o2_p,
    n801_o2_p
  );


  and

  (
    g387_p,
    n724_o2_n,
    n725_o2_n
  );


  or

  (
    g387_n,
    n724_o2_p,
    n725_o2_p
  );


  and

  (
    g388_p,
    n761_o2_n,
    n762_o2_n
  );


  or

  (
    g388_n,
    n761_o2_p,
    n762_o2_p
  );


  or

  (
    g389_n,
    g381_p,
    g382_n_spl_0
  );


  or

  (
    g390_n,
    g383_n_spl_0,
    g384_p
  );


  or

  (
    g391_n,
    g385_p_spl_0,
    g388_p_spl_0
  );


  and

  (
    g392_p,
    g385_p_spl_0,
    g388_p_spl_0
  );


  or

  (
    g392_n,
    g385_n_spl_0,
    g388_n_spl_0
  );


  or

  (
    g393_n,
    g386_p_spl_0,
    g387_p_spl_0
  );


  or

  (
    g394_n,
    g381_n_spl_0,
    g390_n_spl_
  );


  or

  (
    g395_n,
    g381_n_spl_0,
    g384_n_spl_0
  );


  or

  (
    g396_n,
    g382_p,
    g395_n_spl_
  );


  or

  (
    g397_n,
    g384_n_spl_0,
    g389_n_spl_
  );


  and

  (
    g398_p,
    g386_p_spl_0,
    g387_p_spl_0
  );


  or

  (
    g398_n,
    g386_n_spl_0,
    g387_n_spl_0
  );


  or

  (
    g399_n,
    g383_p,
    g395_n_spl_
  );


  and

  (
    g400_p,
    g394_n_spl_,
    g399_n
  );


  or

  (
    g401_n,
    g382_n_spl_0,
    g400_p
  );


  and

  (
    g402_p,
    g396_n_spl_,
    g397_n_spl_
  );


  or

  (
    g403_n,
    g383_n_spl_0,
    g402_p
  );


  and

  (
    g404_p,
    g385_n_spl_0,
    g386_p_spl_
  );


  and

  (
    g405_p,
    g385_p_spl_,
    g386_n_spl_0
  );


  and

  (
    g406_p,
    g387_n_spl_0,
    g388_p_spl_
  );


  and

  (
    g407_p,
    g387_p_spl_,
    g388_n_spl_0
  );


  and

  (
    g408_p,
    g391_n_spl_,
    g392_n_spl_
  );


  or

  (
    g409_n,
    g398_n_spl_,
    g408_p
  );


  and

  (
    g410_p,
    g392_p,
    g393_n_spl_
  );


  or

  (
    g411_n,
    g398_p,
    g410_p
  );


  and

  (
    g412_p,
    g409_n,
    g411_n
  );


  and

  (
    g413_p,
    lo002_buf_o2_p_spl_0,
    lo018_buf_o2_n_spl_
  );


  or

  (
    g413_n,
    lo002_buf_o2_n_spl_,
    lo018_buf_o2_p_spl_0
  );


  and

  (
    g414_p,
    lo002_buf_o2_n_spl_,
    lo018_buf_o2_p_spl_0
  );


  or

  (
    g414_n,
    lo002_buf_o2_p_spl_0,
    lo018_buf_o2_n_spl_
  );


  and

  (
    g415_p,
    g413_n,
    g414_n
  );


  or

  (
    g415_n,
    g413_p,
    g414_p
  );


  and

  (
    g416_p,
    lo034_buf_o2_p_spl_0,
    lo050_buf_o2_n_spl_
  );


  or

  (
    g416_n,
    lo034_buf_o2_n_spl_,
    lo050_buf_o2_p_spl_0
  );


  and

  (
    g417_p,
    lo034_buf_o2_n_spl_,
    lo050_buf_o2_p_spl_0
  );


  or

  (
    g417_n,
    lo034_buf_o2_p_spl_0,
    lo050_buf_o2_n_spl_
  );


  and

  (
    g418_p,
    g416_n,
    g417_n
  );


  or

  (
    g418_n,
    g416_p,
    g417_p
  );


  and

  (
    g419_p,
    g415_p,
    g418_n
  );


  and

  (
    g420_p,
    g415_n,
    g418_p
  );


  or

  (
    g421_n,
    g419_p,
    g420_p
  );


  and

  (
    g422_p,
    lo129_buf_o2_p,
    lo161_buf_o2_p_spl_00
  );


  or

  (
    g422_n,
    lo129_buf_o2_n,
    lo161_buf_o2_n_spl_00
  );


  and

  (
    g423_p,
    n584_o2_n_spl_0,
    n593_o2_p_spl_0
  );


  or

  (
    g423_n,
    n584_o2_p_spl_0,
    n593_o2_n_spl_0
  );


  and

  (
    g424_p,
    n584_o2_p_spl_0,
    n593_o2_n_spl_0
  );


  or

  (
    g424_n,
    n584_o2_n_spl_0,
    n593_o2_p_spl_0
  );


  and

  (
    g425_p,
    g423_n,
    g424_n
  );


  or

  (
    g425_n,
    g423_p,
    g424_p
  );


  or

  (
    g426_n,
    g422_p,
    g425_p
  );


  or

  (
    g427_n,
    g422_n,
    g425_n
  );


  and

  (
    g428_p,
    g426_n,
    g427_n
  );


  or

  (
    g429_n,
    g421_n_spl_,
    g428_p_spl_
  );


  and

  (
    g430_p,
    g421_n_spl_,
    g428_p_spl_
  );


  and

  (
    g431_p,
    lo006_buf_o2_p_spl_0,
    lo022_buf_o2_n_spl_
  );


  or

  (
    g431_n,
    lo006_buf_o2_n_spl_,
    lo022_buf_o2_p_spl_0
  );


  and

  (
    g432_p,
    lo006_buf_o2_n_spl_,
    lo022_buf_o2_p_spl_0
  );


  or

  (
    g432_n,
    lo006_buf_o2_p_spl_0,
    lo022_buf_o2_n_spl_
  );


  and

  (
    g433_p,
    g431_n,
    g432_n
  );


  or

  (
    g433_n,
    g431_p,
    g432_p
  );


  and

  (
    g434_p,
    lo038_buf_o2_p_spl_0,
    lo054_buf_o2_n_spl_
  );


  or

  (
    g434_n,
    lo038_buf_o2_n_spl_,
    lo054_buf_o2_p_spl_0
  );


  and

  (
    g435_p,
    lo038_buf_o2_n_spl_,
    lo054_buf_o2_p_spl_0
  );


  or

  (
    g435_n,
    lo038_buf_o2_p_spl_0,
    lo054_buf_o2_n_spl_
  );


  and

  (
    g436_p,
    g434_n,
    g435_n
  );


  or

  (
    g436_n,
    g434_p,
    g435_p
  );


  and

  (
    g437_p,
    g433_p,
    g436_n
  );


  and

  (
    g438_p,
    g433_n,
    g436_p
  );


  or

  (
    g439_n,
    g437_p,
    g438_p
  );


  and

  (
    g440_p,
    lo133_buf_o2_p,
    lo161_buf_o2_p_spl_00
  );


  or

  (
    g440_n,
    lo133_buf_o2_n,
    lo161_buf_o2_n_spl_00
  );


  and

  (
    g441_p,
    n630_o2_p_spl_0,
    n621_o2_n_spl_0
  );


  or

  (
    g441_n,
    n630_o2_n_spl_0,
    n621_o2_p_spl_0
  );


  and

  (
    g442_p,
    n630_o2_n_spl_0,
    n621_o2_p_spl_0
  );


  or

  (
    g442_n,
    n630_o2_p_spl_0,
    n621_o2_n_spl_0
  );


  and

  (
    g443_p,
    g441_n,
    g442_n
  );


  or

  (
    g443_n,
    g441_p,
    g442_p
  );


  or

  (
    g444_n,
    g440_p,
    g443_p
  );


  or

  (
    g445_n,
    g440_n,
    g443_n
  );


  and

  (
    g446_p,
    g444_n,
    g445_n
  );


  or

  (
    g447_n,
    g439_n_spl_,
    g446_p_spl_
  );


  and

  (
    g448_p,
    g439_n_spl_,
    g446_p_spl_
  );


  and

  (
    g449_p,
    lo010_buf_o2_p_spl_0,
    lo026_buf_o2_n_spl_
  );


  or

  (
    g449_n,
    lo010_buf_o2_n_spl_,
    lo026_buf_o2_p_spl_0
  );


  and

  (
    g450_p,
    lo010_buf_o2_n_spl_,
    lo026_buf_o2_p_spl_0
  );


  or

  (
    g450_n,
    lo010_buf_o2_p_spl_0,
    lo026_buf_o2_n_spl_
  );


  and

  (
    g451_p,
    g449_n,
    g450_n
  );


  or

  (
    g451_n,
    g449_p,
    g450_p
  );


  and

  (
    g452_p,
    lo042_buf_o2_p_spl_0,
    lo058_buf_o2_n_spl_
  );


  or

  (
    g452_n,
    lo042_buf_o2_n_spl_,
    lo058_buf_o2_p_spl_0
  );


  and

  (
    g453_p,
    lo042_buf_o2_n_spl_,
    lo058_buf_o2_p_spl_0
  );


  or

  (
    g453_n,
    lo042_buf_o2_p_spl_0,
    lo058_buf_o2_n_spl_
  );


  and

  (
    g454_p,
    g452_n,
    g453_n
  );


  or

  (
    g454_n,
    g452_p,
    g453_p
  );


  and

  (
    g455_p,
    g451_p,
    g454_n
  );


  and

  (
    g456_p,
    g451_n,
    g454_p
  );


  or

  (
    g457_n,
    g455_p,
    g456_p
  );


  and

  (
    g458_p,
    lo137_buf_o2_p,
    lo161_buf_o2_p_spl_01
  );


  or

  (
    g458_n,
    lo137_buf_o2_n,
    lo161_buf_o2_n_spl_01
  );


  and

  (
    g459_p,
    n584_o2_n_spl_1,
    n630_o2_p_spl_1
  );


  or

  (
    g459_n,
    n584_o2_p_spl_1,
    n630_o2_n_spl_1
  );


  and

  (
    g460_p,
    n584_o2_p_spl_1,
    n630_o2_n_spl_1
  );


  or

  (
    g460_n,
    n584_o2_n_spl_1,
    n630_o2_p_spl_1
  );


  and

  (
    g461_p,
    g459_n,
    g460_n
  );


  or

  (
    g461_n,
    g459_p,
    g460_p
  );


  or

  (
    g462_n,
    g458_p,
    g461_p
  );


  or

  (
    g463_n,
    g458_n,
    g461_n
  );


  and

  (
    g464_p,
    g462_n,
    g463_n
  );


  or

  (
    g465_n,
    g457_n_spl_,
    g464_p_spl_
  );


  and

  (
    g466_p,
    g457_n_spl_,
    g464_p_spl_
  );


  and

  (
    g467_p,
    lo014_buf_o2_p_spl_0,
    lo030_buf_o2_n_spl_
  );


  or

  (
    g467_n,
    lo014_buf_o2_n_spl_,
    lo030_buf_o2_p_spl_0
  );


  and

  (
    g468_p,
    lo014_buf_o2_n_spl_,
    lo030_buf_o2_p_spl_0
  );


  or

  (
    g468_n,
    lo014_buf_o2_p_spl_0,
    lo030_buf_o2_n_spl_
  );


  and

  (
    g469_p,
    g467_n,
    g468_n
  );


  or

  (
    g469_n,
    g467_p,
    g468_p
  );


  and

  (
    g470_p,
    lo046_buf_o2_p_spl_0,
    lo062_buf_o2_n_spl_
  );


  or

  (
    g470_n,
    lo046_buf_o2_n_spl_,
    lo062_buf_o2_p_spl_0
  );


  and

  (
    g471_p,
    lo046_buf_o2_n_spl_,
    lo062_buf_o2_p_spl_0
  );


  or

  (
    g471_n,
    lo046_buf_o2_p_spl_0,
    lo062_buf_o2_n_spl_
  );


  and

  (
    g472_p,
    g470_n,
    g471_n
  );


  or

  (
    g472_n,
    g470_p,
    g471_p
  );


  and

  (
    g473_p,
    g469_p,
    g472_n
  );


  and

  (
    g474_p,
    g469_n,
    g472_p
  );


  or

  (
    g475_n,
    g473_p,
    g474_p
  );


  and

  (
    g476_p,
    lo141_buf_o2_p,
    lo161_buf_o2_p_spl_01
  );


  or

  (
    g476_n,
    lo141_buf_o2_n,
    lo161_buf_o2_n_spl_01
  );


  and

  (
    g477_p,
    n593_o2_n_spl_1,
    n621_o2_p_spl_1
  );


  or

  (
    g477_n,
    n593_o2_p_spl_1,
    n621_o2_n_spl_1
  );


  and

  (
    g478_p,
    n593_o2_p_spl_1,
    n621_o2_n_spl_1
  );


  or

  (
    g478_n,
    n593_o2_n_spl_1,
    n621_o2_p_spl_1
  );


  and

  (
    g479_p,
    g477_n,
    g478_n
  );


  or

  (
    g479_n,
    g477_p,
    g478_p
  );


  or

  (
    g480_n,
    g476_p,
    g479_p
  );


  or

  (
    g481_n,
    g476_n,
    g479_n
  );


  and

  (
    g482_p,
    g480_n,
    g481_n
  );


  or

  (
    g483_n,
    g475_n_spl_,
    g482_p_spl_
  );


  and

  (
    g484_p,
    g475_n_spl_,
    g482_p_spl_
  );


  and

  (
    g485_p,
    lo066_buf_o2_p_spl_0,
    lo082_buf_o2_n_spl_
  );


  or

  (
    g485_n,
    lo066_buf_o2_n_spl_,
    lo082_buf_o2_p_spl_0
  );


  and

  (
    g486_p,
    lo066_buf_o2_n_spl_,
    lo082_buf_o2_p_spl_0
  );


  or

  (
    g486_n,
    lo066_buf_o2_p_spl_0,
    lo082_buf_o2_n_spl_
  );


  and

  (
    g487_p,
    g485_n,
    g486_n
  );


  or

  (
    g487_n,
    g485_p,
    g486_p
  );


  and

  (
    g488_p,
    lo098_buf_o2_p_spl_0,
    lo114_buf_o2_n_spl_
  );


  or

  (
    g488_n,
    lo098_buf_o2_n_spl_,
    lo114_buf_o2_p_spl_0
  );


  and

  (
    g489_p,
    lo098_buf_o2_n_spl_,
    lo114_buf_o2_p_spl_0
  );


  or

  (
    g489_n,
    lo098_buf_o2_p_spl_0,
    lo114_buf_o2_n_spl_
  );


  and

  (
    g490_p,
    g488_n,
    g489_n
  );


  or

  (
    g490_n,
    g488_p,
    g489_p
  );


  and

  (
    g491_p,
    g487_p,
    g490_n
  );


  and

  (
    g492_p,
    g487_n,
    g490_p
  );


  or

  (
    g493_n,
    g491_p,
    g492_p
  );


  and

  (
    g494_p,
    lo145_buf_o2_p,
    lo161_buf_o2_p_spl_10
  );


  or

  (
    g494_n,
    lo145_buf_o2_n,
    lo161_buf_o2_n_spl_10
  );


  and

  (
    g495_p,
    n708_o2_n_spl_0,
    n745_o2_p_spl_0
  );


  or

  (
    g495_n,
    n708_o2_p_spl_0,
    n745_o2_n_spl_0
  );


  and

  (
    g496_p,
    n708_o2_p_spl_0,
    n745_o2_n_spl_0
  );


  or

  (
    g496_n,
    n708_o2_n_spl_0,
    n745_o2_p_spl_0
  );


  and

  (
    g497_p,
    g495_n,
    g496_n
  );


  or

  (
    g497_n,
    g495_p,
    g496_p
  );


  or

  (
    g498_n,
    g494_p,
    g497_p
  );


  or

  (
    g499_n,
    g494_n,
    g497_n
  );


  and

  (
    g500_p,
    g498_n,
    g499_n
  );


  or

  (
    g501_n,
    g493_n_spl_,
    g500_p_spl_
  );


  and

  (
    g502_p,
    g493_n_spl_,
    g500_p_spl_
  );


  and

  (
    g503_p,
    lo070_buf_o2_p_spl_0,
    lo086_buf_o2_n_spl_
  );


  or

  (
    g503_n,
    lo070_buf_o2_n_spl_,
    lo086_buf_o2_p_spl_0
  );


  and

  (
    g504_p,
    lo070_buf_o2_n_spl_,
    lo086_buf_o2_p_spl_0
  );


  or

  (
    g504_n,
    lo070_buf_o2_p_spl_0,
    lo086_buf_o2_n_spl_
  );


  and

  (
    g505_p,
    g503_n,
    g504_n
  );


  or

  (
    g505_n,
    g503_p,
    g504_p
  );


  and

  (
    g506_p,
    lo102_buf_o2_p_spl_0,
    lo118_buf_o2_n_spl_
  );


  or

  (
    g506_n,
    lo102_buf_o2_n_spl_,
    lo118_buf_o2_p_spl_0
  );


  and

  (
    g507_p,
    lo102_buf_o2_n_spl_,
    lo118_buf_o2_p_spl_0
  );


  or

  (
    g507_n,
    lo102_buf_o2_p_spl_0,
    lo118_buf_o2_n_spl_
  );


  and

  (
    g508_p,
    g506_n,
    g507_n
  );


  or

  (
    g508_n,
    g506_p,
    g507_p
  );


  and

  (
    g509_p,
    g505_p,
    g508_n
  );


  and

  (
    g510_p,
    g505_n,
    g508_p
  );


  or

  (
    g511_n,
    g509_p,
    g510_p
  );


  and

  (
    g512_p,
    lo149_buf_o2_p,
    lo161_buf_o2_p_spl_10
  );


  or

  (
    g512_n,
    lo149_buf_o2_n,
    lo161_buf_o2_n_spl_10
  );


  and

  (
    g513_p,
    n717_o2_n_spl_0,
    n754_o2_p_spl_0
  );


  or

  (
    g513_n,
    n717_o2_p_spl_0,
    n754_o2_n_spl_0
  );


  and

  (
    g514_p,
    n717_o2_p_spl_0,
    n754_o2_n_spl_0
  );


  or

  (
    g514_n,
    n717_o2_n_spl_0,
    n754_o2_p_spl_0
  );


  and

  (
    g515_p,
    g513_n,
    g514_n
  );


  or

  (
    g515_n,
    g513_p,
    g514_p
  );


  or

  (
    g516_n,
    g512_p,
    g515_p
  );


  or

  (
    g517_n,
    g512_n,
    g515_n
  );


  and

  (
    g518_p,
    g516_n,
    g517_n
  );


  or

  (
    g519_n,
    g511_n_spl_,
    g518_p_spl_
  );


  and

  (
    g520_p,
    g511_n_spl_,
    g518_p_spl_
  );


  and

  (
    g521_p,
    lo074_buf_o2_p_spl_0,
    lo090_buf_o2_n_spl_
  );


  or

  (
    g521_n,
    lo074_buf_o2_n_spl_,
    lo090_buf_o2_p_spl_0
  );


  and

  (
    g522_p,
    lo074_buf_o2_n_spl_,
    lo090_buf_o2_p_spl_0
  );


  or

  (
    g522_n,
    lo074_buf_o2_p_spl_0,
    lo090_buf_o2_n_spl_
  );


  and

  (
    g523_p,
    g521_n,
    g522_n
  );


  or

  (
    g523_n,
    g521_p,
    g522_p
  );


  and

  (
    g524_p,
    lo106_buf_o2_p_spl_0,
    lo122_buf_o2_n_spl_
  );


  or

  (
    g524_n,
    lo106_buf_o2_n_spl_,
    lo122_buf_o2_p_spl_0
  );


  and

  (
    g525_p,
    lo106_buf_o2_n_spl_,
    lo122_buf_o2_p_spl_0
  );


  or

  (
    g525_n,
    lo106_buf_o2_p_spl_0,
    lo122_buf_o2_n_spl_
  );


  and

  (
    g526_p,
    g524_n,
    g525_n
  );


  or

  (
    g526_n,
    g524_p,
    g525_p
  );


  and

  (
    g527_p,
    g523_p,
    g526_n
  );


  and

  (
    g528_p,
    g523_n,
    g526_p
  );


  or

  (
    g529_n,
    g527_p,
    g528_p
  );


  and

  (
    g530_p,
    lo153_buf_o2_p,
    lo161_buf_o2_p_spl_11
  );


  or

  (
    g530_n,
    lo153_buf_o2_n,
    lo161_buf_o2_n_spl_11
  );


  and

  (
    g531_p,
    n708_o2_n_spl_1,
    n717_o2_p_spl_1
  );


  or

  (
    g531_n,
    n708_o2_p_spl_1,
    n717_o2_n_spl_1
  );


  and

  (
    g532_p,
    n708_o2_p_spl_1,
    n717_o2_n_spl_1
  );


  or

  (
    g532_n,
    n708_o2_n_spl_1,
    n717_o2_p_spl_1
  );


  and

  (
    g533_p,
    g531_n,
    g532_n
  );


  or

  (
    g533_n,
    g531_p,
    g532_p
  );


  or

  (
    g534_n,
    g530_p,
    g533_p
  );


  or

  (
    g535_n,
    g530_n,
    g533_n
  );


  and

  (
    g536_p,
    g534_n,
    g535_n
  );


  or

  (
    g537_n,
    g529_n_spl_,
    g536_p_spl_
  );


  and

  (
    g538_p,
    g529_n_spl_,
    g536_p_spl_
  );


  and

  (
    g539_p,
    lo078_buf_o2_p_spl_0,
    lo094_buf_o2_n_spl_
  );


  or

  (
    g539_n,
    lo078_buf_o2_n_spl_,
    lo094_buf_o2_p_spl_0
  );


  and

  (
    g540_p,
    lo078_buf_o2_n_spl_,
    lo094_buf_o2_p_spl_0
  );


  or

  (
    g540_n,
    lo078_buf_o2_p_spl_0,
    lo094_buf_o2_n_spl_
  );


  and

  (
    g541_p,
    g539_n,
    g540_n
  );


  or

  (
    g541_n,
    g539_p,
    g540_p
  );


  and

  (
    g542_p,
    lo110_buf_o2_p_spl_0,
    lo126_buf_o2_n_spl_
  );


  or

  (
    g542_n,
    lo110_buf_o2_n_spl_,
    lo126_buf_o2_p_spl_0
  );


  and

  (
    g543_p,
    lo110_buf_o2_n_spl_,
    lo126_buf_o2_p_spl_0
  );


  or

  (
    g543_n,
    lo110_buf_o2_p_spl_0,
    lo126_buf_o2_n_spl_
  );


  and

  (
    g544_p,
    g542_n,
    g543_n
  );


  or

  (
    g544_n,
    g542_p,
    g543_p
  );


  and

  (
    g545_p,
    g541_p,
    g544_n
  );


  and

  (
    g546_p,
    g541_n,
    g544_p
  );


  or

  (
    g547_n,
    g545_p,
    g546_p
  );


  and

  (
    g548_p,
    lo157_buf_o2_p,
    lo161_buf_o2_p_spl_11
  );


  or

  (
    g548_n,
    lo157_buf_o2_n,
    lo161_buf_o2_n_spl_11
  );


  and

  (
    g549_p,
    n745_o2_n_spl_1,
    n754_o2_p_spl_1
  );


  or

  (
    g549_n,
    n745_o2_p_spl_1,
    n754_o2_n_spl_1
  );


  and

  (
    g550_p,
    n745_o2_p_spl_1,
    n754_o2_n_spl_1
  );


  or

  (
    g550_n,
    n745_o2_n_spl_1,
    n754_o2_p_spl_1
  );


  and

  (
    g551_p,
    g549_n,
    g550_n
  );


  or

  (
    g551_n,
    g549_p,
    g550_p
  );


  or

  (
    g552_n,
    g548_p,
    g551_p
  );


  or

  (
    g553_n,
    g548_n,
    g551_n
  );


  and

  (
    g554_p,
    g552_n,
    g553_n
  );


  or

  (
    g555_n,
    g547_n_spl_,
    g554_p_spl_
  );


  and

  (
    g556_p,
    g547_n_spl_,
    g554_p_spl_
  );


  and

  (
    g557_p,
    lo001_buf_o2_p_spl_0,
    lo005_buf_o2_n_spl_
  );


  or

  (
    g557_n,
    lo001_buf_o2_n_spl_,
    lo005_buf_o2_p_spl_0
  );


  and

  (
    g558_p,
    lo001_buf_o2_n_spl_,
    lo005_buf_o2_p_spl_0
  );


  or

  (
    g558_n,
    lo001_buf_o2_p_spl_0,
    lo005_buf_o2_n_spl_
  );


  and

  (
    g559_p,
    g557_n,
    g558_n
  );


  or

  (
    g559_n,
    g557_p,
    g558_p
  );


  and

  (
    g560_p,
    lo009_buf_o2_p_spl_0,
    lo013_buf_o2_n_spl_
  );


  or

  (
    g560_n,
    lo009_buf_o2_n_spl_,
    lo013_buf_o2_p_spl_0
  );


  and

  (
    g561_p,
    lo009_buf_o2_n_spl_,
    lo013_buf_o2_p_spl_0
  );


  or

  (
    g561_n,
    lo009_buf_o2_p_spl_0,
    lo013_buf_o2_n_spl_
  );


  and

  (
    g562_p,
    g560_n,
    g561_n
  );


  or

  (
    g562_n,
    g560_p,
    g561_p
  );


  and

  (
    g563_p,
    g559_p,
    g562_n
  );


  and

  (
    g564_p,
    g559_n,
    g562_p
  );


  or

  (
    g565_n,
    g563_p,
    g564_p
  );


  and

  (
    g566_p,
    lo017_buf_o2_p_spl_0,
    lo021_buf_o2_n_spl_
  );


  or

  (
    g566_n,
    lo017_buf_o2_n_spl_,
    lo021_buf_o2_p_spl_0
  );


  and

  (
    g567_p,
    lo017_buf_o2_n_spl_,
    lo021_buf_o2_p_spl_0
  );


  or

  (
    g567_n,
    lo017_buf_o2_p_spl_0,
    lo021_buf_o2_n_spl_
  );


  and

  (
    g568_p,
    g566_n,
    g567_n
  );


  or

  (
    g568_n,
    g566_p,
    g567_p
  );


  and

  (
    g569_p,
    lo025_buf_o2_p_spl_0,
    lo029_buf_o2_n_spl_
  );


  or

  (
    g569_n,
    lo025_buf_o2_n_spl_,
    lo029_buf_o2_p_spl_0
  );


  and

  (
    g570_p,
    lo025_buf_o2_n_spl_,
    lo029_buf_o2_p_spl_0
  );


  or

  (
    g570_n,
    lo025_buf_o2_p_spl_0,
    lo029_buf_o2_n_spl_
  );


  and

  (
    g571_p,
    g569_n,
    g570_n
  );


  or

  (
    g571_n,
    g569_p,
    g570_p
  );


  and

  (
    g572_p,
    g568_p,
    g571_n
  );


  and

  (
    g573_p,
    g568_n,
    g571_p
  );


  or

  (
    g574_n,
    g572_p,
    g573_p
  );


  and

  (
    g575_p,
    lo033_buf_o2_p_spl_0,
    lo037_buf_o2_n_spl_
  );


  or

  (
    g575_n,
    lo033_buf_o2_n_spl_,
    lo037_buf_o2_p_spl_0
  );


  and

  (
    g576_p,
    lo033_buf_o2_n_spl_,
    lo037_buf_o2_p_spl_0
  );


  or

  (
    g576_n,
    lo033_buf_o2_p_spl_0,
    lo037_buf_o2_n_spl_
  );


  and

  (
    g577_p,
    g575_n,
    g576_n
  );


  or

  (
    g577_n,
    g575_p,
    g576_p
  );


  and

  (
    g578_p,
    lo041_buf_o2_p_spl_0,
    lo045_buf_o2_n_spl_
  );


  or

  (
    g578_n,
    lo041_buf_o2_n_spl_,
    lo045_buf_o2_p_spl_0
  );


  and

  (
    g579_p,
    lo041_buf_o2_n_spl_,
    lo045_buf_o2_p_spl_0
  );


  or

  (
    g579_n,
    lo041_buf_o2_p_spl_0,
    lo045_buf_o2_n_spl_
  );


  and

  (
    g580_p,
    g578_n,
    g579_n
  );


  or

  (
    g580_n,
    g578_p,
    g579_p
  );


  and

  (
    g581_p,
    g577_p,
    g580_n
  );


  and

  (
    g582_p,
    g577_n,
    g580_p
  );


  or

  (
    g583_n,
    g581_p,
    g582_p
  );


  and

  (
    g584_p,
    lo049_buf_o2_p_spl_0,
    lo053_buf_o2_n_spl_
  );


  or

  (
    g584_n,
    lo049_buf_o2_n_spl_,
    lo053_buf_o2_p_spl_0
  );


  and

  (
    g585_p,
    lo049_buf_o2_n_spl_,
    lo053_buf_o2_p_spl_0
  );


  or

  (
    g585_n,
    lo049_buf_o2_p_spl_0,
    lo053_buf_o2_n_spl_
  );


  and

  (
    g586_p,
    g584_n,
    g585_n
  );


  or

  (
    g586_n,
    g584_p,
    g585_p
  );


  and

  (
    g587_p,
    lo057_buf_o2_p_spl_0,
    lo061_buf_o2_n_spl_
  );


  or

  (
    g587_n,
    lo057_buf_o2_n_spl_,
    lo061_buf_o2_p_spl_0
  );


  and

  (
    g588_p,
    lo057_buf_o2_n_spl_,
    lo061_buf_o2_p_spl_0
  );


  or

  (
    g588_n,
    lo057_buf_o2_p_spl_0,
    lo061_buf_o2_n_spl_
  );


  and

  (
    g589_p,
    g587_n,
    g588_n
  );


  or

  (
    g589_n,
    g587_p,
    g588_p
  );


  and

  (
    g590_p,
    g586_p,
    g589_n
  );


  and

  (
    g591_p,
    g586_n,
    g589_p
  );


  or

  (
    g592_n,
    g590_p,
    g591_p
  );


  and

  (
    g593_p,
    lo065_buf_o2_p_spl_0,
    lo069_buf_o2_n_spl_
  );


  or

  (
    g593_n,
    lo065_buf_o2_n_spl_,
    lo069_buf_o2_p_spl_0
  );


  and

  (
    g594_p,
    lo065_buf_o2_n_spl_,
    lo069_buf_o2_p_spl_0
  );


  or

  (
    g594_n,
    lo065_buf_o2_p_spl_0,
    lo069_buf_o2_n_spl_
  );


  and

  (
    g595_p,
    g593_n,
    g594_n
  );


  or

  (
    g595_n,
    g593_p,
    g594_p
  );


  and

  (
    g596_p,
    lo073_buf_o2_p_spl_0,
    lo077_buf_o2_n_spl_
  );


  or

  (
    g596_n,
    lo073_buf_o2_n_spl_,
    lo077_buf_o2_p_spl_0
  );


  and

  (
    g597_p,
    lo073_buf_o2_n_spl_,
    lo077_buf_o2_p_spl_0
  );


  or

  (
    g597_n,
    lo073_buf_o2_p_spl_0,
    lo077_buf_o2_n_spl_
  );


  and

  (
    g598_p,
    g596_n,
    g597_n
  );


  or

  (
    g598_n,
    g596_p,
    g597_p
  );


  and

  (
    g599_p,
    g595_p,
    g598_n
  );


  and

  (
    g600_p,
    g595_n,
    g598_p
  );


  or

  (
    g601_n,
    g599_p,
    g600_p
  );


  and

  (
    g602_p,
    lo081_buf_o2_p_spl_0,
    lo085_buf_o2_n_spl_
  );


  or

  (
    g602_n,
    lo081_buf_o2_n_spl_,
    lo085_buf_o2_p_spl_0
  );


  and

  (
    g603_p,
    lo081_buf_o2_n_spl_,
    lo085_buf_o2_p_spl_0
  );


  or

  (
    g603_n,
    lo081_buf_o2_p_spl_0,
    lo085_buf_o2_n_spl_
  );


  and

  (
    g604_p,
    g602_n,
    g603_n
  );


  or

  (
    g604_n,
    g602_p,
    g603_p
  );


  and

  (
    g605_p,
    lo089_buf_o2_p_spl_0,
    lo093_buf_o2_n_spl_
  );


  or

  (
    g605_n,
    lo089_buf_o2_n_spl_,
    lo093_buf_o2_p_spl_0
  );


  and

  (
    g606_p,
    lo089_buf_o2_n_spl_,
    lo093_buf_o2_p_spl_0
  );


  or

  (
    g606_n,
    lo089_buf_o2_p_spl_0,
    lo093_buf_o2_n_spl_
  );


  and

  (
    g607_p,
    g605_n,
    g606_n
  );


  or

  (
    g607_n,
    g605_p,
    g606_p
  );


  and

  (
    g608_p,
    g604_p,
    g607_n
  );


  and

  (
    g609_p,
    g604_n,
    g607_p
  );


  or

  (
    g610_n,
    g608_p,
    g609_p
  );


  and

  (
    g611_p,
    lo097_buf_o2_p_spl_0,
    lo101_buf_o2_n_spl_
  );


  or

  (
    g611_n,
    lo097_buf_o2_n_spl_,
    lo101_buf_o2_p_spl_0
  );


  and

  (
    g612_p,
    lo097_buf_o2_n_spl_,
    lo101_buf_o2_p_spl_0
  );


  or

  (
    g612_n,
    lo097_buf_o2_p_spl_0,
    lo101_buf_o2_n_spl_
  );


  and

  (
    g613_p,
    g611_n,
    g612_n
  );


  or

  (
    g613_n,
    g611_p,
    g612_p
  );


  and

  (
    g614_p,
    lo105_buf_o2_p_spl_0,
    lo109_buf_o2_n_spl_
  );


  or

  (
    g614_n,
    lo105_buf_o2_n_spl_,
    lo109_buf_o2_p_spl_0
  );


  and

  (
    g615_p,
    lo105_buf_o2_n_spl_,
    lo109_buf_o2_p_spl_0
  );


  or

  (
    g615_n,
    lo105_buf_o2_p_spl_0,
    lo109_buf_o2_n_spl_
  );


  and

  (
    g616_p,
    g614_n,
    g615_n
  );


  or

  (
    g616_n,
    g614_p,
    g615_p
  );


  and

  (
    g617_p,
    g613_p,
    g616_n
  );


  and

  (
    g618_p,
    g613_n,
    g616_p
  );


  or

  (
    g619_n,
    g617_p,
    g618_p
  );


  and

  (
    g620_p,
    lo113_buf_o2_p_spl_0,
    lo117_buf_o2_n_spl_
  );


  or

  (
    g620_n,
    lo113_buf_o2_n_spl_,
    lo117_buf_o2_p_spl_0
  );


  and

  (
    g621_p,
    lo113_buf_o2_n_spl_,
    lo117_buf_o2_p_spl_0
  );


  or

  (
    g621_n,
    lo113_buf_o2_p_spl_0,
    lo117_buf_o2_n_spl_
  );


  and

  (
    g622_p,
    g620_n,
    g621_n
  );


  or

  (
    g622_n,
    g620_p,
    g621_p
  );


  and

  (
    g623_p,
    lo121_buf_o2_p_spl_0,
    lo125_buf_o2_n_spl_
  );


  or

  (
    g623_n,
    lo121_buf_o2_n_spl_,
    lo125_buf_o2_p_spl_0
  );


  and

  (
    g624_p,
    lo121_buf_o2_n_spl_,
    lo125_buf_o2_p_spl_0
  );


  or

  (
    g624_n,
    lo121_buf_o2_p_spl_0,
    lo125_buf_o2_n_spl_
  );


  and

  (
    g625_p,
    g623_n,
    g624_n
  );


  or

  (
    g625_n,
    g623_p,
    g624_p
  );


  and

  (
    g626_p,
    g622_p,
    g625_n
  );


  and

  (
    g627_p,
    g622_n,
    g625_p
  );


  or

  (
    g628_n,
    g626_p,
    g627_p
  );


  buf

  (
    G468,
    g242_n
  );


  buf

  (
    G469,
    g246_n
  );


  buf

  (
    G470,
    g250_n
  );


  buf

  (
    G471,
    g254_n
  );


  buf

  (
    G472,
    g260_n
  );


  buf

  (
    G473,
    g264_n
  );


  buf

  (
    G474,
    g268_n
  );


  buf

  (
    G475,
    g272_n
  );


  buf

  (
    G476,
    g278_n
  );


  buf

  (
    G477,
    g282_n
  );


  buf

  (
    G478,
    g286_n
  );


  buf

  (
    G479,
    g290_n
  );


  buf

  (
    G480,
    g296_n
  );


  buf

  (
    G481,
    g300_n
  );


  buf

  (
    G482,
    g304_n
  );


  buf

  (
    G483,
    g308_n
  );


  buf

  (
    G484,
    g314_n
  );


  buf

  (
    G485,
    g318_n
  );


  buf

  (
    G486,
    g322_n
  );


  buf

  (
    G487,
    g326_n
  );


  buf

  (
    G488,
    g332_n
  );


  buf

  (
    G489,
    g336_n
  );


  buf

  (
    G490,
    g340_n
  );


  buf

  (
    G491,
    g344_n
  );


  buf

  (
    G492,
    g350_n
  );


  buf

  (
    G493,
    g354_n
  );


  buf

  (
    G494,
    g358_n
  );


  buf

  (
    G495,
    g362_n
  );


  buf

  (
    G496,
    g368_n
  );


  buf

  (
    G497,
    g372_n
  );


  buf

  (
    G498,
    g376_n
  );


  buf

  (
    G499,
    g380_n
  );


  buf

  (
    n1020_li003_li003,
    n1589_o2_p
  );


  buf

  (
    n1032_li007_li007,
    n1590_o2_p
  );


  buf

  (
    n1044_li011_li011,
    n1591_o2_p
  );


  buf

  (
    n1056_li015_li015,
    n1592_o2_p
  );


  buf

  (
    n1068_li019_li019,
    n1593_o2_p
  );


  buf

  (
    n1080_li023_li023,
    n1594_o2_p
  );


  buf

  (
    n1092_li027_li027,
    n1595_o2_p
  );


  buf

  (
    n1104_li031_li031,
    n1596_o2_p
  );


  buf

  (
    n1116_li035_li035,
    n1597_o2_p
  );


  buf

  (
    n1128_li039_li039,
    n1598_o2_p
  );


  buf

  (
    n1140_li043_li043,
    n1599_o2_p
  );


  buf

  (
    n1152_li047_li047,
    n1600_o2_p
  );


  buf

  (
    n1164_li051_li051,
    n1601_o2_p
  );


  buf

  (
    n1176_li055_li055,
    n1602_o2_p
  );


  buf

  (
    n1188_li059_li059,
    n1603_o2_p
  );


  buf

  (
    n1200_li063_li063,
    n1604_o2_p
  );


  buf

  (
    n1212_li067_li067,
    n1605_o2_p
  );


  buf

  (
    n1224_li071_li071,
    n1606_o2_p
  );


  buf

  (
    n1236_li075_li075,
    n1607_o2_p
  );


  buf

  (
    n1248_li079_li079,
    n1608_o2_p
  );


  buf

  (
    n1260_li083_li083,
    n1609_o2_p
  );


  buf

  (
    n1272_li087_li087,
    n1610_o2_p
  );


  buf

  (
    n1284_li091_li091,
    n1611_o2_p
  );


  buf

  (
    n1296_li095_li095,
    n1612_o2_p
  );


  buf

  (
    n1308_li099_li099,
    n1613_o2_p
  );


  buf

  (
    n1320_li103_li103,
    n1614_o2_p
  );


  buf

  (
    n1332_li107_li107,
    n1615_o2_p
  );


  buf

  (
    n1344_li111_li111,
    n1616_o2_p
  );


  buf

  (
    n1356_li115_li115,
    n1617_o2_p
  );


  buf

  (
    n1368_li119_li119,
    n1618_o2_p
  );


  buf

  (
    n1380_li123_li123,
    n1619_o2_p
  );


  buf

  (
    n1392_li127_li127,
    n1620_o2_p
  );


  buf

  (
    n1395_li128_li128,
    G33_p
  );


  buf

  (
    n1407_li132_li132,
    G34_p
  );


  buf

  (
    n1419_li136_li136,
    G35_p
  );


  buf

  (
    n1431_li140_li140,
    G36_p
  );


  buf

  (
    n1443_li144_li144,
    G37_p
  );


  buf

  (
    n1455_li148_li148,
    G38_p
  );


  buf

  (
    n1467_li152_li152,
    G39_p
  );


  buf

  (
    n1479_li156_li156,
    G40_p
  );


  buf

  (
    n1491_li160_li160,
    G41_p
  );


  buf

  (
    n1589_i2,
    lo002_buf_o2_p_spl_
  );


  buf

  (
    n1590_i2,
    lo006_buf_o2_p_spl_
  );


  buf

  (
    n1591_i2,
    lo010_buf_o2_p_spl_
  );


  buf

  (
    n1592_i2,
    lo014_buf_o2_p_spl_
  );


  buf

  (
    n1593_i2,
    lo018_buf_o2_p_spl_
  );


  buf

  (
    n1594_i2,
    lo022_buf_o2_p_spl_
  );


  buf

  (
    n1595_i2,
    lo026_buf_o2_p_spl_
  );


  buf

  (
    n1596_i2,
    lo030_buf_o2_p_spl_
  );


  buf

  (
    n1597_i2,
    lo034_buf_o2_p_spl_
  );


  buf

  (
    n1598_i2,
    lo038_buf_o2_p_spl_
  );


  buf

  (
    n1599_i2,
    lo042_buf_o2_p_spl_
  );


  buf

  (
    n1600_i2,
    lo046_buf_o2_p_spl_
  );


  buf

  (
    n1601_i2,
    lo050_buf_o2_p_spl_
  );


  buf

  (
    n1602_i2,
    lo054_buf_o2_p_spl_
  );


  buf

  (
    n1603_i2,
    lo058_buf_o2_p_spl_
  );


  buf

  (
    n1604_i2,
    lo062_buf_o2_p_spl_
  );


  buf

  (
    n1605_i2,
    lo066_buf_o2_p_spl_
  );


  buf

  (
    n1606_i2,
    lo070_buf_o2_p_spl_
  );


  buf

  (
    n1607_i2,
    lo074_buf_o2_p_spl_
  );


  buf

  (
    n1608_i2,
    lo078_buf_o2_p_spl_
  );


  buf

  (
    n1609_i2,
    lo082_buf_o2_p_spl_
  );


  buf

  (
    n1610_i2,
    lo086_buf_o2_p_spl_
  );


  buf

  (
    n1611_i2,
    lo090_buf_o2_p_spl_
  );


  buf

  (
    n1612_i2,
    lo094_buf_o2_p_spl_
  );


  buf

  (
    n1613_i2,
    lo098_buf_o2_p_spl_
  );


  buf

  (
    n1614_i2,
    lo102_buf_o2_p_spl_
  );


  buf

  (
    n1615_i2,
    lo106_buf_o2_p_spl_
  );


  buf

  (
    n1616_i2,
    lo110_buf_o2_p_spl_
  );


  buf

  (
    n1617_i2,
    lo114_buf_o2_p_spl_
  );


  buf

  (
    n1618_i2,
    lo118_buf_o2_p_spl_
  );


  buf

  (
    n1619_i2,
    lo122_buf_o2_p_spl_
  );


  buf

  (
    n1620_i2,
    lo126_buf_o2_p_spl_
  );


  buf

  (
    n602_i2,
    g381_n_spl_
  );


  buf

  (
    n639_i2,
    g382_n_spl_
  );


  buf

  (
    n678_i2,
    g383_n_spl_
  );


  buf

  (
    n658_i2,
    g384_n_spl_
  );


  buf

  (
    n783_i2,
    g385_n_spl_
  );


  buf

  (
    n802_i2,
    g386_n_spl_
  );


  buf

  (
    n726_i2,
    g387_n_spl_
  );


  buf

  (
    n763_i2,
    g388_n_spl_
  );


  not

  (
    n685_i2,
    g389_n_spl_
  );


  not

  (
    n680_i2,
    g390_n_spl_
  );


  not

  (
    n822_i2,
    g391_n_spl_
  );


  buf

  (
    n843_i2,
    g392_n_spl_
  );


  not

  (
    n842_i2,
    g393_n_spl_
  );


  not

  (
    n681_i2,
    g394_n_spl_
  );


  not

  (
    n684_i2,
    g396_n_spl_
  );


  not

  (
    n686_i2,
    g397_n_spl_
  );


  buf

  (
    n823_i2,
    g398_n_spl_
  );


  buf

  (
    lo002_buf_i2,
    lo001_buf_o2_p_spl_
  );


  buf

  (
    lo006_buf_i2,
    lo005_buf_o2_p_spl_
  );


  buf

  (
    lo010_buf_i2,
    lo009_buf_o2_p_spl_
  );


  buf

  (
    lo014_buf_i2,
    lo013_buf_o2_p_spl_
  );


  buf

  (
    lo018_buf_i2,
    lo017_buf_o2_p_spl_
  );


  buf

  (
    lo022_buf_i2,
    lo021_buf_o2_p_spl_
  );


  buf

  (
    lo026_buf_i2,
    lo025_buf_o2_p_spl_
  );


  buf

  (
    lo030_buf_i2,
    lo029_buf_o2_p_spl_
  );


  buf

  (
    lo034_buf_i2,
    lo033_buf_o2_p_spl_
  );


  buf

  (
    lo038_buf_i2,
    lo037_buf_o2_p_spl_
  );


  buf

  (
    lo042_buf_i2,
    lo041_buf_o2_p_spl_
  );


  buf

  (
    lo046_buf_i2,
    lo045_buf_o2_p_spl_
  );


  buf

  (
    lo050_buf_i2,
    lo049_buf_o2_p_spl_
  );


  buf

  (
    lo054_buf_i2,
    lo053_buf_o2_p_spl_
  );


  buf

  (
    lo058_buf_i2,
    lo057_buf_o2_p_spl_
  );


  buf

  (
    lo062_buf_i2,
    lo061_buf_o2_p_spl_
  );


  buf

  (
    lo066_buf_i2,
    lo065_buf_o2_p_spl_
  );


  buf

  (
    lo070_buf_i2,
    lo069_buf_o2_p_spl_
  );


  buf

  (
    lo074_buf_i2,
    lo073_buf_o2_p_spl_
  );


  buf

  (
    lo078_buf_i2,
    lo077_buf_o2_p_spl_
  );


  buf

  (
    lo082_buf_i2,
    lo081_buf_o2_p_spl_
  );


  buf

  (
    lo086_buf_i2,
    lo085_buf_o2_p_spl_
  );


  buf

  (
    lo090_buf_i2,
    lo089_buf_o2_p_spl_
  );


  buf

  (
    lo094_buf_i2,
    lo093_buf_o2_p_spl_
  );


  buf

  (
    lo098_buf_i2,
    lo097_buf_o2_p_spl_
  );


  buf

  (
    lo102_buf_i2,
    lo101_buf_o2_p_spl_
  );


  buf

  (
    lo106_buf_i2,
    lo105_buf_o2_p_spl_
  );


  buf

  (
    lo110_buf_i2,
    lo109_buf_o2_p_spl_
  );


  buf

  (
    lo114_buf_i2,
    lo113_buf_o2_p_spl_
  );


  buf

  (
    lo118_buf_i2,
    lo117_buf_o2_p_spl_
  );


  buf

  (
    lo122_buf_i2,
    lo121_buf_o2_p_spl_
  );


  buf

  (
    lo126_buf_i2,
    lo125_buf_o2_p_spl_
  );


  not

  (
    n683_i2,
    g401_n
  );


  not

  (
    n688_i2,
    g403_n
  );


  buf

  (
    n803_i2,
    g404_p
  );


  buf

  (
    n862_i2,
    g405_p
  );


  buf

  (
    n764_i2,
    g406_p
  );


  buf

  (
    n863_i2,
    g407_p
  );


  buf

  (
    n886_i2,
    g412_p
  );


  not

  (
    n600_i2,
    g429_n
  );


  buf

  (
    n601_i2,
    g430_p
  );


  not

  (
    n637_i2,
    g447_n
  );


  buf

  (
    n638_i2,
    g448_p
  );


  not

  (
    n676_i2,
    g465_n
  );


  buf

  (
    n677_i2,
    g466_p
  );


  not

  (
    n656_i2,
    g483_n
  );


  buf

  (
    n657_i2,
    g484_p
  );


  not

  (
    n781_i2,
    g501_n
  );


  buf

  (
    n782_i2,
    g502_p
  );


  not

  (
    n800_i2,
    g519_n
  );


  buf

  (
    n801_i2,
    g520_p
  );


  not

  (
    n724_i2,
    g537_n
  );


  buf

  (
    n725_i2,
    g538_p
  );


  not

  (
    n761_i2,
    g555_n
  );


  buf

  (
    n762_i2,
    g556_p
  );


  buf

  (
    lo129_buf_i2,
    n661_lo_p
  );


  buf

  (
    lo133_buf_i2,
    n673_lo_p
  );


  buf

  (
    lo137_buf_i2,
    n685_lo_p
  );


  buf

  (
    lo141_buf_i2,
    n697_lo_p
  );


  buf

  (
    lo145_buf_i2,
    n709_lo_p
  );


  buf

  (
    lo149_buf_i2,
    n721_lo_p
  );


  buf

  (
    lo153_buf_i2,
    n733_lo_p
  );


  buf

  (
    lo157_buf_i2,
    n745_lo_p
  );


  buf

  (
    lo161_buf_i2,
    n757_lo_p
  );


  buf

  (
    n708_i2,
    g565_n
  );


  buf

  (
    n745_i2,
    g574_n
  );


  buf

  (
    n717_i2,
    g583_n
  );


  buf

  (
    n754_i2,
    g592_n
  );


  buf

  (
    n584_i2,
    g601_n
  );


  buf

  (
    n593_i2,
    g610_n
  );


  buf

  (
    n630_i2,
    g619_n
  );


  buf

  (
    n621_i2,
    g628_n
  );


  buf

  (
    lo001_buf_i2,
    G1_p
  );


  buf

  (
    lo005_buf_i2,
    G2_p
  );


  buf

  (
    lo009_buf_i2,
    G3_p
  );


  buf

  (
    lo013_buf_i2,
    G4_p
  );


  buf

  (
    lo017_buf_i2,
    G5_p
  );


  buf

  (
    lo021_buf_i2,
    G6_p
  );


  buf

  (
    lo025_buf_i2,
    G7_p
  );


  buf

  (
    lo029_buf_i2,
    G8_p
  );


  buf

  (
    lo033_buf_i2,
    G9_p
  );


  buf

  (
    lo037_buf_i2,
    G10_p
  );


  buf

  (
    lo041_buf_i2,
    G11_p
  );


  buf

  (
    lo045_buf_i2,
    G12_p
  );


  buf

  (
    lo049_buf_i2,
    G13_p
  );


  buf

  (
    lo053_buf_i2,
    G14_p
  );


  buf

  (
    lo057_buf_i2,
    G15_p
  );


  buf

  (
    lo061_buf_i2,
    G16_p
  );


  buf

  (
    lo065_buf_i2,
    G17_p
  );


  buf

  (
    lo069_buf_i2,
    G18_p
  );


  buf

  (
    lo073_buf_i2,
    G19_p
  );


  buf

  (
    lo077_buf_i2,
    G20_p
  );


  buf

  (
    lo081_buf_i2,
    G21_p
  );


  buf

  (
    lo085_buf_i2,
    G22_p
  );


  buf

  (
    lo089_buf_i2,
    G23_p
  );


  buf

  (
    lo093_buf_i2,
    G24_p
  );


  buf

  (
    lo097_buf_i2,
    G25_p
  );


  buf

  (
    lo101_buf_i2,
    G26_p
  );


  buf

  (
    lo105_buf_i2,
    G27_p
  );


  buf

  (
    lo109_buf_i2,
    G28_p
  );


  buf

  (
    lo113_buf_i2,
    G29_p
  );


  buf

  (
    lo117_buf_i2,
    G30_p
  );


  buf

  (
    lo121_buf_i2,
    G31_p
  );


  buf

  (
    lo125_buf_i2,
    G32_p
  );


  buf

  (
    g236_n_spl_,
    g236_n
  );


  buf

  (
    g236_n_spl_0,
    g236_n_spl_
  );


  buf

  (
    g236_n_spl_1,
    g236_n_spl_
  );


  buf

  (
    g236_p_spl_,
    g236_p
  );


  buf

  (
    g236_p_spl_0,
    g236_p_spl_
  );


  buf

  (
    g236_p_spl_1,
    g236_p_spl_
  );


  buf

  (
    n602_o2_p_spl_,
    n602_o2_p
  );


  buf

  (
    n602_o2_p_spl_0,
    n602_o2_p_spl_
  );


  buf

  (
    n602_o2_p_spl_1,
    n602_o2_p_spl_
  );


  buf

  (
    g238_p_spl_,
    g238_p
  );


  buf

  (
    g238_p_spl_0,
    g238_p_spl_
  );


  buf

  (
    g238_p_spl_1,
    g238_p_spl_
  );


  buf

  (
    n602_o2_n_spl_,
    n602_o2_n
  );


  buf

  (
    n602_o2_n_spl_0,
    n602_o2_n_spl_
  );


  buf

  (
    n602_o2_n_spl_1,
    n602_o2_n_spl_
  );


  buf

  (
    g238_n_spl_,
    g238_n
  );


  buf

  (
    g238_n_spl_0,
    g238_n_spl_
  );


  buf

  (
    g238_n_spl_1,
    g238_n_spl_
  );


  buf

  (
    n639_o2_p_spl_,
    n639_o2_p
  );


  buf

  (
    n639_o2_p_spl_0,
    n639_o2_p_spl_
  );


  buf

  (
    n639_o2_p_spl_00,
    n639_o2_p_spl_0
  );


  buf

  (
    n639_o2_p_spl_1,
    n639_o2_p_spl_
  );


  buf

  (
    n639_o2_n_spl_,
    n639_o2_n
  );


  buf

  (
    n639_o2_n_spl_0,
    n639_o2_n_spl_
  );


  buf

  (
    n639_o2_n_spl_00,
    n639_o2_n_spl_0
  );


  buf

  (
    n639_o2_n_spl_1,
    n639_o2_n_spl_
  );


  buf

  (
    n678_o2_p_spl_,
    n678_o2_p
  );


  buf

  (
    n678_o2_p_spl_0,
    n678_o2_p_spl_
  );


  buf

  (
    n678_o2_p_spl_00,
    n678_o2_p_spl_0
  );


  buf

  (
    n678_o2_p_spl_01,
    n678_o2_p_spl_0
  );


  buf

  (
    n678_o2_p_spl_1,
    n678_o2_p_spl_
  );


  buf

  (
    n678_o2_n_spl_,
    n678_o2_n
  );


  buf

  (
    n678_o2_n_spl_0,
    n678_o2_n_spl_
  );


  buf

  (
    n678_o2_n_spl_00,
    n678_o2_n_spl_0
  );


  buf

  (
    n678_o2_n_spl_01,
    n678_o2_n_spl_0
  );


  buf

  (
    n678_o2_n_spl_1,
    n678_o2_n_spl_
  );


  buf

  (
    n658_o2_p_spl_,
    n658_o2_p
  );


  buf

  (
    n658_o2_p_spl_0,
    n658_o2_p_spl_
  );


  buf

  (
    n658_o2_p_spl_1,
    n658_o2_p_spl_
  );


  buf

  (
    n658_o2_n_spl_,
    n658_o2_n
  );


  buf

  (
    n658_o2_n_spl_0,
    n658_o2_n_spl_
  );


  buf

  (
    n658_o2_n_spl_1,
    n658_o2_n_spl_
  );


  buf

  (
    g256_p_spl_,
    g256_p
  );


  buf

  (
    g256_p_spl_0,
    g256_p_spl_
  );


  buf

  (
    g256_p_spl_1,
    g256_p_spl_
  );


  buf

  (
    g256_n_spl_,
    g256_n
  );


  buf

  (
    g256_n_spl_0,
    g256_n_spl_
  );


  buf

  (
    g256_n_spl_1,
    g256_n_spl_
  );


  buf

  (
    g274_p_spl_,
    g274_p
  );


  buf

  (
    g274_p_spl_0,
    g274_p_spl_
  );


  buf

  (
    g274_p_spl_1,
    g274_p_spl_
  );


  buf

  (
    g274_n_spl_,
    g274_n
  );


  buf

  (
    g274_n_spl_0,
    g274_n_spl_
  );


  buf

  (
    g274_n_spl_1,
    g274_n_spl_
  );


  buf

  (
    g292_p_spl_,
    g292_p
  );


  buf

  (
    g292_p_spl_0,
    g292_p_spl_
  );


  buf

  (
    g292_p_spl_1,
    g292_p_spl_
  );


  buf

  (
    g292_n_spl_,
    g292_n
  );


  buf

  (
    g292_n_spl_0,
    g292_n_spl_
  );


  buf

  (
    g292_n_spl_1,
    g292_n_spl_
  );


  buf

  (
    n886_o2_p_spl_,
    n886_o2_p
  );


  buf

  (
    n886_o2_p_spl_0,
    n886_o2_p_spl_
  );


  buf

  (
    n886_o2_p_spl_1,
    n886_o2_p_spl_
  );


  buf

  (
    n886_o2_n_spl_,
    n886_o2_n
  );


  buf

  (
    n886_o2_n_spl_0,
    n886_o2_n_spl_
  );


  buf

  (
    n886_o2_n_spl_1,
    n886_o2_n_spl_
  );


  buf

  (
    n783_o2_p_spl_,
    n783_o2_p
  );


  buf

  (
    n783_o2_p_spl_0,
    n783_o2_p_spl_
  );


  buf

  (
    n783_o2_p_spl_1,
    n783_o2_p_spl_
  );


  buf

  (
    g310_p_spl_,
    g310_p
  );


  buf

  (
    g310_p_spl_0,
    g310_p_spl_
  );


  buf

  (
    g310_p_spl_1,
    g310_p_spl_
  );


  buf

  (
    n783_o2_n_spl_,
    n783_o2_n
  );


  buf

  (
    n783_o2_n_spl_0,
    n783_o2_n_spl_
  );


  buf

  (
    n783_o2_n_spl_1,
    n783_o2_n_spl_
  );


  buf

  (
    g310_n_spl_,
    g310_n
  );


  buf

  (
    g310_n_spl_0,
    g310_n_spl_
  );


  buf

  (
    g310_n_spl_1,
    g310_n_spl_
  );


  buf

  (
    n802_o2_p_spl_,
    n802_o2_p
  );


  buf

  (
    n802_o2_p_spl_0,
    n802_o2_p_spl_
  );


  buf

  (
    n802_o2_p_spl_1,
    n802_o2_p_spl_
  );


  buf

  (
    n802_o2_n_spl_,
    n802_o2_n
  );


  buf

  (
    n802_o2_n_spl_0,
    n802_o2_n_spl_
  );


  buf

  (
    n802_o2_n_spl_1,
    n802_o2_n_spl_
  );


  buf

  (
    n726_o2_p_spl_,
    n726_o2_p
  );


  buf

  (
    n726_o2_p_spl_0,
    n726_o2_p_spl_
  );


  buf

  (
    n726_o2_p_spl_1,
    n726_o2_p_spl_
  );


  buf

  (
    n726_o2_n_spl_,
    n726_o2_n
  );


  buf

  (
    n726_o2_n_spl_0,
    n726_o2_n_spl_
  );


  buf

  (
    n726_o2_n_spl_1,
    n726_o2_n_spl_
  );


  buf

  (
    n763_o2_p_spl_,
    n763_o2_p
  );


  buf

  (
    n763_o2_p_spl_0,
    n763_o2_p_spl_
  );


  buf

  (
    n763_o2_p_spl_1,
    n763_o2_p_spl_
  );


  buf

  (
    n763_o2_n_spl_,
    n763_o2_n
  );


  buf

  (
    n763_o2_n_spl_0,
    n763_o2_n_spl_
  );


  buf

  (
    n763_o2_n_spl_1,
    n763_o2_n_spl_
  );


  buf

  (
    g328_p_spl_,
    g328_p
  );


  buf

  (
    g328_p_spl_0,
    g328_p_spl_
  );


  buf

  (
    g328_p_spl_1,
    g328_p_spl_
  );


  buf

  (
    g328_n_spl_,
    g328_n
  );


  buf

  (
    g328_n_spl_0,
    g328_n_spl_
  );


  buf

  (
    g328_n_spl_1,
    g328_n_spl_
  );


  buf

  (
    g346_p_spl_,
    g346_p
  );


  buf

  (
    g346_p_spl_0,
    g346_p_spl_
  );


  buf

  (
    g346_p_spl_1,
    g346_p_spl_
  );


  buf

  (
    g346_n_spl_,
    g346_n
  );


  buf

  (
    g346_n_spl_0,
    g346_n_spl_
  );


  buf

  (
    g346_n_spl_1,
    g346_n_spl_
  );


  buf

  (
    g364_p_spl_,
    g364_p
  );


  buf

  (
    g364_p_spl_0,
    g364_p_spl_
  );


  buf

  (
    g364_p_spl_1,
    g364_p_spl_
  );


  buf

  (
    g364_n_spl_,
    g364_n
  );


  buf

  (
    g364_n_spl_0,
    g364_n_spl_
  );


  buf

  (
    g364_n_spl_1,
    g364_n_spl_
  );


  buf

  (
    g382_n_spl_,
    g382_n
  );


  buf

  (
    g382_n_spl_0,
    g382_n_spl_
  );


  buf

  (
    g383_n_spl_,
    g383_n
  );


  buf

  (
    g383_n_spl_0,
    g383_n_spl_
  );


  buf

  (
    g385_p_spl_,
    g385_p
  );


  buf

  (
    g385_p_spl_0,
    g385_p_spl_
  );


  buf

  (
    g388_p_spl_,
    g388_p
  );


  buf

  (
    g388_p_spl_0,
    g388_p_spl_
  );


  buf

  (
    g385_n_spl_,
    g385_n
  );


  buf

  (
    g385_n_spl_0,
    g385_n_spl_
  );


  buf

  (
    g388_n_spl_,
    g388_n
  );


  buf

  (
    g388_n_spl_0,
    g388_n_spl_
  );


  buf

  (
    g386_p_spl_,
    g386_p
  );


  buf

  (
    g386_p_spl_0,
    g386_p_spl_
  );


  buf

  (
    g387_p_spl_,
    g387_p
  );


  buf

  (
    g387_p_spl_0,
    g387_p_spl_
  );


  buf

  (
    g381_n_spl_,
    g381_n
  );


  buf

  (
    g381_n_spl_0,
    g381_n_spl_
  );


  buf

  (
    g390_n_spl_,
    g390_n
  );


  buf

  (
    g384_n_spl_,
    g384_n
  );


  buf

  (
    g384_n_spl_0,
    g384_n_spl_
  );


  buf

  (
    g395_n_spl_,
    g395_n
  );


  buf

  (
    g389_n_spl_,
    g389_n
  );


  buf

  (
    g386_n_spl_,
    g386_n
  );


  buf

  (
    g386_n_spl_0,
    g386_n_spl_
  );


  buf

  (
    g387_n_spl_,
    g387_n
  );


  buf

  (
    g387_n_spl_0,
    g387_n_spl_
  );


  buf

  (
    g394_n_spl_,
    g394_n
  );


  buf

  (
    g396_n_spl_,
    g396_n
  );


  buf

  (
    g397_n_spl_,
    g397_n
  );


  buf

  (
    g391_n_spl_,
    g391_n
  );


  buf

  (
    g392_n_spl_,
    g392_n
  );


  buf

  (
    g398_n_spl_,
    g398_n
  );


  buf

  (
    g393_n_spl_,
    g393_n
  );


  buf

  (
    lo002_buf_o2_p_spl_,
    lo002_buf_o2_p
  );


  buf

  (
    lo002_buf_o2_p_spl_0,
    lo002_buf_o2_p_spl_
  );


  buf

  (
    lo018_buf_o2_n_spl_,
    lo018_buf_o2_n
  );


  buf

  (
    lo002_buf_o2_n_spl_,
    lo002_buf_o2_n
  );


  buf

  (
    lo018_buf_o2_p_spl_,
    lo018_buf_o2_p
  );


  buf

  (
    lo018_buf_o2_p_spl_0,
    lo018_buf_o2_p_spl_
  );


  buf

  (
    lo034_buf_o2_p_spl_,
    lo034_buf_o2_p
  );


  buf

  (
    lo034_buf_o2_p_spl_0,
    lo034_buf_o2_p_spl_
  );


  buf

  (
    lo050_buf_o2_n_spl_,
    lo050_buf_o2_n
  );


  buf

  (
    lo034_buf_o2_n_spl_,
    lo034_buf_o2_n
  );


  buf

  (
    lo050_buf_o2_p_spl_,
    lo050_buf_o2_p
  );


  buf

  (
    lo050_buf_o2_p_spl_0,
    lo050_buf_o2_p_spl_
  );


  buf

  (
    lo161_buf_o2_p_spl_,
    lo161_buf_o2_p
  );


  buf

  (
    lo161_buf_o2_p_spl_0,
    lo161_buf_o2_p_spl_
  );


  buf

  (
    lo161_buf_o2_p_spl_00,
    lo161_buf_o2_p_spl_0
  );


  buf

  (
    lo161_buf_o2_p_spl_01,
    lo161_buf_o2_p_spl_0
  );


  buf

  (
    lo161_buf_o2_p_spl_1,
    lo161_buf_o2_p_spl_
  );


  buf

  (
    lo161_buf_o2_p_spl_10,
    lo161_buf_o2_p_spl_1
  );


  buf

  (
    lo161_buf_o2_p_spl_11,
    lo161_buf_o2_p_spl_1
  );


  buf

  (
    lo161_buf_o2_n_spl_,
    lo161_buf_o2_n
  );


  buf

  (
    lo161_buf_o2_n_spl_0,
    lo161_buf_o2_n_spl_
  );


  buf

  (
    lo161_buf_o2_n_spl_00,
    lo161_buf_o2_n_spl_0
  );


  buf

  (
    lo161_buf_o2_n_spl_01,
    lo161_buf_o2_n_spl_0
  );


  buf

  (
    lo161_buf_o2_n_spl_1,
    lo161_buf_o2_n_spl_
  );


  buf

  (
    lo161_buf_o2_n_spl_10,
    lo161_buf_o2_n_spl_1
  );


  buf

  (
    lo161_buf_o2_n_spl_11,
    lo161_buf_o2_n_spl_1
  );


  buf

  (
    n584_o2_n_spl_,
    n584_o2_n
  );


  buf

  (
    n584_o2_n_spl_0,
    n584_o2_n_spl_
  );


  buf

  (
    n584_o2_n_spl_1,
    n584_o2_n_spl_
  );


  buf

  (
    n593_o2_p_spl_,
    n593_o2_p
  );


  buf

  (
    n593_o2_p_spl_0,
    n593_o2_p_spl_
  );


  buf

  (
    n593_o2_p_spl_1,
    n593_o2_p_spl_
  );


  buf

  (
    n584_o2_p_spl_,
    n584_o2_p
  );


  buf

  (
    n584_o2_p_spl_0,
    n584_o2_p_spl_
  );


  buf

  (
    n584_o2_p_spl_1,
    n584_o2_p_spl_
  );


  buf

  (
    n593_o2_n_spl_,
    n593_o2_n
  );


  buf

  (
    n593_o2_n_spl_0,
    n593_o2_n_spl_
  );


  buf

  (
    n593_o2_n_spl_1,
    n593_o2_n_spl_
  );


  buf

  (
    g421_n_spl_,
    g421_n
  );


  buf

  (
    g428_p_spl_,
    g428_p
  );


  buf

  (
    lo006_buf_o2_p_spl_,
    lo006_buf_o2_p
  );


  buf

  (
    lo006_buf_o2_p_spl_0,
    lo006_buf_o2_p_spl_
  );


  buf

  (
    lo022_buf_o2_n_spl_,
    lo022_buf_o2_n
  );


  buf

  (
    lo006_buf_o2_n_spl_,
    lo006_buf_o2_n
  );


  buf

  (
    lo022_buf_o2_p_spl_,
    lo022_buf_o2_p
  );


  buf

  (
    lo022_buf_o2_p_spl_0,
    lo022_buf_o2_p_spl_
  );


  buf

  (
    lo038_buf_o2_p_spl_,
    lo038_buf_o2_p
  );


  buf

  (
    lo038_buf_o2_p_spl_0,
    lo038_buf_o2_p_spl_
  );


  buf

  (
    lo054_buf_o2_n_spl_,
    lo054_buf_o2_n
  );


  buf

  (
    lo038_buf_o2_n_spl_,
    lo038_buf_o2_n
  );


  buf

  (
    lo054_buf_o2_p_spl_,
    lo054_buf_o2_p
  );


  buf

  (
    lo054_buf_o2_p_spl_0,
    lo054_buf_o2_p_spl_
  );


  buf

  (
    n630_o2_p_spl_,
    n630_o2_p
  );


  buf

  (
    n630_o2_p_spl_0,
    n630_o2_p_spl_
  );


  buf

  (
    n630_o2_p_spl_1,
    n630_o2_p_spl_
  );


  buf

  (
    n621_o2_n_spl_,
    n621_o2_n
  );


  buf

  (
    n621_o2_n_spl_0,
    n621_o2_n_spl_
  );


  buf

  (
    n621_o2_n_spl_1,
    n621_o2_n_spl_
  );


  buf

  (
    n630_o2_n_spl_,
    n630_o2_n
  );


  buf

  (
    n630_o2_n_spl_0,
    n630_o2_n_spl_
  );


  buf

  (
    n630_o2_n_spl_1,
    n630_o2_n_spl_
  );


  buf

  (
    n621_o2_p_spl_,
    n621_o2_p
  );


  buf

  (
    n621_o2_p_spl_0,
    n621_o2_p_spl_
  );


  buf

  (
    n621_o2_p_spl_1,
    n621_o2_p_spl_
  );


  buf

  (
    g439_n_spl_,
    g439_n
  );


  buf

  (
    g446_p_spl_,
    g446_p
  );


  buf

  (
    lo010_buf_o2_p_spl_,
    lo010_buf_o2_p
  );


  buf

  (
    lo010_buf_o2_p_spl_0,
    lo010_buf_o2_p_spl_
  );


  buf

  (
    lo026_buf_o2_n_spl_,
    lo026_buf_o2_n
  );


  buf

  (
    lo010_buf_o2_n_spl_,
    lo010_buf_o2_n
  );


  buf

  (
    lo026_buf_o2_p_spl_,
    lo026_buf_o2_p
  );


  buf

  (
    lo026_buf_o2_p_spl_0,
    lo026_buf_o2_p_spl_
  );


  buf

  (
    lo042_buf_o2_p_spl_,
    lo042_buf_o2_p
  );


  buf

  (
    lo042_buf_o2_p_spl_0,
    lo042_buf_o2_p_spl_
  );


  buf

  (
    lo058_buf_o2_n_spl_,
    lo058_buf_o2_n
  );


  buf

  (
    lo042_buf_o2_n_spl_,
    lo042_buf_o2_n
  );


  buf

  (
    lo058_buf_o2_p_spl_,
    lo058_buf_o2_p
  );


  buf

  (
    lo058_buf_o2_p_spl_0,
    lo058_buf_o2_p_spl_
  );


  buf

  (
    g457_n_spl_,
    g457_n
  );


  buf

  (
    g464_p_spl_,
    g464_p
  );


  buf

  (
    lo014_buf_o2_p_spl_,
    lo014_buf_o2_p
  );


  buf

  (
    lo014_buf_o2_p_spl_0,
    lo014_buf_o2_p_spl_
  );


  buf

  (
    lo030_buf_o2_n_spl_,
    lo030_buf_o2_n
  );


  buf

  (
    lo014_buf_o2_n_spl_,
    lo014_buf_o2_n
  );


  buf

  (
    lo030_buf_o2_p_spl_,
    lo030_buf_o2_p
  );


  buf

  (
    lo030_buf_o2_p_spl_0,
    lo030_buf_o2_p_spl_
  );


  buf

  (
    lo046_buf_o2_p_spl_,
    lo046_buf_o2_p
  );


  buf

  (
    lo046_buf_o2_p_spl_0,
    lo046_buf_o2_p_spl_
  );


  buf

  (
    lo062_buf_o2_n_spl_,
    lo062_buf_o2_n
  );


  buf

  (
    lo046_buf_o2_n_spl_,
    lo046_buf_o2_n
  );


  buf

  (
    lo062_buf_o2_p_spl_,
    lo062_buf_o2_p
  );


  buf

  (
    lo062_buf_o2_p_spl_0,
    lo062_buf_o2_p_spl_
  );


  buf

  (
    g475_n_spl_,
    g475_n
  );


  buf

  (
    g482_p_spl_,
    g482_p
  );


  buf

  (
    lo066_buf_o2_p_spl_,
    lo066_buf_o2_p
  );


  buf

  (
    lo066_buf_o2_p_spl_0,
    lo066_buf_o2_p_spl_
  );


  buf

  (
    lo082_buf_o2_n_spl_,
    lo082_buf_o2_n
  );


  buf

  (
    lo066_buf_o2_n_spl_,
    lo066_buf_o2_n
  );


  buf

  (
    lo082_buf_o2_p_spl_,
    lo082_buf_o2_p
  );


  buf

  (
    lo082_buf_o2_p_spl_0,
    lo082_buf_o2_p_spl_
  );


  buf

  (
    lo098_buf_o2_p_spl_,
    lo098_buf_o2_p
  );


  buf

  (
    lo098_buf_o2_p_spl_0,
    lo098_buf_o2_p_spl_
  );


  buf

  (
    lo114_buf_o2_n_spl_,
    lo114_buf_o2_n
  );


  buf

  (
    lo098_buf_o2_n_spl_,
    lo098_buf_o2_n
  );


  buf

  (
    lo114_buf_o2_p_spl_,
    lo114_buf_o2_p
  );


  buf

  (
    lo114_buf_o2_p_spl_0,
    lo114_buf_o2_p_spl_
  );


  buf

  (
    n708_o2_n_spl_,
    n708_o2_n
  );


  buf

  (
    n708_o2_n_spl_0,
    n708_o2_n_spl_
  );


  buf

  (
    n708_o2_n_spl_1,
    n708_o2_n_spl_
  );


  buf

  (
    n745_o2_p_spl_,
    n745_o2_p
  );


  buf

  (
    n745_o2_p_spl_0,
    n745_o2_p_spl_
  );


  buf

  (
    n745_o2_p_spl_1,
    n745_o2_p_spl_
  );


  buf

  (
    n708_o2_p_spl_,
    n708_o2_p
  );


  buf

  (
    n708_o2_p_spl_0,
    n708_o2_p_spl_
  );


  buf

  (
    n708_o2_p_spl_1,
    n708_o2_p_spl_
  );


  buf

  (
    n745_o2_n_spl_,
    n745_o2_n
  );


  buf

  (
    n745_o2_n_spl_0,
    n745_o2_n_spl_
  );


  buf

  (
    n745_o2_n_spl_1,
    n745_o2_n_spl_
  );


  buf

  (
    g493_n_spl_,
    g493_n
  );


  buf

  (
    g500_p_spl_,
    g500_p
  );


  buf

  (
    lo070_buf_o2_p_spl_,
    lo070_buf_o2_p
  );


  buf

  (
    lo070_buf_o2_p_spl_0,
    lo070_buf_o2_p_spl_
  );


  buf

  (
    lo086_buf_o2_n_spl_,
    lo086_buf_o2_n
  );


  buf

  (
    lo070_buf_o2_n_spl_,
    lo070_buf_o2_n
  );


  buf

  (
    lo086_buf_o2_p_spl_,
    lo086_buf_o2_p
  );


  buf

  (
    lo086_buf_o2_p_spl_0,
    lo086_buf_o2_p_spl_
  );


  buf

  (
    lo102_buf_o2_p_spl_,
    lo102_buf_o2_p
  );


  buf

  (
    lo102_buf_o2_p_spl_0,
    lo102_buf_o2_p_spl_
  );


  buf

  (
    lo118_buf_o2_n_spl_,
    lo118_buf_o2_n
  );


  buf

  (
    lo102_buf_o2_n_spl_,
    lo102_buf_o2_n
  );


  buf

  (
    lo118_buf_o2_p_spl_,
    lo118_buf_o2_p
  );


  buf

  (
    lo118_buf_o2_p_spl_0,
    lo118_buf_o2_p_spl_
  );


  buf

  (
    n717_o2_n_spl_,
    n717_o2_n
  );


  buf

  (
    n717_o2_n_spl_0,
    n717_o2_n_spl_
  );


  buf

  (
    n717_o2_n_spl_1,
    n717_o2_n_spl_
  );


  buf

  (
    n754_o2_p_spl_,
    n754_o2_p
  );


  buf

  (
    n754_o2_p_spl_0,
    n754_o2_p_spl_
  );


  buf

  (
    n754_o2_p_spl_1,
    n754_o2_p_spl_
  );


  buf

  (
    n717_o2_p_spl_,
    n717_o2_p
  );


  buf

  (
    n717_o2_p_spl_0,
    n717_o2_p_spl_
  );


  buf

  (
    n717_o2_p_spl_1,
    n717_o2_p_spl_
  );


  buf

  (
    n754_o2_n_spl_,
    n754_o2_n
  );


  buf

  (
    n754_o2_n_spl_0,
    n754_o2_n_spl_
  );


  buf

  (
    n754_o2_n_spl_1,
    n754_o2_n_spl_
  );


  buf

  (
    g511_n_spl_,
    g511_n
  );


  buf

  (
    g518_p_spl_,
    g518_p
  );


  buf

  (
    lo074_buf_o2_p_spl_,
    lo074_buf_o2_p
  );


  buf

  (
    lo074_buf_o2_p_spl_0,
    lo074_buf_o2_p_spl_
  );


  buf

  (
    lo090_buf_o2_n_spl_,
    lo090_buf_o2_n
  );


  buf

  (
    lo074_buf_o2_n_spl_,
    lo074_buf_o2_n
  );


  buf

  (
    lo090_buf_o2_p_spl_,
    lo090_buf_o2_p
  );


  buf

  (
    lo090_buf_o2_p_spl_0,
    lo090_buf_o2_p_spl_
  );


  buf

  (
    lo106_buf_o2_p_spl_,
    lo106_buf_o2_p
  );


  buf

  (
    lo106_buf_o2_p_spl_0,
    lo106_buf_o2_p_spl_
  );


  buf

  (
    lo122_buf_o2_n_spl_,
    lo122_buf_o2_n
  );


  buf

  (
    lo106_buf_o2_n_spl_,
    lo106_buf_o2_n
  );


  buf

  (
    lo122_buf_o2_p_spl_,
    lo122_buf_o2_p
  );


  buf

  (
    lo122_buf_o2_p_spl_0,
    lo122_buf_o2_p_spl_
  );


  buf

  (
    g529_n_spl_,
    g529_n
  );


  buf

  (
    g536_p_spl_,
    g536_p
  );


  buf

  (
    lo078_buf_o2_p_spl_,
    lo078_buf_o2_p
  );


  buf

  (
    lo078_buf_o2_p_spl_0,
    lo078_buf_o2_p_spl_
  );


  buf

  (
    lo094_buf_o2_n_spl_,
    lo094_buf_o2_n
  );


  buf

  (
    lo078_buf_o2_n_spl_,
    lo078_buf_o2_n
  );


  buf

  (
    lo094_buf_o2_p_spl_,
    lo094_buf_o2_p
  );


  buf

  (
    lo094_buf_o2_p_spl_0,
    lo094_buf_o2_p_spl_
  );


  buf

  (
    lo110_buf_o2_p_spl_,
    lo110_buf_o2_p
  );


  buf

  (
    lo110_buf_o2_p_spl_0,
    lo110_buf_o2_p_spl_
  );


  buf

  (
    lo126_buf_o2_n_spl_,
    lo126_buf_o2_n
  );


  buf

  (
    lo110_buf_o2_n_spl_,
    lo110_buf_o2_n
  );


  buf

  (
    lo126_buf_o2_p_spl_,
    lo126_buf_o2_p
  );


  buf

  (
    lo126_buf_o2_p_spl_0,
    lo126_buf_o2_p_spl_
  );


  buf

  (
    g547_n_spl_,
    g547_n
  );


  buf

  (
    g554_p_spl_,
    g554_p
  );


  buf

  (
    lo001_buf_o2_p_spl_,
    lo001_buf_o2_p
  );


  buf

  (
    lo001_buf_o2_p_spl_0,
    lo001_buf_o2_p_spl_
  );


  buf

  (
    lo005_buf_o2_n_spl_,
    lo005_buf_o2_n
  );


  buf

  (
    lo001_buf_o2_n_spl_,
    lo001_buf_o2_n
  );


  buf

  (
    lo005_buf_o2_p_spl_,
    lo005_buf_o2_p
  );


  buf

  (
    lo005_buf_o2_p_spl_0,
    lo005_buf_o2_p_spl_
  );


  buf

  (
    lo009_buf_o2_p_spl_,
    lo009_buf_o2_p
  );


  buf

  (
    lo009_buf_o2_p_spl_0,
    lo009_buf_o2_p_spl_
  );


  buf

  (
    lo013_buf_o2_n_spl_,
    lo013_buf_o2_n
  );


  buf

  (
    lo009_buf_o2_n_spl_,
    lo009_buf_o2_n
  );


  buf

  (
    lo013_buf_o2_p_spl_,
    lo013_buf_o2_p
  );


  buf

  (
    lo013_buf_o2_p_spl_0,
    lo013_buf_o2_p_spl_
  );


  buf

  (
    lo017_buf_o2_p_spl_,
    lo017_buf_o2_p
  );


  buf

  (
    lo017_buf_o2_p_spl_0,
    lo017_buf_o2_p_spl_
  );


  buf

  (
    lo021_buf_o2_n_spl_,
    lo021_buf_o2_n
  );


  buf

  (
    lo017_buf_o2_n_spl_,
    lo017_buf_o2_n
  );


  buf

  (
    lo021_buf_o2_p_spl_,
    lo021_buf_o2_p
  );


  buf

  (
    lo021_buf_o2_p_spl_0,
    lo021_buf_o2_p_spl_
  );


  buf

  (
    lo025_buf_o2_p_spl_,
    lo025_buf_o2_p
  );


  buf

  (
    lo025_buf_o2_p_spl_0,
    lo025_buf_o2_p_spl_
  );


  buf

  (
    lo029_buf_o2_n_spl_,
    lo029_buf_o2_n
  );


  buf

  (
    lo025_buf_o2_n_spl_,
    lo025_buf_o2_n
  );


  buf

  (
    lo029_buf_o2_p_spl_,
    lo029_buf_o2_p
  );


  buf

  (
    lo029_buf_o2_p_spl_0,
    lo029_buf_o2_p_spl_
  );


  buf

  (
    lo033_buf_o2_p_spl_,
    lo033_buf_o2_p
  );


  buf

  (
    lo033_buf_o2_p_spl_0,
    lo033_buf_o2_p_spl_
  );


  buf

  (
    lo037_buf_o2_n_spl_,
    lo037_buf_o2_n
  );


  buf

  (
    lo033_buf_o2_n_spl_,
    lo033_buf_o2_n
  );


  buf

  (
    lo037_buf_o2_p_spl_,
    lo037_buf_o2_p
  );


  buf

  (
    lo037_buf_o2_p_spl_0,
    lo037_buf_o2_p_spl_
  );


  buf

  (
    lo041_buf_o2_p_spl_,
    lo041_buf_o2_p
  );


  buf

  (
    lo041_buf_o2_p_spl_0,
    lo041_buf_o2_p_spl_
  );


  buf

  (
    lo045_buf_o2_n_spl_,
    lo045_buf_o2_n
  );


  buf

  (
    lo041_buf_o2_n_spl_,
    lo041_buf_o2_n
  );


  buf

  (
    lo045_buf_o2_p_spl_,
    lo045_buf_o2_p
  );


  buf

  (
    lo045_buf_o2_p_spl_0,
    lo045_buf_o2_p_spl_
  );


  buf

  (
    lo049_buf_o2_p_spl_,
    lo049_buf_o2_p
  );


  buf

  (
    lo049_buf_o2_p_spl_0,
    lo049_buf_o2_p_spl_
  );


  buf

  (
    lo053_buf_o2_n_spl_,
    lo053_buf_o2_n
  );


  buf

  (
    lo049_buf_o2_n_spl_,
    lo049_buf_o2_n
  );


  buf

  (
    lo053_buf_o2_p_spl_,
    lo053_buf_o2_p
  );


  buf

  (
    lo053_buf_o2_p_spl_0,
    lo053_buf_o2_p_spl_
  );


  buf

  (
    lo057_buf_o2_p_spl_,
    lo057_buf_o2_p
  );


  buf

  (
    lo057_buf_o2_p_spl_0,
    lo057_buf_o2_p_spl_
  );


  buf

  (
    lo061_buf_o2_n_spl_,
    lo061_buf_o2_n
  );


  buf

  (
    lo057_buf_o2_n_spl_,
    lo057_buf_o2_n
  );


  buf

  (
    lo061_buf_o2_p_spl_,
    lo061_buf_o2_p
  );


  buf

  (
    lo061_buf_o2_p_spl_0,
    lo061_buf_o2_p_spl_
  );


  buf

  (
    lo065_buf_o2_p_spl_,
    lo065_buf_o2_p
  );


  buf

  (
    lo065_buf_o2_p_spl_0,
    lo065_buf_o2_p_spl_
  );


  buf

  (
    lo069_buf_o2_n_spl_,
    lo069_buf_o2_n
  );


  buf

  (
    lo065_buf_o2_n_spl_,
    lo065_buf_o2_n
  );


  buf

  (
    lo069_buf_o2_p_spl_,
    lo069_buf_o2_p
  );


  buf

  (
    lo069_buf_o2_p_spl_0,
    lo069_buf_o2_p_spl_
  );


  buf

  (
    lo073_buf_o2_p_spl_,
    lo073_buf_o2_p
  );


  buf

  (
    lo073_buf_o2_p_spl_0,
    lo073_buf_o2_p_spl_
  );


  buf

  (
    lo077_buf_o2_n_spl_,
    lo077_buf_o2_n
  );


  buf

  (
    lo073_buf_o2_n_spl_,
    lo073_buf_o2_n
  );


  buf

  (
    lo077_buf_o2_p_spl_,
    lo077_buf_o2_p
  );


  buf

  (
    lo077_buf_o2_p_spl_0,
    lo077_buf_o2_p_spl_
  );


  buf

  (
    lo081_buf_o2_p_spl_,
    lo081_buf_o2_p
  );


  buf

  (
    lo081_buf_o2_p_spl_0,
    lo081_buf_o2_p_spl_
  );


  buf

  (
    lo085_buf_o2_n_spl_,
    lo085_buf_o2_n
  );


  buf

  (
    lo081_buf_o2_n_spl_,
    lo081_buf_o2_n
  );


  buf

  (
    lo085_buf_o2_p_spl_,
    lo085_buf_o2_p
  );


  buf

  (
    lo085_buf_o2_p_spl_0,
    lo085_buf_o2_p_spl_
  );


  buf

  (
    lo089_buf_o2_p_spl_,
    lo089_buf_o2_p
  );


  buf

  (
    lo089_buf_o2_p_spl_0,
    lo089_buf_o2_p_spl_
  );


  buf

  (
    lo093_buf_o2_n_spl_,
    lo093_buf_o2_n
  );


  buf

  (
    lo089_buf_o2_n_spl_,
    lo089_buf_o2_n
  );


  buf

  (
    lo093_buf_o2_p_spl_,
    lo093_buf_o2_p
  );


  buf

  (
    lo093_buf_o2_p_spl_0,
    lo093_buf_o2_p_spl_
  );


  buf

  (
    lo097_buf_o2_p_spl_,
    lo097_buf_o2_p
  );


  buf

  (
    lo097_buf_o2_p_spl_0,
    lo097_buf_o2_p_spl_
  );


  buf

  (
    lo101_buf_o2_n_spl_,
    lo101_buf_o2_n
  );


  buf

  (
    lo097_buf_o2_n_spl_,
    lo097_buf_o2_n
  );


  buf

  (
    lo101_buf_o2_p_spl_,
    lo101_buf_o2_p
  );


  buf

  (
    lo101_buf_o2_p_spl_0,
    lo101_buf_o2_p_spl_
  );


  buf

  (
    lo105_buf_o2_p_spl_,
    lo105_buf_o2_p
  );


  buf

  (
    lo105_buf_o2_p_spl_0,
    lo105_buf_o2_p_spl_
  );


  buf

  (
    lo109_buf_o2_n_spl_,
    lo109_buf_o2_n
  );


  buf

  (
    lo105_buf_o2_n_spl_,
    lo105_buf_o2_n
  );


  buf

  (
    lo109_buf_o2_p_spl_,
    lo109_buf_o2_p
  );


  buf

  (
    lo109_buf_o2_p_spl_0,
    lo109_buf_o2_p_spl_
  );


  buf

  (
    lo113_buf_o2_p_spl_,
    lo113_buf_o2_p
  );


  buf

  (
    lo113_buf_o2_p_spl_0,
    lo113_buf_o2_p_spl_
  );


  buf

  (
    lo117_buf_o2_n_spl_,
    lo117_buf_o2_n
  );


  buf

  (
    lo113_buf_o2_n_spl_,
    lo113_buf_o2_n
  );


  buf

  (
    lo117_buf_o2_p_spl_,
    lo117_buf_o2_p
  );


  buf

  (
    lo117_buf_o2_p_spl_0,
    lo117_buf_o2_p_spl_
  );


  buf

  (
    lo121_buf_o2_p_spl_,
    lo121_buf_o2_p
  );


  buf

  (
    lo121_buf_o2_p_spl_0,
    lo121_buf_o2_p_spl_
  );


  buf

  (
    lo125_buf_o2_n_spl_,
    lo125_buf_o2_n
  );


  buf

  (
    lo121_buf_o2_n_spl_,
    lo121_buf_o2_n
  );


  buf

  (
    lo125_buf_o2_p_spl_,
    lo125_buf_o2_p
  );


  buf

  (
    lo125_buf_o2_p_spl_0,
    lo125_buf_o2_p_spl_
  );


endmodule
