// Benchmark "c3540" written by ABC on Sun Oct 29 22:18:02 2023

module c3540 ( 
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50,
    G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528,
    G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538,
    G3539, G3540  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50;
  output G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528,
    G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538,
    G3539, G3540;
  wire new_n73_, new_n74_, new_n76_, new_n78_, new_n79_, new_n80_, new_n81_,
    new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_,
    new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_,
    new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n133_,
    new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_,
    new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_,
    new_n146_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_;
  nor1 g000(.dina(G7), .dinb(G8), .dout(new_n73_));
  anb1 g001(.dina(new_n73_), .dinb(G9), .dout(new_n74_));
  anb1 g002(.dina(new_n74_), .dinb(G10), .dout(G3519));
  nor1 g003(.dina(G12), .dinb(G13), .dout(new_n76_));
  anb2 g004(.dina(new_n76_), .dinb(G11), .dout(G3520));
  nor1 g005(.dina(G1), .dinb(G3), .dout(new_n78_));
  anb1 g006(.dina(G34), .dinb(G11), .dout(new_n79_));
  anb2 g007(.dina(G9), .dinb(G32), .dout(new_n80_));
  anb2 g008(.dina(new_n79_), .dinb(new_n80_), .dout(new_n81_));
  anb2 g009(.dina(G7), .dinb(G30), .dout(new_n82_));
  anb1 g010(.dina(G33), .dinb(G10), .dout(new_n83_));
  anb1 g011(.dina(new_n82_), .dinb(new_n83_), .dout(new_n84_));
  anb2 g012(.dina(new_n81_), .dinb(new_n84_), .dout(new_n85_));
  anb2 g013(.dina(G14), .dinb(G37), .dout(new_n86_));
  anb1 g014(.dina(G31), .dinb(G8), .dout(new_n87_));
  anb1 g015(.dina(new_n86_), .dinb(new_n87_), .dout(new_n88_));
  anb1 g016(.dina(G35), .dinb(G12), .dout(new_n89_));
  anb2 g017(.dina(G13), .dinb(G36), .dout(new_n90_));
  anb2 g018(.dina(new_n89_), .dinb(new_n90_), .dout(new_n91_));
  anb1 g019(.dina(new_n88_), .dinb(new_n91_), .dout(new_n92_));
  anb2 g020(.dina(new_n85_), .dinb(new_n92_), .dout(new_n93_));
  anb2 g021(.dina(new_n78_), .dinb(new_n93_), .dout(new_n94_));
  anb2 g022(.dina(G1), .dinb(G2), .dout(new_n95_));
  nor1 g023(.dina(G3), .dinb(new_n95_), .dout(new_n96_));
  and2 g024(.dina(G8), .dinb(G9), .dout(new_n97_));
  nab1 g025(.dina(G7), .dinb(new_n97_), .dout(new_n98_));
  and1 g026(.dina(new_n96_), .dinb(new_n98_), .dout(new_n99_));
  and2 g027(.dina(G1), .dinb(G2), .dout(new_n100_));
  and2 g028(.dina(G3), .dinb(new_n100_), .dout(new_n101_));
  nor1 g029(.dina(G35), .dinb(G36), .dout(new_n102_));
  anb1 g030(.dina(G34), .dinb(new_n102_), .dout(new_n103_));
  anb2 g031(.dina(new_n101_), .dinb(new_n103_), .dout(new_n104_));
  anb2 g032(.dina(new_n99_), .dinb(new_n104_), .dout(new_n105_));
  anb1 g033(.dina(new_n94_), .dinb(new_n105_), .dout(G3521));
  anb2 g034(.dina(G37), .dinb(G36), .dout(new_n107_));
  anb1 g035(.dina(G37), .dinb(G36), .dout(new_n108_));
  anb1 g036(.dina(new_n107_), .dinb(new_n108_), .dout(new_n109_));
  anb2 g037(.dina(G35), .dinb(G34), .dout(new_n110_));
  anb1 g038(.dina(G35), .dinb(G34), .dout(new_n111_));
  anb1 g039(.dina(new_n110_), .dinb(new_n111_), .dout(new_n112_));
  anb2 g040(.dina(new_n109_), .dinb(new_n112_), .dout(new_n113_));
  anb1 g041(.dina(new_n109_), .dinb(new_n112_), .dout(new_n114_));
  anb1 g042(.dina(new_n113_), .dinb(new_n114_), .dout(new_n115_));
  anb2 g043(.dina(G33), .dinb(G32), .dout(new_n116_));
  anb1 g044(.dina(G33), .dinb(G32), .dout(new_n117_));
  anb1 g045(.dina(new_n116_), .dinb(new_n117_), .dout(new_n118_));
  anb2 g046(.dina(G31), .dinb(G30), .dout(new_n119_));
  anb1 g047(.dina(G31), .dinb(G30), .dout(new_n120_));
  anb1 g048(.dina(new_n119_), .dinb(new_n120_), .dout(new_n121_));
  anb1 g049(.dina(new_n118_), .dinb(new_n121_), .dout(new_n122_));
  anb2 g050(.dina(new_n118_), .dinb(new_n121_), .dout(new_n123_));
  anb2 g051(.dina(new_n122_), .dinb(new_n123_), .dout(new_n124_));
  anb2 g052(.dina(new_n115_), .dinb(new_n124_), .dout(new_n125_));
  anb1 g053(.dina(new_n115_), .dinb(new_n124_), .dout(new_n126_));
  anb1 g054(.dina(new_n125_), .dinb(new_n126_), .dout(G3522));
  and2 g055(.dina(G11), .dinb(G12), .dout(new_n128_));
  and1 g056(.dina(G11), .dinb(G12), .dout(new_n129_));
  anb1 g057(.dina(new_n128_), .dinb(new_n129_), .dout(new_n130_));
  anb1 g058(.dina(G13), .dinb(G14), .dout(new_n131_));
  anb2 g059(.dina(G13), .dinb(G14), .dout(new_n132_));
  anb2 g060(.dina(new_n131_), .dinb(new_n132_), .dout(new_n133_));
  anb1 g061(.dina(new_n130_), .dinb(new_n133_), .dout(new_n134_));
  anb2 g062(.dina(new_n130_), .dinb(new_n133_), .dout(new_n135_));
  anb2 g063(.dina(new_n134_), .dinb(new_n135_), .dout(new_n136_));
  nor2 g064(.dina(G7), .dinb(G8), .dout(new_n137_));
  anb2 g065(.dina(new_n73_), .dinb(new_n137_), .dout(new_n138_));
  nor1 g066(.dina(G9), .dinb(G10), .dout(new_n139_));
  nor2 g067(.dina(G9), .dinb(G10), .dout(new_n140_));
  anb2 g068(.dina(new_n139_), .dinb(new_n140_), .dout(new_n141_));
  anb2 g069(.dina(new_n138_), .dinb(new_n141_), .dout(new_n142_));
  anb1 g070(.dina(new_n138_), .dinb(new_n141_), .dout(new_n143_));
  nab2 g071(.dina(new_n142_), .dinb(new_n143_), .dout(new_n144_));
  anb1 g072(.dina(new_n136_), .dinb(new_n144_), .dout(new_n145_));
  anb2 g073(.dina(new_n136_), .dinb(new_n144_), .dout(new_n146_));
  anb2 g074(.dina(new_n145_), .dinb(new_n146_), .dout(G3523));
  nor2 g075(.dina(G1), .dinb(G2), .dout(new_n148_));
  nor2 g076(.dina(G1), .dinb(G3), .dout(new_n149_));
  anb1 g077(.dina(G4), .dinb(new_n149_), .dout(new_n150_));
  anb1 g078(.dina(new_n148_), .dinb(new_n150_), .dout(new_n151_));
  anb1 g079(.dina(G4), .dinb(G3), .dout(new_n152_));
  anb2 g080(.dina(G3), .dinb(G4), .dout(new_n153_));
  nor1 g081(.dina(G3), .dinb(G4), .dout(new_n154_));
  and2 g082(.dina(G3), .dinb(G4), .dout(new_n155_));
  anb1 g083(.dina(new_n154_), .dinb(G12), .dout(new_n156_));
  nab2 g084(.dina(G39), .dinb(new_n153_), .dout(new_n157_));
  anb2 g085(.dina(new_n156_), .dinb(new_n157_), .dout(new_n158_));
  nab1 g086(.dina(new_n151_), .dinb(new_n158_), .dout(new_n159_));
  nab2 g087(.dina(G3), .dinb(new_n95_), .dout(new_n160_));
  nab1 g088(.dina(G14), .dinb(new_n160_), .dout(new_n161_));
  and1 g089(.dina(new_n151_), .dinb(new_n160_), .dout(new_n162_));
  anb1 g090(.dina(G4), .dinb(G1), .dout(new_n163_));
  anb1 g091(.dina(new_n162_), .dinb(new_n163_), .dout(new_n164_));
  anb1 g092(.dina(G3), .dinb(new_n151_), .dout(new_n165_));
  anb1 g093(.dina(G14), .dinb(new_n165_), .dout(new_n166_));
  anb2 g094(.dina(new_n164_), .dinb(new_n166_), .dout(new_n167_));
  anb2 g095(.dina(new_n161_), .dinb(new_n167_), .dout(new_n168_));
  anb2 g096(.dina(new_n159_), .dinb(new_n168_), .dout(new_n169_));
  and1 g097(.dina(G4), .dinb(G5), .dout(new_n170_));
  nor1 g098(.dina(new_n148_), .dinb(new_n170_), .dout(new_n171_));
  anb2 g099(.dina(new_n171_), .dinb(G38), .dout(new_n172_));
  nor1 g100(.dina(G1), .dinb(G6), .dout(new_n173_));
  anb1 g101(.dina(new_n173_), .dinb(G5), .dout(new_n174_));
  nab1 g102(.dina(new_n172_), .dinb(new_n174_), .dout(new_n175_));
  anb1 g103(.dina(G37), .dinb(new_n174_), .dout(new_n176_));
  nor1 g104(.dina(G4), .dinb(G41), .dout(new_n177_));
  anb2 g105(.dina(G36), .dinb(G4), .dout(new_n178_));
  anb2 g106(.dina(new_n177_), .dinb(new_n178_), .dout(new_n179_));
  and2 g107(.dina(G4), .dinb(G49), .dout(new_n180_));
  anb1 g108(.dina(G35), .dinb(new_n180_), .dout(new_n181_));
  anb1 g109(.dina(new_n179_), .dinb(new_n181_), .dout(new_n182_));
  anb2 g110(.dina(new_n176_), .dinb(new_n182_), .dout(new_n183_));
  anb2 g111(.dina(new_n171_), .dinb(new_n183_), .dout(new_n184_));
  anb2 g112(.dina(new_n175_), .dinb(new_n184_), .dout(new_n185_));
  nor1 g113(.dina(G25), .dinb(G26), .dout(new_n186_));
  and2 g114(.dina(new_n185_), .dinb(new_n186_), .dout(new_n187_));
  anb2 g115(.dina(new_n169_), .dinb(new_n187_), .dout(new_n188_));
  and2 g116(.dina(G23), .dinb(G24), .dout(new_n189_));
  anb2 g117(.dina(new_n185_), .dinb(new_n189_), .dout(new_n190_));
  anb2 g118(.dina(new_n190_), .dinb(new_n169_), .dout(new_n191_));
  and1 g119(.dina(new_n188_), .dinb(new_n191_), .dout(new_n192_));
  anb1 g120(.dina(new_n154_), .dinb(G11), .dout(new_n193_));
  nab2 g121(.dina(G14), .dinb(new_n153_), .dout(new_n194_));
  anb2 g122(.dina(new_n193_), .dinb(new_n194_), .dout(new_n195_));
  anb2 g123(.dina(new_n151_), .dinb(new_n195_), .dout(new_n196_));
  nab2 g124(.dina(new_n160_), .dinb(new_n165_), .dout(new_n197_));
  and1 g125(.dina(G13), .dinb(new_n164_), .dout(new_n198_));
  nab1 g126(.dina(G13), .dinb(new_n197_), .dout(new_n199_));
  anb1 g127(.dina(new_n196_), .dinb(new_n198_), .dout(new_n200_));
  anb2 g128(.dina(new_n199_), .dinb(new_n200_), .dout(new_n201_));
  anb1 g129(.dina(G36), .dinb(new_n174_), .dout(new_n202_));
  nor1 g130(.dina(G4), .dinb(G40), .dout(new_n203_));
  anb2 g131(.dina(G35), .dinb(G4), .dout(new_n204_));
  anb2 g132(.dina(new_n203_), .dinb(new_n204_), .dout(new_n205_));
  anb1 g133(.dina(G34), .dinb(new_n180_), .dout(new_n206_));
  anb1 g134(.dina(new_n205_), .dinb(new_n206_), .dout(new_n207_));
  anb2 g135(.dina(new_n202_), .dinb(new_n207_), .dout(new_n208_));
  anb2 g136(.dina(new_n171_), .dinb(new_n208_), .dout(new_n209_));
  nab1 g137(.dina(new_n175_), .dinb(new_n209_), .dout(new_n210_));
  anb2 g138(.dina(new_n186_), .dinb(new_n210_), .dout(new_n211_));
  anb1 g139(.dina(new_n211_), .dinb(new_n201_), .dout(new_n212_));
  nor2 g140(.dina(new_n189_), .dinb(new_n210_), .dout(new_n213_));
  anb2 g141(.dina(new_n213_), .dinb(new_n201_), .dout(new_n214_));
  anb2 g142(.dina(new_n212_), .dinb(new_n214_), .dout(new_n215_));
  anb2 g143(.dina(new_n164_), .dinb(G11), .dout(new_n216_));
  nab1 g144(.dina(G11), .dinb(new_n160_), .dout(new_n217_));
  anb1 g145(.dina(new_n216_), .dinb(new_n217_), .dout(new_n218_));
  anb1 g146(.dina(new_n154_), .dinb(G9), .dout(new_n219_));
  anb2 g147(.dina(G12), .dinb(new_n152_), .dout(new_n220_));
  nor1 g148(.dina(G13), .dinb(new_n128_), .dout(new_n221_));
  anb1 g149(.dina(G3), .dinb(new_n221_), .dout(new_n222_));
  anb1 g150(.dina(new_n220_), .dinb(new_n222_), .dout(new_n223_));
  anb2 g151(.dina(new_n219_), .dinb(new_n223_), .dout(new_n224_));
  anb2 g152(.dina(new_n151_), .dinb(new_n224_), .dout(new_n225_));
  anb2 g153(.dina(new_n218_), .dinb(new_n225_), .dout(new_n226_));
  anb2 g154(.dina(new_n172_), .dinb(new_n173_), .dout(new_n227_));
  anb1 g155(.dina(G32), .dinb(new_n180_), .dout(new_n228_));
  nor2 g156(.dina(G4), .dinb(G33), .dout(new_n229_));
  anb1 g157(.dina(G14), .dinb(G4), .dout(new_n230_));
  anb1 g158(.dina(new_n229_), .dinb(new_n230_), .dout(new_n231_));
  anb1 g159(.dina(G34), .dinb(new_n173_), .dout(new_n232_));
  anb1 g160(.dina(new_n231_), .dinb(new_n232_), .dout(new_n233_));
  anb2 g161(.dina(new_n228_), .dinb(new_n233_), .dout(new_n234_));
  nab1 g162(.dina(new_n171_), .dinb(new_n234_), .dout(new_n235_));
  anb1 g163(.dina(new_n227_), .dinb(new_n235_), .dout(new_n236_));
  anb2 g164(.dina(new_n186_), .dinb(new_n236_), .dout(new_n237_));
  anb2 g165(.dina(new_n226_), .dinb(new_n237_), .dout(new_n238_));
  nor2 g166(.dina(new_n189_), .dinb(new_n236_), .dout(new_n239_));
  anb2 g167(.dina(new_n239_), .dinb(new_n226_), .dout(new_n240_));
  and1 g168(.dina(new_n238_), .dinb(new_n240_), .dout(new_n241_));
  anb1 g169(.dina(G12), .dinb(new_n164_), .dout(new_n242_));
  anb2 g170(.dina(G12), .dinb(new_n160_), .dout(new_n243_));
  anb2 g171(.dina(new_n242_), .dinb(new_n243_), .dout(new_n244_));
  anb1 g172(.dina(G10), .dinb(new_n155_), .dout(new_n245_));
  nab2 g173(.dina(G13), .dinb(new_n153_), .dout(new_n246_));
  nor2 g174(.dina(G12), .dinb(G13), .dout(new_n247_));
  anb2 g175(.dina(new_n76_), .dinb(new_n247_), .dout(new_n248_));
  anb1 g176(.dina(G3), .dinb(new_n248_), .dout(new_n249_));
  anb1 g177(.dina(new_n246_), .dinb(new_n249_), .dout(new_n250_));
  anb2 g178(.dina(new_n245_), .dinb(new_n250_), .dout(new_n251_));
  nab1 g179(.dina(new_n151_), .dinb(new_n251_), .dout(new_n252_));
  anb1 g180(.dina(new_n244_), .dinb(new_n252_), .dout(new_n253_));
  anb1 g181(.dina(G35), .dinb(new_n174_), .dout(new_n254_));
  nor1 g182(.dina(G4), .dinb(G39), .dout(new_n255_));
  anb2 g183(.dina(G34), .dinb(G4), .dout(new_n256_));
  anb2 g184(.dina(new_n255_), .dinb(new_n256_), .dout(new_n257_));
  anb1 g185(.dina(G33), .dinb(new_n180_), .dout(new_n258_));
  anb1 g186(.dina(new_n257_), .dinb(new_n258_), .dout(new_n259_));
  anb2 g187(.dina(new_n254_), .dinb(new_n259_), .dout(new_n260_));
  anb2 g188(.dina(new_n171_), .dinb(new_n260_), .dout(new_n261_));
  anb2 g189(.dina(new_n175_), .dinb(new_n261_), .dout(new_n262_));
  nor1 g190(.dina(new_n186_), .dinb(new_n262_), .dout(new_n263_));
  anb2 g191(.dina(new_n263_), .dinb(new_n253_), .dout(new_n264_));
  anb1 g192(.dina(new_n189_), .dinb(new_n262_), .dout(new_n265_));
  anb2 g193(.dina(new_n253_), .dinb(new_n265_), .dout(new_n266_));
  and1 g194(.dina(new_n264_), .dinb(new_n266_), .dout(new_n267_));
  nor2 g195(.dina(new_n241_), .dinb(new_n267_), .dout(new_n268_));
  and2 g196(.dina(new_n215_), .dinb(new_n268_), .dout(new_n269_));
  anb1 g197(.dina(new_n192_), .dinb(new_n269_), .dout(new_n270_));
  anb1 g198(.dina(new_n154_), .dinb(G8), .dout(new_n271_));
  anb2 g199(.dina(G11), .dinb(new_n152_), .dout(new_n272_));
  anb2 g200(.dina(new_n271_), .dinb(new_n272_), .dout(new_n273_));
  anb2 g201(.dina(new_n151_), .dinb(new_n273_), .dout(new_n274_));
  anb2 g202(.dina(G10), .dinb(new_n160_), .dout(new_n275_));
  anb1 g203(.dina(G3), .dinb(G1), .dout(new_n276_));
  anb1 g204(.dina(new_n162_), .dinb(new_n276_), .dout(new_n277_));
  anb1 g205(.dina(G10), .dinb(new_n165_), .dout(new_n278_));
  anb1 g206(.dina(new_n278_), .dinb(new_n277_), .dout(new_n279_));
  anb1 g207(.dina(new_n275_), .dinb(new_n279_), .dout(new_n280_));
  anb1 g208(.dina(new_n274_), .dinb(new_n280_), .dout(new_n281_));
  and2 g209(.dina(G5), .dinb(G6), .dout(new_n282_));
  nab1 g210(.dina(G1), .dinb(new_n282_), .dout(new_n283_));
  anb2 g211(.dina(new_n172_), .dinb(new_n283_), .dout(new_n284_));
  anb1 g212(.dina(G33), .dinb(new_n283_), .dout(new_n285_));
  nor1 g213(.dina(G4), .dinb(G13), .dout(new_n286_));
  anb2 g214(.dina(G32), .dinb(G4), .dout(new_n287_));
  anb2 g215(.dina(new_n286_), .dinb(new_n287_), .dout(new_n288_));
  anb1 g216(.dina(G31), .dinb(new_n180_), .dout(new_n289_));
  anb1 g217(.dina(new_n288_), .dinb(new_n289_), .dout(new_n290_));
  anb2 g218(.dina(new_n285_), .dinb(new_n290_), .dout(new_n291_));
  nab1 g219(.dina(new_n171_), .dinb(new_n291_), .dout(new_n292_));
  anb1 g220(.dina(new_n284_), .dinb(new_n292_), .dout(new_n293_));
  anb1 g221(.dina(new_n293_), .dinb(new_n186_), .dout(new_n294_));
  anb1 g222(.dina(new_n281_), .dinb(new_n294_), .dout(new_n295_));
  nab2 g223(.dina(new_n189_), .dinb(new_n281_), .dout(new_n296_));
  nab2 g224(.dina(new_n293_), .dinb(new_n296_), .dout(new_n297_));
  anb2 g225(.dina(new_n295_), .dinb(new_n297_), .dout(new_n298_));
  anb1 g226(.dina(G7), .dinb(new_n155_), .dout(new_n299_));
  nab2 g227(.dina(G10), .dinb(new_n153_), .dout(new_n300_));
  anb2 g228(.dina(new_n299_), .dinb(new_n300_), .dout(new_n301_));
  anb2 g229(.dina(new_n151_), .dinb(new_n301_), .dout(new_n302_));
  and1 g230(.dina(G9), .dinb(new_n277_), .dout(new_n303_));
  nab1 g231(.dina(G9), .dinb(new_n197_), .dout(new_n304_));
  anb1 g232(.dina(new_n302_), .dinb(new_n303_), .dout(new_n305_));
  anb2 g233(.dina(new_n304_), .dinb(new_n305_), .dout(new_n306_));
  anb1 g234(.dina(G32), .dinb(new_n283_), .dout(new_n307_));
  nor1 g235(.dina(G4), .dinb(G12), .dout(new_n308_));
  anb2 g236(.dina(G31), .dinb(G4), .dout(new_n309_));
  anb2 g237(.dina(new_n308_), .dinb(new_n309_), .dout(new_n310_));
  anb1 g238(.dina(G30), .dinb(new_n180_), .dout(new_n311_));
  anb1 g239(.dina(new_n310_), .dinb(new_n311_), .dout(new_n312_));
  anb2 g240(.dina(new_n307_), .dinb(new_n312_), .dout(new_n313_));
  nab1 g241(.dina(new_n171_), .dinb(new_n313_), .dout(new_n314_));
  anb1 g242(.dina(new_n284_), .dinb(new_n314_), .dout(new_n315_));
  anb2 g243(.dina(new_n186_), .dinb(new_n315_), .dout(new_n316_));
  anb2 g244(.dina(new_n306_), .dinb(new_n316_), .dout(new_n317_));
  nor2 g245(.dina(new_n189_), .dinb(new_n315_), .dout(new_n318_));
  anb1 g246(.dina(new_n306_), .dinb(new_n318_), .dout(new_n319_));
  anb1 g247(.dina(new_n317_), .dinb(new_n319_), .dout(new_n320_));
  anb2 g248(.dina(new_n277_), .dinb(G7), .dout(new_n321_));
  nab1 g249(.dina(G7), .dinb(new_n160_), .dout(new_n322_));
  anb1 g250(.dina(new_n321_), .dinb(new_n322_), .dout(new_n323_));
  anb1 g251(.dina(G21), .dinb(new_n155_), .dout(new_n324_));
  anb2 g252(.dina(G8), .dinb(new_n152_), .dout(new_n325_));
  anb1 g253(.dina(G3), .dinb(new_n74_), .dout(new_n326_));
  anb1 g254(.dina(new_n325_), .dinb(new_n326_), .dout(new_n327_));
  anb2 g255(.dina(new_n324_), .dinb(new_n327_), .dout(new_n328_));
  anb2 g256(.dina(new_n151_), .dinb(new_n328_), .dout(new_n329_));
  anb2 g257(.dina(new_n323_), .dinb(new_n329_), .dout(new_n330_));
  anb1 g258(.dina(G30), .dinb(new_n283_), .dout(new_n331_));
  nor1 g259(.dina(G4), .dinb(G10), .dout(new_n332_));
  anb2 g260(.dina(G29), .dinb(G4), .dout(new_n333_));
  anb2 g261(.dina(new_n332_), .dinb(new_n333_), .dout(new_n334_));
  anb1 g262(.dina(G28), .dinb(new_n180_), .dout(new_n335_));
  anb1 g263(.dina(new_n334_), .dinb(new_n335_), .dout(new_n336_));
  anb2 g264(.dina(new_n331_), .dinb(new_n336_), .dout(new_n337_));
  nab1 g265(.dina(new_n171_), .dinb(new_n337_), .dout(new_n338_));
  anb1 g266(.dina(new_n284_), .dinb(new_n338_), .dout(new_n339_));
  anb2 g267(.dina(new_n186_), .dinb(new_n339_), .dout(new_n340_));
  anb2 g268(.dina(new_n330_), .dinb(new_n340_), .dout(new_n341_));
  nor2 g269(.dina(new_n189_), .dinb(new_n330_), .dout(new_n342_));
  nab2 g270(.dina(new_n339_), .dinb(new_n342_), .dout(new_n343_));
  and1 g271(.dina(new_n341_), .dinb(new_n343_), .dout(new_n344_));
  anb2 g272(.dina(new_n277_), .dinb(G8), .dout(new_n345_));
  nab1 g273(.dina(G8), .dinb(new_n160_), .dout(new_n346_));
  anb1 g274(.dina(new_n345_), .dinb(new_n346_), .dout(new_n347_));
  anb1 g275(.dina(G22), .dinb(new_n155_), .dout(new_n348_));
  anb2 g276(.dina(G9), .dinb(new_n152_), .dout(new_n349_));
  and1 g277(.dina(G8), .dinb(G9), .dout(new_n350_));
  nab2 g278(.dina(new_n97_), .dinb(new_n350_), .dout(new_n351_));
  anb1 g279(.dina(G3), .dinb(new_n351_), .dout(new_n352_));
  anb1 g280(.dina(new_n349_), .dinb(new_n352_), .dout(new_n353_));
  anb2 g281(.dina(new_n348_), .dinb(new_n353_), .dout(new_n354_));
  anb2 g282(.dina(new_n151_), .dinb(new_n354_), .dout(new_n355_));
  anb2 g283(.dina(new_n347_), .dinb(new_n355_), .dout(new_n356_));
  anb1 g284(.dina(G31), .dinb(new_n283_), .dout(new_n357_));
  nor1 g285(.dina(G4), .dinb(G11), .dout(new_n358_));
  anb2 g286(.dina(G30), .dinb(G4), .dout(new_n359_));
  anb2 g287(.dina(new_n358_), .dinb(new_n359_), .dout(new_n360_));
  anb1 g288(.dina(G29), .dinb(new_n180_), .dout(new_n361_));
  anb1 g289(.dina(new_n360_), .dinb(new_n361_), .dout(new_n362_));
  anb2 g290(.dina(new_n357_), .dinb(new_n362_), .dout(new_n363_));
  nab1 g291(.dina(new_n171_), .dinb(new_n363_), .dout(new_n364_));
  anb1 g292(.dina(new_n284_), .dinb(new_n364_), .dout(new_n365_));
  anb2 g293(.dina(new_n186_), .dinb(new_n365_), .dout(new_n366_));
  anb1 g294(.dina(new_n366_), .dinb(new_n356_), .dout(new_n367_));
  nor2 g295(.dina(new_n189_), .dinb(new_n365_), .dout(new_n368_));
  anb2 g296(.dina(new_n368_), .dinb(new_n356_), .dout(new_n369_));
  anb2 g297(.dina(new_n367_), .dinb(new_n369_), .dout(new_n370_));
  nab2 g298(.dina(new_n344_), .dinb(new_n370_), .dout(new_n371_));
  anb1 g299(.dina(new_n320_), .dinb(new_n371_), .dout(new_n372_));
  anb2 g300(.dina(new_n298_), .dinb(new_n372_), .dout(new_n373_));
  anb1 g301(.dina(new_n270_), .dinb(new_n373_), .dout(G3524));
  and2 g302(.dina(new_n191_), .dinb(new_n269_), .dout(new_n375_));
  nor1 g303(.dina(new_n214_), .dinb(new_n268_), .dout(new_n376_));
  anb1 g304(.dina(new_n241_), .dinb(new_n266_), .dout(new_n377_));
  anb1 g305(.dina(new_n240_), .dinb(new_n377_), .dout(new_n378_));
  anb2 g306(.dina(new_n376_), .dinb(new_n378_), .dout(new_n379_));
  anb1 g307(.dina(new_n375_), .dinb(new_n379_), .dout(new_n380_));
  nor1 g308(.dina(new_n373_), .dinb(new_n380_), .dout(new_n381_));
  anb2 g309(.dina(new_n297_), .dinb(new_n372_), .dout(new_n382_));
  anb1 g310(.dina(new_n319_), .dinb(new_n371_), .dout(new_n383_));
  anb1 g311(.dina(new_n344_), .dinb(new_n369_), .dout(new_n384_));
  anb1 g312(.dina(new_n343_), .dinb(new_n384_), .dout(new_n385_));
  anb2 g313(.dina(new_n383_), .dinb(new_n385_), .dout(new_n386_));
  anb1 g314(.dina(new_n382_), .dinb(new_n386_), .dout(new_n387_));
  anb2 g315(.dina(new_n381_), .dinb(new_n387_), .dout(G3525));
  nab2 g316(.dina(G27), .dinb(new_n101_), .dout(new_n389_));
  nab2 g317(.dina(G48), .dinb(new_n389_), .dout(new_n390_));
  anb1 g318(.dina(new_n201_), .dinb(new_n390_), .dout(new_n391_));
  anb1 g319(.dina(new_n215_), .dinb(new_n391_), .dout(new_n392_));
  anb2 g320(.dina(new_n215_), .dinb(new_n391_), .dout(new_n393_));
  anb2 g321(.dina(new_n392_), .dinb(new_n393_), .dout(new_n394_));
  anb2 g322(.dina(new_n390_), .dinb(new_n169_), .dout(new_n395_));
  anb2 g323(.dina(new_n192_), .dinb(new_n395_), .dout(new_n396_));
  anb1 g324(.dina(new_n192_), .dinb(new_n395_), .dout(new_n397_));
  anb1 g325(.dina(new_n396_), .dinb(new_n397_), .dout(new_n398_));
  nor2 g326(.dina(G47), .dinb(new_n398_), .dout(new_n399_));
  anb1 g327(.dina(new_n394_), .dinb(new_n399_), .dout(G3526));
  anb1 g328(.dina(G5), .dinb(new_n101_), .dout(new_n401_));
  anb1 g329(.dina(new_n98_), .dinb(new_n401_), .dout(new_n402_));
  nab1 g330(.dina(new_n380_), .dinb(new_n390_), .dout(new_n403_));
  anb2 g331(.dina(G1), .dinb(new_n403_), .dout(new_n404_));
  anb2 g332(.dina(new_n402_), .dinb(new_n404_), .dout(G3527));
  anb1 g333(.dina(new_n398_), .dinb(G47), .dout(new_n406_));
  and2 g334(.dina(G2), .dinb(G3), .dout(new_n407_));
  nab2 g335(.dina(G6), .dinb(new_n407_), .dout(new_n408_));
  anb2 g336(.dina(G1), .dinb(new_n408_), .dout(new_n409_));
  nab2 g337(.dina(new_n401_), .dinb(new_n409_), .dout(new_n410_));
  anb2 g338(.dina(new_n398_), .dinb(G47), .dout(new_n411_));
  anb2 g339(.dina(new_n406_), .dinb(new_n411_), .dout(new_n412_));
  anb1 g340(.dina(new_n410_), .dinb(new_n412_), .dout(new_n413_));
  nab2 g341(.dina(G4), .dinb(new_n407_), .dout(new_n414_));
  anb1 g342(.dina(new_n398_), .dinb(new_n414_), .dout(new_n415_));
  anb2 g343(.dina(G23), .dinb(G3), .dout(new_n416_));
  anb1 g344(.dina(new_n416_), .dinb(new_n95_), .dout(new_n417_));
  nor1 g345(.dina(G4), .dinb(new_n101_), .dout(new_n418_));
  anb2 g346(.dina(new_n418_), .dinb(G14), .dout(new_n419_));
  anb2 g347(.dina(G6), .dinb(new_n144_), .dout(new_n420_));
  anb1 g348(.dina(G6), .dinb(new_n98_), .dout(new_n421_));
  nab1 g349(.dina(G3520), .dinb(new_n418_), .dout(new_n422_));
  anb2 g350(.dina(new_n421_), .dinb(new_n422_), .dout(new_n423_));
  anb1 g351(.dina(new_n420_), .dinb(new_n423_), .dout(new_n424_));
  anb1 g352(.dina(new_n419_), .dinb(new_n424_), .dout(new_n425_));
  anb1 g353(.dina(new_n417_), .dinb(new_n425_), .dout(new_n426_));
  nor2 g354(.dina(G3), .dinb(G25), .dout(new_n427_));
  and1 g355(.dina(G3), .dinb(G24), .dout(new_n428_));
  anb2 g356(.dina(new_n428_), .dinb(G26), .dout(new_n429_));
  anb1 g357(.dina(new_n427_), .dinb(new_n429_), .dout(new_n430_));
  anb1 g358(.dina(G45), .dinb(new_n430_), .dout(new_n431_));
  and2 g359(.dina(G26), .dinb(new_n428_), .dout(new_n432_));
  nor1 g360(.dina(new_n427_), .dinb(new_n432_), .dout(new_n433_));
  anb2 g361(.dina(new_n433_), .dinb(G46), .dout(new_n434_));
  anb1 g362(.dina(new_n427_), .dinb(new_n432_), .dout(new_n435_));
  anb2 g363(.dina(new_n435_), .dinb(G44), .dout(new_n436_));
  and2 g364(.dina(new_n427_), .dinb(new_n429_), .dout(new_n437_));
  and1 g365(.dina(G43), .dinb(new_n437_), .dout(new_n438_));
  nor2 g366(.dina(G3), .dinb(new_n430_), .dout(new_n439_));
  and1 g367(.dina(G41), .dinb(new_n439_), .dout(new_n440_));
  anb1 g368(.dina(G42), .dinb(new_n433_), .dout(new_n441_));
  nor2 g369(.dina(G39), .dinb(new_n437_), .dout(new_n442_));
  anb2 g370(.dina(new_n441_), .dinb(new_n442_), .dout(new_n443_));
  anb2 g371(.dina(new_n186_), .dinb(G3), .dout(new_n444_));
  anb2 g372(.dina(new_n428_), .dinb(new_n444_), .dout(new_n445_));
  nor2 g373(.dina(G40), .dinb(new_n445_), .dout(new_n446_));
  anb2 g374(.dina(new_n431_), .dinb(new_n436_), .dout(new_n447_));
  anb1 g375(.dina(new_n434_), .dinb(new_n438_), .dout(new_n448_));
  nab1 g376(.dina(new_n443_), .dinb(new_n448_), .dout(new_n449_));
  anb2 g377(.dina(new_n447_), .dinb(new_n449_), .dout(new_n450_));
  anb2 g378(.dina(new_n440_), .dinb(G4), .dout(new_n451_));
  anb1 g379(.dina(new_n446_), .dinb(new_n451_), .dout(new_n452_));
  anb2 g380(.dina(new_n450_), .dinb(new_n452_), .dout(new_n453_));
  nor1 g381(.dina(G8), .dinb(new_n435_), .dout(new_n454_));
  nab1 g382(.dina(G12), .dinb(new_n445_), .dout(new_n455_));
  nab1 g383(.dina(G13), .dinb(new_n437_), .dout(new_n456_));
  anb2 g384(.dina(new_n433_), .dinb(G22), .dout(new_n457_));
  anb2 g385(.dina(G9), .dinb(new_n437_), .dout(new_n458_));
  nab1 g386(.dina(G4), .dinb(new_n458_), .dout(new_n459_));
  nab1 g387(.dina(G11), .dinb(new_n439_), .dout(new_n460_));
  and2 g388(.dina(G10), .dinb(new_n433_), .dout(new_n461_));
  and2 g389(.dina(G7), .dinb(new_n430_), .dout(new_n462_));
  anb2 g390(.dina(new_n454_), .dinb(new_n462_), .dout(new_n463_));
  anb2 g391(.dina(new_n455_), .dinb(new_n457_), .dout(new_n464_));
  nab1 g392(.dina(new_n456_), .dinb(new_n461_), .dout(new_n465_));
  anb1 g393(.dina(new_n465_), .dinb(new_n460_), .dout(new_n466_));
  anb1 g394(.dina(new_n459_), .dinb(new_n464_), .dout(new_n467_));
  anb2 g395(.dina(new_n463_), .dinb(new_n467_), .dout(new_n468_));
  anb1 g396(.dina(new_n466_), .dinb(new_n468_), .dout(new_n469_));
  anb1 g397(.dina(new_n453_), .dinb(new_n469_), .dout(new_n470_));
  anb2 g398(.dina(new_n417_), .dinb(new_n470_), .dout(new_n471_));
  anb2 g399(.dina(new_n426_), .dinb(new_n471_), .dout(new_n472_));
  anb1 g400(.dina(new_n472_), .dinb(new_n410_), .dout(new_n473_));
  anb2 g401(.dina(new_n415_), .dinb(new_n473_), .dout(new_n474_));
  anb2 g402(.dina(new_n413_), .dinb(new_n474_), .dout(G3528));
  anb2 g403(.dina(G2), .dinb(G4), .dout(new_n476_));
  nor1 g404(.dina(new_n281_), .dinb(new_n390_), .dout(new_n477_));
  anb1 g405(.dina(new_n298_), .dinb(new_n477_), .dout(new_n478_));
  anb2 g406(.dina(new_n298_), .dinb(new_n477_), .dout(new_n479_));
  anb2 g407(.dina(new_n478_), .dinb(new_n479_), .dout(new_n480_));
  and2 g408(.dina(new_n476_), .dinb(new_n480_), .dout(new_n481_));
  anb2 g409(.dina(new_n433_), .dinb(G18), .dout(new_n482_));
  anb1 g410(.dina(G19), .dinb(new_n430_), .dout(new_n483_));
  anb1 g411(.dina(new_n482_), .dinb(new_n483_), .dout(new_n484_));
  nab1 g412(.dina(G8), .dinb(new_n445_), .dout(new_n485_));
  anb1 g413(.dina(G20), .dinb(new_n435_), .dout(new_n486_));
  nab1 g414(.dina(G7), .dinb(new_n439_), .dout(new_n487_));
  nor2 g415(.dina(G21), .dinb(new_n437_), .dout(new_n488_));
  anb2 g416(.dina(new_n486_), .dinb(new_n488_), .dout(new_n489_));
  anb1 g417(.dina(new_n484_), .dinb(new_n489_), .dout(new_n490_));
  anb1 g418(.dina(new_n457_), .dinb(new_n485_), .dout(new_n491_));
  and1 g419(.dina(new_n459_), .dinb(new_n491_), .dout(new_n492_));
  anb2 g420(.dina(new_n487_), .dinb(new_n492_), .dout(new_n493_));
  anb1 g421(.dina(new_n490_), .dinb(new_n493_), .dout(new_n494_));
  nor1 g422(.dina(G14), .dinb(new_n433_), .dout(new_n495_));
  anb2 g423(.dina(new_n430_), .dinb(G41), .dout(new_n496_));
  anb2 g424(.dina(new_n495_), .dinb(new_n496_), .dout(new_n497_));
  anb2 g425(.dina(new_n435_), .dinb(G40), .dout(new_n498_));
  nab1 g426(.dina(G11), .dinb(new_n437_), .dout(new_n499_));
  anb1 g427(.dina(new_n498_), .dinb(new_n499_), .dout(new_n500_));
  anb2 g428(.dina(new_n497_), .dinb(new_n500_), .dout(new_n501_));
  anb2 g429(.dina(G13), .dinb(new_n439_), .dout(new_n502_));
  anb1 g430(.dina(G4), .dinb(new_n455_), .dout(new_n503_));
  anb2 g431(.dina(new_n443_), .dinb(new_n503_), .dout(new_n504_));
  anb1 g432(.dina(new_n502_), .dinb(new_n504_), .dout(new_n505_));
  anb2 g433(.dina(new_n501_), .dinb(new_n505_), .dout(new_n506_));
  anb2 g434(.dina(new_n494_), .dinb(new_n506_), .dout(new_n507_));
  anb2 g435(.dina(new_n417_), .dinb(new_n507_), .dout(new_n508_));
  anb2 g436(.dina(new_n410_), .dinb(new_n508_), .dout(new_n509_));
  anb1 g437(.dina(new_n481_), .dinb(new_n509_), .dout(new_n510_));
  anb1 g438(.dina(new_n185_), .dinb(new_n210_), .dout(new_n511_));
  anb2 g439(.dina(new_n236_), .dinb(new_n262_), .dout(new_n512_));
  anb1 g440(.dina(new_n511_), .dinb(new_n512_), .dout(new_n513_));
  anb1 g441(.dina(G24), .dinb(new_n513_), .dout(new_n514_));
  anb2 g442(.dina(new_n185_), .dinb(new_n210_), .dout(new_n515_));
  anb1 g443(.dina(new_n236_), .dinb(new_n262_), .dout(new_n516_));
  anb2 g444(.dina(new_n515_), .dinb(new_n516_), .dout(new_n517_));
  anb2 g445(.dina(G24), .dinb(new_n517_), .dout(new_n518_));
  anb2 g446(.dina(new_n514_), .dinb(new_n518_), .dout(new_n519_));
  nab2 g447(.dina(new_n390_), .dinb(new_n519_), .dout(new_n520_));
  anb1 g448(.dina(new_n270_), .dinb(new_n390_), .dout(new_n521_));
  anb1 g449(.dina(new_n520_), .dinb(new_n521_), .dout(new_n522_));
  anb1 g450(.dina(G47), .dinb(new_n522_), .dout(new_n523_));
  and1 g451(.dina(new_n403_), .dinb(new_n480_), .dout(new_n524_));
  and2 g452(.dina(new_n403_), .dinb(new_n480_), .dout(new_n525_));
  anb2 g453(.dina(new_n524_), .dinb(new_n525_), .dout(new_n526_));
  nab2 g454(.dina(new_n523_), .dinb(new_n526_), .dout(new_n527_));
  nab1 g455(.dina(new_n523_), .dinb(new_n526_), .dout(new_n528_));
  anb1 g456(.dina(new_n527_), .dinb(new_n528_), .dout(new_n529_));
  nab2 g457(.dina(new_n410_), .dinb(new_n529_), .dout(new_n530_));
  anb2 g458(.dina(new_n510_), .dinb(new_n530_), .dout(G3529));
  anb2 g459(.dina(new_n390_), .dinb(new_n306_), .dout(new_n532_));
  anb2 g460(.dina(new_n320_), .dinb(new_n532_), .dout(new_n533_));
  anb1 g461(.dina(new_n320_), .dinb(new_n532_), .dout(new_n534_));
  anb1 g462(.dina(new_n533_), .dinb(new_n534_), .dout(new_n535_));
  anb1 g463(.dina(new_n356_), .dinb(new_n389_), .dout(new_n536_));
  nab2 g464(.dina(new_n370_), .dinb(new_n536_), .dout(new_n537_));
  nab1 g465(.dina(new_n370_), .dinb(new_n536_), .dout(new_n538_));
  anb1 g466(.dina(new_n537_), .dinb(new_n538_), .dout(new_n539_));
  and1 g467(.dina(new_n535_), .dinb(new_n539_), .dout(new_n540_));
  anb2 g468(.dina(new_n480_), .dinb(new_n522_), .dout(new_n541_));
  anb1 g469(.dina(new_n540_), .dinb(new_n541_), .dout(new_n542_));
  and1 g470(.dina(new_n373_), .dinb(new_n522_), .dout(new_n543_));
  anb2 g471(.dina(new_n542_), .dinb(new_n543_), .dout(new_n544_));
  anb1 g472(.dina(new_n542_), .dinb(new_n543_), .dout(new_n545_));
  anb1 g473(.dina(new_n544_), .dinb(new_n545_), .dout(new_n546_));
  anb1 g474(.dina(G47), .dinb(new_n546_), .dout(new_n547_));
  anb1 g475(.dina(new_n373_), .dinb(new_n403_), .dout(new_n548_));
  anb1 g476(.dina(new_n387_), .dinb(new_n548_), .dout(new_n549_));
  anb1 g477(.dina(new_n390_), .dinb(new_n297_), .dout(new_n550_));
  anb2 g478(.dina(new_n550_), .dinb(new_n540_), .dout(new_n551_));
  nor2 g479(.dina(new_n319_), .dinb(new_n390_), .dout(new_n552_));
  anb1 g480(.dina(new_n539_), .dinb(new_n552_), .dout(new_n553_));
  anb2 g481(.dina(new_n369_), .dinb(new_n389_), .dout(new_n554_));
  anb2 g482(.dina(new_n553_), .dinb(new_n554_), .dout(new_n555_));
  anb1 g483(.dina(new_n551_), .dinb(new_n555_), .dout(new_n556_));
  anb1 g484(.dina(new_n549_), .dinb(new_n556_), .dout(new_n557_));
  anb2 g485(.dina(new_n549_), .dinb(new_n556_), .dout(new_n558_));
  anb2 g486(.dina(new_n557_), .dinb(new_n558_), .dout(new_n559_));
  anb1 g487(.dina(new_n547_), .dinb(new_n559_), .dout(new_n560_));
  anb2 g488(.dina(new_n547_), .dinb(new_n559_), .dout(new_n561_));
  anb2 g489(.dina(new_n560_), .dinb(new_n561_), .dout(new_n562_));
  anb2 g490(.dina(new_n96_), .dinb(new_n100_), .dout(new_n563_));
  anb1 g491(.dina(new_n562_), .dinb(new_n563_), .dout(new_n564_));
  anb2 g492(.dina(G14), .dinb(new_n96_), .dout(new_n565_));
  anb2 g493(.dina(new_n565_), .dinb(new_n248_), .dout(new_n566_));
  anb2 g494(.dina(G10), .dinb(new_n351_), .dout(new_n567_));
  anb2 g495(.dina(G7), .dinb(new_n567_), .dout(new_n568_));
  nor2 g496(.dina(G7), .dinb(G9), .dout(new_n569_));
  anb2 g497(.dina(new_n100_), .dinb(new_n569_), .dout(new_n570_));
  anb1 g498(.dina(new_n568_), .dinb(new_n570_), .dout(new_n571_));
  anb1 g499(.dina(new_n566_), .dinb(new_n571_), .dout(new_n572_));
  anb2 g500(.dina(new_n564_), .dinb(new_n572_), .dout(G3530));
  anb2 g501(.dina(new_n390_), .dinb(new_n226_), .dout(new_n574_));
  nab1 g502(.dina(new_n241_), .dinb(new_n574_), .dout(new_n575_));
  nab2 g503(.dina(new_n241_), .dinb(new_n574_), .dout(new_n576_));
  anb2 g504(.dina(new_n575_), .dinb(new_n576_), .dout(new_n577_));
  and2 g505(.dina(new_n414_), .dinb(new_n577_), .dout(new_n578_));
  and2 g506(.dina(G39), .dinb(G43), .dout(new_n579_));
  anb2 g507(.dina(new_n433_), .dinb(new_n579_), .dout(new_n580_));
  nab1 g508(.dina(G13), .dinb(new_n445_), .dout(new_n581_));
  anb2 g509(.dina(new_n430_), .dinb(G42), .dout(new_n582_));
  anb2 g510(.dina(G40), .dinb(G12), .dout(new_n583_));
  and1 g511(.dina(new_n437_), .dinb(new_n583_), .dout(new_n584_));
  anb1 g512(.dina(new_n580_), .dinb(new_n584_), .dout(new_n585_));
  anb2 g513(.dina(new_n581_), .dinb(new_n582_), .dout(new_n586_));
  anb1 g514(.dina(new_n585_), .dinb(new_n586_), .dout(new_n587_));
  nab1 g515(.dina(G14), .dinb(new_n439_), .dout(new_n588_));
  anb1 g516(.dina(G41), .dinb(new_n435_), .dout(new_n589_));
  anb1 g517(.dina(G4), .dinb(new_n589_), .dout(new_n590_));
  anb2 g518(.dina(new_n588_), .dinb(new_n590_), .dout(new_n591_));
  anb1 g519(.dina(new_n587_), .dinb(new_n591_), .dout(new_n592_));
  anb1 g520(.dina(G20), .dinb(new_n430_), .dout(new_n593_));
  anb1 g521(.dina(G7), .dinb(G19), .dout(new_n594_));
  and2 g522(.dina(new_n433_), .dinb(new_n594_), .dout(new_n595_));
  anb2 g523(.dina(new_n593_), .dinb(new_n595_), .dout(new_n596_));
  anb2 g524(.dina(new_n435_), .dinb(G21), .dout(new_n597_));
  anb1 g525(.dina(G10), .dinb(G22), .dout(new_n598_));
  anb1 g526(.dina(new_n437_), .dinb(new_n598_), .dout(new_n599_));
  anb1 g527(.dina(new_n597_), .dinb(new_n599_), .dout(new_n600_));
  anb2 g528(.dina(new_n596_), .dinb(new_n600_), .dout(new_n601_));
  anb2 g529(.dina(G8), .dinb(new_n439_), .dout(new_n602_));
  nab1 g530(.dina(G9), .dinb(new_n445_), .dout(new_n603_));
  and2 g531(.dina(G4), .dinb(new_n603_), .dout(new_n604_));
  anb1 g532(.dina(new_n602_), .dinb(new_n604_), .dout(new_n605_));
  anb2 g533(.dina(new_n601_), .dinb(new_n605_), .dout(new_n606_));
  anb2 g534(.dina(new_n592_), .dinb(new_n606_), .dout(new_n607_));
  anb2 g535(.dina(new_n417_), .dinb(new_n607_), .dout(new_n608_));
  anb2 g536(.dina(new_n410_), .dinb(new_n608_), .dout(new_n609_));
  anb1 g537(.dina(new_n578_), .dinb(new_n609_), .dout(new_n610_));
  and2 g538(.dina(new_n253_), .dinb(new_n390_), .dout(new_n611_));
  anb2 g539(.dina(new_n267_), .dinb(new_n611_), .dout(new_n612_));
  anb1 g540(.dina(new_n267_), .dinb(new_n611_), .dout(new_n613_));
  anb1 g541(.dina(new_n612_), .dinb(new_n613_), .dout(new_n614_));
  anb1 g542(.dina(G3526), .dinb(new_n614_), .dout(new_n615_));
  anb1 g543(.dina(new_n390_), .dinb(new_n266_), .dout(new_n616_));
  anb1 g544(.dina(new_n390_), .dinb(new_n191_), .dout(new_n617_));
  anb1 g545(.dina(new_n394_), .dinb(new_n617_), .dout(new_n618_));
  anb2 g546(.dina(new_n214_), .dinb(new_n390_), .dout(new_n619_));
  anb2 g547(.dina(new_n618_), .dinb(new_n619_), .dout(new_n620_));
  anb2 g548(.dina(new_n614_), .dinb(new_n620_), .dout(new_n621_));
  anb2 g549(.dina(new_n616_), .dinb(new_n621_), .dout(new_n622_));
  anb1 g550(.dina(new_n577_), .dinb(new_n622_), .dout(new_n623_));
  anb2 g551(.dina(new_n577_), .dinb(new_n622_), .dout(new_n624_));
  anb2 g552(.dina(new_n623_), .dinb(new_n624_), .dout(new_n625_));
  anb2 g553(.dina(new_n615_), .dinb(new_n625_), .dout(new_n626_));
  anb1 g554(.dina(new_n615_), .dinb(new_n625_), .dout(new_n627_));
  anb1 g555(.dina(new_n626_), .dinb(new_n627_), .dout(new_n628_));
  anb2 g556(.dina(new_n394_), .dinb(new_n617_), .dout(new_n629_));
  nab1 g557(.dina(new_n618_), .dinb(new_n629_), .dout(new_n630_));
  anb1 g558(.dina(new_n411_), .dinb(new_n630_), .dout(new_n631_));
  anb2 g559(.dina(new_n411_), .dinb(new_n630_), .dout(new_n632_));
  anb2 g560(.dina(new_n631_), .dinb(new_n632_), .dout(new_n633_));
  anb2 g561(.dina(G3526), .dinb(new_n620_), .dout(new_n634_));
  nab2 g562(.dina(new_n614_), .dinb(new_n634_), .dout(new_n635_));
  nab1 g563(.dina(new_n614_), .dinb(new_n634_), .dout(new_n636_));
  anb1 g564(.dina(new_n635_), .dinb(new_n636_), .dout(new_n637_));
  anb1 g565(.dina(new_n633_), .dinb(new_n637_), .dout(new_n638_));
  anb2 g566(.dina(new_n638_), .dinb(new_n403_), .dout(new_n639_));
  anb2 g567(.dina(new_n401_), .dinb(new_n639_), .dout(new_n640_));
  anb2 g568(.dina(new_n409_), .dinb(new_n640_), .dout(new_n641_));
  anb2 g569(.dina(new_n628_), .dinb(new_n641_), .dout(new_n642_));
  anb2 g570(.dina(new_n610_), .dinb(new_n642_), .dout(G3531));
  nor1 g571(.dina(new_n394_), .dinb(new_n414_), .dout(new_n644_));
  anb1 g572(.dina(G14), .dinb(G42), .dout(new_n645_));
  nab2 g573(.dina(new_n437_), .dinb(new_n645_), .dout(new_n646_));
  anb1 g574(.dina(G43), .dinb(new_n435_), .dout(new_n647_));
  and2 g575(.dina(G41), .dinb(G45), .dout(new_n648_));
  nab1 g576(.dina(new_n433_), .dinb(new_n648_), .dout(new_n649_));
  and1 g577(.dina(G39), .dinb(new_n445_), .dout(new_n650_));
  and1 g578(.dina(G40), .dinb(new_n439_), .dout(new_n651_));
  anb2 g579(.dina(new_n430_), .dinb(G44), .dout(new_n652_));
  anb1 g580(.dina(new_n646_), .dinb(new_n649_), .dout(new_n653_));
  anb2 g581(.dina(new_n647_), .dinb(new_n652_), .dout(new_n654_));
  anb1 g582(.dina(new_n653_), .dinb(new_n654_), .dout(new_n655_));
  anb1 g583(.dina(G4), .dinb(new_n650_), .dout(new_n656_));
  anb2 g584(.dina(new_n651_), .dinb(new_n656_), .dout(new_n657_));
  anb1 g585(.dina(new_n655_), .dinb(new_n657_), .dout(new_n658_));
  nab1 g586(.dina(G10), .dinb(new_n439_), .dout(new_n659_));
  anb2 g587(.dina(G12), .dinb(new_n437_), .dout(new_n660_));
  nab1 g588(.dina(G4), .dinb(new_n660_), .dout(new_n661_));
  anb2 g589(.dina(new_n659_), .dinb(new_n661_), .dout(new_n662_));
  anb2 g590(.dina(G11), .dinb(new_n445_), .dout(new_n663_));
  nab1 g591(.dina(G8), .dinb(new_n437_), .dout(new_n664_));
  anb1 g592(.dina(new_n663_), .dinb(new_n664_), .dout(new_n665_));
  nor1 g593(.dina(G7), .dinb(new_n435_), .dout(new_n666_));
  anb2 g594(.dina(new_n430_), .dinb(G22), .dout(new_n667_));
  anb2 g595(.dina(new_n666_), .dinb(new_n667_), .dout(new_n668_));
  anb2 g596(.dina(G21), .dinb(G9), .dout(new_n669_));
  anb2 g597(.dina(new_n433_), .dinb(new_n669_), .dout(new_n670_));
  anb2 g598(.dina(new_n668_), .dinb(new_n670_), .dout(new_n671_));
  anb1 g599(.dina(new_n665_), .dinb(new_n671_), .dout(new_n672_));
  anb2 g600(.dina(new_n662_), .dinb(new_n672_), .dout(new_n673_));
  anb2 g601(.dina(new_n658_), .dinb(new_n673_), .dout(new_n674_));
  anb2 g602(.dina(new_n417_), .dinb(new_n674_), .dout(new_n675_));
  anb1 g603(.dina(new_n675_), .dinb(new_n410_), .dout(new_n676_));
  anb2 g604(.dina(new_n644_), .dinb(new_n676_), .dout(new_n677_));
  nab2 g605(.dina(new_n403_), .dinb(new_n633_), .dout(new_n678_));
  and1 g606(.dina(new_n409_), .dinb(new_n633_), .dout(new_n679_));
  nab1 g607(.dina(new_n403_), .dinb(new_n633_), .dout(new_n680_));
  anb1 g608(.dina(new_n678_), .dinb(new_n680_), .dout(new_n681_));
  anb1 g609(.dina(new_n681_), .dinb(new_n401_), .dout(new_n682_));
  anb1 g610(.dina(new_n677_), .dinb(new_n679_), .dout(new_n683_));
  anb2 g611(.dina(new_n682_), .dinb(new_n683_), .dout(G3532));
  anb1 g612(.dina(new_n637_), .dinb(new_n680_), .dout(new_n685_));
  anb2 g613(.dina(new_n637_), .dinb(new_n680_), .dout(new_n686_));
  anb2 g614(.dina(new_n685_), .dinb(new_n686_), .dout(new_n687_));
  nab1 g615(.dina(new_n401_), .dinb(new_n687_), .dout(new_n688_));
  nab2 g616(.dina(new_n409_), .dinb(new_n637_), .dout(new_n689_));
  anb2 g617(.dina(new_n414_), .dinb(new_n614_), .dout(new_n690_));
  and2 g618(.dina(G40), .dinb(G44), .dout(new_n691_));
  anb2 g619(.dina(new_n433_), .dinb(new_n691_), .dout(new_n692_));
  anb2 g620(.dina(G41), .dinb(G13), .dout(new_n693_));
  nab1 g621(.dina(G14), .dinb(new_n445_), .dout(new_n694_));
  anb1 g622(.dina(G42), .dinb(new_n435_), .dout(new_n695_));
  and1 g623(.dina(G39), .dinb(new_n439_), .dout(new_n696_));
  anb2 g624(.dina(new_n430_), .dinb(G43), .dout(new_n697_));
  nor2 g625(.dina(G41), .dinb(new_n437_), .dout(new_n698_));
  anb2 g626(.dina(new_n695_), .dinb(new_n698_), .dout(new_n699_));
  anb1 g627(.dina(new_n692_), .dinb(new_n699_), .dout(new_n700_));
  anb1 g628(.dina(G4), .dinb(new_n456_), .dout(new_n701_));
  anb2 g629(.dina(new_n694_), .dinb(new_n697_), .dout(new_n702_));
  anb1 g630(.dina(new_n701_), .dinb(new_n702_), .dout(new_n703_));
  anb2 g631(.dina(new_n696_), .dinb(new_n703_), .dout(new_n704_));
  anb1 g632(.dina(new_n700_), .dinb(new_n704_), .dout(new_n705_));
  anb1 g633(.dina(G22), .dinb(new_n435_), .dout(new_n706_));
  and1 g634(.dina(G7), .dinb(G11), .dout(new_n707_));
  nab2 g635(.dina(new_n437_), .dinb(new_n707_), .dout(new_n708_));
  anb2 g636(.dina(new_n430_), .dinb(G21), .dout(new_n709_));
  nab1 g637(.dina(G10), .dinb(new_n445_), .dout(new_n710_));
  anb2 g638(.dina(G9), .dinb(new_n439_), .dout(new_n711_));
  anb2 g639(.dina(G20), .dinb(G8), .dout(new_n712_));
  anb2 g640(.dina(new_n433_), .dinb(new_n712_), .dout(new_n713_));
  anb2 g641(.dina(new_n710_), .dinb(new_n713_), .dout(new_n714_));
  anb2 g642(.dina(new_n706_), .dinb(new_n709_), .dout(new_n715_));
  nab1 g643(.dina(G4), .dinb(new_n711_), .dout(new_n716_));
  anb2 g644(.dina(new_n715_), .dinb(new_n716_), .dout(new_n717_));
  anb1 g645(.dina(new_n708_), .dinb(new_n714_), .dout(new_n718_));
  anb2 g646(.dina(new_n717_), .dinb(new_n718_), .dout(new_n719_));
  anb2 g647(.dina(new_n705_), .dinb(new_n719_), .dout(new_n720_));
  anb2 g648(.dina(new_n417_), .dinb(new_n720_), .dout(new_n721_));
  anb2 g649(.dina(new_n410_), .dinb(new_n721_), .dout(new_n722_));
  anb1 g650(.dina(new_n690_), .dinb(new_n722_), .dout(new_n723_));
  anb1 g651(.dina(new_n689_), .dinb(new_n723_), .dout(new_n724_));
  anb2 g652(.dina(new_n688_), .dinb(new_n724_), .dout(G3533));
  nab2 g653(.dina(G47), .dinb(new_n541_), .dout(new_n726_));
  anb1 g654(.dina(new_n535_), .dinb(new_n726_), .dout(new_n727_));
  anb1 g655(.dina(new_n535_), .dinb(new_n550_), .dout(new_n728_));
  nab2 g656(.dina(new_n552_), .dinb(new_n728_), .dout(new_n729_));
  anb1 g657(.dina(new_n539_), .dinb(new_n729_), .dout(new_n730_));
  anb2 g658(.dina(new_n539_), .dinb(new_n729_), .dout(new_n731_));
  anb2 g659(.dina(new_n730_), .dinb(new_n731_), .dout(new_n732_));
  anb1 g660(.dina(new_n727_), .dinb(new_n732_), .dout(new_n733_));
  anb2 g661(.dina(new_n727_), .dinb(new_n732_), .dout(new_n734_));
  nab1 g662(.dina(new_n733_), .dinb(new_n734_), .dout(new_n735_));
  nab2 g663(.dina(new_n525_), .dinb(new_n550_), .dout(new_n736_));
  anb2 g664(.dina(new_n535_), .dinb(new_n726_), .dout(new_n737_));
  anb2 g665(.dina(new_n727_), .dinb(new_n737_), .dout(new_n738_));
  anb2 g666(.dina(new_n736_), .dinb(new_n738_), .dout(new_n739_));
  anb1 g667(.dina(new_n736_), .dinb(new_n738_), .dout(new_n740_));
  anb1 g668(.dina(new_n739_), .dinb(new_n740_), .dout(new_n741_));
  and1 g669(.dina(G47), .dinb(new_n543_), .dout(new_n742_));
  anb2 g670(.dina(new_n549_), .dinb(new_n742_), .dout(new_n743_));
  nab1 g671(.dina(new_n741_), .dinb(new_n743_), .dout(new_n744_));
  anb1 g672(.dina(new_n735_), .dinb(new_n744_), .dout(new_n745_));
  anb2 g673(.dina(new_n735_), .dinb(new_n744_), .dout(new_n746_));
  anb2 g674(.dina(new_n745_), .dinb(new_n746_), .dout(new_n747_));
  nab1 g675(.dina(new_n401_), .dinb(new_n747_), .dout(new_n748_));
  nab1 g676(.dina(new_n476_), .dinb(new_n539_), .dout(new_n749_));
  nor1 g677(.dina(G14), .dinb(new_n435_), .dout(new_n750_));
  anb2 g678(.dina(new_n430_), .dinb(G39), .dout(new_n751_));
  anb2 g679(.dina(new_n433_), .dinb(new_n583_), .dout(new_n752_));
  anb2 g680(.dina(new_n750_), .dinb(new_n751_), .dout(new_n753_));
  anb1 g681(.dina(new_n752_), .dinb(new_n753_), .dout(new_n754_));
  nab2 g682(.dina(new_n458_), .dinb(new_n710_), .dout(new_n755_));
  anb1 g683(.dina(new_n701_), .dinb(new_n755_), .dout(new_n756_));
  anb2 g684(.dina(new_n460_), .dinb(new_n756_), .dout(new_n757_));
  anb1 g685(.dina(new_n754_), .dinb(new_n757_), .dout(new_n758_));
  anb1 g686(.dina(G18), .dinb(new_n435_), .dout(new_n759_));
  and2 g687(.dina(G16), .dinb(G20), .dout(new_n760_));
  anb2 g688(.dina(new_n433_), .dinb(new_n760_), .dout(new_n761_));
  nor2 g689(.dina(G22), .dinb(new_n445_), .dout(new_n762_));
  anb1 g690(.dina(new_n437_), .dinb(new_n594_), .dout(new_n763_));
  anb1 g691(.dina(new_n761_), .dinb(new_n763_), .dout(new_n764_));
  and1 g692(.dina(G21), .dinb(new_n439_), .dout(new_n765_));
  anb2 g693(.dina(new_n430_), .dinb(G17), .dout(new_n766_));
  anb2 g694(.dina(new_n765_), .dinb(new_n766_), .dout(new_n767_));
  nab1 g695(.dina(G4), .dinb(new_n762_), .dout(new_n768_));
  anb2 g696(.dina(new_n759_), .dinb(new_n764_), .dout(new_n769_));
  anb1 g697(.dina(new_n768_), .dinb(new_n769_), .dout(new_n770_));
  anb2 g698(.dina(new_n767_), .dinb(new_n770_), .dout(new_n771_));
  anb2 g699(.dina(new_n758_), .dinb(new_n771_), .dout(new_n772_));
  anb2 g700(.dina(new_n417_), .dinb(new_n772_), .dout(new_n773_));
  anb1 g701(.dina(new_n773_), .dinb(new_n410_), .dout(new_n774_));
  anb2 g702(.dina(new_n749_), .dinb(new_n774_), .dout(new_n775_));
  anb1 g703(.dina(new_n409_), .dinb(new_n735_), .dout(new_n776_));
  anb1 g704(.dina(new_n775_), .dinb(new_n776_), .dout(new_n777_));
  anb1 g705(.dina(new_n777_), .dinb(new_n748_), .dout(new_n778_));
  anb2 g706(.dina(new_n748_), .dinb(new_n777_), .dout(G3534));
  anb2 g707(.dina(new_n389_), .dinb(new_n330_), .dout(new_n780_));
  nab1 g708(.dina(new_n344_), .dinb(new_n780_), .dout(new_n781_));
  nab2 g709(.dina(new_n344_), .dinb(new_n780_), .dout(new_n782_));
  anb2 g710(.dina(new_n781_), .dinb(new_n782_), .dout(new_n783_));
  and2 g711(.dina(new_n476_), .dinb(new_n783_), .dout(new_n784_));
  nor1 g712(.dina(G5), .dinb(G7), .dout(new_n785_));
  anb1 g713(.dina(G17), .dinb(new_n435_), .dout(new_n786_));
  nor1 g714(.dina(G18), .dinb(G22), .dout(new_n787_));
  anb1 g715(.dina(new_n437_), .dinb(new_n787_), .dout(new_n788_));
  and2 g716(.dina(G15), .dinb(G19), .dout(new_n789_));
  anb2 g717(.dina(new_n433_), .dinb(new_n789_), .dout(new_n790_));
  nor2 g718(.dina(G21), .dinb(new_n445_), .dout(new_n791_));
  and1 g719(.dina(G20), .dinb(new_n439_), .dout(new_n792_));
  anb1 g720(.dina(G16), .dinb(new_n430_), .dout(new_n793_));
  anb2 g721(.dina(new_n788_), .dinb(new_n790_), .dout(new_n794_));
  anb1 g722(.dina(new_n791_), .dinb(new_n793_), .dout(new_n795_));
  anb2 g723(.dina(new_n794_), .dinb(new_n795_), .dout(new_n796_));
  anb1 g724(.dina(new_n170_), .dinb(new_n786_), .dout(new_n797_));
  anb1 g725(.dina(new_n797_), .dinb(new_n792_), .dout(new_n798_));
  anb2 g726(.dina(new_n796_), .dinb(new_n798_), .dout(new_n799_));
  anb2 g727(.dina(new_n785_), .dinb(new_n799_), .dout(new_n800_));
  anb1 g728(.dina(G5), .dinb(new_n603_), .dout(new_n801_));
  nor1 g729(.dina(G13), .dinb(new_n435_), .dout(new_n802_));
  anb2 g730(.dina(G39), .dinb(G11), .dout(new_n803_));
  anb2 g731(.dina(new_n433_), .dinb(new_n803_), .dout(new_n804_));
  and2 g732(.dina(G14), .dinb(new_n430_), .dout(new_n805_));
  anb2 g733(.dina(new_n802_), .dinb(new_n805_), .dout(new_n806_));
  anb2 g734(.dina(new_n664_), .dinb(new_n804_), .dout(new_n807_));
  and2 g735(.dina(new_n806_), .dinb(new_n807_), .dout(new_n808_));
  anb1 g736(.dina(new_n801_), .dinb(new_n808_), .dout(new_n809_));
  anb2 g737(.dina(new_n662_), .dinb(new_n809_), .dout(new_n810_));
  anb2 g738(.dina(new_n800_), .dinb(new_n810_), .dout(new_n811_));
  anb2 g739(.dina(new_n417_), .dinb(new_n811_), .dout(new_n812_));
  anb2 g740(.dina(new_n410_), .dinb(new_n812_), .dout(new_n813_));
  anb1 g741(.dina(new_n784_), .dinb(new_n813_), .dout(new_n814_));
  nab1 g742(.dina(new_n556_), .dinb(new_n783_), .dout(new_n815_));
  nab2 g743(.dina(new_n556_), .dinb(new_n783_), .dout(new_n816_));
  anb2 g744(.dina(new_n815_), .dinb(new_n816_), .dout(new_n817_));
  anb2 g745(.dina(new_n733_), .dinb(new_n817_), .dout(new_n818_));
  anb1 g746(.dina(new_n733_), .dinb(new_n817_), .dout(new_n819_));
  anb1 g747(.dina(new_n818_), .dinb(new_n819_), .dout(new_n820_));
  and2 g748(.dina(new_n735_), .dinb(new_n741_), .dout(new_n821_));
  anb2 g749(.dina(new_n743_), .dinb(new_n821_), .dout(new_n822_));
  anb2 g750(.dina(new_n401_), .dinb(new_n822_), .dout(new_n823_));
  anb2 g751(.dina(new_n409_), .dinb(new_n823_), .dout(new_n824_));
  anb2 g752(.dina(new_n820_), .dinb(new_n824_), .dout(new_n825_));
  anb2 g753(.dina(new_n814_), .dinb(new_n825_), .dout(G3535));
  anb2 g754(.dina(new_n476_), .dinb(new_n535_), .dout(new_n827_));
  anb2 g755(.dina(new_n435_), .dinb(G19), .dout(new_n828_));
  nab1 g756(.dina(G7), .dinb(new_n445_), .dout(new_n829_));
  nor2 g757(.dina(new_n437_), .dinb(new_n712_), .dout(new_n830_));
  anb1 g758(.dina(G18), .dinb(new_n430_), .dout(new_n831_));
  anb1 g759(.dina(new_n828_), .dinb(new_n831_), .dout(new_n832_));
  anb2 g760(.dina(new_n829_), .dinb(new_n830_), .dout(new_n833_));
  anb1 g761(.dina(new_n832_), .dinb(new_n833_), .dout(new_n834_));
  and1 g762(.dina(G22), .dinb(new_n439_), .dout(new_n835_));
  and2 g763(.dina(G17), .dinb(G21), .dout(new_n836_));
  anb2 g764(.dina(new_n433_), .dinb(new_n836_), .dout(new_n837_));
  nab1 g765(.dina(G4), .dinb(new_n837_), .dout(new_n838_));
  anb2 g766(.dina(new_n835_), .dinb(new_n838_), .dout(new_n839_));
  anb1 g767(.dina(new_n834_), .dinb(new_n839_), .dout(new_n840_));
  and1 g768(.dina(G10), .dinb(G14), .dout(new_n841_));
  anb1 g769(.dina(new_n437_), .dinb(new_n841_), .dout(new_n842_));
  anb2 g770(.dina(new_n430_), .dinb(G40), .dout(new_n843_));
  anb2 g771(.dina(new_n433_), .dinb(new_n693_), .dout(new_n844_));
  anb1 g772(.dina(G39), .dinb(new_n435_), .dout(new_n845_));
  anb2 g773(.dina(new_n842_), .dinb(new_n844_), .dout(new_n846_));
  nab1 g774(.dina(G12), .dinb(new_n439_), .dout(new_n847_));
  anb1 g775(.dina(new_n663_), .dinb(new_n846_), .dout(new_n848_));
  anb2 g776(.dina(new_n845_), .dinb(G4), .dout(new_n849_));
  anb1 g777(.dina(new_n843_), .dinb(new_n847_), .dout(new_n850_));
  anb2 g778(.dina(new_n849_), .dinb(new_n850_), .dout(new_n851_));
  anb1 g779(.dina(new_n848_), .dinb(new_n851_), .dout(new_n852_));
  and2 g780(.dina(new_n840_), .dinb(new_n852_), .dout(new_n853_));
  anb2 g781(.dina(new_n417_), .dinb(new_n853_), .dout(new_n854_));
  anb2 g782(.dina(new_n410_), .dinb(new_n854_), .dout(new_n855_));
  anb1 g783(.dina(new_n827_), .dinb(new_n855_), .dout(new_n856_));
  anb1 g784(.dina(new_n741_), .dinb(new_n743_), .dout(new_n857_));
  anb1 g785(.dina(new_n409_), .dinb(new_n741_), .dout(new_n858_));
  and2 g786(.dina(new_n401_), .dinb(new_n744_), .dout(new_n859_));
  anb2 g787(.dina(new_n858_), .dinb(new_n859_), .dout(new_n860_));
  anb2 g788(.dina(new_n857_), .dinb(new_n860_), .dout(new_n861_));
  anb2 g789(.dina(new_n856_), .dinb(new_n861_), .dout(G3536));
  anb1 g790(.dina(new_n778_), .dinb(G3535), .dout(new_n863_));
  and2 g791(.dina(G3529), .dinb(G3536), .dout(new_n864_));
  nor1 g792(.dina(G3531), .dinb(G3533), .dout(new_n865_));
  and2 g793(.dina(G3528), .dinb(G3532), .dout(new_n866_));
  anb1 g794(.dina(new_n865_), .dinb(new_n866_), .dout(new_n867_));
  anb2 g795(.dina(new_n864_), .dinb(new_n867_), .dout(new_n868_));
  nab2 g796(.dina(new_n863_), .dinb(new_n868_), .dout(G3537));
  nor2 g797(.dina(G27), .dinb(G48), .dout(new_n870_));
  anb1 g798(.dina(new_n863_), .dinb(new_n870_), .dout(new_n871_));
  and1 g799(.dina(G27), .dinb(G3537), .dout(new_n872_));
  anb2 g800(.dina(new_n871_), .dinb(new_n872_), .dout(G3538));
  and1 g801(.dina(G3528), .dinb(G3532), .dout(new_n874_));
  nab2 g802(.dina(new_n866_), .dinb(new_n874_), .dout(new_n875_));
  nor2 g803(.dina(G3531), .dinb(G3533), .dout(new_n876_));
  anb2 g804(.dina(new_n865_), .dinb(new_n876_), .dout(new_n877_));
  anb2 g805(.dina(new_n875_), .dinb(new_n877_), .dout(new_n878_));
  anb1 g806(.dina(new_n875_), .dinb(new_n877_), .dout(new_n879_));
  anb1 g807(.dina(new_n878_), .dinb(new_n879_), .dout(new_n880_));
  and1 g808(.dina(G3529), .dinb(G3536), .dout(new_n881_));
  nab2 g809(.dina(new_n864_), .dinb(new_n881_), .dout(new_n882_));
  anb2 g810(.dina(new_n778_), .dinb(G3535), .dout(new_n883_));
  anb2 g811(.dina(new_n863_), .dinb(new_n883_), .dout(new_n884_));
  anb1 g812(.dina(G50), .dinb(new_n884_), .dout(new_n885_));
  nab1 g813(.dina(G50), .dinb(new_n884_), .dout(new_n886_));
  anb1 g814(.dina(new_n870_), .dinb(new_n885_), .dout(new_n887_));
  anb2 g815(.dina(new_n886_), .dinb(new_n887_), .dout(new_n888_));
  anb2 g816(.dina(new_n882_), .dinb(new_n888_), .dout(new_n889_));
  anb1 g817(.dina(new_n882_), .dinb(new_n888_), .dout(new_n890_));
  anb1 g818(.dina(new_n889_), .dinb(new_n890_), .dout(new_n891_));
  anb2 g819(.dina(new_n880_), .dinb(new_n891_), .dout(new_n892_));
  anb1 g820(.dina(new_n880_), .dinb(new_n891_), .dout(new_n893_));
  nab2 g821(.dina(new_n892_), .dinb(new_n893_), .dout(G3539));
  anb2 g822(.dina(new_n882_), .dinb(new_n884_), .dout(new_n895_));
  anb1 g823(.dina(new_n882_), .dinb(new_n884_), .dout(new_n896_));
  anb1 g824(.dina(new_n895_), .dinb(new_n896_), .dout(new_n897_));
  anb2 g825(.dina(new_n880_), .dinb(new_n897_), .dout(new_n898_));
  anb1 g826(.dina(new_n880_), .dinb(new_n897_), .dout(new_n899_));
  anb1 g827(.dina(new_n898_), .dinb(new_n899_), .dout(G3540));
endmodule


