
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  G42,
  G43,
  G44,
  G45,
  G46,
  G47,
  G48,
  G49,
  G50,
  G51,
  G52,
  G53,
  G54,
  G55,
  G56,
  G57,
  G58,
  G59,
  G60,
  G61,
  G62,
  G63,
  G64,
  G65,
  G66,
  G67,
  G68,
  G69,
  G70,
  G71,
  G72,
  G73,
  G74,
  G75,
  G76,
  G77,
  G78,
  G79,
  G80,
  G81,
  G82,
  G83,
  G84,
  G85,
  G86,
  G87,
  G88,
  G89,
  G90,
  G91,
  G92,
  G93,
  G94,
  G95,
  G96,
  G97,
  G98,
  G99,
  G100,
  G101,
  G102,
  G103,
  G104,
  G105,
  G106,
  G107,
  G108,
  G109,
  G110,
  G111,
  G112,
  G113,
  G114,
  G115,
  G116,
  G117,
  G118,
  G119,
  G120,
  G121,
  G122,
  G123,
  G124,
  G125,
  G126,
  G127,
  G128,
  G129,
  G130,
  G131,
  G132,
  G133,
  G134,
  G135,
  G136,
  G137,
  G138,
  G139,
  G140,
  G141,
  G142,
  G143,
  G144,
  G145,
  G146,
  G147,
  G148,
  G149,
  G150,
  G151,
  G152,
  G153,
  G154,
  G155,
  G156,
  G157,
  n1416_lo,
  n1419_lo,
  n1422_lo,
  n1425_lo,
  n1428_lo,
  n1431_lo,
  n1434_lo,
  n1437_lo,
  n1440_lo,
  n1443_lo,
  n1446_lo,
  n1449_lo,
  n1452_lo,
  n1455_lo,
  n1458_lo,
  n1464_lo,
  n1467_lo,
  n1470_lo,
  n1476_lo,
  n1479_lo,
  n1482_lo,
  n1488_lo,
  n1491_lo,
  n1494_lo,
  n1497_lo,
  n1500_lo,
  n1503_lo,
  n1512_lo,
  n1515_lo,
  n1518_lo,
  n1521_lo,
  n1524_lo,
  n1527_lo,
  n1530_lo,
  n1533_lo,
  n1536_lo,
  n1539_lo,
  n1542_lo,
  n1545_lo,
  n1548_lo,
  n1551_lo,
  n1554_lo,
  n1560_lo,
  n1563_lo,
  n1566_lo,
  n1572_lo,
  n1575_lo,
  n1578_lo,
  n1584_lo,
  n1587_lo,
  n1590_lo,
  n1596_lo,
  n1599_lo,
  n1602_lo,
  n1608_lo,
  n1611_lo,
  n1614_lo,
  n1620_lo,
  n1623_lo,
  n1626_lo,
  n1632_lo,
  n1635_lo,
  n1638_lo,
  n1644_lo,
  n1647_lo,
  n1650_lo,
  n1656_lo,
  n1659_lo,
  n1662_lo,
  n1668_lo,
  n1671_lo,
  n1674_lo,
  n1680_lo,
  n1683_lo,
  n1686_lo,
  n1692_lo,
  n1695_lo,
  n1698_lo,
  n1704_lo,
  n1707_lo,
  n1710_lo,
  n1716_lo,
  n1719_lo,
  n1722_lo,
  n1728_lo,
  n1731_lo,
  n1734_lo,
  n1740_lo,
  n1743_lo,
  n1746_lo,
  n1749_lo,
  n1752_lo,
  n1755_lo,
  n1758_lo,
  n1761_lo,
  n1764_lo,
  n1776_lo,
  n1788_lo,
  n1791_lo,
  n1794_lo,
  n1797_lo,
  n1800_lo,
  n1803_lo,
  n1812_lo,
  n1815_lo,
  n1824_lo,
  n1827_lo,
  n1836_lo,
  n1839_lo,
  n1848_lo,
  n1851_lo,
  n1860_lo,
  n1872_lo,
  n1875_lo,
  n1884_lo,
  n1896_lo,
  n1899_lo,
  n1908_lo,
  n1920_lo,
  n1923_lo,
  n1926_lo,
  n1929_lo,
  n1932_lo,
  n1935_lo,
  n1944_lo,
  n1947_lo,
  n1956_lo,
  n1959_lo,
  n1962_lo,
  n1968_lo,
  n1971_lo,
  n1980_lo,
  n1983_lo,
  n1992_lo,
  n1995_lo,
  n2004_lo,
  n2016_lo,
  n2019_lo,
  n2028_lo,
  n2040_lo,
  n2043_lo,
  n2046_lo,
  n2049_lo,
  n2052_lo,
  n2055_lo,
  n2064_lo,
  n2067_lo,
  n2076_lo,
  n2079_lo,
  n2088_lo,
  n2091_lo,
  n2100_lo,
  n2103_lo,
  n2112_lo,
  n2115_lo,
  n2124_lo,
  n2127_lo,
  n2136_lo,
  n2148_lo,
  n2151_lo,
  n2160_lo,
  n2172_lo,
  n2175_lo,
  n2178_lo,
  n2181_lo,
  n2184_lo,
  n2187_lo,
  n2196_lo,
  n2199_lo,
  n2208_lo,
  n2211_lo,
  n2220_lo,
  n2223_lo,
  n2232_lo,
  n2235_lo,
  n2244_lo,
  n2247_lo,
  n2256_lo,
  n2259_lo,
  n2268_lo,
  n2280_lo,
  n2283_lo,
  n2292_lo,
  n2295_lo,
  n2298_lo,
  n2301_lo,
  n2304_lo,
  n2307_lo,
  n2316_lo,
  n2319_lo,
  n2322_lo,
  n2325_lo,
  n2328_lo,
  n2331_lo,
  n2340_lo,
  n2343_lo,
  n2376_lo,
  n2379_lo,
  n2388_lo,
  n2391_lo,
  n2400_lo,
  n2403_lo,
  n2412_lo,
  n2415_lo,
  n2424_lo,
  n2427_lo,
  n2436_lo,
  n2439_lo,
  n2442_lo,
  n2445_lo,
  n2448_lo,
  n2451_lo,
  n2460_lo,
  n2463_lo,
  n2496_lo,
  n2499_lo,
  n2508_lo,
  n2511_lo,
  n2520_lo,
  n2523_lo,
  n2532_lo,
  n2535_lo,
  n2544_lo,
  n2547_lo,
  n2556_lo,
  n2559_lo,
  n2562_lo,
  n2565_lo,
  n2568_lo,
  n2571_lo,
  n2580_lo,
  n2583_lo,
  n2616_lo,
  n2619_lo,
  n2628_lo,
  n2631_lo,
  n2640_lo,
  n2643_lo,
  n2652_lo,
  n2655_lo,
  n2664_lo,
  n2667_lo,
  n2676_lo,
  n2679_lo,
  n2682_lo,
  n2685_lo,
  n2688_lo,
  n2691_lo,
  n2700_lo,
  n2703_lo,
  n2736_lo,
  n2739_lo,
  n2748_lo,
  n2751_lo,
  n2760_lo,
  n2763_lo,
  n2772_lo,
  n2775_lo,
  n2784_lo,
  n2787_lo,
  n2790_lo,
  n2793_lo,
  n2796_lo,
  n2799_lo,
  n2802_lo,
  n2805_lo,
  n2808_lo,
  n2820_lo,
  n2823_lo,
  n2826_lo,
  n2829_lo,
  n2832_lo,
  n2835_lo,
  n2838_lo,
  n2841_lo,
  n2844_lo,
  n2856_lo,
  n2859_lo,
  n2862_lo,
  n2865_lo,
  n2868_lo,
  n2871_lo,
  n2874_lo,
  n2877_lo,
  n2880_lo,
  n2883_lo,
  n2886_lo,
  n2889_lo,
  n2892_lo,
  n2895_lo,
  n2898_lo,
  n2901_lo,
  n2904_lo,
  n2907_lo,
  n2916_lo,
  n2919_lo,
  n2925_lo,
  n2928_lo,
  n2940_lo,
  n2943_lo,
  n2952_lo,
  n2955_lo,
  n2961_lo,
  n2964_lo,
  n2967_lo,
  n2970_lo,
  n2976_lo,
  n2979_lo,
  n2982_lo,
  n2988_lo,
  n2991_lo,
  n2994_lo,
  n2997_lo,
  n3000_lo,
  n3003_lo,
  n3006_lo,
  n3012_lo,
  n3015_lo,
  n3018_lo,
  n3021_lo,
  n3024_lo,
  n3027_lo,
  n3030_lo,
  n3033_lo,
  n3036_lo,
  n3039_lo,
  n3045_lo,
  n3048_lo,
  n3051_lo,
  n3054_lo,
  n3057_lo,
  n3060_lo,
  n3063_lo,
  n3069_lo,
  n3072_lo,
  n3075_lo,
  n3081_lo,
  n3084_lo,
  n3087_lo,
  n3093_lo,
  n3096_lo,
  n3099_lo,
  n3102_lo,
  n3105_lo,
  n3108_lo,
  n3111_lo,
  n3114_lo,
  n3117_lo,
  n3120_lo,
  n3123_lo,
  n3126_lo,
  n3129_lo,
  n3132_lo,
  n3135_lo,
  n3138_lo,
  n3141_lo,
  n3156_lo,
  n3168_lo,
  n3171_lo,
  n3174_lo,
  n3177_lo,
  n3180_lo,
  n3183_lo,
  n3192_lo,
  n3195_lo,
  n3204_lo,
  n3207_lo,
  n3210_lo,
  n3216_lo,
  n3219_lo,
  n3222_lo,
  n3228_lo,
  n3231_lo,
  n3240_lo,
  n3243_lo,
  n3252_lo,
  n3255_lo,
  n3258_lo,
  n3264_lo,
  n3267_lo,
  n3270_lo,
  n3276_lo,
  n3279_lo,
  n3282_lo,
  n3288_lo,
  n3291_lo,
  n3294_lo,
  n3603_o2,
  n3604_o2,
  n1391_inv,
  n3798_o2,
  n3846_o2,
  n4019_o2,
  n4017_o2,
  n2177_o2,
  n2150_o2,
  n2154_o2,
  n2184_o2,
  n2515_o2,
  n3837_o2,
  n2167_o2,
  n2118_o2,
  n2186_o2,
  n2174_o2,
  n3964_o2,
  n4005_o2,
  n4006_o2,
  n1445_inv,
  n2176_o2,
  n2227_o2,
  n2236_o2,
  n2245_o2,
  n2518_o2,
  n4023_o2,
  n1466_inv,
  n4038_o2,
  n4039_o2,
  n1475_inv,
  n2119_o2,
  n2275_o2,
  n2595_o2,
  n2594_o2,
  lo498_buf_o2,
  lo502_buf_o2,
  lo550_buf_o2,
  n2596_o2,
  n2593_o2,
  n2668_o2,
  lo542_buf_o2,
  n2667_o2,
  n2404_o2,
  n2410_o2,
  n2419_o2,
  n2392_o2,
  n2369_o2,
  n2397_o2,
  n2601_o2,
  n2658_o2,
  n2574_o2,
  n2205_o2,
  lo510_buf_o2,
  lo514_buf_o2,
  lo554_buf_o2,
  lo558_buf_o2,
  lo578_buf_o2,
  n2254_o2,
  n2421_o2,
  n2422_o2,
  n2130_o2,
  n2127_o2,
  n2131_o2,
  n2128_o2,
  n2264_o2,
  n2467_o2,
  n2471_o2,
  n2488_o2,
  n2478_o2,
  n2486_o2,
  n2485_o2,
  n2498_o2,
  n2495_o2,
  n2496_o2,
  n2458_o2,
  n2643_o2,
  n2462_o2,
  n2468_o2,
  n2639_o2,
  n2499_o2,
  n2472_o2,
  n2474_o2,
  n2489_o2,
  n2321_o2,
  n2322_o2,
  n2640_o2,
  n2642_o2,
  n2187_o2,
  n2373_o2,
  n2603_o2,
  n2388_o2,
  n2437_o2,
  n2356_o2,
  n2452_o2,
  n2347_o2,
  n2329_o2,
  n2669_o2,
  n2332_o2,
  n2664_o2,
  n2665_o2,
  n2653_o2,
  n2654_o2,
  n2636_o2,
  n2660_o2,
  n2318_o2,
  n2319_o2,
  n2586_o2,
  n2587_o2,
  n2288_o2,
  n2344_o2,
  n2530_o2,
  n2303_o2,
  n2566_o2,
  n2567_o2,
  n2554_o2,
  n2194_o2,
  lo582_buf_o2,
  lo030_buf_o2,
  lo174_buf_o2,
  lo178_buf_o2,
  lo186_buf_o2,
  lo266_buf_o2,
  lo306_buf_o2,
  lo346_buf_o2,
  lo386_buf_o2,
  lo426_buf_o2,
  lo590_buf_o2,
  lo594_buf_o2,
  lo606_buf_o2,
  lo610_buf_o2,
  n2238_o2,
  n2229_o2,
  n2242_o2,
  n2233_o2,
  n2168_o2,
  n2237_o2,
  n2228_o2,
  n2172_o2,
  n2223_o2,
  n2222_o2,
  n2170_o2,
  n2181_o2,
  n2510_o2,
  n2621_o2,
  lo466_buf_o2,
  lo478_buf_o2,
  n2149_o2,
  n2429_o2,
  n2444_o2,
  n2153_o2,
  n2433_o2,
  n2448_o2,
  n2367_o2,
  n2386_o2,
  n2539_o2,
  n2183_o2,
  n2220_o2,
  n2514_o2,
  n2196_o2,
  n2616_o2,
  n2612_o2,
  n2627_o2,
  n2140_o2,
  n1877_inv,
  lo149_buf_o2,
  lo197_buf_o2,
  lo118_buf_o2,
  lo158_buf_o2,
  lo166_buf_o2,
  lo242_buf_o2,
  lo286_buf_o2,
  lo506_buf_o2,
  n2198_o2,
  n2202_o2,
  n2197_o2,
  n1913_inv,
  n2146_o2,
  n1919_inv,
  lo312_buf_o2,
  lo316_buf_o2,
  lo352_buf_o2,
  lo356_buf_o2,
  lo392_buf_o2,
  lo396_buf_o2,
  lo432_buf_o2,
  lo436_buf_o2,
  lo576_buf_o2,
  G2531,
  G2532,
  G2533,
  G2534,
  G2535,
  G2536,
  G2537,
  G2538,
  G2539,
  G2540,
  G2541,
  G2542,
  G2543,
  G2544,
  G2545,
  G2546,
  G2547,
  G2548,
  G2549,
  G2550,
  G2551,
  G2552,
  G2553,
  G2554,
  G2555,
  G2556,
  G2557,
  G2558,
  G2559,
  G2560,
  G2561,
  G2562,
  G2563,
  G2564,
  G2565,
  G2566,
  G2567,
  G2568,
  G2569,
  G2570,
  G2571,
  G2572,
  G2573,
  G2574,
  G2575,
  G2576,
  G2577,
  G2578,
  G2579,
  G2580,
  G2581,
  G2582,
  G2583,
  G2584,
  G2585,
  G2586,
  G2587,
  G2588,
  G2589,
  G2590,
  G2591,
  G2592,
  G2593,
  G2594,
  n4649_li000_li000,
  n4652_li001_li001,
  n4655_li002_li002,
  n4658_li003_li003,
  n4661_li004_li004,
  n4664_li005_li005,
  n4667_li006_li006,
  n4670_li007_li007,
  n4673_li008_li008,
  n4676_li009_li009,
  n4679_li010_li010,
  n4682_li011_li011,
  n4685_li012_li012,
  n4688_li013_li013,
  n4691_li014_li014,
  n4697_li016_li016,
  n4700_li017_li017,
  n4703_li018_li018,
  n4709_li020_li020,
  n4712_li021_li021,
  n4715_li022_li022,
  n4721_li024_li024,
  n4724_li025_li025,
  n4727_li026_li026,
  n4730_li027_li027,
  n4733_li028_li028,
  n4736_li029_li029,
  n4745_li032_li032,
  n4748_li033_li033,
  n4751_li034_li034,
  n4754_li035_li035,
  n4757_li036_li036,
  n4760_li037_li037,
  n4763_li038_li038,
  n4766_li039_li039,
  n4769_li040_li040,
  n4772_li041_li041,
  n4775_li042_li042,
  n4778_li043_li043,
  n4781_li044_li044,
  n4784_li045_li045,
  n4787_li046_li046,
  n4793_li048_li048,
  n4796_li049_li049,
  n4799_li050_li050,
  n4805_li052_li052,
  n4808_li053_li053,
  n4811_li054_li054,
  n4817_li056_li056,
  n4820_li057_li057,
  n4823_li058_li058,
  n4829_li060_li060,
  n4832_li061_li061,
  n4835_li062_li062,
  n4841_li064_li064,
  n4844_li065_li065,
  n4847_li066_li066,
  n4853_li068_li068,
  n4856_li069_li069,
  n4859_li070_li070,
  n4865_li072_li072,
  n4868_li073_li073,
  n4871_li074_li074,
  n4877_li076_li076,
  n4880_li077_li077,
  n4883_li078_li078,
  n4889_li080_li080,
  n4892_li081_li081,
  n4895_li082_li082,
  n4901_li084_li084,
  n4904_li085_li085,
  n4907_li086_li086,
  n4913_li088_li088,
  n4916_li089_li089,
  n4919_li090_li090,
  n4925_li092_li092,
  n4928_li093_li093,
  n4931_li094_li094,
  n4937_li096_li096,
  n4940_li097_li097,
  n4943_li098_li098,
  n4949_li100_li100,
  n4952_li101_li101,
  n4955_li102_li102,
  n4961_li104_li104,
  n4964_li105_li105,
  n4967_li106_li106,
  n4973_li108_li108,
  n4976_li109_li109,
  n4979_li110_li110,
  n4982_li111_li111,
  n4985_li112_li112,
  n4988_li113_li113,
  n4991_li114_li114,
  n4994_li115_li115,
  n4997_li116_li116,
  n5009_li120_li120,
  n5021_li124_li124,
  n5024_li125_li125,
  n5027_li126_li126,
  n5030_li127_li127,
  n5033_li128_li128,
  n5036_li129_li129,
  n5045_li132_li132,
  n5048_li133_li133,
  n5057_li136_li136,
  n5060_li137_li137,
  n5069_li140_li140,
  n5072_li141_li141,
  n5081_li144_li144,
  n5084_li145_li145,
  n5093_li148_li148,
  n5105_li152_li152,
  n5108_li153_li153,
  n5117_li156_li156,
  n5129_li160_li160,
  n5132_li161_li161,
  n5141_li164_li164,
  n5153_li168_li168,
  n5156_li169_li169,
  n5159_li170_li170,
  n5162_li171_li171,
  n5165_li172_li172,
  n5168_li173_li173,
  n5177_li176_li176,
  n5180_li177_li177,
  n5189_li180_li180,
  n5192_li181_li181,
  n5195_li182_li182,
  n5201_li184_li184,
  n5204_li185_li185,
  n5213_li188_li188,
  n5216_li189_li189,
  n5225_li192_li192,
  n5228_li193_li193,
  n5237_li196_li196,
  n5249_li200_li200,
  n5252_li201_li201,
  n5261_li204_li204,
  n5273_li208_li208,
  n5276_li209_li209,
  n5279_li210_li210,
  n5282_li211_li211,
  n5285_li212_li212,
  n5288_li213_li213,
  n5297_li216_li216,
  n5300_li217_li217,
  n5309_li220_li220,
  n5312_li221_li221,
  n5321_li224_li224,
  n5324_li225_li225,
  n5333_li228_li228,
  n5336_li229_li229,
  n5345_li232_li232,
  n5348_li233_li233,
  n5357_li236_li236,
  n5360_li237_li237,
  n5369_li240_li240,
  n5381_li244_li244,
  n5384_li245_li245,
  n5393_li248_li248,
  n5405_li252_li252,
  n5408_li253_li253,
  n5411_li254_li254,
  n5414_li255_li255,
  n5417_li256_li256,
  n5420_li257_li257,
  n5429_li260_li260,
  n5432_li261_li261,
  n5441_li264_li264,
  n5444_li265_li265,
  n5453_li268_li268,
  n5456_li269_li269,
  n5465_li272_li272,
  n5468_li273_li273,
  n5477_li276_li276,
  n5480_li277_li277,
  n5489_li280_li280,
  n5492_li281_li281,
  n5501_li284_li284,
  n5513_li288_li288,
  n5516_li289_li289,
  n5525_li292_li292,
  n5528_li293_li293,
  n5531_li294_li294,
  n5534_li295_li295,
  n5537_li296_li296,
  n5540_li297_li297,
  n5549_li300_li300,
  n5552_li301_li301,
  n5555_li302_li302,
  n5558_li303_li303,
  n5561_li304_li304,
  n5564_li305_li305,
  n5573_li308_li308,
  n5576_li309_li309,
  n5609_li320_li320,
  n5612_li321_li321,
  n5621_li324_li324,
  n5624_li325_li325,
  n5633_li328_li328,
  n5636_li329_li329,
  n5645_li332_li332,
  n5648_li333_li333,
  n5657_li336_li336,
  n5660_li337_li337,
  n5669_li340_li340,
  n5672_li341_li341,
  n5675_li342_li342,
  n5678_li343_li343,
  n5681_li344_li344,
  n5684_li345_li345,
  n5693_li348_li348,
  n5696_li349_li349,
  n5729_li360_li360,
  n5732_li361_li361,
  n5741_li364_li364,
  n5744_li365_li365,
  n5753_li368_li368,
  n5756_li369_li369,
  n5765_li372_li372,
  n5768_li373_li373,
  n5777_li376_li376,
  n5780_li377_li377,
  n5789_li380_li380,
  n5792_li381_li381,
  n5795_li382_li382,
  n5798_li383_li383,
  n5801_li384_li384,
  n5804_li385_li385,
  n5813_li388_li388,
  n5816_li389_li389,
  n5849_li400_li400,
  n5852_li401_li401,
  n5861_li404_li404,
  n5864_li405_li405,
  n5873_li408_li408,
  n5876_li409_li409,
  n5885_li412_li412,
  n5888_li413_li413,
  n5897_li416_li416,
  n5900_li417_li417,
  n5909_li420_li420,
  n5912_li421_li421,
  n5915_li422_li422,
  n5918_li423_li423,
  n5921_li424_li424,
  n5924_li425_li425,
  n5933_li428_li428,
  n5936_li429_li429,
  n5969_li440_li440,
  n5972_li441_li441,
  n5981_li444_li444,
  n5984_li445_li445,
  n5993_li448_li448,
  n5996_li449_li449,
  n6005_li452_li452,
  n6008_li453_li453,
  n6017_li456_li456,
  n6020_li457_li457,
  n6023_li458_li458,
  n6026_li459_li459,
  n6029_li460_li460,
  n6032_li461_li461,
  n6035_li462_li462,
  n6038_li463_li463,
  n6041_li464_li464,
  n6053_li468_li468,
  n6056_li469_li469,
  n6059_li470_li470,
  n6062_li471_li471,
  n6065_li472_li472,
  n6068_li473_li473,
  n6071_li474_li474,
  n6074_li475_li475,
  n6077_li476_li476,
  n6089_li480_li480,
  n6092_li481_li481,
  n6095_li482_li482,
  n6098_li483_li483,
  n6101_li484_li484,
  n6104_li485_li485,
  n6107_li486_li486,
  n6110_li487_li487,
  n6113_li488_li488,
  n6116_li489_li489,
  n6119_li490_li490,
  n6122_li491_li491,
  n6125_li492_li492,
  n6128_li493_li493,
  n6131_li494_li494,
  n6134_li495_li495,
  n6137_li496_li496,
  n6140_li497_li497,
  n6149_li500_li500,
  n6152_li501_li501,
  n6158_li503_li503,
  n6161_li504_li504,
  n6173_li508_li508,
  n6176_li509_li509,
  n6185_li512_li512,
  n6188_li513_li513,
  n6194_li515_li515,
  n6197_li516_li516,
  n6200_li517_li517,
  n6203_li518_li518,
  n6209_li520_li520,
  n6212_li521_li521,
  n6215_li522_li522,
  n6221_li524_li524,
  n6224_li525_li525,
  n6227_li526_li526,
  n6230_li527_li527,
  n6233_li528_li528,
  n6236_li529_li529,
  n6239_li530_li530,
  n6245_li532_li532,
  n6248_li533_li533,
  n6251_li534_li534,
  n6254_li535_li535,
  n6257_li536_li536,
  n6260_li537_li537,
  n6263_li538_li538,
  n6266_li539_li539,
  n6269_li540_li540,
  n6272_li541_li541,
  n6278_li543_li543,
  n6281_li544_li544,
  n6284_li545_li545,
  n6287_li546_li546,
  n6290_li547_li547,
  n6293_li548_li548,
  n6296_li549_li549,
  n6302_li551_li551,
  n6305_li552_li552,
  n6308_li553_li553,
  n6314_li555_li555,
  n6317_li556_li556,
  n6320_li557_li557,
  n6326_li559_li559,
  n6329_li560_li560,
  n6332_li561_li561,
  n6335_li562_li562,
  n6338_li563_li563,
  n6341_li564_li564,
  n6344_li565_li565,
  n6347_li566_li566,
  n6350_li567_li567,
  n6353_li568_li568,
  n6356_li569_li569,
  n6359_li570_li570,
  n6362_li571_li571,
  n6365_li572_li572,
  n6368_li573_li573,
  n6371_li574_li574,
  n6374_li575_li575,
  n6389_li580_li580,
  n6401_li584_li584,
  n6404_li585_li585,
  n6407_li586_li586,
  n6410_li587_li587,
  n6413_li588_li588,
  n6416_li589_li589,
  n6425_li592_li592,
  n6428_li593_li593,
  n6437_li596_li596,
  n6440_li597_li597,
  n6443_li598_li598,
  n6449_li600_li600,
  n6452_li601_li601,
  n6455_li602_li602,
  n6461_li604_li604,
  n6464_li605_li605,
  n6473_li608_li608,
  n6476_li609_li609,
  n6485_li612_li612,
  n6488_li613_li613,
  n6491_li614_li614,
  n6497_li616_li616,
  n6500_li617_li617,
  n6503_li618_li618,
  n6509_li620_li620,
  n6512_li621_li621,
  n6515_li622_li622,
  n6521_li624_li624,
  n6524_li625_li625,
  n6527_li626_li626,
  n3603_i2,
  n3604_i2,
  n3618_i2,
  n3798_i2,
  n3846_i2,
  n4019_i2,
  n4017_i2,
  n2177_i2,
  n2150_i2,
  n2154_i2,
  n2184_i2,
  n2515_i2,
  n3837_i2,
  n2167_i2,
  n2118_i2,
  n2186_i2,
  n2174_i2,
  n3964_i2,
  n4005_i2,
  n4006_i2,
  n2195_i2,
  n2176_i2,
  n2227_i2,
  n2236_i2,
  n2245_i2,
  n2518_i2,
  n4023_i2,
  n4024_i2,
  n4038_i2,
  n4039_i2,
  n4040_i2,
  n2119_i2,
  n2275_i2,
  n2595_i2,
  n2594_i2,
  lo498_buf_i2,
  lo502_buf_i2,
  lo550_buf_i2,
  n2596_i2,
  n2593_i2,
  n2668_i2,
  lo542_buf_i2,
  n2667_i2,
  n2404_i2,
  n2410_i2,
  n2419_i2,
  n2392_i2,
  n2369_i2,
  n2397_i2,
  n2601_i2,
  n2658_i2,
  n2574_i2,
  n2205_i2,
  lo510_buf_i2,
  lo514_buf_i2,
  lo554_buf_i2,
  lo558_buf_i2,
  lo578_buf_i2,
  n2254_i2,
  n2421_i2,
  n2422_i2,
  n2130_i2,
  n2127_i2,
  n2131_i2,
  n2128_i2,
  n2264_i2,
  n2467_i2,
  n2471_i2,
  n2488_i2,
  n2478_i2,
  n2486_i2,
  n2485_i2,
  n2498_i2,
  n2495_i2,
  n2496_i2,
  n2458_i2,
  n2643_i2,
  n2462_i2,
  n2468_i2,
  n2639_i2,
  n2499_i2,
  n2472_i2,
  n2474_i2,
  n2489_i2,
  n2321_i2,
  n2322_i2,
  n2640_i2,
  n2642_i2,
  n2187_i2,
  n2373_i2,
  n2603_i2,
  n2388_i2,
  n2437_i2,
  n2356_i2,
  n2452_i2,
  n2347_i2,
  n2329_i2,
  n2669_i2,
  n2332_i2,
  n2664_i2,
  n2665_i2,
  n2653_i2,
  n2654_i2,
  n2636_i2,
  n2660_i2,
  n2318_i2,
  n2319_i2,
  n2586_i2,
  n2587_i2,
  n2288_i2,
  n2344_i2,
  n2530_i2,
  n2303_i2,
  n2566_i2,
  n2567_i2,
  n2554_i2,
  n2194_i2,
  lo582_buf_i2,
  lo030_buf_i2,
  lo174_buf_i2,
  lo178_buf_i2,
  lo186_buf_i2,
  lo266_buf_i2,
  lo306_buf_i2,
  lo346_buf_i2,
  lo386_buf_i2,
  lo426_buf_i2,
  lo590_buf_i2,
  lo594_buf_i2,
  lo606_buf_i2,
  lo610_buf_i2,
  n2238_i2,
  n2229_i2,
  n2242_i2,
  n2233_i2,
  n2168_i2,
  n2237_i2,
  n2228_i2,
  n2172_i2,
  n2223_i2,
  n2222_i2,
  n2170_i2,
  n2181_i2,
  n2510_i2,
  n2621_i2,
  lo466_buf_i2,
  lo478_buf_i2,
  n2149_i2,
  n2429_i2,
  n2444_i2,
  n2153_i2,
  n2433_i2,
  n2448_i2,
  n2367_i2,
  n2386_i2,
  n2539_i2,
  n2183_i2,
  n2220_i2,
  n2514_i2,
  n2196_i2,
  n2616_i2,
  n2612_i2,
  n2627_i2,
  n2140_i2,
  n2144_i2,
  lo149_buf_i2,
  lo197_buf_i2,
  lo118_buf_i2,
  lo158_buf_i2,
  lo166_buf_i2,
  lo242_buf_i2,
  lo286_buf_i2,
  lo506_buf_i2,
  n2198_i2,
  n2202_i2,
  n2197_i2,
  n2166_i2,
  n2146_i2,
  n2165_i2,
  lo312_buf_i2,
  lo316_buf_i2,
  lo352_buf_i2,
  lo356_buf_i2,
  lo392_buf_i2,
  lo396_buf_i2,
  lo432_buf_i2,
  lo436_buf_i2,
  lo576_buf_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input G42;input G43;input G44;input G45;input G46;input G47;input G48;input G49;input G50;input G51;input G52;input G53;input G54;input G55;input G56;input G57;input G58;input G59;input G60;input G61;input G62;input G63;input G64;input G65;input G66;input G67;input G68;input G69;input G70;input G71;input G72;input G73;input G74;input G75;input G76;input G77;input G78;input G79;input G80;input G81;input G82;input G83;input G84;input G85;input G86;input G87;input G88;input G89;input G90;input G91;input G92;input G93;input G94;input G95;input G96;input G97;input G98;input G99;input G100;input G101;input G102;input G103;input G104;input G105;input G106;input G107;input G108;input G109;input G110;input G111;input G112;input G113;input G114;input G115;input G116;input G117;input G118;input G119;input G120;input G121;input G122;input G123;input G124;input G125;input G126;input G127;input G128;input G129;input G130;input G131;input G132;input G133;input G134;input G135;input G136;input G137;input G138;input G139;input G140;input G141;input G142;input G143;input G144;input G145;input G146;input G147;input G148;input G149;input G150;input G151;input G152;input G153;input G154;input G155;input G156;input G157;input n1416_lo;input n1419_lo;input n1422_lo;input n1425_lo;input n1428_lo;input n1431_lo;input n1434_lo;input n1437_lo;input n1440_lo;input n1443_lo;input n1446_lo;input n1449_lo;input n1452_lo;input n1455_lo;input n1458_lo;input n1464_lo;input n1467_lo;input n1470_lo;input n1476_lo;input n1479_lo;input n1482_lo;input n1488_lo;input n1491_lo;input n1494_lo;input n1497_lo;input n1500_lo;input n1503_lo;input n1512_lo;input n1515_lo;input n1518_lo;input n1521_lo;input n1524_lo;input n1527_lo;input n1530_lo;input n1533_lo;input n1536_lo;input n1539_lo;input n1542_lo;input n1545_lo;input n1548_lo;input n1551_lo;input n1554_lo;input n1560_lo;input n1563_lo;input n1566_lo;input n1572_lo;input n1575_lo;input n1578_lo;input n1584_lo;input n1587_lo;input n1590_lo;input n1596_lo;input n1599_lo;input n1602_lo;input n1608_lo;input n1611_lo;input n1614_lo;input n1620_lo;input n1623_lo;input n1626_lo;input n1632_lo;input n1635_lo;input n1638_lo;input n1644_lo;input n1647_lo;input n1650_lo;input n1656_lo;input n1659_lo;input n1662_lo;input n1668_lo;input n1671_lo;input n1674_lo;input n1680_lo;input n1683_lo;input n1686_lo;input n1692_lo;input n1695_lo;input n1698_lo;input n1704_lo;input n1707_lo;input n1710_lo;input n1716_lo;input n1719_lo;input n1722_lo;input n1728_lo;input n1731_lo;input n1734_lo;input n1740_lo;input n1743_lo;input n1746_lo;input n1749_lo;input n1752_lo;input n1755_lo;input n1758_lo;input n1761_lo;input n1764_lo;input n1776_lo;input n1788_lo;input n1791_lo;input n1794_lo;input n1797_lo;input n1800_lo;input n1803_lo;input n1812_lo;input n1815_lo;input n1824_lo;input n1827_lo;input n1836_lo;input n1839_lo;input n1848_lo;input n1851_lo;input n1860_lo;input n1872_lo;input n1875_lo;input n1884_lo;input n1896_lo;input n1899_lo;input n1908_lo;input n1920_lo;input n1923_lo;input n1926_lo;input n1929_lo;input n1932_lo;input n1935_lo;input n1944_lo;input n1947_lo;input n1956_lo;input n1959_lo;input n1962_lo;input n1968_lo;input n1971_lo;input n1980_lo;input n1983_lo;input n1992_lo;input n1995_lo;input n2004_lo;input n2016_lo;input n2019_lo;input n2028_lo;input n2040_lo;input n2043_lo;input n2046_lo;input n2049_lo;input n2052_lo;input n2055_lo;input n2064_lo;input n2067_lo;input n2076_lo;input n2079_lo;input n2088_lo;input n2091_lo;input n2100_lo;input n2103_lo;input n2112_lo;input n2115_lo;input n2124_lo;input n2127_lo;input n2136_lo;input n2148_lo;input n2151_lo;input n2160_lo;input n2172_lo;input n2175_lo;input n2178_lo;input n2181_lo;input n2184_lo;input n2187_lo;input n2196_lo;input n2199_lo;input n2208_lo;input n2211_lo;input n2220_lo;input n2223_lo;input n2232_lo;input n2235_lo;input n2244_lo;input n2247_lo;input n2256_lo;input n2259_lo;input n2268_lo;input n2280_lo;input n2283_lo;input n2292_lo;input n2295_lo;input n2298_lo;input n2301_lo;input n2304_lo;input n2307_lo;input n2316_lo;input n2319_lo;input n2322_lo;input n2325_lo;input n2328_lo;input n2331_lo;input n2340_lo;input n2343_lo;input n2376_lo;input n2379_lo;input n2388_lo;input n2391_lo;input n2400_lo;input n2403_lo;input n2412_lo;input n2415_lo;input n2424_lo;input n2427_lo;input n2436_lo;input n2439_lo;input n2442_lo;input n2445_lo;input n2448_lo;input n2451_lo;input n2460_lo;input n2463_lo;input n2496_lo;input n2499_lo;input n2508_lo;input n2511_lo;input n2520_lo;input n2523_lo;input n2532_lo;input n2535_lo;input n2544_lo;input n2547_lo;input n2556_lo;input n2559_lo;input n2562_lo;input n2565_lo;input n2568_lo;input n2571_lo;input n2580_lo;input n2583_lo;input n2616_lo;input n2619_lo;input n2628_lo;input n2631_lo;input n2640_lo;input n2643_lo;input n2652_lo;input n2655_lo;input n2664_lo;input n2667_lo;input n2676_lo;input n2679_lo;input n2682_lo;input n2685_lo;input n2688_lo;input n2691_lo;input n2700_lo;input n2703_lo;input n2736_lo;input n2739_lo;input n2748_lo;input n2751_lo;input n2760_lo;input n2763_lo;input n2772_lo;input n2775_lo;input n2784_lo;input n2787_lo;input n2790_lo;input n2793_lo;input n2796_lo;input n2799_lo;input n2802_lo;input n2805_lo;input n2808_lo;input n2820_lo;input n2823_lo;input n2826_lo;input n2829_lo;input n2832_lo;input n2835_lo;input n2838_lo;input n2841_lo;input n2844_lo;input n2856_lo;input n2859_lo;input n2862_lo;input n2865_lo;input n2868_lo;input n2871_lo;input n2874_lo;input n2877_lo;input n2880_lo;input n2883_lo;input n2886_lo;input n2889_lo;input n2892_lo;input n2895_lo;input n2898_lo;input n2901_lo;input n2904_lo;input n2907_lo;input n2916_lo;input n2919_lo;input n2925_lo;input n2928_lo;input n2940_lo;input n2943_lo;input n2952_lo;input n2955_lo;input n2961_lo;input n2964_lo;input n2967_lo;input n2970_lo;input n2976_lo;input n2979_lo;input n2982_lo;input n2988_lo;input n2991_lo;input n2994_lo;input n2997_lo;input n3000_lo;input n3003_lo;input n3006_lo;input n3012_lo;input n3015_lo;input n3018_lo;input n3021_lo;input n3024_lo;input n3027_lo;input n3030_lo;input n3033_lo;input n3036_lo;input n3039_lo;input n3045_lo;input n3048_lo;input n3051_lo;input n3054_lo;input n3057_lo;input n3060_lo;input n3063_lo;input n3069_lo;input n3072_lo;input n3075_lo;input n3081_lo;input n3084_lo;input n3087_lo;input n3093_lo;input n3096_lo;input n3099_lo;input n3102_lo;input n3105_lo;input n3108_lo;input n3111_lo;input n3114_lo;input n3117_lo;input n3120_lo;input n3123_lo;input n3126_lo;input n3129_lo;input n3132_lo;input n3135_lo;input n3138_lo;input n3141_lo;input n3156_lo;input n3168_lo;input n3171_lo;input n3174_lo;input n3177_lo;input n3180_lo;input n3183_lo;input n3192_lo;input n3195_lo;input n3204_lo;input n3207_lo;input n3210_lo;input n3216_lo;input n3219_lo;input n3222_lo;input n3228_lo;input n3231_lo;input n3240_lo;input n3243_lo;input n3252_lo;input n3255_lo;input n3258_lo;input n3264_lo;input n3267_lo;input n3270_lo;input n3276_lo;input n3279_lo;input n3282_lo;input n3288_lo;input n3291_lo;input n3294_lo;input n3603_o2;input n3604_o2;input n1391_inv;input n3798_o2;input n3846_o2;input n4019_o2;input n4017_o2;input n2177_o2;input n2150_o2;input n2154_o2;input n2184_o2;input n2515_o2;input n3837_o2;input n2167_o2;input n2118_o2;input n2186_o2;input n2174_o2;input n3964_o2;input n4005_o2;input n4006_o2;input n1445_inv;input n2176_o2;input n2227_o2;input n2236_o2;input n2245_o2;input n2518_o2;input n4023_o2;input n1466_inv;input n4038_o2;input n4039_o2;input n1475_inv;input n2119_o2;input n2275_o2;input n2595_o2;input n2594_o2;input lo498_buf_o2;input lo502_buf_o2;input lo550_buf_o2;input n2596_o2;input n2593_o2;input n2668_o2;input lo542_buf_o2;input n2667_o2;input n2404_o2;input n2410_o2;input n2419_o2;input n2392_o2;input n2369_o2;input n2397_o2;input n2601_o2;input n2658_o2;input n2574_o2;input n2205_o2;input lo510_buf_o2;input lo514_buf_o2;input lo554_buf_o2;input lo558_buf_o2;input lo578_buf_o2;input n2254_o2;input n2421_o2;input n2422_o2;input n2130_o2;input n2127_o2;input n2131_o2;input n2128_o2;input n2264_o2;input n2467_o2;input n2471_o2;input n2488_o2;input n2478_o2;input n2486_o2;input n2485_o2;input n2498_o2;input n2495_o2;input n2496_o2;input n2458_o2;input n2643_o2;input n2462_o2;input n2468_o2;input n2639_o2;input n2499_o2;input n2472_o2;input n2474_o2;input n2489_o2;input n2321_o2;input n2322_o2;input n2640_o2;input n2642_o2;input n2187_o2;input n2373_o2;input n2603_o2;input n2388_o2;input n2437_o2;input n2356_o2;input n2452_o2;input n2347_o2;input n2329_o2;input n2669_o2;input n2332_o2;input n2664_o2;input n2665_o2;input n2653_o2;input n2654_o2;input n2636_o2;input n2660_o2;input n2318_o2;input n2319_o2;input n2586_o2;input n2587_o2;input n2288_o2;input n2344_o2;input n2530_o2;input n2303_o2;input n2566_o2;input n2567_o2;input n2554_o2;input n2194_o2;input lo582_buf_o2;input lo030_buf_o2;input lo174_buf_o2;input lo178_buf_o2;input lo186_buf_o2;input lo266_buf_o2;input lo306_buf_o2;input lo346_buf_o2;input lo386_buf_o2;input lo426_buf_o2;input lo590_buf_o2;input lo594_buf_o2;input lo606_buf_o2;input lo610_buf_o2;input n2238_o2;input n2229_o2;input n2242_o2;input n2233_o2;input n2168_o2;input n2237_o2;input n2228_o2;input n2172_o2;input n2223_o2;input n2222_o2;input n2170_o2;input n2181_o2;input n2510_o2;input n2621_o2;input lo466_buf_o2;input lo478_buf_o2;input n2149_o2;input n2429_o2;input n2444_o2;input n2153_o2;input n2433_o2;input n2448_o2;input n2367_o2;input n2386_o2;input n2539_o2;input n2183_o2;input n2220_o2;input n2514_o2;input n2196_o2;input n2616_o2;input n2612_o2;input n2627_o2;input n2140_o2;input n1877_inv;input lo149_buf_o2;input lo197_buf_o2;input lo118_buf_o2;input lo158_buf_o2;input lo166_buf_o2;input lo242_buf_o2;input lo286_buf_o2;input lo506_buf_o2;input n2198_o2;input n2202_o2;input n2197_o2;input n1913_inv;input n2146_o2;input n1919_inv;input lo312_buf_o2;input lo316_buf_o2;input lo352_buf_o2;input lo356_buf_o2;input lo392_buf_o2;input lo396_buf_o2;input lo432_buf_o2;input lo436_buf_o2;input lo576_buf_o2;
  output G2531;output G2532;output G2533;output G2534;output G2535;output G2536;output G2537;output G2538;output G2539;output G2540;output G2541;output G2542;output G2543;output G2544;output G2545;output G2546;output G2547;output G2548;output G2549;output G2550;output G2551;output G2552;output G2553;output G2554;output G2555;output G2556;output G2557;output G2558;output G2559;output G2560;output G2561;output G2562;output G2563;output G2564;output G2565;output G2566;output G2567;output G2568;output G2569;output G2570;output G2571;output G2572;output G2573;output G2574;output G2575;output G2576;output G2577;output G2578;output G2579;output G2580;output G2581;output G2582;output G2583;output G2584;output G2585;output G2586;output G2587;output G2588;output G2589;output G2590;output G2591;output G2592;output G2593;output G2594;output n4649_li000_li000;output n4652_li001_li001;output n4655_li002_li002;output n4658_li003_li003;output n4661_li004_li004;output n4664_li005_li005;output n4667_li006_li006;output n4670_li007_li007;output n4673_li008_li008;output n4676_li009_li009;output n4679_li010_li010;output n4682_li011_li011;output n4685_li012_li012;output n4688_li013_li013;output n4691_li014_li014;output n4697_li016_li016;output n4700_li017_li017;output n4703_li018_li018;output n4709_li020_li020;output n4712_li021_li021;output n4715_li022_li022;output n4721_li024_li024;output n4724_li025_li025;output n4727_li026_li026;output n4730_li027_li027;output n4733_li028_li028;output n4736_li029_li029;output n4745_li032_li032;output n4748_li033_li033;output n4751_li034_li034;output n4754_li035_li035;output n4757_li036_li036;output n4760_li037_li037;output n4763_li038_li038;output n4766_li039_li039;output n4769_li040_li040;output n4772_li041_li041;output n4775_li042_li042;output n4778_li043_li043;output n4781_li044_li044;output n4784_li045_li045;output n4787_li046_li046;output n4793_li048_li048;output n4796_li049_li049;output n4799_li050_li050;output n4805_li052_li052;output n4808_li053_li053;output n4811_li054_li054;output n4817_li056_li056;output n4820_li057_li057;output n4823_li058_li058;output n4829_li060_li060;output n4832_li061_li061;output n4835_li062_li062;output n4841_li064_li064;output n4844_li065_li065;output n4847_li066_li066;output n4853_li068_li068;output n4856_li069_li069;output n4859_li070_li070;output n4865_li072_li072;output n4868_li073_li073;output n4871_li074_li074;output n4877_li076_li076;output n4880_li077_li077;output n4883_li078_li078;output n4889_li080_li080;output n4892_li081_li081;output n4895_li082_li082;output n4901_li084_li084;output n4904_li085_li085;output n4907_li086_li086;output n4913_li088_li088;output n4916_li089_li089;output n4919_li090_li090;output n4925_li092_li092;output n4928_li093_li093;output n4931_li094_li094;output n4937_li096_li096;output n4940_li097_li097;output n4943_li098_li098;output n4949_li100_li100;output n4952_li101_li101;output n4955_li102_li102;output n4961_li104_li104;output n4964_li105_li105;output n4967_li106_li106;output n4973_li108_li108;output n4976_li109_li109;output n4979_li110_li110;output n4982_li111_li111;output n4985_li112_li112;output n4988_li113_li113;output n4991_li114_li114;output n4994_li115_li115;output n4997_li116_li116;output n5009_li120_li120;output n5021_li124_li124;output n5024_li125_li125;output n5027_li126_li126;output n5030_li127_li127;output n5033_li128_li128;output n5036_li129_li129;output n5045_li132_li132;output n5048_li133_li133;output n5057_li136_li136;output n5060_li137_li137;output n5069_li140_li140;output n5072_li141_li141;output n5081_li144_li144;output n5084_li145_li145;output n5093_li148_li148;output n5105_li152_li152;output n5108_li153_li153;output n5117_li156_li156;output n5129_li160_li160;output n5132_li161_li161;output n5141_li164_li164;output n5153_li168_li168;output n5156_li169_li169;output n5159_li170_li170;output n5162_li171_li171;output n5165_li172_li172;output n5168_li173_li173;output n5177_li176_li176;output n5180_li177_li177;output n5189_li180_li180;output n5192_li181_li181;output n5195_li182_li182;output n5201_li184_li184;output n5204_li185_li185;output n5213_li188_li188;output n5216_li189_li189;output n5225_li192_li192;output n5228_li193_li193;output n5237_li196_li196;output n5249_li200_li200;output n5252_li201_li201;output n5261_li204_li204;output n5273_li208_li208;output n5276_li209_li209;output n5279_li210_li210;output n5282_li211_li211;output n5285_li212_li212;output n5288_li213_li213;output n5297_li216_li216;output n5300_li217_li217;output n5309_li220_li220;output n5312_li221_li221;output n5321_li224_li224;output n5324_li225_li225;output n5333_li228_li228;output n5336_li229_li229;output n5345_li232_li232;output n5348_li233_li233;output n5357_li236_li236;output n5360_li237_li237;output n5369_li240_li240;output n5381_li244_li244;output n5384_li245_li245;output n5393_li248_li248;output n5405_li252_li252;output n5408_li253_li253;output n5411_li254_li254;output n5414_li255_li255;output n5417_li256_li256;output n5420_li257_li257;output n5429_li260_li260;output n5432_li261_li261;output n5441_li264_li264;output n5444_li265_li265;output n5453_li268_li268;output n5456_li269_li269;output n5465_li272_li272;output n5468_li273_li273;output n5477_li276_li276;output n5480_li277_li277;output n5489_li280_li280;output n5492_li281_li281;output n5501_li284_li284;output n5513_li288_li288;output n5516_li289_li289;output n5525_li292_li292;output n5528_li293_li293;output n5531_li294_li294;output n5534_li295_li295;output n5537_li296_li296;output n5540_li297_li297;output n5549_li300_li300;output n5552_li301_li301;output n5555_li302_li302;output n5558_li303_li303;output n5561_li304_li304;output n5564_li305_li305;output n5573_li308_li308;output n5576_li309_li309;output n5609_li320_li320;output n5612_li321_li321;output n5621_li324_li324;output n5624_li325_li325;output n5633_li328_li328;output n5636_li329_li329;output n5645_li332_li332;output n5648_li333_li333;output n5657_li336_li336;output n5660_li337_li337;output n5669_li340_li340;output n5672_li341_li341;output n5675_li342_li342;output n5678_li343_li343;output n5681_li344_li344;output n5684_li345_li345;output n5693_li348_li348;output n5696_li349_li349;output n5729_li360_li360;output n5732_li361_li361;output n5741_li364_li364;output n5744_li365_li365;output n5753_li368_li368;output n5756_li369_li369;output n5765_li372_li372;output n5768_li373_li373;output n5777_li376_li376;output n5780_li377_li377;output n5789_li380_li380;output n5792_li381_li381;output n5795_li382_li382;output n5798_li383_li383;output n5801_li384_li384;output n5804_li385_li385;output n5813_li388_li388;output n5816_li389_li389;output n5849_li400_li400;output n5852_li401_li401;output n5861_li404_li404;output n5864_li405_li405;output n5873_li408_li408;output n5876_li409_li409;output n5885_li412_li412;output n5888_li413_li413;output n5897_li416_li416;output n5900_li417_li417;output n5909_li420_li420;output n5912_li421_li421;output n5915_li422_li422;output n5918_li423_li423;output n5921_li424_li424;output n5924_li425_li425;output n5933_li428_li428;output n5936_li429_li429;output n5969_li440_li440;output n5972_li441_li441;output n5981_li444_li444;output n5984_li445_li445;output n5993_li448_li448;output n5996_li449_li449;output n6005_li452_li452;output n6008_li453_li453;output n6017_li456_li456;output n6020_li457_li457;output n6023_li458_li458;output n6026_li459_li459;output n6029_li460_li460;output n6032_li461_li461;output n6035_li462_li462;output n6038_li463_li463;output n6041_li464_li464;output n6053_li468_li468;output n6056_li469_li469;output n6059_li470_li470;output n6062_li471_li471;output n6065_li472_li472;output n6068_li473_li473;output n6071_li474_li474;output n6074_li475_li475;output n6077_li476_li476;output n6089_li480_li480;output n6092_li481_li481;output n6095_li482_li482;output n6098_li483_li483;output n6101_li484_li484;output n6104_li485_li485;output n6107_li486_li486;output n6110_li487_li487;output n6113_li488_li488;output n6116_li489_li489;output n6119_li490_li490;output n6122_li491_li491;output n6125_li492_li492;output n6128_li493_li493;output n6131_li494_li494;output n6134_li495_li495;output n6137_li496_li496;output n6140_li497_li497;output n6149_li500_li500;output n6152_li501_li501;output n6158_li503_li503;output n6161_li504_li504;output n6173_li508_li508;output n6176_li509_li509;output n6185_li512_li512;output n6188_li513_li513;output n6194_li515_li515;output n6197_li516_li516;output n6200_li517_li517;output n6203_li518_li518;output n6209_li520_li520;output n6212_li521_li521;output n6215_li522_li522;output n6221_li524_li524;output n6224_li525_li525;output n6227_li526_li526;output n6230_li527_li527;output n6233_li528_li528;output n6236_li529_li529;output n6239_li530_li530;output n6245_li532_li532;output n6248_li533_li533;output n6251_li534_li534;output n6254_li535_li535;output n6257_li536_li536;output n6260_li537_li537;output n6263_li538_li538;output n6266_li539_li539;output n6269_li540_li540;output n6272_li541_li541;output n6278_li543_li543;output n6281_li544_li544;output n6284_li545_li545;output n6287_li546_li546;output n6290_li547_li547;output n6293_li548_li548;output n6296_li549_li549;output n6302_li551_li551;output n6305_li552_li552;output n6308_li553_li553;output n6314_li555_li555;output n6317_li556_li556;output n6320_li557_li557;output n6326_li559_li559;output n6329_li560_li560;output n6332_li561_li561;output n6335_li562_li562;output n6338_li563_li563;output n6341_li564_li564;output n6344_li565_li565;output n6347_li566_li566;output n6350_li567_li567;output n6353_li568_li568;output n6356_li569_li569;output n6359_li570_li570;output n6362_li571_li571;output n6365_li572_li572;output n6368_li573_li573;output n6371_li574_li574;output n6374_li575_li575;output n6389_li580_li580;output n6401_li584_li584;output n6404_li585_li585;output n6407_li586_li586;output n6410_li587_li587;output n6413_li588_li588;output n6416_li589_li589;output n6425_li592_li592;output n6428_li593_li593;output n6437_li596_li596;output n6440_li597_li597;output n6443_li598_li598;output n6449_li600_li600;output n6452_li601_li601;output n6455_li602_li602;output n6461_li604_li604;output n6464_li605_li605;output n6473_li608_li608;output n6476_li609_li609;output n6485_li612_li612;output n6488_li613_li613;output n6491_li614_li614;output n6497_li616_li616;output n6500_li617_li617;output n6503_li618_li618;output n6509_li620_li620;output n6512_li621_li621;output n6515_li622_li622;output n6521_li624_li624;output n6524_li625_li625;output n6527_li626_li626;output n3603_i2;output n3604_i2;output n3618_i2;output n3798_i2;output n3846_i2;output n4019_i2;output n4017_i2;output n2177_i2;output n2150_i2;output n2154_i2;output n2184_i2;output n2515_i2;output n3837_i2;output n2167_i2;output n2118_i2;output n2186_i2;output n2174_i2;output n3964_i2;output n4005_i2;output n4006_i2;output n2195_i2;output n2176_i2;output n2227_i2;output n2236_i2;output n2245_i2;output n2518_i2;output n4023_i2;output n4024_i2;output n4038_i2;output n4039_i2;output n4040_i2;output n2119_i2;output n2275_i2;output n2595_i2;output n2594_i2;output lo498_buf_i2;output lo502_buf_i2;output lo550_buf_i2;output n2596_i2;output n2593_i2;output n2668_i2;output lo542_buf_i2;output n2667_i2;output n2404_i2;output n2410_i2;output n2419_i2;output n2392_i2;output n2369_i2;output n2397_i2;output n2601_i2;output n2658_i2;output n2574_i2;output n2205_i2;output lo510_buf_i2;output lo514_buf_i2;output lo554_buf_i2;output lo558_buf_i2;output lo578_buf_i2;output n2254_i2;output n2421_i2;output n2422_i2;output n2130_i2;output n2127_i2;output n2131_i2;output n2128_i2;output n2264_i2;output n2467_i2;output n2471_i2;output n2488_i2;output n2478_i2;output n2486_i2;output n2485_i2;output n2498_i2;output n2495_i2;output n2496_i2;output n2458_i2;output n2643_i2;output n2462_i2;output n2468_i2;output n2639_i2;output n2499_i2;output n2472_i2;output n2474_i2;output n2489_i2;output n2321_i2;output n2322_i2;output n2640_i2;output n2642_i2;output n2187_i2;output n2373_i2;output n2603_i2;output n2388_i2;output n2437_i2;output n2356_i2;output n2452_i2;output n2347_i2;output n2329_i2;output n2669_i2;output n2332_i2;output n2664_i2;output n2665_i2;output n2653_i2;output n2654_i2;output n2636_i2;output n2660_i2;output n2318_i2;output n2319_i2;output n2586_i2;output n2587_i2;output n2288_i2;output n2344_i2;output n2530_i2;output n2303_i2;output n2566_i2;output n2567_i2;output n2554_i2;output n2194_i2;output lo582_buf_i2;output lo030_buf_i2;output lo174_buf_i2;output lo178_buf_i2;output lo186_buf_i2;output lo266_buf_i2;output lo306_buf_i2;output lo346_buf_i2;output lo386_buf_i2;output lo426_buf_i2;output lo590_buf_i2;output lo594_buf_i2;output lo606_buf_i2;output lo610_buf_i2;output n2238_i2;output n2229_i2;output n2242_i2;output n2233_i2;output n2168_i2;output n2237_i2;output n2228_i2;output n2172_i2;output n2223_i2;output n2222_i2;output n2170_i2;output n2181_i2;output n2510_i2;output n2621_i2;output lo466_buf_i2;output lo478_buf_i2;output n2149_i2;output n2429_i2;output n2444_i2;output n2153_i2;output n2433_i2;output n2448_i2;output n2367_i2;output n2386_i2;output n2539_i2;output n2183_i2;output n2220_i2;output n2514_i2;output n2196_i2;output n2616_i2;output n2612_i2;output n2627_i2;output n2140_i2;output n2144_i2;output lo149_buf_i2;output lo197_buf_i2;output lo118_buf_i2;output lo158_buf_i2;output lo166_buf_i2;output lo242_buf_i2;output lo286_buf_i2;output lo506_buf_i2;output n2198_i2;output n2202_i2;output n2197_i2;output n2166_i2;output n2146_i2;output n2165_i2;output lo312_buf_i2;output lo316_buf_i2;output lo352_buf_i2;output lo356_buf_i2;output lo392_buf_i2;output lo396_buf_i2;output lo432_buf_i2;output lo436_buf_i2;output lo576_buf_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire G42_p;
  wire G42_n;
  wire G43_p;
  wire G43_n;
  wire G44_p;
  wire G44_n;
  wire G45_p;
  wire G45_n;
  wire G46_p;
  wire G46_n;
  wire G47_p;
  wire G47_n;
  wire G48_p;
  wire G48_n;
  wire G49_p;
  wire G49_n;
  wire G50_p;
  wire G50_n;
  wire G51_p;
  wire G51_n;
  wire G52_p;
  wire G52_n;
  wire G53_p;
  wire G53_n;
  wire G54_p;
  wire G54_n;
  wire G55_p;
  wire G55_n;
  wire G56_p;
  wire G56_n;
  wire G57_p;
  wire G57_n;
  wire G58_p;
  wire G58_n;
  wire G59_p;
  wire G59_n;
  wire G60_p;
  wire G60_n;
  wire G61_p;
  wire G61_n;
  wire G62_p;
  wire G62_n;
  wire G63_p;
  wire G63_n;
  wire G64_p;
  wire G64_n;
  wire G65_p;
  wire G65_n;
  wire G66_p;
  wire G66_n;
  wire G67_p;
  wire G67_n;
  wire G68_p;
  wire G68_n;
  wire G69_p;
  wire G69_n;
  wire G70_p;
  wire G70_n;
  wire G71_p;
  wire G71_n;
  wire G72_p;
  wire G72_n;
  wire G73_p;
  wire G73_n;
  wire G74_p;
  wire G74_n;
  wire G75_p;
  wire G75_n;
  wire G76_p;
  wire G76_n;
  wire G77_p;
  wire G77_n;
  wire G78_p;
  wire G78_n;
  wire G79_p;
  wire G79_n;
  wire G80_p;
  wire G80_n;
  wire G81_p;
  wire G81_n;
  wire G82_p;
  wire G82_n;
  wire G83_p;
  wire G83_n;
  wire G84_p;
  wire G84_n;
  wire G85_p;
  wire G85_n;
  wire G86_p;
  wire G86_n;
  wire G87_p;
  wire G87_n;
  wire G88_p;
  wire G88_n;
  wire G89_p;
  wire G89_n;
  wire G90_p;
  wire G90_n;
  wire G91_p;
  wire G91_n;
  wire G92_p;
  wire G92_n;
  wire G93_p;
  wire G93_n;
  wire G94_p;
  wire G94_n;
  wire G95_p;
  wire G95_n;
  wire G96_p;
  wire G96_n;
  wire G97_p;
  wire G97_n;
  wire G98_p;
  wire G98_n;
  wire G99_p;
  wire G99_n;
  wire G100_p;
  wire G100_n;
  wire G101_p;
  wire G101_n;
  wire G102_p;
  wire G102_n;
  wire G103_p;
  wire G103_n;
  wire G104_p;
  wire G104_n;
  wire G105_p;
  wire G105_n;
  wire G106_p;
  wire G106_n;
  wire G107_p;
  wire G107_n;
  wire G108_p;
  wire G108_n;
  wire G109_p;
  wire G109_n;
  wire G110_p;
  wire G110_n;
  wire G111_p;
  wire G111_n;
  wire G112_p;
  wire G112_n;
  wire G113_p;
  wire G113_n;
  wire G114_p;
  wire G114_n;
  wire G115_p;
  wire G115_n;
  wire G116_p;
  wire G116_n;
  wire G117_p;
  wire G117_n;
  wire G118_p;
  wire G118_n;
  wire G119_p;
  wire G119_n;
  wire G120_p;
  wire G120_n;
  wire G121_p;
  wire G121_n;
  wire G122_p;
  wire G122_n;
  wire G123_p;
  wire G123_n;
  wire G124_p;
  wire G124_n;
  wire G125_p;
  wire G125_n;
  wire G126_p;
  wire G126_n;
  wire G127_p;
  wire G127_n;
  wire G128_p;
  wire G128_n;
  wire G129_p;
  wire G129_n;
  wire G130_p;
  wire G130_n;
  wire G131_p;
  wire G131_n;
  wire G132_p;
  wire G132_n;
  wire G133_p;
  wire G133_n;
  wire G134_p;
  wire G134_n;
  wire G135_p;
  wire G135_n;
  wire G136_p;
  wire G136_n;
  wire G137_p;
  wire G137_n;
  wire G138_p;
  wire G138_n;
  wire G139_p;
  wire G139_n;
  wire G140_p;
  wire G140_n;
  wire G141_p;
  wire G141_n;
  wire G142_p;
  wire G142_n;
  wire G143_p;
  wire G143_n;
  wire G144_p;
  wire G144_n;
  wire G145_p;
  wire G145_n;
  wire G146_p;
  wire G146_n;
  wire G147_p;
  wire G147_n;
  wire G148_p;
  wire G148_n;
  wire G149_p;
  wire G149_n;
  wire G150_p;
  wire G150_n;
  wire G151_p;
  wire G151_n;
  wire G152_p;
  wire G152_n;
  wire G153_p;
  wire G153_n;
  wire G154_p;
  wire G154_n;
  wire G155_p;
  wire G155_n;
  wire G156_p;
  wire G156_n;
  wire G157_p;
  wire G157_n;
  wire n1416_lo_p;
  wire n1416_lo_n;
  wire n1419_lo_p;
  wire n1419_lo_n;
  wire n1422_lo_p;
  wire n1422_lo_n;
  wire n1425_lo_p;
  wire n1425_lo_n;
  wire n1428_lo_p;
  wire n1428_lo_n;
  wire n1431_lo_p;
  wire n1431_lo_n;
  wire n1434_lo_p;
  wire n1434_lo_n;
  wire n1437_lo_p;
  wire n1437_lo_n;
  wire n1440_lo_p;
  wire n1440_lo_n;
  wire n1443_lo_p;
  wire n1443_lo_n;
  wire n1446_lo_p;
  wire n1446_lo_n;
  wire n1449_lo_p;
  wire n1449_lo_n;
  wire n1452_lo_p;
  wire n1452_lo_n;
  wire n1455_lo_p;
  wire n1455_lo_n;
  wire n1458_lo_p;
  wire n1458_lo_n;
  wire n1464_lo_p;
  wire n1464_lo_n;
  wire n1467_lo_p;
  wire n1467_lo_n;
  wire n1470_lo_p;
  wire n1470_lo_n;
  wire n1476_lo_p;
  wire n1476_lo_n;
  wire n1479_lo_p;
  wire n1479_lo_n;
  wire n1482_lo_p;
  wire n1482_lo_n;
  wire n1488_lo_p;
  wire n1488_lo_n;
  wire n1491_lo_p;
  wire n1491_lo_n;
  wire n1494_lo_p;
  wire n1494_lo_n;
  wire n1497_lo_p;
  wire n1497_lo_n;
  wire n1500_lo_p;
  wire n1500_lo_n;
  wire n1503_lo_p;
  wire n1503_lo_n;
  wire n1512_lo_p;
  wire n1512_lo_n;
  wire n1515_lo_p;
  wire n1515_lo_n;
  wire n1518_lo_p;
  wire n1518_lo_n;
  wire n1521_lo_p;
  wire n1521_lo_n;
  wire n1524_lo_p;
  wire n1524_lo_n;
  wire n1527_lo_p;
  wire n1527_lo_n;
  wire n1530_lo_p;
  wire n1530_lo_n;
  wire n1533_lo_p;
  wire n1533_lo_n;
  wire n1536_lo_p;
  wire n1536_lo_n;
  wire n1539_lo_p;
  wire n1539_lo_n;
  wire n1542_lo_p;
  wire n1542_lo_n;
  wire n1545_lo_p;
  wire n1545_lo_n;
  wire n1548_lo_p;
  wire n1548_lo_n;
  wire n1551_lo_p;
  wire n1551_lo_n;
  wire n1554_lo_p;
  wire n1554_lo_n;
  wire n1560_lo_p;
  wire n1560_lo_n;
  wire n1563_lo_p;
  wire n1563_lo_n;
  wire n1566_lo_p;
  wire n1566_lo_n;
  wire n1572_lo_p;
  wire n1572_lo_n;
  wire n1575_lo_p;
  wire n1575_lo_n;
  wire n1578_lo_p;
  wire n1578_lo_n;
  wire n1584_lo_p;
  wire n1584_lo_n;
  wire n1587_lo_p;
  wire n1587_lo_n;
  wire n1590_lo_p;
  wire n1590_lo_n;
  wire n1596_lo_p;
  wire n1596_lo_n;
  wire n1599_lo_p;
  wire n1599_lo_n;
  wire n1602_lo_p;
  wire n1602_lo_n;
  wire n1608_lo_p;
  wire n1608_lo_n;
  wire n1611_lo_p;
  wire n1611_lo_n;
  wire n1614_lo_p;
  wire n1614_lo_n;
  wire n1620_lo_p;
  wire n1620_lo_n;
  wire n1623_lo_p;
  wire n1623_lo_n;
  wire n1626_lo_p;
  wire n1626_lo_n;
  wire n1632_lo_p;
  wire n1632_lo_n;
  wire n1635_lo_p;
  wire n1635_lo_n;
  wire n1638_lo_p;
  wire n1638_lo_n;
  wire n1644_lo_p;
  wire n1644_lo_n;
  wire n1647_lo_p;
  wire n1647_lo_n;
  wire n1650_lo_p;
  wire n1650_lo_n;
  wire n1656_lo_p;
  wire n1656_lo_n;
  wire n1659_lo_p;
  wire n1659_lo_n;
  wire n1662_lo_p;
  wire n1662_lo_n;
  wire n1668_lo_p;
  wire n1668_lo_n;
  wire n1671_lo_p;
  wire n1671_lo_n;
  wire n1674_lo_p;
  wire n1674_lo_n;
  wire n1680_lo_p;
  wire n1680_lo_n;
  wire n1683_lo_p;
  wire n1683_lo_n;
  wire n1686_lo_p;
  wire n1686_lo_n;
  wire n1692_lo_p;
  wire n1692_lo_n;
  wire n1695_lo_p;
  wire n1695_lo_n;
  wire n1698_lo_p;
  wire n1698_lo_n;
  wire n1704_lo_p;
  wire n1704_lo_n;
  wire n1707_lo_p;
  wire n1707_lo_n;
  wire n1710_lo_p;
  wire n1710_lo_n;
  wire n1716_lo_p;
  wire n1716_lo_n;
  wire n1719_lo_p;
  wire n1719_lo_n;
  wire n1722_lo_p;
  wire n1722_lo_n;
  wire n1728_lo_p;
  wire n1728_lo_n;
  wire n1731_lo_p;
  wire n1731_lo_n;
  wire n1734_lo_p;
  wire n1734_lo_n;
  wire n1740_lo_p;
  wire n1740_lo_n;
  wire n1743_lo_p;
  wire n1743_lo_n;
  wire n1746_lo_p;
  wire n1746_lo_n;
  wire n1749_lo_p;
  wire n1749_lo_n;
  wire n1752_lo_p;
  wire n1752_lo_n;
  wire n1755_lo_p;
  wire n1755_lo_n;
  wire n1758_lo_p;
  wire n1758_lo_n;
  wire n1761_lo_p;
  wire n1761_lo_n;
  wire n1764_lo_p;
  wire n1764_lo_n;
  wire n1776_lo_p;
  wire n1776_lo_n;
  wire n1788_lo_p;
  wire n1788_lo_n;
  wire n1791_lo_p;
  wire n1791_lo_n;
  wire n1794_lo_p;
  wire n1794_lo_n;
  wire n1797_lo_p;
  wire n1797_lo_n;
  wire n1800_lo_p;
  wire n1800_lo_n;
  wire n1803_lo_p;
  wire n1803_lo_n;
  wire n1812_lo_p;
  wire n1812_lo_n;
  wire n1815_lo_p;
  wire n1815_lo_n;
  wire n1824_lo_p;
  wire n1824_lo_n;
  wire n1827_lo_p;
  wire n1827_lo_n;
  wire n1836_lo_p;
  wire n1836_lo_n;
  wire n1839_lo_p;
  wire n1839_lo_n;
  wire n1848_lo_p;
  wire n1848_lo_n;
  wire n1851_lo_p;
  wire n1851_lo_n;
  wire n1860_lo_p;
  wire n1860_lo_n;
  wire n1872_lo_p;
  wire n1872_lo_n;
  wire n1875_lo_p;
  wire n1875_lo_n;
  wire n1884_lo_p;
  wire n1884_lo_n;
  wire n1896_lo_p;
  wire n1896_lo_n;
  wire n1899_lo_p;
  wire n1899_lo_n;
  wire n1908_lo_p;
  wire n1908_lo_n;
  wire n1920_lo_p;
  wire n1920_lo_n;
  wire n1923_lo_p;
  wire n1923_lo_n;
  wire n1926_lo_p;
  wire n1926_lo_n;
  wire n1929_lo_p;
  wire n1929_lo_n;
  wire n1932_lo_p;
  wire n1932_lo_n;
  wire n1935_lo_p;
  wire n1935_lo_n;
  wire n1944_lo_p;
  wire n1944_lo_n;
  wire n1947_lo_p;
  wire n1947_lo_n;
  wire n1956_lo_p;
  wire n1956_lo_n;
  wire n1959_lo_p;
  wire n1959_lo_n;
  wire n1962_lo_p;
  wire n1962_lo_n;
  wire n1968_lo_p;
  wire n1968_lo_n;
  wire n1971_lo_p;
  wire n1971_lo_n;
  wire n1980_lo_p;
  wire n1980_lo_n;
  wire n1983_lo_p;
  wire n1983_lo_n;
  wire n1992_lo_p;
  wire n1992_lo_n;
  wire n1995_lo_p;
  wire n1995_lo_n;
  wire n2004_lo_p;
  wire n2004_lo_n;
  wire n2016_lo_p;
  wire n2016_lo_n;
  wire n2019_lo_p;
  wire n2019_lo_n;
  wire n2028_lo_p;
  wire n2028_lo_n;
  wire n2040_lo_p;
  wire n2040_lo_n;
  wire n2043_lo_p;
  wire n2043_lo_n;
  wire n2046_lo_p;
  wire n2046_lo_n;
  wire n2049_lo_p;
  wire n2049_lo_n;
  wire n2052_lo_p;
  wire n2052_lo_n;
  wire n2055_lo_p;
  wire n2055_lo_n;
  wire n2064_lo_p;
  wire n2064_lo_n;
  wire n2067_lo_p;
  wire n2067_lo_n;
  wire n2076_lo_p;
  wire n2076_lo_n;
  wire n2079_lo_p;
  wire n2079_lo_n;
  wire n2088_lo_p;
  wire n2088_lo_n;
  wire n2091_lo_p;
  wire n2091_lo_n;
  wire n2100_lo_p;
  wire n2100_lo_n;
  wire n2103_lo_p;
  wire n2103_lo_n;
  wire n2112_lo_p;
  wire n2112_lo_n;
  wire n2115_lo_p;
  wire n2115_lo_n;
  wire n2124_lo_p;
  wire n2124_lo_n;
  wire n2127_lo_p;
  wire n2127_lo_n;
  wire n2136_lo_p;
  wire n2136_lo_n;
  wire n2148_lo_p;
  wire n2148_lo_n;
  wire n2151_lo_p;
  wire n2151_lo_n;
  wire n2160_lo_p;
  wire n2160_lo_n;
  wire n2172_lo_p;
  wire n2172_lo_n;
  wire n2175_lo_p;
  wire n2175_lo_n;
  wire n2178_lo_p;
  wire n2178_lo_n;
  wire n2181_lo_p;
  wire n2181_lo_n;
  wire n2184_lo_p;
  wire n2184_lo_n;
  wire n2187_lo_p;
  wire n2187_lo_n;
  wire n2196_lo_p;
  wire n2196_lo_n;
  wire n2199_lo_p;
  wire n2199_lo_n;
  wire n2208_lo_p;
  wire n2208_lo_n;
  wire n2211_lo_p;
  wire n2211_lo_n;
  wire n2220_lo_p;
  wire n2220_lo_n;
  wire n2223_lo_p;
  wire n2223_lo_n;
  wire n2232_lo_p;
  wire n2232_lo_n;
  wire n2235_lo_p;
  wire n2235_lo_n;
  wire n2244_lo_p;
  wire n2244_lo_n;
  wire n2247_lo_p;
  wire n2247_lo_n;
  wire n2256_lo_p;
  wire n2256_lo_n;
  wire n2259_lo_p;
  wire n2259_lo_n;
  wire n2268_lo_p;
  wire n2268_lo_n;
  wire n2280_lo_p;
  wire n2280_lo_n;
  wire n2283_lo_p;
  wire n2283_lo_n;
  wire n2292_lo_p;
  wire n2292_lo_n;
  wire n2295_lo_p;
  wire n2295_lo_n;
  wire n2298_lo_p;
  wire n2298_lo_n;
  wire n2301_lo_p;
  wire n2301_lo_n;
  wire n2304_lo_p;
  wire n2304_lo_n;
  wire n2307_lo_p;
  wire n2307_lo_n;
  wire n2316_lo_p;
  wire n2316_lo_n;
  wire n2319_lo_p;
  wire n2319_lo_n;
  wire n2322_lo_p;
  wire n2322_lo_n;
  wire n2325_lo_p;
  wire n2325_lo_n;
  wire n2328_lo_p;
  wire n2328_lo_n;
  wire n2331_lo_p;
  wire n2331_lo_n;
  wire n2340_lo_p;
  wire n2340_lo_n;
  wire n2343_lo_p;
  wire n2343_lo_n;
  wire n2376_lo_p;
  wire n2376_lo_n;
  wire n2379_lo_p;
  wire n2379_lo_n;
  wire n2388_lo_p;
  wire n2388_lo_n;
  wire n2391_lo_p;
  wire n2391_lo_n;
  wire n2400_lo_p;
  wire n2400_lo_n;
  wire n2403_lo_p;
  wire n2403_lo_n;
  wire n2412_lo_p;
  wire n2412_lo_n;
  wire n2415_lo_p;
  wire n2415_lo_n;
  wire n2424_lo_p;
  wire n2424_lo_n;
  wire n2427_lo_p;
  wire n2427_lo_n;
  wire n2436_lo_p;
  wire n2436_lo_n;
  wire n2439_lo_p;
  wire n2439_lo_n;
  wire n2442_lo_p;
  wire n2442_lo_n;
  wire n2445_lo_p;
  wire n2445_lo_n;
  wire n2448_lo_p;
  wire n2448_lo_n;
  wire n2451_lo_p;
  wire n2451_lo_n;
  wire n2460_lo_p;
  wire n2460_lo_n;
  wire n2463_lo_p;
  wire n2463_lo_n;
  wire n2496_lo_p;
  wire n2496_lo_n;
  wire n2499_lo_p;
  wire n2499_lo_n;
  wire n2508_lo_p;
  wire n2508_lo_n;
  wire n2511_lo_p;
  wire n2511_lo_n;
  wire n2520_lo_p;
  wire n2520_lo_n;
  wire n2523_lo_p;
  wire n2523_lo_n;
  wire n2532_lo_p;
  wire n2532_lo_n;
  wire n2535_lo_p;
  wire n2535_lo_n;
  wire n2544_lo_p;
  wire n2544_lo_n;
  wire n2547_lo_p;
  wire n2547_lo_n;
  wire n2556_lo_p;
  wire n2556_lo_n;
  wire n2559_lo_p;
  wire n2559_lo_n;
  wire n2562_lo_p;
  wire n2562_lo_n;
  wire n2565_lo_p;
  wire n2565_lo_n;
  wire n2568_lo_p;
  wire n2568_lo_n;
  wire n2571_lo_p;
  wire n2571_lo_n;
  wire n2580_lo_p;
  wire n2580_lo_n;
  wire n2583_lo_p;
  wire n2583_lo_n;
  wire n2616_lo_p;
  wire n2616_lo_n;
  wire n2619_lo_p;
  wire n2619_lo_n;
  wire n2628_lo_p;
  wire n2628_lo_n;
  wire n2631_lo_p;
  wire n2631_lo_n;
  wire n2640_lo_p;
  wire n2640_lo_n;
  wire n2643_lo_p;
  wire n2643_lo_n;
  wire n2652_lo_p;
  wire n2652_lo_n;
  wire n2655_lo_p;
  wire n2655_lo_n;
  wire n2664_lo_p;
  wire n2664_lo_n;
  wire n2667_lo_p;
  wire n2667_lo_n;
  wire n2676_lo_p;
  wire n2676_lo_n;
  wire n2679_lo_p;
  wire n2679_lo_n;
  wire n2682_lo_p;
  wire n2682_lo_n;
  wire n2685_lo_p;
  wire n2685_lo_n;
  wire n2688_lo_p;
  wire n2688_lo_n;
  wire n2691_lo_p;
  wire n2691_lo_n;
  wire n2700_lo_p;
  wire n2700_lo_n;
  wire n2703_lo_p;
  wire n2703_lo_n;
  wire n2736_lo_p;
  wire n2736_lo_n;
  wire n2739_lo_p;
  wire n2739_lo_n;
  wire n2748_lo_p;
  wire n2748_lo_n;
  wire n2751_lo_p;
  wire n2751_lo_n;
  wire n2760_lo_p;
  wire n2760_lo_n;
  wire n2763_lo_p;
  wire n2763_lo_n;
  wire n2772_lo_p;
  wire n2772_lo_n;
  wire n2775_lo_p;
  wire n2775_lo_n;
  wire n2784_lo_p;
  wire n2784_lo_n;
  wire n2787_lo_p;
  wire n2787_lo_n;
  wire n2790_lo_p;
  wire n2790_lo_n;
  wire n2793_lo_p;
  wire n2793_lo_n;
  wire n2796_lo_p;
  wire n2796_lo_n;
  wire n2799_lo_p;
  wire n2799_lo_n;
  wire n2802_lo_p;
  wire n2802_lo_n;
  wire n2805_lo_p;
  wire n2805_lo_n;
  wire n2808_lo_p;
  wire n2808_lo_n;
  wire n2820_lo_p;
  wire n2820_lo_n;
  wire n2823_lo_p;
  wire n2823_lo_n;
  wire n2826_lo_p;
  wire n2826_lo_n;
  wire n2829_lo_p;
  wire n2829_lo_n;
  wire n2832_lo_p;
  wire n2832_lo_n;
  wire n2835_lo_p;
  wire n2835_lo_n;
  wire n2838_lo_p;
  wire n2838_lo_n;
  wire n2841_lo_p;
  wire n2841_lo_n;
  wire n2844_lo_p;
  wire n2844_lo_n;
  wire n2856_lo_p;
  wire n2856_lo_n;
  wire n2859_lo_p;
  wire n2859_lo_n;
  wire n2862_lo_p;
  wire n2862_lo_n;
  wire n2865_lo_p;
  wire n2865_lo_n;
  wire n2868_lo_p;
  wire n2868_lo_n;
  wire n2871_lo_p;
  wire n2871_lo_n;
  wire n2874_lo_p;
  wire n2874_lo_n;
  wire n2877_lo_p;
  wire n2877_lo_n;
  wire n2880_lo_p;
  wire n2880_lo_n;
  wire n2883_lo_p;
  wire n2883_lo_n;
  wire n2886_lo_p;
  wire n2886_lo_n;
  wire n2889_lo_p;
  wire n2889_lo_n;
  wire n2892_lo_p;
  wire n2892_lo_n;
  wire n2895_lo_p;
  wire n2895_lo_n;
  wire n2898_lo_p;
  wire n2898_lo_n;
  wire n2901_lo_p;
  wire n2901_lo_n;
  wire n2904_lo_p;
  wire n2904_lo_n;
  wire n2907_lo_p;
  wire n2907_lo_n;
  wire n2916_lo_p;
  wire n2916_lo_n;
  wire n2919_lo_p;
  wire n2919_lo_n;
  wire n2925_lo_p;
  wire n2925_lo_n;
  wire n2928_lo_p;
  wire n2928_lo_n;
  wire n2940_lo_p;
  wire n2940_lo_n;
  wire n2943_lo_p;
  wire n2943_lo_n;
  wire n2952_lo_p;
  wire n2952_lo_n;
  wire n2955_lo_p;
  wire n2955_lo_n;
  wire n2961_lo_p;
  wire n2961_lo_n;
  wire n2964_lo_p;
  wire n2964_lo_n;
  wire n2967_lo_p;
  wire n2967_lo_n;
  wire n2970_lo_p;
  wire n2970_lo_n;
  wire n2976_lo_p;
  wire n2976_lo_n;
  wire n2979_lo_p;
  wire n2979_lo_n;
  wire n2982_lo_p;
  wire n2982_lo_n;
  wire n2988_lo_p;
  wire n2988_lo_n;
  wire n2991_lo_p;
  wire n2991_lo_n;
  wire n2994_lo_p;
  wire n2994_lo_n;
  wire n2997_lo_p;
  wire n2997_lo_n;
  wire n3000_lo_p;
  wire n3000_lo_n;
  wire n3003_lo_p;
  wire n3003_lo_n;
  wire n3006_lo_p;
  wire n3006_lo_n;
  wire n3012_lo_p;
  wire n3012_lo_n;
  wire n3015_lo_p;
  wire n3015_lo_n;
  wire n3018_lo_p;
  wire n3018_lo_n;
  wire n3021_lo_p;
  wire n3021_lo_n;
  wire n3024_lo_p;
  wire n3024_lo_n;
  wire n3027_lo_p;
  wire n3027_lo_n;
  wire n3030_lo_p;
  wire n3030_lo_n;
  wire n3033_lo_p;
  wire n3033_lo_n;
  wire n3036_lo_p;
  wire n3036_lo_n;
  wire n3039_lo_p;
  wire n3039_lo_n;
  wire n3045_lo_p;
  wire n3045_lo_n;
  wire n3048_lo_p;
  wire n3048_lo_n;
  wire n3051_lo_p;
  wire n3051_lo_n;
  wire n3054_lo_p;
  wire n3054_lo_n;
  wire n3057_lo_p;
  wire n3057_lo_n;
  wire n3060_lo_p;
  wire n3060_lo_n;
  wire n3063_lo_p;
  wire n3063_lo_n;
  wire n3069_lo_p;
  wire n3069_lo_n;
  wire n3072_lo_p;
  wire n3072_lo_n;
  wire n3075_lo_p;
  wire n3075_lo_n;
  wire n3081_lo_p;
  wire n3081_lo_n;
  wire n3084_lo_p;
  wire n3084_lo_n;
  wire n3087_lo_p;
  wire n3087_lo_n;
  wire n3093_lo_p;
  wire n3093_lo_n;
  wire n3096_lo_p;
  wire n3096_lo_n;
  wire n3099_lo_p;
  wire n3099_lo_n;
  wire n3102_lo_p;
  wire n3102_lo_n;
  wire n3105_lo_p;
  wire n3105_lo_n;
  wire n3108_lo_p;
  wire n3108_lo_n;
  wire n3111_lo_p;
  wire n3111_lo_n;
  wire n3114_lo_p;
  wire n3114_lo_n;
  wire n3117_lo_p;
  wire n3117_lo_n;
  wire n3120_lo_p;
  wire n3120_lo_n;
  wire n3123_lo_p;
  wire n3123_lo_n;
  wire n3126_lo_p;
  wire n3126_lo_n;
  wire n3129_lo_p;
  wire n3129_lo_n;
  wire n3132_lo_p;
  wire n3132_lo_n;
  wire n3135_lo_p;
  wire n3135_lo_n;
  wire n3138_lo_p;
  wire n3138_lo_n;
  wire n3141_lo_p;
  wire n3141_lo_n;
  wire n3156_lo_p;
  wire n3156_lo_n;
  wire n3168_lo_p;
  wire n3168_lo_n;
  wire n3171_lo_p;
  wire n3171_lo_n;
  wire n3174_lo_p;
  wire n3174_lo_n;
  wire n3177_lo_p;
  wire n3177_lo_n;
  wire n3180_lo_p;
  wire n3180_lo_n;
  wire n3183_lo_p;
  wire n3183_lo_n;
  wire n3192_lo_p;
  wire n3192_lo_n;
  wire n3195_lo_p;
  wire n3195_lo_n;
  wire n3204_lo_p;
  wire n3204_lo_n;
  wire n3207_lo_p;
  wire n3207_lo_n;
  wire n3210_lo_p;
  wire n3210_lo_n;
  wire n3216_lo_p;
  wire n3216_lo_n;
  wire n3219_lo_p;
  wire n3219_lo_n;
  wire n3222_lo_p;
  wire n3222_lo_n;
  wire n3228_lo_p;
  wire n3228_lo_n;
  wire n3231_lo_p;
  wire n3231_lo_n;
  wire n3240_lo_p;
  wire n3240_lo_n;
  wire n3243_lo_p;
  wire n3243_lo_n;
  wire n3252_lo_p;
  wire n3252_lo_n;
  wire n3255_lo_p;
  wire n3255_lo_n;
  wire n3258_lo_p;
  wire n3258_lo_n;
  wire n3264_lo_p;
  wire n3264_lo_n;
  wire n3267_lo_p;
  wire n3267_lo_n;
  wire n3270_lo_p;
  wire n3270_lo_n;
  wire n3276_lo_p;
  wire n3276_lo_n;
  wire n3279_lo_p;
  wire n3279_lo_n;
  wire n3282_lo_p;
  wire n3282_lo_n;
  wire n3288_lo_p;
  wire n3288_lo_n;
  wire n3291_lo_p;
  wire n3291_lo_n;
  wire n3294_lo_p;
  wire n3294_lo_n;
  wire n3603_o2_p;
  wire n3603_o2_n;
  wire n3604_o2_p;
  wire n3604_o2_n;
  wire n1391_inv_p;
  wire n1391_inv_n;
  wire n3798_o2_p;
  wire n3798_o2_n;
  wire n3846_o2_p;
  wire n3846_o2_n;
  wire n4019_o2_p;
  wire n4019_o2_n;
  wire n4017_o2_p;
  wire n4017_o2_n;
  wire n2177_o2_p;
  wire n2177_o2_n;
  wire n2150_o2_p;
  wire n2150_o2_n;
  wire n2154_o2_p;
  wire n2154_o2_n;
  wire n2184_o2_p;
  wire n2184_o2_n;
  wire n2515_o2_p;
  wire n2515_o2_n;
  wire n3837_o2_p;
  wire n3837_o2_n;
  wire n2167_o2_p;
  wire n2167_o2_n;
  wire n2118_o2_p;
  wire n2118_o2_n;
  wire n2186_o2_p;
  wire n2186_o2_n;
  wire n2174_o2_p;
  wire n2174_o2_n;
  wire n3964_o2_p;
  wire n3964_o2_n;
  wire n4005_o2_p;
  wire n4005_o2_n;
  wire n4006_o2_p;
  wire n4006_o2_n;
  wire n1445_inv_p;
  wire n1445_inv_n;
  wire n2176_o2_p;
  wire n2176_o2_n;
  wire n2227_o2_p;
  wire n2227_o2_n;
  wire n2236_o2_p;
  wire n2236_o2_n;
  wire n2245_o2_p;
  wire n2245_o2_n;
  wire n2518_o2_p;
  wire n2518_o2_n;
  wire n4023_o2_p;
  wire n4023_o2_n;
  wire n1466_inv_p;
  wire n1466_inv_n;
  wire n4038_o2_p;
  wire n4038_o2_n;
  wire n4039_o2_p;
  wire n4039_o2_n;
  wire n1475_inv_p;
  wire n1475_inv_n;
  wire n2119_o2_p;
  wire n2119_o2_n;
  wire n2275_o2_p;
  wire n2275_o2_n;
  wire n2595_o2_p;
  wire n2595_o2_n;
  wire n2594_o2_p;
  wire n2594_o2_n;
  wire lo498_buf_o2_p;
  wire lo498_buf_o2_n;
  wire lo502_buf_o2_p;
  wire lo502_buf_o2_n;
  wire lo550_buf_o2_p;
  wire lo550_buf_o2_n;
  wire n2596_o2_p;
  wire n2596_o2_n;
  wire n2593_o2_p;
  wire n2593_o2_n;
  wire n2668_o2_p;
  wire n2668_o2_n;
  wire lo542_buf_o2_p;
  wire lo542_buf_o2_n;
  wire n2667_o2_p;
  wire n2667_o2_n;
  wire n2404_o2_p;
  wire n2404_o2_n;
  wire n2410_o2_p;
  wire n2410_o2_n;
  wire n2419_o2_p;
  wire n2419_o2_n;
  wire n2392_o2_p;
  wire n2392_o2_n;
  wire n2369_o2_p;
  wire n2369_o2_n;
  wire n2397_o2_p;
  wire n2397_o2_n;
  wire n2601_o2_p;
  wire n2601_o2_n;
  wire n2658_o2_p;
  wire n2658_o2_n;
  wire n2574_o2_p;
  wire n2574_o2_n;
  wire n2205_o2_p;
  wire n2205_o2_n;
  wire lo510_buf_o2_p;
  wire lo510_buf_o2_n;
  wire lo514_buf_o2_p;
  wire lo514_buf_o2_n;
  wire lo554_buf_o2_p;
  wire lo554_buf_o2_n;
  wire lo558_buf_o2_p;
  wire lo558_buf_o2_n;
  wire lo578_buf_o2_p;
  wire lo578_buf_o2_n;
  wire n2254_o2_p;
  wire n2254_o2_n;
  wire n2421_o2_p;
  wire n2421_o2_n;
  wire n2422_o2_p;
  wire n2422_o2_n;
  wire n2130_o2_p;
  wire n2130_o2_n;
  wire n2127_o2_p;
  wire n2127_o2_n;
  wire n2131_o2_p;
  wire n2131_o2_n;
  wire n2128_o2_p;
  wire n2128_o2_n;
  wire n2264_o2_p;
  wire n2264_o2_n;
  wire n2467_o2_p;
  wire n2467_o2_n;
  wire n2471_o2_p;
  wire n2471_o2_n;
  wire n2488_o2_p;
  wire n2488_o2_n;
  wire n2478_o2_p;
  wire n2478_o2_n;
  wire n2486_o2_p;
  wire n2486_o2_n;
  wire n2485_o2_p;
  wire n2485_o2_n;
  wire n2498_o2_p;
  wire n2498_o2_n;
  wire n2495_o2_p;
  wire n2495_o2_n;
  wire n2496_o2_p;
  wire n2496_o2_n;
  wire n2458_o2_p;
  wire n2458_o2_n;
  wire n2643_o2_p;
  wire n2643_o2_n;
  wire n2462_o2_p;
  wire n2462_o2_n;
  wire n2468_o2_p;
  wire n2468_o2_n;
  wire n2639_o2_p;
  wire n2639_o2_n;
  wire n2499_o2_p;
  wire n2499_o2_n;
  wire n2472_o2_p;
  wire n2472_o2_n;
  wire n2474_o2_p;
  wire n2474_o2_n;
  wire n2489_o2_p;
  wire n2489_o2_n;
  wire n2321_o2_p;
  wire n2321_o2_n;
  wire n2322_o2_p;
  wire n2322_o2_n;
  wire n2640_o2_p;
  wire n2640_o2_n;
  wire n2642_o2_p;
  wire n2642_o2_n;
  wire n2187_o2_p;
  wire n2187_o2_n;
  wire n2373_o2_p;
  wire n2373_o2_n;
  wire n2603_o2_p;
  wire n2603_o2_n;
  wire n2388_o2_p;
  wire n2388_o2_n;
  wire n2437_o2_p;
  wire n2437_o2_n;
  wire n2356_o2_p;
  wire n2356_o2_n;
  wire n2452_o2_p;
  wire n2452_o2_n;
  wire n2347_o2_p;
  wire n2347_o2_n;
  wire n2329_o2_p;
  wire n2329_o2_n;
  wire n2669_o2_p;
  wire n2669_o2_n;
  wire n2332_o2_p;
  wire n2332_o2_n;
  wire n2664_o2_p;
  wire n2664_o2_n;
  wire n2665_o2_p;
  wire n2665_o2_n;
  wire n2653_o2_p;
  wire n2653_o2_n;
  wire n2654_o2_p;
  wire n2654_o2_n;
  wire n2636_o2_p;
  wire n2636_o2_n;
  wire n2660_o2_p;
  wire n2660_o2_n;
  wire n2318_o2_p;
  wire n2318_o2_n;
  wire n2319_o2_p;
  wire n2319_o2_n;
  wire n2586_o2_p;
  wire n2586_o2_n;
  wire n2587_o2_p;
  wire n2587_o2_n;
  wire n2288_o2_p;
  wire n2288_o2_n;
  wire n2344_o2_p;
  wire n2344_o2_n;
  wire n2530_o2_p;
  wire n2530_o2_n;
  wire n2303_o2_p;
  wire n2303_o2_n;
  wire n2566_o2_p;
  wire n2566_o2_n;
  wire n2567_o2_p;
  wire n2567_o2_n;
  wire n2554_o2_p;
  wire n2554_o2_n;
  wire n2194_o2_p;
  wire n2194_o2_n;
  wire lo582_buf_o2_p;
  wire lo582_buf_o2_n;
  wire lo030_buf_o2_p;
  wire lo030_buf_o2_n;
  wire lo174_buf_o2_p;
  wire lo174_buf_o2_n;
  wire lo178_buf_o2_p;
  wire lo178_buf_o2_n;
  wire lo186_buf_o2_p;
  wire lo186_buf_o2_n;
  wire lo266_buf_o2_p;
  wire lo266_buf_o2_n;
  wire lo306_buf_o2_p;
  wire lo306_buf_o2_n;
  wire lo346_buf_o2_p;
  wire lo346_buf_o2_n;
  wire lo386_buf_o2_p;
  wire lo386_buf_o2_n;
  wire lo426_buf_o2_p;
  wire lo426_buf_o2_n;
  wire lo590_buf_o2_p;
  wire lo590_buf_o2_n;
  wire lo594_buf_o2_p;
  wire lo594_buf_o2_n;
  wire lo606_buf_o2_p;
  wire lo606_buf_o2_n;
  wire lo610_buf_o2_p;
  wire lo610_buf_o2_n;
  wire n2238_o2_p;
  wire n2238_o2_n;
  wire n2229_o2_p;
  wire n2229_o2_n;
  wire n2242_o2_p;
  wire n2242_o2_n;
  wire n2233_o2_p;
  wire n2233_o2_n;
  wire n2168_o2_p;
  wire n2168_o2_n;
  wire n2237_o2_p;
  wire n2237_o2_n;
  wire n2228_o2_p;
  wire n2228_o2_n;
  wire n2172_o2_p;
  wire n2172_o2_n;
  wire n2223_o2_p;
  wire n2223_o2_n;
  wire n2222_o2_p;
  wire n2222_o2_n;
  wire n2170_o2_p;
  wire n2170_o2_n;
  wire n2181_o2_p;
  wire n2181_o2_n;
  wire n2510_o2_p;
  wire n2510_o2_n;
  wire n2621_o2_p;
  wire n2621_o2_n;
  wire lo466_buf_o2_p;
  wire lo466_buf_o2_n;
  wire lo478_buf_o2_p;
  wire lo478_buf_o2_n;
  wire n2149_o2_p;
  wire n2149_o2_n;
  wire n2429_o2_p;
  wire n2429_o2_n;
  wire n2444_o2_p;
  wire n2444_o2_n;
  wire n2153_o2_p;
  wire n2153_o2_n;
  wire n2433_o2_p;
  wire n2433_o2_n;
  wire n2448_o2_p;
  wire n2448_o2_n;
  wire n2367_o2_p;
  wire n2367_o2_n;
  wire n2386_o2_p;
  wire n2386_o2_n;
  wire n2539_o2_p;
  wire n2539_o2_n;
  wire n2183_o2_p;
  wire n2183_o2_n;
  wire n2220_o2_p;
  wire n2220_o2_n;
  wire n2514_o2_p;
  wire n2514_o2_n;
  wire n2196_o2_p;
  wire n2196_o2_n;
  wire n2616_o2_p;
  wire n2616_o2_n;
  wire n2612_o2_p;
  wire n2612_o2_n;
  wire n2627_o2_p;
  wire n2627_o2_n;
  wire n2140_o2_p;
  wire n2140_o2_n;
  wire n1877_inv_p;
  wire n1877_inv_n;
  wire lo149_buf_o2_p;
  wire lo149_buf_o2_n;
  wire lo197_buf_o2_p;
  wire lo197_buf_o2_n;
  wire lo118_buf_o2_p;
  wire lo118_buf_o2_n;
  wire lo158_buf_o2_p;
  wire lo158_buf_o2_n;
  wire lo166_buf_o2_p;
  wire lo166_buf_o2_n;
  wire lo242_buf_o2_p;
  wire lo242_buf_o2_n;
  wire lo286_buf_o2_p;
  wire lo286_buf_o2_n;
  wire lo506_buf_o2_p;
  wire lo506_buf_o2_n;
  wire n2198_o2_p;
  wire n2198_o2_n;
  wire n2202_o2_p;
  wire n2202_o2_n;
  wire n2197_o2_p;
  wire n2197_o2_n;
  wire n1913_inv_p;
  wire n1913_inv_n;
  wire n2146_o2_p;
  wire n2146_o2_n;
  wire n1919_inv_p;
  wire n1919_inv_n;
  wire lo312_buf_o2_p;
  wire lo312_buf_o2_n;
  wire lo316_buf_o2_p;
  wire lo316_buf_o2_n;
  wire lo352_buf_o2_p;
  wire lo352_buf_o2_n;
  wire lo356_buf_o2_p;
  wire lo356_buf_o2_n;
  wire lo392_buf_o2_p;
  wire lo392_buf_o2_n;
  wire lo396_buf_o2_p;
  wire lo396_buf_o2_n;
  wire lo432_buf_o2_p;
  wire lo432_buf_o2_n;
  wire lo436_buf_o2_p;
  wire lo436_buf_o2_n;
  wire lo576_buf_o2_p;
  wire lo576_buf_o2_n;
  wire g733_p;
  wire g733_n;
  wire g734_p;
  wire g734_n;
  wire g735_p;
  wire g735_n;
  wire g736_p;
  wire g736_n;
  wire g737_p;
  wire g737_n;
  wire g738_p;
  wire g738_n;
  wire g739_p;
  wire g739_n;
  wire g740_p;
  wire g740_n;
  wire g741_p;
  wire g741_n;
  wire g742_p;
  wire g742_n;
  wire g743_p;
  wire g743_n;
  wire g744_p;
  wire g744_n;
  wire g745_p;
  wire g745_n;
  wire g746_p;
  wire g746_n;
  wire g747_p;
  wire g747_n;
  wire g748_p;
  wire g748_n;
  wire g749_p;
  wire g749_n;
  wire g750_p;
  wire g750_n;
  wire g751_p;
  wire g751_n;
  wire g752_p;
  wire g752_n;
  wire g753_p;
  wire g753_n;
  wire g754_p;
  wire g754_n;
  wire g755_p;
  wire g755_n;
  wire g756_p;
  wire g756_n;
  wire g757_p;
  wire g757_n;
  wire g758_p;
  wire g758_n;
  wire g759_p;
  wire g759_n;
  wire g760_p;
  wire g760_n;
  wire g761_p;
  wire g761_n;
  wire g762_p;
  wire g762_n;
  wire g763_p;
  wire g763_n;
  wire g764_p;
  wire g764_n;
  wire g765_p;
  wire g765_n;
  wire g766_p;
  wire g766_n;
  wire g767_p;
  wire g767_n;
  wire g768_p;
  wire g768_n;
  wire g769_p;
  wire g769_n;
  wire g770_p;
  wire g770_n;
  wire g771_p;
  wire g771_n;
  wire g772_p;
  wire g772_n;
  wire g773_p;
  wire g773_n;
  wire g774_p;
  wire g774_n;
  wire g775_p;
  wire g775_n;
  wire g776_p;
  wire g776_n;
  wire g777_p;
  wire g777_n;
  wire g778_p;
  wire g778_n;
  wire g779_p;
  wire g779_n;
  wire g780_p;
  wire g780_n;
  wire g781_p;
  wire g781_n;
  wire g782_p;
  wire g782_n;
  wire g783_p;
  wire g783_n;
  wire g784_p;
  wire g784_n;
  wire g785_p;
  wire g785_n;
  wire g786_p;
  wire g786_n;
  wire g787_p;
  wire g787_n;
  wire g788_p;
  wire g788_n;
  wire g789_p;
  wire g789_n;
  wire g790_p;
  wire g790_n;
  wire g791_p;
  wire g791_n;
  wire g792_p;
  wire g792_n;
  wire g793_p;
  wire g793_n;
  wire g794_p;
  wire g794_n;
  wire g795_p;
  wire g795_n;
  wire g796_p;
  wire g796_n;
  wire g797_p;
  wire g797_n;
  wire g798_p;
  wire g798_n;
  wire g799_p;
  wire g799_n;
  wire g800_p;
  wire g800_n;
  wire g801_p;
  wire g801_n;
  wire g802_p;
  wire g802_n;
  wire g803_p;
  wire g803_n;
  wire g804_p;
  wire g804_n;
  wire g805_p;
  wire g805_n;
  wire g806_p;
  wire g806_n;
  wire g807_p;
  wire g807_n;
  wire g808_p;
  wire g808_n;
  wire g809_p;
  wire g809_n;
  wire g810_p;
  wire g810_n;
  wire g811_p;
  wire g811_n;
  wire g812_p;
  wire g812_n;
  wire g813_p;
  wire g813_n;
  wire g814_p;
  wire g814_n;
  wire g815_p;
  wire g815_n;
  wire g816_p;
  wire g816_n;
  wire g817_p;
  wire g817_n;
  wire g818_p;
  wire g818_n;
  wire g819_p;
  wire g819_n;
  wire g820_p;
  wire g820_n;
  wire g821_p;
  wire g821_n;
  wire g822_p;
  wire g822_n;
  wire g823_p;
  wire g823_n;
  wire g824_p;
  wire g824_n;
  wire g825_p;
  wire g825_n;
  wire g826_p;
  wire g826_n;
  wire g827_p;
  wire g827_n;
  wire g828_p;
  wire g828_n;
  wire g829_p;
  wire g829_n;
  wire g830_p;
  wire g830_n;
  wire g831_p;
  wire g831_n;
  wire g832_p;
  wire g832_n;
  wire g833_p;
  wire g833_n;
  wire g834_p;
  wire g834_n;
  wire g835_p;
  wire g835_n;
  wire g836_p;
  wire g836_n;
  wire g837_p;
  wire g837_n;
  wire g838_p;
  wire g838_n;
  wire g839_p;
  wire g839_n;
  wire g840_p;
  wire g840_n;
  wire g841_p;
  wire g841_n;
  wire g842_p;
  wire g842_n;
  wire g843_p;
  wire g843_n;
  wire g844_p;
  wire g844_n;
  wire g845_p;
  wire g845_n;
  wire g846_p;
  wire g846_n;
  wire g847_p;
  wire g847_n;
  wire g848_p;
  wire g848_n;
  wire g849_p;
  wire g849_n;
  wire g850_p;
  wire g850_n;
  wire g851_p;
  wire g851_n;
  wire g852_p;
  wire g852_n;
  wire g853_p;
  wire g853_n;
  wire g854_p;
  wire g854_n;
  wire g855_p;
  wire g855_n;
  wire g856_p;
  wire g856_n;
  wire g857_p;
  wire g857_n;
  wire g858_p;
  wire g858_n;
  wire g859_p;
  wire g859_n;
  wire g860_p;
  wire g860_n;
  wire g861_p;
  wire g861_n;
  wire g862_p;
  wire g862_n;
  wire g863_p;
  wire g863_n;
  wire g864_p;
  wire g864_n;
  wire g865_p;
  wire g865_n;
  wire g866_p;
  wire g866_n;
  wire g867_p;
  wire g867_n;
  wire g868_p;
  wire g868_n;
  wire g869_p;
  wire g869_n;
  wire g870_p;
  wire g870_n;
  wire g871_p;
  wire g871_n;
  wire g872_p;
  wire g872_n;
  wire g873_p;
  wire g873_n;
  wire g874_p;
  wire g874_n;
  wire g875_p;
  wire g875_n;
  wire g876_p;
  wire g876_n;
  wire g877_p;
  wire g877_n;
  wire g878_p;
  wire g878_n;
  wire g879_p;
  wire g879_n;
  wire g880_p;
  wire g880_n;
  wire g881_p;
  wire g881_n;
  wire g882_p;
  wire g882_n;
  wire g883_p;
  wire g883_n;
  wire g884_p;
  wire g884_n;
  wire g885_p;
  wire g885_n;
  wire g886_p;
  wire g886_n;
  wire g887_p;
  wire g887_n;
  wire g888_p;
  wire g888_n;
  wire g889_p;
  wire g889_n;
  wire g890_p;
  wire g890_n;
  wire g891_p;
  wire g891_n;
  wire g892_p;
  wire g892_n;
  wire g893_p;
  wire g893_n;
  wire g894_p;
  wire g894_n;
  wire g895_p;
  wire g895_n;
  wire g896_p;
  wire g896_n;
  wire g897_p;
  wire g897_n;
  wire g898_p;
  wire g898_n;
  wire g899_p;
  wire g899_n;
  wire g900_p;
  wire g900_n;
  wire g901_p;
  wire g901_n;
  wire g902_p;
  wire g902_n;
  wire g903_p;
  wire g903_n;
  wire g904_p;
  wire g904_n;
  wire g905_p;
  wire g905_n;
  wire g906_p;
  wire g906_n;
  wire g907_p;
  wire g907_n;
  wire g908_p;
  wire g908_n;
  wire g909_p;
  wire g909_n;
  wire g910_p;
  wire g910_n;
  wire g911_p;
  wire g911_n;
  wire g912_p;
  wire g912_n;
  wire g913_p;
  wire g913_n;
  wire g914_p;
  wire g914_n;
  wire g915_p;
  wire g915_n;
  wire g916_p;
  wire g916_n;
  wire g917_p;
  wire g917_n;
  wire g918_p;
  wire g918_n;
  wire g919_p;
  wire g919_n;
  wire g920_p;
  wire g920_n;
  wire g921_p;
  wire g921_n;
  wire g922_p;
  wire g922_n;
  wire g923_p;
  wire g923_n;
  wire g924_p;
  wire g924_n;
  wire g925_p;
  wire g925_n;
  wire g926_p;
  wire g926_n;
  wire g927_p;
  wire g927_n;
  wire g928_p;
  wire g928_n;
  wire g929_p;
  wire g929_n;
  wire g930_p;
  wire g930_n;
  wire g931_p;
  wire g931_n;
  wire g932_p;
  wire g932_n;
  wire g933_p;
  wire g933_n;
  wire g934_p;
  wire g934_n;
  wire g935_p;
  wire g935_n;
  wire g936_p;
  wire g936_n;
  wire g937_p;
  wire g937_n;
  wire g938_p;
  wire g938_n;
  wire g939_p;
  wire g939_n;
  wire g940_p;
  wire g940_n;
  wire g941_p;
  wire g941_n;
  wire g942_p;
  wire g942_n;
  wire g943_p;
  wire g943_n;
  wire g944_p;
  wire g944_n;
  wire g945_p;
  wire g945_n;
  wire g946_p;
  wire g946_n;
  wire g947_p;
  wire g947_n;
  wire g948_p;
  wire g948_n;
  wire g949_p;
  wire g949_n;
  wire g950_p;
  wire g950_n;
  wire g951_p;
  wire g951_n;
  wire g952_p;
  wire g952_n;
  wire g953_p;
  wire g953_n;
  wire g954_p;
  wire g954_n;
  wire g955_p;
  wire g955_n;
  wire g956_p;
  wire g956_n;
  wire g957_p;
  wire g957_n;
  wire g958_p;
  wire g958_n;
  wire g959_p;
  wire g959_n;
  wire g960_p;
  wire g960_n;
  wire g961_p;
  wire g961_n;
  wire g962_p;
  wire g962_n;
  wire g963_p;
  wire g963_n;
  wire g964_p;
  wire g964_n;
  wire g965_p;
  wire g965_n;
  wire g966_p;
  wire g966_n;
  wire g967_p;
  wire g967_n;
  wire g968_p;
  wire g968_n;
  wire g969_p;
  wire g969_n;
  wire g970_p;
  wire g970_n;
  wire g971_p;
  wire g971_n;
  wire g972_p;
  wire g972_n;
  wire g973_p;
  wire g973_n;
  wire g974_p;
  wire g974_n;
  wire g975_p;
  wire g975_n;
  wire g976_p;
  wire g976_n;
  wire g977_p;
  wire g977_n;
  wire g978_p;
  wire g978_n;
  wire g979_p;
  wire g979_n;
  wire g980_p;
  wire g980_n;
  wire g981_p;
  wire g981_n;
  wire g982_p;
  wire g982_n;
  wire g983_p;
  wire g983_n;
  wire g984_p;
  wire g984_n;
  wire g985_p;
  wire g985_n;
  wire g986_p;
  wire g986_n;
  wire g987_p;
  wire g987_n;
  wire g988_p;
  wire g988_n;
  wire g989_p;
  wire g989_n;
  wire g990_p;
  wire g990_n;
  wire g991_p;
  wire g991_n;
  wire g992_p;
  wire g992_n;
  wire g993_p;
  wire g993_n;
  wire g994_p;
  wire g994_n;
  wire g995_p;
  wire g995_n;
  wire g996_p;
  wire g996_n;
  wire g997_p;
  wire g997_n;
  wire g998_p;
  wire g998_n;
  wire g999_p;
  wire g999_n;
  wire g1000_p;
  wire g1000_n;
  wire g1001_p;
  wire g1001_n;
  wire g1002_p;
  wire g1002_n;
  wire g1003_p;
  wire g1003_n;
  wire g1004_p;
  wire g1004_n;
  wire g1005_p;
  wire g1005_n;
  wire g1006_p;
  wire g1006_n;
  wire g1007_p;
  wire g1007_n;
  wire g1008_p;
  wire g1008_n;
  wire g1009_p;
  wire g1009_n;
  wire g1010_p;
  wire g1010_n;
  wire g1011_p;
  wire g1011_n;
  wire g1012_p;
  wire g1012_n;
  wire g1013_p;
  wire g1013_n;
  wire g1014_p;
  wire g1014_n;
  wire g1015_p;
  wire g1015_n;
  wire g1016_p;
  wire g1016_n;
  wire g1017_p;
  wire g1017_n;
  wire g1018_p;
  wire g1018_n;
  wire g1019_p;
  wire g1019_n;
  wire g1020_p;
  wire g1020_n;
  wire g1021_p;
  wire g1021_n;
  wire g1022_p;
  wire g1022_n;
  wire g1023_p;
  wire g1023_n;
  wire g1024_p;
  wire g1024_n;
  wire g1025_p;
  wire g1025_n;
  wire g1026_p;
  wire g1026_n;
  wire g1027_p;
  wire g1027_n;
  wire g1028_p;
  wire g1028_n;
  wire g1029_p;
  wire g1029_n;
  wire g1030_p;
  wire g1030_n;
  wire g1031_p;
  wire g1031_n;
  wire g1032_p;
  wire g1032_n;
  wire g1033_p;
  wire g1033_n;
  wire g1034_p;
  wire g1034_n;
  wire g1035_p;
  wire g1035_n;
  wire g1036_p;
  wire g1036_n;
  wire g1037_p;
  wire g1037_n;
  wire g1038_p;
  wire g1038_n;
  wire g1039_p;
  wire g1039_n;
  wire g1040_p;
  wire g1040_n;
  wire g1041_p;
  wire g1041_n;
  wire g1042_p;
  wire g1042_n;
  wire g1043_p;
  wire g1043_n;
  wire g1044_p;
  wire g1044_n;
  wire g1045_p;
  wire g1045_n;
  wire g1046_p;
  wire g1046_n;
  wire g1047_p;
  wire g1047_n;
  wire g1048_p;
  wire g1048_n;
  wire g1049_p;
  wire g1049_n;
  wire g1050_p;
  wire g1050_n;
  wire g1051_p;
  wire g1051_n;
  wire g1052_p;
  wire g1052_n;
  wire g1053_p;
  wire g1053_n;
  wire g1054_p;
  wire g1054_n;
  wire g1055_p;
  wire g1055_n;
  wire g1056_p;
  wire g1056_n;
  wire g1057_p;
  wire g1057_n;
  wire g1058_p;
  wire g1058_n;
  wire g1059_p;
  wire g1059_n;
  wire g1060_p;
  wire g1060_n;
  wire g1061_p;
  wire g1061_n;
  wire g1062_p;
  wire g1062_n;
  wire g1063_p;
  wire g1063_n;
  wire g1064_p;
  wire g1064_n;
  wire g1065_p;
  wire g1065_n;
  wire g1066_p;
  wire g1066_n;
  wire g1067_p;
  wire g1067_n;
  wire g1068_p;
  wire g1068_n;
  wire g1069_p;
  wire g1069_n;
  wire g1070_p;
  wire g1070_n;
  wire g1071_p;
  wire g1071_n;
  wire g1072_p;
  wire g1072_n;
  wire g1073_p;
  wire g1073_n;
  wire g1074_p;
  wire g1074_n;
  wire g1075_p;
  wire g1075_n;
  wire g1076_p;
  wire g1076_n;
  wire g1077_p;
  wire g1077_n;
  wire g1078_p;
  wire g1078_n;
  wire g1079_p;
  wire g1079_n;
  wire g1080_p;
  wire g1080_n;
  wire g1081_p;
  wire g1081_n;
  wire g1082_p;
  wire g1082_n;
  wire g1083_p;
  wire g1083_n;
  wire g1084_p;
  wire g1084_n;
  wire g1085_p;
  wire g1085_n;
  wire g1086_p;
  wire g1086_n;
  wire g1087_p;
  wire g1087_n;
  wire g1088_p;
  wire g1088_n;
  wire g1089_p;
  wire g1089_n;
  wire g1090_p;
  wire g1090_n;
  wire g1091_p;
  wire g1091_n;
  wire g1092_p;
  wire g1092_n;
  wire g1093_p;
  wire g1093_n;
  wire g1094_p;
  wire g1094_n;
  wire g1095_p;
  wire g1095_n;
  wire g1096_p;
  wire g1096_n;
  wire g1097_p;
  wire g1097_n;
  wire g1098_p;
  wire g1098_n;
  wire g1099_p;
  wire g1099_n;
  wire g1100_p;
  wire g1100_n;
  wire g1101_p;
  wire g1101_n;
  wire g1102_p;
  wire g1102_n;
  wire g1103_p;
  wire g1103_n;
  wire g1104_p;
  wire g1104_n;
  wire g1105_p;
  wire g1105_n;
  wire g1106_p;
  wire g1106_n;
  wire g1107_p;
  wire g1107_n;
  wire g1108_p;
  wire g1108_n;
  wire g1109_p;
  wire g1109_n;
  wire g1110_p;
  wire g1110_n;
  wire g1111_p;
  wire g1111_n;
  wire g1112_p;
  wire g1112_n;
  wire g1113_p;
  wire g1113_n;
  wire g1114_p;
  wire g1114_n;
  wire g1115_p;
  wire g1115_n;
  wire g1116_p;
  wire g1116_n;
  wire g1117_p;
  wire g1117_n;
  wire g1118_p;
  wire g1118_n;
  wire g1119_p;
  wire g1119_n;
  wire g1120_p;
  wire g1120_n;
  wire g1121_p;
  wire g1121_n;
  wire g1122_p;
  wire g1122_n;
  wire g1123_p;
  wire g1123_n;
  wire g1124_p;
  wire g1124_n;
  wire g1125_p;
  wire g1125_n;
  wire g1126_p;
  wire g1126_n;
  wire g1127_p;
  wire g1127_n;
  wire g1128_p;
  wire g1128_n;
  wire g1129_p;
  wire g1129_n;
  wire g1130_p;
  wire g1130_n;
  wire g1131_p;
  wire g1131_n;
  wire g1132_p;
  wire g1132_n;
  wire g1133_p;
  wire g1133_n;
  wire g1134_p;
  wire g1134_n;
  wire g1135_p;
  wire g1135_n;
  wire g1136_p;
  wire g1136_n;
  wire g1137_p;
  wire g1137_n;
  wire g1138_p;
  wire g1138_n;
  wire g1139_p;
  wire g1139_n;
  wire g1140_p;
  wire g1140_n;
  wire g1141_p;
  wire g1141_n;
  wire g1142_p;
  wire g1142_n;
  wire g1143_p;
  wire g1143_n;
  wire g1144_p;
  wire g1144_n;
  wire g1145_p;
  wire g1145_n;
  wire g1146_p;
  wire g1146_n;
  wire g1147_p;
  wire g1147_n;
  wire g1148_p;
  wire g1148_n;
  wire g1149_p;
  wire g1149_n;
  wire g1150_p;
  wire g1150_n;
  wire g1151_p;
  wire g1151_n;
  wire g1152_p;
  wire g1152_n;
  wire g1153_p;
  wire g1153_n;
  wire g1154_p;
  wire g1154_n;
  wire g1155_p;
  wire g1155_n;
  wire g1156_p;
  wire g1156_n;
  wire g1157_p;
  wire g1157_n;
  wire g1158_p;
  wire g1158_n;
  wire g1159_p;
  wire g1159_n;
  wire g1160_p;
  wire g1160_n;
  wire g1161_p;
  wire g1161_n;
  wire g1162_p;
  wire g1162_n;
  wire g1163_p;
  wire g1163_n;
  wire g1164_p;
  wire g1164_n;
  wire g1165_p;
  wire g1165_n;
  wire g1166_p;
  wire g1166_n;
  wire g1167_p;
  wire g1167_n;
  wire g1168_p;
  wire g1168_n;
  wire g1169_p;
  wire g1169_n;
  wire g1170_p;
  wire g1170_n;
  wire g1171_p;
  wire g1171_n;
  wire g1172_p;
  wire g1172_n;
  wire g1173_p;
  wire g1173_n;
  wire g1174_p;
  wire g1174_n;
  wire g1175_p;
  wire g1175_n;
  wire g1176_p;
  wire g1176_n;
  wire g1177_p;
  wire g1177_n;
  wire g1178_p;
  wire g1178_n;
  wire g1179_p;
  wire g1179_n;
  wire g1180_p;
  wire g1180_n;
  wire g1181_p;
  wire g1181_n;
  wire g1182_p;
  wire g1182_n;
  wire g1183_p;
  wire g1183_n;
  wire g1184_p;
  wire g1184_n;
  wire g1185_p;
  wire g1185_n;
  wire g1186_p;
  wire g1186_n;
  wire g1187_p;
  wire g1187_n;
  wire g1188_p;
  wire g1188_n;
  wire g1189_p;
  wire g1189_n;
  wire g1190_p;
  wire g1190_n;
  wire g1191_p;
  wire g1191_n;
  wire g1192_p;
  wire g1192_n;
  wire g1193_p;
  wire g1193_n;
  wire g1194_p;
  wire g1194_n;
  wire g1195_p;
  wire g1195_n;
  wire g1196_p;
  wire g1196_n;
  wire g1197_p;
  wire g1197_n;
  wire g1198_p;
  wire g1198_n;
  wire g1199_p;
  wire g1199_n;
  wire g1200_p;
  wire g1200_n;
  wire g1201_p;
  wire g1201_n;
  wire g1202_p;
  wire g1202_n;
  wire g1203_p;
  wire g1203_n;
  wire g1204_p;
  wire g1204_n;
  wire g1205_p;
  wire g1205_n;
  wire g1206_p;
  wire g1206_n;
  wire g1207_p;
  wire g1207_n;
  wire g1208_p;
  wire g1208_n;
  wire g1209_p;
  wire g1209_n;
  wire g1210_p;
  wire g1210_n;
  wire g1211_p;
  wire g1211_n;
  wire g1212_p;
  wire g1212_n;
  wire g1213_p;
  wire g1213_n;
  wire g1214_p;
  wire g1214_n;
  wire g1215_p;
  wire g1215_n;
  wire g1216_p;
  wire g1216_n;
  wire g1217_p;
  wire g1217_n;
  wire g1218_p;
  wire g1218_n;
  wire g1219_p;
  wire g1219_n;
  wire g1220_p;
  wire g1220_n;
  wire g1221_p;
  wire g1221_n;
  wire g1222_p;
  wire g1222_n;
  wire g1223_p;
  wire g1223_n;
  wire g1224_p;
  wire g1224_n;
  wire g1225_p;
  wire g1225_n;
  wire g1226_p;
  wire g1226_n;
  wire g1227_p;
  wire g1227_n;
  wire g1228_p;
  wire g1228_n;
  wire g1229_p;
  wire g1229_n;
  wire g1230_p;
  wire g1230_n;
  wire g1231_p;
  wire g1231_n;
  wire g1232_p;
  wire g1232_n;
  wire g1233_p;
  wire g1233_n;
  wire g1234_p;
  wire g1234_n;
  wire g1235_p;
  wire g1235_n;
  wire g1236_p;
  wire g1236_n;
  wire g1237_p;
  wire g1237_n;
  wire g1238_p;
  wire g1238_n;
  wire g1239_p;
  wire g1239_n;
  wire g1240_p;
  wire g1240_n;
  wire g1241_p;
  wire g1241_n;
  wire g1242_p;
  wire g1242_n;
  wire g1243_p;
  wire g1243_n;
  wire g1244_p;
  wire g1244_n;
  wire g1245_p;
  wire g1245_n;
  wire g1246_p;
  wire g1246_n;
  wire g1247_p;
  wire g1247_n;
  wire g1248_p;
  wire g1248_n;
  wire g1249_p;
  wire g1249_n;
  wire g1250_p;
  wire g1250_n;
  wire g1251_p;
  wire g1251_n;
  wire g1252_p;
  wire g1252_n;
  wire g1253_p;
  wire g1253_n;
  wire g1254_p;
  wire g1254_n;
  wire g1255_p;
  wire g1255_n;
  wire g1256_p;
  wire g1256_n;
  wire g1257_p;
  wire g1257_n;
  wire g1258_p;
  wire g1258_n;
  wire g1259_p;
  wire g1259_n;
  wire g1260_p;
  wire g1260_n;
  wire g1261_p;
  wire g1261_n;
  wire g1262_p;
  wire g1262_n;
  wire g1263_p;
  wire g1263_n;
  wire g1264_p;
  wire g1264_n;
  wire g1265_p;
  wire g1265_n;
  wire g1266_p;
  wire g1266_n;
  wire g1267_p;
  wire g1267_n;
  wire g1268_p;
  wire g1268_n;
  wire g1269_p;
  wire g1269_n;
  wire g1270_p;
  wire g1270_n;
  wire g1271_p;
  wire g1271_n;
  wire g1272_p;
  wire g1272_n;
  wire g1273_p;
  wire g1273_n;
  wire g1274_p;
  wire g1274_n;
  wire g1275_p;
  wire g1275_n;
  wire g1276_p;
  wire g1276_n;
  wire g1277_p;
  wire g1277_n;
  wire g1278_p;
  wire g1278_n;
  wire g1279_p;
  wire g1279_n;
  wire g1280_p;
  wire g1280_n;
  wire g1281_p;
  wire g1281_n;
  wire g1282_p;
  wire g1282_n;
  wire g1283_p;
  wire g1283_n;
  wire g1284_p;
  wire g1284_n;
  wire g1285_p;
  wire g1285_n;
  wire g1286_p;
  wire g1286_n;
  wire g1287_p;
  wire g1287_n;
  wire g1288_p;
  wire g1288_n;
  wire g1289_p;
  wire g1289_n;
  wire g1290_p;
  wire g1290_n;
  wire g1291_p;
  wire g1291_n;
  wire g1292_p;
  wire g1292_n;
  wire g1293_p;
  wire g1293_n;
  wire g1294_p;
  wire g1294_n;
  wire g1295_p;
  wire g1295_n;
  wire g1296_p;
  wire g1296_n;
  wire g1297_p;
  wire g1297_n;
  wire g1298_p;
  wire g1298_n;
  wire g1299_p;
  wire g1299_n;
  wire g1300_p;
  wire g1300_n;
  wire g1301_p;
  wire g1301_n;
  wire g1302_p;
  wire g1302_n;
  wire n2865_lo_n_spl_;
  wire n2793_lo_n_spl_;
  wire n2793_lo_n_spl_0;
  wire n2793_lo_n_spl_1;
  wire g737_n_spl_;
  wire g737_n_spl_0;
  wire g740_n_spl_;
  wire g741_n_spl_;
  wire n2877_lo_n_spl_;
  wire n2877_lo_n_spl_0;
  wire g745_n_spl_;
  wire g745_n_spl_0;
  wire g752_n_spl_;
  wire n2889_lo_p_spl_;
  wire n2889_lo_p_spl_0;
  wire n2889_lo_p_spl_1;
  wire n3846_o2_n_spl_;
  wire n2889_lo_n_spl_;
  wire n2889_lo_n_spl_0;
  wire n2889_lo_n_spl_1;
  wire n4019_o2_p_spl_;
  wire g749_n_spl_;
  wire n2829_lo_p_spl_;
  wire n3846_o2_p_spl_;
  wire n2264_o2_n_spl_;
  wire n2264_o2_n_spl_0;
  wire n2329_o2_p_spl_;
  wire n2332_o2_n_spl_;
  wire n2329_o2_n_spl_;
  wire n2332_o2_p_spl_;
  wire n2347_o2_n_spl_;
  wire n2344_o2_p_spl_;
  wire n2347_o2_p_spl_;
  wire n2344_o2_n_spl_;
  wire n2515_o2_p_spl_;
  wire n1761_lo_n_spl_;
  wire n2574_o2_n_spl_;
  wire n2264_o2_p_spl_;
  wire n2574_o2_p_spl_;
  wire g851_p_spl_;
  wire g851_n_spl_;
  wire g868_n_spl_;
  wire n2660_o2_p_spl_;
  wire g875_n_spl_;
  wire g877_n_spl_;
  wire g876_n_spl_;
  wire g774_p_spl_;
  wire g779_p_spl_;
  wire g788_p_spl_;
  wire g849_p_spl_;
  wire g864_p_spl_;
  wire n4038_o2_p_spl_;
  wire n4038_o2_p_spl_0;
  wire n4038_o2_p_spl_1;
  wire n4038_o2_n_spl_;
  wire n4038_o2_n_spl_0;
  wire n4038_o2_n_spl_1;
  wire n3964_o2_p_spl_;
  wire n3964_o2_p_spl_0;
  wire n3964_o2_p_spl_00;
  wire n3964_o2_p_spl_01;
  wire n3964_o2_p_spl_1;
  wire n3964_o2_p_spl_10;
  wire n3964_o2_p_spl_11;
  wire n3964_o2_n_spl_;
  wire n3964_o2_n_spl_0;
  wire n3964_o2_n_spl_00;
  wire n3964_o2_n_spl_01;
  wire n3964_o2_n_spl_1;
  wire n3964_o2_n_spl_10;
  wire n3964_o2_n_spl_11;
  wire lo554_buf_o2_p_spl_;
  wire lo554_buf_o2_p_spl_0;
  wire lo558_buf_o2_p_spl_;
  wire lo558_buf_o2_p_spl_0;
  wire lo554_buf_o2_n_spl_;
  wire lo554_buf_o2_n_spl_0;
  wire lo558_buf_o2_n_spl_;
  wire lo558_buf_o2_n_spl_0;
  wire g896_p_spl_;
  wire g899_p_spl_;
  wire n4006_o2_n_spl_;
  wire n4006_o2_n_spl_0;
  wire n4006_o2_n_spl_00;
  wire n4006_o2_n_spl_01;
  wire n4006_o2_n_spl_1;
  wire n4006_o2_p_spl_;
  wire n4006_o2_p_spl_0;
  wire n4006_o2_p_spl_00;
  wire n4006_o2_p_spl_01;
  wire n4006_o2_p_spl_1;
  wire g901_p_spl_;
  wire g906_p_spl_;
  wire n4005_o2_n_spl_;
  wire n4005_o2_p_spl_;
  wire n2205_o2_n_spl_;
  wire g900_n_spl_;
  wire g900_n_spl_0;
  wire n2205_o2_p_spl_;
  wire n2205_o2_p_spl_0;
  wire n2205_o2_p_spl_1;
  wire g900_p_spl_;
  wire n3102_lo_n_spl_;
  wire n3102_lo_n_spl_0;
  wire n3114_lo_n_spl_;
  wire n3837_o2_n_spl_;
  wire n3837_o2_n_spl_0;
  wire n3837_o2_n_spl_1;
  wire n3837_o2_p_spl_;
  wire n3837_o2_p_spl_0;
  wire n3837_o2_p_spl_1;
  wire n2146_o2_p_spl_;
  wire n1919_inv_p_spl_;
  wire g939_p_spl_;
  wire g940_p_spl_;
  wire lo030_buf_o2_n_spl_;
  wire g908_n_spl_;
  wire g908_n_spl_0;
  wire g908_n_spl_1;
  wire n3018_lo_p_spl_;
  wire n3018_lo_p_spl_0;
  wire g943_n_spl_;
  wire g943_n_spl_0;
  wire g943_n_spl_00;
  wire g943_n_spl_1;
  wire g925_p_spl_;
  wire g943_p_spl_;
  wire g943_p_spl_0;
  wire g943_p_spl_00;
  wire g943_p_spl_1;
  wire n1554_lo_p_spl_;
  wire n1554_lo_p_spl_0;
  wire n1554_lo_p_spl_00;
  wire n1554_lo_p_spl_000;
  wire n1554_lo_p_spl_01;
  wire n1554_lo_p_spl_1;
  wire n1554_lo_p_spl_10;
  wire n1554_lo_p_spl_11;
  wire n1554_lo_n_spl_;
  wire n1554_lo_n_spl_0;
  wire n1554_lo_n_spl_00;
  wire n1554_lo_n_spl_000;
  wire n1554_lo_n_spl_01;
  wire n1554_lo_n_spl_1;
  wire n1554_lo_n_spl_10;
  wire n1554_lo_n_spl_11;
  wire n2254_o2_p_spl_;
  wire n2254_o2_p_spl_0;
  wire n2254_o2_p_spl_00;
  wire n2254_o2_p_spl_1;
  wire g925_n_spl_;
  wire g925_n_spl_0;
  wire g913_p_spl_;
  wire g913_p_spl_0;
  wire n1686_lo_p_spl_;
  wire n1686_lo_p_spl_0;
  wire n1686_lo_p_spl_00;
  wire n1686_lo_p_spl_01;
  wire n1686_lo_p_spl_1;
  wire n1686_lo_p_spl_10;
  wire n1686_lo_p_spl_11;
  wire n1686_lo_n_spl_;
  wire n1686_lo_n_spl_0;
  wire n1686_lo_n_spl_00;
  wire n1686_lo_n_spl_01;
  wire n1686_lo_n_spl_1;
  wire n1686_lo_n_spl_10;
  wire n1686_lo_n_spl_11;
  wire n1475_inv_p_spl_;
  wire n1475_inv_p_spl_0;
  wire n1475_inv_p_spl_1;
  wire n2367_o2_p_spl_;
  wire n2367_o2_p_spl_0;
  wire n4039_o2_p_spl_;
  wire n4039_o2_p_spl_0;
  wire lo030_buf_o2_p_spl_;
  wire n2982_lo_n_spl_;
  wire n2982_lo_n_spl_0;
  wire n2982_lo_n_spl_00;
  wire n2982_lo_n_spl_1;
  wire g964_p_spl_;
  wire g964_p_spl_0;
  wire g964_p_spl_1;
  wire g966_p_spl_;
  wire g966_p_spl_0;
  wire g966_p_spl_1;
  wire g971_n_spl_;
  wire g971_n_spl_0;
  wire g971_n_spl_1;
  wire g971_p_spl_;
  wire g971_p_spl_0;
  wire lo542_buf_o2_n_spl_;
  wire lo542_buf_o2_p_spl_;
  wire lo542_buf_o2_p_spl_0;
  wire n2220_o2_p_spl_;
  wire n2220_o2_p_spl_0;
  wire n2220_o2_p_spl_00;
  wire n2220_o2_p_spl_01;
  wire n2220_o2_p_spl_1;
  wire n2254_o2_n_spl_;
  wire n2220_o2_n_spl_;
  wire g928_n_spl_;
  wire lo478_buf_o2_p_spl_;
  wire lo478_buf_o2_p_spl_0;
  wire lo478_buf_o2_p_spl_00;
  wire lo478_buf_o2_p_spl_000;
  wire lo478_buf_o2_p_spl_001;
  wire lo478_buf_o2_p_spl_01;
  wire lo478_buf_o2_p_spl_010;
  wire lo478_buf_o2_p_spl_1;
  wire lo478_buf_o2_p_spl_10;
  wire lo478_buf_o2_p_spl_11;
  wire n1913_inv_p_spl_;
  wire n1913_inv_p_spl_0;
  wire n1913_inv_p_spl_00;
  wire n1913_inv_p_spl_1;
  wire lo478_buf_o2_n_spl_;
  wire lo478_buf_o2_n_spl_0;
  wire lo478_buf_o2_n_spl_00;
  wire lo478_buf_o2_n_spl_1;
  wire lo466_buf_o2_p_spl_;
  wire lo466_buf_o2_p_spl_0;
  wire lo466_buf_o2_p_spl_00;
  wire lo466_buf_o2_p_spl_000;
  wire lo466_buf_o2_p_spl_001;
  wire lo466_buf_o2_p_spl_01;
  wire lo466_buf_o2_p_spl_1;
  wire lo466_buf_o2_p_spl_10;
  wire lo466_buf_o2_p_spl_11;
  wire lo466_buf_o2_n_spl_;
  wire lo466_buf_o2_n_spl_0;
  wire lo466_buf_o2_n_spl_00;
  wire lo466_buf_o2_n_spl_000;
  wire lo466_buf_o2_n_spl_001;
  wire lo466_buf_o2_n_spl_01;
  wire lo466_buf_o2_n_spl_010;
  wire lo466_buf_o2_n_spl_011;
  wire lo466_buf_o2_n_spl_1;
  wire lo466_buf_o2_n_spl_10;
  wire lo466_buf_o2_n_spl_100;
  wire lo466_buf_o2_n_spl_101;
  wire lo466_buf_o2_n_spl_11;
  wire lo466_buf_o2_n_spl_110;
  wire g938_n_spl_;
  wire g938_n_spl_0;
  wire n1794_lo_p_spl_;
  wire n2178_lo_p_spl_;
  wire n1926_lo_p_spl_;
  wire n2046_lo_p_spl_;
  wire n2322_lo_p_spl_;
  wire n2682_lo_p_spl_;
  wire n2442_lo_p_spl_;
  wire n2562_lo_p_spl_;
  wire n2826_lo_p_spl_;
  wire lo498_buf_o2_n_spl_;
  wire lo498_buf_o2_n_spl_0;
  wire lo498_buf_o2_n_spl_1;
  wire g1005_n_spl_;
  wire lo502_buf_o2_n_spl_;
  wire lo502_buf_o2_n_spl_0;
  wire g948_n_spl_;
  wire lo510_buf_o2_n_spl_;
  wire lo510_buf_o2_n_spl_0;
  wire lo510_buf_o2_n_spl_1;
  wire g1011_n_spl_;
  wire g903_n_spl_;
  wire g903_n_spl_0;
  wire g903_n_spl_1;
  wire n2970_lo_n_spl_;
  wire n2970_lo_n_spl_0;
  wire n2970_lo_n_spl_1;
  wire g1016_n_spl_;
  wire g1021_n_spl_;
  wire n2994_lo_n_spl_;
  wire n2994_lo_n_spl_0;
  wire n2994_lo_n_spl_1;
  wire g954_n_spl_;
  wire g919_n_spl_;
  wire g919_n_spl_0;
  wire n3006_lo_n_spl_;
  wire n3006_lo_n_spl_0;
  wire n3006_lo_n_spl_1;
  wire g1028_n_spl_;
  wire n3018_lo_n_spl_;
  wire g951_n_spl_;
  wire g960_n_spl_;
  wire g957_n_spl_;
  wire g963_n_spl_;
  wire n3126_lo_p_spl_;
  wire n3138_lo_p_spl_;
  wire g919_p_spl_;
  wire g913_n_spl_;
  wire n2196_o2_p_spl_;
  wire n2196_o2_p_spl_0;
  wire n2196_o2_p_spl_1;
  wire g942_n_spl_;
  wire g968_n_spl_;
  wire n2386_o2_p_spl_;
  wire n2386_o2_p_spl_0;
  wire g1051_n_spl_;
  wire g1051_n_spl_0;
  wire g1051_n_spl_1;
  wire g897_p_spl_;
  wire g898_p_spl_;
  wire g1055_n_spl_;
  wire g1055_n_spl_0;
  wire lo514_buf_o2_p_spl_;
  wire g944_n_spl_;
  wire g945_p_spl_;
  wire n3030_lo_p_spl_;
  wire n3030_lo_n_spl_;
  wire n2386_o2_n_spl_;
  wire n2386_o2_n_spl_0;
  wire g1071_n_spl_;
  wire g1072_p_spl_;
  wire lo550_buf_o2_n_spl_;
  wire lo550_buf_o2_n_spl_0;
  wire g1075_n_spl_;
  wire g1076_p_spl_;
  wire g1079_n_spl_;
  wire g1082_n_spl_;
  wire n2612_o2_n_spl_;
  wire n2616_o2_n_spl_;
  wire g974_n_spl_;
  wire n3102_lo_p_spl_;
  wire n3114_lo_p_spl_;
  wire g929_n_spl_;
  wire g902_p_spl_;
  wire n3294_lo_n_spl_;
  wire n3294_lo_p_spl_;
  wire lo550_buf_o2_p_spl_;
  wire lo550_buf_o2_p_spl_0;
  wire g1099_p_spl_;
  wire g1107_p_spl_;
  wire g907_n_spl_;
  wire g980_n_spl_;
  wire g980_n_spl_0;
  wire g1112_n_spl_;
  wire n3258_lo_p_spl_;
  wire n3270_lo_n_spl_;
  wire n3258_lo_n_spl_;
  wire n3270_lo_p_spl_;
  wire lo498_buf_o2_p_spl_;
  wire lo502_buf_o2_p_spl_;
  wire lo502_buf_o2_p_spl_0;
  wire n2982_lo_p_spl_;
  wire n2994_lo_p_spl_;
  wire n2994_lo_p_spl_0;
  wire n3282_lo_n_spl_;
  wire n3282_lo_p_spl_;
  wire lo510_buf_o2_p_spl_;
  wire n4039_o2_n_spl_;
  wire g1055_p_spl_;
  wire lo606_buf_o2_p_spl_;
  wire lo610_buf_o2_n_spl_;
  wire lo606_buf_o2_n_spl_;
  wire lo610_buf_o2_p_spl_;
  wire lo590_buf_o2_p_spl_;
  wire lo594_buf_o2_n_spl_;
  wire lo590_buf_o2_n_spl_;
  wire lo594_buf_o2_p_spl_;
  wire g1141_p_spl_;
  wire g1144_p_spl_;
  wire g1141_n_spl_;
  wire g1144_n_spl_;
  wire n3210_lo_p_spl_;
  wire n3222_lo_n_spl_;
  wire n3210_lo_n_spl_;
  wire n3222_lo_p_spl_;
  wire g1156_n_spl_;
  wire g1159_p_spl_;
  wire n2539_o2_p_spl_;
  wire n2539_o2_n_spl_;
  wire n1475_inv_n_spl_;
  wire n2367_o2_n_spl_;
  wire g1164_p_spl_;
  wire g1167_p_spl_;
  wire g1164_n_spl_;
  wire g1167_n_spl_;
  wire g1051_p_spl_;
  wire n3063_lo_p_spl_;
  wire g941_n_spl_;
  wire g941_n_spl_0;
  wire g941_n_spl_1;
  wire n2919_lo_p_spl_;
  wire g941_p_spl_;
  wire g941_p_spl_0;
  wire g941_p_spl_00;
  wire g941_p_spl_1;
  wire g995_n_spl_;
  wire g995_n_spl_0;
  wire g1204_p_spl_;
  wire lo578_buf_o2_n_spl_;
  wire lo578_buf_o2_n_spl_0;
  wire lo578_buf_o2_n_spl_00;
  wire lo578_buf_o2_n_spl_000;
  wire lo578_buf_o2_n_spl_001;
  wire lo578_buf_o2_n_spl_01;
  wire lo578_buf_o2_n_spl_010;
  wire lo578_buf_o2_n_spl_011;
  wire lo578_buf_o2_n_spl_1;
  wire lo578_buf_o2_n_spl_10;
  wire lo578_buf_o2_n_spl_11;
  wire lo578_buf_o2_p_spl_;
  wire lo578_buf_o2_p_spl_0;
  wire lo578_buf_o2_p_spl_00;
  wire lo578_buf_o2_p_spl_000;
  wire lo578_buf_o2_p_spl_001;
  wire lo578_buf_o2_p_spl_01;
  wire lo578_buf_o2_p_spl_010;
  wire lo578_buf_o2_p_spl_011;
  wire lo578_buf_o2_p_spl_1;
  wire lo578_buf_o2_p_spl_10;
  wire lo578_buf_o2_p_spl_100;
  wire lo578_buf_o2_p_spl_11;
  wire lo582_buf_o2_p_spl_;
  wire lo582_buf_o2_p_spl_0;
  wire lo582_buf_o2_p_spl_1;
  wire lo582_buf_o2_n_spl_;
  wire lo582_buf_o2_n_spl_0;
  wire g1040_n_spl_;
  wire g1183_n_spl_;
  wire n3075_lo_p_spl_;
  wire n2943_lo_p_spl_;
  wire n3087_lo_p_spl_;
  wire n2955_lo_p_spl_;
  wire n3039_lo_p_spl_;
  wire n2907_lo_p_spl_;
  wire g986_n_spl_;
  wire lo576_buf_o2_p_spl_;
  wire lo576_buf_o2_p_spl_0;
  wire lo576_buf_o2_p_spl_00;
  wire lo576_buf_o2_p_spl_1;
  wire lo576_buf_o2_n_spl_;
  wire lo576_buf_o2_n_spl_0;
  wire lo576_buf_o2_n_spl_1;
  wire n3156_lo_n_spl_;
  wire n3156_lo_p_spl_;
  wire n3156_lo_p_spl_0;
  wire n2808_lo_n_spl_;
  wire n2808_lo_p_spl_;
  wire n2808_lo_p_spl_0;
  wire g1284_n_spl_;
  wire g1288_n_spl_;
  wire n2901_lo_n_spl_;
  wire n3057_lo_n_spl_;
  wire n3057_lo_n_spl_0;
  wire g742_n_spl_;
  wire g758_p_spl_;
  wire g761_n_spl_;
  wire g766_p_spl_;
  wire g838_n_spl_;
  wire g859_p_spl_;
  wire g895_n_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  buf

  (
    G42_p,
    G42
  );


  not

  (
    G42_n,
    G42
  );


  buf

  (
    G43_p,
    G43
  );


  not

  (
    G43_n,
    G43
  );


  buf

  (
    G44_p,
    G44
  );


  not

  (
    G44_n,
    G44
  );


  buf

  (
    G45_p,
    G45
  );


  not

  (
    G45_n,
    G45
  );


  buf

  (
    G46_p,
    G46
  );


  not

  (
    G46_n,
    G46
  );


  buf

  (
    G47_p,
    G47
  );


  not

  (
    G47_n,
    G47
  );


  buf

  (
    G48_p,
    G48
  );


  not

  (
    G48_n,
    G48
  );


  buf

  (
    G49_p,
    G49
  );


  not

  (
    G49_n,
    G49
  );


  buf

  (
    G50_p,
    G50
  );


  not

  (
    G50_n,
    G50
  );


  buf

  (
    G51_p,
    G51
  );


  not

  (
    G51_n,
    G51
  );


  buf

  (
    G52_p,
    G52
  );


  not

  (
    G52_n,
    G52
  );


  buf

  (
    G53_p,
    G53
  );


  not

  (
    G53_n,
    G53
  );


  buf

  (
    G54_p,
    G54
  );


  not

  (
    G54_n,
    G54
  );


  buf

  (
    G55_p,
    G55
  );


  not

  (
    G55_n,
    G55
  );


  buf

  (
    G56_p,
    G56
  );


  not

  (
    G56_n,
    G56
  );


  buf

  (
    G57_p,
    G57
  );


  not

  (
    G57_n,
    G57
  );


  buf

  (
    G58_p,
    G58
  );


  not

  (
    G58_n,
    G58
  );


  buf

  (
    G59_p,
    G59
  );


  not

  (
    G59_n,
    G59
  );


  buf

  (
    G60_p,
    G60
  );


  not

  (
    G60_n,
    G60
  );


  buf

  (
    G61_p,
    G61
  );


  not

  (
    G61_n,
    G61
  );


  buf

  (
    G62_p,
    G62
  );


  not

  (
    G62_n,
    G62
  );


  buf

  (
    G63_p,
    G63
  );


  not

  (
    G63_n,
    G63
  );


  buf

  (
    G64_p,
    G64
  );


  not

  (
    G64_n,
    G64
  );


  buf

  (
    G65_p,
    G65
  );


  not

  (
    G65_n,
    G65
  );


  buf

  (
    G66_p,
    G66
  );


  not

  (
    G66_n,
    G66
  );


  buf

  (
    G67_p,
    G67
  );


  not

  (
    G67_n,
    G67
  );


  buf

  (
    G68_p,
    G68
  );


  not

  (
    G68_n,
    G68
  );


  buf

  (
    G69_p,
    G69
  );


  not

  (
    G69_n,
    G69
  );


  buf

  (
    G70_p,
    G70
  );


  not

  (
    G70_n,
    G70
  );


  buf

  (
    G71_p,
    G71
  );


  not

  (
    G71_n,
    G71
  );


  buf

  (
    G72_p,
    G72
  );


  not

  (
    G72_n,
    G72
  );


  buf

  (
    G73_p,
    G73
  );


  not

  (
    G73_n,
    G73
  );


  buf

  (
    G74_p,
    G74
  );


  not

  (
    G74_n,
    G74
  );


  buf

  (
    G75_p,
    G75
  );


  not

  (
    G75_n,
    G75
  );


  buf

  (
    G76_p,
    G76
  );


  not

  (
    G76_n,
    G76
  );


  buf

  (
    G77_p,
    G77
  );


  not

  (
    G77_n,
    G77
  );


  buf

  (
    G78_p,
    G78
  );


  not

  (
    G78_n,
    G78
  );


  buf

  (
    G79_p,
    G79
  );


  not

  (
    G79_n,
    G79
  );


  buf

  (
    G80_p,
    G80
  );


  not

  (
    G80_n,
    G80
  );


  buf

  (
    G81_p,
    G81
  );


  not

  (
    G81_n,
    G81
  );


  buf

  (
    G82_p,
    G82
  );


  not

  (
    G82_n,
    G82
  );


  buf

  (
    G83_p,
    G83
  );


  not

  (
    G83_n,
    G83
  );


  buf

  (
    G84_p,
    G84
  );


  not

  (
    G84_n,
    G84
  );


  buf

  (
    G85_p,
    G85
  );


  not

  (
    G85_n,
    G85
  );


  buf

  (
    G86_p,
    G86
  );


  not

  (
    G86_n,
    G86
  );


  buf

  (
    G87_p,
    G87
  );


  not

  (
    G87_n,
    G87
  );


  buf

  (
    G88_p,
    G88
  );


  not

  (
    G88_n,
    G88
  );


  buf

  (
    G89_p,
    G89
  );


  not

  (
    G89_n,
    G89
  );


  buf

  (
    G90_p,
    G90
  );


  not

  (
    G90_n,
    G90
  );


  buf

  (
    G91_p,
    G91
  );


  not

  (
    G91_n,
    G91
  );


  buf

  (
    G92_p,
    G92
  );


  not

  (
    G92_n,
    G92
  );


  buf

  (
    G93_p,
    G93
  );


  not

  (
    G93_n,
    G93
  );


  buf

  (
    G94_p,
    G94
  );


  not

  (
    G94_n,
    G94
  );


  buf

  (
    G95_p,
    G95
  );


  not

  (
    G95_n,
    G95
  );


  buf

  (
    G96_p,
    G96
  );


  not

  (
    G96_n,
    G96
  );


  buf

  (
    G97_p,
    G97
  );


  not

  (
    G97_n,
    G97
  );


  buf

  (
    G98_p,
    G98
  );


  not

  (
    G98_n,
    G98
  );


  buf

  (
    G99_p,
    G99
  );


  not

  (
    G99_n,
    G99
  );


  buf

  (
    G100_p,
    G100
  );


  not

  (
    G100_n,
    G100
  );


  buf

  (
    G101_p,
    G101
  );


  not

  (
    G101_n,
    G101
  );


  buf

  (
    G102_p,
    G102
  );


  not

  (
    G102_n,
    G102
  );


  buf

  (
    G103_p,
    G103
  );


  not

  (
    G103_n,
    G103
  );


  buf

  (
    G104_p,
    G104
  );


  not

  (
    G104_n,
    G104
  );


  buf

  (
    G105_p,
    G105
  );


  not

  (
    G105_n,
    G105
  );


  buf

  (
    G106_p,
    G106
  );


  not

  (
    G106_n,
    G106
  );


  buf

  (
    G107_p,
    G107
  );


  not

  (
    G107_n,
    G107
  );


  buf

  (
    G108_p,
    G108
  );


  not

  (
    G108_n,
    G108
  );


  buf

  (
    G109_p,
    G109
  );


  not

  (
    G109_n,
    G109
  );


  buf

  (
    G110_p,
    G110
  );


  not

  (
    G110_n,
    G110
  );


  buf

  (
    G111_p,
    G111
  );


  not

  (
    G111_n,
    G111
  );


  buf

  (
    G112_p,
    G112
  );


  not

  (
    G112_n,
    G112
  );


  buf

  (
    G113_p,
    G113
  );


  not

  (
    G113_n,
    G113
  );


  buf

  (
    G114_p,
    G114
  );


  not

  (
    G114_n,
    G114
  );


  buf

  (
    G115_p,
    G115
  );


  not

  (
    G115_n,
    G115
  );


  buf

  (
    G116_p,
    G116
  );


  not

  (
    G116_n,
    G116
  );


  buf

  (
    G117_p,
    G117
  );


  not

  (
    G117_n,
    G117
  );


  buf

  (
    G118_p,
    G118
  );


  not

  (
    G118_n,
    G118
  );


  buf

  (
    G119_p,
    G119
  );


  not

  (
    G119_n,
    G119
  );


  buf

  (
    G120_p,
    G120
  );


  not

  (
    G120_n,
    G120
  );


  buf

  (
    G121_p,
    G121
  );


  not

  (
    G121_n,
    G121
  );


  buf

  (
    G122_p,
    G122
  );


  not

  (
    G122_n,
    G122
  );


  buf

  (
    G123_p,
    G123
  );


  not

  (
    G123_n,
    G123
  );


  buf

  (
    G124_p,
    G124
  );


  not

  (
    G124_n,
    G124
  );


  buf

  (
    G125_p,
    G125
  );


  not

  (
    G125_n,
    G125
  );


  buf

  (
    G126_p,
    G126
  );


  not

  (
    G126_n,
    G126
  );


  buf

  (
    G127_p,
    G127
  );


  not

  (
    G127_n,
    G127
  );


  buf

  (
    G128_p,
    G128
  );


  not

  (
    G128_n,
    G128
  );


  buf

  (
    G129_p,
    G129
  );


  not

  (
    G129_n,
    G129
  );


  buf

  (
    G130_p,
    G130
  );


  not

  (
    G130_n,
    G130
  );


  buf

  (
    G131_p,
    G131
  );


  not

  (
    G131_n,
    G131
  );


  buf

  (
    G132_p,
    G132
  );


  not

  (
    G132_n,
    G132
  );


  buf

  (
    G133_p,
    G133
  );


  not

  (
    G133_n,
    G133
  );


  buf

  (
    G134_p,
    G134
  );


  not

  (
    G134_n,
    G134
  );


  buf

  (
    G135_p,
    G135
  );


  not

  (
    G135_n,
    G135
  );


  buf

  (
    G136_p,
    G136
  );


  not

  (
    G136_n,
    G136
  );


  buf

  (
    G137_p,
    G137
  );


  not

  (
    G137_n,
    G137
  );


  buf

  (
    G138_p,
    G138
  );


  not

  (
    G138_n,
    G138
  );


  buf

  (
    G139_p,
    G139
  );


  not

  (
    G139_n,
    G139
  );


  buf

  (
    G140_p,
    G140
  );


  not

  (
    G140_n,
    G140
  );


  buf

  (
    G141_p,
    G141
  );


  not

  (
    G141_n,
    G141
  );


  buf

  (
    G142_p,
    G142
  );


  not

  (
    G142_n,
    G142
  );


  buf

  (
    G143_p,
    G143
  );


  not

  (
    G143_n,
    G143
  );


  buf

  (
    G144_p,
    G144
  );


  not

  (
    G144_n,
    G144
  );


  buf

  (
    G145_p,
    G145
  );


  not

  (
    G145_n,
    G145
  );


  buf

  (
    G146_p,
    G146
  );


  not

  (
    G146_n,
    G146
  );


  buf

  (
    G147_p,
    G147
  );


  not

  (
    G147_n,
    G147
  );


  buf

  (
    G148_p,
    G148
  );


  not

  (
    G148_n,
    G148
  );


  buf

  (
    G149_p,
    G149
  );


  not

  (
    G149_n,
    G149
  );


  buf

  (
    G150_p,
    G150
  );


  not

  (
    G150_n,
    G150
  );


  buf

  (
    G151_p,
    G151
  );


  not

  (
    G151_n,
    G151
  );


  buf

  (
    G152_p,
    G152
  );


  not

  (
    G152_n,
    G152
  );


  buf

  (
    G153_p,
    G153
  );


  not

  (
    G153_n,
    G153
  );


  buf

  (
    G154_p,
    G154
  );


  not

  (
    G154_n,
    G154
  );


  buf

  (
    G155_p,
    G155
  );


  not

  (
    G155_n,
    G155
  );


  buf

  (
    G156_p,
    G156
  );


  not

  (
    G156_n,
    G156
  );


  buf

  (
    G157_p,
    G157
  );


  not

  (
    G157_n,
    G157
  );


  buf

  (
    n1416_lo_p,
    n1416_lo
  );


  not

  (
    n1416_lo_n,
    n1416_lo
  );


  buf

  (
    n1419_lo_p,
    n1419_lo
  );


  not

  (
    n1419_lo_n,
    n1419_lo
  );


  buf

  (
    n1422_lo_p,
    n1422_lo
  );


  not

  (
    n1422_lo_n,
    n1422_lo
  );


  buf

  (
    n1425_lo_p,
    n1425_lo
  );


  not

  (
    n1425_lo_n,
    n1425_lo
  );


  buf

  (
    n1428_lo_p,
    n1428_lo
  );


  not

  (
    n1428_lo_n,
    n1428_lo
  );


  buf

  (
    n1431_lo_p,
    n1431_lo
  );


  not

  (
    n1431_lo_n,
    n1431_lo
  );


  buf

  (
    n1434_lo_p,
    n1434_lo
  );


  not

  (
    n1434_lo_n,
    n1434_lo
  );


  buf

  (
    n1437_lo_p,
    n1437_lo
  );


  not

  (
    n1437_lo_n,
    n1437_lo
  );


  buf

  (
    n1440_lo_p,
    n1440_lo
  );


  not

  (
    n1440_lo_n,
    n1440_lo
  );


  buf

  (
    n1443_lo_p,
    n1443_lo
  );


  not

  (
    n1443_lo_n,
    n1443_lo
  );


  buf

  (
    n1446_lo_p,
    n1446_lo
  );


  not

  (
    n1446_lo_n,
    n1446_lo
  );


  buf

  (
    n1449_lo_p,
    n1449_lo
  );


  not

  (
    n1449_lo_n,
    n1449_lo
  );


  buf

  (
    n1452_lo_p,
    n1452_lo
  );


  not

  (
    n1452_lo_n,
    n1452_lo
  );


  buf

  (
    n1455_lo_p,
    n1455_lo
  );


  not

  (
    n1455_lo_n,
    n1455_lo
  );


  buf

  (
    n1458_lo_p,
    n1458_lo
  );


  not

  (
    n1458_lo_n,
    n1458_lo
  );


  buf

  (
    n1464_lo_p,
    n1464_lo
  );


  not

  (
    n1464_lo_n,
    n1464_lo
  );


  buf

  (
    n1467_lo_p,
    n1467_lo
  );


  not

  (
    n1467_lo_n,
    n1467_lo
  );


  buf

  (
    n1470_lo_p,
    n1470_lo
  );


  not

  (
    n1470_lo_n,
    n1470_lo
  );


  buf

  (
    n1476_lo_p,
    n1476_lo
  );


  not

  (
    n1476_lo_n,
    n1476_lo
  );


  buf

  (
    n1479_lo_p,
    n1479_lo
  );


  not

  (
    n1479_lo_n,
    n1479_lo
  );


  buf

  (
    n1482_lo_p,
    n1482_lo
  );


  not

  (
    n1482_lo_n,
    n1482_lo
  );


  buf

  (
    n1488_lo_p,
    n1488_lo
  );


  not

  (
    n1488_lo_n,
    n1488_lo
  );


  buf

  (
    n1491_lo_p,
    n1491_lo
  );


  not

  (
    n1491_lo_n,
    n1491_lo
  );


  buf

  (
    n1494_lo_p,
    n1494_lo
  );


  not

  (
    n1494_lo_n,
    n1494_lo
  );


  buf

  (
    n1497_lo_p,
    n1497_lo
  );


  not

  (
    n1497_lo_n,
    n1497_lo
  );


  buf

  (
    n1500_lo_p,
    n1500_lo
  );


  not

  (
    n1500_lo_n,
    n1500_lo
  );


  buf

  (
    n1503_lo_p,
    n1503_lo
  );


  not

  (
    n1503_lo_n,
    n1503_lo
  );


  buf

  (
    n1512_lo_p,
    n1512_lo
  );


  not

  (
    n1512_lo_n,
    n1512_lo
  );


  buf

  (
    n1515_lo_p,
    n1515_lo
  );


  not

  (
    n1515_lo_n,
    n1515_lo
  );


  buf

  (
    n1518_lo_p,
    n1518_lo
  );


  not

  (
    n1518_lo_n,
    n1518_lo
  );


  buf

  (
    n1521_lo_p,
    n1521_lo
  );


  not

  (
    n1521_lo_n,
    n1521_lo
  );


  buf

  (
    n1524_lo_p,
    n1524_lo
  );


  not

  (
    n1524_lo_n,
    n1524_lo
  );


  buf

  (
    n1527_lo_p,
    n1527_lo
  );


  not

  (
    n1527_lo_n,
    n1527_lo
  );


  buf

  (
    n1530_lo_p,
    n1530_lo
  );


  not

  (
    n1530_lo_n,
    n1530_lo
  );


  buf

  (
    n1533_lo_p,
    n1533_lo
  );


  not

  (
    n1533_lo_n,
    n1533_lo
  );


  buf

  (
    n1536_lo_p,
    n1536_lo
  );


  not

  (
    n1536_lo_n,
    n1536_lo
  );


  buf

  (
    n1539_lo_p,
    n1539_lo
  );


  not

  (
    n1539_lo_n,
    n1539_lo
  );


  buf

  (
    n1542_lo_p,
    n1542_lo
  );


  not

  (
    n1542_lo_n,
    n1542_lo
  );


  buf

  (
    n1545_lo_p,
    n1545_lo
  );


  not

  (
    n1545_lo_n,
    n1545_lo
  );


  buf

  (
    n1548_lo_p,
    n1548_lo
  );


  not

  (
    n1548_lo_n,
    n1548_lo
  );


  buf

  (
    n1551_lo_p,
    n1551_lo
  );


  not

  (
    n1551_lo_n,
    n1551_lo
  );


  buf

  (
    n1554_lo_p,
    n1554_lo
  );


  not

  (
    n1554_lo_n,
    n1554_lo
  );


  buf

  (
    n1560_lo_p,
    n1560_lo
  );


  not

  (
    n1560_lo_n,
    n1560_lo
  );


  buf

  (
    n1563_lo_p,
    n1563_lo
  );


  not

  (
    n1563_lo_n,
    n1563_lo
  );


  buf

  (
    n1566_lo_p,
    n1566_lo
  );


  not

  (
    n1566_lo_n,
    n1566_lo
  );


  buf

  (
    n1572_lo_p,
    n1572_lo
  );


  not

  (
    n1572_lo_n,
    n1572_lo
  );


  buf

  (
    n1575_lo_p,
    n1575_lo
  );


  not

  (
    n1575_lo_n,
    n1575_lo
  );


  buf

  (
    n1578_lo_p,
    n1578_lo
  );


  not

  (
    n1578_lo_n,
    n1578_lo
  );


  buf

  (
    n1584_lo_p,
    n1584_lo
  );


  not

  (
    n1584_lo_n,
    n1584_lo
  );


  buf

  (
    n1587_lo_p,
    n1587_lo
  );


  not

  (
    n1587_lo_n,
    n1587_lo
  );


  buf

  (
    n1590_lo_p,
    n1590_lo
  );


  not

  (
    n1590_lo_n,
    n1590_lo
  );


  buf

  (
    n1596_lo_p,
    n1596_lo
  );


  not

  (
    n1596_lo_n,
    n1596_lo
  );


  buf

  (
    n1599_lo_p,
    n1599_lo
  );


  not

  (
    n1599_lo_n,
    n1599_lo
  );


  buf

  (
    n1602_lo_p,
    n1602_lo
  );


  not

  (
    n1602_lo_n,
    n1602_lo
  );


  buf

  (
    n1608_lo_p,
    n1608_lo
  );


  not

  (
    n1608_lo_n,
    n1608_lo
  );


  buf

  (
    n1611_lo_p,
    n1611_lo
  );


  not

  (
    n1611_lo_n,
    n1611_lo
  );


  buf

  (
    n1614_lo_p,
    n1614_lo
  );


  not

  (
    n1614_lo_n,
    n1614_lo
  );


  buf

  (
    n1620_lo_p,
    n1620_lo
  );


  not

  (
    n1620_lo_n,
    n1620_lo
  );


  buf

  (
    n1623_lo_p,
    n1623_lo
  );


  not

  (
    n1623_lo_n,
    n1623_lo
  );


  buf

  (
    n1626_lo_p,
    n1626_lo
  );


  not

  (
    n1626_lo_n,
    n1626_lo
  );


  buf

  (
    n1632_lo_p,
    n1632_lo
  );


  not

  (
    n1632_lo_n,
    n1632_lo
  );


  buf

  (
    n1635_lo_p,
    n1635_lo
  );


  not

  (
    n1635_lo_n,
    n1635_lo
  );


  buf

  (
    n1638_lo_p,
    n1638_lo
  );


  not

  (
    n1638_lo_n,
    n1638_lo
  );


  buf

  (
    n1644_lo_p,
    n1644_lo
  );


  not

  (
    n1644_lo_n,
    n1644_lo
  );


  buf

  (
    n1647_lo_p,
    n1647_lo
  );


  not

  (
    n1647_lo_n,
    n1647_lo
  );


  buf

  (
    n1650_lo_p,
    n1650_lo
  );


  not

  (
    n1650_lo_n,
    n1650_lo
  );


  buf

  (
    n1656_lo_p,
    n1656_lo
  );


  not

  (
    n1656_lo_n,
    n1656_lo
  );


  buf

  (
    n1659_lo_p,
    n1659_lo
  );


  not

  (
    n1659_lo_n,
    n1659_lo
  );


  buf

  (
    n1662_lo_p,
    n1662_lo
  );


  not

  (
    n1662_lo_n,
    n1662_lo
  );


  buf

  (
    n1668_lo_p,
    n1668_lo
  );


  not

  (
    n1668_lo_n,
    n1668_lo
  );


  buf

  (
    n1671_lo_p,
    n1671_lo
  );


  not

  (
    n1671_lo_n,
    n1671_lo
  );


  buf

  (
    n1674_lo_p,
    n1674_lo
  );


  not

  (
    n1674_lo_n,
    n1674_lo
  );


  buf

  (
    n1680_lo_p,
    n1680_lo
  );


  not

  (
    n1680_lo_n,
    n1680_lo
  );


  buf

  (
    n1683_lo_p,
    n1683_lo
  );


  not

  (
    n1683_lo_n,
    n1683_lo
  );


  buf

  (
    n1686_lo_p,
    n1686_lo
  );


  not

  (
    n1686_lo_n,
    n1686_lo
  );


  buf

  (
    n1692_lo_p,
    n1692_lo
  );


  not

  (
    n1692_lo_n,
    n1692_lo
  );


  buf

  (
    n1695_lo_p,
    n1695_lo
  );


  not

  (
    n1695_lo_n,
    n1695_lo
  );


  buf

  (
    n1698_lo_p,
    n1698_lo
  );


  not

  (
    n1698_lo_n,
    n1698_lo
  );


  buf

  (
    n1704_lo_p,
    n1704_lo
  );


  not

  (
    n1704_lo_n,
    n1704_lo
  );


  buf

  (
    n1707_lo_p,
    n1707_lo
  );


  not

  (
    n1707_lo_n,
    n1707_lo
  );


  buf

  (
    n1710_lo_p,
    n1710_lo
  );


  not

  (
    n1710_lo_n,
    n1710_lo
  );


  buf

  (
    n1716_lo_p,
    n1716_lo
  );


  not

  (
    n1716_lo_n,
    n1716_lo
  );


  buf

  (
    n1719_lo_p,
    n1719_lo
  );


  not

  (
    n1719_lo_n,
    n1719_lo
  );


  buf

  (
    n1722_lo_p,
    n1722_lo
  );


  not

  (
    n1722_lo_n,
    n1722_lo
  );


  buf

  (
    n1728_lo_p,
    n1728_lo
  );


  not

  (
    n1728_lo_n,
    n1728_lo
  );


  buf

  (
    n1731_lo_p,
    n1731_lo
  );


  not

  (
    n1731_lo_n,
    n1731_lo
  );


  buf

  (
    n1734_lo_p,
    n1734_lo
  );


  not

  (
    n1734_lo_n,
    n1734_lo
  );


  buf

  (
    n1740_lo_p,
    n1740_lo
  );


  not

  (
    n1740_lo_n,
    n1740_lo
  );


  buf

  (
    n1743_lo_p,
    n1743_lo
  );


  not

  (
    n1743_lo_n,
    n1743_lo
  );


  buf

  (
    n1746_lo_p,
    n1746_lo
  );


  not

  (
    n1746_lo_n,
    n1746_lo
  );


  buf

  (
    n1749_lo_p,
    n1749_lo
  );


  not

  (
    n1749_lo_n,
    n1749_lo
  );


  buf

  (
    n1752_lo_p,
    n1752_lo
  );


  not

  (
    n1752_lo_n,
    n1752_lo
  );


  buf

  (
    n1755_lo_p,
    n1755_lo
  );


  not

  (
    n1755_lo_n,
    n1755_lo
  );


  buf

  (
    n1758_lo_p,
    n1758_lo
  );


  not

  (
    n1758_lo_n,
    n1758_lo
  );


  buf

  (
    n1761_lo_p,
    n1761_lo
  );


  not

  (
    n1761_lo_n,
    n1761_lo
  );


  buf

  (
    n1764_lo_p,
    n1764_lo
  );


  not

  (
    n1764_lo_n,
    n1764_lo
  );


  buf

  (
    n1776_lo_p,
    n1776_lo
  );


  not

  (
    n1776_lo_n,
    n1776_lo
  );


  buf

  (
    n1788_lo_p,
    n1788_lo
  );


  not

  (
    n1788_lo_n,
    n1788_lo
  );


  buf

  (
    n1791_lo_p,
    n1791_lo
  );


  not

  (
    n1791_lo_n,
    n1791_lo
  );


  buf

  (
    n1794_lo_p,
    n1794_lo
  );


  not

  (
    n1794_lo_n,
    n1794_lo
  );


  buf

  (
    n1797_lo_p,
    n1797_lo
  );


  not

  (
    n1797_lo_n,
    n1797_lo
  );


  buf

  (
    n1800_lo_p,
    n1800_lo
  );


  not

  (
    n1800_lo_n,
    n1800_lo
  );


  buf

  (
    n1803_lo_p,
    n1803_lo
  );


  not

  (
    n1803_lo_n,
    n1803_lo
  );


  buf

  (
    n1812_lo_p,
    n1812_lo
  );


  not

  (
    n1812_lo_n,
    n1812_lo
  );


  buf

  (
    n1815_lo_p,
    n1815_lo
  );


  not

  (
    n1815_lo_n,
    n1815_lo
  );


  buf

  (
    n1824_lo_p,
    n1824_lo
  );


  not

  (
    n1824_lo_n,
    n1824_lo
  );


  buf

  (
    n1827_lo_p,
    n1827_lo
  );


  not

  (
    n1827_lo_n,
    n1827_lo
  );


  buf

  (
    n1836_lo_p,
    n1836_lo
  );


  not

  (
    n1836_lo_n,
    n1836_lo
  );


  buf

  (
    n1839_lo_p,
    n1839_lo
  );


  not

  (
    n1839_lo_n,
    n1839_lo
  );


  buf

  (
    n1848_lo_p,
    n1848_lo
  );


  not

  (
    n1848_lo_n,
    n1848_lo
  );


  buf

  (
    n1851_lo_p,
    n1851_lo
  );


  not

  (
    n1851_lo_n,
    n1851_lo
  );


  buf

  (
    n1860_lo_p,
    n1860_lo
  );


  not

  (
    n1860_lo_n,
    n1860_lo
  );


  buf

  (
    n1872_lo_p,
    n1872_lo
  );


  not

  (
    n1872_lo_n,
    n1872_lo
  );


  buf

  (
    n1875_lo_p,
    n1875_lo
  );


  not

  (
    n1875_lo_n,
    n1875_lo
  );


  buf

  (
    n1884_lo_p,
    n1884_lo
  );


  not

  (
    n1884_lo_n,
    n1884_lo
  );


  buf

  (
    n1896_lo_p,
    n1896_lo
  );


  not

  (
    n1896_lo_n,
    n1896_lo
  );


  buf

  (
    n1899_lo_p,
    n1899_lo
  );


  not

  (
    n1899_lo_n,
    n1899_lo
  );


  buf

  (
    n1908_lo_p,
    n1908_lo
  );


  not

  (
    n1908_lo_n,
    n1908_lo
  );


  buf

  (
    n1920_lo_p,
    n1920_lo
  );


  not

  (
    n1920_lo_n,
    n1920_lo
  );


  buf

  (
    n1923_lo_p,
    n1923_lo
  );


  not

  (
    n1923_lo_n,
    n1923_lo
  );


  buf

  (
    n1926_lo_p,
    n1926_lo
  );


  not

  (
    n1926_lo_n,
    n1926_lo
  );


  buf

  (
    n1929_lo_p,
    n1929_lo
  );


  not

  (
    n1929_lo_n,
    n1929_lo
  );


  buf

  (
    n1932_lo_p,
    n1932_lo
  );


  not

  (
    n1932_lo_n,
    n1932_lo
  );


  buf

  (
    n1935_lo_p,
    n1935_lo
  );


  not

  (
    n1935_lo_n,
    n1935_lo
  );


  buf

  (
    n1944_lo_p,
    n1944_lo
  );


  not

  (
    n1944_lo_n,
    n1944_lo
  );


  buf

  (
    n1947_lo_p,
    n1947_lo
  );


  not

  (
    n1947_lo_n,
    n1947_lo
  );


  buf

  (
    n1956_lo_p,
    n1956_lo
  );


  not

  (
    n1956_lo_n,
    n1956_lo
  );


  buf

  (
    n1959_lo_p,
    n1959_lo
  );


  not

  (
    n1959_lo_n,
    n1959_lo
  );


  buf

  (
    n1962_lo_p,
    n1962_lo
  );


  not

  (
    n1962_lo_n,
    n1962_lo
  );


  buf

  (
    n1968_lo_p,
    n1968_lo
  );


  not

  (
    n1968_lo_n,
    n1968_lo
  );


  buf

  (
    n1971_lo_p,
    n1971_lo
  );


  not

  (
    n1971_lo_n,
    n1971_lo
  );


  buf

  (
    n1980_lo_p,
    n1980_lo
  );


  not

  (
    n1980_lo_n,
    n1980_lo
  );


  buf

  (
    n1983_lo_p,
    n1983_lo
  );


  not

  (
    n1983_lo_n,
    n1983_lo
  );


  buf

  (
    n1992_lo_p,
    n1992_lo
  );


  not

  (
    n1992_lo_n,
    n1992_lo
  );


  buf

  (
    n1995_lo_p,
    n1995_lo
  );


  not

  (
    n1995_lo_n,
    n1995_lo
  );


  buf

  (
    n2004_lo_p,
    n2004_lo
  );


  not

  (
    n2004_lo_n,
    n2004_lo
  );


  buf

  (
    n2016_lo_p,
    n2016_lo
  );


  not

  (
    n2016_lo_n,
    n2016_lo
  );


  buf

  (
    n2019_lo_p,
    n2019_lo
  );


  not

  (
    n2019_lo_n,
    n2019_lo
  );


  buf

  (
    n2028_lo_p,
    n2028_lo
  );


  not

  (
    n2028_lo_n,
    n2028_lo
  );


  buf

  (
    n2040_lo_p,
    n2040_lo
  );


  not

  (
    n2040_lo_n,
    n2040_lo
  );


  buf

  (
    n2043_lo_p,
    n2043_lo
  );


  not

  (
    n2043_lo_n,
    n2043_lo
  );


  buf

  (
    n2046_lo_p,
    n2046_lo
  );


  not

  (
    n2046_lo_n,
    n2046_lo
  );


  buf

  (
    n2049_lo_p,
    n2049_lo
  );


  not

  (
    n2049_lo_n,
    n2049_lo
  );


  buf

  (
    n2052_lo_p,
    n2052_lo
  );


  not

  (
    n2052_lo_n,
    n2052_lo
  );


  buf

  (
    n2055_lo_p,
    n2055_lo
  );


  not

  (
    n2055_lo_n,
    n2055_lo
  );


  buf

  (
    n2064_lo_p,
    n2064_lo
  );


  not

  (
    n2064_lo_n,
    n2064_lo
  );


  buf

  (
    n2067_lo_p,
    n2067_lo
  );


  not

  (
    n2067_lo_n,
    n2067_lo
  );


  buf

  (
    n2076_lo_p,
    n2076_lo
  );


  not

  (
    n2076_lo_n,
    n2076_lo
  );


  buf

  (
    n2079_lo_p,
    n2079_lo
  );


  not

  (
    n2079_lo_n,
    n2079_lo
  );


  buf

  (
    n2088_lo_p,
    n2088_lo
  );


  not

  (
    n2088_lo_n,
    n2088_lo
  );


  buf

  (
    n2091_lo_p,
    n2091_lo
  );


  not

  (
    n2091_lo_n,
    n2091_lo
  );


  buf

  (
    n2100_lo_p,
    n2100_lo
  );


  not

  (
    n2100_lo_n,
    n2100_lo
  );


  buf

  (
    n2103_lo_p,
    n2103_lo
  );


  not

  (
    n2103_lo_n,
    n2103_lo
  );


  buf

  (
    n2112_lo_p,
    n2112_lo
  );


  not

  (
    n2112_lo_n,
    n2112_lo
  );


  buf

  (
    n2115_lo_p,
    n2115_lo
  );


  not

  (
    n2115_lo_n,
    n2115_lo
  );


  buf

  (
    n2124_lo_p,
    n2124_lo
  );


  not

  (
    n2124_lo_n,
    n2124_lo
  );


  buf

  (
    n2127_lo_p,
    n2127_lo
  );


  not

  (
    n2127_lo_n,
    n2127_lo
  );


  buf

  (
    n2136_lo_p,
    n2136_lo
  );


  not

  (
    n2136_lo_n,
    n2136_lo
  );


  buf

  (
    n2148_lo_p,
    n2148_lo
  );


  not

  (
    n2148_lo_n,
    n2148_lo
  );


  buf

  (
    n2151_lo_p,
    n2151_lo
  );


  not

  (
    n2151_lo_n,
    n2151_lo
  );


  buf

  (
    n2160_lo_p,
    n2160_lo
  );


  not

  (
    n2160_lo_n,
    n2160_lo
  );


  buf

  (
    n2172_lo_p,
    n2172_lo
  );


  not

  (
    n2172_lo_n,
    n2172_lo
  );


  buf

  (
    n2175_lo_p,
    n2175_lo
  );


  not

  (
    n2175_lo_n,
    n2175_lo
  );


  buf

  (
    n2178_lo_p,
    n2178_lo
  );


  not

  (
    n2178_lo_n,
    n2178_lo
  );


  buf

  (
    n2181_lo_p,
    n2181_lo
  );


  not

  (
    n2181_lo_n,
    n2181_lo
  );


  buf

  (
    n2184_lo_p,
    n2184_lo
  );


  not

  (
    n2184_lo_n,
    n2184_lo
  );


  buf

  (
    n2187_lo_p,
    n2187_lo
  );


  not

  (
    n2187_lo_n,
    n2187_lo
  );


  buf

  (
    n2196_lo_p,
    n2196_lo
  );


  not

  (
    n2196_lo_n,
    n2196_lo
  );


  buf

  (
    n2199_lo_p,
    n2199_lo
  );


  not

  (
    n2199_lo_n,
    n2199_lo
  );


  buf

  (
    n2208_lo_p,
    n2208_lo
  );


  not

  (
    n2208_lo_n,
    n2208_lo
  );


  buf

  (
    n2211_lo_p,
    n2211_lo
  );


  not

  (
    n2211_lo_n,
    n2211_lo
  );


  buf

  (
    n2220_lo_p,
    n2220_lo
  );


  not

  (
    n2220_lo_n,
    n2220_lo
  );


  buf

  (
    n2223_lo_p,
    n2223_lo
  );


  not

  (
    n2223_lo_n,
    n2223_lo
  );


  buf

  (
    n2232_lo_p,
    n2232_lo
  );


  not

  (
    n2232_lo_n,
    n2232_lo
  );


  buf

  (
    n2235_lo_p,
    n2235_lo
  );


  not

  (
    n2235_lo_n,
    n2235_lo
  );


  buf

  (
    n2244_lo_p,
    n2244_lo
  );


  not

  (
    n2244_lo_n,
    n2244_lo
  );


  buf

  (
    n2247_lo_p,
    n2247_lo
  );


  not

  (
    n2247_lo_n,
    n2247_lo
  );


  buf

  (
    n2256_lo_p,
    n2256_lo
  );


  not

  (
    n2256_lo_n,
    n2256_lo
  );


  buf

  (
    n2259_lo_p,
    n2259_lo
  );


  not

  (
    n2259_lo_n,
    n2259_lo
  );


  buf

  (
    n2268_lo_p,
    n2268_lo
  );


  not

  (
    n2268_lo_n,
    n2268_lo
  );


  buf

  (
    n2280_lo_p,
    n2280_lo
  );


  not

  (
    n2280_lo_n,
    n2280_lo
  );


  buf

  (
    n2283_lo_p,
    n2283_lo
  );


  not

  (
    n2283_lo_n,
    n2283_lo
  );


  buf

  (
    n2292_lo_p,
    n2292_lo
  );


  not

  (
    n2292_lo_n,
    n2292_lo
  );


  buf

  (
    n2295_lo_p,
    n2295_lo
  );


  not

  (
    n2295_lo_n,
    n2295_lo
  );


  buf

  (
    n2298_lo_p,
    n2298_lo
  );


  not

  (
    n2298_lo_n,
    n2298_lo
  );


  buf

  (
    n2301_lo_p,
    n2301_lo
  );


  not

  (
    n2301_lo_n,
    n2301_lo
  );


  buf

  (
    n2304_lo_p,
    n2304_lo
  );


  not

  (
    n2304_lo_n,
    n2304_lo
  );


  buf

  (
    n2307_lo_p,
    n2307_lo
  );


  not

  (
    n2307_lo_n,
    n2307_lo
  );


  buf

  (
    n2316_lo_p,
    n2316_lo
  );


  not

  (
    n2316_lo_n,
    n2316_lo
  );


  buf

  (
    n2319_lo_p,
    n2319_lo
  );


  not

  (
    n2319_lo_n,
    n2319_lo
  );


  buf

  (
    n2322_lo_p,
    n2322_lo
  );


  not

  (
    n2322_lo_n,
    n2322_lo
  );


  buf

  (
    n2325_lo_p,
    n2325_lo
  );


  not

  (
    n2325_lo_n,
    n2325_lo
  );


  buf

  (
    n2328_lo_p,
    n2328_lo
  );


  not

  (
    n2328_lo_n,
    n2328_lo
  );


  buf

  (
    n2331_lo_p,
    n2331_lo
  );


  not

  (
    n2331_lo_n,
    n2331_lo
  );


  buf

  (
    n2340_lo_p,
    n2340_lo
  );


  not

  (
    n2340_lo_n,
    n2340_lo
  );


  buf

  (
    n2343_lo_p,
    n2343_lo
  );


  not

  (
    n2343_lo_n,
    n2343_lo
  );


  buf

  (
    n2376_lo_p,
    n2376_lo
  );


  not

  (
    n2376_lo_n,
    n2376_lo
  );


  buf

  (
    n2379_lo_p,
    n2379_lo
  );


  not

  (
    n2379_lo_n,
    n2379_lo
  );


  buf

  (
    n2388_lo_p,
    n2388_lo
  );


  not

  (
    n2388_lo_n,
    n2388_lo
  );


  buf

  (
    n2391_lo_p,
    n2391_lo
  );


  not

  (
    n2391_lo_n,
    n2391_lo
  );


  buf

  (
    n2400_lo_p,
    n2400_lo
  );


  not

  (
    n2400_lo_n,
    n2400_lo
  );


  buf

  (
    n2403_lo_p,
    n2403_lo
  );


  not

  (
    n2403_lo_n,
    n2403_lo
  );


  buf

  (
    n2412_lo_p,
    n2412_lo
  );


  not

  (
    n2412_lo_n,
    n2412_lo
  );


  buf

  (
    n2415_lo_p,
    n2415_lo
  );


  not

  (
    n2415_lo_n,
    n2415_lo
  );


  buf

  (
    n2424_lo_p,
    n2424_lo
  );


  not

  (
    n2424_lo_n,
    n2424_lo
  );


  buf

  (
    n2427_lo_p,
    n2427_lo
  );


  not

  (
    n2427_lo_n,
    n2427_lo
  );


  buf

  (
    n2436_lo_p,
    n2436_lo
  );


  not

  (
    n2436_lo_n,
    n2436_lo
  );


  buf

  (
    n2439_lo_p,
    n2439_lo
  );


  not

  (
    n2439_lo_n,
    n2439_lo
  );


  buf

  (
    n2442_lo_p,
    n2442_lo
  );


  not

  (
    n2442_lo_n,
    n2442_lo
  );


  buf

  (
    n2445_lo_p,
    n2445_lo
  );


  not

  (
    n2445_lo_n,
    n2445_lo
  );


  buf

  (
    n2448_lo_p,
    n2448_lo
  );


  not

  (
    n2448_lo_n,
    n2448_lo
  );


  buf

  (
    n2451_lo_p,
    n2451_lo
  );


  not

  (
    n2451_lo_n,
    n2451_lo
  );


  buf

  (
    n2460_lo_p,
    n2460_lo
  );


  not

  (
    n2460_lo_n,
    n2460_lo
  );


  buf

  (
    n2463_lo_p,
    n2463_lo
  );


  not

  (
    n2463_lo_n,
    n2463_lo
  );


  buf

  (
    n2496_lo_p,
    n2496_lo
  );


  not

  (
    n2496_lo_n,
    n2496_lo
  );


  buf

  (
    n2499_lo_p,
    n2499_lo
  );


  not

  (
    n2499_lo_n,
    n2499_lo
  );


  buf

  (
    n2508_lo_p,
    n2508_lo
  );


  not

  (
    n2508_lo_n,
    n2508_lo
  );


  buf

  (
    n2511_lo_p,
    n2511_lo
  );


  not

  (
    n2511_lo_n,
    n2511_lo
  );


  buf

  (
    n2520_lo_p,
    n2520_lo
  );


  not

  (
    n2520_lo_n,
    n2520_lo
  );


  buf

  (
    n2523_lo_p,
    n2523_lo
  );


  not

  (
    n2523_lo_n,
    n2523_lo
  );


  buf

  (
    n2532_lo_p,
    n2532_lo
  );


  not

  (
    n2532_lo_n,
    n2532_lo
  );


  buf

  (
    n2535_lo_p,
    n2535_lo
  );


  not

  (
    n2535_lo_n,
    n2535_lo
  );


  buf

  (
    n2544_lo_p,
    n2544_lo
  );


  not

  (
    n2544_lo_n,
    n2544_lo
  );


  buf

  (
    n2547_lo_p,
    n2547_lo
  );


  not

  (
    n2547_lo_n,
    n2547_lo
  );


  buf

  (
    n2556_lo_p,
    n2556_lo
  );


  not

  (
    n2556_lo_n,
    n2556_lo
  );


  buf

  (
    n2559_lo_p,
    n2559_lo
  );


  not

  (
    n2559_lo_n,
    n2559_lo
  );


  buf

  (
    n2562_lo_p,
    n2562_lo
  );


  not

  (
    n2562_lo_n,
    n2562_lo
  );


  buf

  (
    n2565_lo_p,
    n2565_lo
  );


  not

  (
    n2565_lo_n,
    n2565_lo
  );


  buf

  (
    n2568_lo_p,
    n2568_lo
  );


  not

  (
    n2568_lo_n,
    n2568_lo
  );


  buf

  (
    n2571_lo_p,
    n2571_lo
  );


  not

  (
    n2571_lo_n,
    n2571_lo
  );


  buf

  (
    n2580_lo_p,
    n2580_lo
  );


  not

  (
    n2580_lo_n,
    n2580_lo
  );


  buf

  (
    n2583_lo_p,
    n2583_lo
  );


  not

  (
    n2583_lo_n,
    n2583_lo
  );


  buf

  (
    n2616_lo_p,
    n2616_lo
  );


  not

  (
    n2616_lo_n,
    n2616_lo
  );


  buf

  (
    n2619_lo_p,
    n2619_lo
  );


  not

  (
    n2619_lo_n,
    n2619_lo
  );


  buf

  (
    n2628_lo_p,
    n2628_lo
  );


  not

  (
    n2628_lo_n,
    n2628_lo
  );


  buf

  (
    n2631_lo_p,
    n2631_lo
  );


  not

  (
    n2631_lo_n,
    n2631_lo
  );


  buf

  (
    n2640_lo_p,
    n2640_lo
  );


  not

  (
    n2640_lo_n,
    n2640_lo
  );


  buf

  (
    n2643_lo_p,
    n2643_lo
  );


  not

  (
    n2643_lo_n,
    n2643_lo
  );


  buf

  (
    n2652_lo_p,
    n2652_lo
  );


  not

  (
    n2652_lo_n,
    n2652_lo
  );


  buf

  (
    n2655_lo_p,
    n2655_lo
  );


  not

  (
    n2655_lo_n,
    n2655_lo
  );


  buf

  (
    n2664_lo_p,
    n2664_lo
  );


  not

  (
    n2664_lo_n,
    n2664_lo
  );


  buf

  (
    n2667_lo_p,
    n2667_lo
  );


  not

  (
    n2667_lo_n,
    n2667_lo
  );


  buf

  (
    n2676_lo_p,
    n2676_lo
  );


  not

  (
    n2676_lo_n,
    n2676_lo
  );


  buf

  (
    n2679_lo_p,
    n2679_lo
  );


  not

  (
    n2679_lo_n,
    n2679_lo
  );


  buf

  (
    n2682_lo_p,
    n2682_lo
  );


  not

  (
    n2682_lo_n,
    n2682_lo
  );


  buf

  (
    n2685_lo_p,
    n2685_lo
  );


  not

  (
    n2685_lo_n,
    n2685_lo
  );


  buf

  (
    n2688_lo_p,
    n2688_lo
  );


  not

  (
    n2688_lo_n,
    n2688_lo
  );


  buf

  (
    n2691_lo_p,
    n2691_lo
  );


  not

  (
    n2691_lo_n,
    n2691_lo
  );


  buf

  (
    n2700_lo_p,
    n2700_lo
  );


  not

  (
    n2700_lo_n,
    n2700_lo
  );


  buf

  (
    n2703_lo_p,
    n2703_lo
  );


  not

  (
    n2703_lo_n,
    n2703_lo
  );


  buf

  (
    n2736_lo_p,
    n2736_lo
  );


  not

  (
    n2736_lo_n,
    n2736_lo
  );


  buf

  (
    n2739_lo_p,
    n2739_lo
  );


  not

  (
    n2739_lo_n,
    n2739_lo
  );


  buf

  (
    n2748_lo_p,
    n2748_lo
  );


  not

  (
    n2748_lo_n,
    n2748_lo
  );


  buf

  (
    n2751_lo_p,
    n2751_lo
  );


  not

  (
    n2751_lo_n,
    n2751_lo
  );


  buf

  (
    n2760_lo_p,
    n2760_lo
  );


  not

  (
    n2760_lo_n,
    n2760_lo
  );


  buf

  (
    n2763_lo_p,
    n2763_lo
  );


  not

  (
    n2763_lo_n,
    n2763_lo
  );


  buf

  (
    n2772_lo_p,
    n2772_lo
  );


  not

  (
    n2772_lo_n,
    n2772_lo
  );


  buf

  (
    n2775_lo_p,
    n2775_lo
  );


  not

  (
    n2775_lo_n,
    n2775_lo
  );


  buf

  (
    n2784_lo_p,
    n2784_lo
  );


  not

  (
    n2784_lo_n,
    n2784_lo
  );


  buf

  (
    n2787_lo_p,
    n2787_lo
  );


  not

  (
    n2787_lo_n,
    n2787_lo
  );


  buf

  (
    n2790_lo_p,
    n2790_lo
  );


  not

  (
    n2790_lo_n,
    n2790_lo
  );


  buf

  (
    n2793_lo_p,
    n2793_lo
  );


  not

  (
    n2793_lo_n,
    n2793_lo
  );


  buf

  (
    n2796_lo_p,
    n2796_lo
  );


  not

  (
    n2796_lo_n,
    n2796_lo
  );


  buf

  (
    n2799_lo_p,
    n2799_lo
  );


  not

  (
    n2799_lo_n,
    n2799_lo
  );


  buf

  (
    n2802_lo_p,
    n2802_lo
  );


  not

  (
    n2802_lo_n,
    n2802_lo
  );


  buf

  (
    n2805_lo_p,
    n2805_lo
  );


  not

  (
    n2805_lo_n,
    n2805_lo
  );


  buf

  (
    n2808_lo_p,
    n2808_lo
  );


  not

  (
    n2808_lo_n,
    n2808_lo
  );


  buf

  (
    n2820_lo_p,
    n2820_lo
  );


  not

  (
    n2820_lo_n,
    n2820_lo
  );


  buf

  (
    n2823_lo_p,
    n2823_lo
  );


  not

  (
    n2823_lo_n,
    n2823_lo
  );


  buf

  (
    n2826_lo_p,
    n2826_lo
  );


  not

  (
    n2826_lo_n,
    n2826_lo
  );


  buf

  (
    n2829_lo_p,
    n2829_lo
  );


  not

  (
    n2829_lo_n,
    n2829_lo
  );


  buf

  (
    n2832_lo_p,
    n2832_lo
  );


  not

  (
    n2832_lo_n,
    n2832_lo
  );


  buf

  (
    n2835_lo_p,
    n2835_lo
  );


  not

  (
    n2835_lo_n,
    n2835_lo
  );


  buf

  (
    n2838_lo_p,
    n2838_lo
  );


  not

  (
    n2838_lo_n,
    n2838_lo
  );


  buf

  (
    n2841_lo_p,
    n2841_lo
  );


  not

  (
    n2841_lo_n,
    n2841_lo
  );


  buf

  (
    n2844_lo_p,
    n2844_lo
  );


  not

  (
    n2844_lo_n,
    n2844_lo
  );


  buf

  (
    n2856_lo_p,
    n2856_lo
  );


  not

  (
    n2856_lo_n,
    n2856_lo
  );


  buf

  (
    n2859_lo_p,
    n2859_lo
  );


  not

  (
    n2859_lo_n,
    n2859_lo
  );


  buf

  (
    n2862_lo_p,
    n2862_lo
  );


  not

  (
    n2862_lo_n,
    n2862_lo
  );


  buf

  (
    n2865_lo_p,
    n2865_lo
  );


  not

  (
    n2865_lo_n,
    n2865_lo
  );


  buf

  (
    n2868_lo_p,
    n2868_lo
  );


  not

  (
    n2868_lo_n,
    n2868_lo
  );


  buf

  (
    n2871_lo_p,
    n2871_lo
  );


  not

  (
    n2871_lo_n,
    n2871_lo
  );


  buf

  (
    n2874_lo_p,
    n2874_lo
  );


  not

  (
    n2874_lo_n,
    n2874_lo
  );


  buf

  (
    n2877_lo_p,
    n2877_lo
  );


  not

  (
    n2877_lo_n,
    n2877_lo
  );


  buf

  (
    n2880_lo_p,
    n2880_lo
  );


  not

  (
    n2880_lo_n,
    n2880_lo
  );


  buf

  (
    n2883_lo_p,
    n2883_lo
  );


  not

  (
    n2883_lo_n,
    n2883_lo
  );


  buf

  (
    n2886_lo_p,
    n2886_lo
  );


  not

  (
    n2886_lo_n,
    n2886_lo
  );


  buf

  (
    n2889_lo_p,
    n2889_lo
  );


  not

  (
    n2889_lo_n,
    n2889_lo
  );


  buf

  (
    n2892_lo_p,
    n2892_lo
  );


  not

  (
    n2892_lo_n,
    n2892_lo
  );


  buf

  (
    n2895_lo_p,
    n2895_lo
  );


  not

  (
    n2895_lo_n,
    n2895_lo
  );


  buf

  (
    n2898_lo_p,
    n2898_lo
  );


  not

  (
    n2898_lo_n,
    n2898_lo
  );


  buf

  (
    n2901_lo_p,
    n2901_lo
  );


  not

  (
    n2901_lo_n,
    n2901_lo
  );


  buf

  (
    n2904_lo_p,
    n2904_lo
  );


  not

  (
    n2904_lo_n,
    n2904_lo
  );


  buf

  (
    n2907_lo_p,
    n2907_lo
  );


  not

  (
    n2907_lo_n,
    n2907_lo
  );


  buf

  (
    n2916_lo_p,
    n2916_lo
  );


  not

  (
    n2916_lo_n,
    n2916_lo
  );


  buf

  (
    n2919_lo_p,
    n2919_lo
  );


  not

  (
    n2919_lo_n,
    n2919_lo
  );


  buf

  (
    n2925_lo_p,
    n2925_lo
  );


  not

  (
    n2925_lo_n,
    n2925_lo
  );


  buf

  (
    n2928_lo_p,
    n2928_lo
  );


  not

  (
    n2928_lo_n,
    n2928_lo
  );


  buf

  (
    n2940_lo_p,
    n2940_lo
  );


  not

  (
    n2940_lo_n,
    n2940_lo
  );


  buf

  (
    n2943_lo_p,
    n2943_lo
  );


  not

  (
    n2943_lo_n,
    n2943_lo
  );


  buf

  (
    n2952_lo_p,
    n2952_lo
  );


  not

  (
    n2952_lo_n,
    n2952_lo
  );


  buf

  (
    n2955_lo_p,
    n2955_lo
  );


  not

  (
    n2955_lo_n,
    n2955_lo
  );


  buf

  (
    n2961_lo_p,
    n2961_lo
  );


  not

  (
    n2961_lo_n,
    n2961_lo
  );


  buf

  (
    n2964_lo_p,
    n2964_lo
  );


  not

  (
    n2964_lo_n,
    n2964_lo
  );


  buf

  (
    n2967_lo_p,
    n2967_lo
  );


  not

  (
    n2967_lo_n,
    n2967_lo
  );


  buf

  (
    n2970_lo_p,
    n2970_lo
  );


  not

  (
    n2970_lo_n,
    n2970_lo
  );


  buf

  (
    n2976_lo_p,
    n2976_lo
  );


  not

  (
    n2976_lo_n,
    n2976_lo
  );


  buf

  (
    n2979_lo_p,
    n2979_lo
  );


  not

  (
    n2979_lo_n,
    n2979_lo
  );


  buf

  (
    n2982_lo_p,
    n2982_lo
  );


  not

  (
    n2982_lo_n,
    n2982_lo
  );


  buf

  (
    n2988_lo_p,
    n2988_lo
  );


  not

  (
    n2988_lo_n,
    n2988_lo
  );


  buf

  (
    n2991_lo_p,
    n2991_lo
  );


  not

  (
    n2991_lo_n,
    n2991_lo
  );


  buf

  (
    n2994_lo_p,
    n2994_lo
  );


  not

  (
    n2994_lo_n,
    n2994_lo
  );


  buf

  (
    n2997_lo_p,
    n2997_lo
  );


  not

  (
    n2997_lo_n,
    n2997_lo
  );


  buf

  (
    n3000_lo_p,
    n3000_lo
  );


  not

  (
    n3000_lo_n,
    n3000_lo
  );


  buf

  (
    n3003_lo_p,
    n3003_lo
  );


  not

  (
    n3003_lo_n,
    n3003_lo
  );


  buf

  (
    n3006_lo_p,
    n3006_lo
  );


  not

  (
    n3006_lo_n,
    n3006_lo
  );


  buf

  (
    n3012_lo_p,
    n3012_lo
  );


  not

  (
    n3012_lo_n,
    n3012_lo
  );


  buf

  (
    n3015_lo_p,
    n3015_lo
  );


  not

  (
    n3015_lo_n,
    n3015_lo
  );


  buf

  (
    n3018_lo_p,
    n3018_lo
  );


  not

  (
    n3018_lo_n,
    n3018_lo
  );


  buf

  (
    n3021_lo_p,
    n3021_lo
  );


  not

  (
    n3021_lo_n,
    n3021_lo
  );


  buf

  (
    n3024_lo_p,
    n3024_lo
  );


  not

  (
    n3024_lo_n,
    n3024_lo
  );


  buf

  (
    n3027_lo_p,
    n3027_lo
  );


  not

  (
    n3027_lo_n,
    n3027_lo
  );


  buf

  (
    n3030_lo_p,
    n3030_lo
  );


  not

  (
    n3030_lo_n,
    n3030_lo
  );


  buf

  (
    n3033_lo_p,
    n3033_lo
  );


  not

  (
    n3033_lo_n,
    n3033_lo
  );


  buf

  (
    n3036_lo_p,
    n3036_lo
  );


  not

  (
    n3036_lo_n,
    n3036_lo
  );


  buf

  (
    n3039_lo_p,
    n3039_lo
  );


  not

  (
    n3039_lo_n,
    n3039_lo
  );


  buf

  (
    n3045_lo_p,
    n3045_lo
  );


  not

  (
    n3045_lo_n,
    n3045_lo
  );


  buf

  (
    n3048_lo_p,
    n3048_lo
  );


  not

  (
    n3048_lo_n,
    n3048_lo
  );


  buf

  (
    n3051_lo_p,
    n3051_lo
  );


  not

  (
    n3051_lo_n,
    n3051_lo
  );


  buf

  (
    n3054_lo_p,
    n3054_lo
  );


  not

  (
    n3054_lo_n,
    n3054_lo
  );


  buf

  (
    n3057_lo_p,
    n3057_lo
  );


  not

  (
    n3057_lo_n,
    n3057_lo
  );


  buf

  (
    n3060_lo_p,
    n3060_lo
  );


  not

  (
    n3060_lo_n,
    n3060_lo
  );


  buf

  (
    n3063_lo_p,
    n3063_lo
  );


  not

  (
    n3063_lo_n,
    n3063_lo
  );


  buf

  (
    n3069_lo_p,
    n3069_lo
  );


  not

  (
    n3069_lo_n,
    n3069_lo
  );


  buf

  (
    n3072_lo_p,
    n3072_lo
  );


  not

  (
    n3072_lo_n,
    n3072_lo
  );


  buf

  (
    n3075_lo_p,
    n3075_lo
  );


  not

  (
    n3075_lo_n,
    n3075_lo
  );


  buf

  (
    n3081_lo_p,
    n3081_lo
  );


  not

  (
    n3081_lo_n,
    n3081_lo
  );


  buf

  (
    n3084_lo_p,
    n3084_lo
  );


  not

  (
    n3084_lo_n,
    n3084_lo
  );


  buf

  (
    n3087_lo_p,
    n3087_lo
  );


  not

  (
    n3087_lo_n,
    n3087_lo
  );


  buf

  (
    n3093_lo_p,
    n3093_lo
  );


  not

  (
    n3093_lo_n,
    n3093_lo
  );


  buf

  (
    n3096_lo_p,
    n3096_lo
  );


  not

  (
    n3096_lo_n,
    n3096_lo
  );


  buf

  (
    n3099_lo_p,
    n3099_lo
  );


  not

  (
    n3099_lo_n,
    n3099_lo
  );


  buf

  (
    n3102_lo_p,
    n3102_lo
  );


  not

  (
    n3102_lo_n,
    n3102_lo
  );


  buf

  (
    n3105_lo_p,
    n3105_lo
  );


  not

  (
    n3105_lo_n,
    n3105_lo
  );


  buf

  (
    n3108_lo_p,
    n3108_lo
  );


  not

  (
    n3108_lo_n,
    n3108_lo
  );


  buf

  (
    n3111_lo_p,
    n3111_lo
  );


  not

  (
    n3111_lo_n,
    n3111_lo
  );


  buf

  (
    n3114_lo_p,
    n3114_lo
  );


  not

  (
    n3114_lo_n,
    n3114_lo
  );


  buf

  (
    n3117_lo_p,
    n3117_lo
  );


  not

  (
    n3117_lo_n,
    n3117_lo
  );


  buf

  (
    n3120_lo_p,
    n3120_lo
  );


  not

  (
    n3120_lo_n,
    n3120_lo
  );


  buf

  (
    n3123_lo_p,
    n3123_lo
  );


  not

  (
    n3123_lo_n,
    n3123_lo
  );


  buf

  (
    n3126_lo_p,
    n3126_lo
  );


  not

  (
    n3126_lo_n,
    n3126_lo
  );


  buf

  (
    n3129_lo_p,
    n3129_lo
  );


  not

  (
    n3129_lo_n,
    n3129_lo
  );


  buf

  (
    n3132_lo_p,
    n3132_lo
  );


  not

  (
    n3132_lo_n,
    n3132_lo
  );


  buf

  (
    n3135_lo_p,
    n3135_lo
  );


  not

  (
    n3135_lo_n,
    n3135_lo
  );


  buf

  (
    n3138_lo_p,
    n3138_lo
  );


  not

  (
    n3138_lo_n,
    n3138_lo
  );


  buf

  (
    n3141_lo_p,
    n3141_lo
  );


  not

  (
    n3141_lo_n,
    n3141_lo
  );


  buf

  (
    n3156_lo_p,
    n3156_lo
  );


  not

  (
    n3156_lo_n,
    n3156_lo
  );


  buf

  (
    n3168_lo_p,
    n3168_lo
  );


  not

  (
    n3168_lo_n,
    n3168_lo
  );


  buf

  (
    n3171_lo_p,
    n3171_lo
  );


  not

  (
    n3171_lo_n,
    n3171_lo
  );


  buf

  (
    n3174_lo_p,
    n3174_lo
  );


  not

  (
    n3174_lo_n,
    n3174_lo
  );


  buf

  (
    n3177_lo_p,
    n3177_lo
  );


  not

  (
    n3177_lo_n,
    n3177_lo
  );


  buf

  (
    n3180_lo_p,
    n3180_lo
  );


  not

  (
    n3180_lo_n,
    n3180_lo
  );


  buf

  (
    n3183_lo_p,
    n3183_lo
  );


  not

  (
    n3183_lo_n,
    n3183_lo
  );


  buf

  (
    n3192_lo_p,
    n3192_lo
  );


  not

  (
    n3192_lo_n,
    n3192_lo
  );


  buf

  (
    n3195_lo_p,
    n3195_lo
  );


  not

  (
    n3195_lo_n,
    n3195_lo
  );


  buf

  (
    n3204_lo_p,
    n3204_lo
  );


  not

  (
    n3204_lo_n,
    n3204_lo
  );


  buf

  (
    n3207_lo_p,
    n3207_lo
  );


  not

  (
    n3207_lo_n,
    n3207_lo
  );


  buf

  (
    n3210_lo_p,
    n3210_lo
  );


  not

  (
    n3210_lo_n,
    n3210_lo
  );


  buf

  (
    n3216_lo_p,
    n3216_lo
  );


  not

  (
    n3216_lo_n,
    n3216_lo
  );


  buf

  (
    n3219_lo_p,
    n3219_lo
  );


  not

  (
    n3219_lo_n,
    n3219_lo
  );


  buf

  (
    n3222_lo_p,
    n3222_lo
  );


  not

  (
    n3222_lo_n,
    n3222_lo
  );


  buf

  (
    n3228_lo_p,
    n3228_lo
  );


  not

  (
    n3228_lo_n,
    n3228_lo
  );


  buf

  (
    n3231_lo_p,
    n3231_lo
  );


  not

  (
    n3231_lo_n,
    n3231_lo
  );


  buf

  (
    n3240_lo_p,
    n3240_lo
  );


  not

  (
    n3240_lo_n,
    n3240_lo
  );


  buf

  (
    n3243_lo_p,
    n3243_lo
  );


  not

  (
    n3243_lo_n,
    n3243_lo
  );


  buf

  (
    n3252_lo_p,
    n3252_lo
  );


  not

  (
    n3252_lo_n,
    n3252_lo
  );


  buf

  (
    n3255_lo_p,
    n3255_lo
  );


  not

  (
    n3255_lo_n,
    n3255_lo
  );


  buf

  (
    n3258_lo_p,
    n3258_lo
  );


  not

  (
    n3258_lo_n,
    n3258_lo
  );


  buf

  (
    n3264_lo_p,
    n3264_lo
  );


  not

  (
    n3264_lo_n,
    n3264_lo
  );


  buf

  (
    n3267_lo_p,
    n3267_lo
  );


  not

  (
    n3267_lo_n,
    n3267_lo
  );


  buf

  (
    n3270_lo_p,
    n3270_lo
  );


  not

  (
    n3270_lo_n,
    n3270_lo
  );


  buf

  (
    n3276_lo_p,
    n3276_lo
  );


  not

  (
    n3276_lo_n,
    n3276_lo
  );


  buf

  (
    n3279_lo_p,
    n3279_lo
  );


  not

  (
    n3279_lo_n,
    n3279_lo
  );


  buf

  (
    n3282_lo_p,
    n3282_lo
  );


  not

  (
    n3282_lo_n,
    n3282_lo
  );


  buf

  (
    n3288_lo_p,
    n3288_lo
  );


  not

  (
    n3288_lo_n,
    n3288_lo
  );


  buf

  (
    n3291_lo_p,
    n3291_lo
  );


  not

  (
    n3291_lo_n,
    n3291_lo
  );


  buf

  (
    n3294_lo_p,
    n3294_lo
  );


  not

  (
    n3294_lo_n,
    n3294_lo
  );


  buf

  (
    n3603_o2_p,
    n3603_o2
  );


  not

  (
    n3603_o2_n,
    n3603_o2
  );


  buf

  (
    n3604_o2_p,
    n3604_o2
  );


  not

  (
    n3604_o2_n,
    n3604_o2
  );


  buf

  (
    n1391_inv_p,
    n1391_inv
  );


  not

  (
    n1391_inv_n,
    n1391_inv
  );


  buf

  (
    n3798_o2_p,
    n3798_o2
  );


  not

  (
    n3798_o2_n,
    n3798_o2
  );


  buf

  (
    n3846_o2_p,
    n3846_o2
  );


  not

  (
    n3846_o2_n,
    n3846_o2
  );


  buf

  (
    n4019_o2_p,
    n4019_o2
  );


  not

  (
    n4019_o2_n,
    n4019_o2
  );


  buf

  (
    n4017_o2_p,
    n4017_o2
  );


  not

  (
    n4017_o2_n,
    n4017_o2
  );


  buf

  (
    n2177_o2_p,
    n2177_o2
  );


  not

  (
    n2177_o2_n,
    n2177_o2
  );


  buf

  (
    n2150_o2_p,
    n2150_o2
  );


  not

  (
    n2150_o2_n,
    n2150_o2
  );


  buf

  (
    n2154_o2_p,
    n2154_o2
  );


  not

  (
    n2154_o2_n,
    n2154_o2
  );


  buf

  (
    n2184_o2_p,
    n2184_o2
  );


  not

  (
    n2184_o2_n,
    n2184_o2
  );


  buf

  (
    n2515_o2_p,
    n2515_o2
  );


  not

  (
    n2515_o2_n,
    n2515_o2
  );


  buf

  (
    n3837_o2_p,
    n3837_o2
  );


  not

  (
    n3837_o2_n,
    n3837_o2
  );


  buf

  (
    n2167_o2_p,
    n2167_o2
  );


  not

  (
    n2167_o2_n,
    n2167_o2
  );


  buf

  (
    n2118_o2_p,
    n2118_o2
  );


  not

  (
    n2118_o2_n,
    n2118_o2
  );


  buf

  (
    n2186_o2_p,
    n2186_o2
  );


  not

  (
    n2186_o2_n,
    n2186_o2
  );


  buf

  (
    n2174_o2_p,
    n2174_o2
  );


  not

  (
    n2174_o2_n,
    n2174_o2
  );


  buf

  (
    n3964_o2_p,
    n3964_o2
  );


  not

  (
    n3964_o2_n,
    n3964_o2
  );


  buf

  (
    n4005_o2_p,
    n4005_o2
  );


  not

  (
    n4005_o2_n,
    n4005_o2
  );


  buf

  (
    n4006_o2_p,
    n4006_o2
  );


  not

  (
    n4006_o2_n,
    n4006_o2
  );


  buf

  (
    n1445_inv_p,
    n1445_inv
  );


  not

  (
    n1445_inv_n,
    n1445_inv
  );


  buf

  (
    n2176_o2_p,
    n2176_o2
  );


  not

  (
    n2176_o2_n,
    n2176_o2
  );


  buf

  (
    n2227_o2_p,
    n2227_o2
  );


  not

  (
    n2227_o2_n,
    n2227_o2
  );


  buf

  (
    n2236_o2_p,
    n2236_o2
  );


  not

  (
    n2236_o2_n,
    n2236_o2
  );


  buf

  (
    n2245_o2_p,
    n2245_o2
  );


  not

  (
    n2245_o2_n,
    n2245_o2
  );


  buf

  (
    n2518_o2_p,
    n2518_o2
  );


  not

  (
    n2518_o2_n,
    n2518_o2
  );


  buf

  (
    n4023_o2_p,
    n4023_o2
  );


  not

  (
    n4023_o2_n,
    n4023_o2
  );


  buf

  (
    n1466_inv_p,
    n1466_inv
  );


  not

  (
    n1466_inv_n,
    n1466_inv
  );


  buf

  (
    n4038_o2_p,
    n4038_o2
  );


  not

  (
    n4038_o2_n,
    n4038_o2
  );


  buf

  (
    n4039_o2_p,
    n4039_o2
  );


  not

  (
    n4039_o2_n,
    n4039_o2
  );


  buf

  (
    n1475_inv_p,
    n1475_inv
  );


  not

  (
    n1475_inv_n,
    n1475_inv
  );


  buf

  (
    n2119_o2_p,
    n2119_o2
  );


  not

  (
    n2119_o2_n,
    n2119_o2
  );


  buf

  (
    n2275_o2_p,
    n2275_o2
  );


  not

  (
    n2275_o2_n,
    n2275_o2
  );


  buf

  (
    n2595_o2_p,
    n2595_o2
  );


  not

  (
    n2595_o2_n,
    n2595_o2
  );


  buf

  (
    n2594_o2_p,
    n2594_o2
  );


  not

  (
    n2594_o2_n,
    n2594_o2
  );


  buf

  (
    lo498_buf_o2_p,
    lo498_buf_o2
  );


  not

  (
    lo498_buf_o2_n,
    lo498_buf_o2
  );


  buf

  (
    lo502_buf_o2_p,
    lo502_buf_o2
  );


  not

  (
    lo502_buf_o2_n,
    lo502_buf_o2
  );


  buf

  (
    lo550_buf_o2_p,
    lo550_buf_o2
  );


  not

  (
    lo550_buf_o2_n,
    lo550_buf_o2
  );


  buf

  (
    n2596_o2_p,
    n2596_o2
  );


  not

  (
    n2596_o2_n,
    n2596_o2
  );


  buf

  (
    n2593_o2_p,
    n2593_o2
  );


  not

  (
    n2593_o2_n,
    n2593_o2
  );


  buf

  (
    n2668_o2_p,
    n2668_o2
  );


  not

  (
    n2668_o2_n,
    n2668_o2
  );


  buf

  (
    lo542_buf_o2_p,
    lo542_buf_o2
  );


  not

  (
    lo542_buf_o2_n,
    lo542_buf_o2
  );


  buf

  (
    n2667_o2_p,
    n2667_o2
  );


  not

  (
    n2667_o2_n,
    n2667_o2
  );


  buf

  (
    n2404_o2_p,
    n2404_o2
  );


  not

  (
    n2404_o2_n,
    n2404_o2
  );


  buf

  (
    n2410_o2_p,
    n2410_o2
  );


  not

  (
    n2410_o2_n,
    n2410_o2
  );


  buf

  (
    n2419_o2_p,
    n2419_o2
  );


  not

  (
    n2419_o2_n,
    n2419_o2
  );


  buf

  (
    n2392_o2_p,
    n2392_o2
  );


  not

  (
    n2392_o2_n,
    n2392_o2
  );


  buf

  (
    n2369_o2_p,
    n2369_o2
  );


  not

  (
    n2369_o2_n,
    n2369_o2
  );


  buf

  (
    n2397_o2_p,
    n2397_o2
  );


  not

  (
    n2397_o2_n,
    n2397_o2
  );


  buf

  (
    n2601_o2_p,
    n2601_o2
  );


  not

  (
    n2601_o2_n,
    n2601_o2
  );


  buf

  (
    n2658_o2_p,
    n2658_o2
  );


  not

  (
    n2658_o2_n,
    n2658_o2
  );


  buf

  (
    n2574_o2_p,
    n2574_o2
  );


  not

  (
    n2574_o2_n,
    n2574_o2
  );


  buf

  (
    n2205_o2_p,
    n2205_o2
  );


  not

  (
    n2205_o2_n,
    n2205_o2
  );


  buf

  (
    lo510_buf_o2_p,
    lo510_buf_o2
  );


  not

  (
    lo510_buf_o2_n,
    lo510_buf_o2
  );


  buf

  (
    lo514_buf_o2_p,
    lo514_buf_o2
  );


  not

  (
    lo514_buf_o2_n,
    lo514_buf_o2
  );


  buf

  (
    lo554_buf_o2_p,
    lo554_buf_o2
  );


  not

  (
    lo554_buf_o2_n,
    lo554_buf_o2
  );


  buf

  (
    lo558_buf_o2_p,
    lo558_buf_o2
  );


  not

  (
    lo558_buf_o2_n,
    lo558_buf_o2
  );


  buf

  (
    lo578_buf_o2_p,
    lo578_buf_o2
  );


  not

  (
    lo578_buf_o2_n,
    lo578_buf_o2
  );


  buf

  (
    n2254_o2_p,
    n2254_o2
  );


  not

  (
    n2254_o2_n,
    n2254_o2
  );


  buf

  (
    n2421_o2_p,
    n2421_o2
  );


  not

  (
    n2421_o2_n,
    n2421_o2
  );


  buf

  (
    n2422_o2_p,
    n2422_o2
  );


  not

  (
    n2422_o2_n,
    n2422_o2
  );


  buf

  (
    n2130_o2_p,
    n2130_o2
  );


  not

  (
    n2130_o2_n,
    n2130_o2
  );


  buf

  (
    n2127_o2_p,
    n2127_o2
  );


  not

  (
    n2127_o2_n,
    n2127_o2
  );


  buf

  (
    n2131_o2_p,
    n2131_o2
  );


  not

  (
    n2131_o2_n,
    n2131_o2
  );


  buf

  (
    n2128_o2_p,
    n2128_o2
  );


  not

  (
    n2128_o2_n,
    n2128_o2
  );


  buf

  (
    n2264_o2_p,
    n2264_o2
  );


  not

  (
    n2264_o2_n,
    n2264_o2
  );


  buf

  (
    n2467_o2_p,
    n2467_o2
  );


  not

  (
    n2467_o2_n,
    n2467_o2
  );


  buf

  (
    n2471_o2_p,
    n2471_o2
  );


  not

  (
    n2471_o2_n,
    n2471_o2
  );


  buf

  (
    n2488_o2_p,
    n2488_o2
  );


  not

  (
    n2488_o2_n,
    n2488_o2
  );


  buf

  (
    n2478_o2_p,
    n2478_o2
  );


  not

  (
    n2478_o2_n,
    n2478_o2
  );


  buf

  (
    n2486_o2_p,
    n2486_o2
  );


  not

  (
    n2486_o2_n,
    n2486_o2
  );


  buf

  (
    n2485_o2_p,
    n2485_o2
  );


  not

  (
    n2485_o2_n,
    n2485_o2
  );


  buf

  (
    n2498_o2_p,
    n2498_o2
  );


  not

  (
    n2498_o2_n,
    n2498_o2
  );


  buf

  (
    n2495_o2_p,
    n2495_o2
  );


  not

  (
    n2495_o2_n,
    n2495_o2
  );


  buf

  (
    n2496_o2_p,
    n2496_o2
  );


  not

  (
    n2496_o2_n,
    n2496_o2
  );


  buf

  (
    n2458_o2_p,
    n2458_o2
  );


  not

  (
    n2458_o2_n,
    n2458_o2
  );


  buf

  (
    n2643_o2_p,
    n2643_o2
  );


  not

  (
    n2643_o2_n,
    n2643_o2
  );


  buf

  (
    n2462_o2_p,
    n2462_o2
  );


  not

  (
    n2462_o2_n,
    n2462_o2
  );


  buf

  (
    n2468_o2_p,
    n2468_o2
  );


  not

  (
    n2468_o2_n,
    n2468_o2
  );


  buf

  (
    n2639_o2_p,
    n2639_o2
  );


  not

  (
    n2639_o2_n,
    n2639_o2
  );


  buf

  (
    n2499_o2_p,
    n2499_o2
  );


  not

  (
    n2499_o2_n,
    n2499_o2
  );


  buf

  (
    n2472_o2_p,
    n2472_o2
  );


  not

  (
    n2472_o2_n,
    n2472_o2
  );


  buf

  (
    n2474_o2_p,
    n2474_o2
  );


  not

  (
    n2474_o2_n,
    n2474_o2
  );


  buf

  (
    n2489_o2_p,
    n2489_o2
  );


  not

  (
    n2489_o2_n,
    n2489_o2
  );


  buf

  (
    n2321_o2_p,
    n2321_o2
  );


  not

  (
    n2321_o2_n,
    n2321_o2
  );


  buf

  (
    n2322_o2_p,
    n2322_o2
  );


  not

  (
    n2322_o2_n,
    n2322_o2
  );


  buf

  (
    n2640_o2_p,
    n2640_o2
  );


  not

  (
    n2640_o2_n,
    n2640_o2
  );


  buf

  (
    n2642_o2_p,
    n2642_o2
  );


  not

  (
    n2642_o2_n,
    n2642_o2
  );


  buf

  (
    n2187_o2_p,
    n2187_o2
  );


  not

  (
    n2187_o2_n,
    n2187_o2
  );


  buf

  (
    n2373_o2_p,
    n2373_o2
  );


  not

  (
    n2373_o2_n,
    n2373_o2
  );


  buf

  (
    n2603_o2_p,
    n2603_o2
  );


  not

  (
    n2603_o2_n,
    n2603_o2
  );


  buf

  (
    n2388_o2_p,
    n2388_o2
  );


  not

  (
    n2388_o2_n,
    n2388_o2
  );


  buf

  (
    n2437_o2_p,
    n2437_o2
  );


  not

  (
    n2437_o2_n,
    n2437_o2
  );


  buf

  (
    n2356_o2_p,
    n2356_o2
  );


  not

  (
    n2356_o2_n,
    n2356_o2
  );


  buf

  (
    n2452_o2_p,
    n2452_o2
  );


  not

  (
    n2452_o2_n,
    n2452_o2
  );


  buf

  (
    n2347_o2_p,
    n2347_o2
  );


  not

  (
    n2347_o2_n,
    n2347_o2
  );


  buf

  (
    n2329_o2_p,
    n2329_o2
  );


  not

  (
    n2329_o2_n,
    n2329_o2
  );


  buf

  (
    n2669_o2_p,
    n2669_o2
  );


  not

  (
    n2669_o2_n,
    n2669_o2
  );


  buf

  (
    n2332_o2_p,
    n2332_o2
  );


  not

  (
    n2332_o2_n,
    n2332_o2
  );


  buf

  (
    n2664_o2_p,
    n2664_o2
  );


  not

  (
    n2664_o2_n,
    n2664_o2
  );


  buf

  (
    n2665_o2_p,
    n2665_o2
  );


  not

  (
    n2665_o2_n,
    n2665_o2
  );


  buf

  (
    n2653_o2_p,
    n2653_o2
  );


  not

  (
    n2653_o2_n,
    n2653_o2
  );


  buf

  (
    n2654_o2_p,
    n2654_o2
  );


  not

  (
    n2654_o2_n,
    n2654_o2
  );


  buf

  (
    n2636_o2_p,
    n2636_o2
  );


  not

  (
    n2636_o2_n,
    n2636_o2
  );


  buf

  (
    n2660_o2_p,
    n2660_o2
  );


  not

  (
    n2660_o2_n,
    n2660_o2
  );


  buf

  (
    n2318_o2_p,
    n2318_o2
  );


  not

  (
    n2318_o2_n,
    n2318_o2
  );


  buf

  (
    n2319_o2_p,
    n2319_o2
  );


  not

  (
    n2319_o2_n,
    n2319_o2
  );


  buf

  (
    n2586_o2_p,
    n2586_o2
  );


  not

  (
    n2586_o2_n,
    n2586_o2
  );


  buf

  (
    n2587_o2_p,
    n2587_o2
  );


  not

  (
    n2587_o2_n,
    n2587_o2
  );


  buf

  (
    n2288_o2_p,
    n2288_o2
  );


  not

  (
    n2288_o2_n,
    n2288_o2
  );


  buf

  (
    n2344_o2_p,
    n2344_o2
  );


  not

  (
    n2344_o2_n,
    n2344_o2
  );


  buf

  (
    n2530_o2_p,
    n2530_o2
  );


  not

  (
    n2530_o2_n,
    n2530_o2
  );


  buf

  (
    n2303_o2_p,
    n2303_o2
  );


  not

  (
    n2303_o2_n,
    n2303_o2
  );


  buf

  (
    n2566_o2_p,
    n2566_o2
  );


  not

  (
    n2566_o2_n,
    n2566_o2
  );


  buf

  (
    n2567_o2_p,
    n2567_o2
  );


  not

  (
    n2567_o2_n,
    n2567_o2
  );


  buf

  (
    n2554_o2_p,
    n2554_o2
  );


  not

  (
    n2554_o2_n,
    n2554_o2
  );


  buf

  (
    n2194_o2_p,
    n2194_o2
  );


  not

  (
    n2194_o2_n,
    n2194_o2
  );


  buf

  (
    lo582_buf_o2_p,
    lo582_buf_o2
  );


  not

  (
    lo582_buf_o2_n,
    lo582_buf_o2
  );


  buf

  (
    lo030_buf_o2_p,
    lo030_buf_o2
  );


  not

  (
    lo030_buf_o2_n,
    lo030_buf_o2
  );


  buf

  (
    lo174_buf_o2_p,
    lo174_buf_o2
  );


  not

  (
    lo174_buf_o2_n,
    lo174_buf_o2
  );


  buf

  (
    lo178_buf_o2_p,
    lo178_buf_o2
  );


  not

  (
    lo178_buf_o2_n,
    lo178_buf_o2
  );


  buf

  (
    lo186_buf_o2_p,
    lo186_buf_o2
  );


  not

  (
    lo186_buf_o2_n,
    lo186_buf_o2
  );


  buf

  (
    lo266_buf_o2_p,
    lo266_buf_o2
  );


  not

  (
    lo266_buf_o2_n,
    lo266_buf_o2
  );


  buf

  (
    lo306_buf_o2_p,
    lo306_buf_o2
  );


  not

  (
    lo306_buf_o2_n,
    lo306_buf_o2
  );


  buf

  (
    lo346_buf_o2_p,
    lo346_buf_o2
  );


  not

  (
    lo346_buf_o2_n,
    lo346_buf_o2
  );


  buf

  (
    lo386_buf_o2_p,
    lo386_buf_o2
  );


  not

  (
    lo386_buf_o2_n,
    lo386_buf_o2
  );


  buf

  (
    lo426_buf_o2_p,
    lo426_buf_o2
  );


  not

  (
    lo426_buf_o2_n,
    lo426_buf_o2
  );


  buf

  (
    lo590_buf_o2_p,
    lo590_buf_o2
  );


  not

  (
    lo590_buf_o2_n,
    lo590_buf_o2
  );


  buf

  (
    lo594_buf_o2_p,
    lo594_buf_o2
  );


  not

  (
    lo594_buf_o2_n,
    lo594_buf_o2
  );


  buf

  (
    lo606_buf_o2_p,
    lo606_buf_o2
  );


  not

  (
    lo606_buf_o2_n,
    lo606_buf_o2
  );


  buf

  (
    lo610_buf_o2_p,
    lo610_buf_o2
  );


  not

  (
    lo610_buf_o2_n,
    lo610_buf_o2
  );


  buf

  (
    n2238_o2_p,
    n2238_o2
  );


  not

  (
    n2238_o2_n,
    n2238_o2
  );


  buf

  (
    n2229_o2_p,
    n2229_o2
  );


  not

  (
    n2229_o2_n,
    n2229_o2
  );


  buf

  (
    n2242_o2_p,
    n2242_o2
  );


  not

  (
    n2242_o2_n,
    n2242_o2
  );


  buf

  (
    n2233_o2_p,
    n2233_o2
  );


  not

  (
    n2233_o2_n,
    n2233_o2
  );


  buf

  (
    n2168_o2_p,
    n2168_o2
  );


  not

  (
    n2168_o2_n,
    n2168_o2
  );


  buf

  (
    n2237_o2_p,
    n2237_o2
  );


  not

  (
    n2237_o2_n,
    n2237_o2
  );


  buf

  (
    n2228_o2_p,
    n2228_o2
  );


  not

  (
    n2228_o2_n,
    n2228_o2
  );


  buf

  (
    n2172_o2_p,
    n2172_o2
  );


  not

  (
    n2172_o2_n,
    n2172_o2
  );


  buf

  (
    n2223_o2_p,
    n2223_o2
  );


  not

  (
    n2223_o2_n,
    n2223_o2
  );


  buf

  (
    n2222_o2_p,
    n2222_o2
  );


  not

  (
    n2222_o2_n,
    n2222_o2
  );


  buf

  (
    n2170_o2_p,
    n2170_o2
  );


  not

  (
    n2170_o2_n,
    n2170_o2
  );


  buf

  (
    n2181_o2_p,
    n2181_o2
  );


  not

  (
    n2181_o2_n,
    n2181_o2
  );


  buf

  (
    n2510_o2_p,
    n2510_o2
  );


  not

  (
    n2510_o2_n,
    n2510_o2
  );


  buf

  (
    n2621_o2_p,
    n2621_o2
  );


  not

  (
    n2621_o2_n,
    n2621_o2
  );


  buf

  (
    lo466_buf_o2_p,
    lo466_buf_o2
  );


  not

  (
    lo466_buf_o2_n,
    lo466_buf_o2
  );


  buf

  (
    lo478_buf_o2_p,
    lo478_buf_o2
  );


  not

  (
    lo478_buf_o2_n,
    lo478_buf_o2
  );


  buf

  (
    n2149_o2_p,
    n2149_o2
  );


  not

  (
    n2149_o2_n,
    n2149_o2
  );


  buf

  (
    n2429_o2_p,
    n2429_o2
  );


  not

  (
    n2429_o2_n,
    n2429_o2
  );


  buf

  (
    n2444_o2_p,
    n2444_o2
  );


  not

  (
    n2444_o2_n,
    n2444_o2
  );


  buf

  (
    n2153_o2_p,
    n2153_o2
  );


  not

  (
    n2153_o2_n,
    n2153_o2
  );


  buf

  (
    n2433_o2_p,
    n2433_o2
  );


  not

  (
    n2433_o2_n,
    n2433_o2
  );


  buf

  (
    n2448_o2_p,
    n2448_o2
  );


  not

  (
    n2448_o2_n,
    n2448_o2
  );


  buf

  (
    n2367_o2_p,
    n2367_o2
  );


  not

  (
    n2367_o2_n,
    n2367_o2
  );


  buf

  (
    n2386_o2_p,
    n2386_o2
  );


  not

  (
    n2386_o2_n,
    n2386_o2
  );


  buf

  (
    n2539_o2_p,
    n2539_o2
  );


  not

  (
    n2539_o2_n,
    n2539_o2
  );


  buf

  (
    n2183_o2_p,
    n2183_o2
  );


  not

  (
    n2183_o2_n,
    n2183_o2
  );


  buf

  (
    n2220_o2_p,
    n2220_o2
  );


  not

  (
    n2220_o2_n,
    n2220_o2
  );


  buf

  (
    n2514_o2_p,
    n2514_o2
  );


  not

  (
    n2514_o2_n,
    n2514_o2
  );


  buf

  (
    n2196_o2_p,
    n2196_o2
  );


  not

  (
    n2196_o2_n,
    n2196_o2
  );


  buf

  (
    n2616_o2_p,
    n2616_o2
  );


  not

  (
    n2616_o2_n,
    n2616_o2
  );


  buf

  (
    n2612_o2_p,
    n2612_o2
  );


  not

  (
    n2612_o2_n,
    n2612_o2
  );


  buf

  (
    n2627_o2_p,
    n2627_o2
  );


  not

  (
    n2627_o2_n,
    n2627_o2
  );


  buf

  (
    n2140_o2_p,
    n2140_o2
  );


  not

  (
    n2140_o2_n,
    n2140_o2
  );


  buf

  (
    n1877_inv_p,
    n1877_inv
  );


  not

  (
    n1877_inv_n,
    n1877_inv
  );


  buf

  (
    lo149_buf_o2_p,
    lo149_buf_o2
  );


  not

  (
    lo149_buf_o2_n,
    lo149_buf_o2
  );


  buf

  (
    lo197_buf_o2_p,
    lo197_buf_o2
  );


  not

  (
    lo197_buf_o2_n,
    lo197_buf_o2
  );


  buf

  (
    lo118_buf_o2_p,
    lo118_buf_o2
  );


  not

  (
    lo118_buf_o2_n,
    lo118_buf_o2
  );


  buf

  (
    lo158_buf_o2_p,
    lo158_buf_o2
  );


  not

  (
    lo158_buf_o2_n,
    lo158_buf_o2
  );


  buf

  (
    lo166_buf_o2_p,
    lo166_buf_o2
  );


  not

  (
    lo166_buf_o2_n,
    lo166_buf_o2
  );


  buf

  (
    lo242_buf_o2_p,
    lo242_buf_o2
  );


  not

  (
    lo242_buf_o2_n,
    lo242_buf_o2
  );


  buf

  (
    lo286_buf_o2_p,
    lo286_buf_o2
  );


  not

  (
    lo286_buf_o2_n,
    lo286_buf_o2
  );


  buf

  (
    lo506_buf_o2_p,
    lo506_buf_o2
  );


  not

  (
    lo506_buf_o2_n,
    lo506_buf_o2
  );


  buf

  (
    n2198_o2_p,
    n2198_o2
  );


  not

  (
    n2198_o2_n,
    n2198_o2
  );


  buf

  (
    n2202_o2_p,
    n2202_o2
  );


  not

  (
    n2202_o2_n,
    n2202_o2
  );


  buf

  (
    n2197_o2_p,
    n2197_o2
  );


  not

  (
    n2197_o2_n,
    n2197_o2
  );


  buf

  (
    n1913_inv_p,
    n1913_inv
  );


  not

  (
    n1913_inv_n,
    n1913_inv
  );


  buf

  (
    n2146_o2_p,
    n2146_o2
  );


  not

  (
    n2146_o2_n,
    n2146_o2
  );


  buf

  (
    n1919_inv_p,
    n1919_inv
  );


  not

  (
    n1919_inv_n,
    n1919_inv
  );


  buf

  (
    lo312_buf_o2_p,
    lo312_buf_o2
  );


  not

  (
    lo312_buf_o2_n,
    lo312_buf_o2
  );


  buf

  (
    lo316_buf_o2_p,
    lo316_buf_o2
  );


  not

  (
    lo316_buf_o2_n,
    lo316_buf_o2
  );


  buf

  (
    lo352_buf_o2_p,
    lo352_buf_o2
  );


  not

  (
    lo352_buf_o2_n,
    lo352_buf_o2
  );


  buf

  (
    lo356_buf_o2_p,
    lo356_buf_o2
  );


  not

  (
    lo356_buf_o2_n,
    lo356_buf_o2
  );


  buf

  (
    lo392_buf_o2_p,
    lo392_buf_o2
  );


  not

  (
    lo392_buf_o2_n,
    lo392_buf_o2
  );


  buf

  (
    lo396_buf_o2_p,
    lo396_buf_o2
  );


  not

  (
    lo396_buf_o2_n,
    lo396_buf_o2
  );


  buf

  (
    lo432_buf_o2_p,
    lo432_buf_o2
  );


  not

  (
    lo432_buf_o2_n,
    lo432_buf_o2
  );


  buf

  (
    lo436_buf_o2_p,
    lo436_buf_o2
  );


  not

  (
    lo436_buf_o2_n,
    lo436_buf_o2
  );


  buf

  (
    lo576_buf_o2_p,
    lo576_buf_o2
  );


  not

  (
    lo576_buf_o2_n,
    lo576_buf_o2
  );


  or

  (
    g733_n,
    n2118_o2_n,
    n2119_o2_n
  );


  or

  (
    g734_n,
    n1437_lo_n,
    n1545_lo_n
  );


  or

  (
    g735_n,
    n2865_lo_n_spl_,
    g734_n
  );


  and

  (
    g736_p,
    n2301_lo_p,
    n2793_lo_n_spl_0
  );


  or

  (
    g737_n,
    n1497_lo_n,
    n2865_lo_n_spl_
  );


  or

  (
    g738_n,
    n2841_lo_n,
    g737_n_spl_0
  );


  or

  (
    g739_n,
    n3177_lo_n,
    g737_n_spl_0
  );


  or

  (
    g740_n,
    n2127_o2_n,
    n2128_o2_n
  );


  or

  (
    g741_n,
    n2130_o2_n,
    n2131_o2_n
  );


  or

  (
    g742_n,
    g740_n_spl_,
    g741_n_spl_
  );


  and

  (
    g743_p,
    n3177_lo_p,
    g741_n_spl_
  );


  and

  (
    g744_p,
    n2841_lo_p,
    g740_n_spl_
  );


  or

  (
    g745_n,
    g743_p,
    g744_p
  );


  and

  (
    g746_p,
    n3603_o2_n,
    n3604_o2_n
  );


  and

  (
    g747_p,
    n2150_o2_n,
    n2154_o2_n
  );


  and

  (
    g748_p,
    n2167_o2_n,
    n2174_o2_n
  );


  or

  (
    g749_n,
    n2177_o2_p,
    n2184_o2_p
  );


  or

  (
    g750_n,
    n2877_lo_n_spl_0,
    n3798_o2_p
  );


  or

  (
    g751_n,
    n2805_lo_n,
    n2865_lo_p
  );


  or

  (
    g752_n,
    g745_n_spl_0,
    g751_n
  );


  or

  (
    g753_n,
    n1749_lo_n,
    g752_n_spl_
  );


  and

  (
    g754_p,
    n1425_lo_p,
    n1449_lo_p
  );


  or

  (
    g755_n,
    g752_n_spl_,
    g754_p
  );


  or

  (
    g756_n,
    n2889_lo_p_spl_0,
    n3846_o2_n_spl_
  );


  or

  (
    g757_n,
    n2889_lo_n_spl_0,
    n4019_o2_p_spl_
  );


  and

  (
    g758_p,
    g756_n,
    g757_n
  );


  and

  (
    g759_p,
    n2889_lo_n_spl_0,
    n4017_o2_n
  );


  and

  (
    g760_p,
    n2889_lo_p_spl_0,
    g749_n_spl_
  );


  or

  (
    g761_n,
    g759_p,
    g760_p
  );


  and

  (
    g762_p,
    n2829_lo_p_spl_,
    n2877_lo_n_spl_0
  );


  or

  (
    g763_n,
    n3846_o2_p_spl_,
    g762_p
  );


  or

  (
    g764_n,
    n2889_lo_p_spl_1,
    n3798_o2_n
  );


  or

  (
    g765_n,
    n2889_lo_n_spl_1,
    n2264_o2_n_spl_0
  );


  and

  (
    g766_p,
    g764_n,
    g765_n
  );


  or

  (
    g767_n,
    n3129_lo_p,
    n2275_o2_n
  );


  or

  (
    g768_n,
    n3129_lo_n,
    n2275_o2_p
  );


  and

  (
    g769_p,
    g767_n,
    g768_n
  );


  or

  (
    g770_n,
    n3141_lo_p,
    g769_p
  );


  or

  (
    g771_n,
    n2288_o2_n,
    n2303_o2_n
  );


  or

  (
    g772_n,
    n2288_o2_p,
    n2303_o2_p
  );


  and

  (
    g773_p,
    n1533_lo_p,
    g772_n
  );


  and

  (
    g774_p,
    g771_n,
    g773_p
  );


  and

  (
    g775_p,
    n2318_o2_n,
    n2319_o2_n
  );


  or

  (
    g775_n,
    n2318_o2_p,
    n2319_o2_p
  );


  and

  (
    g776_p,
    n2321_o2_n,
    n2322_o2_n
  );


  or

  (
    g776_n,
    n2321_o2_p,
    n2322_o2_p
  );


  or

  (
    g777_n,
    g775_n,
    g776_p
  );


  or

  (
    g778_n,
    g775_p,
    g776_n
  );


  and

  (
    g779_p,
    g777_n,
    g778_n
  );


  and

  (
    g780_p,
    n2329_o2_p_spl_,
    n2332_o2_n_spl_
  );


  or

  (
    g780_n,
    n2329_o2_n_spl_,
    n2332_o2_p_spl_
  );


  and

  (
    g781_p,
    n2329_o2_n_spl_,
    n2332_o2_p_spl_
  );


  or

  (
    g781_n,
    n2329_o2_p_spl_,
    n2332_o2_n_spl_
  );


  and

  (
    g782_p,
    g780_n,
    g781_n
  );


  or

  (
    g782_n,
    g780_p,
    g781_p
  );


  and

  (
    g783_p,
    n2347_o2_n_spl_,
    n2344_o2_p_spl_
  );


  or

  (
    g783_n,
    n2347_o2_p_spl_,
    n2344_o2_n_spl_
  );


  and

  (
    g784_p,
    n2347_o2_p_spl_,
    n2344_o2_n_spl_
  );


  or

  (
    g784_n,
    n2347_o2_n_spl_,
    n2344_o2_p_spl_
  );


  and

  (
    g785_p,
    g783_n,
    g784_n
  );


  or

  (
    g785_n,
    g783_p,
    g784_p
  );


  or

  (
    g786_n,
    g782_p,
    g785_n
  );


  or

  (
    g787_n,
    g782_n,
    g785_p
  );


  and

  (
    g788_p,
    g786_n,
    g787_n
  );


  and

  (
    g789_p,
    n3117_lo_n,
    n2356_o2_p
  );


  and

  (
    g790_p,
    n3081_lo_p,
    n2369_o2_n
  );


  and

  (
    g791_p,
    n2961_lo_n,
    n2373_o2_p
  );


  or

  (
    g792_n,
    g790_p,
    g791_p
  );


  or

  (
    g793_n,
    g789_p,
    g792_n
  );


  and

  (
    g794_p,
    n3033_lo_p,
    n2388_o2_n
  );


  and

  (
    g795_p,
    n3093_lo_n,
    n2392_o2_p
  );


  or

  (
    g796_n,
    g794_p,
    g795_p
  );


  and

  (
    g797_p,
    n3105_lo_p,
    n2397_o2_n
  );


  and

  (
    g798_p,
    n3033_lo_n,
    n2388_o2_p
  );


  or

  (
    g799_n,
    g797_p,
    g798_p
  );


  or

  (
    g800_n,
    g796_n,
    g799_n
  );


  and

  (
    g801_p,
    n2925_lo_n,
    n2404_o2_p
  );


  and

  (
    g802_p,
    n2961_lo_p,
    n2373_o2_n
  );


  or

  (
    g803_n,
    g801_p,
    g802_p
  );


  and

  (
    g804_p,
    n3021_lo_n,
    n2410_o2_p
  );


  and

  (
    g805_p,
    n3117_lo_p,
    n2356_o2_n
  );


  or

  (
    g806_n,
    g804_p,
    g805_p
  );


  or

  (
    g807_n,
    g803_n,
    g806_n
  );


  or

  (
    g808_n,
    g800_n,
    g807_n
  );


  or

  (
    g809_n,
    g793_n,
    g808_n
  );


  and

  (
    g810_p,
    n2997_lo_p,
    n2419_o2_n
  );


  and

  (
    g811_p,
    n2421_o2_n,
    n2422_o2_n
  );


  or

  (
    g812_n,
    n1521_lo_n,
    g811_p
  );


  or

  (
    g813_n,
    g810_p,
    g812_n
  );


  and

  (
    g814_p,
    n3069_lo_n,
    n2437_o2_p
  );


  and

  (
    g815_p,
    n3069_lo_p,
    n2437_o2_n
  );


  or

  (
    g816_n,
    g814_p,
    g815_p
  );


  and

  (
    g817_p,
    n3045_lo_p,
    n2452_o2_n
  );


  and

  (
    g818_p,
    n3045_lo_n,
    n2452_o2_p
  );


  or

  (
    g819_n,
    g817_p,
    g818_p
  );


  or

  (
    g820_n,
    g816_n,
    g819_n
  );


  or

  (
    g821_n,
    g813_n,
    g820_n
  );


  or

  (
    g822_n,
    n2458_o2_p,
    n2462_o2_p
  );


  or

  (
    g823_n,
    n2467_o2_p,
    n2468_o2_p
  );


  or

  (
    g824_n,
    g822_n,
    g823_n
  );


  or

  (
    g825_n,
    n2471_o2_p,
    n2472_o2_p
  );


  or

  (
    g826_n,
    n2478_o2_p,
    n2474_o2_p
  );


  or

  (
    g827_n,
    g825_n,
    g826_n
  );


  or

  (
    g828_n,
    g824_n,
    g827_n
  );


  or

  (
    g829_n,
    n2486_o2_p,
    n2485_o2_p
  );


  or

  (
    g830_n,
    n2488_o2_p,
    n2489_o2_p
  );


  or

  (
    g831_n,
    g829_n,
    g830_n
  );


  or

  (
    g832_n,
    n2495_o2_p,
    n2496_o2_p
  );


  or

  (
    g833_n,
    n2498_o2_p,
    n2499_o2_p
  );


  or

  (
    g834_n,
    g832_n,
    g833_n
  );


  or

  (
    g835_n,
    g831_n,
    g834_n
  );


  or

  (
    g836_n,
    g828_n,
    g835_n
  );


  or

  (
    g837_n,
    g821_n,
    g836_n
  );


  or

  (
    g838_n,
    g809_n,
    g837_n
  );


  and

  (
    g839_p,
    n2829_lo_p_spl_,
    n3846_o2_n_spl_
  );


  or

  (
    g839_n,
    n2829_lo_n,
    n3846_o2_p_spl_
  );


  and

  (
    g840_p,
    n2518_o2_n,
    g839_p
  );


  and

  (
    g841_p,
    n2518_o2_p,
    g839_n
  );


  or

  (
    g842_n,
    g840_p,
    g841_p
  );


  and

  (
    g843_p,
    n2877_lo_n_spl_,
    g842_n
  );


  and

  (
    g844_p,
    n2877_lo_p,
    n2515_o2_p_spl_
  );


  or

  (
    g845_n,
    g843_p,
    g844_p
  );


  or

  (
    g846_n,
    n2530_o2_p,
    n2554_o2_p
  );


  or

  (
    g847_n,
    n2530_o2_n,
    n2554_o2_n
  );


  and

  (
    g848_p,
    n1761_lo_n_spl_,
    g847_n
  );


  and

  (
    g849_p,
    g846_n,
    g848_p
  );


  or

  (
    g850_n,
    n2889_lo_p_spl_1,
    n2515_o2_p_spl_
  );


  and

  (
    g851_p,
    n2566_o2_n,
    n2567_o2_n
  );


  or

  (
    g851_n,
    n2566_o2_p,
    n2567_o2_p
  );


  and

  (
    g852_p,
    n2574_o2_n_spl_,
    n2264_o2_p_spl_
  );


  or

  (
    g852_n,
    n2574_o2_p_spl_,
    n2264_o2_n_spl_0
  );


  and

  (
    g853_p,
    n2574_o2_p_spl_,
    n2264_o2_n_spl_
  );


  or

  (
    g853_n,
    n2574_o2_n_spl_,
    n2264_o2_p_spl_
  );


  and

  (
    g854_p,
    g852_n,
    g853_n
  );


  or

  (
    g854_n,
    g852_p,
    g853_p
  );


  or

  (
    g855_n,
    g851_p_spl_,
    g854_p
  );


  or

  (
    g856_n,
    g851_n_spl_,
    g854_n
  );


  and

  (
    g857_p,
    g855_n,
    g856_n
  );


  or

  (
    g858_n,
    n2889_lo_n_spl_1,
    g857_p
  );


  and

  (
    g859_p,
    g850_n,
    g858_n
  );


  and

  (
    g860_p,
    n2586_o2_p,
    n2587_o2_n
  );


  or

  (
    g860_n,
    n2586_o2_n,
    n2587_o2_p
  );


  or

  (
    g861_n,
    g851_p_spl_,
    g860_n
  );


  or

  (
    g862_n,
    g851_n_spl_,
    g860_p
  );


  and

  (
    g863_p,
    n1761_lo_n_spl_,
    g862_n
  );


  and

  (
    g864_p,
    g861_n,
    g863_p
  );


  or

  (
    g865_n,
    n2593_o2_p,
    n2601_o2_n
  );


  or

  (
    g866_n,
    n2603_o2_p,
    n2636_o2_p
  );


  and

  (
    g867_p,
    g865_n,
    g866_n
  );


  or

  (
    g868_n,
    n2639_o2_p,
    n2640_o2_p
  );


  or

  (
    g869_n,
    n2643_o2_p,
    n2642_o2_p
  );


  or

  (
    g870_n,
    g868_n_spl_,
    g869_n
  );


  or

  (
    g871_n,
    g867_p,
    g870_n
  );


  or

  (
    g872_n,
    n2643_o2_n,
    g868_n_spl_
  );


  and

  (
    g873_p,
    n2639_o2_n,
    g872_n
  );


  and

  (
    g874_p,
    g871_n,
    g873_p
  );


  or

  (
    g875_n,
    n2653_o2_p,
    n2654_o2_p
  );


  or

  (
    g876_n,
    n2660_o2_p_spl_,
    g875_n_spl_
  );


  or

  (
    g877_n,
    n2664_o2_p,
    n2665_o2_p
  );


  and

  (
    g878_p,
    n2668_o2_n,
    n2667_o2_p
  );


  or

  (
    g879_n,
    n2669_o2_p,
    g878_p
  );


  or

  (
    g880_n,
    g877_n_spl_,
    g879_n
  );


  or

  (
    g881_n,
    g876_n_spl_,
    g880_n
  );


  or

  (
    g882_n,
    g874_p,
    g881_n
  );


  or

  (
    g883_n,
    n2669_o2_n,
    n2660_o2_p_spl_
  );


  or

  (
    g884_n,
    g877_n_spl_,
    g883_n
  );


  and

  (
    g885_p,
    n2658_o2_n,
    g884_n
  );


  or

  (
    g886_n,
    g875_n_spl_,
    g885_p
  );


  or

  (
    g887_n,
    n2664_o2_n,
    g876_n_spl_
  );


  and

  (
    g888_p,
    n2653_o2_n,
    g887_n
  );


  and

  (
    g889_p,
    g886_n,
    g888_p
  );


  and

  (
    g890_p,
    g882_n,
    g889_p
  );


  or

  (
    g891_n,
    g774_p_spl_,
    g779_p_spl_
  );


  or

  (
    g892_n,
    g788_p_spl_,
    g891_n
  );


  or

  (
    g893_n,
    g745_n_spl_0,
    g849_p_spl_
  );


  or

  (
    g894_n,
    g864_p_spl_,
    g893_n
  );


  or

  (
    g895_n,
    g892_n,
    g894_n
  );


  and

  (
    g896_p,
    n4038_o2_p_spl_0,
    lo186_buf_o2_p
  );


  or

  (
    g896_n,
    n4038_o2_n_spl_0,
    lo186_buf_o2_n
  );


  and

  (
    g897_p,
    n3964_o2_p_spl_00,
    n2149_o2_p
  );


  or

  (
    g897_n,
    n3964_o2_n_spl_00,
    n2149_o2_n
  );


  and

  (
    g898_p,
    n3964_o2_n_spl_00,
    n2153_o2_p
  );


  or

  (
    g898_n,
    n3964_o2_p_spl_00,
    n2153_o2_n
  );


  and

  (
    g899_p,
    n2181_o2_p,
    n2183_o2_n
  );


  or

  (
    g899_n,
    n2181_o2_n,
    n2183_o2_p
  );


  and

  (
    g900_p,
    n2510_o2_n,
    n2514_o2_n
  );


  or

  (
    g900_n,
    n2510_o2_p,
    n2514_o2_p
  );


  and

  (
    g901_p,
    n1962_lo_p,
    n4038_o2_p_spl_0
  );


  or

  (
    g901_n,
    n1962_lo_n,
    n4038_o2_n_spl_0
  );


  and

  (
    g902_p,
    lo554_buf_o2_p_spl_0,
    lo558_buf_o2_p_spl_0
  );


  or

  (
    g902_n,
    lo554_buf_o2_n_spl_0,
    lo558_buf_o2_n_spl_0
  );


  and

  (
    g903_p,
    g896_n,
    g899_n
  );


  or

  (
    g903_n,
    g896_p_spl_,
    g899_p_spl_
  );


  and

  (
    g904_p,
    n4006_o2_n_spl_00,
    n2168_o2_n
  );


  or

  (
    g904_n,
    n4006_o2_p_spl_00,
    n2168_o2_p
  );


  and

  (
    g905_p,
    n2172_o2_n,
    n2170_o2_n
  );


  or

  (
    g905_n,
    n2172_o2_p,
    n2170_o2_p
  );


  and

  (
    g906_p,
    g904_n,
    g905_p
  );


  or

  (
    g906_n,
    g904_p,
    g905_n
  );


  and

  (
    g907_p,
    n2187_o2_n,
    n2194_o2_n
  );


  or

  (
    g907_n,
    n2187_o2_p,
    n2194_o2_p
  );


  and

  (
    g908_p,
    g901_n,
    g906_n
  );


  or

  (
    g908_n,
    g901_p_spl_,
    g906_p_spl_
  );


  and

  (
    g909_p,
    n2223_o2_n,
    n2222_o2_p
  );


  or

  (
    g909_n,
    n2223_o2_p,
    n2222_o2_n
  );


  and

  (
    g910_p,
    n4005_o2_n_spl_,
    g909_n
  );


  or

  (
    g910_n,
    n4005_o2_p_spl_,
    g909_p
  );


  and

  (
    g911_p,
    n4006_o2_p_spl_00,
    lo266_buf_o2_n
  );


  or

  (
    g911_n,
    n4006_o2_n_spl_00,
    lo266_buf_o2_p
  );


  and

  (
    g912_p,
    n4005_o2_p_spl_,
    g911_p
  );


  or

  (
    g912_n,
    n4005_o2_n_spl_,
    g911_n
  );


  and

  (
    g913_p,
    g910_n,
    g912_n
  );


  or

  (
    g913_n,
    g910_p,
    g912_p
  );


  and

  (
    g914_p,
    n2229_o2_n,
    n2228_o2_n
  );


  or

  (
    g914_n,
    n2229_o2_p,
    n2228_o2_p
  );


  and

  (
    g915_p,
    n4006_o2_p_spl_01,
    g914_n
  );


  or

  (
    g915_n,
    n4006_o2_n_spl_01,
    g914_p
  );


  and

  (
    g916_p,
    n4038_o2_p_spl_1,
    lo178_buf_o2_p
  );


  or

  (
    g916_n,
    n4038_o2_n_spl_1,
    lo178_buf_o2_n
  );


  and

  (
    g917_p,
    n4006_o2_n_spl_01,
    n2233_o2_p
  );


  or

  (
    g917_n,
    n4006_o2_p_spl_01,
    n2233_o2_n
  );


  and

  (
    g918_p,
    g916_n,
    g917_n
  );


  or

  (
    g918_n,
    g916_p,
    g917_p
  );


  and

  (
    g919_p,
    g915_n,
    g918_p
  );


  or

  (
    g919_n,
    g915_p,
    g918_n
  );


  and

  (
    g920_p,
    n2238_o2_n,
    n2237_o2_n
  );


  or

  (
    g920_n,
    n2238_o2_p,
    n2237_o2_p
  );


  and

  (
    g921_p,
    n4006_o2_p_spl_1,
    g920_n
  );


  or

  (
    g921_n,
    n4006_o2_n_spl_1,
    g920_p
  );


  and

  (
    g922_p,
    n4038_o2_p_spl_1,
    lo174_buf_o2_p
  );


  or

  (
    g922_n,
    n4038_o2_n_spl_1,
    lo174_buf_o2_n
  );


  and

  (
    g923_p,
    n4006_o2_n_spl_1,
    n2242_o2_p
  );


  or

  (
    g923_n,
    n4006_o2_p_spl_1,
    n2242_o2_n
  );


  and

  (
    g924_p,
    g922_n,
    g923_n
  );


  or

  (
    g924_n,
    g922_p,
    g923_p
  );


  and

  (
    g925_p,
    g921_n,
    g924_p
  );


  or

  (
    g925_n,
    g921_p,
    g924_n
  );


  and

  (
    g926_p,
    n2205_o2_n_spl_,
    g900_n_spl_0
  );


  or

  (
    g926_n,
    n2205_o2_p_spl_0,
    g900_p_spl_
  );


  and

  (
    g927_p,
    n2205_o2_p_spl_0,
    g900_p_spl_
  );


  or

  (
    g927_n,
    n2205_o2_n_spl_,
    g900_n_spl_0
  );


  and

  (
    g928_p,
    g926_n,
    g927_n
  );


  or

  (
    g928_n,
    g926_p,
    g927_p
  );


  or

  (
    g929_n,
    n3102_lo_n_spl_0,
    n3114_lo_n_spl_
  );


  and

  (
    g930_p,
    n3837_o2_n_spl_0,
    lo306_buf_o2_p
  );


  or

  (
    g930_n,
    n3837_o2_p_spl_0,
    lo306_buf_o2_n
  );


  and

  (
    g931_p,
    n3837_o2_p_spl_0,
    lo426_buf_o2_p
  );


  or

  (
    g931_n,
    n3837_o2_n_spl_0,
    lo426_buf_o2_n
  );


  and

  (
    g932_p,
    g930_n,
    g931_n
  );


  or

  (
    g932_n,
    g930_p,
    g931_p
  );


  and

  (
    g933_p,
    n3964_o2_p_spl_01,
    g932_n
  );


  or

  (
    g933_n,
    n3964_o2_n_spl_01,
    g932_p
  );


  and

  (
    g934_p,
    n3837_o2_n_spl_1,
    lo346_buf_o2_p
  );


  or

  (
    g934_n,
    n3837_o2_p_spl_1,
    lo346_buf_o2_n
  );


  and

  (
    g935_p,
    n3837_o2_p_spl_1,
    lo386_buf_o2_p
  );


  or

  (
    g935_n,
    n3837_o2_n_spl_1,
    lo386_buf_o2_n
  );


  and

  (
    g936_p,
    g934_n,
    g935_n
  );


  or

  (
    g936_n,
    g934_p,
    g935_p
  );


  and

  (
    g937_p,
    n3964_o2_n_spl_01,
    g936_n
  );


  or

  (
    g937_n,
    n3964_o2_p_spl_01,
    g936_p
  );


  and

  (
    g938_p,
    g933_n,
    g937_n
  );


  or

  (
    g938_n,
    g933_p,
    g937_p
  );


  and

  (
    g939_p,
    lo118_buf_o2_p,
    n2146_o2_n
  );


  or

  (
    g939_n,
    lo118_buf_o2_n,
    n2146_o2_p_spl_
  );


  and

  (
    g940_p,
    lo506_buf_o2_n,
    n1919_inv_p_spl_
  );


  or

  (
    g940_n,
    lo506_buf_o2_p,
    n1919_inv_n
  );


  and

  (
    g941_p,
    g939_p_spl_,
    g940_p_spl_
  );


  or

  (
    g941_n,
    g939_n,
    g940_n
  );


  or

  (
    g942_n,
    lo030_buf_o2_n_spl_,
    g908_n_spl_0
  );


  and

  (
    g943_p,
    n2595_o2_p,
    n2594_o2_n
  );


  or

  (
    g943_n,
    n2595_o2_n,
    n2594_o2_p
  );


  or

  (
    g944_n,
    n3018_lo_p_spl_0,
    g943_n_spl_00
  );


  and

  (
    g945_p,
    g925_p_spl_,
    g943_p_spl_00
  );


  and

  (
    g946_p,
    n1458_lo_p,
    n1554_lo_p_spl_000
  );


  and

  (
    g947_p,
    n1554_lo_n_spl_000,
    n2254_o2_p_spl_00
  );


  or

  (
    g948_n,
    g946_p,
    g947_p
  );


  and

  (
    g949_p,
    n1554_lo_p_spl_000,
    n1626_lo_p
  );


  and

  (
    g950_p,
    n1554_lo_n_spl_000,
    g925_n_spl_0
  );


  or

  (
    g951_n,
    g949_p,
    g950_p
  );


  and

  (
    g952_p,
    n1554_lo_p_spl_00,
    n1614_lo_p
  );


  and

  (
    g953_p,
    n1554_lo_n_spl_00,
    g913_p_spl_0
  );


  or

  (
    g954_n,
    g952_p,
    g953_p
  );


  and

  (
    g955_p,
    n1662_lo_p,
    n1686_lo_p_spl_00
  );


  and

  (
    g956_p,
    n1686_lo_n_spl_00,
    n1475_inv_p_spl_0
  );


  or

  (
    g957_n,
    g955_p,
    g956_p
  );


  and

  (
    g958_p,
    n1686_lo_p_spl_00,
    n1710_lo_p
  );


  and

  (
    g959_p,
    n1686_lo_n_spl_00,
    n2367_o2_p_spl_0
  );


  or

  (
    g960_n,
    g958_p,
    g959_p
  );


  and

  (
    g961_p,
    n1686_lo_p_spl_01,
    n1722_lo_p
  );


  and

  (
    g962_p,
    n1686_lo_n_spl_01,
    n4039_o2_p_spl_0
  );


  or

  (
    g963_n,
    g961_p,
    g962_p
  );


  and

  (
    g964_p,
    n2596_o2_n,
    lo030_buf_o2_p_spl_
  );


  and

  (
    g965_p,
    n2982_lo_n_spl_00,
    g964_p_spl_0
  );


  and

  (
    g966_p,
    n2596_o2_p,
    lo030_buf_o2_p_spl_
  );


  and

  (
    g967_p,
    n3114_lo_n_spl_,
    g966_p_spl_0
  );


  or

  (
    g968_n,
    g965_p,
    g967_p
  );


  and

  (
    g969_p,
    n3964_o2_p_spl_10,
    n2444_o2_p
  );


  or

  (
    g969_n,
    n3964_o2_n_spl_10,
    n2444_o2_n
  );


  and

  (
    g970_p,
    n3964_o2_n_spl_10,
    n2448_o2_p
  );


  or

  (
    g970_n,
    n3964_o2_p_spl_10,
    n2448_o2_n
  );


  and

  (
    g971_p,
    g969_n,
    g970_n
  );


  or

  (
    g971_n,
    g969_p,
    g970_p
  );


  and

  (
    g972_p,
    g943_p_spl_00,
    g971_n_spl_0
  );


  or

  (
    g972_n,
    g943_n_spl_00,
    g971_p_spl_0
  );


  and

  (
    g973_p,
    lo542_buf_o2_n_spl_,
    g943_p_spl_0
  );


  or

  (
    g973_n,
    lo542_buf_o2_p_spl_0,
    g943_n_spl_0
  );


  or

  (
    g974_n,
    g972_p,
    g973_n
  );


  and

  (
    g975_p,
    n2254_o2_p_spl_00,
    n2220_o2_p_spl_00
  );


  or

  (
    g975_n,
    n2254_o2_n_spl_,
    n2220_o2_n_spl_
  );


  and

  (
    g976_p,
    n2254_o2_n_spl_,
    n2220_o2_n_spl_
  );


  or

  (
    g976_n,
    n2254_o2_p_spl_0,
    n2220_o2_p_spl_00
  );


  and

  (
    g977_p,
    g975_n,
    g976_n
  );


  or

  (
    g977_n,
    g975_p,
    g976_p
  );


  and

  (
    g978_p,
    g928_n_spl_,
    g977_p
  );


  and

  (
    g979_p,
    g928_p,
    g977_n
  );


  or

  (
    g980_n,
    g978_p,
    g979_p
  );


  or

  (
    g981_n,
    n2198_o2_p,
    n2197_o2_p
  );


  and

  (
    g982_p,
    lo478_buf_o2_p_spl_000,
    g981_n
  );


  and

  (
    g983_p,
    lo166_buf_o2_p,
    n1913_inv_p_spl_00
  );


  and

  (
    g984_p,
    lo478_buf_o2_n_spl_00,
    n2202_o2_p
  );


  or

  (
    g985_n,
    g983_p,
    g984_p
  );


  or

  (
    g986_n,
    g982_p,
    g985_n
  );


  and

  (
    g987_p,
    lo466_buf_o2_p_spl_000,
    lo286_buf_o2_p
  );


  and

  (
    g988_p,
    lo466_buf_o2_n_spl_000,
    lo158_buf_o2_p
  );


  or

  (
    g989_n,
    g987_p,
    g988_p
  );


  and

  (
    g990_p,
    lo478_buf_o2_p_spl_000,
    g989_n
  );


  and

  (
    g991_p,
    lo197_buf_o2_p,
    n1913_inv_p_spl_00
  );


  and

  (
    g992_p,
    lo466_buf_o2_n_spl_000,
    lo242_buf_o2_p
  );


  and

  (
    g993_p,
    lo478_buf_o2_n_spl_00,
    g992_p
  );


  or

  (
    g994_n,
    g991_p,
    g993_p
  );


  or

  (
    g995_n,
    g990_p,
    g994_n
  );


  and

  (
    g996_p,
    n1674_lo_p,
    n1686_lo_p_spl_01
  );


  and

  (
    g997_p,
    n1686_lo_n_spl_01,
    g938_n_spl_0
  );


  and

  (
    g998_p,
    n1794_lo_p_spl_,
    n2178_lo_p_spl_
  );


  and

  (
    g999_p,
    n1926_lo_p_spl_,
    n2046_lo_p_spl_
  );


  and

  (
    g1000_p,
    n2322_lo_p_spl_,
    n2682_lo_p_spl_
  );


  and

  (
    g1001_p,
    n2442_lo_p_spl_,
    n2562_lo_p_spl_
  );


  or

  (
    g1002_n,
    n2826_lo_p_spl_,
    n2254_o2_p_spl_1
  );


  and

  (
    g1003_p,
    n1554_lo_p_spl_01,
    n1566_lo_p
  );


  and

  (
    g1004_p,
    n1554_lo_n_spl_01,
    n2205_o2_p_spl_1
  );


  or

  (
    g1005_n,
    g1003_p,
    g1004_p
  );


  or

  (
    g1006_n,
    lo498_buf_o2_n_spl_0,
    g1005_n_spl_
  );


  and

  (
    g1007_p,
    lo498_buf_o2_n_spl_0,
    g1005_n_spl_
  );


  or

  (
    g1008_n,
    lo502_buf_o2_n_spl_0,
    g948_n_spl_
  );


  and

  (
    g1009_p,
    n1554_lo_p_spl_01,
    n1578_lo_p
  );


  and

  (
    g1010_p,
    n1554_lo_n_spl_01,
    n2220_o2_p_spl_01
  );


  or

  (
    g1011_n,
    g1009_p,
    g1010_p
  );


  or

  (
    g1012_n,
    lo510_buf_o2_n_spl_0,
    g1011_n_spl_
  );


  and

  (
    g1013_p,
    lo510_buf_o2_n_spl_0,
    g1011_n_spl_
  );


  and

  (
    g1014_p,
    n1554_lo_p_spl_10,
    n1590_lo_p
  );


  and

  (
    g1015_p,
    n1554_lo_n_spl_10,
    g903_n_spl_0
  );


  or

  (
    g1016_n,
    g1014_p,
    g1015_p
  );


  and

  (
    g1017_p,
    n2970_lo_n_spl_0,
    g1016_n_spl_
  );


  or

  (
    g1018_n,
    n2970_lo_n_spl_0,
    g1016_n_spl_
  );


  and

  (
    g1019_p,
    n1554_lo_p_spl_10,
    n1602_lo_p
  );


  and

  (
    g1020_p,
    n1554_lo_n_spl_10,
    g908_n_spl_0
  );


  or

  (
    g1021_n,
    g1019_p,
    g1020_p
  );


  and

  (
    g1022_p,
    n2982_lo_n_spl_00,
    g1021_n_spl_
  );


  or

  (
    g1023_n,
    n2982_lo_n_spl_0,
    g1021_n_spl_
  );


  and

  (
    g1024_p,
    n2994_lo_n_spl_0,
    g954_n_spl_
  );


  and

  (
    g1025_p,
    n2994_lo_n_spl_0,
    g964_p_spl_0
  );


  and

  (
    g1026_p,
    n1482_lo_p,
    n1554_lo_p_spl_11
  );


  and

  (
    g1027_p,
    n1554_lo_n_spl_11,
    g919_n_spl_0
  );


  or

  (
    g1028_n,
    g1026_p,
    g1027_p
  );


  and

  (
    g1029_p,
    n3006_lo_n_spl_0,
    g1028_n_spl_
  );


  or

  (
    g1030_n,
    n3006_lo_n_spl_0,
    g1028_n_spl_
  );


  and

  (
    g1031_p,
    n3006_lo_n_spl_1,
    g964_p_spl_1
  );


  or

  (
    g1032_n,
    n3018_lo_n_spl_,
    g951_n_spl_
  );


  and

  (
    g1033_p,
    lo554_buf_o2_n_spl_0,
    g960_n_spl_
  );


  or

  (
    g1034_n,
    lo558_buf_o2_n_spl_0,
    g957_n_spl_
  );


  and

  (
    g1035_p,
    n3102_lo_n_spl_0,
    g963_n_spl_
  );


  and

  (
    g1036_p,
    n3126_lo_p_spl_,
    n3138_lo_n
  );


  and

  (
    g1037_p,
    n3126_lo_n,
    n3138_lo_p_spl_
  );


  and

  (
    g1038_p,
    g919_p_spl_,
    g966_p_spl_0
  );


  and

  (
    g1039_p,
    g913_n_spl_,
    g966_p_spl_1
  );


  or

  (
    g1040_n,
    n1983_lo_n,
    n1913_inv_n
  );


  and

  (
    g1041_p,
    n1470_lo_p,
    n1554_lo_p_spl_11
  );


  and

  (
    g1042_p,
    n1554_lo_n_spl_11,
    n2196_o2_p_spl_0
  );


  or

  (
    g1043_n,
    g1041_p,
    g1042_p
  );


  or

  (
    g1044_n,
    g942_n_spl_,
    g968_n_spl_
  );


  and

  (
    g1045_p,
    n1638_lo_p,
    n1686_lo_p_spl_10
  );


  and

  (
    g1046_p,
    n1686_lo_n_spl_10,
    n2386_o2_p_spl_0
  );


  or

  (
    g1047_n,
    g1045_p,
    g1046_p
  );


  and

  (
    g1048_p,
    n1650_lo_p,
    n1686_lo_p_spl_10
  );


  and

  (
    g1049_p,
    n3964_o2_p_spl_11,
    n2429_o2_p
  );


  or

  (
    g1049_n,
    n3964_o2_n_spl_11,
    n2429_o2_n
  );


  and

  (
    g1050_p,
    n3964_o2_n_spl_11,
    n2433_o2_p
  );


  or

  (
    g1050_n,
    n3964_o2_p_spl_11,
    n2433_o2_n
  );


  and

  (
    g1051_p,
    g1049_n,
    g1050_n
  );


  or

  (
    g1051_n,
    g1049_p,
    g1050_p
  );


  and

  (
    g1052_p,
    n1686_lo_n_spl_10,
    g1051_n_spl_0
  );


  or

  (
    g1053_n,
    g1048_p,
    g1052_p
  );


  and

  (
    g1054_p,
    n1686_lo_p_spl_11,
    n1734_lo_p
  );


  and

  (
    g1055_p,
    g897_n,
    g898_n
  );


  or

  (
    g1055_n,
    g897_p_spl_,
    g898_p_spl_
  );


  and

  (
    g1056_p,
    n1686_lo_n_spl_11,
    g1055_n_spl_0
  );


  or

  (
    g1057_n,
    g1054_p,
    g1056_p
  );


  and

  (
    g1058_p,
    n1686_lo_p_spl_11,
    n1698_lo_p
  );


  and

  (
    g1059_p,
    n1686_lo_n_spl_11,
    g971_n_spl_0
  );


  or

  (
    g1060_n,
    g1058_p,
    g1059_p
  );


  and

  (
    g1061_p,
    n2970_lo_n_spl_1,
    lo514_buf_o2_p_spl_
  );


  and

  (
    g1062_p,
    n2970_lo_p,
    lo514_buf_o2_n
  );


  or

  (
    g1063_n,
    g1061_p,
    g1062_p
  );


  and

  (
    g1064_p,
    n3006_lo_p,
    n3018_lo_n_spl_
  );


  and

  (
    g1065_p,
    n3006_lo_n_spl_1,
    n3018_lo_p_spl_0
  );


  or

  (
    g1066_n,
    g1064_p,
    g1065_p
  );


  or

  (
    g1067_n,
    g944_n_spl_,
    g945_p_spl_
  );


  and

  (
    g1068_p,
    n3030_lo_p_spl_,
    lo542_buf_o2_n_spl_
  );


  and

  (
    g1069_p,
    n3030_lo_n_spl_,
    lo542_buf_o2_p_spl_0
  );


  or

  (
    g1070_n,
    g1068_p,
    g1069_p
  );


  or

  (
    g1071_n,
    n2386_o2_n_spl_0,
    g943_n_spl_1
  );


  and

  (
    g1072_p,
    n3030_lo_n_spl_,
    g943_p_spl_1
  );


  and

  (
    g1073_p,
    g1071_n_spl_,
    g1072_p_spl_
  );


  or

  (
    g1074_n,
    g1071_n_spl_,
    g1072_p_spl_
  );


  or

  (
    g1075_n,
    g943_n_spl_1,
    g1051_n_spl_0
  );


  and

  (
    g1076_p,
    lo550_buf_o2_n_spl_0,
    g943_p_spl_1
  );


  and

  (
    g1077_p,
    g1075_n_spl_,
    g1076_p_spl_
  );


  or

  (
    g1078_n,
    g1075_n_spl_,
    g1076_p_spl_
  );


  or

  (
    g1079_n,
    lo030_buf_o2_n_spl_,
    g903_n_spl_0
  );


  and

  (
    g1080_p,
    n2970_lo_n_spl_1,
    g964_p_spl_1
  );


  and

  (
    g1081_p,
    n3102_lo_n_spl_,
    g966_p_spl_1
  );


  or

  (
    g1082_n,
    g1080_p,
    g1081_p
  );


  and

  (
    g1083_p,
    g1079_n_spl_,
    g1082_n_spl_
  );


  or

  (
    g1084_n,
    g1079_n_spl_,
    g1082_n_spl_
  );


  and

  (
    g1085_p,
    n2196_o2_p_spl_0,
    n2612_o2_n_spl_
  );


  and

  (
    g1086_p,
    n2220_o2_p_spl_01,
    n2616_o2_n_spl_
  );


  and

  (
    g1087_p,
    n2621_o2_n,
    n2627_o2_n
  );


  or

  (
    g1088_n,
    g1086_p,
    g1087_p
  );


  or

  (
    g1089_n,
    n2196_o2_p_spl_1,
    n2612_o2_n_spl_
  );


  or

  (
    g1090_n,
    n2220_o2_p_spl_1,
    n2616_o2_n_spl_
  );


  and

  (
    g1091_p,
    g1089_n,
    g1090_n
  );


  and

  (
    g1092_p,
    g1088_n,
    g1091_p
  );


  or

  (
    g1093_n,
    g1085_p,
    g1092_p
  );


  and

  (
    g1094_p,
    g1084_n,
    g1093_n
  );


  or

  (
    g1095_n,
    g1083_p,
    g1094_p
  );


  or

  (
    g1096_n,
    g972_n,
    g973_p
  );


  and

  (
    g1097_p,
    g974_n_spl_,
    g1096_n
  );


  or

  (
    g1098_n,
    n3102_lo_p_spl_,
    n3114_lo_p_spl_
  );


  and

  (
    g1099_p,
    g929_n_spl_,
    g1098_n
  );


  and

  (
    g1100_p,
    lo554_buf_o2_n_spl_,
    lo558_buf_o2_n_spl_
  );


  or

  (
    g1100_n,
    lo554_buf_o2_p_spl_0,
    lo558_buf_o2_p_spl_0
  );


  and

  (
    g1101_p,
    g902_n,
    g1100_n
  );


  or

  (
    g1101_n,
    g902_p_spl_,
    g1100_p
  );


  and

  (
    g1102_p,
    n3294_lo_n_spl_,
    lo550_buf_o2_n_spl_0
  );


  or

  (
    g1102_n,
    n3294_lo_p_spl_,
    lo550_buf_o2_p_spl_0
  );


  and

  (
    g1103_p,
    n3294_lo_p_spl_,
    lo550_buf_o2_p_spl_0
  );


  or

  (
    g1103_n,
    n3294_lo_n_spl_,
    lo550_buf_o2_n_spl_
  );


  and

  (
    g1104_p,
    g1102_n,
    g1103_n
  );


  or

  (
    g1104_n,
    g1102_p,
    g1103_p
  );


  or

  (
    g1105_n,
    g1101_p,
    g1104_n
  );


  or

  (
    g1106_n,
    g1101_n,
    g1104_p
  );


  and

  (
    g1107_p,
    g1105_n,
    g1106_n
  );


  or

  (
    g1108_n,
    g1099_p_spl_,
    g1107_p_spl_
  );


  and

  (
    g1109_p,
    g1099_p_spl_,
    g1107_p_spl_
  );


  and

  (
    g1110_p,
    g903_n_spl_1,
    g907_n_spl_
  );


  and

  (
    g1111_p,
    g903_p,
    g907_p
  );


  or

  (
    g1112_n,
    g1110_p,
    g1111_p
  );


  and

  (
    g1113_p,
    g980_n_spl_0,
    g1112_n_spl_
  );


  or

  (
    g1114_n,
    g980_n_spl_0,
    g1112_n_spl_
  );


  and

  (
    g1115_p,
    n3258_lo_p_spl_,
    n3270_lo_n_spl_
  );


  or

  (
    g1115_n,
    n3258_lo_n_spl_,
    n3270_lo_p_spl_
  );


  and

  (
    g1116_p,
    n3258_lo_n_spl_,
    n3270_lo_p_spl_
  );


  or

  (
    g1116_n,
    n3258_lo_p_spl_,
    n3270_lo_n_spl_
  );


  and

  (
    g1117_p,
    g1115_n,
    g1116_n
  );


  or

  (
    g1117_n,
    g1115_p,
    g1116_p
  );


  and

  (
    g1118_p,
    lo498_buf_o2_p_spl_,
    lo502_buf_o2_n_spl_0
  );


  or

  (
    g1118_n,
    lo498_buf_o2_n_spl_1,
    lo502_buf_o2_p_spl_0
  );


  and

  (
    g1119_p,
    lo498_buf_o2_n_spl_1,
    lo502_buf_o2_p_spl_0
  );


  or

  (
    g1119_n,
    lo498_buf_o2_p_spl_,
    lo502_buf_o2_n_spl_
  );


  and

  (
    g1120_p,
    g1118_n,
    g1119_n
  );


  or

  (
    g1120_n,
    g1118_p,
    g1119_p
  );


  and

  (
    g1121_p,
    g1117_n,
    g1120_p
  );


  and

  (
    g1122_p,
    g1117_p,
    g1120_n
  );


  or

  (
    g1123_n,
    g1121_p,
    g1122_p
  );


  and

  (
    g1124_p,
    n2982_lo_p_spl_,
    n2994_lo_n_spl_1
  );


  or

  (
    g1124_n,
    n2982_lo_n_spl_1,
    n2994_lo_p_spl_0
  );


  and

  (
    g1125_p,
    n2982_lo_n_spl_1,
    n2994_lo_p_spl_0
  );


  or

  (
    g1125_n,
    n2982_lo_p_spl_,
    n2994_lo_n_spl_1
  );


  and

  (
    g1126_p,
    g1124_n,
    g1125_n
  );


  or

  (
    g1126_n,
    g1124_p,
    g1125_p
  );


  and

  (
    g1127_p,
    n3282_lo_n_spl_,
    lo510_buf_o2_n_spl_1
  );


  or

  (
    g1127_n,
    n3282_lo_p_spl_,
    lo510_buf_o2_p_spl_
  );


  and

  (
    g1128_p,
    n3282_lo_p_spl_,
    lo510_buf_o2_p_spl_
  );


  or

  (
    g1128_n,
    n3282_lo_n_spl_,
    lo510_buf_o2_n_spl_1
  );


  and

  (
    g1129_p,
    g1127_n,
    g1128_n
  );


  or

  (
    g1129_n,
    g1127_p,
    g1128_p
  );


  and

  (
    g1130_p,
    g1126_p,
    g1129_p
  );


  and

  (
    g1131_p,
    g1126_n,
    g1129_n
  );


  or

  (
    g1132_n,
    g1130_p,
    g1131_p
  );


  and

  (
    g1133_p,
    n4039_o2_n_spl_,
    g1055_n_spl_0
  );


  or

  (
    g1133_n,
    n4039_o2_p_spl_0,
    g1055_p_spl_
  );


  and

  (
    g1134_p,
    n4039_o2_p_spl_,
    g1055_p_spl_
  );


  or

  (
    g1134_n,
    n4039_o2_n_spl_,
    g1055_n_spl_
  );


  and

  (
    g1135_p,
    g1133_n,
    g1134_n
  );


  or

  (
    g1135_n,
    g1133_p,
    g1134_p
  );


  or

  (
    g1136_n,
    g938_p,
    g1135_p
  );


  or

  (
    g1137_n,
    g938_n_spl_0,
    g1135_n
  );


  and

  (
    g1138_p,
    g1136_n,
    g1137_n
  );


  and

  (
    g1139_p,
    lo606_buf_o2_p_spl_,
    lo610_buf_o2_n_spl_
  );


  or

  (
    g1139_n,
    lo606_buf_o2_n_spl_,
    lo610_buf_o2_p_spl_
  );


  and

  (
    g1140_p,
    lo606_buf_o2_n_spl_,
    lo610_buf_o2_p_spl_
  );


  or

  (
    g1140_n,
    lo606_buf_o2_p_spl_,
    lo610_buf_o2_n_spl_
  );


  and

  (
    g1141_p,
    g1139_n,
    g1140_n
  );


  or

  (
    g1141_n,
    g1139_p,
    g1140_p
  );


  and

  (
    g1142_p,
    lo590_buf_o2_p_spl_,
    lo594_buf_o2_n_spl_
  );


  or

  (
    g1142_n,
    lo590_buf_o2_n_spl_,
    lo594_buf_o2_p_spl_
  );


  and

  (
    g1143_p,
    lo590_buf_o2_n_spl_,
    lo594_buf_o2_p_spl_
  );


  or

  (
    g1143_n,
    lo590_buf_o2_p_spl_,
    lo594_buf_o2_n_spl_
  );


  and

  (
    g1144_p,
    g1142_n,
    g1143_n
  );


  or

  (
    g1144_n,
    g1142_p,
    g1143_p
  );


  and

  (
    g1145_p,
    g1141_p_spl_,
    g1144_p_spl_
  );


  or

  (
    g1145_n,
    g1141_n_spl_,
    g1144_n_spl_
  );


  and

  (
    g1146_p,
    g1141_n_spl_,
    g1144_n_spl_
  );


  or

  (
    g1146_n,
    g1141_p_spl_,
    g1144_p_spl_
  );


  and

  (
    g1147_p,
    g1145_n,
    g1146_n
  );


  or

  (
    g1147_n,
    g1145_p,
    g1146_p
  );


  and

  (
    g1148_p,
    n3210_lo_p_spl_,
    n3222_lo_n_spl_
  );


  or

  (
    g1148_n,
    n3210_lo_n_spl_,
    n3222_lo_p_spl_
  );


  and

  (
    g1149_p,
    n3210_lo_n_spl_,
    n3222_lo_p_spl_
  );


  or

  (
    g1149_n,
    n3210_lo_p_spl_,
    n3222_lo_n_spl_
  );


  and

  (
    g1150_p,
    g1148_n,
    g1149_n
  );


  or

  (
    g1150_n,
    g1148_p,
    g1149_p
  );


  or

  (
    g1151_n,
    g1147_p,
    g1150_n
  );


  or

  (
    g1152_n,
    g1147_n,
    g1150_p
  );


  and

  (
    g1153_p,
    g1151_n,
    g1152_n
  );


  and

  (
    g1154_p,
    g908_p,
    g913_p_spl_0
  );


  and

  (
    g1155_p,
    g908_n_spl_1,
    g913_n_spl_
  );


  or

  (
    g1156_n,
    g1154_p,
    g1155_p
  );


  or

  (
    g1157_n,
    g919_n_spl_0,
    g925_p_spl_
  );


  or

  (
    g1158_n,
    g919_p_spl_,
    g925_n_spl_0
  );


  and

  (
    g1159_p,
    g1157_n,
    g1158_n
  );


  and

  (
    g1160_p,
    g1156_n_spl_,
    g1159_p_spl_
  );


  or

  (
    g1161_n,
    g1156_n_spl_,
    g1159_p_spl_
  );


  and

  (
    g1162_p,
    n2386_o2_p_spl_0,
    n2539_o2_p_spl_
  );


  or

  (
    g1162_n,
    n2386_o2_n_spl_0,
    n2539_o2_n_spl_
  );


  and

  (
    g1163_p,
    n2386_o2_n_spl_,
    n2539_o2_n_spl_
  );


  or

  (
    g1163_n,
    n2386_o2_p_spl_,
    n2539_o2_p_spl_
  );


  and

  (
    g1164_p,
    g1162_n,
    g1163_n
  );


  or

  (
    g1164_n,
    g1162_p,
    g1163_p
  );


  and

  (
    g1165_p,
    n1475_inv_n_spl_,
    n2367_o2_p_spl_0
  );


  or

  (
    g1165_n,
    n1475_inv_p_spl_0,
    n2367_o2_n_spl_
  );


  and

  (
    g1166_p,
    n1475_inv_p_spl_1,
    n2367_o2_n_spl_
  );


  or

  (
    g1166_n,
    n1475_inv_n_spl_,
    n2367_o2_p_spl_
  );


  and

  (
    g1167_p,
    g1165_n,
    g1166_n
  );


  or

  (
    g1167_n,
    g1165_p,
    g1166_p
  );


  and

  (
    g1168_p,
    g1164_p_spl_,
    g1167_p_spl_
  );


  or

  (
    g1168_n,
    g1164_n_spl_,
    g1167_n_spl_
  );


  and

  (
    g1169_p,
    g1164_n_spl_,
    g1167_n_spl_
  );


  or

  (
    g1169_n,
    g1164_p_spl_,
    g1167_p_spl_
  );


  and

  (
    g1170_p,
    g1168_n,
    g1169_n
  );


  or

  (
    g1170_n,
    g1168_p,
    g1169_p
  );


  and

  (
    g1171_p,
    g971_n_spl_1,
    g1051_p_spl_
  );


  or

  (
    g1171_n,
    g971_p_spl_0,
    g1051_n_spl_1
  );


  and

  (
    g1172_p,
    g971_p_spl_,
    g1051_n_spl_1
  );


  or

  (
    g1172_n,
    g971_n_spl_1,
    g1051_p_spl_
  );


  and

  (
    g1173_p,
    g1171_n,
    g1172_n
  );


  or

  (
    g1173_n,
    g1171_p,
    g1172_p
  );


  and

  (
    g1174_p,
    g1170_n,
    g1173_p
  );


  and

  (
    g1175_p,
    g1170_p,
    g1173_n
  );


  or

  (
    g1176_n,
    g1174_p,
    g1175_p
  );


  or

  (
    g1177_n,
    n2115_lo_n,
    lo466_buf_o2_p_spl_000
  );


  and

  (
    g1178_p,
    lo478_buf_o2_n_spl_0,
    g1177_n
  );


  and

  (
    g1179_p,
    lo466_buf_o2_n_spl_001,
    lo149_buf_o2_n
  );


  and

  (
    g1180_p,
    lo478_buf_o2_p_spl_001,
    g1179_p
  );


  and

  (
    g1181_p,
    n2247_lo_n,
    lo466_buf_o2_p_spl_001
  );


  or

  (
    g1182_n,
    g1180_p,
    g1181_p
  );


  or

  (
    g1183_n,
    g1178_p,
    g1182_n
  );


  and

  (
    g1184_p,
    n1803_lo_p,
    lo466_buf_o2_n_spl_001
  );


  and

  (
    g1185_p,
    n1815_lo_p,
    lo466_buf_o2_n_spl_010
  );


  and

  (
    g1186_p,
    n2055_lo_p,
    lo466_buf_o2_n_spl_010
  );


  and

  (
    g1187_p,
    n2067_lo_p,
    lo466_buf_o2_n_spl_011
  );


  and

  (
    g1188_p,
    n2091_lo_p,
    lo466_buf_o2_n_spl_011
  );


  and

  (
    g1189_p,
    n2187_lo_p,
    lo466_buf_o2_p_spl_001
  );


  and

  (
    g1190_p,
    n2199_lo_p,
    lo466_buf_o2_p_spl_01
  );


  and

  (
    g1191_p,
    n2223_lo_n,
    lo466_buf_o2_p_spl_01
  );


  and

  (
    g1192_p,
    n1827_lo_n,
    lo478_buf_o2_p_spl_001
  );


  or

  (
    g1193_n,
    n2079_lo_p,
    lo478_buf_o2_p_spl_010
  );


  and

  (
    g1194_p,
    n1839_lo_n,
    lo466_buf_o2_n_spl_100
  );


  and

  (
    g1195_p,
    lo478_buf_o2_p_spl_010,
    g1194_p
  );


  and

  (
    g1196_p,
    n2103_lo_p,
    lo466_buf_o2_n_spl_100
  );


  or

  (
    g1197_n,
    lo478_buf_o2_p_spl_01,
    g1196_p
  );


  and

  (
    g1198_p,
    n2283_lo_p,
    lo466_buf_o2_p_spl_10
  );


  and

  (
    g1199_p,
    n1899_lo_p,
    lo466_buf_o2_n_spl_101
  );


  or

  (
    g1200_n,
    g1198_p,
    g1199_p
  );


  and

  (
    g1201_p,
    lo478_buf_o2_p_spl_10,
    g1200_n
  );


  or

  (
    g1202_n,
    n3063_lo_p_spl_,
    g941_n_spl_0
  );


  or

  (
    g1203_n,
    n2919_lo_p_spl_,
    g941_p_spl_00
  );


  and

  (
    g1204_p,
    g1202_n,
    g1203_n
  );


  and

  (
    g1205_p,
    g995_n_spl_0,
    g1204_p_spl_
  );


  and

  (
    g1206_p,
    n2343_lo_p,
    lo578_buf_o2_n_spl_000
  );


  and

  (
    g1207_p,
    n2703_lo_p,
    lo578_buf_o2_p_spl_000
  );


  or

  (
    g1208_n,
    g1206_p,
    g1207_p
  );


  and

  (
    g1209_p,
    n2391_lo_p,
    lo578_buf_o2_n_spl_000
  );


  and

  (
    g1210_p,
    n2751_lo_p,
    lo578_buf_o2_p_spl_000
  );


  or

  (
    g1211_n,
    g1209_p,
    g1210_p
  );


  and

  (
    g1212_p,
    n2403_lo_p,
    lo578_buf_o2_n_spl_001
  );


  and

  (
    g1213_p,
    n2763_lo_p,
    lo578_buf_o2_p_spl_001
  );


  or

  (
    g1214_n,
    g1212_p,
    g1213_p
  );


  and

  (
    g1215_p,
    n2463_lo_p,
    lo578_buf_o2_n_spl_001
  );


  and

  (
    g1216_p,
    n2583_lo_p,
    lo578_buf_o2_p_spl_001
  );


  or

  (
    g1217_n,
    g1215_p,
    g1216_p
  );


  and

  (
    g1218_p,
    n2511_lo_p,
    lo578_buf_o2_n_spl_010
  );


  and

  (
    g1219_p,
    n2631_lo_p,
    lo578_buf_o2_p_spl_010
  );


  or

  (
    g1220_n,
    g1218_p,
    g1219_p
  );


  and

  (
    g1221_p,
    n2523_lo_p,
    lo578_buf_o2_n_spl_010
  );


  and

  (
    g1222_p,
    n2643_lo_p,
    lo578_buf_o2_p_spl_010
  );


  or

  (
    g1223_n,
    g1221_p,
    g1222_p
  );


  and

  (
    g1224_p,
    n2379_lo_p,
    lo578_buf_o2_n_spl_011
  );


  and

  (
    g1225_p,
    n2739_lo_p,
    lo578_buf_o2_p_spl_011
  );


  or

  (
    g1226_n,
    g1224_p,
    g1225_p
  );


  and

  (
    g1227_p,
    lo582_buf_o2_p_spl_0,
    g1226_n
  );


  and

  (
    g1228_p,
    n2499_lo_p,
    lo578_buf_o2_n_spl_011
  );


  and

  (
    g1229_p,
    n2619_lo_p,
    lo578_buf_o2_p_spl_011
  );


  or

  (
    g1230_n,
    g1228_p,
    g1229_p
  );


  and

  (
    g1231_p,
    lo582_buf_o2_n_spl_0,
    g1230_n
  );


  or

  (
    g1232_n,
    g1227_p,
    g1231_p
  );


  and

  (
    g1233_p,
    n2307_lo_p,
    lo578_buf_o2_n_spl_10
  );


  and

  (
    g1234_p,
    n2667_lo_p,
    lo578_buf_o2_p_spl_100
  );


  or

  (
    g1235_n,
    g1233_p,
    g1234_p
  );


  and

  (
    g1236_p,
    lo582_buf_o2_p_spl_0,
    g1235_n
  );


  and

  (
    g1237_p,
    n2427_lo_p,
    lo578_buf_o2_n_spl_10
  );


  and

  (
    g1238_p,
    n2547_lo_p,
    lo578_buf_o2_p_spl_100
  );


  or

  (
    g1239_n,
    g1237_p,
    g1238_p
  );


  and

  (
    g1240_p,
    lo582_buf_o2_n_spl_0,
    g1239_n
  );


  or

  (
    g1241_n,
    g1236_p,
    g1240_p
  );


  and

  (
    g1242_p,
    n2415_lo_p,
    lo578_buf_o2_n_spl_11
  );


  and

  (
    g1243_p,
    n2775_lo_p,
    lo578_buf_o2_p_spl_10
  );


  or

  (
    g1244_n,
    g1242_p,
    g1243_p
  );


  and

  (
    g1245_p,
    lo582_buf_o2_p_spl_1,
    g1244_n
  );


  and

  (
    g1246_p,
    n2535_lo_p,
    lo578_buf_o2_n_spl_11
  );


  and

  (
    g1247_p,
    n2655_lo_p,
    lo578_buf_o2_p_spl_11
  );


  or

  (
    g1248_n,
    g1246_p,
    g1247_p
  );


  and

  (
    g1249_p,
    lo582_buf_o2_n_spl_,
    g1248_n
  );


  or

  (
    g1250_n,
    g1245_p,
    g1249_p
  );


  and

  (
    g1251_p,
    n1851_lo_n,
    lo466_buf_o2_n_spl_101
  );


  and

  (
    g1252_p,
    lo478_buf_o2_p_spl_10,
    g1251_p
  );


  and

  (
    g1253_p,
    n2235_lo_n,
    lo466_buf_o2_p_spl_10
  );


  or

  (
    g1254_n,
    g1252_p,
    g1253_p
  );


  and

  (
    g1255_p,
    n2259_lo_p,
    lo466_buf_o2_p_spl_11
  );


  and

  (
    g1256_p,
    n1875_lo_p,
    lo466_buf_o2_n_spl_110
  );


  or

  (
    g1257_n,
    g1255_p,
    g1256_p
  );


  and

  (
    g1258_p,
    lo478_buf_o2_p_spl_11,
    g1257_n
  );


  and

  (
    g1259_p,
    n1995_lo_p,
    n1913_inv_p_spl_0
  );


  and

  (
    g1260_p,
    n2127_lo_p,
    lo466_buf_o2_n_spl_110
  );


  and

  (
    g1261_p,
    lo478_buf_o2_n_spl_1,
    g1260_p
  );


  or

  (
    g1262_n,
    g1259_p,
    g1261_p
  );


  or

  (
    g1263_n,
    g1258_p,
    g1262_n
  );


  and

  (
    g1264_p,
    n2019_lo_p,
    n1913_inv_p_spl_1
  );


  and

  (
    g1265_p,
    n2151_lo_p,
    lo466_buf_o2_n_spl_11
  );


  and

  (
    g1266_p,
    lo478_buf_o2_n_spl_1,
    g1265_p
  );


  or

  (
    g1267_n,
    g1264_p,
    g1266_p
  );


  and

  (
    g1268_p,
    g1040_n_spl_,
    g1183_n_spl_
  );


  or

  (
    g1269_n,
    n3075_lo_p_spl_,
    g941_n_spl_0
  );


  or

  (
    g1270_n,
    n2943_lo_p_spl_,
    g941_p_spl_00
  );


  and

  (
    g1271_p,
    g1269_n,
    g1270_n
  );


  or

  (
    g1272_n,
    n3087_lo_p_spl_,
    g941_n_spl_1
  );


  or

  (
    g1273_n,
    n2955_lo_p_spl_,
    g941_p_spl_0
  );


  and

  (
    g1274_p,
    g1272_n,
    g1273_n
  );


  or

  (
    g1275_n,
    g995_n_spl_0,
    g1204_p_spl_
  );


  and

  (
    g1276_p,
    n3039_lo_p_spl_,
    g941_p_spl_1
  );


  and

  (
    g1277_p,
    n2907_lo_p_spl_,
    g941_n_spl_1
  );


  or

  (
    g1278_n,
    g986_n_spl_,
    g1277_p
  );


  or

  (
    g1279_n,
    g1276_p,
    g1278_n
  );


  and

  (
    g1280_p,
    g1275_n,
    g1279_n
  );


  or

  (
    g1281_n,
    lo312_buf_o2_n,
    lo576_buf_o2_p_spl_00
  );


  or

  (
    g1282_n,
    lo432_buf_o2_n,
    lo576_buf_o2_n_spl_0
  );


  and

  (
    g1283_p,
    g1281_n,
    g1282_n
  );


  or

  (
    g1284_n,
    n3156_lo_n_spl_,
    g1283_p
  );


  or

  (
    g1285_n,
    lo352_buf_o2_n,
    lo576_buf_o2_p_spl_00
  );


  or

  (
    g1286_n,
    lo392_buf_o2_n,
    lo576_buf_o2_n_spl_0
  );


  and

  (
    g1287_p,
    g1285_n,
    g1286_n
  );


  or

  (
    g1288_n,
    n3156_lo_p_spl_0,
    g1287_p
  );


  and

  (
    g1289_p,
    n1776_lo_p,
    n2808_lo_n_spl_
  );


  and

  (
    g1290_p,
    n2028_lo_p,
    n2808_lo_n_spl_
  );


  and

  (
    g1291_p,
    n2160_lo_p,
    n2808_lo_p_spl_0
  );


  and

  (
    g1292_p,
    n2808_lo_p_spl_0,
    n2844_lo_n
  );


  and

  (
    g1293_p,
    g1284_n_spl_,
    g1288_n_spl_
  );


  and

  (
    g1294_p,
    lo316_buf_o2_p,
    lo576_buf_o2_n_spl_1
  );


  and

  (
    g1295_p,
    lo436_buf_o2_p,
    lo576_buf_o2_p_spl_0
  );


  or

  (
    g1296_n,
    g1294_p,
    g1295_p
  );


  and

  (
    g1297_p,
    n3156_lo_p_spl_0,
    g1296_n
  );


  and

  (
    g1298_p,
    lo356_buf_o2_p,
    lo576_buf_o2_n_spl_1
  );


  and

  (
    g1299_p,
    lo396_buf_o2_p,
    lo576_buf_o2_p_spl_1
  );


  or

  (
    g1300_n,
    g1298_p,
    g1299_p
  );


  and

  (
    g1301_p,
    n3156_lo_n_spl_,
    g1300_n
  );


  or

  (
    g1302_n,
    g1297_p,
    g1301_p
  );


  buf

  (
    G2531,
    n2793_lo_n_spl_0
  );


  buf

  (
    G2532,
    n2793_lo_n_spl_1
  );


  buf

  (
    G2533,
    n2793_lo_n_spl_1
  );


  buf

  (
    G2534,
    n2901_lo_n_spl_
  );


  buf

  (
    G2535,
    n2901_lo_n_spl_
  );


  buf

  (
    G2536,
    n3057_lo_n_spl_0
  );


  buf

  (
    G2537,
    n3057_lo_n_spl_0
  );


  buf

  (
    G2538,
    n3057_lo_n_spl_
  );


  buf

  (
    G2539,
    n1797_lo_n
  );


  buf

  (
    G2540,
    n2685_lo_n
  );


  buf

  (
    G2541,
    n2181_lo_n
  );


  buf

  (
    G2542,
    n2325_lo_n
  );


  buf

  (
    G2543,
    n2049_lo_n
  );


  buf

  (
    G2544,
    n2565_lo_n
  );


  buf

  (
    G2545,
    n1929_lo_n
  );


  buf

  (
    G2546,
    n2445_lo_n
  );


  buf

  (
    G2547,
    g733_n
  );


  buf

  (
    G2548,
    g735_n
  );


  buf

  (
    G2549,
    n2793_lo_p
  );


  buf

  (
    G2550,
    g736_p
  );


  buf

  (
    G2551,
    g737_n_spl_
  );


  buf

  (
    G2552,
    g738_n
  );


  buf

  (
    G2553,
    g739_n
  );


  buf

  (
    G2554,
    g742_n_spl_
  );


  buf

  (
    G2555,
    g742_n_spl_
  );


  buf

  (
    G2556,
    g745_n_spl_
  );


  buf

  (
    G2557,
    g746_p
  );


  buf

  (
    G2558,
    g747_p
  );


  buf

  (
    G2559,
    n1391_inv_n
  );


  buf

  (
    G2560,
    g748_p
  );


  not

  (
    G2561,
    g749_n_spl_
  );


  buf

  (
    G2562,
    n1445_inv_n
  );


  buf

  (
    G2563,
    g750_n
  );


  buf

  (
    G2564,
    g753_n
  );


  buf

  (
    G2565,
    g755_n
  );


  buf

  (
    G2566,
    n4017_o2_p
  );


  buf

  (
    G2567,
    n4019_o2_p_spl_
  );


  buf

  (
    G2568,
    n2186_o2_p
  );


  buf

  (
    G2569,
    n2176_o2_p
  );


  buf

  (
    G2570,
    n2227_o2_p
  );


  buf

  (
    G2571,
    n2236_o2_p
  );


  buf

  (
    G2572,
    n2245_o2_p
  );


  buf

  (
    G2573,
    g758_p_spl_
  );


  buf

  (
    G2574,
    g758_p_spl_
  );


  not

  (
    G2575,
    g761_n_spl_
  );


  not

  (
    G2576,
    g761_n_spl_
  );


  buf

  (
    G2577,
    g763_n
  );


  buf

  (
    G2578,
    g766_p_spl_
  );


  buf

  (
    G2579,
    g766_p_spl_
  );


  buf

  (
    G2580,
    g770_n
  );


  not

  (
    G2581,
    g774_p_spl_
  );


  buf

  (
    G2582,
    g779_p_spl_
  );


  buf

  (
    G2583,
    g788_p_spl_
  );


  buf

  (
    G2584,
    g838_n_spl_
  );


  buf

  (
    G2585,
    g838_n_spl_
  );


  buf

  (
    G2586,
    g845_n
  );


  not

  (
    G2587,
    g849_p_spl_
  );


  buf

  (
    G2588,
    g859_p_spl_
  );


  buf

  (
    G2589,
    g859_p_spl_
  );


  not

  (
    G2590,
    g864_p_spl_
  );


  buf

  (
    G2591,
    g890_p
  );


  buf

  (
    G2592,
    1'b0
  );


  buf

  (
    G2593,
    g895_n_spl_
  );


  buf

  (
    G2594,
    g895_n_spl_
  );


  buf

  (
    n4649_li000_li000,
    G1_p
  );


  buf

  (
    n4652_li001_li001,
    n1416_lo_p
  );


  buf

  (
    n4655_li002_li002,
    n1419_lo_p
  );


  buf

  (
    n4658_li003_li003,
    n1422_lo_p
  );


  buf

  (
    n4661_li004_li004,
    G2_p
  );


  buf

  (
    n4664_li005_li005,
    n1428_lo_p
  );


  buf

  (
    n4667_li006_li006,
    n1431_lo_p
  );


  buf

  (
    n4670_li007_li007,
    n1434_lo_p
  );


  buf

  (
    n4673_li008_li008,
    G3_p
  );


  buf

  (
    n4676_li009_li009,
    n1440_lo_p
  );


  buf

  (
    n4679_li010_li010,
    n1443_lo_p
  );


  buf

  (
    n4682_li011_li011,
    n1446_lo_p
  );


  buf

  (
    n4685_li012_li012,
    G4_p
  );


  buf

  (
    n4688_li013_li013,
    n1452_lo_p
  );


  buf

  (
    n4691_li014_li014,
    n1455_lo_p
  );


  buf

  (
    n4697_li016_li016,
    G5_p
  );


  buf

  (
    n4700_li017_li017,
    n1464_lo_p
  );


  buf

  (
    n4703_li018_li018,
    n1467_lo_p
  );


  buf

  (
    n4709_li020_li020,
    G6_p
  );


  buf

  (
    n4712_li021_li021,
    n1476_lo_p
  );


  buf

  (
    n4715_li022_li022,
    n1479_lo_p
  );


  buf

  (
    n4721_li024_li024,
    G7_p
  );


  buf

  (
    n4724_li025_li025,
    n1488_lo_p
  );


  buf

  (
    n4727_li026_li026,
    n1491_lo_p
  );


  buf

  (
    n4730_li027_li027,
    n1494_lo_p
  );


  buf

  (
    n4733_li028_li028,
    G8_p
  );


  buf

  (
    n4736_li029_li029,
    n1500_lo_p
  );


  buf

  (
    n4745_li032_li032,
    G9_p
  );


  buf

  (
    n4748_li033_li033,
    n1512_lo_p
  );


  buf

  (
    n4751_li034_li034,
    n1515_lo_p
  );


  buf

  (
    n4754_li035_li035,
    n1518_lo_p
  );


  buf

  (
    n4757_li036_li036,
    G10_p
  );


  buf

  (
    n4760_li037_li037,
    n1524_lo_p
  );


  buf

  (
    n4763_li038_li038,
    n1527_lo_p
  );


  buf

  (
    n4766_li039_li039,
    n1530_lo_p
  );


  buf

  (
    n4769_li040_li040,
    G11_p
  );


  buf

  (
    n4772_li041_li041,
    n1536_lo_p
  );


  buf

  (
    n4775_li042_li042,
    n1539_lo_p
  );


  buf

  (
    n4778_li043_li043,
    n1542_lo_p
  );


  buf

  (
    n4781_li044_li044,
    G12_p
  );


  buf

  (
    n4784_li045_li045,
    n1548_lo_p
  );


  buf

  (
    n4787_li046_li046,
    n1551_lo_p
  );


  buf

  (
    n4793_li048_li048,
    G13_p
  );


  buf

  (
    n4796_li049_li049,
    n1560_lo_p
  );


  buf

  (
    n4799_li050_li050,
    n1563_lo_p
  );


  buf

  (
    n4805_li052_li052,
    G14_p
  );


  buf

  (
    n4808_li053_li053,
    n1572_lo_p
  );


  buf

  (
    n4811_li054_li054,
    n1575_lo_p
  );


  buf

  (
    n4817_li056_li056,
    G15_p
  );


  buf

  (
    n4820_li057_li057,
    n1584_lo_p
  );


  buf

  (
    n4823_li058_li058,
    n1587_lo_p
  );


  buf

  (
    n4829_li060_li060,
    G16_p
  );


  buf

  (
    n4832_li061_li061,
    n1596_lo_p
  );


  buf

  (
    n4835_li062_li062,
    n1599_lo_p
  );


  buf

  (
    n4841_li064_li064,
    G17_p
  );


  buf

  (
    n4844_li065_li065,
    n1608_lo_p
  );


  buf

  (
    n4847_li066_li066,
    n1611_lo_p
  );


  buf

  (
    n4853_li068_li068,
    G18_p
  );


  buf

  (
    n4856_li069_li069,
    n1620_lo_p
  );


  buf

  (
    n4859_li070_li070,
    n1623_lo_p
  );


  buf

  (
    n4865_li072_li072,
    G19_p
  );


  buf

  (
    n4868_li073_li073,
    n1632_lo_p
  );


  buf

  (
    n4871_li074_li074,
    n1635_lo_p
  );


  buf

  (
    n4877_li076_li076,
    G20_p
  );


  buf

  (
    n4880_li077_li077,
    n1644_lo_p
  );


  buf

  (
    n4883_li078_li078,
    n1647_lo_p
  );


  buf

  (
    n4889_li080_li080,
    G21_p
  );


  buf

  (
    n4892_li081_li081,
    n1656_lo_p
  );


  buf

  (
    n4895_li082_li082,
    n1659_lo_p
  );


  buf

  (
    n4901_li084_li084,
    G22_p
  );


  buf

  (
    n4904_li085_li085,
    n1668_lo_p
  );


  buf

  (
    n4907_li086_li086,
    n1671_lo_p
  );


  buf

  (
    n4913_li088_li088,
    G23_p
  );


  buf

  (
    n4916_li089_li089,
    n1680_lo_p
  );


  buf

  (
    n4919_li090_li090,
    n1683_lo_p
  );


  buf

  (
    n4925_li092_li092,
    G24_p
  );


  buf

  (
    n4928_li093_li093,
    n1692_lo_p
  );


  buf

  (
    n4931_li094_li094,
    n1695_lo_p
  );


  buf

  (
    n4937_li096_li096,
    G25_p
  );


  buf

  (
    n4940_li097_li097,
    n1704_lo_p
  );


  buf

  (
    n4943_li098_li098,
    n1707_lo_p
  );


  buf

  (
    n4949_li100_li100,
    G26_p
  );


  buf

  (
    n4952_li101_li101,
    n1716_lo_p
  );


  buf

  (
    n4955_li102_li102,
    n1719_lo_p
  );


  buf

  (
    n4961_li104_li104,
    G27_p
  );


  buf

  (
    n4964_li105_li105,
    n1728_lo_p
  );


  buf

  (
    n4967_li106_li106,
    n1731_lo_p
  );


  buf

  (
    n4973_li108_li108,
    G28_p
  );


  buf

  (
    n4976_li109_li109,
    n1740_lo_p
  );


  buf

  (
    n4979_li110_li110,
    n1743_lo_p
  );


  buf

  (
    n4982_li111_li111,
    n1746_lo_p
  );


  buf

  (
    n4985_li112_li112,
    G29_p
  );


  buf

  (
    n4988_li113_li113,
    n1752_lo_p
  );


  buf

  (
    n4991_li114_li114,
    n1755_lo_p
  );


  buf

  (
    n4994_li115_li115,
    n1758_lo_p
  );


  buf

  (
    n4997_li116_li116,
    G30_p
  );


  buf

  (
    n5009_li120_li120,
    G31_p
  );


  buf

  (
    n5021_li124_li124,
    G32_p
  );


  buf

  (
    n5024_li125_li125,
    n1788_lo_p
  );


  buf

  (
    n5027_li126_li126,
    n1791_lo_p
  );


  buf

  (
    n5030_li127_li127,
    n1794_lo_p_spl_
  );


  buf

  (
    n5033_li128_li128,
    G33_p
  );


  buf

  (
    n5036_li129_li129,
    n1800_lo_p
  );


  buf

  (
    n5045_li132_li132,
    G34_p
  );


  buf

  (
    n5048_li133_li133,
    n1812_lo_p
  );


  buf

  (
    n5057_li136_li136,
    G35_p
  );


  buf

  (
    n5060_li137_li137,
    n1824_lo_p
  );


  buf

  (
    n5069_li140_li140,
    G36_p
  );


  buf

  (
    n5072_li141_li141,
    n1836_lo_p
  );


  buf

  (
    n5081_li144_li144,
    G37_p
  );


  buf

  (
    n5084_li145_li145,
    n1848_lo_p
  );


  buf

  (
    n5093_li148_li148,
    G38_p
  );


  buf

  (
    n5105_li152_li152,
    G39_p
  );


  buf

  (
    n5108_li153_li153,
    n1872_lo_p
  );


  buf

  (
    n5117_li156_li156,
    G40_p
  );


  buf

  (
    n5129_li160_li160,
    G41_p
  );


  buf

  (
    n5132_li161_li161,
    n1896_lo_p
  );


  buf

  (
    n5141_li164_li164,
    G42_p
  );


  buf

  (
    n5153_li168_li168,
    G43_p
  );


  buf

  (
    n5156_li169_li169,
    n1920_lo_p
  );


  buf

  (
    n5159_li170_li170,
    n1923_lo_p
  );


  buf

  (
    n5162_li171_li171,
    n1926_lo_p_spl_
  );


  buf

  (
    n5165_li172_li172,
    G44_p
  );


  buf

  (
    n5168_li173_li173,
    n1932_lo_p
  );


  buf

  (
    n5177_li176_li176,
    G45_p
  );


  buf

  (
    n5180_li177_li177,
    n1944_lo_p
  );


  buf

  (
    n5189_li180_li180,
    G46_p
  );


  buf

  (
    n5192_li181_li181,
    n1956_lo_p
  );


  buf

  (
    n5195_li182_li182,
    n1959_lo_p
  );


  buf

  (
    n5201_li184_li184,
    G47_p
  );


  buf

  (
    n5204_li185_li185,
    n1968_lo_p
  );


  buf

  (
    n5213_li188_li188,
    G48_p
  );


  buf

  (
    n5216_li189_li189,
    n1980_lo_p
  );


  buf

  (
    n5225_li192_li192,
    G49_p
  );


  buf

  (
    n5228_li193_li193,
    n1992_lo_p
  );


  buf

  (
    n5237_li196_li196,
    G50_p
  );


  buf

  (
    n5249_li200_li200,
    G51_p
  );


  buf

  (
    n5252_li201_li201,
    n2016_lo_p
  );


  buf

  (
    n5261_li204_li204,
    G52_p
  );


  buf

  (
    n5273_li208_li208,
    G53_p
  );


  buf

  (
    n5276_li209_li209,
    n2040_lo_p
  );


  buf

  (
    n5279_li210_li210,
    n2043_lo_p
  );


  buf

  (
    n5282_li211_li211,
    n2046_lo_p_spl_
  );


  buf

  (
    n5285_li212_li212,
    G54_p
  );


  buf

  (
    n5288_li213_li213,
    n2052_lo_p
  );


  buf

  (
    n5297_li216_li216,
    G55_p
  );


  buf

  (
    n5300_li217_li217,
    n2064_lo_p
  );


  buf

  (
    n5309_li220_li220,
    G56_p
  );


  buf

  (
    n5312_li221_li221,
    n2076_lo_p
  );


  buf

  (
    n5321_li224_li224,
    G57_p
  );


  buf

  (
    n5324_li225_li225,
    n2088_lo_p
  );


  buf

  (
    n5333_li228_li228,
    G58_p
  );


  buf

  (
    n5336_li229_li229,
    n2100_lo_p
  );


  buf

  (
    n5345_li232_li232,
    G59_p
  );


  buf

  (
    n5348_li233_li233,
    n2112_lo_p
  );


  buf

  (
    n5357_li236_li236,
    G60_p
  );


  buf

  (
    n5360_li237_li237,
    n2124_lo_p
  );


  buf

  (
    n5369_li240_li240,
    G61_p
  );


  buf

  (
    n5381_li244_li244,
    G62_p
  );


  buf

  (
    n5384_li245_li245,
    n2148_lo_p
  );


  buf

  (
    n5393_li248_li248,
    G63_p
  );


  buf

  (
    n5405_li252_li252,
    G64_p
  );


  buf

  (
    n5408_li253_li253,
    n2172_lo_p
  );


  buf

  (
    n5411_li254_li254,
    n2175_lo_p
  );


  buf

  (
    n5414_li255_li255,
    n2178_lo_p_spl_
  );


  buf

  (
    n5417_li256_li256,
    G65_p
  );


  buf

  (
    n5420_li257_li257,
    n2184_lo_p
  );


  buf

  (
    n5429_li260_li260,
    G66_p
  );


  buf

  (
    n5432_li261_li261,
    n2196_lo_p
  );


  buf

  (
    n5441_li264_li264,
    G67_p
  );


  buf

  (
    n5444_li265_li265,
    n2208_lo_p
  );


  buf

  (
    n5453_li268_li268,
    G68_p
  );


  buf

  (
    n5456_li269_li269,
    n2220_lo_p
  );


  buf

  (
    n5465_li272_li272,
    G69_p
  );


  buf

  (
    n5468_li273_li273,
    n2232_lo_p
  );


  buf

  (
    n5477_li276_li276,
    G70_p
  );


  buf

  (
    n5480_li277_li277,
    n2244_lo_p
  );


  buf

  (
    n5489_li280_li280,
    G71_p
  );


  buf

  (
    n5492_li281_li281,
    n2256_lo_p
  );


  buf

  (
    n5501_li284_li284,
    G72_p
  );


  buf

  (
    n5513_li288_li288,
    G73_p
  );


  buf

  (
    n5516_li289_li289,
    n2280_lo_p
  );


  buf

  (
    n5525_li292_li292,
    G74_p
  );


  buf

  (
    n5528_li293_li293,
    n2292_lo_p
  );


  buf

  (
    n5531_li294_li294,
    n2295_lo_p
  );


  buf

  (
    n5534_li295_li295,
    n2298_lo_p
  );


  buf

  (
    n5537_li296_li296,
    G75_p
  );


  buf

  (
    n5540_li297_li297,
    n2304_lo_p
  );


  buf

  (
    n5549_li300_li300,
    G76_p
  );


  buf

  (
    n5552_li301_li301,
    n2316_lo_p
  );


  buf

  (
    n5555_li302_li302,
    n2319_lo_p
  );


  buf

  (
    n5558_li303_li303,
    n2322_lo_p_spl_
  );


  buf

  (
    n5561_li304_li304,
    G77_p
  );


  buf

  (
    n5564_li305_li305,
    n2328_lo_p
  );


  buf

  (
    n5573_li308_li308,
    G78_p
  );


  buf

  (
    n5576_li309_li309,
    n2340_lo_p
  );


  buf

  (
    n5609_li320_li320,
    G81_p
  );


  buf

  (
    n5612_li321_li321,
    n2376_lo_p
  );


  buf

  (
    n5621_li324_li324,
    G82_p
  );


  buf

  (
    n5624_li325_li325,
    n2388_lo_p
  );


  buf

  (
    n5633_li328_li328,
    G83_p
  );


  buf

  (
    n5636_li329_li329,
    n2400_lo_p
  );


  buf

  (
    n5645_li332_li332,
    G84_p
  );


  buf

  (
    n5648_li333_li333,
    n2412_lo_p
  );


  buf

  (
    n5657_li336_li336,
    G85_p
  );


  buf

  (
    n5660_li337_li337,
    n2424_lo_p
  );


  buf

  (
    n5669_li340_li340,
    G86_p
  );


  buf

  (
    n5672_li341_li341,
    n2436_lo_p
  );


  buf

  (
    n5675_li342_li342,
    n2439_lo_p
  );


  buf

  (
    n5678_li343_li343,
    n2442_lo_p_spl_
  );


  buf

  (
    n5681_li344_li344,
    G87_p
  );


  buf

  (
    n5684_li345_li345,
    n2448_lo_p
  );


  buf

  (
    n5693_li348_li348,
    G88_p
  );


  buf

  (
    n5696_li349_li349,
    n2460_lo_p
  );


  buf

  (
    n5729_li360_li360,
    G91_p
  );


  buf

  (
    n5732_li361_li361,
    n2496_lo_p
  );


  buf

  (
    n5741_li364_li364,
    G92_p
  );


  buf

  (
    n5744_li365_li365,
    n2508_lo_p
  );


  buf

  (
    n5753_li368_li368,
    G93_p
  );


  buf

  (
    n5756_li369_li369,
    n2520_lo_p
  );


  buf

  (
    n5765_li372_li372,
    G94_p
  );


  buf

  (
    n5768_li373_li373,
    n2532_lo_p
  );


  buf

  (
    n5777_li376_li376,
    G95_p
  );


  buf

  (
    n5780_li377_li377,
    n2544_lo_p
  );


  buf

  (
    n5789_li380_li380,
    G96_p
  );


  buf

  (
    n5792_li381_li381,
    n2556_lo_p
  );


  buf

  (
    n5795_li382_li382,
    n2559_lo_p
  );


  buf

  (
    n5798_li383_li383,
    n2562_lo_p_spl_
  );


  buf

  (
    n5801_li384_li384,
    G97_p
  );


  buf

  (
    n5804_li385_li385,
    n2568_lo_p
  );


  buf

  (
    n5813_li388_li388,
    G98_p
  );


  buf

  (
    n5816_li389_li389,
    n2580_lo_p
  );


  buf

  (
    n5849_li400_li400,
    G101_p
  );


  buf

  (
    n5852_li401_li401,
    n2616_lo_p
  );


  buf

  (
    n5861_li404_li404,
    G102_p
  );


  buf

  (
    n5864_li405_li405,
    n2628_lo_p
  );


  buf

  (
    n5873_li408_li408,
    G103_p
  );


  buf

  (
    n5876_li409_li409,
    n2640_lo_p
  );


  buf

  (
    n5885_li412_li412,
    G104_p
  );


  buf

  (
    n5888_li413_li413,
    n2652_lo_p
  );


  buf

  (
    n5897_li416_li416,
    G105_p
  );


  buf

  (
    n5900_li417_li417,
    n2664_lo_p
  );


  buf

  (
    n5909_li420_li420,
    G106_p
  );


  buf

  (
    n5912_li421_li421,
    n2676_lo_p
  );


  buf

  (
    n5915_li422_li422,
    n2679_lo_p
  );


  buf

  (
    n5918_li423_li423,
    n2682_lo_p_spl_
  );


  buf

  (
    n5921_li424_li424,
    G107_p
  );


  buf

  (
    n5924_li425_li425,
    n2688_lo_p
  );


  buf

  (
    n5933_li428_li428,
    G108_p
  );


  buf

  (
    n5936_li429_li429,
    n2700_lo_p
  );


  buf

  (
    n5969_li440_li440,
    G111_p
  );


  buf

  (
    n5972_li441_li441,
    n2736_lo_p
  );


  buf

  (
    n5981_li444_li444,
    G112_p
  );


  buf

  (
    n5984_li445_li445,
    n2748_lo_p
  );


  buf

  (
    n5993_li448_li448,
    G113_p
  );


  buf

  (
    n5996_li449_li449,
    n2760_lo_p
  );


  buf

  (
    n6005_li452_li452,
    G114_p
  );


  buf

  (
    n6008_li453_li453,
    n2772_lo_p
  );


  buf

  (
    n6017_li456_li456,
    G115_p
  );


  buf

  (
    n6020_li457_li457,
    n2784_lo_p
  );


  buf

  (
    n6023_li458_li458,
    n2787_lo_p
  );


  buf

  (
    n6026_li459_li459,
    n2790_lo_p
  );


  buf

  (
    n6029_li460_li460,
    G116_p
  );


  buf

  (
    n6032_li461_li461,
    n2796_lo_p
  );


  buf

  (
    n6035_li462_li462,
    n2799_lo_p
  );


  buf

  (
    n6038_li463_li463,
    n2802_lo_p
  );


  buf

  (
    n6041_li464_li464,
    G117_p
  );


  buf

  (
    n6053_li468_li468,
    G118_p
  );


  buf

  (
    n6056_li469_li469,
    n2820_lo_p
  );


  buf

  (
    n6059_li470_li470,
    n2823_lo_p
  );


  buf

  (
    n6062_li471_li471,
    n2826_lo_p_spl_
  );


  buf

  (
    n6065_li472_li472,
    G119_p
  );


  buf

  (
    n6068_li473_li473,
    n2832_lo_p
  );


  buf

  (
    n6071_li474_li474,
    n2835_lo_p
  );


  buf

  (
    n6074_li475_li475,
    n2838_lo_p
  );


  buf

  (
    n6077_li476_li476,
    G120_p
  );


  buf

  (
    n6089_li480_li480,
    G121_p
  );


  buf

  (
    n6092_li481_li481,
    n2856_lo_p
  );


  buf

  (
    n6095_li482_li482,
    n2859_lo_p
  );


  buf

  (
    n6098_li483_li483,
    n2862_lo_p
  );


  buf

  (
    n6101_li484_li484,
    G122_p
  );


  buf

  (
    n6104_li485_li485,
    n2868_lo_p
  );


  buf

  (
    n6107_li486_li486,
    n2871_lo_p
  );


  buf

  (
    n6110_li487_li487,
    n2874_lo_p
  );


  buf

  (
    n6113_li488_li488,
    G123_p
  );


  buf

  (
    n6116_li489_li489,
    n2880_lo_p
  );


  buf

  (
    n6119_li490_li490,
    n2883_lo_p
  );


  buf

  (
    n6122_li491_li491,
    n2886_lo_p
  );


  buf

  (
    n6125_li492_li492,
    G124_p
  );


  buf

  (
    n6128_li493_li493,
    n2892_lo_p
  );


  buf

  (
    n6131_li494_li494,
    n2895_lo_p
  );


  buf

  (
    n6134_li495_li495,
    n2898_lo_p
  );


  buf

  (
    n6137_li496_li496,
    G125_p
  );


  buf

  (
    n6140_li497_li497,
    n2904_lo_p
  );


  buf

  (
    n6149_li500_li500,
    G126_p
  );


  buf

  (
    n6152_li501_li501,
    n2916_lo_p
  );


  buf

  (
    n6158_li503_li503,
    lo502_buf_o2_p_spl_
  );


  buf

  (
    n6161_li504_li504,
    G127_p
  );


  buf

  (
    n6173_li508_li508,
    G128_p
  );


  buf

  (
    n6176_li509_li509,
    n2940_lo_p
  );


  buf

  (
    n6185_li512_li512,
    G129_p
  );


  buf

  (
    n6188_li513_li513,
    n2952_lo_p
  );


  buf

  (
    n6194_li515_li515,
    lo514_buf_o2_p_spl_
  );


  buf

  (
    n6197_li516_li516,
    G130_p
  );


  buf

  (
    n6200_li517_li517,
    n2964_lo_p
  );


  buf

  (
    n6203_li518_li518,
    n2967_lo_p
  );


  buf

  (
    n6209_li520_li520,
    G131_p
  );


  buf

  (
    n6212_li521_li521,
    n2976_lo_p
  );


  buf

  (
    n6215_li522_li522,
    n2979_lo_p
  );


  buf

  (
    n6221_li524_li524,
    G132_p
  );


  buf

  (
    n6224_li525_li525,
    n2988_lo_p
  );


  buf

  (
    n6227_li526_li526,
    n2991_lo_p
  );


  buf

  (
    n6230_li527_li527,
    n2994_lo_p_spl_
  );


  buf

  (
    n6233_li528_li528,
    G133_p
  );


  buf

  (
    n6236_li529_li529,
    n3000_lo_p
  );


  buf

  (
    n6239_li530_li530,
    n3003_lo_p
  );


  buf

  (
    n6245_li532_li532,
    G134_p
  );


  buf

  (
    n6248_li533_li533,
    n3012_lo_p
  );


  buf

  (
    n6251_li534_li534,
    n3015_lo_p
  );


  buf

  (
    n6254_li535_li535,
    n3018_lo_p_spl_
  );


  buf

  (
    n6257_li536_li536,
    G135_p
  );


  buf

  (
    n6260_li537_li537,
    n3024_lo_p
  );


  buf

  (
    n6263_li538_li538,
    n3027_lo_p
  );


  buf

  (
    n6266_li539_li539,
    n3030_lo_p_spl_
  );


  buf

  (
    n6269_li540_li540,
    G136_p
  );


  buf

  (
    n6272_li541_li541,
    n3036_lo_p
  );


  buf

  (
    n6278_li543_li543,
    lo542_buf_o2_p_spl_
  );


  buf

  (
    n6281_li544_li544,
    G137_p
  );


  buf

  (
    n6284_li545_li545,
    n3048_lo_p
  );


  buf

  (
    n6287_li546_li546,
    n3051_lo_p
  );


  buf

  (
    n6290_li547_li547,
    n3054_lo_p
  );


  buf

  (
    n6293_li548_li548,
    G138_p
  );


  buf

  (
    n6296_li549_li549,
    n3060_lo_p
  );


  buf

  (
    n6302_li551_li551,
    lo550_buf_o2_p_spl_
  );


  buf

  (
    n6305_li552_li552,
    G139_p
  );


  buf

  (
    n6308_li553_li553,
    n3072_lo_p
  );


  buf

  (
    n6314_li555_li555,
    lo554_buf_o2_p_spl_
  );


  buf

  (
    n6317_li556_li556,
    G140_p
  );


  buf

  (
    n6320_li557_li557,
    n3084_lo_p
  );


  buf

  (
    n6326_li559_li559,
    lo558_buf_o2_p_spl_
  );


  buf

  (
    n6329_li560_li560,
    G141_p
  );


  buf

  (
    n6332_li561_li561,
    n3096_lo_p
  );


  buf

  (
    n6335_li562_li562,
    n3099_lo_p
  );


  buf

  (
    n6338_li563_li563,
    n3102_lo_p_spl_
  );


  buf

  (
    n6341_li564_li564,
    G142_p
  );


  buf

  (
    n6344_li565_li565,
    n3108_lo_p
  );


  buf

  (
    n6347_li566_li566,
    n3111_lo_p
  );


  buf

  (
    n6350_li567_li567,
    n3114_lo_p_spl_
  );


  buf

  (
    n6353_li568_li568,
    G143_p
  );


  buf

  (
    n6356_li569_li569,
    n3120_lo_p
  );


  buf

  (
    n6359_li570_li570,
    n3123_lo_p
  );


  buf

  (
    n6362_li571_li571,
    n3126_lo_p_spl_
  );


  buf

  (
    n6365_li572_li572,
    G144_p
  );


  buf

  (
    n6368_li573_li573,
    n3132_lo_p
  );


  buf

  (
    n6371_li574_li574,
    n3135_lo_p
  );


  buf

  (
    n6374_li575_li575,
    n3138_lo_p_spl_
  );


  buf

  (
    n6389_li580_li580,
    G146_p
  );


  buf

  (
    n6401_li584_li584,
    G147_p
  );


  buf

  (
    n6404_li585_li585,
    n3168_lo_p
  );


  buf

  (
    n6407_li586_li586,
    n3171_lo_p
  );


  buf

  (
    n6410_li587_li587,
    n3174_lo_p
  );


  buf

  (
    n6413_li588_li588,
    G148_p
  );


  buf

  (
    n6416_li589_li589,
    n3180_lo_p
  );


  buf

  (
    n6425_li592_li592,
    G149_p
  );


  buf

  (
    n6428_li593_li593,
    n3192_lo_p
  );


  buf

  (
    n6437_li596_li596,
    G150_p
  );


  buf

  (
    n6440_li597_li597,
    n3204_lo_p
  );


  buf

  (
    n6443_li598_li598,
    n3207_lo_p
  );


  buf

  (
    n6449_li600_li600,
    G151_p
  );


  buf

  (
    n6452_li601_li601,
    n3216_lo_p
  );


  buf

  (
    n6455_li602_li602,
    n3219_lo_p
  );


  buf

  (
    n6461_li604_li604,
    G152_p
  );


  buf

  (
    n6464_li605_li605,
    n3228_lo_p
  );


  buf

  (
    n6473_li608_li608,
    G153_p
  );


  buf

  (
    n6476_li609_li609,
    n3240_lo_p
  );


  buf

  (
    n6485_li612_li612,
    G154_p
  );


  buf

  (
    n6488_li613_li613,
    n3252_lo_p
  );


  buf

  (
    n6491_li614_li614,
    n3255_lo_p
  );


  buf

  (
    n6497_li616_li616,
    G155_p
  );


  buf

  (
    n6500_li617_li617,
    n3264_lo_p
  );


  buf

  (
    n6503_li618_li618,
    n3267_lo_p
  );


  buf

  (
    n6509_li620_li620,
    G156_p
  );


  buf

  (
    n6512_li621_li621,
    n3276_lo_p
  );


  buf

  (
    n6515_li622_li622,
    n3279_lo_p
  );


  buf

  (
    n6521_li624_li624,
    G157_p
  );


  buf

  (
    n6524_li625_li625,
    n3288_lo_p
  );


  buf

  (
    n6527_li626_li626,
    n3291_lo_p
  );


  buf

  (
    n3603_i2,
    n4023_o2_p
  );


  buf

  (
    n3604_i2,
    n1466_inv_p
  );


  buf

  (
    n3618_i2,
    n1475_inv_p_spl_1
  );


  buf

  (
    n3798_i2,
    n2205_o2_p_spl_1
  );


  buf

  (
    n3846_i2,
    n2254_o2_p_spl_1
  );


  buf

  (
    n4019_i2,
    n2196_o2_p_spl_1
  );


  buf

  (
    n4017_i2,
    n2220_o2_p_spl_1
  );


  buf

  (
    n2177_i2,
    g896_p_spl_
  );


  buf

  (
    n2150_i2,
    g897_p_spl_
  );


  buf

  (
    n2154_i2,
    g898_p_spl_
  );


  buf

  (
    n2184_i2,
    g899_p_spl_
  );


  buf

  (
    n2515_i2,
    g900_n_spl_
  );


  buf

  (
    n3837_i2,
    lo578_buf_o2_p_spl_11
  );


  buf

  (
    n2167_i2,
    g901_p_spl_
  );


  buf

  (
    n2118_i2,
    g902_p_spl_
  );


  buf

  (
    n2186_i2,
    g903_n_spl_1
  );


  buf

  (
    n2174_i2,
    g906_p_spl_
  );


  buf

  (
    n3964_i2,
    lo582_buf_o2_p_spl_1
  );


  buf

  (
    n4005_i2,
    lo466_buf_o2_p_spl_11
  );


  buf

  (
    n4006_i2,
    lo478_buf_o2_p_spl_11
  );


  buf

  (
    n2195_i2,
    g907_n_spl_
  );


  buf

  (
    n2176_i2,
    g908_n_spl_1
  );


  buf

  (
    n2227_i2,
    g913_p_spl_
  );


  buf

  (
    n2236_i2,
    g919_n_spl_
  );


  buf

  (
    n2245_i2,
    g925_n_spl_
  );


  buf

  (
    n2518_i2,
    g928_n_spl_
  );


  buf

  (
    n4023_i2,
    n2140_o2_p
  );


  buf

  (
    n4024_i2,
    n1877_inv_p
  );


  buf

  (
    n4038_i2,
    n1913_inv_p_spl_1
  );


  buf

  (
    n4039_i2,
    n2146_o2_p_spl_
  );


  buf

  (
    n4040_i2,
    n1919_inv_p_spl_
  );


  not

  (
    n2119_i2,
    g929_n_spl_
  );


  buf

  (
    n2275_i2,
    g938_n_spl_
  );


  buf

  (
    n2595_i2,
    g939_p_spl_
  );


  buf

  (
    n2594_i2,
    g940_p_spl_
  );


  buf

  (
    lo498_buf_i2,
    n2907_lo_p_spl_
  );


  buf

  (
    lo502_buf_i2,
    n2919_lo_p_spl_
  );


  buf

  (
    lo550_buf_i2,
    n3063_lo_p_spl_
  );


  buf

  (
    n2596_i2,
    g941_p_spl_1
  );


  not

  (
    n2593_i2,
    g942_n_spl_
  );


  not

  (
    n2668_i2,
    g944_n_spl_
  );


  buf

  (
    lo542_buf_i2,
    n3039_lo_p_spl_
  );


  buf

  (
    n2667_i2,
    g945_p_spl_
  );


  buf

  (
    n2404_i2,
    g948_n_spl_
  );


  buf

  (
    n2410_i2,
    g951_n_spl_
  );


  buf

  (
    n2419_i2,
    g954_n_spl_
  );


  buf

  (
    n2392_i2,
    g957_n_spl_
  );


  buf

  (
    n2369_i2,
    g960_n_spl_
  );


  buf

  (
    n2397_i2,
    g963_n_spl_
  );


  buf

  (
    n2601_i2,
    g968_n_spl_
  );


  not

  (
    n2658_i2,
    g974_n_spl_
  );


  not

  (
    n2574_i2,
    g980_n_spl_
  );


  buf

  (
    n2205_i2,
    g986_n_spl_
  );


  buf

  (
    lo510_buf_i2,
    n2943_lo_p_spl_
  );


  buf

  (
    lo514_buf_i2,
    n2955_lo_p_spl_
  );


  buf

  (
    lo554_buf_i2,
    n3075_lo_p_spl_
  );


  buf

  (
    lo558_buf_i2,
    n3087_lo_p_spl_
  );


  buf

  (
    lo578_buf_i2,
    lo576_buf_o2_p_spl_1
  );


  buf

  (
    n2254_i2,
    g995_n_spl_
  );


  buf

  (
    n2421_i2,
    g996_p
  );


  buf

  (
    n2422_i2,
    g997_p
  );


  buf

  (
    n2130_i2,
    g998_p
  );


  buf

  (
    n2127_i2,
    g999_p
  );


  buf

  (
    n2131_i2,
    g1000_p
  );


  buf

  (
    n2128_i2,
    g1001_p
  );


  buf

  (
    n2264_i2,
    g1002_n
  );


  not

  (
    n2467_i2,
    g1006_n
  );


  buf

  (
    n2471_i2,
    g1007_p
  );


  not

  (
    n2488_i2,
    g1008_n
  );


  not

  (
    n2478_i2,
    g1012_n
  );


  buf

  (
    n2486_i2,
    g1013_p
  );


  buf

  (
    n2485_i2,
    g1017_p
  );


  not

  (
    n2498_i2,
    g1018_n
  );


  buf

  (
    n2495_i2,
    g1022_p
  );


  not

  (
    n2496_i2,
    g1023_n
  );


  buf

  (
    n2458_i2,
    g1024_p
  );


  buf

  (
    n2643_i2,
    g1025_p
  );


  buf

  (
    n2462_i2,
    g1029_p
  );


  not

  (
    n2468_i2,
    g1030_n
  );


  buf

  (
    n2639_i2,
    g1031_p
  );


  not

  (
    n2499_i2,
    g1032_n
  );


  buf

  (
    n2472_i2,
    g1033_p
  );


  not

  (
    n2474_i2,
    g1034_n
  );


  buf

  (
    n2489_i2,
    g1035_p
  );


  buf

  (
    n2321_i2,
    g1036_p
  );


  buf

  (
    n2322_i2,
    g1037_p
  );


  buf

  (
    n2640_i2,
    g1038_p
  );


  buf

  (
    n2642_i2,
    g1039_p
  );


  not

  (
    n2187_i2,
    g1040_n_spl_
  );


  buf

  (
    n2373_i2,
    g1043_n
  );


  not

  (
    n2603_i2,
    g1044_n
  );


  buf

  (
    n2388_i2,
    g1047_n
  );


  buf

  (
    n2437_i2,
    g1053_n
  );


  buf

  (
    n2356_i2,
    g1057_n
  );


  buf

  (
    n2452_i2,
    g1060_n
  );


  buf

  (
    n2347_i2,
    g1063_n
  );


  buf

  (
    n2329_i2,
    g1066_n
  );


  not

  (
    n2669_i2,
    g1067_n
  );


  buf

  (
    n2332_i2,
    g1070_n
  );


  buf

  (
    n2664_i2,
    g1073_p
  );


  not

  (
    n2665_i2,
    g1074_n
  );


  buf

  (
    n2653_i2,
    g1077_p
  );


  not

  (
    n2654_i2,
    g1078_n
  );


  not

  (
    n2636_i2,
    g1095_n
  );


  not

  (
    n2660_i2,
    g1097_p
  );


  not

  (
    n2318_i2,
    g1108_n
  );


  buf

  (
    n2319_i2,
    g1109_p
  );


  not

  (
    n2586_i2,
    g1113_p
  );


  not

  (
    n2587_i2,
    g1114_n
  );


  buf

  (
    n2288_i2,
    g1123_n
  );


  buf

  (
    n2344_i2,
    g1132_n
  );


  buf

  (
    n2530_i2,
    g1138_p
  );


  buf

  (
    n2303_i2,
    g1153_p
  );


  buf

  (
    n2566_i2,
    g1160_p
  );


  not

  (
    n2567_i2,
    g1161_n
  );


  buf

  (
    n2554_i2,
    g1176_n
  );


  not

  (
    n2194_i2,
    g1183_n_spl_
  );


  buf

  (
    lo582_buf_i2,
    n3156_lo_p_spl_
  );


  buf

  (
    lo030_buf_i2,
    n1503_lo_p
  );


  buf

  (
    lo174_buf_i2,
    n1935_lo_p
  );


  buf

  (
    lo178_buf_i2,
    n1947_lo_p
  );


  buf

  (
    lo186_buf_i2,
    n1971_lo_p
  );


  buf

  (
    lo266_buf_i2,
    n2211_lo_p
  );


  buf

  (
    lo306_buf_i2,
    n2331_lo_p
  );


  buf

  (
    lo346_buf_i2,
    n2451_lo_p
  );


  buf

  (
    lo386_buf_i2,
    n2571_lo_p
  );


  buf

  (
    lo426_buf_i2,
    n2691_lo_p
  );


  buf

  (
    lo590_buf_i2,
    n3183_lo_p
  );


  buf

  (
    lo594_buf_i2,
    n3195_lo_p
  );


  buf

  (
    lo606_buf_i2,
    n3231_lo_p
  );


  buf

  (
    lo610_buf_i2,
    n3243_lo_p
  );


  buf

  (
    n2238_i2,
    g1184_p
  );


  buf

  (
    n2229_i2,
    g1185_p
  );


  buf

  (
    n2242_i2,
    g1186_p
  );


  buf

  (
    n2233_i2,
    g1187_p
  );


  buf

  (
    n2168_i2,
    g1188_p
  );


  buf

  (
    n2237_i2,
    g1189_p
  );


  buf

  (
    n2228_i2,
    g1190_p
  );


  buf

  (
    n2172_i2,
    g1191_p
  );


  buf

  (
    n2223_i2,
    g1192_p
  );


  buf

  (
    n2222_i2,
    g1193_n
  );


  buf

  (
    n2170_i2,
    g1195_p
  );


  buf

  (
    n2181_i2,
    g1197_n
  );


  buf

  (
    n2510_i2,
    g1201_p
  );


  buf

  (
    n2621_i2,
    g1205_p
  );


  buf

  (
    lo466_buf_i2,
    n2808_lo_p_spl_
  );


  buf

  (
    lo478_buf_i2,
    n2844_lo_p
  );


  buf

  (
    n2149_i2,
    g1208_n
  );


  buf

  (
    n2429_i2,
    g1211_n
  );


  buf

  (
    n2444_i2,
    g1214_n
  );


  buf

  (
    n2153_i2,
    g1217_n
  );


  buf

  (
    n2433_i2,
    g1220_n
  );


  buf

  (
    n2448_i2,
    g1223_n
  );


  buf

  (
    n2367_i2,
    g1232_n
  );


  buf

  (
    n2386_i2,
    g1241_n
  );


  buf

  (
    n2539_i2,
    g1250_n
  );


  buf

  (
    n2183_i2,
    g1254_n
  );


  buf

  (
    n2220_i2,
    g1263_n
  );


  buf

  (
    n2514_i2,
    g1267_n
  );


  not

  (
    n2196_i2,
    g1268_p
  );


  buf

  (
    n2616_i2,
    g1271_p
  );


  buf

  (
    n2612_i2,
    g1274_p
  );


  buf

  (
    n2627_i2,
    g1280_p
  );


  not

  (
    n2140_i2,
    g1284_n_spl_
  );


  not

  (
    n2144_i2,
    g1288_n_spl_
  );


  buf

  (
    lo149_buf_i2,
    n1860_lo_p
  );


  buf

  (
    lo197_buf_i2,
    n2004_lo_p
  );


  buf

  (
    lo118_buf_i2,
    n1764_lo_p
  );


  buf

  (
    lo158_buf_i2,
    n1884_lo_p
  );


  buf

  (
    lo166_buf_i2,
    n1908_lo_p
  );


  buf

  (
    lo242_buf_i2,
    n2136_lo_p
  );


  buf

  (
    lo286_buf_i2,
    n2268_lo_p
  );


  buf

  (
    lo506_buf_i2,
    n2928_lo_p
  );


  buf

  (
    n2198_i2,
    g1289_p
  );


  buf

  (
    n2202_i2,
    g1290_p
  );


  buf

  (
    n2197_i2,
    g1291_p
  );


  buf

  (
    n2166_i2,
    g1292_p
  );


  not

  (
    n2146_i2,
    g1293_p
  );


  buf

  (
    n2165_i2,
    g1302_n
  );


  buf

  (
    lo312_buf_i2,
    G79_p
  );


  buf

  (
    lo316_buf_i2,
    G80_p
  );


  buf

  (
    lo352_buf_i2,
    G89_p
  );


  buf

  (
    lo356_buf_i2,
    G90_p
  );


  buf

  (
    lo392_buf_i2,
    G99_p
  );


  buf

  (
    lo396_buf_i2,
    G100_p
  );


  buf

  (
    lo432_buf_i2,
    G109_p
  );


  buf

  (
    lo436_buf_i2,
    G110_p
  );


  buf

  (
    lo576_buf_i2,
    G145_p
  );


  buf

  (
    n2865_lo_n_spl_,
    n2865_lo_n
  );


  buf

  (
    n2793_lo_n_spl_,
    n2793_lo_n
  );


  buf

  (
    n2793_lo_n_spl_0,
    n2793_lo_n_spl_
  );


  buf

  (
    n2793_lo_n_spl_1,
    n2793_lo_n_spl_
  );


  buf

  (
    g737_n_spl_,
    g737_n
  );


  buf

  (
    g737_n_spl_0,
    g737_n_spl_
  );


  buf

  (
    g740_n_spl_,
    g740_n
  );


  buf

  (
    g741_n_spl_,
    g741_n
  );


  buf

  (
    n2877_lo_n_spl_,
    n2877_lo_n
  );


  buf

  (
    n2877_lo_n_spl_0,
    n2877_lo_n_spl_
  );


  buf

  (
    g745_n_spl_,
    g745_n
  );


  buf

  (
    g745_n_spl_0,
    g745_n_spl_
  );


  buf

  (
    g752_n_spl_,
    g752_n
  );


  buf

  (
    n2889_lo_p_spl_,
    n2889_lo_p
  );


  buf

  (
    n2889_lo_p_spl_0,
    n2889_lo_p_spl_
  );


  buf

  (
    n2889_lo_p_spl_1,
    n2889_lo_p_spl_
  );


  buf

  (
    n3846_o2_n_spl_,
    n3846_o2_n
  );


  buf

  (
    n2889_lo_n_spl_,
    n2889_lo_n
  );


  buf

  (
    n2889_lo_n_spl_0,
    n2889_lo_n_spl_
  );


  buf

  (
    n2889_lo_n_spl_1,
    n2889_lo_n_spl_
  );


  buf

  (
    n4019_o2_p_spl_,
    n4019_o2_p
  );


  buf

  (
    g749_n_spl_,
    g749_n
  );


  buf

  (
    n2829_lo_p_spl_,
    n2829_lo_p
  );


  buf

  (
    n3846_o2_p_spl_,
    n3846_o2_p
  );


  buf

  (
    n2264_o2_n_spl_,
    n2264_o2_n
  );


  buf

  (
    n2264_o2_n_spl_0,
    n2264_o2_n_spl_
  );


  buf

  (
    n2329_o2_p_spl_,
    n2329_o2_p
  );


  buf

  (
    n2332_o2_n_spl_,
    n2332_o2_n
  );


  buf

  (
    n2329_o2_n_spl_,
    n2329_o2_n
  );


  buf

  (
    n2332_o2_p_spl_,
    n2332_o2_p
  );


  buf

  (
    n2347_o2_n_spl_,
    n2347_o2_n
  );


  buf

  (
    n2344_o2_p_spl_,
    n2344_o2_p
  );


  buf

  (
    n2347_o2_p_spl_,
    n2347_o2_p
  );


  buf

  (
    n2344_o2_n_spl_,
    n2344_o2_n
  );


  buf

  (
    n2515_o2_p_spl_,
    n2515_o2_p
  );


  buf

  (
    n1761_lo_n_spl_,
    n1761_lo_n
  );


  buf

  (
    n2574_o2_n_spl_,
    n2574_o2_n
  );


  buf

  (
    n2264_o2_p_spl_,
    n2264_o2_p
  );


  buf

  (
    n2574_o2_p_spl_,
    n2574_o2_p
  );


  buf

  (
    g851_p_spl_,
    g851_p
  );


  buf

  (
    g851_n_spl_,
    g851_n
  );


  buf

  (
    g868_n_spl_,
    g868_n
  );


  buf

  (
    n2660_o2_p_spl_,
    n2660_o2_p
  );


  buf

  (
    g875_n_spl_,
    g875_n
  );


  buf

  (
    g877_n_spl_,
    g877_n
  );


  buf

  (
    g876_n_spl_,
    g876_n
  );


  buf

  (
    g774_p_spl_,
    g774_p
  );


  buf

  (
    g779_p_spl_,
    g779_p
  );


  buf

  (
    g788_p_spl_,
    g788_p
  );


  buf

  (
    g849_p_spl_,
    g849_p
  );


  buf

  (
    g864_p_spl_,
    g864_p
  );


  buf

  (
    n4038_o2_p_spl_,
    n4038_o2_p
  );


  buf

  (
    n4038_o2_p_spl_0,
    n4038_o2_p_spl_
  );


  buf

  (
    n4038_o2_p_spl_1,
    n4038_o2_p_spl_
  );


  buf

  (
    n4038_o2_n_spl_,
    n4038_o2_n
  );


  buf

  (
    n4038_o2_n_spl_0,
    n4038_o2_n_spl_
  );


  buf

  (
    n4038_o2_n_spl_1,
    n4038_o2_n_spl_
  );


  buf

  (
    n3964_o2_p_spl_,
    n3964_o2_p
  );


  buf

  (
    n3964_o2_p_spl_0,
    n3964_o2_p_spl_
  );


  buf

  (
    n3964_o2_p_spl_00,
    n3964_o2_p_spl_0
  );


  buf

  (
    n3964_o2_p_spl_01,
    n3964_o2_p_spl_0
  );


  buf

  (
    n3964_o2_p_spl_1,
    n3964_o2_p_spl_
  );


  buf

  (
    n3964_o2_p_spl_10,
    n3964_o2_p_spl_1
  );


  buf

  (
    n3964_o2_p_spl_11,
    n3964_o2_p_spl_1
  );


  buf

  (
    n3964_o2_n_spl_,
    n3964_o2_n
  );


  buf

  (
    n3964_o2_n_spl_0,
    n3964_o2_n_spl_
  );


  buf

  (
    n3964_o2_n_spl_00,
    n3964_o2_n_spl_0
  );


  buf

  (
    n3964_o2_n_spl_01,
    n3964_o2_n_spl_0
  );


  buf

  (
    n3964_o2_n_spl_1,
    n3964_o2_n_spl_
  );


  buf

  (
    n3964_o2_n_spl_10,
    n3964_o2_n_spl_1
  );


  buf

  (
    n3964_o2_n_spl_11,
    n3964_o2_n_spl_1
  );


  buf

  (
    lo554_buf_o2_p_spl_,
    lo554_buf_o2_p
  );


  buf

  (
    lo554_buf_o2_p_spl_0,
    lo554_buf_o2_p_spl_
  );


  buf

  (
    lo558_buf_o2_p_spl_,
    lo558_buf_o2_p
  );


  buf

  (
    lo558_buf_o2_p_spl_0,
    lo558_buf_o2_p_spl_
  );


  buf

  (
    lo554_buf_o2_n_spl_,
    lo554_buf_o2_n
  );


  buf

  (
    lo554_buf_o2_n_spl_0,
    lo554_buf_o2_n_spl_
  );


  buf

  (
    lo558_buf_o2_n_spl_,
    lo558_buf_o2_n
  );


  buf

  (
    lo558_buf_o2_n_spl_0,
    lo558_buf_o2_n_spl_
  );


  buf

  (
    g896_p_spl_,
    g896_p
  );


  buf

  (
    g899_p_spl_,
    g899_p
  );


  buf

  (
    n4006_o2_n_spl_,
    n4006_o2_n
  );


  buf

  (
    n4006_o2_n_spl_0,
    n4006_o2_n_spl_
  );


  buf

  (
    n4006_o2_n_spl_00,
    n4006_o2_n_spl_0
  );


  buf

  (
    n4006_o2_n_spl_01,
    n4006_o2_n_spl_0
  );


  buf

  (
    n4006_o2_n_spl_1,
    n4006_o2_n_spl_
  );


  buf

  (
    n4006_o2_p_spl_,
    n4006_o2_p
  );


  buf

  (
    n4006_o2_p_spl_0,
    n4006_o2_p_spl_
  );


  buf

  (
    n4006_o2_p_spl_00,
    n4006_o2_p_spl_0
  );


  buf

  (
    n4006_o2_p_spl_01,
    n4006_o2_p_spl_0
  );


  buf

  (
    n4006_o2_p_spl_1,
    n4006_o2_p_spl_
  );


  buf

  (
    g901_p_spl_,
    g901_p
  );


  buf

  (
    g906_p_spl_,
    g906_p
  );


  buf

  (
    n4005_o2_n_spl_,
    n4005_o2_n
  );


  buf

  (
    n4005_o2_p_spl_,
    n4005_o2_p
  );


  buf

  (
    n2205_o2_n_spl_,
    n2205_o2_n
  );


  buf

  (
    g900_n_spl_,
    g900_n
  );


  buf

  (
    g900_n_spl_0,
    g900_n_spl_
  );


  buf

  (
    n2205_o2_p_spl_,
    n2205_o2_p
  );


  buf

  (
    n2205_o2_p_spl_0,
    n2205_o2_p_spl_
  );


  buf

  (
    n2205_o2_p_spl_1,
    n2205_o2_p_spl_
  );


  buf

  (
    g900_p_spl_,
    g900_p
  );


  buf

  (
    n3102_lo_n_spl_,
    n3102_lo_n
  );


  buf

  (
    n3102_lo_n_spl_0,
    n3102_lo_n_spl_
  );


  buf

  (
    n3114_lo_n_spl_,
    n3114_lo_n
  );


  buf

  (
    n3837_o2_n_spl_,
    n3837_o2_n
  );


  buf

  (
    n3837_o2_n_spl_0,
    n3837_o2_n_spl_
  );


  buf

  (
    n3837_o2_n_spl_1,
    n3837_o2_n_spl_
  );


  buf

  (
    n3837_o2_p_spl_,
    n3837_o2_p
  );


  buf

  (
    n3837_o2_p_spl_0,
    n3837_o2_p_spl_
  );


  buf

  (
    n3837_o2_p_spl_1,
    n3837_o2_p_spl_
  );


  buf

  (
    n2146_o2_p_spl_,
    n2146_o2_p
  );


  buf

  (
    n1919_inv_p_spl_,
    n1919_inv_p
  );


  buf

  (
    g939_p_spl_,
    g939_p
  );


  buf

  (
    g940_p_spl_,
    g940_p
  );


  buf

  (
    lo030_buf_o2_n_spl_,
    lo030_buf_o2_n
  );


  buf

  (
    g908_n_spl_,
    g908_n
  );


  buf

  (
    g908_n_spl_0,
    g908_n_spl_
  );


  buf

  (
    g908_n_spl_1,
    g908_n_spl_
  );


  buf

  (
    n3018_lo_p_spl_,
    n3018_lo_p
  );


  buf

  (
    n3018_lo_p_spl_0,
    n3018_lo_p_spl_
  );


  buf

  (
    g943_n_spl_,
    g943_n
  );


  buf

  (
    g943_n_spl_0,
    g943_n_spl_
  );


  buf

  (
    g943_n_spl_00,
    g943_n_spl_0
  );


  buf

  (
    g943_n_spl_1,
    g943_n_spl_
  );


  buf

  (
    g925_p_spl_,
    g925_p
  );


  buf

  (
    g943_p_spl_,
    g943_p
  );


  buf

  (
    g943_p_spl_0,
    g943_p_spl_
  );


  buf

  (
    g943_p_spl_00,
    g943_p_spl_0
  );


  buf

  (
    g943_p_spl_1,
    g943_p_spl_
  );


  buf

  (
    n1554_lo_p_spl_,
    n1554_lo_p
  );


  buf

  (
    n1554_lo_p_spl_0,
    n1554_lo_p_spl_
  );


  buf

  (
    n1554_lo_p_spl_00,
    n1554_lo_p_spl_0
  );


  buf

  (
    n1554_lo_p_spl_000,
    n1554_lo_p_spl_00
  );


  buf

  (
    n1554_lo_p_spl_01,
    n1554_lo_p_spl_0
  );


  buf

  (
    n1554_lo_p_spl_1,
    n1554_lo_p_spl_
  );


  buf

  (
    n1554_lo_p_spl_10,
    n1554_lo_p_spl_1
  );


  buf

  (
    n1554_lo_p_spl_11,
    n1554_lo_p_spl_1
  );


  buf

  (
    n1554_lo_n_spl_,
    n1554_lo_n
  );


  buf

  (
    n1554_lo_n_spl_0,
    n1554_lo_n_spl_
  );


  buf

  (
    n1554_lo_n_spl_00,
    n1554_lo_n_spl_0
  );


  buf

  (
    n1554_lo_n_spl_000,
    n1554_lo_n_spl_00
  );


  buf

  (
    n1554_lo_n_spl_01,
    n1554_lo_n_spl_0
  );


  buf

  (
    n1554_lo_n_spl_1,
    n1554_lo_n_spl_
  );


  buf

  (
    n1554_lo_n_spl_10,
    n1554_lo_n_spl_1
  );


  buf

  (
    n1554_lo_n_spl_11,
    n1554_lo_n_spl_1
  );


  buf

  (
    n2254_o2_p_spl_,
    n2254_o2_p
  );


  buf

  (
    n2254_o2_p_spl_0,
    n2254_o2_p_spl_
  );


  buf

  (
    n2254_o2_p_spl_00,
    n2254_o2_p_spl_0
  );


  buf

  (
    n2254_o2_p_spl_1,
    n2254_o2_p_spl_
  );


  buf

  (
    g925_n_spl_,
    g925_n
  );


  buf

  (
    g925_n_spl_0,
    g925_n_spl_
  );


  buf

  (
    g913_p_spl_,
    g913_p
  );


  buf

  (
    g913_p_spl_0,
    g913_p_spl_
  );


  buf

  (
    n1686_lo_p_spl_,
    n1686_lo_p
  );


  buf

  (
    n1686_lo_p_spl_0,
    n1686_lo_p_spl_
  );


  buf

  (
    n1686_lo_p_spl_00,
    n1686_lo_p_spl_0
  );


  buf

  (
    n1686_lo_p_spl_01,
    n1686_lo_p_spl_0
  );


  buf

  (
    n1686_lo_p_spl_1,
    n1686_lo_p_spl_
  );


  buf

  (
    n1686_lo_p_spl_10,
    n1686_lo_p_spl_1
  );


  buf

  (
    n1686_lo_p_spl_11,
    n1686_lo_p_spl_1
  );


  buf

  (
    n1686_lo_n_spl_,
    n1686_lo_n
  );


  buf

  (
    n1686_lo_n_spl_0,
    n1686_lo_n_spl_
  );


  buf

  (
    n1686_lo_n_spl_00,
    n1686_lo_n_spl_0
  );


  buf

  (
    n1686_lo_n_spl_01,
    n1686_lo_n_spl_0
  );


  buf

  (
    n1686_lo_n_spl_1,
    n1686_lo_n_spl_
  );


  buf

  (
    n1686_lo_n_spl_10,
    n1686_lo_n_spl_1
  );


  buf

  (
    n1686_lo_n_spl_11,
    n1686_lo_n_spl_1
  );


  buf

  (
    n1475_inv_p_spl_,
    n1475_inv_p
  );


  buf

  (
    n1475_inv_p_spl_0,
    n1475_inv_p_spl_
  );


  buf

  (
    n1475_inv_p_spl_1,
    n1475_inv_p_spl_
  );


  buf

  (
    n2367_o2_p_spl_,
    n2367_o2_p
  );


  buf

  (
    n2367_o2_p_spl_0,
    n2367_o2_p_spl_
  );


  buf

  (
    n4039_o2_p_spl_,
    n4039_o2_p
  );


  buf

  (
    n4039_o2_p_spl_0,
    n4039_o2_p_spl_
  );


  buf

  (
    lo030_buf_o2_p_spl_,
    lo030_buf_o2_p
  );


  buf

  (
    n2982_lo_n_spl_,
    n2982_lo_n
  );


  buf

  (
    n2982_lo_n_spl_0,
    n2982_lo_n_spl_
  );


  buf

  (
    n2982_lo_n_spl_00,
    n2982_lo_n_spl_0
  );


  buf

  (
    n2982_lo_n_spl_1,
    n2982_lo_n_spl_
  );


  buf

  (
    g964_p_spl_,
    g964_p
  );


  buf

  (
    g964_p_spl_0,
    g964_p_spl_
  );


  buf

  (
    g964_p_spl_1,
    g964_p_spl_
  );


  buf

  (
    g966_p_spl_,
    g966_p
  );


  buf

  (
    g966_p_spl_0,
    g966_p_spl_
  );


  buf

  (
    g966_p_spl_1,
    g966_p_spl_
  );


  buf

  (
    g971_n_spl_,
    g971_n
  );


  buf

  (
    g971_n_spl_0,
    g971_n_spl_
  );


  buf

  (
    g971_n_spl_1,
    g971_n_spl_
  );


  buf

  (
    g971_p_spl_,
    g971_p
  );


  buf

  (
    g971_p_spl_0,
    g971_p_spl_
  );


  buf

  (
    lo542_buf_o2_n_spl_,
    lo542_buf_o2_n
  );


  buf

  (
    lo542_buf_o2_p_spl_,
    lo542_buf_o2_p
  );


  buf

  (
    lo542_buf_o2_p_spl_0,
    lo542_buf_o2_p_spl_
  );


  buf

  (
    n2220_o2_p_spl_,
    n2220_o2_p
  );


  buf

  (
    n2220_o2_p_spl_0,
    n2220_o2_p_spl_
  );


  buf

  (
    n2220_o2_p_spl_00,
    n2220_o2_p_spl_0
  );


  buf

  (
    n2220_o2_p_spl_01,
    n2220_o2_p_spl_0
  );


  buf

  (
    n2220_o2_p_spl_1,
    n2220_o2_p_spl_
  );


  buf

  (
    n2254_o2_n_spl_,
    n2254_o2_n
  );


  buf

  (
    n2220_o2_n_spl_,
    n2220_o2_n
  );


  buf

  (
    g928_n_spl_,
    g928_n
  );


  buf

  (
    lo478_buf_o2_p_spl_,
    lo478_buf_o2_p
  );


  buf

  (
    lo478_buf_o2_p_spl_0,
    lo478_buf_o2_p_spl_
  );


  buf

  (
    lo478_buf_o2_p_spl_00,
    lo478_buf_o2_p_spl_0
  );


  buf

  (
    lo478_buf_o2_p_spl_000,
    lo478_buf_o2_p_spl_00
  );


  buf

  (
    lo478_buf_o2_p_spl_001,
    lo478_buf_o2_p_spl_00
  );


  buf

  (
    lo478_buf_o2_p_spl_01,
    lo478_buf_o2_p_spl_0
  );


  buf

  (
    lo478_buf_o2_p_spl_010,
    lo478_buf_o2_p_spl_01
  );


  buf

  (
    lo478_buf_o2_p_spl_1,
    lo478_buf_o2_p_spl_
  );


  buf

  (
    lo478_buf_o2_p_spl_10,
    lo478_buf_o2_p_spl_1
  );


  buf

  (
    lo478_buf_o2_p_spl_11,
    lo478_buf_o2_p_spl_1
  );


  buf

  (
    n1913_inv_p_spl_,
    n1913_inv_p
  );


  buf

  (
    n1913_inv_p_spl_0,
    n1913_inv_p_spl_
  );


  buf

  (
    n1913_inv_p_spl_00,
    n1913_inv_p_spl_0
  );


  buf

  (
    n1913_inv_p_spl_1,
    n1913_inv_p_spl_
  );


  buf

  (
    lo478_buf_o2_n_spl_,
    lo478_buf_o2_n
  );


  buf

  (
    lo478_buf_o2_n_spl_0,
    lo478_buf_o2_n_spl_
  );


  buf

  (
    lo478_buf_o2_n_spl_00,
    lo478_buf_o2_n_spl_0
  );


  buf

  (
    lo478_buf_o2_n_spl_1,
    lo478_buf_o2_n_spl_
  );


  buf

  (
    lo466_buf_o2_p_spl_,
    lo466_buf_o2_p
  );


  buf

  (
    lo466_buf_o2_p_spl_0,
    lo466_buf_o2_p_spl_
  );


  buf

  (
    lo466_buf_o2_p_spl_00,
    lo466_buf_o2_p_spl_0
  );


  buf

  (
    lo466_buf_o2_p_spl_000,
    lo466_buf_o2_p_spl_00
  );


  buf

  (
    lo466_buf_o2_p_spl_001,
    lo466_buf_o2_p_spl_00
  );


  buf

  (
    lo466_buf_o2_p_spl_01,
    lo466_buf_o2_p_spl_0
  );


  buf

  (
    lo466_buf_o2_p_spl_1,
    lo466_buf_o2_p_spl_
  );


  buf

  (
    lo466_buf_o2_p_spl_10,
    lo466_buf_o2_p_spl_1
  );


  buf

  (
    lo466_buf_o2_p_spl_11,
    lo466_buf_o2_p_spl_1
  );


  buf

  (
    lo466_buf_o2_n_spl_,
    lo466_buf_o2_n
  );


  buf

  (
    lo466_buf_o2_n_spl_0,
    lo466_buf_o2_n_spl_
  );


  buf

  (
    lo466_buf_o2_n_spl_00,
    lo466_buf_o2_n_spl_0
  );


  buf

  (
    lo466_buf_o2_n_spl_000,
    lo466_buf_o2_n_spl_00
  );


  buf

  (
    lo466_buf_o2_n_spl_001,
    lo466_buf_o2_n_spl_00
  );


  buf

  (
    lo466_buf_o2_n_spl_01,
    lo466_buf_o2_n_spl_0
  );


  buf

  (
    lo466_buf_o2_n_spl_010,
    lo466_buf_o2_n_spl_01
  );


  buf

  (
    lo466_buf_o2_n_spl_011,
    lo466_buf_o2_n_spl_01
  );


  buf

  (
    lo466_buf_o2_n_spl_1,
    lo466_buf_o2_n_spl_
  );


  buf

  (
    lo466_buf_o2_n_spl_10,
    lo466_buf_o2_n_spl_1
  );


  buf

  (
    lo466_buf_o2_n_spl_100,
    lo466_buf_o2_n_spl_10
  );


  buf

  (
    lo466_buf_o2_n_spl_101,
    lo466_buf_o2_n_spl_10
  );


  buf

  (
    lo466_buf_o2_n_spl_11,
    lo466_buf_o2_n_spl_1
  );


  buf

  (
    lo466_buf_o2_n_spl_110,
    lo466_buf_o2_n_spl_11
  );


  buf

  (
    g938_n_spl_,
    g938_n
  );


  buf

  (
    g938_n_spl_0,
    g938_n_spl_
  );


  buf

  (
    n1794_lo_p_spl_,
    n1794_lo_p
  );


  buf

  (
    n2178_lo_p_spl_,
    n2178_lo_p
  );


  buf

  (
    n1926_lo_p_spl_,
    n1926_lo_p
  );


  buf

  (
    n2046_lo_p_spl_,
    n2046_lo_p
  );


  buf

  (
    n2322_lo_p_spl_,
    n2322_lo_p
  );


  buf

  (
    n2682_lo_p_spl_,
    n2682_lo_p
  );


  buf

  (
    n2442_lo_p_spl_,
    n2442_lo_p
  );


  buf

  (
    n2562_lo_p_spl_,
    n2562_lo_p
  );


  buf

  (
    n2826_lo_p_spl_,
    n2826_lo_p
  );


  buf

  (
    lo498_buf_o2_n_spl_,
    lo498_buf_o2_n
  );


  buf

  (
    lo498_buf_o2_n_spl_0,
    lo498_buf_o2_n_spl_
  );


  buf

  (
    lo498_buf_o2_n_spl_1,
    lo498_buf_o2_n_spl_
  );


  buf

  (
    g1005_n_spl_,
    g1005_n
  );


  buf

  (
    lo502_buf_o2_n_spl_,
    lo502_buf_o2_n
  );


  buf

  (
    lo502_buf_o2_n_spl_0,
    lo502_buf_o2_n_spl_
  );


  buf

  (
    g948_n_spl_,
    g948_n
  );


  buf

  (
    lo510_buf_o2_n_spl_,
    lo510_buf_o2_n
  );


  buf

  (
    lo510_buf_o2_n_spl_0,
    lo510_buf_o2_n_spl_
  );


  buf

  (
    lo510_buf_o2_n_spl_1,
    lo510_buf_o2_n_spl_
  );


  buf

  (
    g1011_n_spl_,
    g1011_n
  );


  buf

  (
    g903_n_spl_,
    g903_n
  );


  buf

  (
    g903_n_spl_0,
    g903_n_spl_
  );


  buf

  (
    g903_n_spl_1,
    g903_n_spl_
  );


  buf

  (
    n2970_lo_n_spl_,
    n2970_lo_n
  );


  buf

  (
    n2970_lo_n_spl_0,
    n2970_lo_n_spl_
  );


  buf

  (
    n2970_lo_n_spl_1,
    n2970_lo_n_spl_
  );


  buf

  (
    g1016_n_spl_,
    g1016_n
  );


  buf

  (
    g1021_n_spl_,
    g1021_n
  );


  buf

  (
    n2994_lo_n_spl_,
    n2994_lo_n
  );


  buf

  (
    n2994_lo_n_spl_0,
    n2994_lo_n_spl_
  );


  buf

  (
    n2994_lo_n_spl_1,
    n2994_lo_n_spl_
  );


  buf

  (
    g954_n_spl_,
    g954_n
  );


  buf

  (
    g919_n_spl_,
    g919_n
  );


  buf

  (
    g919_n_spl_0,
    g919_n_spl_
  );


  buf

  (
    n3006_lo_n_spl_,
    n3006_lo_n
  );


  buf

  (
    n3006_lo_n_spl_0,
    n3006_lo_n_spl_
  );


  buf

  (
    n3006_lo_n_spl_1,
    n3006_lo_n_spl_
  );


  buf

  (
    g1028_n_spl_,
    g1028_n
  );


  buf

  (
    n3018_lo_n_spl_,
    n3018_lo_n
  );


  buf

  (
    g951_n_spl_,
    g951_n
  );


  buf

  (
    g960_n_spl_,
    g960_n
  );


  buf

  (
    g957_n_spl_,
    g957_n
  );


  buf

  (
    g963_n_spl_,
    g963_n
  );


  buf

  (
    n3126_lo_p_spl_,
    n3126_lo_p
  );


  buf

  (
    n3138_lo_p_spl_,
    n3138_lo_p
  );


  buf

  (
    g919_p_spl_,
    g919_p
  );


  buf

  (
    g913_n_spl_,
    g913_n
  );


  buf

  (
    n2196_o2_p_spl_,
    n2196_o2_p
  );


  buf

  (
    n2196_o2_p_spl_0,
    n2196_o2_p_spl_
  );


  buf

  (
    n2196_o2_p_spl_1,
    n2196_o2_p_spl_
  );


  buf

  (
    g942_n_spl_,
    g942_n
  );


  buf

  (
    g968_n_spl_,
    g968_n
  );


  buf

  (
    n2386_o2_p_spl_,
    n2386_o2_p
  );


  buf

  (
    n2386_o2_p_spl_0,
    n2386_o2_p_spl_
  );


  buf

  (
    g1051_n_spl_,
    g1051_n
  );


  buf

  (
    g1051_n_spl_0,
    g1051_n_spl_
  );


  buf

  (
    g1051_n_spl_1,
    g1051_n_spl_
  );


  buf

  (
    g897_p_spl_,
    g897_p
  );


  buf

  (
    g898_p_spl_,
    g898_p
  );


  buf

  (
    g1055_n_spl_,
    g1055_n
  );


  buf

  (
    g1055_n_spl_0,
    g1055_n_spl_
  );


  buf

  (
    lo514_buf_o2_p_spl_,
    lo514_buf_o2_p
  );


  buf

  (
    g944_n_spl_,
    g944_n
  );


  buf

  (
    g945_p_spl_,
    g945_p
  );


  buf

  (
    n3030_lo_p_spl_,
    n3030_lo_p
  );


  buf

  (
    n3030_lo_n_spl_,
    n3030_lo_n
  );


  buf

  (
    n2386_o2_n_spl_,
    n2386_o2_n
  );


  buf

  (
    n2386_o2_n_spl_0,
    n2386_o2_n_spl_
  );


  buf

  (
    g1071_n_spl_,
    g1071_n
  );


  buf

  (
    g1072_p_spl_,
    g1072_p
  );


  buf

  (
    lo550_buf_o2_n_spl_,
    lo550_buf_o2_n
  );


  buf

  (
    lo550_buf_o2_n_spl_0,
    lo550_buf_o2_n_spl_
  );


  buf

  (
    g1075_n_spl_,
    g1075_n
  );


  buf

  (
    g1076_p_spl_,
    g1076_p
  );


  buf

  (
    g1079_n_spl_,
    g1079_n
  );


  buf

  (
    g1082_n_spl_,
    g1082_n
  );


  buf

  (
    n2612_o2_n_spl_,
    n2612_o2_n
  );


  buf

  (
    n2616_o2_n_spl_,
    n2616_o2_n
  );


  buf

  (
    g974_n_spl_,
    g974_n
  );


  buf

  (
    n3102_lo_p_spl_,
    n3102_lo_p
  );


  buf

  (
    n3114_lo_p_spl_,
    n3114_lo_p
  );


  buf

  (
    g929_n_spl_,
    g929_n
  );


  buf

  (
    g902_p_spl_,
    g902_p
  );


  buf

  (
    n3294_lo_n_spl_,
    n3294_lo_n
  );


  buf

  (
    n3294_lo_p_spl_,
    n3294_lo_p
  );


  buf

  (
    lo550_buf_o2_p_spl_,
    lo550_buf_o2_p
  );


  buf

  (
    lo550_buf_o2_p_spl_0,
    lo550_buf_o2_p_spl_
  );


  buf

  (
    g1099_p_spl_,
    g1099_p
  );


  buf

  (
    g1107_p_spl_,
    g1107_p
  );


  buf

  (
    g907_n_spl_,
    g907_n
  );


  buf

  (
    g980_n_spl_,
    g980_n
  );


  buf

  (
    g980_n_spl_0,
    g980_n_spl_
  );


  buf

  (
    g1112_n_spl_,
    g1112_n
  );


  buf

  (
    n3258_lo_p_spl_,
    n3258_lo_p
  );


  buf

  (
    n3270_lo_n_spl_,
    n3270_lo_n
  );


  buf

  (
    n3258_lo_n_spl_,
    n3258_lo_n
  );


  buf

  (
    n3270_lo_p_spl_,
    n3270_lo_p
  );


  buf

  (
    lo498_buf_o2_p_spl_,
    lo498_buf_o2_p
  );


  buf

  (
    lo502_buf_o2_p_spl_,
    lo502_buf_o2_p
  );


  buf

  (
    lo502_buf_o2_p_spl_0,
    lo502_buf_o2_p_spl_
  );


  buf

  (
    n2982_lo_p_spl_,
    n2982_lo_p
  );


  buf

  (
    n2994_lo_p_spl_,
    n2994_lo_p
  );


  buf

  (
    n2994_lo_p_spl_0,
    n2994_lo_p_spl_
  );


  buf

  (
    n3282_lo_n_spl_,
    n3282_lo_n
  );


  buf

  (
    n3282_lo_p_spl_,
    n3282_lo_p
  );


  buf

  (
    lo510_buf_o2_p_spl_,
    lo510_buf_o2_p
  );


  buf

  (
    n4039_o2_n_spl_,
    n4039_o2_n
  );


  buf

  (
    g1055_p_spl_,
    g1055_p
  );


  buf

  (
    lo606_buf_o2_p_spl_,
    lo606_buf_o2_p
  );


  buf

  (
    lo610_buf_o2_n_spl_,
    lo610_buf_o2_n
  );


  buf

  (
    lo606_buf_o2_n_spl_,
    lo606_buf_o2_n
  );


  buf

  (
    lo610_buf_o2_p_spl_,
    lo610_buf_o2_p
  );


  buf

  (
    lo590_buf_o2_p_spl_,
    lo590_buf_o2_p
  );


  buf

  (
    lo594_buf_o2_n_spl_,
    lo594_buf_o2_n
  );


  buf

  (
    lo590_buf_o2_n_spl_,
    lo590_buf_o2_n
  );


  buf

  (
    lo594_buf_o2_p_spl_,
    lo594_buf_o2_p
  );


  buf

  (
    g1141_p_spl_,
    g1141_p
  );


  buf

  (
    g1144_p_spl_,
    g1144_p
  );


  buf

  (
    g1141_n_spl_,
    g1141_n
  );


  buf

  (
    g1144_n_spl_,
    g1144_n
  );


  buf

  (
    n3210_lo_p_spl_,
    n3210_lo_p
  );


  buf

  (
    n3222_lo_n_spl_,
    n3222_lo_n
  );


  buf

  (
    n3210_lo_n_spl_,
    n3210_lo_n
  );


  buf

  (
    n3222_lo_p_spl_,
    n3222_lo_p
  );


  buf

  (
    g1156_n_spl_,
    g1156_n
  );


  buf

  (
    g1159_p_spl_,
    g1159_p
  );


  buf

  (
    n2539_o2_p_spl_,
    n2539_o2_p
  );


  buf

  (
    n2539_o2_n_spl_,
    n2539_o2_n
  );


  buf

  (
    n1475_inv_n_spl_,
    n1475_inv_n
  );


  buf

  (
    n2367_o2_n_spl_,
    n2367_o2_n
  );


  buf

  (
    g1164_p_spl_,
    g1164_p
  );


  buf

  (
    g1167_p_spl_,
    g1167_p
  );


  buf

  (
    g1164_n_spl_,
    g1164_n
  );


  buf

  (
    g1167_n_spl_,
    g1167_n
  );


  buf

  (
    g1051_p_spl_,
    g1051_p
  );


  buf

  (
    n3063_lo_p_spl_,
    n3063_lo_p
  );


  buf

  (
    g941_n_spl_,
    g941_n
  );


  buf

  (
    g941_n_spl_0,
    g941_n_spl_
  );


  buf

  (
    g941_n_spl_1,
    g941_n_spl_
  );


  buf

  (
    n2919_lo_p_spl_,
    n2919_lo_p
  );


  buf

  (
    g941_p_spl_,
    g941_p
  );


  buf

  (
    g941_p_spl_0,
    g941_p_spl_
  );


  buf

  (
    g941_p_spl_00,
    g941_p_spl_0
  );


  buf

  (
    g941_p_spl_1,
    g941_p_spl_
  );


  buf

  (
    g995_n_spl_,
    g995_n
  );


  buf

  (
    g995_n_spl_0,
    g995_n_spl_
  );


  buf

  (
    g1204_p_spl_,
    g1204_p
  );


  buf

  (
    lo578_buf_o2_n_spl_,
    lo578_buf_o2_n
  );


  buf

  (
    lo578_buf_o2_n_spl_0,
    lo578_buf_o2_n_spl_
  );


  buf

  (
    lo578_buf_o2_n_spl_00,
    lo578_buf_o2_n_spl_0
  );


  buf

  (
    lo578_buf_o2_n_spl_000,
    lo578_buf_o2_n_spl_00
  );


  buf

  (
    lo578_buf_o2_n_spl_001,
    lo578_buf_o2_n_spl_00
  );


  buf

  (
    lo578_buf_o2_n_spl_01,
    lo578_buf_o2_n_spl_0
  );


  buf

  (
    lo578_buf_o2_n_spl_010,
    lo578_buf_o2_n_spl_01
  );


  buf

  (
    lo578_buf_o2_n_spl_011,
    lo578_buf_o2_n_spl_01
  );


  buf

  (
    lo578_buf_o2_n_spl_1,
    lo578_buf_o2_n_spl_
  );


  buf

  (
    lo578_buf_o2_n_spl_10,
    lo578_buf_o2_n_spl_1
  );


  buf

  (
    lo578_buf_o2_n_spl_11,
    lo578_buf_o2_n_spl_1
  );


  buf

  (
    lo578_buf_o2_p_spl_,
    lo578_buf_o2_p
  );


  buf

  (
    lo578_buf_o2_p_spl_0,
    lo578_buf_o2_p_spl_
  );


  buf

  (
    lo578_buf_o2_p_spl_00,
    lo578_buf_o2_p_spl_0
  );


  buf

  (
    lo578_buf_o2_p_spl_000,
    lo578_buf_o2_p_spl_00
  );


  buf

  (
    lo578_buf_o2_p_spl_001,
    lo578_buf_o2_p_spl_00
  );


  buf

  (
    lo578_buf_o2_p_spl_01,
    lo578_buf_o2_p_spl_0
  );


  buf

  (
    lo578_buf_o2_p_spl_010,
    lo578_buf_o2_p_spl_01
  );


  buf

  (
    lo578_buf_o2_p_spl_011,
    lo578_buf_o2_p_spl_01
  );


  buf

  (
    lo578_buf_o2_p_spl_1,
    lo578_buf_o2_p_spl_
  );


  buf

  (
    lo578_buf_o2_p_spl_10,
    lo578_buf_o2_p_spl_1
  );


  buf

  (
    lo578_buf_o2_p_spl_100,
    lo578_buf_o2_p_spl_10
  );


  buf

  (
    lo578_buf_o2_p_spl_11,
    lo578_buf_o2_p_spl_1
  );


  buf

  (
    lo582_buf_o2_p_spl_,
    lo582_buf_o2_p
  );


  buf

  (
    lo582_buf_o2_p_spl_0,
    lo582_buf_o2_p_spl_
  );


  buf

  (
    lo582_buf_o2_p_spl_1,
    lo582_buf_o2_p_spl_
  );


  buf

  (
    lo582_buf_o2_n_spl_,
    lo582_buf_o2_n
  );


  buf

  (
    lo582_buf_o2_n_spl_0,
    lo582_buf_o2_n_spl_
  );


  buf

  (
    g1040_n_spl_,
    g1040_n
  );


  buf

  (
    g1183_n_spl_,
    g1183_n
  );


  buf

  (
    n3075_lo_p_spl_,
    n3075_lo_p
  );


  buf

  (
    n2943_lo_p_spl_,
    n2943_lo_p
  );


  buf

  (
    n3087_lo_p_spl_,
    n3087_lo_p
  );


  buf

  (
    n2955_lo_p_spl_,
    n2955_lo_p
  );


  buf

  (
    n3039_lo_p_spl_,
    n3039_lo_p
  );


  buf

  (
    n2907_lo_p_spl_,
    n2907_lo_p
  );


  buf

  (
    g986_n_spl_,
    g986_n
  );


  buf

  (
    lo576_buf_o2_p_spl_,
    lo576_buf_o2_p
  );


  buf

  (
    lo576_buf_o2_p_spl_0,
    lo576_buf_o2_p_spl_
  );


  buf

  (
    lo576_buf_o2_p_spl_00,
    lo576_buf_o2_p_spl_0
  );


  buf

  (
    lo576_buf_o2_p_spl_1,
    lo576_buf_o2_p_spl_
  );


  buf

  (
    lo576_buf_o2_n_spl_,
    lo576_buf_o2_n
  );


  buf

  (
    lo576_buf_o2_n_spl_0,
    lo576_buf_o2_n_spl_
  );


  buf

  (
    lo576_buf_o2_n_spl_1,
    lo576_buf_o2_n_spl_
  );


  buf

  (
    n3156_lo_n_spl_,
    n3156_lo_n
  );


  buf

  (
    n3156_lo_p_spl_,
    n3156_lo_p
  );


  buf

  (
    n3156_lo_p_spl_0,
    n3156_lo_p_spl_
  );


  buf

  (
    n2808_lo_n_spl_,
    n2808_lo_n
  );


  buf

  (
    n2808_lo_p_spl_,
    n2808_lo_p
  );


  buf

  (
    n2808_lo_p_spl_0,
    n2808_lo_p_spl_
  );


  buf

  (
    g1284_n_spl_,
    g1284_n
  );


  buf

  (
    g1288_n_spl_,
    g1288_n
  );


  buf

  (
    n2901_lo_n_spl_,
    n2901_lo_n
  );


  buf

  (
    n3057_lo_n_spl_,
    n3057_lo_n
  );


  buf

  (
    n3057_lo_n_spl_0,
    n3057_lo_n_spl_
  );


  buf

  (
    g742_n_spl_,
    g742_n
  );


  buf

  (
    g758_p_spl_,
    g758_p
  );


  buf

  (
    g761_n_spl_,
    g761_n
  );


  buf

  (
    g766_p_spl_,
    g766_p
  );


  buf

  (
    g838_n_spl_,
    g838_n
  );


  buf

  (
    g859_p_spl_,
    g859_p
  );


  buf

  (
    g895_n_spl_,
    g895_n
  );


endmodule
