// Benchmark "mymod" written by ABC on Sun Oct 29 23:44:40 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G58,
    G59, G60,
    G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, G865, G866,
    G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, G877, G878,
    G879, G880  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G58, G59, G60;
  output G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, G865,
    G866, G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, G877,
    G878, G879, G880;
  reg n492_lo, n495_lo, n498_lo, n501_lo, n516_lo, n528_lo, n540_lo,
    n543_lo, n546_lo, n549_lo, n552_lo, n564_lo, n600_lo, n603_lo, n606_lo,
    n609_lo, n615_lo, n618_lo, n621_lo, n627_lo, n630_lo, n633_lo, n639_lo,
    n642_lo, n645_lo, n648_lo, n660_lo, n672_lo, n675_lo, n678_lo, n681_lo,
    n684_lo, n687_lo, n690_lo, n693_lo, n696_lo, n699_lo, n702_lo, n705_lo,
    n708_lo, n711_lo, n714_lo, n717_lo, n720_lo, n723_lo, n726_lo, n729_lo,
    n732_lo, n735_lo, n738_lo, n741_lo, n744_lo, n747_lo, n750_lo, n753_lo,
    n756_lo, n759_lo, n762_lo, n765_lo, n768_lo, n771_lo, n774_lo, n777_lo,
    n780_lo, n783_lo, n786_lo, n792_lo, n795_lo, n798_lo, n807_lo, n816_lo,
    n819_lo, n828_lo, n831_lo, n843_lo, n846_lo, n849_lo, n852_lo, n855_lo,
    n858_lo, n861_lo, n864_lo, n867_lo, n870_lo, n879_lo, n882_lo, n891_lo,
    n903_lo, n915_lo, n918_lo, n951_lo, n954_lo, n957_lo, n960_lo, n963_lo,
    n966_lo, n969_lo, n972_lo, n975_lo, n978_lo, n981_lo, n984_lo, n987_lo,
    n990_lo, n993_lo, n996_lo, n999_lo, n1002_lo, n1008_lo, n1011_lo,
    n1014_lo, n1020_lo, n1023_lo, n1032_lo, n1035_lo, n1044_lo, n1047_lo,
    n1050_lo, n1053_lo, n1056_lo, n1059_lo, n1062_lo, n1065_lo, n1068_lo,
    n1071_lo, n1074_lo, n1077_lo, n1080_lo, n1083_lo, n1086_lo, n1089_lo,
    n1092_lo, n1095_lo, n1098_lo, n1101_lo, n1104_lo, n1107_lo, n1110_lo,
    n1113_lo, n1116_lo, n1119_lo, n1122_lo, n1125_lo, n1128_lo, n1131_lo,
    n1134_lo, n1137_lo, n1143_lo, n1146_lo, n1149_lo, n1152_lo, n1155_lo,
    n1164_lo, n1167_lo, n1170_lo, n1173_lo, n1176_lo, n1188_lo, n563_inv,
    n1429_o2, n1427_o2, n1471_o2, n1476_o2, n1499_o2, n1500_o2, n1501_o2,
    n1516_o2, n1517_o2, n1562_o2, n1563_o2, n1564_o2, n1582_o2, n1583_o2,
    n1618_o2, n1622_o2, n1502_o2, n1503_o2, n1504_o2, n1505_o2, n1506_o2,
    n1512_o2, n1513_o2, n1514_o2, n1515_o2, n1644_o2, n1647_o2, n1527_o2,
    n650_inv, n653_inv, n656_inv, n1567_o2, n955_o2, n1568_o2, n1037_o2,
    n960_o2, n1587_o2, n1040_o2, n1039_o2, n1589_o2, n1624_o2, n1643_o2,
    n1038_o2, n1645_o2, n1029_o2, n701_inv, n1662_o2, n1663_o2, n710_inv,
    n813_o2, lo114_buf_o2, n1031_o2, lo186_buf_o2, n1042_o2, n728_inv,
    n917_o2, n734_inv, n1649_o2, n1650_o2, n1651_o2, n1652_o2, n1653_o2,
    lo138_buf_o2, n1664_o2, n1665_o2, n1666_o2, n1667_o2, n944_o2,
    n770_inv, n1672_o2, n776_inv, n1679_o2, n782_inv, n785_inv,
    lo110_buf_o2, lo134_buf_o2, n1030_o2, lo182_buf_o2, n830_o2, n1021_o2,
    n806_inv, n809_inv, n946_o2, lo038_buf_o2, lo238_buf_o2, n1010_o2,
    n1006_o2, n907_o2, n902_o2, lo154_buf_o2, n836_inv, n839_inv,
    lo122_buf_o2, n845_inv, n904_o2, lo106_buf_o2, n980_o2, n1023_o2,
    lo178_buf_o2, n981_o2, n837_o2, n1013_o2, n840_o2, n849_o2, n852_o2,
    n864_o2, n867_o2, n1044_o2, n876_o2, n893_inv, n879_o2, n925_o2,
    n902_inv, lo146_buf_o2, n1026_o2, n1032_o2, lo118_buf_o2, n917_inv,
    lo190_buf_o2, n1036_o2, n926_inv, n929_inv, lo002_buf_o2, lo014_buf_o2,
    lo030_buf_o2, lo034_buf_o2, lo042_buf_o2, lo113_buf_o2, lo185_buf_o2,
    n939_o2, n941_o2, lo142_buf_o2, lo230_buf_o2, lo006_buf_o2,
    lo018_buf_o2, lo022_buf_o2, lo066_buf_o2, n977_inv, n826_o2, n892_o2,
    lo152_buf_o2, n896_o2, n905_o2, n995_inv, lo037_buf_o2, lo237_buf_o2,
    lo062_buf_o2, n1007_inv, n1010_inv, n891_o2;
  wire new_new_n705__, new_new_n706__, new_new_n707__, new_new_n709__,
    new_new_n711__, new_new_n712__, new_new_n713__, new_new_n714__,
    new_new_n715__, new_new_n717__, new_new_n719__, new_new_n720__,
    new_new_n721__, new_new_n722__, new_new_n723__, new_new_n725__,
    new_new_n726__, new_new_n727__, new_new_n729__, new_new_n731__,
    new_new_n733__, new_new_n735__, new_new_n737__, new_new_n739__,
    new_new_n741__, new_new_n743__, new_new_n745__, new_new_n747__,
    new_new_n749__, new_new_n751__, new_new_n753__, new_new_n755__,
    new_new_n757__, new_new_n759__, new_new_n761__, new_new_n763__,
    new_new_n765__, new_new_n767__, new_new_n769__, new_new_n771__,
    new_new_n773__, new_new_n775__, new_new_n777__, new_new_n779__,
    new_new_n781__, new_new_n784__, new_new_n785__, new_new_n787__,
    new_new_n789__, new_new_n791__, new_new_n793__, new_new_n795__,
    new_new_n797__, new_new_n799__, new_new_n801__, new_new_n803__,
    new_new_n805__, new_new_n807__, new_new_n809__, new_new_n811__,
    new_new_n813__, new_new_n815__, new_new_n817__, new_new_n819__,
    new_new_n821__, new_new_n823__, new_new_n826__, new_new_n827__,
    new_new_n829__, new_new_n832__, new_new_n834__, new_new_n836__,
    new_new_n837__, new_new_n838__, new_new_n839__, new_new_n841__,
    new_new_n843__, new_new_n845__, new_new_n846__, new_new_n847__,
    new_new_n848__, new_new_n850__, new_new_n851__, new_new_n853__,
    new_new_n856__, new_new_n857__, new_new_n859__, new_new_n862__,
    new_new_n863__, new_new_n865__, new_new_n868__, new_new_n869__,
    new_new_n871__, new_new_n873__, new_new_n876__, new_new_n878__,
    new_new_n880__, new_new_n881__, new_new_n883__, new_new_n885__,
    new_new_n888__, new_new_n889__, new_new_n891__, new_new_n893__,
    new_new_n896__, new_new_n897__, new_new_n899__, new_new_n901__,
    new_new_n903__, new_new_n905__, new_new_n907__, new_new_n909__,
    new_new_n911__, new_new_n913__, new_new_n915__, new_new_n917__,
    new_new_n919__, new_new_n921__, new_new_n923__, new_new_n925__,
    new_new_n927__, new_new_n929__, new_new_n931__, new_new_n933__,
    new_new_n934__, new_new_n936__, new_new_n937__, new_new_n939__,
    new_new_n941__, new_new_n942__, new_new_n944__, new_new_n945__,
    new_new_n947__, new_new_n949__, new_new_n950__, new_new_n952__,
    new_new_n953__, new_new_n955__, new_new_n958__, new_new_n959__,
    new_new_n961__, new_new_n963__, new_new_n966__, new_new_n967__,
    new_new_n970__, new_new_n971__, new_new_n973__, new_new_n975__,
    new_new_n977__, new_new_n979__, new_new_n980__, new_new_n981__,
    new_new_n983__, new_new_n985__, new_new_n987__, new_new_n988__,
    new_new_n989__, new_new_n991__, new_new_n992__, new_new_n993__,
    new_new_n995__, new_new_n997__, new_new_n999__, new_new_n1001__,
    new_new_n1004__, new_new_n1005__, new_new_n1007__, new_new_n1009__,
    new_new_n1010__, new_new_n1011__, new_new_n1012__, new_new_n1013__,
    new_new_n1015__, new_new_n1017__, new_new_n1018__, new_new_n1019__,
    new_new_n1020__, new_new_n1021__, new_new_n1023__, new_new_n1025__,
    new_new_n1026__, new_new_n1028__, new_new_n1029__, new_new_n1031__,
    new_new_n1033__, new_new_n1034__, new_new_n1036__, new_new_n1037__,
    new_new_n1039__, new_new_n1042__, new_new_n1043__, new_new_n1045__,
    new_new_n1046__, new_new_n1048__, new_new_n1049__, new_new_n1052__,
    new_new_n1053__, new_new_n1056__, new_new_n1057__, new_new_n1059__,
    new_new_n1061__, new_new_n1063__, new_new_n1064__, new_new_n1065__,
    new_new_n1067__, new_new_n1069__, new_new_n1072__, new_new_n1073__,
    new_new_n1075__, new_new_n1077__, new_new_n1080__, new_new_n1081__,
    new_new_n1083__, new_new_n1085__, new_new_n1088__, new_new_n1089__,
    new_new_n1091__, new_new_n1093__, new_new_n1096__, new_new_n1097__,
    new_new_n1099__, new_new_n1101__, new_new_n1104__, new_new_n1105__,
    new_new_n1107__, new_new_n1109__, new_new_n1112__, new_new_n1113__,
    new_new_n1115__, new_new_n1117__, new_new_n1119__, new_new_n1121__,
    new_new_n1123__, new_new_n1126__, new_new_n1127__, new_new_n1130__,
    new_new_n1131__, new_new_n1133__, new_new_n1135__, new_new_n1138__,
    new_new_n1140__, new_new_n1142__, new_new_n1144__, new_new_n1145__,
    new_new_n1148__, new_new_n1150__, new_new_n1151__, new_new_n1152__,
    new_new_n1153__, new_new_n1156__, new_new_n1158__, new_new_n1160__,
    new_new_n1161__, new_new_n1162__, new_new_n1164__, new_new_n1165__,
    new_new_n1167__, new_new_n1168__, new_new_n1169__, new_new_n1170__,
    new_new_n1171__, new_new_n1172__, new_new_n1174__, new_new_n1176__,
    new_new_n1177__, new_new_n1179__, new_new_n1181__, new_new_n1183__,
    new_new_n1185__, new_new_n1186__, new_new_n1187__, new_new_n1189__,
    new_new_n1191__, new_new_n1194__, new_new_n1196__, new_new_n1197__,
    new_new_n1199__, new_new_n1200__, new_new_n1201__, new_new_n1203__,
    new_new_n1206__, new_new_n1207__, new_new_n1208__, new_new_n1209__,
    new_new_n1212__, new_new_n1213__, new_new_n1215__, new_new_n1216__,
    new_new_n1217__, new_new_n1218__, new_new_n1219__, new_new_n1220__,
    new_new_n1221__, new_new_n1222__, new_new_n1224__, new_new_n1225__,
    new_new_n1226__, new_new_n1227__, new_new_n1228__, new_new_n1229__,
    new_new_n1230__, new_new_n1232__, new_new_n1233__, new_new_n1235__,
    new_new_n1237__, new_new_n1239__, new_new_n1242__, new_new_n1243__,
    new_new_n1244__, new_new_n1245__, new_new_n1246__, new_new_n1247__,
    new_new_n1248__, new_new_n1249__, new_new_n1250__, new_new_n1251__,
    new_new_n1253__, new_new_n1255__, new_new_n1257__, new_new_n1259__,
    new_new_n1260__, new_new_n1261__, new_new_n1263__, new_new_n1265__,
    new_new_n1267__, new_new_n1269__, new_new_n1271__, new_new_n1273__,
    new_new_n1275__, new_new_n1277__, new_new_n1279__, new_new_n1281__,
    new_new_n1283__, new_new_n1285__, new_new_n1287__, new_new_n1288__,
    new_new_n1289__, new_new_n1291__, new_new_n1292__, new_new_n1293__,
    new_new_n1295__, new_new_n1296__, new_new_n1297__, new_new_n1298__,
    new_new_n1300__, new_new_n1301__, new_new_n1302__, new_new_n1303__,
    new_new_n1305__, new_new_n1307__, new_new_n1309__, new_new_n1310__,
    new_new_n1311__, new_new_n1313__, new_new_n1314__, new_new_n1315__,
    new_new_n1316__, new_new_n1317__, new_new_n1318__, new_new_n1320__,
    new_new_n1322__, new_new_n1323__, new_new_n1325__, new_new_n1327__,
    new_new_n1329__, new_new_n1330__, new_new_n1331__, new_new_n1332__,
    new_new_n1333__, new_new_n1334__, new_new_n1336__, new_new_n1337__,
    new_new_n1338__, new_new_n1339__, new_new_n1340__, new_new_n1342__,
    new_new_n1343__, new_new_n1344__, new_new_n1345__, new_new_n1346__,
    new_new_n1347__, new_new_n1348__, new_new_n1349__, new_new_n1350__,
    new_new_n1351__, new_new_n1352__, new_new_n1353__, new_new_n1354__,
    new_new_n1355__, new_new_n1356__, new_new_n1357__, new_new_n1358__,
    new_new_n1359__, new_new_n1360__, new_new_n1361__, new_new_n1363__,
    new_new_n1364__, new_new_n1366__, new_new_n1367__, new_new_n1368__,
    new_new_n1369__, new_new_n1372__, new_new_n1374__, new_new_n1375__,
    new_new_n1377__, new_new_n1378__, new_new_n1379__, new_new_n1380__,
    new_new_n1382__, new_new_n1383__, new_new_n1384__, new_new_n1385__,
    new_new_n1386__, new_new_n1387__, new_new_n1388__, new_new_n1389__,
    new_new_n1391__, new_new_n1393__, new_new_n1395__, new_new_n1397__,
    new_new_n1398__, new_new_n1399__, new_new_n1400__, new_new_n1402__,
    new_new_n1404__, new_new_n1405__, new_new_n1406__, new_new_n1407__,
    new_new_n1408__, new_new_n1409__, new_new_n1411__, new_new_n1413__,
    new_new_n1415__, new_new_n1417__, new_new_n1418__, new_new_n1419__,
    new_new_n1421__, new_new_n1423__, new_new_n1425__, new_new_n1427__,
    new_new_n1429__, new_new_n1430__, new_new_n1431__, new_new_n1433__,
    new_new_n1434__, new_new_n1435__, new_new_n1436__, new_new_n1437__,
    new_new_n1439__, new_new_n1441__, new_new_n1443__, new_new_n1444__,
    new_new_n1445__, new_new_n1446__, new_new_n1447__, new_new_n1448__,
    new_new_n1449__, new_new_n1450__, new_new_n1451__, new_new_n1452__,
    new_new_n1453__, new_new_n1454__, new_new_n1455__, new_new_n1456__,
    new_new_n1457__, new_new_n1458__, new_new_n1459__, new_new_n1460__,
    new_new_n1461__, new_new_n1462__, new_new_n1463__, new_new_n1464__,
    new_new_n1465__, new_new_n1466__, new_new_n1467__, new_new_n1468__,
    new_new_n1469__, new_new_n1470__, new_new_n1471__, new_new_n1472__,
    new_new_n1473__, new_new_n1474__, new_new_n1475__, new_new_n1476__,
    new_new_n1477__, new_new_n1478__, new_new_n1479__, new_new_n1480__,
    new_new_n1481__, new_new_n1482__, new_new_n1483__, new_new_n1484__,
    new_new_n1485__, new_new_n1486__, new_new_n1487__, new_new_n1488__,
    new_new_n1489__, new_new_n1490__, new_new_n1491__, new_new_n1492__,
    new_new_n1493__, new_new_n1494__, new_new_n1495__, new_new_n1496__,
    new_new_n1497__, new_new_n1498__, new_new_n1499__, new_new_n1500__,
    new_new_n1501__, new_new_n1502__, new_new_n1503__, new_new_n1504__,
    new_new_n1505__, new_new_n1506__, new_new_n1507__, new_new_n1508__,
    new_new_n1509__, new_new_n1510__, new_new_n1511__, new_new_n1512__,
    new_new_n1513__, new_new_n1514__, new_new_n1515__, new_new_n1516__,
    new_new_n1517__, new_new_n1518__, new_new_n1519__, new_new_n1520__,
    new_new_n1521__, new_new_n1522__, new_new_n1523__, new_new_n1524__,
    new_new_n1525__, new_new_n1526__, new_new_n1527__, new_new_n1528__,
    new_new_n1529__, new_new_n1530__, new_new_n1531__, new_new_n1532__,
    new_new_n1533__, new_new_n1534__, new_new_n1535__, new_new_n1536__,
    new_new_n1537__, new_new_n1538__, new_new_n1539__, new_new_n1540__,
    new_new_n1541__, new_new_n1542__, new_new_n1543__, new_new_n1544__,
    new_new_n1545__, new_new_n1546__, new_new_n1547__, new_new_n1548__,
    new_new_n1549__, new_new_n1550__, new_new_n1551__, new_new_n1552__,
    new_new_n1553__, new_new_n1554__, new_new_n1555__, new_new_n1556__,
    new_new_n1557__, new_new_n1558__, new_new_n1559__, new_new_n1560__,
    new_new_n1561__, new_new_n1562__, new_new_n1563__, new_new_n1564__,
    new_new_n1565__, new_new_n1566__, new_new_n1567__, new_new_n1568__,
    new_new_n1569__, new_new_n1570__, new_new_n1571__, new_new_n1572__,
    new_new_n1573__, new_new_n1574__, new_new_n1575__, new_new_n1576__,
    new_new_n1577__, new_new_n1578__, new_new_n1579__, new_new_n1580__,
    new_new_n1581__, new_new_n1582__, new_new_n1583__, new_new_n1584__,
    new_new_n1585__, new_new_n1586__, new_new_n1587__, new_new_n1588__,
    new_new_n1589__, new_new_n1590__, new_new_n1591__, new_new_n1592__,
    new_new_n1593__, new_new_n1594__, new_new_n1595__, new_new_n1596__,
    new_new_n1597__, new_new_n1598__, new_new_n1599__, new_new_n1600__,
    new_new_n1601__, new_new_n1602__, new_new_n1603__, new_new_n1604__,
    new_new_n1605__, new_new_n1606__, new_new_n1607__, new_new_n1608__,
    new_new_n1609__, new_new_n1610__, new_new_n1611__, new_new_n1612__,
    new_new_n1613__, new_new_n1614__, new_new_n1615__, new_new_n1616__,
    new_new_n1617__, new_new_n1618__, new_new_n1619__, new_new_n1620__,
    new_new_n1621__, new_new_n1622__, new_new_n1623__, new_new_n1624__,
    new_new_n1625__, new_new_n1626__, new_new_n1627__, new_new_n1628__,
    new_new_n1629__, new_new_n1630__, new_new_n1631__, new_new_n1632__,
    new_new_n1633__, new_new_n1634__, new_new_n1635__, new_new_n1636__,
    new_new_n1637__, new_new_n1638__, new_new_n1639__, new_new_n1640__,
    new_new_n1641__, new_new_n1642__, new_new_n1643__, new_new_n1644__,
    new_new_n1645__, new_new_n1646__, new_new_n1647__, new_new_n1648__,
    new_new_n1649__, new_new_n1650__, new_new_n1651__, new_new_n1652__,
    new_new_n1653__, new_new_n1654__, new_new_n1655__, new_new_n1656__,
    new_new_n1657__, new_new_n1658__, new_new_n1659__, new_new_n1660__,
    new_new_n1661__, new_new_n1662__, new_new_n1663__, new_new_n1664__,
    new_new_n1665__, new_new_n1666__, new_new_n1667__, new_new_n1668__,
    new_new_n1669__, new_new_n1670__, new_new_n1671__, new_new_n1672__,
    new_new_n1673__, new_new_n1674__, new_new_n1675__, new_new_n1676__,
    new_new_n1677__, new_new_n1678__, new_new_n1679__, new_new_n1680__,
    new_new_n1681__, new_new_n1682__, new_new_n1683__, new_new_n1684__,
    new_new_n1685__, new_new_n1686__, new_new_n1687__, new_new_n1688__,
    new_new_n1689__, new_new_n1690__, new_new_n1691__, new_new_n1692__,
    new_new_n1693__, new_new_n1694__, new_new_n1695__, new_new_n1696__,
    new_new_n1697__, new_new_n1698__, new_new_n1699__, new_new_n1700__,
    new_new_n1701__, new_new_n1702__, new_new_n1703__, new_new_n1704__,
    new_new_n1705__, new_new_n1706__, new_new_n1707__, new_new_n1708__,
    new_new_n1709__, new_new_n1710__, new_new_n1711__, new_new_n1712__,
    new_new_n1713__, new_new_n1714__, new_new_n1715__, new_new_n1716__,
    new_new_n1717__, new_new_n1718__, new_new_n1719__, new_new_n1720__,
    new_new_n1721__, new_new_n1722__, new_new_n1723__, new_new_n1724__,
    new_new_n1725__, new_new_n1726__, new_new_n1727__, new_new_n1728__,
    new_new_n1729__, new_new_n1730__, new_new_n1731__, new_new_n1732__,
    new_new_n1733__, new_new_n1734__, new_new_n1735__, new_new_n1736__,
    new_new_n1737__, new_new_n1738__, new_new_n1739__, new_new_n1740__,
    new_new_n1741__, new_new_n1742__, new_new_n1743__, new_new_n1744__,
    new_new_n1745__, new_new_n1746__, new_new_n1747__, new_new_n1748__,
    new_new_n1749__, new_new_n1750__, new_new_n1751__, new_new_n1752__,
    new_new_n1753__, new_new_n1754__, new_new_n1755__, new_new_n1756__,
    new_new_n1757__, new_new_n1758__, new_new_n1759__, new_new_n1760__,
    new_new_n1761__, new_new_n1762__, new_new_n1763__, new_new_n1764__,
    new_new_n1765__, new_new_n1766__, new_new_n1767__, new_new_n1768__,
    new_new_n1769__, new_new_n1770__, new_new_n1771__, new_new_n1772__,
    new_new_n1773__, new_new_n1774__, new_new_n1775__, new_new_n1776__,
    new_new_n1777__, new_new_n1778__, new_new_n1779__, new_new_n1780__,
    new_new_n2116__, new_new_n2117__, new_new_n2118__, new_new_n2119__,
    new_new_n2120__, new_new_n2121__, new_new_n2122__, new_new_n2123__,
    new_new_n2124__, new_new_n2125__, new_new_n2126__, new_new_n2127__,
    new_new_n2128__, new_new_n2129__, new_new_n2130__, new_new_n2131__,
    new_new_n2132__, new_new_n2133__, new_new_n2134__, new_new_n2135__,
    new_new_n2136__, new_new_n2137__, new_new_n2138__, new_new_n2139__,
    new_new_n2140__, new_new_n2141__, new_new_n2142__, new_new_n2143__,
    new_new_n2144__, new_new_n2145__, new_new_n2146__, new_new_n2147__,
    new_new_n2148__, new_new_n2149__, new_new_n2150__, new_new_n2151__,
    new_new_n2152__, new_new_n2153__, new_new_n2154__, new_new_n2155__,
    new_new_n2156__, new_new_n2157__, new_new_n2158__, new_new_n2159__,
    new_new_n2160__, new_new_n2161__, new_new_n2162__, new_new_n2163__,
    new_new_n2164__, new_new_n2165__, new_new_n2166__, new_new_n2167__,
    new_new_n2168__, new_new_n2169__, new_new_n2170__, new_new_n2171__,
    new_new_n2172__, new_new_n2173__, new_new_n2174__, new_new_n2175__,
    new_new_n2176__, new_new_n2177__, new_new_n2178__, new_new_n2179__,
    new_new_n2180__, new_new_n2181__, new_new_n2182__, new_new_n2183__,
    new_new_n2184__, new_new_n2185__, new_new_n2186__, new_new_n2187__,
    new_new_n2188__, new_new_n2189__, new_new_n2190__, new_new_n2191__,
    new_new_n2192__, new_new_n2193__, new_new_n2194__, new_new_n2195__,
    new_new_n2196__, new_new_n2197__, new_new_n2198__, new_new_n2199__,
    new_new_n2200__, new_new_n2201__, new_new_n2202__, new_new_n2203__,
    new_new_n2204__, new_new_n2205__, new_new_n2206__, new_new_n2207__,
    new_new_n2208__, new_new_n2209__, new_new_n2210__, new_new_n2211__,
    new_new_n2212__, new_new_n2213__, new_new_n2214__, new_new_n2215__,
    new_new_n2216__, new_new_n2217__, new_new_n2218__, new_new_n2219__,
    new_new_n2220__, new_new_n2221__, new_new_n2222__, new_new_n2223__,
    new_new_n2224__, new_new_n2225__, new_new_n2226__, new_new_n2227__,
    new_new_n2228__, new_new_n2229__, new_new_n2230__, new_new_n2231__,
    new_new_n2232__, new_new_n2233__, new_new_n2234__, new_new_n2235__,
    new_new_n2236__, new_new_n2237__, new_new_n2238__, new_new_n2239__,
    new_new_n2240__, new_new_n2241__, new_new_n2242__, new_new_n2243__,
    new_new_n2244__, new_new_n2245__, new_new_n2246__, new_new_n2247__,
    new_new_n2248__, new_new_n2249__, new_new_n2250__, new_new_n2251__,
    new_new_n2252__, new_new_n2253__, new_new_n2254__, new_new_n2255__,
    new_new_n2256__, new_new_n2257__, new_new_n2258__, new_new_n2259__,
    new_new_n2260__, new_new_n2261__, new_new_n2262__, new_new_n2263__,
    new_new_n2264__, new_new_n2265__, new_new_n2266__, new_new_n2267__,
    new_new_n2268__, new_new_n2269__, new_new_n2270__, new_new_n2271__,
    new_new_n2272__, new_new_n2273__, new_new_n2274__, new_new_n2275__,
    new_new_n2276__, new_new_n2277__, new_new_n2278__, new_new_n2279__,
    new_new_n2280__, new_new_n2281__, new_new_n2282__, new_new_n2283__,
    new_new_n2284__, new_new_n2285__, new_new_n2286__, new_new_n2287__,
    new_new_n2288__, new_new_n2289__, new_new_n2290__, new_new_n2291__,
    new_new_n2292__, new_new_n2293__, new_new_n2294__, new_new_n2295__,
    new_new_n2296__, new_new_n2297__, new_new_n2298__, new_new_n2299__,
    new_new_n2300__, new_new_n2301__, new_new_n2302__, new_new_n2303__,
    new_new_n2304__, new_new_n2305__, new_new_n2306__, new_new_n2307__,
    new_new_n2308__, new_new_n2309__, new_new_n2310__, new_new_n2311__,
    new_new_n2312__, new_new_n2313__, new_new_n2314__, new_new_n2315__,
    new_new_n2316__, new_new_n2317__, new_new_n2318__, new_new_n2319__,
    new_new_n2320__, new_new_n2321__, new_new_n2322__, new_new_n2323__,
    new_new_n2324__, new_new_n2325__, new_new_n2326__, new_new_n2327__,
    new_new_n2328__, new_new_n2329__, new_new_n2330__, new_new_n2331__,
    new_new_n2332__, new_new_n2333__, new_new_n2334__, new_new_n2335__,
    new_new_n2336__, new_new_n2337__, new_new_n2338__, n3148, n3151, n3154,
    n3157, n3160, n3163, n3166, n3169, n3172, n3175, n3178, n3181, n3184,
    n3187, n3190, n3193, n3196, n3199, n3202, n3205, n3208, n3211, n3214,
    n3217, n3220, n3223, n3226, n3229, n3232, n3235, n3238, n3241, n3244,
    n3247, n3250, n3253, n3256, n3259, n3262, n3265, n3268, n3271, n3274,
    n3277, n3280, n3283, n3286, n3289, n3292, n3295, n3298, n3301, n3304,
    n3307, n3310, n3313, n3316, n3319, n3322, n3325, n3328, n3331, n3334,
    n3337, n3340, n3343, n3346, n3349, n3352, n3355, n3358, n3361, n3364,
    n3367, n3370, n3373, n3376, n3379, n3382, n3385, n3388, n3391, n3394,
    n3397, n3400, n3403, n3406, n3409, n3412, n3415, n3418, n3421, n3424,
    n3427, n3430, n3433, n3436, n3439, n3442, n3445, n3448, n3451, n3454,
    n3457, n3460, n3463, n3466, n3469, n3472, n3475, n3478, n3481, n3484,
    n3487, n3490, n3493, n3496, n3499, n3502, n3505, n3508, n3511, n3514,
    n3517, n3520, n3523, n3526, n3529, n3532, n3535, n3538, n3541, n3544,
    n3547, n3550, n3553, n3556, n3559, n3562, n3565, n3568, n3571, n3574,
    n3577, n3580, n3583, n3586, n3589, n3592, n3595, n3598, n3601, n3604,
    n3607, n3610, n3613, n3616, n3619, n3622, n3625, n3628, n3631, n3634,
    n3637, n3640, n3643, n3646, n3649, n3652, n3655, n3658, n3661, n3664,
    n3667, n3670, n3673, n3676, n3679, n3682, n3685, n3688, n3691, n3694,
    n3697, n3700, n3703, n3706, n3709, n3712, n3715, n3718, n3721, n3724,
    n3727, n3730, n3733, n3736, n3739, n3742, n3745, n3748, n3751, n3754,
    n3757, n3760, n3763, n3766, n3769, n3772, n3775, n3778, n3781, n3784,
    n3787, n3790, n3793, n3796, n3799, n3802, n3805, n3808, n3811, n3814,
    n3817, n3820, n3823, n3826, n3829, n3832, n3835, n3838, n3841, n3844,
    n3847, n3850, n3853, n3856, n3859, n3862, n3865, n3868, n3871, n3874,
    n3877, n3880, n3883, n3886, n3889, n3892, n3895, n3898, n3901, n3904,
    n3907, n3910, n3913, n3916, n3919, n3922, n3925, n3928, n3931, n3934,
    n3937, n3940, n3943, n3946, n3949, n3952, n3955, n3958, n3961, n3964,
    n3967, n3970, n3973, n3976, n3979, n3982, n3985, n3988, n3991, n3994,
    n3997, n4000, n4003, n4006, n4009, n4012, n4015, n4018, n4021, n4024,
    n4027, n4030, n4033, n4036, n4039, n4042, n4045, n4048, n4051, n4054,
    n4057, n4060, n4063, n4066, n4069, n4072;
  buf1  g0000(.din(G1), .dout(new_new_n705__));
  not1  g0001(.din(G1), .dout(new_new_n706__));
  buf1  g0002(.din(G2), .dout(new_new_n707__));
  buf1  g0003(.din(G3), .dout(new_new_n709__));
  buf1  g0004(.din(G4), .dout(new_new_n711__));
  not1  g0005(.din(G4), .dout(new_new_n712__));
  buf1  g0006(.din(G5), .dout(new_new_n713__));
  not1  g0007(.din(G5), .dout(new_new_n714__));
  buf1  g0008(.din(G6), .dout(new_new_n715__));
  buf1  g0009(.din(G7), .dout(new_new_n717__));
  buf1  g0010(.din(G8), .dout(new_new_n719__));
  not1  g0011(.din(G8), .dout(new_new_n720__));
  buf1  g0012(.din(G9), .dout(new_new_n721__));
  not1  g0013(.din(G9), .dout(new_new_n722__));
  buf1  g0014(.din(G10), .dout(new_new_n723__));
  buf1  g0015(.din(G11), .dout(new_new_n725__));
  not1  g0016(.din(G11), .dout(new_new_n726__));
  buf1  g0017(.din(G12), .dout(new_new_n727__));
  buf1  g0018(.din(G13), .dout(new_new_n729__));
  buf1  g0019(.din(G14), .dout(new_new_n731__));
  buf1  g0020(.din(G15), .dout(new_new_n733__));
  buf1  g0021(.din(G16), .dout(new_new_n735__));
  buf1  g0022(.din(G17), .dout(new_new_n737__));
  buf1  g0023(.din(G18), .dout(new_new_n739__));
  buf1  g0024(.din(G19), .dout(new_new_n741__));
  buf1  g0025(.din(G20), .dout(new_new_n743__));
  buf1  g0026(.din(G21), .dout(new_new_n745__));
  buf1  g0027(.din(G22), .dout(new_new_n747__));
  buf1  g0028(.din(G23), .dout(new_new_n749__));
  buf1  g0029(.din(G24), .dout(new_new_n751__));
  buf1  g0030(.din(G25), .dout(new_new_n753__));
  buf1  g0031(.din(G26), .dout(new_new_n755__));
  buf1  g0032(.din(G27), .dout(new_new_n757__));
  buf1  g0033(.din(G28), .dout(new_new_n759__));
  buf1  g0034(.din(G29), .dout(new_new_n761__));
  buf1  g0035(.din(G30), .dout(new_new_n763__));
  buf1  g0036(.din(G31), .dout(new_new_n765__));
  buf1  g0037(.din(G32), .dout(new_new_n767__));
  buf1  g0038(.din(G33), .dout(new_new_n769__));
  buf1  g0039(.din(G34), .dout(new_new_n771__));
  buf1  g0040(.din(G35), .dout(new_new_n773__));
  buf1  g0041(.din(G36), .dout(new_new_n775__));
  buf1  g0042(.din(G37), .dout(new_new_n777__));
  buf1  g0043(.din(G38), .dout(new_new_n779__));
  buf1  g0044(.din(G39), .dout(new_new_n781__));
  not1  g0045(.din(G40), .dout(new_new_n784__));
  buf1  g0046(.din(G41), .dout(new_new_n785__));
  buf1  g0047(.din(G42), .dout(new_new_n787__));
  buf1  g0048(.din(G43), .dout(new_new_n789__));
  buf1  g0049(.din(G44), .dout(new_new_n791__));
  buf1  g0050(.din(G45), .dout(new_new_n793__));
  buf1  g0051(.din(G46), .dout(new_new_n795__));
  buf1  g0052(.din(G47), .dout(new_new_n797__));
  buf1  g0053(.din(G48), .dout(new_new_n799__));
  buf1  g0054(.din(G49), .dout(new_new_n801__));
  buf1  g0055(.din(G50), .dout(new_new_n803__));
  buf1  g0056(.din(G51), .dout(new_new_n805__));
  buf1  g0057(.din(G52), .dout(new_new_n807__));
  buf1  g0058(.din(G53), .dout(new_new_n809__));
  buf1  g0059(.din(G54), .dout(new_new_n811__));
  buf1  g0060(.din(G55), .dout(new_new_n813__));
  buf1  g0061(.din(G56), .dout(new_new_n815__));
  buf1  g0062(.din(G57), .dout(new_new_n817__));
  buf1  g0063(.din(G58), .dout(new_new_n819__));
  buf1  g0064(.din(G59), .dout(new_new_n821__));
  buf1  g0065(.din(G60), .dout(new_new_n823__));
  not1  g0066(.din(n492_lo), .dout(new_new_n826__));
  buf1  g0067(.din(n495_lo), .dout(new_new_n827__));
  buf1  g0068(.din(n498_lo), .dout(new_new_n829__));
  not1  g0069(.din(n501_lo), .dout(new_new_n832__));
  not1  g0070(.din(n516_lo), .dout(new_new_n834__));
  not1  g0071(.din(n528_lo), .dout(new_new_n836__));
  buf1  g0072(.din(n540_lo), .dout(new_new_n837__));
  not1  g0073(.din(n540_lo), .dout(new_new_n838__));
  buf1  g0074(.din(n543_lo), .dout(new_new_n839__));
  buf1  g0075(.din(n546_lo), .dout(new_new_n841__));
  buf1  g0076(.din(n549_lo), .dout(new_new_n843__));
  buf1  g0077(.din(n552_lo), .dout(new_new_n845__));
  not1  g0078(.din(n552_lo), .dout(new_new_n846__));
  buf1  g0079(.din(n564_lo), .dout(new_new_n847__));
  not1  g0080(.din(n564_lo), .dout(new_new_n848__));
  not1  g0081(.din(n600_lo), .dout(new_new_n850__));
  buf1  g0082(.din(n603_lo), .dout(new_new_n851__));
  buf1  g0083(.din(n606_lo), .dout(new_new_n853__));
  not1  g0084(.din(n609_lo), .dout(new_new_n856__));
  buf1  g0085(.din(n615_lo), .dout(new_new_n857__));
  buf1  g0086(.din(n618_lo), .dout(new_new_n859__));
  not1  g0087(.din(n621_lo), .dout(new_new_n862__));
  buf1  g0088(.din(n627_lo), .dout(new_new_n863__));
  buf1  g0089(.din(n630_lo), .dout(new_new_n865__));
  not1  g0090(.din(n633_lo), .dout(new_new_n868__));
  buf1  g0091(.din(n639_lo), .dout(new_new_n869__));
  buf1  g0092(.din(n642_lo), .dout(new_new_n871__));
  buf1  g0093(.din(n645_lo), .dout(new_new_n873__));
  not1  g0094(.din(n648_lo), .dout(new_new_n876__));
  not1  g0095(.din(n660_lo), .dout(new_new_n878__));
  not1  g0096(.din(n672_lo), .dout(new_new_n880__));
  buf1  g0097(.din(n675_lo), .dout(new_new_n881__));
  buf1  g0098(.din(n678_lo), .dout(new_new_n883__));
  buf1  g0099(.din(n681_lo), .dout(new_new_n885__));
  not1  g0100(.din(n684_lo), .dout(new_new_n888__));
  buf1  g0101(.din(n687_lo), .dout(new_new_n889__));
  buf1  g0102(.din(n690_lo), .dout(new_new_n891__));
  buf1  g0103(.din(n693_lo), .dout(new_new_n893__));
  not1  g0104(.din(n696_lo), .dout(new_new_n896__));
  buf1  g0105(.din(n699_lo), .dout(new_new_n897__));
  buf1  g0106(.din(n702_lo), .dout(new_new_n899__));
  buf1  g0107(.din(n705_lo), .dout(new_new_n901__));
  buf1  g0108(.din(n708_lo), .dout(new_new_n903__));
  buf1  g0109(.din(n711_lo), .dout(new_new_n905__));
  buf1  g0110(.din(n714_lo), .dout(new_new_n907__));
  buf1  g0111(.din(n717_lo), .dout(new_new_n909__));
  buf1  g0112(.din(n720_lo), .dout(new_new_n911__));
  buf1  g0113(.din(n723_lo), .dout(new_new_n913__));
  buf1  g0114(.din(n726_lo), .dout(new_new_n915__));
  buf1  g0115(.din(n729_lo), .dout(new_new_n917__));
  buf1  g0116(.din(n732_lo), .dout(new_new_n919__));
  buf1  g0117(.din(n735_lo), .dout(new_new_n921__));
  buf1  g0118(.din(n738_lo), .dout(new_new_n923__));
  buf1  g0119(.din(n741_lo), .dout(new_new_n925__));
  buf1  g0120(.din(n744_lo), .dout(new_new_n927__));
  buf1  g0121(.din(n747_lo), .dout(new_new_n929__));
  buf1  g0122(.din(n750_lo), .dout(new_new_n931__));
  buf1  g0123(.din(n753_lo), .dout(new_new_n933__));
  not1  g0124(.din(n753_lo), .dout(new_new_n934__));
  not1  g0125(.din(n756_lo), .dout(new_new_n936__));
  buf1  g0126(.din(n759_lo), .dout(new_new_n937__));
  buf1  g0127(.din(n762_lo), .dout(new_new_n939__));
  buf1  g0128(.din(n765_lo), .dout(new_new_n941__));
  not1  g0129(.din(n765_lo), .dout(new_new_n942__));
  not1  g0130(.din(n768_lo), .dout(new_new_n944__));
  buf1  g0131(.din(n771_lo), .dout(new_new_n945__));
  buf1  g0132(.din(n774_lo), .dout(new_new_n947__));
  buf1  g0133(.din(n777_lo), .dout(new_new_n949__));
  not1  g0134(.din(n777_lo), .dout(new_new_n950__));
  not1  g0135(.din(n780_lo), .dout(new_new_n952__));
  buf1  g0136(.din(n783_lo), .dout(new_new_n953__));
  buf1  g0137(.din(n786_lo), .dout(new_new_n955__));
  not1  g0138(.din(n792_lo), .dout(new_new_n958__));
  buf1  g0139(.din(n795_lo), .dout(new_new_n959__));
  buf1  g0140(.din(n798_lo), .dout(new_new_n961__));
  buf1  g0141(.din(n807_lo), .dout(new_new_n963__));
  not1  g0142(.din(n816_lo), .dout(new_new_n966__));
  buf1  g0143(.din(n819_lo), .dout(new_new_n967__));
  not1  g0144(.din(n828_lo), .dout(new_new_n970__));
  buf1  g0145(.din(n831_lo), .dout(new_new_n971__));
  buf1  g0146(.din(n843_lo), .dout(new_new_n973__));
  buf1  g0147(.din(n846_lo), .dout(new_new_n975__));
  buf1  g0148(.din(n849_lo), .dout(new_new_n977__));
  buf1  g0149(.din(n852_lo), .dout(new_new_n979__));
  not1  g0150(.din(n852_lo), .dout(new_new_n980__));
  buf1  g0151(.din(n855_lo), .dout(new_new_n981__));
  buf1  g0152(.din(n858_lo), .dout(new_new_n983__));
  buf1  g0153(.din(n861_lo), .dout(new_new_n985__));
  buf1  g0154(.din(n864_lo), .dout(new_new_n987__));
  not1  g0155(.din(n864_lo), .dout(new_new_n988__));
  buf1  g0156(.din(n867_lo), .dout(new_new_n989__));
  buf1  g0157(.din(n870_lo), .dout(new_new_n991__));
  not1  g0158(.din(n870_lo), .dout(new_new_n992__));
  buf1  g0159(.din(n879_lo), .dout(new_new_n993__));
  buf1  g0160(.din(n882_lo), .dout(new_new_n995__));
  buf1  g0161(.din(n891_lo), .dout(new_new_n997__));
  buf1  g0162(.din(n903_lo), .dout(new_new_n999__));
  buf1  g0163(.din(n915_lo), .dout(new_new_n1001__));
  not1  g0164(.din(n918_lo), .dout(new_new_n1004__));
  buf1  g0165(.din(n951_lo), .dout(new_new_n1005__));
  buf1  g0166(.din(n954_lo), .dout(new_new_n1007__));
  buf1  g0167(.din(n957_lo), .dout(new_new_n1009__));
  not1  g0168(.din(n957_lo), .dout(new_new_n1010__));
  buf1  g0169(.din(n960_lo), .dout(new_new_n1011__));
  not1  g0170(.din(n960_lo), .dout(new_new_n1012__));
  buf1  g0171(.din(n963_lo), .dout(new_new_n1013__));
  buf1  g0172(.din(n966_lo), .dout(new_new_n1015__));
  buf1  g0173(.din(n969_lo), .dout(new_new_n1017__));
  not1  g0174(.din(n969_lo), .dout(new_new_n1018__));
  buf1  g0175(.din(n972_lo), .dout(new_new_n1019__));
  not1  g0176(.din(n972_lo), .dout(new_new_n1020__));
  buf1  g0177(.din(n975_lo), .dout(new_new_n1021__));
  buf1  g0178(.din(n978_lo), .dout(new_new_n1023__));
  buf1  g0179(.din(n981_lo), .dout(new_new_n1025__));
  not1  g0180(.din(n981_lo), .dout(new_new_n1026__));
  not1  g0181(.din(n984_lo), .dout(new_new_n1028__));
  buf1  g0182(.din(n987_lo), .dout(new_new_n1029__));
  buf1  g0183(.din(n990_lo), .dout(new_new_n1031__));
  buf1  g0184(.din(n993_lo), .dout(new_new_n1033__));
  not1  g0185(.din(n993_lo), .dout(new_new_n1034__));
  not1  g0186(.din(n996_lo), .dout(new_new_n1036__));
  buf1  g0187(.din(n999_lo), .dout(new_new_n1037__));
  buf1  g0188(.din(n1002_lo), .dout(new_new_n1039__));
  not1  g0189(.din(n1008_lo), .dout(new_new_n1042__));
  buf1  g0190(.din(n1011_lo), .dout(new_new_n1043__));
  buf1  g0191(.din(n1014_lo), .dout(new_new_n1045__));
  not1  g0192(.din(n1014_lo), .dout(new_new_n1046__));
  not1  g0193(.din(n1020_lo), .dout(new_new_n1048__));
  buf1  g0194(.din(n1023_lo), .dout(new_new_n1049__));
  not1  g0195(.din(n1032_lo), .dout(new_new_n1052__));
  buf1  g0196(.din(n1035_lo), .dout(new_new_n1053__));
  not1  g0197(.din(n1044_lo), .dout(new_new_n1056__));
  buf1  g0198(.din(n1047_lo), .dout(new_new_n1057__));
  buf1  g0199(.din(n1050_lo), .dout(new_new_n1059__));
  buf1  g0200(.din(n1053_lo), .dout(new_new_n1061__));
  buf1  g0201(.din(n1056_lo), .dout(new_new_n1063__));
  not1  g0202(.din(n1056_lo), .dout(new_new_n1064__));
  buf1  g0203(.din(n1059_lo), .dout(new_new_n1065__));
  buf1  g0204(.din(n1062_lo), .dout(new_new_n1067__));
  buf1  g0205(.din(n1065_lo), .dout(new_new_n1069__));
  not1  g0206(.din(n1068_lo), .dout(new_new_n1072__));
  buf1  g0207(.din(n1071_lo), .dout(new_new_n1073__));
  buf1  g0208(.din(n1074_lo), .dout(new_new_n1075__));
  buf1  g0209(.din(n1077_lo), .dout(new_new_n1077__));
  not1  g0210(.din(n1080_lo), .dout(new_new_n1080__));
  buf1  g0211(.din(n1083_lo), .dout(new_new_n1081__));
  buf1  g0212(.din(n1086_lo), .dout(new_new_n1083__));
  buf1  g0213(.din(n1089_lo), .dout(new_new_n1085__));
  not1  g0214(.din(n1092_lo), .dout(new_new_n1088__));
  buf1  g0215(.din(n1095_lo), .dout(new_new_n1089__));
  buf1  g0216(.din(n1098_lo), .dout(new_new_n1091__));
  buf1  g0217(.din(n1101_lo), .dout(new_new_n1093__));
  not1  g0218(.din(n1104_lo), .dout(new_new_n1096__));
  buf1  g0219(.din(n1107_lo), .dout(new_new_n1097__));
  buf1  g0220(.din(n1110_lo), .dout(new_new_n1099__));
  buf1  g0221(.din(n1113_lo), .dout(new_new_n1101__));
  not1  g0222(.din(n1116_lo), .dout(new_new_n1104__));
  buf1  g0223(.din(n1119_lo), .dout(new_new_n1105__));
  buf1  g0224(.din(n1122_lo), .dout(new_new_n1107__));
  buf1  g0225(.din(n1125_lo), .dout(new_new_n1109__));
  not1  g0226(.din(n1128_lo), .dout(new_new_n1112__));
  buf1  g0227(.din(n1131_lo), .dout(new_new_n1113__));
  buf1  g0228(.din(n1134_lo), .dout(new_new_n1115__));
  buf1  g0229(.din(n1137_lo), .dout(new_new_n1117__));
  buf1  g0230(.din(n1143_lo), .dout(new_new_n1119__));
  buf1  g0231(.din(n1146_lo), .dout(new_new_n1121__));
  buf1  g0232(.din(n1149_lo), .dout(new_new_n1123__));
  not1  g0233(.din(n1152_lo), .dout(new_new_n1126__));
  buf1  g0234(.din(n1155_lo), .dout(new_new_n1127__));
  not1  g0235(.din(n1164_lo), .dout(new_new_n1130__));
  buf1  g0236(.din(n1167_lo), .dout(new_new_n1131__));
  buf1  g0237(.din(n1170_lo), .dout(new_new_n1133__));
  buf1  g0238(.din(n1173_lo), .dout(new_new_n1135__));
  not1  g0239(.din(n1176_lo), .dout(new_new_n1138__));
  not1  g0240(.din(n1188_lo), .dout(new_new_n1140__));
  not1  g0241(.din(n563_inv), .dout(new_new_n1142__));
  not1  g0242(.din(n1429_o2), .dout(new_new_n1144__));
  buf1  g0243(.din(n1427_o2), .dout(new_new_n1145__));
  not1  g0244(.din(n1471_o2), .dout(new_new_n1148__));
  not1  g0245(.din(n1476_o2), .dout(new_new_n1150__));
  buf1  g0246(.din(n1499_o2), .dout(new_new_n1151__));
  not1  g0247(.din(n1499_o2), .dout(new_new_n1152__));
  buf1  g0248(.din(n1500_o2), .dout(new_new_n1153__));
  not1  g0249(.din(n1501_o2), .dout(new_new_n1156__));
  not1  g0250(.din(n1516_o2), .dout(new_new_n1158__));
  not1  g0251(.din(n1517_o2), .dout(new_new_n1160__));
  buf1  g0252(.din(n1562_o2), .dout(new_new_n1161__));
  not1  g0253(.din(n1562_o2), .dout(new_new_n1162__));
  not1  g0254(.din(n1563_o2), .dout(new_new_n1164__));
  buf1  g0255(.din(n1564_o2), .dout(new_new_n1165__));
  buf1  g0256(.din(n1582_o2), .dout(new_new_n1167__));
  not1  g0257(.din(n1582_o2), .dout(new_new_n1168__));
  buf1  g0258(.din(n1583_o2), .dout(new_new_n1169__));
  not1  g0259(.din(n1583_o2), .dout(new_new_n1170__));
  buf1  g0260(.din(n1618_o2), .dout(new_new_n1171__));
  not1  g0261(.din(n1618_o2), .dout(new_new_n1172__));
  not1  g0262(.din(n1622_o2), .dout(new_new_n1174__));
  not1  g0263(.din(n1502_o2), .dout(new_new_n1176__));
  buf1  g0264(.din(n1503_o2), .dout(new_new_n1177__));
  buf1  g0265(.din(n1504_o2), .dout(new_new_n1179__));
  buf1  g0266(.din(n1505_o2), .dout(new_new_n1181__));
  buf1  g0267(.din(n1506_o2), .dout(new_new_n1183__));
  buf1  g0268(.din(n1512_o2), .dout(new_new_n1185__));
  not1  g0269(.din(n1512_o2), .dout(new_new_n1186__));
  buf1  g0270(.din(n1513_o2), .dout(new_new_n1187__));
  buf1  g0271(.din(n1514_o2), .dout(new_new_n1189__));
  buf1  g0272(.din(n1515_o2), .dout(new_new_n1191__));
  not1  g0273(.din(n1644_o2), .dout(new_new_n1194__));
  not1  g0274(.din(n1647_o2), .dout(new_new_n1196__));
  buf1  g0275(.din(n1527_o2), .dout(new_new_n1197__));
  buf1  g0276(.din(n650_inv), .dout(new_new_n1199__));
  not1  g0277(.din(n650_inv), .dout(new_new_n1200__));
  buf1  g0278(.din(n653_inv), .dout(new_new_n1201__));
  buf1  g0279(.din(n656_inv), .dout(new_new_n1203__));
  not1  g0280(.din(n1567_o2), .dout(new_new_n1206__));
  buf1  g0281(.din(n955_o2), .dout(new_new_n1207__));
  not1  g0282(.din(n955_o2), .dout(new_new_n1208__));
  buf1  g0283(.din(n1568_o2), .dout(new_new_n1209__));
  not1  g0284(.din(n1037_o2), .dout(new_new_n1212__));
  buf1  g0285(.din(n960_o2), .dout(new_new_n1213__));
  buf1  g0286(.din(n1587_o2), .dout(new_new_n1215__));
  not1  g0287(.din(n1587_o2), .dout(new_new_n1216__));
  buf1  g0288(.din(n1040_o2), .dout(new_new_n1217__));
  not1  g0289(.din(n1040_o2), .dout(new_new_n1218__));
  buf1  g0290(.din(n1039_o2), .dout(new_new_n1219__));
  not1  g0291(.din(n1039_o2), .dout(new_new_n1220__));
  buf1  g0292(.din(n1589_o2), .dout(new_new_n1221__));
  not1  g0293(.din(n1589_o2), .dout(new_new_n1222__));
  not1  g0294(.din(n1624_o2), .dout(new_new_n1224__));
  buf1  g0295(.din(n1643_o2), .dout(new_new_n1225__));
  not1  g0296(.din(n1643_o2), .dout(new_new_n1226__));
  buf1  g0297(.din(n1038_o2), .dout(new_new_n1227__));
  not1  g0298(.din(n1038_o2), .dout(new_new_n1228__));
  buf1  g0299(.din(n1645_o2), .dout(new_new_n1229__));
  not1  g0300(.din(n1645_o2), .dout(new_new_n1230__));
  not1  g0301(.din(n1029_o2), .dout(new_new_n1232__));
  buf1  g0302(.din(n701_inv), .dout(new_new_n1233__));
  buf1  g0303(.din(n1662_o2), .dout(new_new_n1235__));
  buf1  g0304(.din(n1663_o2), .dout(new_new_n1237__));
  buf1  g0305(.din(n710_inv), .dout(new_new_n1239__));
  not1  g0306(.din(n813_o2), .dout(new_new_n1242__));
  buf1  g0307(.din(lo114_buf_o2), .dout(new_new_n1243__));
  not1  g0308(.din(lo114_buf_o2), .dout(new_new_n1244__));
  buf1  g0309(.din(n1031_o2), .dout(new_new_n1245__));
  not1  g0310(.din(n1031_o2), .dout(new_new_n1246__));
  buf1  g0311(.din(lo186_buf_o2), .dout(new_new_n1247__));
  not1  g0312(.din(lo186_buf_o2), .dout(new_new_n1248__));
  buf1  g0313(.din(n1042_o2), .dout(new_new_n1249__));
  not1  g0314(.din(n1042_o2), .dout(new_new_n1250__));
  buf1  g0315(.din(n728_inv), .dout(new_new_n1251__));
  buf1  g0316(.din(n917_o2), .dout(new_new_n1253__));
  buf1  g0317(.din(n734_inv), .dout(new_new_n1255__));
  buf1  g0318(.din(n1649_o2), .dout(new_new_n1257__));
  buf1  g0319(.din(n1650_o2), .dout(new_new_n1259__));
  not1  g0320(.din(n1650_o2), .dout(new_new_n1260__));
  buf1  g0321(.din(n1651_o2), .dout(new_new_n1261__));
  buf1  g0322(.din(n1652_o2), .dout(new_new_n1263__));
  buf1  g0323(.din(n1653_o2), .dout(new_new_n1265__));
  buf1  g0324(.din(lo138_buf_o2), .dout(new_new_n1267__));
  buf1  g0325(.din(n1664_o2), .dout(new_new_n1269__));
  buf1  g0326(.din(n1665_o2), .dout(new_new_n1271__));
  buf1  g0327(.din(n1666_o2), .dout(new_new_n1273__));
  buf1  g0328(.din(n1667_o2), .dout(new_new_n1275__));
  buf1  g0329(.din(n944_o2), .dout(new_new_n1277__));
  buf1  g0330(.din(n770_inv), .dout(new_new_n1279__));
  buf1  g0331(.din(n1672_o2), .dout(new_new_n1281__));
  buf1  g0332(.din(n776_inv), .dout(new_new_n1283__));
  buf1  g0333(.din(n1679_o2), .dout(new_new_n1285__));
  buf1  g0334(.din(n782_inv), .dout(new_new_n1287__));
  not1  g0335(.din(n782_inv), .dout(new_new_n1288__));
  buf1  g0336(.din(n785_inv), .dout(new_new_n1289__));
  buf1  g0337(.din(lo110_buf_o2), .dout(new_new_n1291__));
  not1  g0338(.din(lo110_buf_o2), .dout(new_new_n1292__));
  buf1  g0339(.din(lo134_buf_o2), .dout(new_new_n1293__));
  buf1  g0340(.din(n1030_o2), .dout(new_new_n1295__));
  not1  g0341(.din(n1030_o2), .dout(new_new_n1296__));
  buf1  g0342(.din(lo182_buf_o2), .dout(new_new_n1297__));
  not1  g0343(.din(lo182_buf_o2), .dout(new_new_n1298__));
  not1  g0344(.din(n830_o2), .dout(new_new_n1300__));
  buf1  g0345(.din(n1021_o2), .dout(new_new_n1301__));
  not1  g0346(.din(n1021_o2), .dout(new_new_n1302__));
  buf1  g0347(.din(n806_inv), .dout(new_new_n1303__));
  buf1  g0348(.din(n809_inv), .dout(new_new_n1305__));
  buf1  g0349(.din(n946_o2), .dout(new_new_n1307__));
  buf1  g0350(.din(lo038_buf_o2), .dout(new_new_n1309__));
  not1  g0351(.din(lo038_buf_o2), .dout(new_new_n1310__));
  buf1  g0352(.din(lo238_buf_o2), .dout(new_new_n1311__));
  buf1  g0353(.din(n1010_o2), .dout(new_new_n1313__));
  not1  g0354(.din(n1010_o2), .dout(new_new_n1314__));
  buf1  g0355(.din(n1006_o2), .dout(new_new_n1315__));
  not1  g0356(.din(n1006_o2), .dout(new_new_n1316__));
  buf1  g0357(.din(n907_o2), .dout(new_new_n1317__));
  not1  g0358(.din(n907_o2), .dout(new_new_n1318__));
  not1  g0359(.din(n902_o2), .dout(new_new_n1320__));
  not1  g0360(.din(lo154_buf_o2), .dout(new_new_n1322__));
  buf1  g0361(.din(n836_inv), .dout(new_new_n1323__));
  buf1  g0362(.din(n839_inv), .dout(new_new_n1325__));
  buf1  g0363(.din(lo122_buf_o2), .dout(new_new_n1327__));
  buf1  g0364(.din(n845_inv), .dout(new_new_n1329__));
  not1  g0365(.din(n845_inv), .dout(new_new_n1330__));
  buf1  g0366(.din(n904_o2), .dout(new_new_n1331__));
  not1  g0367(.din(n904_o2), .dout(new_new_n1332__));
  buf1  g0368(.din(lo106_buf_o2), .dout(new_new_n1333__));
  not1  g0369(.din(lo106_buf_o2), .dout(new_new_n1334__));
  not1  g0370(.din(n980_o2), .dout(new_new_n1336__));
  buf1  g0371(.din(n1023_o2), .dout(new_new_n1337__));
  not1  g0372(.din(n1023_o2), .dout(new_new_n1338__));
  buf1  g0373(.din(lo178_buf_o2), .dout(new_new_n1339__));
  not1  g0374(.din(lo178_buf_o2), .dout(new_new_n1340__));
  not1  g0375(.din(n981_o2), .dout(new_new_n1342__));
  buf1  g0376(.din(n837_o2), .dout(new_new_n1343__));
  not1  g0377(.din(n837_o2), .dout(new_new_n1344__));
  buf1  g0378(.din(n1013_o2), .dout(new_new_n1345__));
  not1  g0379(.din(n1013_o2), .dout(new_new_n1346__));
  buf1  g0380(.din(n840_o2), .dout(new_new_n1347__));
  not1  g0381(.din(n840_o2), .dout(new_new_n1348__));
  buf1  g0382(.din(n849_o2), .dout(new_new_n1349__));
  not1  g0383(.din(n849_o2), .dout(new_new_n1350__));
  buf1  g0384(.din(n852_o2), .dout(new_new_n1351__));
  not1  g0385(.din(n852_o2), .dout(new_new_n1352__));
  buf1  g0386(.din(n864_o2), .dout(new_new_n1353__));
  not1  g0387(.din(n864_o2), .dout(new_new_n1354__));
  buf1  g0388(.din(n867_o2), .dout(new_new_n1355__));
  not1  g0389(.din(n867_o2), .dout(new_new_n1356__));
  buf1  g0390(.din(n1044_o2), .dout(new_new_n1357__));
  not1  g0391(.din(n1044_o2), .dout(new_new_n1358__));
  buf1  g0392(.din(n876_o2), .dout(new_new_n1359__));
  not1  g0393(.din(n876_o2), .dout(new_new_n1360__));
  buf1  g0394(.din(n893_inv), .dout(new_new_n1361__));
  buf1  g0395(.din(n879_o2), .dout(new_new_n1363__));
  not1  g0396(.din(n879_o2), .dout(new_new_n1364__));
  not1  g0397(.din(n925_o2), .dout(new_new_n1366__));
  buf1  g0398(.din(n902_inv), .dout(new_new_n1367__));
  not1  g0399(.din(n902_inv), .dout(new_new_n1368__));
  buf1  g0400(.din(lo146_buf_o2), .dout(new_new_n1369__));
  not1  g0401(.din(n1026_o2), .dout(new_new_n1372__));
  not1  g0402(.din(n1032_o2), .dout(new_new_n1374__));
  buf1  g0403(.din(lo118_buf_o2), .dout(new_new_n1375__));
  buf1  g0404(.din(n917_inv), .dout(new_new_n1377__));
  not1  g0405(.din(n917_inv), .dout(new_new_n1378__));
  buf1  g0406(.din(lo190_buf_o2), .dout(new_new_n1379__));
  not1  g0407(.din(lo190_buf_o2), .dout(new_new_n1380__));
  not1  g0408(.din(n1036_o2), .dout(new_new_n1382__));
  buf1  g0409(.din(n926_inv), .dout(new_new_n1383__));
  not1  g0410(.din(n926_inv), .dout(new_new_n1384__));
  buf1  g0411(.din(n929_inv), .dout(new_new_n1385__));
  not1  g0412(.din(n929_inv), .dout(new_new_n1386__));
  buf1  g0413(.din(lo002_buf_o2), .dout(new_new_n1387__));
  not1  g0414(.din(lo002_buf_o2), .dout(new_new_n1388__));
  buf1  g0415(.din(lo014_buf_o2), .dout(new_new_n1389__));
  buf1  g0416(.din(lo030_buf_o2), .dout(new_new_n1391__));
  buf1  g0417(.din(lo034_buf_o2), .dout(new_new_n1393__));
  buf1  g0418(.din(lo042_buf_o2), .dout(new_new_n1395__));
  buf1  g0419(.din(lo113_buf_o2), .dout(new_new_n1397__));
  not1  g0420(.din(lo113_buf_o2), .dout(new_new_n1398__));
  buf1  g0421(.din(lo185_buf_o2), .dout(new_new_n1399__));
  not1  g0422(.din(lo185_buf_o2), .dout(new_new_n1400__));
  not1  g0423(.din(n939_o2), .dout(new_new_n1402__));
  not1  g0424(.din(n941_o2), .dout(new_new_n1404__));
  buf1  g0425(.din(lo142_buf_o2), .dout(new_new_n1405__));
  not1  g0426(.din(lo142_buf_o2), .dout(new_new_n1406__));
  buf1  g0427(.din(lo230_buf_o2), .dout(new_new_n1407__));
  not1  g0428(.din(lo230_buf_o2), .dout(new_new_n1408__));
  buf1  g0429(.din(lo006_buf_o2), .dout(new_new_n1409__));
  buf1  g0430(.din(lo018_buf_o2), .dout(new_new_n1411__));
  buf1  g0431(.din(lo022_buf_o2), .dout(new_new_n1413__));
  buf1  g0432(.din(lo066_buf_o2), .dout(new_new_n1415__));
  buf1  g0433(.din(n977_inv), .dout(new_new_n1417__));
  not1  g0434(.din(n977_inv), .dout(new_new_n1418__));
  buf1  g0435(.din(n826_o2), .dout(new_new_n1419__));
  buf1  g0436(.din(n892_o2), .dout(new_new_n1421__));
  buf1  g0437(.din(lo152_buf_o2), .dout(new_new_n1423__));
  buf1  g0438(.din(n896_o2), .dout(new_new_n1425__));
  buf1  g0439(.din(n905_o2), .dout(new_new_n1427__));
  buf1  g0440(.din(n995_inv), .dout(new_new_n1429__));
  not1  g0441(.din(n995_inv), .dout(new_new_n1430__));
  buf1  g0442(.din(lo037_buf_o2), .dout(new_new_n1431__));
  buf1  g0443(.din(lo237_buf_o2), .dout(new_new_n1433__));
  not1  g0444(.din(lo237_buf_o2), .dout(new_new_n1434__));
  buf1  g0445(.din(lo062_buf_o2), .dout(new_new_n1435__));
  not1  g0446(.din(lo062_buf_o2), .dout(new_new_n1436__));
  buf1  g0447(.din(n1007_inv), .dout(new_new_n1437__));
  buf1  g0448(.din(n1010_inv), .dout(new_new_n1439__));
  buf1  g0449(.din(n891_o2), .dout(new_new_n1441__));
  and1  g0450(.dina(new_new_n847__), .dinb(new_new_n837__), .dout(new_new_n1443__));
  or1   g0451(.dina(new_new_n848__), .dinb(new_new_n2116__), .dout(new_new_n1444__));
  or1   g0452(.dina(new_new_n2117__), .dinb(new_new_n2118__), .dout(new_new_n1445__));
  or1   g0453(.dina(new_new_n1144__), .dinb(new_new_n2120__), .dout(new_new_n1446__));
  and1  g0454(.dina(new_new_n1443__), .dinb(new_new_n2121__), .dout(new_new_n1447__));
  or1   g0455(.dina(new_new_n2117__), .dinb(new_new_n2120__), .dout(new_new_n1448__));
  or1   g0456(.dina(new_new_n896__), .dinb(new_new_n888__), .dout(new_new_n1449__));
  or1   g0457(.dina(new_new_n1242__), .dinb(new_new_n834__), .dout(new_new_n1450__));
  or1   g0458(.dina(new_new_n2122__), .dinb(new_new_n826__), .dout(new_new_n1451__));
  or1   g0459(.dina(new_new_n2122__), .dinb(new_new_n836__), .dout(new_new_n1452__));
  or1   g0460(.dina(new_new_n2123__), .dinb(new_new_n1447__), .dout(new_new_n1453__));
  or1   g0461(.dina(new_new_n880__), .dinb(new_new_n2124__), .dout(new_new_n1454__));
  or1   g0462(.dina(new_new_n2125__), .dinb(new_new_n2118__), .dout(new_new_n1455__));
  or1   g0463(.dina(new_new_n2125__), .dinb(new_new_n2119__), .dout(new_new_n1456__));
  and1  g0464(.dina(new_new_n1145__), .dinb(new_new_n2121__), .dout(new_new_n1457__));
  or1   g0465(.dina(new_new_n911__), .dinb(new_new_n903__), .dout(new_new_n1458__));
  and1  g0466(.dina(new_new_n2126__), .dinb(new_new_n927__), .dout(new_new_n1459__));
  or1   g0467(.dina(new_new_n2123__), .dinb(new_new_n2127__), .dout(new_new_n1460__));
  or1   g0468(.dina(new_new_n2128__), .dinb(new_new_n2116__), .dout(new_new_n1461__));
  or1   g0469(.dina(new_new_n876__), .dinb(new_new_n2124__), .dout(new_new_n1462__));
  or1   g0470(.dina(new_new_n1462__), .dinb(new_new_n2128__), .dout(new_new_n1463__));
  and1  g0471(.dina(new_new_n2126__), .dinb(new_new_n919__), .dout(new_new_n1464__));
  and1  g0472(.dina(new_new_n2129__), .dinb(new_new_n2130__), .dout(new_new_n1465__));
  or1   g0473(.dina(new_new_n2131__), .dinb(new_new_n2132__), .dout(new_new_n1466__));
  and1  g0474(.dina(new_new_n2131__), .dinb(new_new_n2132__), .dout(new_new_n1467__));
  or1   g0475(.dina(new_new_n2129__), .dinb(new_new_n2130__), .dout(new_new_n1468__));
  and1  g0476(.dina(new_new_n1468__), .dinb(new_new_n1466__), .dout(new_new_n1469__));
  or1   g0477(.dina(new_new_n1467__), .dinb(new_new_n1465__), .dout(new_new_n1470__));
  and1  g0478(.dina(new_new_n2133__), .dinb(new_new_n2135__), .dout(new_new_n1471__));
  or1   g0479(.dina(new_new_n2137__), .dinb(new_new_n2139__), .dout(new_new_n1472__));
  and1  g0480(.dina(new_new_n2137__), .dinb(new_new_n2139__), .dout(new_new_n1473__));
  or1   g0481(.dina(new_new_n2133__), .dinb(new_new_n2135__), .dout(new_new_n1474__));
  and1  g0482(.dina(new_new_n1474__), .dinb(new_new_n1472__), .dout(new_new_n1475__));
  or1   g0483(.dina(new_new_n1473__), .dinb(new_new_n1471__), .dout(new_new_n1476__));
  and1  g0484(.dina(new_new_n2141__), .dinb(new_new_n2142__), .dout(new_new_n1477__));
  or1   g0485(.dina(new_new_n2143__), .dinb(new_new_n2144__), .dout(new_new_n1478__));
  and1  g0486(.dina(new_new_n2143__), .dinb(new_new_n2144__), .dout(new_new_n1479__));
  or1   g0487(.dina(new_new_n2141__), .dinb(new_new_n2142__), .dout(new_new_n1480__));
  and1  g0488(.dina(new_new_n1480__), .dinb(new_new_n1478__), .dout(new_new_n1481__));
  or1   g0489(.dina(new_new_n1479__), .dinb(new_new_n1477__), .dout(new_new_n1482__));
  and1  g0490(.dina(new_new_n2145__), .dinb(new_new_n2146__), .dout(new_new_n1483__));
  or1   g0491(.dina(new_new_n2147__), .dinb(new_new_n2148__), .dout(new_new_n1484__));
  and1  g0492(.dina(new_new_n2147__), .dinb(new_new_n2148__), .dout(new_new_n1485__));
  or1   g0493(.dina(new_new_n2145__), .dinb(new_new_n2146__), .dout(new_new_n1486__));
  and1  g0494(.dina(new_new_n1486__), .dinb(new_new_n1484__), .dout(new_new_n1487__));
  or1   g0495(.dina(new_new_n1485__), .dinb(new_new_n1483__), .dout(new_new_n1488__));
  and1  g0496(.dina(new_new_n1488__), .dinb(new_new_n1476__), .dout(new_new_n1489__));
  and1  g0497(.dina(new_new_n1487__), .dinb(new_new_n1475__), .dout(new_new_n1490__));
  or1   g0498(.dina(new_new_n1490__), .dinb(new_new_n1489__), .dout(new_new_n1491__));
  and1  g0499(.dina(new_new_n2149__), .dinb(new_new_n2150__), .dout(new_new_n1492__));
  or1   g0500(.dina(new_new_n2151__), .dinb(new_new_n2152__), .dout(new_new_n1493__));
  and1  g0501(.dina(new_new_n2151__), .dinb(new_new_n2152__), .dout(new_new_n1494__));
  or1   g0502(.dina(new_new_n2149__), .dinb(new_new_n2150__), .dout(new_new_n1495__));
  and1  g0503(.dina(new_new_n1495__), .dinb(new_new_n1493__), .dout(new_new_n1496__));
  or1   g0504(.dina(new_new_n1494__), .dinb(new_new_n1492__), .dout(new_new_n1497__));
  and1  g0505(.dina(new_new_n2153__), .dinb(new_new_n2136__), .dout(new_new_n1498__));
  or1   g0506(.dina(new_new_n2154__), .dinb(new_new_n2140__), .dout(new_new_n1499__));
  and1  g0507(.dina(new_new_n2154__), .dinb(new_new_n2140__), .dout(new_new_n1500__));
  or1   g0508(.dina(new_new_n2153__), .dinb(new_new_n2136__), .dout(new_new_n1501__));
  and1  g0509(.dina(new_new_n1501__), .dinb(new_new_n1499__), .dout(new_new_n1502__));
  or1   g0510(.dina(new_new_n1500__), .dinb(new_new_n1498__), .dout(new_new_n1503__));
  and1  g0511(.dina(new_new_n2155__), .dinb(new_new_n2156__), .dout(new_new_n1504__));
  or1   g0512(.dina(new_new_n2157__), .dinb(new_new_n2158__), .dout(new_new_n1505__));
  and1  g0513(.dina(new_new_n2157__), .dinb(new_new_n2158__), .dout(new_new_n1506__));
  or1   g0514(.dina(new_new_n2155__), .dinb(new_new_n2156__), .dout(new_new_n1507__));
  and1  g0515(.dina(new_new_n1507__), .dinb(new_new_n1505__), .dout(new_new_n1508__));
  or1   g0516(.dina(new_new_n1506__), .dinb(new_new_n1504__), .dout(new_new_n1509__));
  and1  g0517(.dina(new_new_n2159__), .dinb(new_new_n2160__), .dout(new_new_n1510__));
  or1   g0518(.dina(new_new_n2161__), .dinb(new_new_n2162__), .dout(new_new_n1511__));
  and1  g0519(.dina(new_new_n2161__), .dinb(new_new_n2162__), .dout(new_new_n1512__));
  or1   g0520(.dina(new_new_n2159__), .dinb(new_new_n2160__), .dout(new_new_n1513__));
  and1  g0521(.dina(new_new_n1513__), .dinb(new_new_n1511__), .dout(new_new_n1514__));
  or1   g0522(.dina(new_new_n1512__), .dinb(new_new_n1510__), .dout(new_new_n1515__));
  and1  g0523(.dina(new_new_n1515__), .dinb(new_new_n1503__), .dout(new_new_n1516__));
  and1  g0524(.dina(new_new_n1514__), .dinb(new_new_n1502__), .dout(new_new_n1517__));
  or1   g0525(.dina(new_new_n1517__), .dinb(new_new_n1516__), .dout(new_new_n1518__));
  and1  g0526(.dina(new_new_n1151__), .dinb(new_new_n2165__), .dout(new_new_n1519__));
  or1   g0527(.dina(new_new_n1519__), .dinb(new_new_n1150__), .dout(new_new_n1520__));
  or1   g0528(.dina(new_new_n1130__), .dinb(new_new_n2173__), .dout(new_new_n1521__));
  and1  g0529(.dina(new_new_n1521__), .dinb(new_new_n1520__), .dout(new_new_n1522__));
  or1   g0530(.dina(new_new_n1153__), .dinb(new_new_n2173__), .dout(new_new_n1523__));
  and1  g0531(.dina(new_new_n1152__), .dinb(new_new_n2182__), .dout(new_new_n1524__));
  and1  g0532(.dina(new_new_n1524__), .dinb(new_new_n1523__), .dout(new_new_n1525__));
  or1   g0533(.dina(new_new_n1525__), .dinb(new_new_n1522__), .dout(new_new_n1526__));
  or1   g0534(.dina(new_new_n1148__), .dinb(new_new_n2189__), .dout(new_new_n1527__));
  or1   g0535(.dina(new_new_n2196__), .dinb(new_new_n1056__), .dout(new_new_n1528__));
  or1   g0536(.dina(new_new_n2203__), .dinb(new_new_n970__), .dout(new_new_n1529__));
  or1   g0537(.dina(new_new_n1138__), .dinb(new_new_n2207__), .dout(new_new_n1530__));
  and1  g0538(.dina(new_new_n1530__), .dinb(new_new_n1529__), .dout(new_new_n1531__));
  and1  g0539(.dina(new_new_n1531__), .dinb(new_new_n1528__), .dout(new_new_n1532__));
  and1  g0540(.dina(new_new_n1532__), .dinb(new_new_n1527__), .dout(new_new_n1533__));
  and1  g0541(.dina(new_new_n1533__), .dinb(new_new_n1526__), .dout(new_new_n1534__));
  or1   g0542(.dina(new_new_n1196__), .dinb(new_new_n2174__), .dout(new_new_n1535__));
  and1  g0543(.dina(new_new_n1207__), .dinb(new_new_n2165__), .dout(new_new_n1536__));
  or1   g0544(.dina(new_new_n1536__), .dinb(new_new_n1194__), .dout(new_new_n1537__));
  and1  g0545(.dina(new_new_n1537__), .dinb(new_new_n1535__), .dout(new_new_n1538__));
  or1   g0546(.dina(new_new_n1213__), .dinb(new_new_n2174__), .dout(new_new_n1539__));
  and1  g0547(.dina(new_new_n1208__), .dinb(new_new_n2182__), .dout(new_new_n1540__));
  and1  g0548(.dina(new_new_n1540__), .dinb(new_new_n1539__), .dout(new_new_n1541__));
  or1   g0549(.dina(new_new_n1541__), .dinb(new_new_n1538__), .dout(new_new_n1542__));
  or1   g0550(.dina(new_new_n1174__), .dinb(new_new_n2189__), .dout(new_new_n1543__));
  or1   g0551(.dina(new_new_n2203__), .dinb(new_new_n958__), .dout(new_new_n1544__));
  or1   g0552(.dina(new_new_n2196__), .dinb(new_new_n1042__), .dout(new_new_n1545__));
  and1  g0553(.dina(new_new_n1545__), .dinb(new_new_n1544__), .dout(new_new_n1546__));
  and1  g0554(.dina(new_new_n1546__), .dinb(new_new_n1543__), .dout(new_new_n1547__));
  and1  g0555(.dina(new_new_n1547__), .dinb(new_new_n1542__), .dout(new_new_n1548__));
  and1  g0556(.dina(new_new_n1171__), .dinb(new_new_n2208__), .dout(new_new_n1549__));
  or1   g0557(.dina(new_new_n1172__), .dinb(new_new_n1167__), .dout(new_new_n1550__));
  or1   g0558(.dina(new_new_n1549__), .dinb(new_new_n1170__), .dout(new_new_n1551__));
  or1   g0559(.dina(new_new_n2209__), .dinb(new_new_n1169__), .dout(new_new_n1552__));
  and1  g0560(.dina(new_new_n1552__), .dinb(new_new_n1551__), .dout(new_new_n1553__));
  or1   g0561(.dina(new_new_n1553__), .dinb(new_new_n2176__), .dout(new_new_n1554__));
  or1   g0562(.dina(new_new_n2209__), .dinb(new_new_n2183__), .dout(new_new_n1555__));
  or1   g0563(.dina(new_new_n2208__), .dinb(new_new_n2166__), .dout(new_new_n1556__));
  or1   g0564(.dina(new_new_n1164__), .dinb(new_new_n2190__), .dout(new_new_n1557__));
  or1   g0565(.dina(new_new_n2197__), .dinb(new_new_n1048__), .dout(new_new_n1558__));
  and1  g0566(.dina(new_new_n1342__), .dinb(new_new_n1336__), .dout(new_new_n1559__));
  and1  g0567(.dina(new_new_n1559__), .dinb(new_new_n1558__), .dout(new_new_n1560__));
  and1  g0568(.dina(new_new_n1560__), .dinb(new_new_n1557__), .dout(new_new_n1561__));
  and1  g0569(.dina(new_new_n1561__), .dinb(new_new_n1556__), .dout(new_new_n1562__));
  and1  g0570(.dina(new_new_n1562__), .dinb(new_new_n1555__), .dout(new_new_n1563__));
  and1  g0571(.dina(new_new_n1563__), .dinb(new_new_n1554__), .dout(new_new_n1564__));
  and1  g0572(.dina(new_new_n1161__), .dinb(new_new_n2166__), .dout(new_new_n1565__));
  or1   g0573(.dina(new_new_n1565__), .dinb(new_new_n1158__), .dout(new_new_n1566__));
  or1   g0574(.dina(new_new_n1160__), .dinb(new_new_n2176__), .dout(new_new_n1567__));
  and1  g0575(.dina(new_new_n1567__), .dinb(new_new_n1566__), .dout(new_new_n1568__));
  or1   g0576(.dina(new_new_n1165__), .dinb(new_new_n2175__), .dout(new_new_n1569__));
  and1  g0577(.dina(new_new_n1162__), .dinb(new_new_n2183__), .dout(new_new_n1570__));
  and1  g0578(.dina(new_new_n1570__), .dinb(new_new_n1569__), .dout(new_new_n1571__));
  or1   g0579(.dina(new_new_n1571__), .dinb(new_new_n1568__), .dout(new_new_n1572__));
  or1   g0580(.dina(new_new_n1156__), .dinb(new_new_n2190__), .dout(new_new_n1573__));
  or1   g0581(.dina(new_new_n2197__), .dinb(new_new_n1052__), .dout(new_new_n1574__));
  or1   g0582(.dina(new_new_n2204__), .dinb(new_new_n966__), .dout(new_new_n1575__));
  or1   g0583(.dina(new_new_n1126__), .dinb(new_new_n2207__), .dout(new_new_n1576__));
  and1  g0584(.dina(new_new_n1576__), .dinb(new_new_n1575__), .dout(new_new_n1577__));
  and1  g0585(.dina(new_new_n1577__), .dinb(new_new_n1574__), .dout(new_new_n1578__));
  and1  g0586(.dina(new_new_n1578__), .dinb(new_new_n1573__), .dout(new_new_n1579__));
  and1  g0587(.dina(new_new_n1579__), .dinb(new_new_n1572__), .dout(new_new_n1580__));
  and1  g0588(.dina(new_new_n2210__), .dinb(new_new_n2211__), .dout(new_new_n1581__));
  or1   g0589(.dina(new_new_n2213__), .dinb(new_new_n2215__), .dout(new_new_n1582__));
  and1  g0590(.dina(new_new_n2213__), .dinb(new_new_n2215__), .dout(new_new_n1583__));
  or1   g0591(.dina(new_new_n2210__), .dinb(new_new_n2211__), .dout(new_new_n1584__));
  and1  g0592(.dina(new_new_n2216__), .dinb(new_new_n2217__), .dout(new_new_n1585__));
  or1   g0593(.dina(new_new_n1301__), .dinb(new_new_n1019__), .dout(new_new_n1586__));
  and1  g0594(.dina(new_new_n2218__), .dinb(new_new_n2220__), .dout(new_new_n1587__));
  or1   g0595(.dina(new_new_n2221__), .dinb(new_new_n2222__), .dout(new_new_n1588__));
  and1  g0596(.dina(new_new_n1588__), .dinb(new_new_n2223__), .dout(new_new_n1589__));
  or1   g0597(.dina(new_new_n1587__), .dinb(new_new_n2224__), .dout(new_new_n1590__));
  or1   g0598(.dina(new_new_n2225__), .dinb(new_new_n2226__), .dout(new_new_n1591__));
  and1  g0599(.dina(new_new_n1591__), .dinb(new_new_n2228__), .dout(new_new_n1592__));
  and1  g0600(.dina(new_new_n2229__), .dinb(new_new_n1217__), .dout(new_new_n1593__));
  or1   g0601(.dina(new_new_n1227__), .dinb(new_new_n1218__), .dout(new_new_n1594__));
  or1   g0602(.dina(new_new_n1593__), .dinb(new_new_n1220__), .dout(new_new_n1595__));
  or1   g0603(.dina(new_new_n2230__), .dinb(new_new_n1219__), .dout(new_new_n1596__));
  and1  g0604(.dina(new_new_n1596__), .dinb(new_new_n1595__), .dout(new_new_n1597__));
  or1   g0605(.dina(new_new_n1597__), .dinb(new_new_n2178__), .dout(new_new_n1598__));
  or1   g0606(.dina(new_new_n2230__), .dinb(new_new_n2185__), .dout(new_new_n1599__));
  or1   g0607(.dina(new_new_n2229__), .dinb(new_new_n2168__), .dout(new_new_n1600__));
  or1   g0608(.dina(new_new_n1212__), .dinb(new_new_n2192__), .dout(new_new_n1601__));
  or1   g0609(.dina(new_new_n2199__), .dinb(new_new_n1036__), .dout(new_new_n1602__));
  or1   g0610(.dina(new_new_n2204__), .dinb(new_new_n952__), .dout(new_new_n1603__));
  and1  g0611(.dina(new_new_n1603__), .dinb(new_new_n1602__), .dout(new_new_n1604__));
  and1  g0612(.dina(new_new_n1604__), .dinb(new_new_n1601__), .dout(new_new_n1605__));
  and1  g0613(.dina(new_new_n1605__), .dinb(new_new_n1600__), .dout(new_new_n1606__));
  and1  g0614(.dina(new_new_n1606__), .dinb(new_new_n1599__), .dout(new_new_n1607__));
  and1  g0615(.dina(new_new_n1607__), .dinb(new_new_n1598__), .dout(new_new_n1608__));
  and1  g0616(.dina(new_new_n1584__), .dinb(new_new_n2228__), .dout(new_new_n1609__));
  or1   g0617(.dina(new_new_n2226__), .dinb(new_new_n1581__), .dout(new_new_n1610__));
  and1  g0618(.dina(new_new_n1609__), .dinb(new_new_n1589__), .dout(new_new_n1611__));
  and1  g0619(.dina(new_new_n2231__), .dinb(new_new_n2225__), .dout(new_new_n1612__));
  or1   g0620(.dina(new_new_n1612__), .dinb(new_new_n2178__), .dout(new_new_n1613__));
  or1   g0621(.dina(new_new_n1613__), .dinb(new_new_n1611__), .dout(new_new_n1614__));
  or1   g0622(.dina(new_new_n2231__), .dinb(new_new_n2185__), .dout(new_new_n1615__));
  or1   g0623(.dina(new_new_n2227__), .dinb(new_new_n2168__), .dout(new_new_n1616__));
  or1   g0624(.dina(new_new_n2212__), .dinb(new_new_n2192__), .dout(new_new_n1617__));
  or1   g0625(.dina(new_new_n1140__), .dinb(new_new_n2206__), .dout(new_new_n1618__));
  or1   g0626(.dina(new_new_n2199__), .dinb(new_new_n2214__), .dout(new_new_n1619__));
  and1  g0627(.dina(new_new_n1619__), .dinb(new_new_n1618__), .dout(new_new_n1620__));
  and1  g0628(.dina(new_new_n1620__), .dinb(new_new_n1617__), .dout(new_new_n1621__));
  and1  g0629(.dina(new_new_n1621__), .dinb(new_new_n1616__), .dout(new_new_n1622__));
  and1  g0630(.dina(new_new_n1622__), .dinb(new_new_n1615__), .dout(new_new_n1623__));
  and1  g0631(.dina(new_new_n1623__), .dinb(new_new_n1614__), .dout(new_new_n1624__));
  and1  g0632(.dina(new_new_n2223__), .dinb(new_new_n2220__), .dout(new_new_n1625__));
  or1   g0633(.dina(new_new_n2224__), .dinb(new_new_n2222__), .dout(new_new_n1626__));
  and1  g0634(.dina(new_new_n1625__), .dinb(new_new_n2221__), .dout(new_new_n1627__));
  and1  g0635(.dina(new_new_n2232__), .dinb(new_new_n2218__), .dout(new_new_n1628__));
  or1   g0636(.dina(new_new_n1628__), .dinb(new_new_n2179__), .dout(new_new_n1629__));
  or1   g0637(.dina(new_new_n1629__), .dinb(new_new_n1627__), .dout(new_new_n1630__));
  or1   g0638(.dina(new_new_n2232__), .dinb(new_new_n2186__), .dout(new_new_n1631__));
  or1   g0639(.dina(new_new_n2219__), .dinb(new_new_n2169__), .dout(new_new_n1632__));
  or1   g0640(.dina(new_new_n2216__), .dinb(new_new_n2193__), .dout(new_new_n1633__));
  or1   g0641(.dina(new_new_n2206__), .dinb(new_new_n936__), .dout(new_new_n1634__));
  or1   g0642(.dina(new_new_n2200__), .dinb(new_new_n2217__), .dout(new_new_n1635__));
  and1  g0643(.dina(new_new_n1635__), .dinb(new_new_n1634__), .dout(new_new_n1636__));
  and1  g0644(.dina(new_new_n1636__), .dinb(new_new_n1633__), .dout(new_new_n1637__));
  and1  g0645(.dina(new_new_n1637__), .dinb(new_new_n1632__), .dout(new_new_n1638__));
  and1  g0646(.dina(new_new_n1638__), .dinb(new_new_n1631__), .dout(new_new_n1639__));
  and1  g0647(.dina(new_new_n1639__), .dinb(new_new_n1630__), .dout(new_new_n1640__));
  and1  g0648(.dina(new_new_n2233__), .dinb(new_new_n1245__), .dout(new_new_n1641__));
  or1   g0649(.dina(new_new_n1295__), .dinb(new_new_n1246__), .dout(new_new_n1642__));
  and1  g0650(.dina(new_new_n2234__), .dinb(new_new_n1250__), .dout(new_new_n1643__));
  and1  g0651(.dina(new_new_n1641__), .dinb(new_new_n1249__), .dout(new_new_n1644__));
  or1   g0652(.dina(new_new_n1644__), .dinb(new_new_n2179__), .dout(new_new_n1645__));
  or1   g0653(.dina(new_new_n1645__), .dinb(new_new_n1643__), .dout(new_new_n1646__));
  or1   g0654(.dina(new_new_n2234__), .dinb(new_new_n2186__), .dout(new_new_n1647__));
  or1   g0655(.dina(new_new_n2233__), .dinb(new_new_n2169__), .dout(new_new_n1648__));
  or1   g0656(.dina(new_new_n1232__), .dinb(new_new_n2193__), .dout(new_new_n1649__));
  or1   g0657(.dina(new_new_n2205__), .dinb(new_new_n944__), .dout(new_new_n1650__));
  or1   g0658(.dina(new_new_n2200__), .dinb(new_new_n1028__), .dout(new_new_n1651__));
  and1  g0659(.dina(new_new_n1651__), .dinb(new_new_n1650__), .dout(new_new_n1652__));
  and1  g0660(.dina(new_new_n1652__), .dinb(new_new_n1649__), .dout(new_new_n1653__));
  and1  g0661(.dina(new_new_n1653__), .dinb(new_new_n1648__), .dout(new_new_n1654__));
  and1  g0662(.dina(new_new_n1654__), .dinb(new_new_n1647__), .dout(new_new_n1655__));
  and1  g0663(.dina(new_new_n1655__), .dinb(new_new_n1646__), .dout(new_new_n1656__));
  or1   g0664(.dina(new_new_n1368__), .dinb(new_new_n2235__), .dout(new_new_n1657__));
  and1  g0665(.dina(new_new_n1382__), .dinb(new_new_n1374__), .dout(new_new_n1658__));
  or1   g0666(.dina(new_new_n1384__), .dinb(new_new_n1378__), .dout(new_new_n1659__));
  and1  g0667(.dina(new_new_n2237__), .dinb(new_new_n2239__), .dout(new_new_n1660__));
  and1  g0668(.dina(new_new_n2240__), .dinb(new_new_n2241__), .dout(new_new_n1661__));
  or1   g0669(.dina(new_new_n2237__), .dinb(new_new_n2239__), .dout(new_new_n1662__));
  or1   g0670(.dina(new_new_n1222__), .dinb(new_new_n2242__), .dout(new_new_n1663__));
  or1   g0671(.dina(new_new_n1314__), .dinb(new_new_n1224__), .dout(new_new_n1664__));
  and1  g0672(.dina(new_new_n1372__), .dinb(new_new_n1316__), .dout(new_new_n1665__));
  and1  g0673(.dina(new_new_n1665__), .dinb(new_new_n1664__), .dout(new_new_n1666__));
  and1  g0674(.dina(new_new_n1666__), .dinb(new_new_n1663__), .dout(new_new_n1667__));
  or1   g0675(.dina(new_new_n1176__), .dinb(new_new_n832__), .dout(new_new_n1668__));
  and1  g0676(.dina(new_new_n2244__), .dinb(new_new_n2246__), .dout(new_new_n1669__));
  or1   g0677(.dina(new_new_n2247__), .dinb(new_new_n2248__), .dout(new_new_n1670__));
  and1  g0678(.dina(new_new_n1670__), .dinb(new_new_n2249__), .dout(new_new_n1671__));
  or1   g0679(.dina(new_new_n1386__), .dinb(new_new_n1380__), .dout(new_new_n1672__));
  or1   g0680(.dina(new_new_n1418__), .dinb(new_new_n1408__), .dout(new_new_n1673__));
  and1  g0681(.dina(new_new_n1404__), .dinb(new_new_n1402__), .dout(new_new_n1674__));
  and1  g0682(.dina(new_new_n2251__), .dinb(new_new_n2252__), .dout(new_new_n1675__));
  and1  g0683(.dina(new_new_n2253__), .dinb(new_new_n2254__), .dout(new_new_n1676__));
  or1   g0684(.dina(new_new_n2244__), .dinb(new_new_n2246__), .dout(new_new_n1677__));
  or1   g0685(.dina(new_new_n1206__), .dinb(new_new_n1186__), .dout(new_new_n1678__));
  or1   g0686(.dina(new_new_n1678__), .dinb(new_new_n856__), .dout(new_new_n1679__));
  or1   g0687(.dina(new_new_n1679__), .dinb(new_new_n2255__), .dout(new_new_n1680__));
  and1  g0688(.dina(new_new_n2256__), .dinb(new_new_n2258__), .dout(new_new_n1681__));
  and1  g0689(.dina(new_new_n2259__), .dinb(new_new_n1235__), .dout(new_new_n1682__));
  and1  g0690(.dina(new_new_n2260__), .dinb(new_new_n1181__), .dout(new_new_n1683__));
  or1   g0691(.dina(new_new_n1683__), .dinb(new_new_n2261__), .dout(new_new_n1684__));
  or1   g0692(.dina(new_new_n1684__), .dinb(new_new_n1682__), .dout(new_new_n1685__));
  or1   g0693(.dina(new_new_n1685__), .dinb(new_new_n1681__), .dout(new_new_n1686__));
  or1   g0694(.dina(new_new_n2251__), .dinb(new_new_n2252__), .dout(new_new_n1687__));
  or1   g0695(.dina(new_new_n1398__), .dinb(new_new_n1330__), .dout(new_new_n1688__));
  or1   g0696(.dina(new_new_n1406__), .dinb(new_new_n1317__), .dout(new_new_n1689__));
  and1  g0697(.dina(new_new_n1689__), .dinb(new_new_n1332__), .dout(new_new_n1690__));
  and1  g0698(.dina(new_new_n1690__), .dinb(new_new_n1688__), .dout(new_new_n1691__));
  or1   g0699(.dina(new_new_n2262__), .dinb(new_new_n2263__), .dout(new_new_n1692__));
  or1   g0700(.dina(new_new_n1310__), .dinb(new_new_n1281__), .dout(new_new_n1693__));
  or1   g0701(.dina(new_new_n1693__), .dinb(new_new_n1288__), .dout(new_new_n1694__));
  or1   g0702(.dina(new_new_n2264__), .dinb(new_new_n1260__), .dout(new_new_n1695__));
  or1   g0703(.dina(new_new_n1695__), .dinb(new_new_n1320__), .dout(new_new_n1696__));
  and1  g0704(.dina(new_new_n2266__), .dinb(new_new_n1427__), .dout(new_new_n1697__));
  or1   g0705(.dina(new_new_n1697__), .dinb(new_new_n1388__), .dout(new_new_n1698__));
  and1  g0706(.dina(new_new_n2268__), .dinb(new_new_n2269__), .dout(new_new_n1699__));
  and1  g0707(.dina(new_new_n1699__), .dinb(new_new_n2266__), .dout(new_new_n1700__));
  or1   g0708(.dina(new_new_n2271__), .dinb(new_new_n2272__), .dout(new_new_n1701__));
  and1  g0709(.dina(new_new_n2273__), .dinb(new_new_n2274__), .dout(new_new_n1702__));
  and1  g0710(.dina(new_new_n1441__), .dinb(new_new_n2275__), .dout(new_new_n1703__));
  and1  g0711(.dina(new_new_n1703__), .dinb(new_new_n2267__), .dout(new_new_n1704__));
  or1   g0712(.dina(new_new_n1436__), .dinb(new_new_n1430__), .dout(new_new_n1705__));
  and1  g0713(.dina(new_new_n1425__), .dinb(new_new_n1419__), .dout(new_new_n1706__));
  and1  g0714(.dina(new_new_n1706__), .dinb(new_new_n1705__), .dout(new_new_n1707__));
  or1   g0715(.dina(new_new_n1707__), .dinb(new_new_n1704__), .dout(new_new_n1708__));
  and1  g0716(.dina(new_new_n1434__), .dinb(new_new_n2276__), .dout(new_new_n1709__));
  and1  g0717(.dina(new_new_n1709__), .dinb(new_new_n2277__), .dout(new_new_n1710__));
  and1  g0718(.dina(new_new_n2278__), .dinb(new_new_n2279__), .dout(new_new_n1711__));
  and1  g0719(.dina(new_new_n2280__), .dinb(new_new_n2282__), .dout(new_new_n1712__));
  and1  g0720(.dina(new_new_n1117__), .dinb(new_new_n2283__), .dout(new_new_n1713__));
  or1   g0721(.dina(new_new_n2258__), .dinb(new_new_n2285__), .dout(new_new_n1714__));
  or1   g0722(.dina(new_new_n942__), .dinb(new_new_n934__), .dout(new_new_n1715__));
  and1  g0723(.dina(new_new_n1715__), .dinb(new_new_n1714__), .dout(new_new_n1716__));
  and1  g0724(.dina(new_new_n2256__), .dinb(new_new_n2285__), .dout(new_new_n1717__));
  and1  g0725(.dina(new_new_n2260__), .dinb(new_new_n2286__), .dout(new_new_n1718__));
  or1   g0726(.dina(new_new_n1718__), .dinb(new_new_n2261__), .dout(new_new_n1719__));
  and1  g0727(.dina(new_new_n2259__), .dinb(new_new_n1267__), .dout(new_new_n1720__));
  or1   g0728(.dina(new_new_n1720__), .dinb(new_new_n1719__), .dout(new_new_n1721__));
  or1   g0729(.dina(new_new_n1721__), .dinb(new_new_n1717__), .dout(new_new_n1722__));
  or1   g0730(.dina(new_new_n2287__), .dinb(new_new_n2288__), .dout(new_new_n1723__));
  or1   g0731(.dina(new_new_n1334__), .dinb(new_new_n2242__), .dout(new_new_n1724__));
  and1  g0732(.dina(new_new_n1724__), .dinb(new_new_n1723__), .dout(new_new_n1725__));
  or1   g0733(.dina(new_new_n2278__), .dinb(new_new_n2289__), .dout(new_new_n1726__));
  or1   g0734(.dina(new_new_n1292__), .dinb(new_new_n1244__), .dout(new_new_n1727__));
  and1  g0735(.dina(new_new_n1727__), .dinb(new_new_n1726__), .dout(new_new_n1728__));
  or1   g0736(.dina(new_new_n2290__), .dinb(new_new_n1215__), .dout(new_new_n1729__));
  or1   g0737(.dina(new_new_n1226__), .dinb(new_new_n1216__), .dout(new_new_n1730__));
  and1  g0738(.dina(new_new_n1730__), .dinb(new_new_n1729__), .dout(new_new_n1731__));
  or1   g0739(.dina(new_new_n2282__), .dinb(new_new_n2291__), .dout(new_new_n1732__));
  or1   g0740(.dina(new_new_n1018__), .dinb(new_new_n1010__), .dout(new_new_n1733__));
  and1  g0741(.dina(new_new_n1733__), .dinb(new_new_n1732__), .dout(new_new_n1734__));
  or1   g0742(.dina(new_new_n2292__), .dinb(new_new_n2293__), .dout(new_new_n1735__));
  or1   g0743(.dina(new_new_n2238__), .dinb(new_new_n2245__), .dout(new_new_n1736__));
  and1  g0744(.dina(new_new_n1736__), .dinb(new_new_n1735__), .dout(new_new_n1737__));
  or1   g0745(.dina(new_new_n2294__), .dinb(new_new_n2295__), .dout(new_new_n1738__));
  and1  g0746(.dina(new_new_n1738__), .dinb(new_new_n2296__), .dout(new_new_n1739__));
  or1   g0747(.dina(new_new_n2297__), .dinb(new_new_n2298__), .dout(new_new_n1740__));
  or1   g0748(.dina(new_new_n2235__), .dinb(new_new_n1298__), .dout(new_new_n1741__));
  and1  g0749(.dina(new_new_n1741__), .dinb(new_new_n1740__), .dout(new_new_n1742__));
  and1  g0750(.dina(new_new_n2271__), .dinb(new_new_n2272__), .dout(new_new_n1743__));
  or1   g0751(.dina(new_new_n2299__), .dinb(new_new_n2300__), .dout(new_new_n1744__));
  or1   g0752(.dina(new_new_n1248__), .dinb(new_new_n1230__), .dout(new_new_n1745__));
  and1  g0753(.dina(new_new_n1745__), .dinb(new_new_n1744__), .dout(new_new_n1746__));
  or1   g0754(.dina(new_new_n868__), .dinb(new_new_n862__), .dout(new_new_n1747__));
  or1   g0755(.dina(new_new_n1747__), .dinb(new_new_n1200__), .dout(new_new_n1748__));
  or1   g0756(.dina(new_new_n1748__), .dinb(new_new_n2301__), .dout(new_new_n1749__));
  and1  g0757(.dina(new_new_n2303__), .dinb(new_new_n2304__), .dout(new_new_n1750__));
  and1  g0758(.dina(new_new_n1318__), .dinb(new_new_n2305__), .dout(new_new_n1751__));
  or1   g0759(.dina(new_new_n1751__), .dinb(new_new_n1331__), .dout(new_new_n1752__));
  or1   g0760(.dina(new_new_n1752__), .dinb(new_new_n1750__), .dout(new_new_n1753__));
  and1  g0761(.dina(new_new_n2306__), .dinb(new_new_n2307__), .dout(new_new_n1754__));
  and1  g0762(.dina(new_new_n2303__), .dinb(new_new_n2308__), .dout(new_new_n1755__));
  or1   g0763(.dina(new_new_n2309__), .dinb(new_new_n2310__), .dout(new_new_n1756__));
  or1   g0764(.dina(new_new_n2311__), .dinb(new_new_n1322__), .dout(new_new_n1757__));
  or1   g0765(.dina(new_new_n1004__), .dinb(new_new_n992__), .dout(new_new_n1758__));
  and1  g0766(.dina(new_new_n1758__), .dinb(new_new_n2312__), .dout(new_new_n1759__));
  and1  g0767(.dina(new_new_n1759__), .dinb(new_new_n1757__), .dout(new_new_n1760__));
  and1  g0768(.dina(new_new_n2313__), .dinb(new_new_n2314__), .dout(new_new_n1761__));
  or1   g0769(.dina(new_new_n1761__), .dinb(new_new_n2315__), .dout(new_new_n1762__));
  and1  g0770(.dina(new_new_n2317__), .dinb(new_new_n2318__), .dout(new_new_n1763__));
  and1  g0771(.dina(new_new_n2320__), .dinb(new_new_n2321__), .dout(new_new_n1764__));
  or1   g0772(.dina(new_new_n1764__), .dinb(new_new_n2323__), .dout(new_new_n1765__));
  or1   g0773(.dina(new_new_n1765__), .dinb(new_new_n1763__), .dout(new_new_n1766__));
  and1  g0774(.dina(new_new_n2317__), .dinb(new_new_n2324__), .dout(new_new_n1767__));
  and1  g0775(.dina(new_new_n2320__), .dinb(new_new_n2325__), .dout(new_new_n1768__));
  or1   g0776(.dina(new_new_n1768__), .dinb(new_new_n2323__), .dout(new_new_n1769__));
  or1   g0777(.dina(new_new_n2326__), .dinb(new_new_n2327__), .dout(new_new_n1770__));
  or1   g0778(.dina(new_new_n722__), .dinb(new_new_n706__), .dout(new_new_n1771__));
  or1   g0779(.dina(new_new_n784__), .dinb(new_new_n726__), .dout(new_new_n1772__));
  and1  g0780(.dina(new_new_n2329__), .dinb(new_new_n2331__), .dout(new_new_n1773__));
  and1  g0781(.dina(new_new_n2332__), .dinb(new_new_n2329__), .dout(new_new_n1774__));
  and1  g0782(.dina(new_new_n2333__), .dinb(new_new_n2335__), .dout(new_new_n1775__));
  or1   g0783(.dina(new_new_n2336__), .dinb(new_new_n714__), .dout(new_new_n1776__));
  and1  g0784(.dina(new_new_n2337__), .dinb(new_new_n2338__), .dout(new_new_n1777__));
  and1  g0785(.dina(new_new_n720__), .dinb(new_new_n2330__), .dout(new_new_n1778__));
  and1  g0786(.dina(new_new_n2335__), .dinb(new_new_n712__), .dout(new_new_n1779__));
  or1   g0787(.dina(new_new_n1779__), .dinb(new_new_n1778__), .dout(new_new_n1780__));
  buf1  g0788(.din(new_new_n1445__), .dout(G855));
  buf1  g0789(.din(new_new_n1446__), .dout(G856));
  buf1  g0790(.din(new_new_n2127__), .dout(G857));
  buf1  g0791(.din(new_new_n1449__), .dout(G858));
  buf1  g0792(.din(new_new_n1451__), .dout(G859));
  not1  g0793(.din(new_new_n1453__), .dout(G860));
  not1  g0794(.din(new_new_n1455__), .dout(G861));
  not1  g0795(.din(new_new_n1456__), .dout(G862));
  buf1  g0796(.din(new_new_n1457__), .dout(G863));
  not1  g0797(.din(new_new_n1459__), .dout(G864));
  not1  g0798(.din(new_new_n1460__), .dout(G865));
  buf1  g0799(.din(new_new_n1142__), .dout(G866));
  buf1  g0800(.din(new_new_n1461__), .dout(G867));
  buf1  g0801(.din(new_new_n1463__), .dout(G868));
  not1  g0802(.din(new_new_n1464__), .dout(G869));
  buf1  g0803(.din(new_new_n1491__), .dout(G870));
  buf1  g0804(.din(new_new_n1518__), .dout(G871));
  buf1  g0805(.din(new_new_n1534__), .dout(G872));
  buf1  g0806(.din(new_new_n1548__), .dout(G873));
  buf1  g0807(.din(new_new_n1564__), .dout(G874));
  buf1  g0808(.din(new_new_n1580__), .dout(G875));
  buf1  g0809(.din(new_new_n1592__), .dout(G876));
  buf1  g0810(.din(new_new_n1608__), .dout(G877));
  buf1  g0811(.din(new_new_n1624__), .dout(G878));
  buf1  g0812(.din(new_new_n1640__), .dout(G879));
  buf1  g0813(.din(new_new_n1656__), .dout(G880));
  buf1  g0814(.din(new_new_n2286__), .dout(n3148));
  buf1  g0815(.din(new_new_n709__), .dout(n3151));
  buf1  g0816(.din(new_new_n827__), .dout(n3154));
  buf1  g0817(.din(new_new_n829__), .dout(n3157));
  buf1  g0818(.din(new_new_n1177__), .dout(n3160));
  buf1  g0819(.din(new_new_n1187__), .dout(n3163));
  buf1  g0820(.din(new_new_n1189__), .dout(n3166));
  buf1  g0821(.din(new_new_n717__), .dout(n3169));
  buf1  g0822(.din(new_new_n839__), .dout(n3172));
  buf1  g0823(.din(new_new_n841__), .dout(n3175));
  buf1  g0824(.din(new_new_n843__), .dout(n3178));
  buf1  g0825(.din(new_new_n1179__), .dout(n3181));
  buf1  g0826(.din(new_new_n1183__), .dout(n3184));
  buf1  g0827(.din(new_new_n727__), .dout(n3187));
  buf1  g0828(.din(new_new_n851__), .dout(n3190));
  buf1  g0829(.din(new_new_n853__), .dout(n3193));
  buf1  g0830(.din(new_new_n729__), .dout(n3196));
  buf1  g0831(.din(new_new_n857__), .dout(n3199));
  buf1  g0832(.din(new_new_n859__), .dout(n3202));
  buf1  g0833(.din(new_new_n731__), .dout(n3205));
  buf1  g0834(.din(new_new_n863__), .dout(n3208));
  buf1  g0835(.din(new_new_n865__), .dout(n3211));
  buf1  g0836(.din(new_new_n733__), .dout(n3214));
  buf1  g0837(.din(new_new_n869__), .dout(n3217));
  buf1  g0838(.din(new_new_n871__), .dout(n3220));
  buf1  g0839(.din(new_new_n873__), .dout(n3223));
  buf1  g0840(.din(new_new_n1197__), .dout(n3226));
  buf1  g0841(.din(new_new_n1191__), .dout(n3229));
  buf1  g0842(.din(new_new_n739__), .dout(n3232));
  buf1  g0843(.din(new_new_n881__), .dout(n3235));
  buf1  g0844(.din(new_new_n883__), .dout(n3238));
  buf1  g0845(.din(new_new_n885__), .dout(n3241));
  buf1  g0846(.din(new_new_n741__), .dout(n3244));
  buf1  g0847(.din(new_new_n889__), .dout(n3247));
  buf1  g0848(.din(new_new_n891__), .dout(n3250));
  buf1  g0849(.din(new_new_n893__), .dout(n3253));
  buf1  g0850(.din(new_new_n743__), .dout(n3256));
  buf1  g0851(.din(new_new_n897__), .dout(n3259));
  buf1  g0852(.din(new_new_n899__), .dout(n3262));
  buf1  g0853(.din(new_new_n901__), .dout(n3265));
  buf1  g0854(.din(new_new_n745__), .dout(n3268));
  buf1  g0855(.din(new_new_n905__), .dout(n3271));
  buf1  g0856(.din(new_new_n907__), .dout(n3274));
  buf1  g0857(.din(new_new_n909__), .dout(n3277));
  buf1  g0858(.din(new_new_n747__), .dout(n3280));
  buf1  g0859(.din(new_new_n913__), .dout(n3283));
  buf1  g0860(.din(new_new_n915__), .dout(n3286));
  buf1  g0861(.din(new_new_n917__), .dout(n3289));
  buf1  g0862(.din(new_new_n749__), .dout(n3292));
  buf1  g0863(.din(new_new_n921__), .dout(n3295));
  buf1  g0864(.din(new_new_n923__), .dout(n3298));
  buf1  g0865(.din(new_new_n925__), .dout(n3301));
  buf1  g0866(.din(new_new_n751__), .dout(n3304));
  buf1  g0867(.din(new_new_n929__), .dout(n3307));
  buf1  g0868(.din(new_new_n931__), .dout(n3310));
  buf1  g0869(.din(new_new_n2284__), .dout(n3313));
  buf1  g0870(.din(new_new_n753__), .dout(n3316));
  buf1  g0871(.din(new_new_n937__), .dout(n3319));
  buf1  g0872(.din(new_new_n939__), .dout(n3322));
  buf1  g0873(.din(new_new_n2257__), .dout(n3325));
  buf1  g0874(.din(new_new_n755__), .dout(n3328));
  buf1  g0875(.din(new_new_n945__), .dout(n3331));
  buf1  g0876(.din(new_new_n947__), .dout(n3334));
  buf1  g0877(.din(new_new_n2288__), .dout(n3337));
  buf1  g0878(.din(new_new_n757__), .dout(n3340));
  buf1  g0879(.din(new_new_n953__), .dout(n3343));
  buf1  g0880(.din(new_new_n2287__), .dout(n3346));
  buf1  g0881(.din(new_new_n759__), .dout(n3349));
  buf1  g0882(.din(new_new_n959__), .dout(n3352));
  buf1  g0883(.din(new_new_n761__), .dout(n3355));
  buf1  g0884(.din(new_new_n2289__), .dout(n3358));
  buf1  g0885(.din(new_new_n763__), .dout(n3361));
  buf1  g0886(.din(new_new_n2290__), .dout(n3364));
  buf1  g0887(.din(new_new_n765__), .dout(n3367));
  buf1  g0888(.din(new_new_n767__), .dout(n3370));
  buf1  g0889(.din(new_new_n973__), .dout(n3373));
  buf1  g0890(.din(new_new_n975__), .dout(n3376));
  buf1  g0891(.din(new_new_n977__), .dout(n3379));
  buf1  g0892(.din(new_new_n769__), .dout(n3382));
  buf1  g0893(.din(new_new_n981__), .dout(n3385));
  buf1  g0894(.din(new_new_n983__), .dout(n3388));
  buf1  g0895(.din(new_new_n985__), .dout(n3391));
  buf1  g0896(.din(new_new_n771__), .dout(n3394));
  buf1  g0897(.din(new_new_n989__), .dout(n3397));
  buf1  g0898(.din(new_new_n773__), .dout(n3400));
  buf1  g0899(.din(new_new_n993__), .dout(n3403));
  buf1  g0900(.din(new_new_n775__), .dout(n3406));
  buf1  g0901(.din(new_new_n777__), .dout(n3409));
  buf1  g0902(.din(new_new_n779__), .dout(n3412));
  buf1  g0903(.din(new_new_n1001__), .dout(n3415));
  buf1  g0904(.din(new_new_n785__), .dout(n3418));
  buf1  g0905(.din(new_new_n1005__), .dout(n3421));
  buf1  g0906(.din(new_new_n1007__), .dout(n3424));
  buf1  g0907(.din(new_new_n2291__), .dout(n3427));
  buf1  g0908(.din(new_new_n787__), .dout(n3430));
  buf1  g0909(.din(new_new_n1013__), .dout(n3433));
  buf1  g0910(.din(new_new_n1015__), .dout(n3436));
  buf1  g0911(.din(new_new_n2281__), .dout(n3439));
  buf1  g0912(.din(new_new_n789__), .dout(n3442));
  buf1  g0913(.din(new_new_n1021__), .dout(n3445));
  buf1  g0914(.din(new_new_n1023__), .dout(n3448));
  buf1  g0915(.din(new_new_n2293__), .dout(n3451));
  buf1  g0916(.din(new_new_n791__), .dout(n3454));
  buf1  g0917(.din(new_new_n1029__), .dout(n3457));
  buf1  g0918(.din(new_new_n1031__), .dout(n3460));
  buf1  g0919(.din(new_new_n2292__), .dout(n3463));
  buf1  g0920(.din(new_new_n793__), .dout(n3466));
  buf1  g0921(.din(new_new_n1037__), .dout(n3469));
  buf1  g0922(.din(new_new_n2297__), .dout(n3472));
  buf1  g0923(.din(new_new_n795__), .dout(n3475));
  buf1  g0924(.din(new_new_n1043__), .dout(n3478));
  buf1  g0925(.din(new_new_n2298__), .dout(n3481));
  buf1  g0926(.din(new_new_n797__), .dout(n3484));
  buf1  g0927(.din(new_new_n2299__), .dout(n3487));
  buf1  g0928(.din(new_new_n799__), .dout(n3490));
  buf1  g0929(.din(new_new_n2300__), .dout(n3493));
  buf1  g0930(.din(new_new_n801__), .dout(n3496));
  buf1  g0931(.din(new_new_n1057__), .dout(n3499));
  buf1  g0932(.din(new_new_n1059__), .dout(n3502));
  buf1  g0933(.din(new_new_n1061__), .dout(n3505));
  buf1  g0934(.din(new_new_n803__), .dout(n3508));
  buf1  g0935(.din(new_new_n1065__), .dout(n3511));
  buf1  g0936(.din(new_new_n1067__), .dout(n3514));
  buf1  g0937(.din(new_new_n2279__), .dout(n3517));
  buf1  g0938(.din(new_new_n805__), .dout(n3520));
  buf1  g0939(.din(new_new_n1073__), .dout(n3523));
  buf1  g0940(.din(new_new_n1075__), .dout(n3526));
  buf1  g0941(.din(new_new_n1077__), .dout(n3529));
  buf1  g0942(.din(new_new_n807__), .dout(n3532));
  buf1  g0943(.din(new_new_n1081__), .dout(n3535));
  buf1  g0944(.din(new_new_n1083__), .dout(n3538));
  buf1  g0945(.din(new_new_n1085__), .dout(n3541));
  buf1  g0946(.din(new_new_n809__), .dout(n3544));
  buf1  g0947(.din(new_new_n1089__), .dout(n3547));
  buf1  g0948(.din(new_new_n1091__), .dout(n3550));
  buf1  g0949(.din(new_new_n1093__), .dout(n3553));
  buf1  g0950(.din(new_new_n811__), .dout(n3556));
  buf1  g0951(.din(new_new_n1097__), .dout(n3559));
  buf1  g0952(.din(new_new_n1099__), .dout(n3562));
  buf1  g0953(.din(new_new_n1101__), .dout(n3565));
  buf1  g0954(.din(new_new_n813__), .dout(n3568));
  buf1  g0955(.din(new_new_n1105__), .dout(n3571));
  buf1  g0956(.din(new_new_n1107__), .dout(n3574));
  buf1  g0957(.din(new_new_n2283__), .dout(n3577));
  buf1  g0958(.din(new_new_n815__), .dout(n3580));
  buf1  g0959(.din(new_new_n1113__), .dout(n3583));
  buf1  g0960(.din(new_new_n1115__), .dout(n3586));
  buf1  g0961(.din(new_new_n817__), .dout(n3589));
  buf1  g0962(.din(new_new_n1119__), .dout(n3592));
  buf1  g0963(.din(new_new_n1121__), .dout(n3595));
  buf1  g0964(.din(new_new_n1123__), .dout(n3598));
  buf1  g0965(.din(new_new_n819__), .dout(n3601));
  buf1  g0966(.din(new_new_n1237__), .dout(n3604));
  buf1  g0967(.din(new_new_n821__), .dout(n3607));
  buf1  g0968(.din(new_new_n1131__), .dout(n3610));
  buf1  g0969(.din(new_new_n1133__), .dout(n3613));
  buf1  g0970(.din(new_new_n1135__), .dout(n3616));
  buf1  g0971(.din(new_new_n1209__), .dout(n3619));
  buf1  g0972(.din(new_new_n1201__), .dout(n3622));
  buf1  g0973(.din(new_new_n1203__), .dout(n3625));
  buf1  g0974(.din(new_new_n1199__), .dout(n3628));
  buf1  g0975(.din(new_new_n1233__), .dout(n3631));
  buf1  g0976(.din(new_new_n1239__), .dout(n3634));
  buf1  g0977(.din(new_new_n1251__), .dout(n3637));
  buf1  g0978(.din(new_new_n1253__), .dout(n3640));
  buf1  g0979(.din(new_new_n1255__), .dout(n3643));
  buf1  g0980(.din(new_new_n1277__), .dout(n3646));
  buf1  g0981(.din(new_new_n1279__), .dout(n3649));
  buf1  g0982(.din(new_new_n1303__), .dout(n3652));
  buf1  g0983(.din(new_new_n1305__), .dout(n3655));
  buf1  g0984(.din(new_new_n1307__), .dout(n3658));
  buf1  g0985(.din(new_new_n1323__), .dout(n3661));
  buf1  g0986(.din(new_new_n1325__), .dout(n3664));
  buf1  g0987(.din(new_new_n1361__), .dout(n3667));
  buf1  g0988(.din(new_new_n1367__), .dout(n3670));
  buf1  g0989(.din(new_new_n1257__), .dout(n3673));
  buf1  g0990(.din(new_new_n2306__), .dout(n3676));
  buf1  g0991(.din(new_new_n1261__), .dout(n3679));
  buf1  g0992(.din(new_new_n1263__), .dout(n3682));
  buf1  g0993(.din(new_new_n1265__), .dout(n3685));
  buf1  g0994(.din(new_new_n1269__), .dout(n3688));
  buf1  g0995(.din(new_new_n1271__), .dout(n3691));
  buf1  g0996(.din(new_new_n1273__), .dout(n3694));
  buf1  g0997(.din(new_new_n1275__), .dout(n3697));
  buf1  g0998(.din(new_new_n1377__), .dout(n3700));
  buf1  g0999(.din(new_new_n1383__), .dout(n3703));
  buf1  g1000(.din(new_new_n1285__), .dout(n3706));
  buf1  g1001(.din(new_new_n1283__), .dout(n3709));
  buf1  g1002(.din(new_new_n1287__), .dout(n3712));
  buf1  g1003(.din(new_new_n1289__), .dout(n3715));
  buf1  g1004(.din(new_new_n1309__), .dout(n3718));
  not1  g1005(.din(new_new_n2241__), .dout(n3721));
  buf1  g1006(.din(new_new_n2264__), .dout(n3724));
  not1  g1007(.din(new_new_n2236__), .dout(n3727));
  not1  g1008(.din(new_new_n2240__), .dout(n3730));
  buf1  g1009(.din(new_new_n1327__), .dout(n3733));
  not1  g1010(.din(new_new_n2248__), .dout(n3736));
  not1  g1011(.din(new_new_n2247__), .dout(n3739));
  buf1  g1012(.din(new_new_n2302__), .dout(n3742));
  buf1  g1013(.din(new_new_n1369__), .dout(n3745));
  buf1  g1014(.din(new_new_n1375__), .dout(n3748));
  not1  g1015(.din(new_new_n2249__), .dout(n3751));
  buf1  g1016(.din(new_new_n1379__), .dout(n3754));
  not1  g1017(.din(new_new_n2243__), .dout(n3757));
  buf1  g1018(.din(new_new_n1385__), .dout(n3760));
  buf1  g1019(.din(new_new_n1405__), .dout(n3763));
  buf1  g1020(.din(new_new_n1407__), .dout(n3766));
  buf1  g1021(.din(new_new_n1417__), .dout(n3769));
  not1  g1022(.din(new_new_n2255__), .dout(n3772));
  buf1  g1023(.din(new_new_n1397__), .dout(n3775));
  not1  g1024(.din(new_new_n2295__), .dout(n3778));
  buf1  g1025(.din(new_new_n1399__), .dout(n3781));
  not1  g1026(.din(new_new_n2294__), .dout(n3784));
  not1  g1027(.din(new_new_n2254__), .dout(n3787));
  not1  g1028(.din(new_new_n2253__), .dout(n3790));
  not1  g1029(.din(new_new_n2250__), .dout(n3793));
  buf1  g1030(.din(new_new_n1387__), .dout(n3796));
  buf1  g1031(.din(new_new_n1389__), .dout(n3799));
  buf1  g1032(.din(new_new_n1391__), .dout(n3802));
  buf1  g1033(.din(new_new_n1393__), .dout(n3805));
  buf1  g1034(.din(new_new_n1395__), .dout(n3808));
  buf1  g1035(.din(new_new_n2305__), .dout(n3811));
  buf1  g1036(.din(new_new_n1409__), .dout(n3814));
  buf1  g1037(.din(new_new_n1411__), .dout(n3817));
  buf1  g1038(.din(new_new_n1413__), .dout(n3820));
  buf1  g1039(.din(new_new_n1415__), .dout(n3823));
  not1  g1040(.din(new_new_n2263__), .dout(n3826));
  not1  g1041(.din(new_new_n2262__), .dout(n3829));
  buf1  g1042(.din(new_new_n2275__), .dout(n3832));
  buf1  g1043(.din(new_new_n1429__), .dout(n3835));
  buf1  g1044(.din(new_new_n2269__), .dout(n3838));
  buf1  g1045(.din(new_new_n2267__), .dout(n3841));
  buf1  g1046(.din(new_new_n2268__), .dout(n3844));
  buf1  g1047(.din(new_new_n2304__), .dout(n3847));
  buf1  g1048(.din(new_new_n2307__), .dout(n3850));
  not1  g1049(.din(new_new_n2296__), .dout(n3853));
  buf1  g1050(.din(new_new_n1045__), .dout(n3856));
  not1  g1051(.din(new_new_n2301__), .dout(n3859));
  buf1  g1052(.din(new_new_n2280__), .dout(n3862));
  not1  g1053(.din(new_new_n2274__), .dout(n3865));
  not1  g1054(.din(new_new_n2270__), .dout(n3868));
  not1  g1055(.din(new_new_n2273__), .dout(n3871));
  buf1  g1056(.din(new_new_n2276__), .dout(n3874));
  buf1  g1057(.din(new_new_n1433__), .dout(n3877));
  not1  g1058(.din(new_new_n2311__), .dout(n3880));
  not1  g1059(.din(new_new_n2312__), .dout(n3883));
  not1  g1060(.din(new_new_n2319__), .dout(n3886));
  buf1  g1061(.din(new_new_n2277__), .dout(n3889));
  buf1  g1062(.din(new_new_n2321__), .dout(n3892));
  not1  g1063(.din(new_new_n2314__), .dout(n3895));
  not1  g1064(.din(new_new_n2313__), .dout(n3898));
  buf1  g1065(.din(new_new_n2318__), .dout(n3901));
  buf1  g1066(.din(new_new_n2316__), .dout(n3904));
  buf1  g1067(.din(new_new_n2322__), .dout(n3907));
  buf1  g1068(.din(new_new_n2308__), .dout(n3910));
  buf1  g1069(.din(new_new_n1711__), .dout(n3913));
  buf1  g1070(.din(new_new_n1712__), .dout(n3916));
  buf1  g1071(.din(new_new_n2310__), .dout(n3919));
  buf1  g1072(.din(new_new_n1713__), .dout(n3922));
  buf1  g1073(.din(new_new_n1716__), .dout(n3925));
  buf1  g1074(.din(new_new_n1722__), .dout(n3928));
  buf1  g1075(.din(new_new_n1725__), .dout(n3931));
  buf1  g1076(.din(new_new_n1728__), .dout(n3934));
  buf1  g1077(.din(new_new_n1731__), .dout(n3937));
  buf1  g1078(.din(new_new_n1734__), .dout(n3940));
  buf1  g1079(.din(new_new_n1737__), .dout(n3943));
  not1  g1080(.din(new_new_n1739__), .dout(n3946));
  buf1  g1081(.din(new_new_n1742__), .dout(n3949));
  not1  g1082(.din(new_new_n2315__), .dout(n3952));
  buf1  g1083(.din(new_new_n1746__), .dout(n3955));
  not1  g1084(.din(new_new_n1749__), .dout(n3958));
  buf1  g1085(.din(new_new_n2309__), .dout(n3961));
  buf1  g1086(.din(new_new_n2325__), .dout(n3964));
  buf1  g1087(.din(new_new_n1754__), .dout(n3967));
  buf1  g1088(.din(new_new_n1755__), .dout(n3970));
  buf1  g1089(.din(new_new_n2324__), .dout(n3973));
  buf1  g1090(.din(new_new_n1756__), .dout(n3976));
  buf1  g1091(.din(new_new_n2327__), .dout(n3979));
  not1  g1092(.din(new_new_n1760__), .dout(n3982));
  not1  g1093(.din(new_new_n1762__), .dout(n3985));
  buf1  g1094(.din(new_new_n2326__), .dout(n3988));
  buf1  g1095(.din(new_new_n705__), .dout(n3991));
  buf1  g1096(.din(new_new_n2330__), .dout(n3994));
  buf1  g1097(.din(new_new_n2334__), .dout(n3997));
  buf1  g1098(.din(new_new_n721__), .dout(n4000));
  buf1  g1099(.din(new_new_n2333__), .dout(n4003));
  buf1  g1100(.din(new_new_n963__), .dout(n4006));
  buf1  g1101(.din(new_new_n1049__), .dout(n4009));
  buf1  g1102(.din(new_new_n1767__), .dout(n4012));
  buf1  g1103(.din(new_new_n1769__), .dout(n4015));
  buf1  g1104(.din(new_new_n997__), .dout(n4018));
  buf1  g1105(.din(new_new_n1127__), .dout(n4021));
  buf1  g1106(.din(new_new_n2331__), .dout(n4024));
  buf1  g1107(.din(new_new_n713__), .dout(n4027));
  buf1  g1108(.din(new_new_n2338__), .dout(n4030));
  buf1  g1109(.din(new_new_n2337__), .dout(n4033));
  buf1  g1110(.din(new_new_n1770__), .dout(n4036));
  not1  g1111(.din(new_new_n2336__), .dout(n4039));
  not1  g1112(.din(new_new_n2332__), .dout(n4042));
  buf1  g1113(.din(new_new_n781__), .dout(n4045));
  buf1  g1114(.din(new_new_n1773__), .dout(n4048));
  buf1  g1115(.din(new_new_n1774__), .dout(n4051));
  buf1  g1116(.din(new_new_n1775__), .dout(n4054));
  buf1  g1117(.din(new_new_n723__), .dout(n4057));
  buf1  g1118(.din(new_new_n823__), .dout(n4060));
  buf1  g1119(.din(new_new_n735__), .dout(n4063));
  not1  g1120(.din(new_new_n1776__), .dout(n4066));
  buf1  g1121(.din(new_new_n1777__), .dout(n4069));
  buf1  g1122(.din(new_new_n1780__), .dout(n4072));
  buf1  g1123(.din(new_new_n838__), .dout(new_new_n2116__));
  buf1  g1124(.din(new_new_n1444__), .dout(new_new_n2117__));
  buf1  g1125(.din(new_new_n878__), .dout(new_new_n2118__));
  buf1  g1126(.din(new_new_n846__), .dout(new_new_n2119__));
  buf1  g1127(.din(new_new_n2119__), .dout(new_new_n2120__));
  buf1  g1128(.din(new_new_n845__), .dout(new_new_n2121__));
  buf1  g1129(.din(new_new_n1450__), .dout(new_new_n2122__));
  buf1  g1130(.din(new_new_n1452__), .dout(new_new_n2123__));
  buf1  g1131(.din(new_new_n850__), .dout(new_new_n2124__));
  buf1  g1132(.din(new_new_n1454__), .dout(new_new_n2125__));
  buf1  g1133(.din(new_new_n1458__), .dout(new_new_n2126__));
  buf1  g1134(.din(new_new_n1448__), .dout(new_new_n2127__));
  buf1  g1135(.din(new_new_n1300__), .dout(new_new_n2128__));
  buf1  g1136(.din(new_new_n1348__), .dout(new_new_n2129__));
  buf1  g1137(.din(new_new_n1344__), .dout(new_new_n2130__));
  buf1  g1138(.din(new_new_n1347__), .dout(new_new_n2131__));
  buf1  g1139(.din(new_new_n1343__), .dout(new_new_n2132__));
  buf1  g1140(.din(new_new_n1469__), .dout(new_new_n2133__));
  buf1  g1141(.din(new_new_n979__), .dout(new_new_n2134__));
  buf1  g1142(.din(new_new_n2134__), .dout(new_new_n2135__));
  buf1  g1143(.din(new_new_n2134__), .dout(new_new_n2136__));
  buf1  g1144(.din(new_new_n1470__), .dout(new_new_n2137__));
  buf1  g1145(.din(new_new_n980__), .dout(new_new_n2138__));
  buf1  g1146(.din(new_new_n2138__), .dout(new_new_n2139__));
  buf1  g1147(.din(new_new_n2138__), .dout(new_new_n2140__));
  buf1  g1148(.din(new_new_n1352__), .dout(new_new_n2141__));
  buf1  g1149(.din(new_new_n1350__), .dout(new_new_n2142__));
  buf1  g1150(.din(new_new_n1351__), .dout(new_new_n2143__));
  buf1  g1151(.din(new_new_n1349__), .dout(new_new_n2144__));
  buf1  g1152(.din(new_new_n1481__), .dout(new_new_n2145__));
  buf1  g1153(.din(new_new_n987__), .dout(new_new_n2146__));
  buf1  g1154(.din(new_new_n1482__), .dout(new_new_n2147__));
  buf1  g1155(.din(new_new_n988__), .dout(new_new_n2148__));
  buf1  g1156(.din(new_new_n1356__), .dout(new_new_n2149__));
  buf1  g1157(.din(new_new_n1354__), .dout(new_new_n2150__));
  buf1  g1158(.din(new_new_n1355__), .dout(new_new_n2151__));
  buf1  g1159(.din(new_new_n1353__), .dout(new_new_n2152__));
  buf1  g1160(.din(new_new_n1496__), .dout(new_new_n2153__));
  buf1  g1161(.din(new_new_n1497__), .dout(new_new_n2154__));
  buf1  g1162(.din(new_new_n1364__), .dout(new_new_n2155__));
  buf1  g1163(.din(new_new_n1360__), .dout(new_new_n2156__));
  buf1  g1164(.din(new_new_n1363__), .dout(new_new_n2157__));
  buf1  g1165(.din(new_new_n1359__), .dout(new_new_n2158__));
  buf1  g1166(.din(new_new_n1508__), .dout(new_new_n2159__));
  buf1  g1167(.din(new_new_n1063__), .dout(new_new_n2160__));
  buf1  g1168(.din(new_new_n1509__), .dout(new_new_n2161__));
  buf1  g1169(.din(new_new_n1064__), .dout(new_new_n2162__));
  buf1  g1170(.din(new_new_n1096__), .dout(new_new_n2163__));
  buf1  g1171(.din(new_new_n2163__), .dout(new_new_n2164__));
  buf1  g1172(.din(new_new_n2164__), .dout(new_new_n2165__));
  buf1  g1173(.din(new_new_n2164__), .dout(new_new_n2166__));
  buf1  g1174(.din(new_new_n2163__), .dout(new_new_n2167__));
  buf1  g1175(.din(new_new_n2167__), .dout(new_new_n2168__));
  buf1  g1176(.din(new_new_n2167__), .dout(new_new_n2169__));
  buf1  g1177(.din(new_new_n1080__), .dout(new_new_n2170__));
  buf1  g1178(.din(new_new_n2170__), .dout(new_new_n2171__));
  buf1  g1179(.din(new_new_n2171__), .dout(new_new_n2172__));
  buf1  g1180(.din(new_new_n2172__), .dout(new_new_n2173__));
  buf1  g1181(.din(new_new_n2172__), .dout(new_new_n2174__));
  buf1  g1182(.din(new_new_n2171__), .dout(new_new_n2175__));
  buf1  g1183(.din(new_new_n2175__), .dout(new_new_n2176__));
  buf1  g1184(.din(new_new_n2170__), .dout(new_new_n2177__));
  buf1  g1185(.din(new_new_n2177__), .dout(new_new_n2178__));
  buf1  g1186(.din(new_new_n2177__), .dout(new_new_n2179__));
  buf1  g1187(.din(new_new_n1088__), .dout(new_new_n2180__));
  buf1  g1188(.din(new_new_n2180__), .dout(new_new_n2181__));
  buf1  g1189(.din(new_new_n2181__), .dout(new_new_n2182__));
  buf1  g1190(.din(new_new_n2181__), .dout(new_new_n2183__));
  buf1  g1191(.din(new_new_n2180__), .dout(new_new_n2184__));
  buf1  g1192(.din(new_new_n2184__), .dout(new_new_n2185__));
  buf1  g1193(.din(new_new_n2184__), .dout(new_new_n2186__));
  buf1  g1194(.din(new_new_n1104__), .dout(new_new_n2187__));
  buf1  g1195(.din(new_new_n2187__), .dout(new_new_n2188__));
  buf1  g1196(.din(new_new_n2188__), .dout(new_new_n2189__));
  buf1  g1197(.din(new_new_n2188__), .dout(new_new_n2190__));
  buf1  g1198(.din(new_new_n2187__), .dout(new_new_n2191__));
  buf1  g1199(.din(new_new_n2191__), .dout(new_new_n2192__));
  buf1  g1200(.din(new_new_n2191__), .dout(new_new_n2193__));
  buf1  g1201(.din(new_new_n1366__), .dout(new_new_n2194__));
  buf1  g1202(.din(new_new_n2194__), .dout(new_new_n2195__));
  buf1  g1203(.din(new_new_n2195__), .dout(new_new_n2196__));
  buf1  g1204(.din(new_new_n2195__), .dout(new_new_n2197__));
  buf1  g1205(.din(new_new_n2194__), .dout(new_new_n2198__));
  buf1  g1206(.din(new_new_n2198__), .dout(new_new_n2199__));
  buf1  g1207(.din(new_new_n2198__), .dout(new_new_n2200__));
  buf1  g1208(.din(new_new_n1072__), .dout(new_new_n2201__));
  buf1  g1209(.din(new_new_n2201__), .dout(new_new_n2202__));
  buf1  g1210(.din(new_new_n2202__), .dout(new_new_n2203__));
  buf1  g1211(.din(new_new_n2202__), .dout(new_new_n2204__));
  buf1  g1212(.din(new_new_n2201__), .dout(new_new_n2205__));
  buf1  g1213(.din(new_new_n2205__), .dout(new_new_n2206__));
  buf1  g1214(.din(new_new_n1112__), .dout(new_new_n2207__));
  buf1  g1215(.din(new_new_n1168__), .dout(new_new_n2208__));
  buf1  g1216(.din(new_new_n1550__), .dout(new_new_n2209__));
  buf1  g1217(.din(new_new_n1345__), .dout(new_new_n2210__));
  buf1  g1218(.din(new_new_n1011__), .dout(new_new_n2211__));
  buf1  g1219(.din(new_new_n1346__), .dout(new_new_n2212__));
  buf1  g1220(.din(new_new_n2212__), .dout(new_new_n2213__));
  buf1  g1221(.din(new_new_n1012__), .dout(new_new_n2214__));
  buf1  g1222(.din(new_new_n2214__), .dout(new_new_n2215__));
  buf1  g1223(.din(new_new_n1302__), .dout(new_new_n2216__));
  buf1  g1224(.din(new_new_n1020__), .dout(new_new_n2217__));
  buf1  g1225(.din(new_new_n1358__), .dout(new_new_n2218__));
  buf1  g1226(.din(new_new_n1338__), .dout(new_new_n2219__));
  buf1  g1227(.din(new_new_n2219__), .dout(new_new_n2220__));
  buf1  g1228(.din(new_new_n1357__), .dout(new_new_n2221__));
  buf1  g1229(.din(new_new_n1337__), .dout(new_new_n2222__));
  buf1  g1230(.din(new_new_n1586__), .dout(new_new_n2223__));
  buf1  g1231(.din(new_new_n1585__), .dout(new_new_n2224__));
  buf1  g1232(.din(new_new_n1590__), .dout(new_new_n2225__));
  buf1  g1233(.din(new_new_n1583__), .dout(new_new_n2226__));
  buf1  g1234(.din(new_new_n1582__), .dout(new_new_n2227__));
  buf1  g1235(.din(new_new_n2227__), .dout(new_new_n2228__));
  buf1  g1236(.din(new_new_n1228__), .dout(new_new_n2229__));
  buf1  g1237(.din(new_new_n1594__), .dout(new_new_n2230__));
  buf1  g1238(.din(new_new_n1610__), .dout(new_new_n2231__));
  buf1  g1239(.din(new_new_n1626__), .dout(new_new_n2232__));
  buf1  g1240(.din(new_new_n1296__), .dout(new_new_n2233__));
  buf1  g1241(.din(new_new_n1642__), .dout(new_new_n2234__));
  buf1  g1242(.din(new_new_n1340__), .dout(new_new_n2235__));
  buf1  g1243(.din(new_new_n1658__), .dout(new_new_n2236__));
  buf1  g1244(.din(new_new_n2236__), .dout(new_new_n2237__));
  buf1  g1245(.din(new_new_n1034__), .dout(new_new_n2238__));
  buf1  g1246(.din(new_new_n2238__), .dout(new_new_n2239__));
  buf1  g1247(.din(new_new_n1659__), .dout(new_new_n2240__));
  buf1  g1248(.din(new_new_n1657__), .dout(new_new_n2241__));
  buf1  g1249(.din(new_new_n950__), .dout(new_new_n2242__));
  buf1  g1250(.din(new_new_n1667__), .dout(new_new_n2243__));
  buf1  g1251(.din(new_new_n2243__), .dout(new_new_n2244__));
  buf1  g1252(.din(new_new_n1026__), .dout(new_new_n2245__));
  buf1  g1253(.din(new_new_n2245__), .dout(new_new_n2246__));
  buf1  g1254(.din(new_new_n1661__), .dout(new_new_n2247__));
  buf1  g1255(.din(new_new_n1660__), .dout(new_new_n2248__));
  buf1  g1256(.din(new_new_n1662__), .dout(new_new_n2249__));
  buf1  g1257(.din(new_new_n1674__), .dout(new_new_n2250__));
  buf1  g1258(.din(new_new_n2250__), .dout(new_new_n2251__));
  buf1  g1259(.din(new_new_n1400__), .dout(new_new_n2252__));
  buf1  g1260(.din(new_new_n1673__), .dout(new_new_n2253__));
  buf1  g1261(.din(new_new_n1672__), .dout(new_new_n2254__));
  buf1  g1262(.din(new_new_n1668__), .dout(new_new_n2255__));
  buf1  g1263(.din(new_new_n1221__), .dout(new_new_n2256__));
  buf1  g1264(.din(new_new_n941__), .dout(new_new_n2257__));
  buf1  g1265(.din(new_new_n2257__), .dout(new_new_n2258__));
  buf1  g1266(.din(new_new_n1313__), .dout(new_new_n2259__));
  buf1  g1267(.din(new_new_n1293__), .dout(new_new_n2260__));
  buf1  g1268(.din(new_new_n1315__), .dout(new_new_n2261__));
  buf1  g1269(.din(new_new_n1676__), .dout(new_new_n2262__));
  buf1  g1270(.din(new_new_n1675__), .dout(new_new_n2263__));
  buf1  g1271(.din(new_new_n1311__), .dout(new_new_n2264__));
  buf1  g1272(.din(new_new_n1437__), .dout(new_new_n2265__));
  buf1  g1273(.din(new_new_n2265__), .dout(new_new_n2266__));
  buf1  g1274(.din(new_new_n2265__), .dout(new_new_n2267__));
  buf1  g1275(.din(new_new_n1439__), .dout(new_new_n2268__));
  buf1  g1276(.din(new_new_n1435__), .dout(new_new_n2269__));
  buf1  g1277(.din(new_new_n1691__), .dout(new_new_n2270__));
  buf1  g1278(.din(new_new_n2270__), .dout(new_new_n2271__));
  buf1  g1279(.din(new_new_n1046__), .dout(new_new_n2272__));
  buf1  g1280(.din(new_new_n1692__), .dout(new_new_n2273__));
  buf1  g1281(.din(new_new_n1687__), .dout(new_new_n2274__));
  buf1  g1282(.din(new_new_n1421__), .dout(new_new_n2275__));
  buf1  g1283(.din(new_new_n1431__), .dout(new_new_n2276__));
  buf1  g1284(.din(new_new_n1700__), .dout(new_new_n2277__));
  buf1  g1285(.din(new_new_n1291__), .dout(new_new_n2278__));
  buf1  g1286(.din(new_new_n1069__), .dout(new_new_n2279__));
  buf1  g1287(.din(new_new_n1686__), .dout(new_new_n2280__));
  buf1  g1288(.din(new_new_n1017__), .dout(new_new_n2281__));
  buf1  g1289(.din(new_new_n2281__), .dout(new_new_n2282__));
  buf1  g1290(.din(new_new_n1109__), .dout(new_new_n2283__));
  buf1  g1291(.din(new_new_n933__), .dout(new_new_n2284__));
  buf1  g1292(.din(new_new_n2284__), .dout(new_new_n2285__));
  buf1  g1293(.din(new_new_n1185__), .dout(new_new_n2286__));
  buf1  g1294(.din(new_new_n1333__), .dout(new_new_n2287__));
  buf1  g1295(.din(new_new_n949__), .dout(new_new_n2288__));
  buf1  g1296(.din(new_new_n1243__), .dout(new_new_n2289__));
  buf1  g1297(.din(new_new_n1225__), .dout(new_new_n2290__));
  buf1  g1298(.din(new_new_n1009__), .dout(new_new_n2291__));
  buf1  g1299(.din(new_new_n1033__), .dout(new_new_n2292__));
  buf1  g1300(.din(new_new_n1025__), .dout(new_new_n2293__));
  buf1  g1301(.din(new_new_n1671__), .dout(new_new_n2294__));
  buf1  g1302(.din(new_new_n1669__), .dout(new_new_n2295__));
  buf1  g1303(.din(new_new_n1677__), .dout(new_new_n2296__));
  buf1  g1304(.din(new_new_n1339__), .dout(new_new_n2297__));
  buf1  g1305(.din(new_new_n1297__), .dout(new_new_n2298__));
  buf1  g1306(.din(new_new_n1247__), .dout(new_new_n2299__));
  buf1  g1307(.din(new_new_n1229__), .dout(new_new_n2300__));
  buf1  g1308(.din(new_new_n1680__), .dout(new_new_n2301__));
  buf1  g1309(.din(new_new_n1329__), .dout(new_new_n2302__));
  buf1  g1310(.din(new_new_n2302__), .dout(new_new_n2303__));
  buf1  g1311(.din(new_new_n961__), .dout(new_new_n2304__));
  buf1  g1312(.din(new_new_n995__), .dout(new_new_n2305__));
  buf1  g1313(.din(new_new_n1259__), .dout(new_new_n2306__));
  buf1  g1314(.din(new_new_n991__), .dout(new_new_n2307__));
  buf1  g1315(.din(new_new_n955__), .dout(new_new_n2308__));
  buf1  g1316(.din(new_new_n1753__), .dout(new_new_n2309__));
  buf1  g1317(.din(new_new_n1039__), .dout(new_new_n2310__));
  buf1  g1318(.din(new_new_n1694__), .dout(new_new_n2311__));
  buf1  g1319(.din(new_new_n1696__), .dout(new_new_n2312__));
  buf1  g1320(.din(new_new_n1702__), .dout(new_new_n2313__));
  buf1  g1321(.din(new_new_n1701__), .dout(new_new_n2314__));
  buf1  g1322(.din(new_new_n1743__), .dout(new_new_n2315__));
  buf1  g1323(.din(new_new_n1708__), .dout(new_new_n2316__));
  buf1  g1324(.din(new_new_n2316__), .dout(new_new_n2317__));
  buf1  g1325(.din(new_new_n971__), .dout(new_new_n2318__));
  buf1  g1326(.din(new_new_n1698__), .dout(new_new_n2319__));
  buf1  g1327(.din(new_new_n2319__), .dout(new_new_n2320__));
  buf1  g1328(.din(new_new_n1423__), .dout(new_new_n2321__));
  buf1  g1329(.din(new_new_n1710__), .dout(new_new_n2322__));
  buf1  g1330(.din(new_new_n2322__), .dout(new_new_n2323__));
  buf1  g1331(.din(new_new_n967__), .dout(new_new_n2324__));
  buf1  g1332(.din(new_new_n999__), .dout(new_new_n2325__));
  buf1  g1333(.din(new_new_n1766__), .dout(new_new_n2326__));
  buf1  g1334(.din(new_new_n1053__), .dout(new_new_n2327__));
  buf1  g1335(.din(new_new_n711__), .dout(new_new_n2328__));
  buf1  g1336(.din(new_new_n2328__), .dout(new_new_n2329__));
  buf1  g1337(.din(new_new_n2328__), .dout(new_new_n2330__));
  buf1  g1338(.din(new_new_n707__), .dout(new_new_n2331__));
  buf1  g1339(.din(new_new_n1772__), .dout(new_new_n2332__));
  buf1  g1340(.din(new_new_n725__), .dout(new_new_n2333__));
  buf1  g1341(.din(new_new_n719__), .dout(new_new_n2334__));
  buf1  g1342(.din(new_new_n2334__), .dout(new_new_n2335__));
  buf1  g1343(.din(new_new_n1771__), .dout(new_new_n2336__));
  buf1  g1344(.din(new_new_n737__), .dout(new_new_n2337__));
  buf1  g1345(.din(new_new_n715__), .dout(new_new_n2338__));
  always @ (posedge clock) begin
    n492_lo <= n3148;
    n495_lo <= n3151;
    n498_lo <= n3154;
    n501_lo <= n3157;
    n516_lo <= n3160;
    n528_lo <= n3163;
    n540_lo <= n3166;
    n543_lo <= n3169;
    n546_lo <= n3172;
    n549_lo <= n3175;
    n552_lo <= n3178;
    n564_lo <= n3181;
    n600_lo <= n3184;
    n603_lo <= n3187;
    n606_lo <= n3190;
    n609_lo <= n3193;
    n615_lo <= n3196;
    n618_lo <= n3199;
    n621_lo <= n3202;
    n627_lo <= n3205;
    n630_lo <= n3208;
    n633_lo <= n3211;
    n639_lo <= n3214;
    n642_lo <= n3217;
    n645_lo <= n3220;
    n648_lo <= n3223;
    n660_lo <= n3226;
    n672_lo <= n3229;
    n675_lo <= n3232;
    n678_lo <= n3235;
    n681_lo <= n3238;
    n684_lo <= n3241;
    n687_lo <= n3244;
    n690_lo <= n3247;
    n693_lo <= n3250;
    n696_lo <= n3253;
    n699_lo <= n3256;
    n702_lo <= n3259;
    n705_lo <= n3262;
    n708_lo <= n3265;
    n711_lo <= n3268;
    n714_lo <= n3271;
    n717_lo <= n3274;
    n720_lo <= n3277;
    n723_lo <= n3280;
    n726_lo <= n3283;
    n729_lo <= n3286;
    n732_lo <= n3289;
    n735_lo <= n3292;
    n738_lo <= n3295;
    n741_lo <= n3298;
    n744_lo <= n3301;
    n747_lo <= n3304;
    n750_lo <= n3307;
    n753_lo <= n3310;
    n756_lo <= n3313;
    n759_lo <= n3316;
    n762_lo <= n3319;
    n765_lo <= n3322;
    n768_lo <= n3325;
    n771_lo <= n3328;
    n774_lo <= n3331;
    n777_lo <= n3334;
    n780_lo <= n3337;
    n783_lo <= n3340;
    n786_lo <= n3343;
    n792_lo <= n3346;
    n795_lo <= n3349;
    n798_lo <= n3352;
    n807_lo <= n3355;
    n816_lo <= n3358;
    n819_lo <= n3361;
    n828_lo <= n3364;
    n831_lo <= n3367;
    n843_lo <= n3370;
    n846_lo <= n3373;
    n849_lo <= n3376;
    n852_lo <= n3379;
    n855_lo <= n3382;
    n858_lo <= n3385;
    n861_lo <= n3388;
    n864_lo <= n3391;
    n867_lo <= n3394;
    n870_lo <= n3397;
    n879_lo <= n3400;
    n882_lo <= n3403;
    n891_lo <= n3406;
    n903_lo <= n3409;
    n915_lo <= n3412;
    n918_lo <= n3415;
    n951_lo <= n3418;
    n954_lo <= n3421;
    n957_lo <= n3424;
    n960_lo <= n3427;
    n963_lo <= n3430;
    n966_lo <= n3433;
    n969_lo <= n3436;
    n972_lo <= n3439;
    n975_lo <= n3442;
    n978_lo <= n3445;
    n981_lo <= n3448;
    n984_lo <= n3451;
    n987_lo <= n3454;
    n990_lo <= n3457;
    n993_lo <= n3460;
    n996_lo <= n3463;
    n999_lo <= n3466;
    n1002_lo <= n3469;
    n1008_lo <= n3472;
    n1011_lo <= n3475;
    n1014_lo <= n3478;
    n1020_lo <= n3481;
    n1023_lo <= n3484;
    n1032_lo <= n3487;
    n1035_lo <= n3490;
    n1044_lo <= n3493;
    n1047_lo <= n3496;
    n1050_lo <= n3499;
    n1053_lo <= n3502;
    n1056_lo <= n3505;
    n1059_lo <= n3508;
    n1062_lo <= n3511;
    n1065_lo <= n3514;
    n1068_lo <= n3517;
    n1071_lo <= n3520;
    n1074_lo <= n3523;
    n1077_lo <= n3526;
    n1080_lo <= n3529;
    n1083_lo <= n3532;
    n1086_lo <= n3535;
    n1089_lo <= n3538;
    n1092_lo <= n3541;
    n1095_lo <= n3544;
    n1098_lo <= n3547;
    n1101_lo <= n3550;
    n1104_lo <= n3553;
    n1107_lo <= n3556;
    n1110_lo <= n3559;
    n1113_lo <= n3562;
    n1116_lo <= n3565;
    n1119_lo <= n3568;
    n1122_lo <= n3571;
    n1125_lo <= n3574;
    n1128_lo <= n3577;
    n1131_lo <= n3580;
    n1134_lo <= n3583;
    n1137_lo <= n3586;
    n1143_lo <= n3589;
    n1146_lo <= n3592;
    n1149_lo <= n3595;
    n1152_lo <= n3598;
    n1155_lo <= n3601;
    n1164_lo <= n3604;
    n1167_lo <= n3607;
    n1170_lo <= n3610;
    n1173_lo <= n3613;
    n1176_lo <= n3616;
    n1188_lo <= n3619;
    n563_inv <= n3622;
    n1429_o2 <= n3625;
    n1427_o2 <= n3628;
    n1471_o2 <= n3631;
    n1476_o2 <= n3634;
    n1499_o2 <= n3637;
    n1500_o2 <= n3640;
    n1501_o2 <= n3643;
    n1516_o2 <= n3646;
    n1517_o2 <= n3649;
    n1562_o2 <= n3652;
    n1563_o2 <= n3655;
    n1564_o2 <= n3658;
    n1582_o2 <= n3661;
    n1583_o2 <= n3664;
    n1618_o2 <= n3667;
    n1622_o2 <= n3670;
    n1502_o2 <= n3673;
    n1503_o2 <= n3676;
    n1504_o2 <= n3679;
    n1505_o2 <= n3682;
    n1506_o2 <= n3685;
    n1512_o2 <= n3688;
    n1513_o2 <= n3691;
    n1514_o2 <= n3694;
    n1515_o2 <= n3697;
    n1644_o2 <= n3700;
    n1647_o2 <= n3703;
    n1527_o2 <= n3706;
    n650_inv <= n3709;
    n653_inv <= n3712;
    n656_inv <= n3715;
    n1567_o2 <= n3718;
    n955_o2 <= n3721;
    n1568_o2 <= n3724;
    n1037_o2 <= n3727;
    n960_o2 <= n3730;
    n1587_o2 <= n3733;
    n1040_o2 <= n3736;
    n1039_o2 <= n3739;
    n1589_o2 <= n3742;
    n1624_o2 <= n3745;
    n1643_o2 <= n3748;
    n1038_o2 <= n3751;
    n1645_o2 <= n3754;
    n1029_o2 <= n3757;
    n701_inv <= n3760;
    n1662_o2 <= n3763;
    n1663_o2 <= n3766;
    n710_inv <= n3769;
    n813_o2 <= n3772;
    lo114_buf_o2 <= n3775;
    n1031_o2 <= n3778;
    lo186_buf_o2 <= n3781;
    n1042_o2 <= n3784;
    n728_inv <= n3787;
    n917_o2 <= n3790;
    n734_inv <= n3793;
    n1649_o2 <= n3796;
    n1650_o2 <= n3799;
    n1651_o2 <= n3802;
    n1652_o2 <= n3805;
    n1653_o2 <= n3808;
    lo138_buf_o2 <= n3811;
    n1664_o2 <= n3814;
    n1665_o2 <= n3817;
    n1666_o2 <= n3820;
    n1667_o2 <= n3823;
    n944_o2 <= n3826;
    n770_inv <= n3829;
    n1672_o2 <= n3832;
    n776_inv <= n3835;
    n1679_o2 <= n3838;
    n782_inv <= n3841;
    n785_inv <= n3844;
    lo110_buf_o2 <= n3847;
    lo134_buf_o2 <= n3850;
    n1030_o2 <= n3853;
    lo182_buf_o2 <= n3856;
    n830_o2 <= n3859;
    n1021_o2 <= n3862;
    n806_inv <= n3865;
    n809_inv <= n3868;
    n946_o2 <= n3871;
    lo038_buf_o2 <= n3874;
    lo238_buf_o2 <= n3877;
    n1010_o2 <= n3880;
    n1006_o2 <= n3883;
    n907_o2 <= n3886;
    n902_o2 <= n3889;
    lo154_buf_o2 <= n3892;
    n836_inv <= n3895;
    n839_inv <= n3898;
    lo122_buf_o2 <= n3901;
    n845_inv <= n3904;
    n904_o2 <= n3907;
    lo106_buf_o2 <= n3910;
    n980_o2 <= n3913;
    n1023_o2 <= n3916;
    lo178_buf_o2 <= n3919;
    n981_o2 <= n3922;
    n837_o2 <= n3925;
    n1013_o2 <= n3928;
    n840_o2 <= n3931;
    n849_o2 <= n3934;
    n852_o2 <= n3937;
    n864_o2 <= n3940;
    n867_o2 <= n3943;
    n1044_o2 <= n3946;
    n876_o2 <= n3949;
    n893_inv <= n3952;
    n879_o2 <= n3955;
    n925_o2 <= n3958;
    n902_inv <= n3961;
    lo146_buf_o2 <= n3964;
    n1026_o2 <= n3967;
    n1032_o2 <= n3970;
    lo118_buf_o2 <= n3973;
    n917_inv <= n3976;
    lo190_buf_o2 <= n3979;
    n1036_o2 <= n3982;
    n926_inv <= n3985;
    n929_inv <= n3988;
    lo002_buf_o2 <= n3991;
    lo014_buf_o2 <= n3994;
    lo030_buf_o2 <= n3997;
    lo034_buf_o2 <= n4000;
    lo042_buf_o2 <= n4003;
    lo113_buf_o2 <= n4006;
    lo185_buf_o2 <= n4009;
    n939_o2 <= n4012;
    n941_o2 <= n4015;
    lo142_buf_o2 <= n4018;
    lo230_buf_o2 <= n4021;
    lo006_buf_o2 <= n4024;
    lo018_buf_o2 <= n4027;
    lo022_buf_o2 <= n4030;
    lo066_buf_o2 <= n4033;
    n977_inv <= n4036;
    n826_o2 <= n4039;
    n892_o2 <= n4042;
    lo152_buf_o2 <= n4045;
    n896_o2 <= n4048;
    n905_o2 <= n4051;
    n995_inv <= n4054;
    lo037_buf_o2 <= n4057;
    lo237_buf_o2 <= n4060;
    lo062_buf_o2 <= n4063;
    n1007_inv <= n4066;
    n1010_inv <= n4069;
    n891_o2 <= n4072;
  end
  initial begin
    n492_lo <= 1'b0;
    n495_lo <= 1'b0;
    n498_lo <= 1'b0;
    n501_lo <= 1'b0;
    n516_lo <= 1'b0;
    n528_lo <= 1'b0;
    n540_lo <= 1'b0;
    n543_lo <= 1'b0;
    n546_lo <= 1'b0;
    n549_lo <= 1'b0;
    n552_lo <= 1'b0;
    n564_lo <= 1'b0;
    n600_lo <= 1'b0;
    n603_lo <= 1'b0;
    n606_lo <= 1'b0;
    n609_lo <= 1'b0;
    n615_lo <= 1'b0;
    n618_lo <= 1'b0;
    n621_lo <= 1'b0;
    n627_lo <= 1'b0;
    n630_lo <= 1'b0;
    n633_lo <= 1'b0;
    n639_lo <= 1'b0;
    n642_lo <= 1'b0;
    n645_lo <= 1'b0;
    n648_lo <= 1'b0;
    n660_lo <= 1'b0;
    n672_lo <= 1'b0;
    n675_lo <= 1'b0;
    n678_lo <= 1'b0;
    n681_lo <= 1'b0;
    n684_lo <= 1'b0;
    n687_lo <= 1'b0;
    n690_lo <= 1'b0;
    n693_lo <= 1'b0;
    n696_lo <= 1'b0;
    n699_lo <= 1'b0;
    n702_lo <= 1'b0;
    n705_lo <= 1'b0;
    n708_lo <= 1'b0;
    n711_lo <= 1'b0;
    n714_lo <= 1'b0;
    n717_lo <= 1'b0;
    n720_lo <= 1'b0;
    n723_lo <= 1'b0;
    n726_lo <= 1'b0;
    n729_lo <= 1'b0;
    n732_lo <= 1'b0;
    n735_lo <= 1'b0;
    n738_lo <= 1'b0;
    n741_lo <= 1'b0;
    n744_lo <= 1'b0;
    n747_lo <= 1'b0;
    n750_lo <= 1'b0;
    n753_lo <= 1'b0;
    n756_lo <= 1'b0;
    n759_lo <= 1'b0;
    n762_lo <= 1'b0;
    n765_lo <= 1'b0;
    n768_lo <= 1'b0;
    n771_lo <= 1'b0;
    n774_lo <= 1'b0;
    n777_lo <= 1'b0;
    n780_lo <= 1'b0;
    n783_lo <= 1'b0;
    n786_lo <= 1'b0;
    n792_lo <= 1'b0;
    n795_lo <= 1'b0;
    n798_lo <= 1'b0;
    n807_lo <= 1'b0;
    n816_lo <= 1'b0;
    n819_lo <= 1'b0;
    n828_lo <= 1'b0;
    n831_lo <= 1'b0;
    n843_lo <= 1'b0;
    n846_lo <= 1'b0;
    n849_lo <= 1'b0;
    n852_lo <= 1'b0;
    n855_lo <= 1'b0;
    n858_lo <= 1'b0;
    n861_lo <= 1'b0;
    n864_lo <= 1'b0;
    n867_lo <= 1'b0;
    n870_lo <= 1'b0;
    n879_lo <= 1'b0;
    n882_lo <= 1'b0;
    n891_lo <= 1'b0;
    n903_lo <= 1'b0;
    n915_lo <= 1'b0;
    n918_lo <= 1'b0;
    n951_lo <= 1'b0;
    n954_lo <= 1'b0;
    n957_lo <= 1'b0;
    n960_lo <= 1'b0;
    n963_lo <= 1'b0;
    n966_lo <= 1'b0;
    n969_lo <= 1'b0;
    n972_lo <= 1'b0;
    n975_lo <= 1'b0;
    n978_lo <= 1'b0;
    n981_lo <= 1'b0;
    n984_lo <= 1'b0;
    n987_lo <= 1'b0;
    n990_lo <= 1'b0;
    n993_lo <= 1'b0;
    n996_lo <= 1'b0;
    n999_lo <= 1'b0;
    n1002_lo <= 1'b0;
    n1008_lo <= 1'b0;
    n1011_lo <= 1'b0;
    n1014_lo <= 1'b0;
    n1020_lo <= 1'b0;
    n1023_lo <= 1'b0;
    n1032_lo <= 1'b0;
    n1035_lo <= 1'b0;
    n1044_lo <= 1'b0;
    n1047_lo <= 1'b0;
    n1050_lo <= 1'b0;
    n1053_lo <= 1'b0;
    n1056_lo <= 1'b0;
    n1059_lo <= 1'b0;
    n1062_lo <= 1'b0;
    n1065_lo <= 1'b0;
    n1068_lo <= 1'b0;
    n1071_lo <= 1'b0;
    n1074_lo <= 1'b0;
    n1077_lo <= 1'b0;
    n1080_lo <= 1'b0;
    n1083_lo <= 1'b0;
    n1086_lo <= 1'b0;
    n1089_lo <= 1'b0;
    n1092_lo <= 1'b0;
    n1095_lo <= 1'b0;
    n1098_lo <= 1'b0;
    n1101_lo <= 1'b0;
    n1104_lo <= 1'b0;
    n1107_lo <= 1'b0;
    n1110_lo <= 1'b0;
    n1113_lo <= 1'b0;
    n1116_lo <= 1'b0;
    n1119_lo <= 1'b0;
    n1122_lo <= 1'b0;
    n1125_lo <= 1'b0;
    n1128_lo <= 1'b0;
    n1131_lo <= 1'b0;
    n1134_lo <= 1'b0;
    n1137_lo <= 1'b0;
    n1143_lo <= 1'b0;
    n1146_lo <= 1'b0;
    n1149_lo <= 1'b0;
    n1152_lo <= 1'b0;
    n1155_lo <= 1'b0;
    n1164_lo <= 1'b0;
    n1167_lo <= 1'b0;
    n1170_lo <= 1'b0;
    n1173_lo <= 1'b0;
    n1176_lo <= 1'b0;
    n1188_lo <= 1'b0;
    n563_inv <= 1'b0;
    n1429_o2 <= 1'b0;
    n1427_o2 <= 1'b0;
    n1471_o2 <= 1'b0;
    n1476_o2 <= 1'b0;
    n1499_o2 <= 1'b0;
    n1500_o2 <= 1'b0;
    n1501_o2 <= 1'b0;
    n1516_o2 <= 1'b0;
    n1517_o2 <= 1'b0;
    n1562_o2 <= 1'b0;
    n1563_o2 <= 1'b0;
    n1564_o2 <= 1'b0;
    n1582_o2 <= 1'b0;
    n1583_o2 <= 1'b0;
    n1618_o2 <= 1'b0;
    n1622_o2 <= 1'b0;
    n1502_o2 <= 1'b0;
    n1503_o2 <= 1'b0;
    n1504_o2 <= 1'b0;
    n1505_o2 <= 1'b0;
    n1506_o2 <= 1'b0;
    n1512_o2 <= 1'b0;
    n1513_o2 <= 1'b0;
    n1514_o2 <= 1'b0;
    n1515_o2 <= 1'b0;
    n1644_o2 <= 1'b0;
    n1647_o2 <= 1'b0;
    n1527_o2 <= 1'b0;
    n650_inv <= 1'b0;
    n653_inv <= 1'b0;
    n656_inv <= 1'b0;
    n1567_o2 <= 1'b0;
    n955_o2 <= 1'b0;
    n1568_o2 <= 1'b0;
    n1037_o2 <= 1'b0;
    n960_o2 <= 1'b0;
    n1587_o2 <= 1'b0;
    n1040_o2 <= 1'b0;
    n1039_o2 <= 1'b0;
    n1589_o2 <= 1'b0;
    n1624_o2 <= 1'b0;
    n1643_o2 <= 1'b0;
    n1038_o2 <= 1'b0;
    n1645_o2 <= 1'b0;
    n1029_o2 <= 1'b0;
    n701_inv <= 1'b0;
    n1662_o2 <= 1'b0;
    n1663_o2 <= 1'b0;
    n710_inv <= 1'b0;
    n813_o2 <= 1'b0;
    lo114_buf_o2 <= 1'b0;
    n1031_o2 <= 1'b0;
    lo186_buf_o2 <= 1'b0;
    n1042_o2 <= 1'b0;
    n728_inv <= 1'b0;
    n917_o2 <= 1'b0;
    n734_inv <= 1'b0;
    n1649_o2 <= 1'b0;
    n1650_o2 <= 1'b0;
    n1651_o2 <= 1'b0;
    n1652_o2 <= 1'b0;
    n1653_o2 <= 1'b0;
    lo138_buf_o2 <= 1'b0;
    n1664_o2 <= 1'b0;
    n1665_o2 <= 1'b0;
    n1666_o2 <= 1'b0;
    n1667_o2 <= 1'b0;
    n944_o2 <= 1'b0;
    n770_inv <= 1'b0;
    n1672_o2 <= 1'b0;
    n776_inv <= 1'b0;
    n1679_o2 <= 1'b0;
    n782_inv <= 1'b0;
    n785_inv <= 1'b0;
    lo110_buf_o2 <= 1'b0;
    lo134_buf_o2 <= 1'b0;
    n1030_o2 <= 1'b0;
    lo182_buf_o2 <= 1'b0;
    n830_o2 <= 1'b0;
    n1021_o2 <= 1'b0;
    n806_inv <= 1'b0;
    n809_inv <= 1'b0;
    n946_o2 <= 1'b0;
    lo038_buf_o2 <= 1'b0;
    lo238_buf_o2 <= 1'b0;
    n1010_o2 <= 1'b0;
    n1006_o2 <= 1'b0;
    n907_o2 <= 1'b0;
    n902_o2 <= 1'b0;
    lo154_buf_o2 <= 1'b0;
    n836_inv <= 1'b0;
    n839_inv <= 1'b0;
    lo122_buf_o2 <= 1'b0;
    n845_inv <= 1'b0;
    n904_o2 <= 1'b0;
    lo106_buf_o2 <= 1'b0;
    n980_o2 <= 1'b0;
    n1023_o2 <= 1'b0;
    lo178_buf_o2 <= 1'b0;
    n981_o2 <= 1'b0;
    n837_o2 <= 1'b0;
    n1013_o2 <= 1'b0;
    n840_o2 <= 1'b0;
    n849_o2 <= 1'b0;
    n852_o2 <= 1'b0;
    n864_o2 <= 1'b0;
    n867_o2 <= 1'b0;
    n1044_o2 <= 1'b0;
    n876_o2 <= 1'b0;
    n893_inv <= 1'b0;
    n879_o2 <= 1'b0;
    n925_o2 <= 1'b0;
    n902_inv <= 1'b0;
    lo146_buf_o2 <= 1'b0;
    n1026_o2 <= 1'b0;
    n1032_o2 <= 1'b0;
    lo118_buf_o2 <= 1'b0;
    n917_inv <= 1'b0;
    lo190_buf_o2 <= 1'b0;
    n1036_o2 <= 1'b0;
    n926_inv <= 1'b0;
    n929_inv <= 1'b0;
    lo002_buf_o2 <= 1'b0;
    lo014_buf_o2 <= 1'b0;
    lo030_buf_o2 <= 1'b0;
    lo034_buf_o2 <= 1'b0;
    lo042_buf_o2 <= 1'b0;
    lo113_buf_o2 <= 1'b0;
    lo185_buf_o2 <= 1'b0;
    n939_o2 <= 1'b0;
    n941_o2 <= 1'b0;
    lo142_buf_o2 <= 1'b0;
    lo230_buf_o2 <= 1'b0;
    lo006_buf_o2 <= 1'b0;
    lo018_buf_o2 <= 1'b0;
    lo022_buf_o2 <= 1'b0;
    lo066_buf_o2 <= 1'b0;
    n977_inv <= 1'b0;
    n826_o2 <= 1'b0;
    n892_o2 <= 1'b0;
    lo152_buf_o2 <= 1'b0;
    n896_o2 <= 1'b0;
    n905_o2 <= 1'b0;
    n995_inv <= 1'b0;
    lo037_buf_o2 <= 1'b0;
    lo237_buf_o2 <= 1'b0;
    lo062_buf_o2 <= 1'b0;
    n1007_inv <= 1'b0;
    n1010_inv <= 1'b0;
    n891_o2 <= 1'b0;
  end
endmodule


