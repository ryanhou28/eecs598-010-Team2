// Benchmark "c499" written by ABC on Sun Oct 29 22:18:03 2023

module c499 ( 
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41,
    G468, G469, G470, G471, G472, G473, G474, G475, G476, G477, G478, G479,
    G480, G481, G482, G483, G484, G485, G486, G487, G488, G489, G490, G491,
    G492, G493, G494, G495, G496, G497, G498, G499  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41;
  output G468, G469, G470, G471, G472, G473, G474, G475, G476, G477, G478,
    G479, G480, G481, G482, G483, G484, G485, G486, G487, G488, G489, G490,
    G491, G492, G493, G494, G495, G496, G497, G498, G499;
  wire new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_,
    new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n318_,
    new_n319_, new_n320_, new_n322_, new_n323_, new_n324_, new_n326_,
    new_n327_, new_n328_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n337_, new_n338_, new_n339_, new_n341_,
    new_n342_, new_n343_, new_n345_, new_n346_, new_n347_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n355_, new_n356_,
    new_n357_, new_n359_, new_n360_, new_n361_, new_n363_, new_n364_,
    new_n365_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n373_, new_n374_, new_n375_, new_n377_, new_n378_, new_n379_,
    new_n381_, new_n382_, new_n383_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n398_, new_n399_, new_n400_,
    new_n402_, new_n403_, new_n404_, new_n406_, new_n407_, new_n408_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n416_,
    new_n417_, new_n418_, new_n420_, new_n421_, new_n422_, new_n424_,
    new_n425_, new_n426_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n434_, new_n435_, new_n436_, new_n438_, new_n439_,
    new_n440_, new_n442_, new_n443_, new_n444_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n451_, new_n452_, new_n453_, new_n455_,
    new_n456_, new_n457_, new_n459_, new_n460_, new_n461_;
  anb1 g000(.dina(G1), .dinb(G5), .dout(new_n74_));
  anb2 g001(.dina(G1), .dinb(G5), .dout(new_n75_));
  anb2 g002(.dina(new_n74_), .dinb(new_n75_), .dout(new_n76_));
  anb1 g003(.dina(G9), .dinb(G13), .dout(new_n77_));
  anb2 g004(.dina(G9), .dinb(G13), .dout(new_n78_));
  anb2 g005(.dina(new_n77_), .dinb(new_n78_), .dout(new_n79_));
  anb2 g006(.dina(new_n76_), .dinb(new_n79_), .dout(new_n80_));
  anb1 g007(.dina(new_n76_), .dinb(new_n79_), .dout(new_n81_));
  anb1 g008(.dina(new_n80_), .dinb(new_n81_), .dout(new_n82_));
  and1 g009(.dina(G33), .dinb(G41), .dout(new_n83_));
  anb1 g010(.dina(G17), .dinb(G18), .dout(new_n84_));
  anb2 g011(.dina(G17), .dinb(G18), .dout(new_n85_));
  anb2 g012(.dina(new_n84_), .dinb(new_n85_), .dout(new_n86_));
  anb1 g013(.dina(G19), .dinb(G20), .dout(new_n87_));
  anb2 g014(.dina(G19), .dinb(G20), .dout(new_n88_));
  anb2 g015(.dina(new_n87_), .dinb(new_n88_), .dout(new_n89_));
  anb2 g016(.dina(new_n86_), .dinb(new_n89_), .dout(new_n90_));
  anb1 g017(.dina(new_n86_), .dinb(new_n89_), .dout(new_n91_));
  anb1 g018(.dina(new_n90_), .dinb(new_n91_), .dout(new_n92_));
  anb1 g019(.dina(G21), .dinb(G22), .dout(new_n93_));
  anb2 g020(.dina(G21), .dinb(G22), .dout(new_n94_));
  anb2 g021(.dina(new_n93_), .dinb(new_n94_), .dout(new_n95_));
  anb1 g022(.dina(G23), .dinb(G24), .dout(new_n96_));
  anb2 g023(.dina(G23), .dinb(G24), .dout(new_n97_));
  anb2 g024(.dina(new_n96_), .dinb(new_n97_), .dout(new_n98_));
  anb2 g025(.dina(new_n95_), .dinb(new_n98_), .dout(new_n99_));
  anb1 g026(.dina(new_n95_), .dinb(new_n98_), .dout(new_n100_));
  anb1 g027(.dina(new_n99_), .dinb(new_n100_), .dout(new_n101_));
  anb1 g028(.dina(new_n92_), .dinb(new_n101_), .dout(new_n102_));
  anb2 g029(.dina(new_n92_), .dinb(new_n101_), .dout(new_n103_));
  anb2 g030(.dina(new_n102_), .dinb(new_n103_), .dout(new_n104_));
  anb2 g031(.dina(new_n83_), .dinb(new_n104_), .dout(new_n105_));
  anb1 g032(.dina(new_n83_), .dinb(new_n104_), .dout(new_n106_));
  anb1 g033(.dina(new_n105_), .dinb(new_n106_), .dout(new_n107_));
  anb1 g034(.dina(new_n82_), .dinb(new_n107_), .dout(new_n108_));
  anb2 g035(.dina(new_n82_), .dinb(new_n107_), .dout(new_n109_));
  anb2 g036(.dina(new_n108_), .dinb(new_n109_), .dout(new_n110_));
  anb1 g037(.dina(G17), .dinb(G21), .dout(new_n111_));
  anb2 g038(.dina(G17), .dinb(G21), .dout(new_n112_));
  anb2 g039(.dina(new_n111_), .dinb(new_n112_), .dout(new_n113_));
  anb1 g040(.dina(G25), .dinb(G29), .dout(new_n114_));
  anb2 g041(.dina(G25), .dinb(G29), .dout(new_n115_));
  anb2 g042(.dina(new_n114_), .dinb(new_n115_), .dout(new_n116_));
  anb2 g043(.dina(new_n113_), .dinb(new_n116_), .dout(new_n117_));
  anb1 g044(.dina(new_n113_), .dinb(new_n116_), .dout(new_n118_));
  anb1 g045(.dina(new_n117_), .dinb(new_n118_), .dout(new_n119_));
  and1 g046(.dina(G37), .dinb(G41), .dout(new_n120_));
  anb1 g047(.dina(G5), .dinb(G6), .dout(new_n121_));
  anb2 g048(.dina(G5), .dinb(G6), .dout(new_n122_));
  anb2 g049(.dina(new_n121_), .dinb(new_n122_), .dout(new_n123_));
  anb1 g050(.dina(G7), .dinb(G8), .dout(new_n124_));
  anb2 g051(.dina(G7), .dinb(G8), .dout(new_n125_));
  anb2 g052(.dina(new_n124_), .dinb(new_n125_), .dout(new_n126_));
  anb2 g053(.dina(new_n123_), .dinb(new_n126_), .dout(new_n127_));
  anb1 g054(.dina(new_n123_), .dinb(new_n126_), .dout(new_n128_));
  anb1 g055(.dina(new_n127_), .dinb(new_n128_), .dout(new_n129_));
  anb1 g056(.dina(G1), .dinb(G2), .dout(new_n130_));
  anb2 g057(.dina(G1), .dinb(G2), .dout(new_n131_));
  anb2 g058(.dina(new_n130_), .dinb(new_n131_), .dout(new_n132_));
  anb1 g059(.dina(G3), .dinb(G4), .dout(new_n133_));
  anb2 g060(.dina(G3), .dinb(G4), .dout(new_n134_));
  anb2 g061(.dina(new_n133_), .dinb(new_n134_), .dout(new_n135_));
  anb2 g062(.dina(new_n132_), .dinb(new_n135_), .dout(new_n136_));
  anb1 g063(.dina(new_n132_), .dinb(new_n135_), .dout(new_n137_));
  anb1 g064(.dina(new_n136_), .dinb(new_n137_), .dout(new_n138_));
  anb1 g065(.dina(new_n129_), .dinb(new_n138_), .dout(new_n139_));
  anb2 g066(.dina(new_n129_), .dinb(new_n138_), .dout(new_n140_));
  anb2 g067(.dina(new_n139_), .dinb(new_n140_), .dout(new_n141_));
  anb2 g068(.dina(new_n120_), .dinb(new_n141_), .dout(new_n142_));
  anb1 g069(.dina(new_n120_), .dinb(new_n141_), .dout(new_n143_));
  anb1 g070(.dina(new_n142_), .dinb(new_n143_), .dout(new_n144_));
  anb1 g071(.dina(new_n119_), .dinb(new_n144_), .dout(new_n145_));
  anb2 g072(.dina(new_n119_), .dinb(new_n144_), .dout(new_n146_));
  anb2 g073(.dina(new_n145_), .dinb(new_n146_), .dout(new_n147_));
  anb1 g074(.dina(G18), .dinb(G22), .dout(new_n148_));
  anb2 g075(.dina(G18), .dinb(G22), .dout(new_n149_));
  anb2 g076(.dina(new_n148_), .dinb(new_n149_), .dout(new_n150_));
  anb1 g077(.dina(G26), .dinb(G30), .dout(new_n151_));
  anb2 g078(.dina(G26), .dinb(G30), .dout(new_n152_));
  anb2 g079(.dina(new_n151_), .dinb(new_n152_), .dout(new_n153_));
  anb2 g080(.dina(new_n150_), .dinb(new_n153_), .dout(new_n154_));
  anb1 g081(.dina(new_n150_), .dinb(new_n153_), .dout(new_n155_));
  anb1 g082(.dina(new_n154_), .dinb(new_n155_), .dout(new_n156_));
  and1 g083(.dina(G38), .dinb(G41), .dout(new_n157_));
  anb1 g084(.dina(G13), .dinb(G14), .dout(new_n158_));
  anb2 g085(.dina(G13), .dinb(G14), .dout(new_n159_));
  anb2 g086(.dina(new_n158_), .dinb(new_n159_), .dout(new_n160_));
  anb1 g087(.dina(G15), .dinb(G16), .dout(new_n161_));
  anb2 g088(.dina(G15), .dinb(G16), .dout(new_n162_));
  anb2 g089(.dina(new_n161_), .dinb(new_n162_), .dout(new_n163_));
  anb2 g090(.dina(new_n160_), .dinb(new_n163_), .dout(new_n164_));
  anb1 g091(.dina(new_n160_), .dinb(new_n163_), .dout(new_n165_));
  anb1 g092(.dina(new_n164_), .dinb(new_n165_), .dout(new_n166_));
  anb1 g093(.dina(G9), .dinb(G10), .dout(new_n167_));
  anb2 g094(.dina(G9), .dinb(G10), .dout(new_n168_));
  anb2 g095(.dina(new_n167_), .dinb(new_n168_), .dout(new_n169_));
  anb1 g096(.dina(G11), .dinb(G12), .dout(new_n170_));
  anb2 g097(.dina(G11), .dinb(G12), .dout(new_n171_));
  anb2 g098(.dina(new_n170_), .dinb(new_n171_), .dout(new_n172_));
  anb2 g099(.dina(new_n169_), .dinb(new_n172_), .dout(new_n173_));
  anb1 g100(.dina(new_n169_), .dinb(new_n172_), .dout(new_n174_));
  anb1 g101(.dina(new_n173_), .dinb(new_n174_), .dout(new_n175_));
  anb1 g102(.dina(new_n166_), .dinb(new_n175_), .dout(new_n176_));
  anb2 g103(.dina(new_n166_), .dinb(new_n175_), .dout(new_n177_));
  anb2 g104(.dina(new_n176_), .dinb(new_n177_), .dout(new_n178_));
  anb2 g105(.dina(new_n157_), .dinb(new_n178_), .dout(new_n179_));
  anb1 g106(.dina(new_n157_), .dinb(new_n178_), .dout(new_n180_));
  anb1 g107(.dina(new_n179_), .dinb(new_n180_), .dout(new_n181_));
  anb1 g108(.dina(new_n156_), .dinb(new_n181_), .dout(new_n182_));
  anb2 g109(.dina(new_n156_), .dinb(new_n181_), .dout(new_n183_));
  anb2 g110(.dina(new_n182_), .dinb(new_n183_), .dout(new_n184_));
  anb2 g111(.dina(new_n184_), .dinb(new_n147_), .dout(new_n185_));
  anb1 g112(.dina(G20), .dinb(G24), .dout(new_n186_));
  anb2 g113(.dina(G20), .dinb(G24), .dout(new_n187_));
  anb2 g114(.dina(new_n186_), .dinb(new_n187_), .dout(new_n188_));
  anb1 g115(.dina(G28), .dinb(G32), .dout(new_n189_));
  anb2 g116(.dina(G28), .dinb(G32), .dout(new_n190_));
  anb2 g117(.dina(new_n189_), .dinb(new_n190_), .dout(new_n191_));
  anb2 g118(.dina(new_n188_), .dinb(new_n191_), .dout(new_n192_));
  anb1 g119(.dina(new_n188_), .dinb(new_n191_), .dout(new_n193_));
  anb1 g120(.dina(new_n192_), .dinb(new_n193_), .dout(new_n194_));
  and1 g121(.dina(G40), .dinb(G41), .dout(new_n195_));
  anb1 g122(.dina(new_n129_), .dinb(new_n166_), .dout(new_n196_));
  anb2 g123(.dina(new_n129_), .dinb(new_n166_), .dout(new_n197_));
  anb2 g124(.dina(new_n196_), .dinb(new_n197_), .dout(new_n198_));
  anb2 g125(.dina(new_n195_), .dinb(new_n198_), .dout(new_n199_));
  anb1 g126(.dina(new_n195_), .dinb(new_n198_), .dout(new_n200_));
  anb1 g127(.dina(new_n199_), .dinb(new_n200_), .dout(new_n201_));
  anb1 g128(.dina(new_n194_), .dinb(new_n201_), .dout(new_n202_));
  anb2 g129(.dina(new_n194_), .dinb(new_n201_), .dout(new_n203_));
  anb2 g130(.dina(new_n202_), .dinb(new_n203_), .dout(new_n204_));
  anb1 g131(.dina(G19), .dinb(G23), .dout(new_n205_));
  anb2 g132(.dina(G19), .dinb(G23), .dout(new_n206_));
  anb2 g133(.dina(new_n205_), .dinb(new_n206_), .dout(new_n207_));
  anb1 g134(.dina(G27), .dinb(G31), .dout(new_n208_));
  anb2 g135(.dina(G27), .dinb(G31), .dout(new_n209_));
  anb2 g136(.dina(new_n208_), .dinb(new_n209_), .dout(new_n210_));
  anb2 g137(.dina(new_n207_), .dinb(new_n210_), .dout(new_n211_));
  anb1 g138(.dina(new_n207_), .dinb(new_n210_), .dout(new_n212_));
  anb1 g139(.dina(new_n211_), .dinb(new_n212_), .dout(new_n213_));
  and1 g140(.dina(G39), .dinb(G41), .dout(new_n214_));
  anb1 g141(.dina(new_n138_), .dinb(new_n175_), .dout(new_n215_));
  anb2 g142(.dina(new_n138_), .dinb(new_n175_), .dout(new_n216_));
  anb2 g143(.dina(new_n215_), .dinb(new_n216_), .dout(new_n217_));
  anb2 g144(.dina(new_n214_), .dinb(new_n217_), .dout(new_n218_));
  anb1 g145(.dina(new_n214_), .dinb(new_n217_), .dout(new_n219_));
  anb1 g146(.dina(new_n218_), .dinb(new_n219_), .dout(new_n220_));
  anb1 g147(.dina(new_n213_), .dinb(new_n220_), .dout(new_n221_));
  anb2 g148(.dina(new_n213_), .dinb(new_n220_), .dout(new_n222_));
  anb2 g149(.dina(new_n221_), .dinb(new_n222_), .dout(new_n223_));
  anb1 g150(.dina(new_n223_), .dinb(new_n204_), .dout(new_n224_));
  anb1 g151(.dina(G4), .dinb(G8), .dout(new_n225_));
  anb2 g152(.dina(G4), .dinb(G8), .dout(new_n226_));
  anb2 g153(.dina(new_n225_), .dinb(new_n226_), .dout(new_n227_));
  anb1 g154(.dina(G12), .dinb(G16), .dout(new_n228_));
  anb2 g155(.dina(G12), .dinb(G16), .dout(new_n229_));
  anb2 g156(.dina(new_n228_), .dinb(new_n229_), .dout(new_n230_));
  anb2 g157(.dina(new_n227_), .dinb(new_n230_), .dout(new_n231_));
  anb1 g158(.dina(new_n227_), .dinb(new_n230_), .dout(new_n232_));
  anb1 g159(.dina(new_n231_), .dinb(new_n232_), .dout(new_n233_));
  and1 g160(.dina(G36), .dinb(G41), .dout(new_n234_));
  anb1 g161(.dina(G29), .dinb(G30), .dout(new_n235_));
  anb2 g162(.dina(G29), .dinb(G30), .dout(new_n236_));
  anb2 g163(.dina(new_n235_), .dinb(new_n236_), .dout(new_n237_));
  anb1 g164(.dina(G31), .dinb(G32), .dout(new_n238_));
  anb2 g165(.dina(G31), .dinb(G32), .dout(new_n239_));
  anb2 g166(.dina(new_n238_), .dinb(new_n239_), .dout(new_n240_));
  anb2 g167(.dina(new_n237_), .dinb(new_n240_), .dout(new_n241_));
  anb1 g168(.dina(new_n237_), .dinb(new_n240_), .dout(new_n242_));
  anb1 g169(.dina(new_n241_), .dinb(new_n242_), .dout(new_n243_));
  anb1 g170(.dina(new_n101_), .dinb(new_n243_), .dout(new_n244_));
  anb2 g171(.dina(new_n101_), .dinb(new_n243_), .dout(new_n245_));
  anb2 g172(.dina(new_n244_), .dinb(new_n245_), .dout(new_n246_));
  anb2 g173(.dina(new_n234_), .dinb(new_n246_), .dout(new_n247_));
  anb1 g174(.dina(new_n234_), .dinb(new_n246_), .dout(new_n248_));
  anb1 g175(.dina(new_n247_), .dinb(new_n248_), .dout(new_n249_));
  anb1 g176(.dina(new_n233_), .dinb(new_n249_), .dout(new_n250_));
  anb2 g177(.dina(new_n233_), .dinb(new_n249_), .dout(new_n251_));
  anb2 g178(.dina(new_n250_), .dinb(new_n251_), .dout(new_n252_));
  anb1 g179(.dina(G3), .dinb(G7), .dout(new_n253_));
  anb2 g180(.dina(G3), .dinb(G7), .dout(new_n254_));
  anb2 g181(.dina(new_n253_), .dinb(new_n254_), .dout(new_n255_));
  anb1 g182(.dina(G11), .dinb(G15), .dout(new_n256_));
  anb2 g183(.dina(G11), .dinb(G15), .dout(new_n257_));
  anb2 g184(.dina(new_n256_), .dinb(new_n257_), .dout(new_n258_));
  anb2 g185(.dina(new_n255_), .dinb(new_n258_), .dout(new_n259_));
  anb1 g186(.dina(new_n255_), .dinb(new_n258_), .dout(new_n260_));
  anb1 g187(.dina(new_n259_), .dinb(new_n260_), .dout(new_n261_));
  and1 g188(.dina(G35), .dinb(G41), .dout(new_n262_));
  anb1 g189(.dina(G25), .dinb(G26), .dout(new_n263_));
  anb2 g190(.dina(G25), .dinb(G26), .dout(new_n264_));
  anb2 g191(.dina(new_n263_), .dinb(new_n264_), .dout(new_n265_));
  anb1 g192(.dina(G27), .dinb(G28), .dout(new_n266_));
  anb2 g193(.dina(G27), .dinb(G28), .dout(new_n267_));
  anb2 g194(.dina(new_n266_), .dinb(new_n267_), .dout(new_n268_));
  anb2 g195(.dina(new_n265_), .dinb(new_n268_), .dout(new_n269_));
  anb1 g196(.dina(new_n265_), .dinb(new_n268_), .dout(new_n270_));
  anb1 g197(.dina(new_n269_), .dinb(new_n270_), .dout(new_n271_));
  anb1 g198(.dina(new_n92_), .dinb(new_n271_), .dout(new_n272_));
  anb2 g199(.dina(new_n92_), .dinb(new_n271_), .dout(new_n273_));
  anb2 g200(.dina(new_n272_), .dinb(new_n273_), .dout(new_n274_));
  anb2 g201(.dina(new_n262_), .dinb(new_n274_), .dout(new_n275_));
  anb1 g202(.dina(new_n262_), .dinb(new_n274_), .dout(new_n276_));
  anb1 g203(.dina(new_n275_), .dinb(new_n276_), .dout(new_n277_));
  anb1 g204(.dina(new_n261_), .dinb(new_n277_), .dout(new_n278_));
  anb2 g205(.dina(new_n261_), .dinb(new_n277_), .dout(new_n279_));
  anb2 g206(.dina(new_n278_), .dinb(new_n279_), .dout(new_n280_));
  anb1 g207(.dina(G2), .dinb(G6), .dout(new_n281_));
  anb2 g208(.dina(G2), .dinb(G6), .dout(new_n282_));
  anb2 g209(.dina(new_n281_), .dinb(new_n282_), .dout(new_n283_));
  anb1 g210(.dina(G10), .dinb(G14), .dout(new_n284_));
  anb2 g211(.dina(G10), .dinb(G14), .dout(new_n285_));
  anb2 g212(.dina(new_n284_), .dinb(new_n285_), .dout(new_n286_));
  anb2 g213(.dina(new_n283_), .dinb(new_n286_), .dout(new_n287_));
  anb1 g214(.dina(new_n283_), .dinb(new_n286_), .dout(new_n288_));
  anb1 g215(.dina(new_n287_), .dinb(new_n288_), .dout(new_n289_));
  and1 g216(.dina(G34), .dinb(G41), .dout(new_n290_));
  anb1 g217(.dina(new_n243_), .dinb(new_n271_), .dout(new_n291_));
  anb2 g218(.dina(new_n243_), .dinb(new_n271_), .dout(new_n292_));
  anb2 g219(.dina(new_n291_), .dinb(new_n292_), .dout(new_n293_));
  anb2 g220(.dina(new_n290_), .dinb(new_n293_), .dout(new_n294_));
  anb1 g221(.dina(new_n290_), .dinb(new_n293_), .dout(new_n295_));
  anb1 g222(.dina(new_n294_), .dinb(new_n295_), .dout(new_n296_));
  anb1 g223(.dina(new_n289_), .dinb(new_n296_), .dout(new_n297_));
  anb2 g224(.dina(new_n289_), .dinb(new_n296_), .dout(new_n298_));
  anb2 g225(.dina(new_n297_), .dinb(new_n298_), .dout(new_n299_));
  anb1 g226(.dina(new_n110_), .dinb(new_n299_), .dout(new_n300_));
  anb2 g227(.dina(new_n280_), .dinb(new_n300_), .dout(new_n301_));
  anb1 g228(.dina(new_n299_), .dinb(new_n110_), .dout(new_n302_));
  anb2 g229(.dina(new_n280_), .dinb(new_n302_), .dout(new_n303_));
  nor2 g230(.dina(new_n301_), .dinb(new_n303_), .dout(new_n304_));
  anb2 g231(.dina(new_n252_), .dinb(new_n304_), .dout(new_n305_));
  anb2 g232(.dina(new_n252_), .dinb(new_n280_), .dout(new_n306_));
  anb1 g233(.dina(new_n252_), .dinb(new_n280_), .dout(new_n307_));
  nab2 g234(.dina(new_n306_), .dinb(new_n307_), .dout(new_n308_));
  and2 g235(.dina(new_n110_), .dinb(new_n299_), .dout(new_n309_));
  anb1 g236(.dina(new_n308_), .dinb(new_n309_), .dout(new_n310_));
  anb1 g237(.dina(new_n305_), .dinb(new_n310_), .dout(new_n311_));
  anb1 g238(.dina(new_n224_), .dinb(new_n311_), .dout(new_n312_));
  anb2 g239(.dina(new_n185_), .dinb(new_n312_), .dout(new_n313_));
  anb1 g240(.dina(new_n110_), .dinb(new_n313_), .dout(new_n314_));
  anb1 g241(.dina(new_n314_), .dinb(G1), .dout(new_n315_));
  anb2 g242(.dina(new_n314_), .dinb(G1), .dout(new_n316_));
  anb2 g243(.dina(new_n315_), .dinb(new_n316_), .dout(G468));
  anb1 g244(.dina(new_n299_), .dinb(new_n313_), .dout(new_n318_));
  anb1 g245(.dina(new_n318_), .dinb(G2), .dout(new_n319_));
  anb2 g246(.dina(new_n318_), .dinb(G2), .dout(new_n320_));
  anb2 g247(.dina(new_n319_), .dinb(new_n320_), .dout(G469));
  anb1 g248(.dina(new_n280_), .dinb(new_n313_), .dout(new_n322_));
  anb1 g249(.dina(new_n322_), .dinb(G3), .dout(new_n323_));
  anb2 g250(.dina(new_n322_), .dinb(G3), .dout(new_n324_));
  anb2 g251(.dina(new_n323_), .dinb(new_n324_), .dout(G470));
  anb1 g252(.dina(new_n252_), .dinb(new_n313_), .dout(new_n326_));
  anb1 g253(.dina(new_n326_), .dinb(G4), .dout(new_n327_));
  anb2 g254(.dina(new_n326_), .dinb(G4), .dout(new_n328_));
  anb2 g255(.dina(new_n327_), .dinb(new_n328_), .dout(G471));
  and2 g256(.dina(new_n185_), .dinb(new_n223_), .dout(new_n330_));
  anb1 g257(.dina(new_n204_), .dinb(new_n311_), .dout(new_n331_));
  anb2 g258(.dina(new_n330_), .dinb(new_n331_), .dout(new_n332_));
  anb1 g259(.dina(new_n110_), .dinb(new_n332_), .dout(new_n333_));
  anb1 g260(.dina(new_n333_), .dinb(G5), .dout(new_n334_));
  anb2 g261(.dina(new_n333_), .dinb(G5), .dout(new_n335_));
  anb2 g262(.dina(new_n334_), .dinb(new_n335_), .dout(G472));
  anb1 g263(.dina(new_n299_), .dinb(new_n332_), .dout(new_n337_));
  anb1 g264(.dina(new_n337_), .dinb(G6), .dout(new_n338_));
  anb2 g265(.dina(new_n337_), .dinb(G6), .dout(new_n339_));
  anb2 g266(.dina(new_n338_), .dinb(new_n339_), .dout(G473));
  anb1 g267(.dina(new_n280_), .dinb(new_n332_), .dout(new_n341_));
  anb1 g268(.dina(new_n341_), .dinb(G7), .dout(new_n342_));
  anb2 g269(.dina(new_n341_), .dinb(G7), .dout(new_n343_));
  anb2 g270(.dina(new_n342_), .dinb(new_n343_), .dout(G474));
  anb1 g271(.dina(new_n252_), .dinb(new_n332_), .dout(new_n345_));
  anb1 g272(.dina(new_n345_), .dinb(G8), .dout(new_n346_));
  anb2 g273(.dina(new_n345_), .dinb(G8), .dout(new_n347_));
  anb2 g274(.dina(new_n346_), .dinb(new_n347_), .dout(G475));
  anb1 g275(.dina(new_n184_), .dinb(new_n147_), .dout(new_n349_));
  nor2 g276(.dina(new_n312_), .dinb(new_n349_), .dout(new_n350_));
  anb1 g277(.dina(new_n110_), .dinb(new_n350_), .dout(new_n351_));
  anb1 g278(.dina(new_n351_), .dinb(G9), .dout(new_n352_));
  anb2 g279(.dina(new_n351_), .dinb(G9), .dout(new_n353_));
  anb2 g280(.dina(new_n352_), .dinb(new_n353_), .dout(G476));
  anb1 g281(.dina(new_n299_), .dinb(new_n350_), .dout(new_n355_));
  anb1 g282(.dina(new_n355_), .dinb(G10), .dout(new_n356_));
  anb2 g283(.dina(new_n355_), .dinb(G10), .dout(new_n357_));
  anb2 g284(.dina(new_n356_), .dinb(new_n357_), .dout(G477));
  anb1 g285(.dina(new_n280_), .dinb(new_n350_), .dout(new_n359_));
  anb1 g286(.dina(new_n359_), .dinb(G11), .dout(new_n360_));
  anb2 g287(.dina(new_n359_), .dinb(G11), .dout(new_n361_));
  anb2 g288(.dina(new_n360_), .dinb(new_n361_), .dout(G478));
  anb1 g289(.dina(new_n252_), .dinb(new_n350_), .dout(new_n363_));
  anb1 g290(.dina(new_n363_), .dinb(G12), .dout(new_n364_));
  anb2 g291(.dina(new_n363_), .dinb(G12), .dout(new_n365_));
  anb2 g292(.dina(new_n364_), .dinb(new_n365_), .dout(G479));
  nab1 g293(.dina(new_n223_), .dinb(new_n349_), .dout(new_n367_));
  nor2 g294(.dina(new_n331_), .dinb(new_n367_), .dout(new_n368_));
  anb1 g295(.dina(new_n110_), .dinb(new_n368_), .dout(new_n369_));
  anb1 g296(.dina(new_n369_), .dinb(G13), .dout(new_n370_));
  anb2 g297(.dina(new_n369_), .dinb(G13), .dout(new_n371_));
  anb2 g298(.dina(new_n370_), .dinb(new_n371_), .dout(G480));
  anb1 g299(.dina(new_n299_), .dinb(new_n368_), .dout(new_n373_));
  anb1 g300(.dina(new_n373_), .dinb(G14), .dout(new_n374_));
  anb2 g301(.dina(new_n373_), .dinb(G14), .dout(new_n375_));
  anb2 g302(.dina(new_n374_), .dinb(new_n375_), .dout(G481));
  anb1 g303(.dina(new_n280_), .dinb(new_n368_), .dout(new_n377_));
  anb1 g304(.dina(new_n377_), .dinb(G15), .dout(new_n378_));
  anb2 g305(.dina(new_n377_), .dinb(G15), .dout(new_n379_));
  anb2 g306(.dina(new_n378_), .dinb(new_n379_), .dout(G482));
  anb1 g307(.dina(new_n252_), .dinb(new_n368_), .dout(new_n381_));
  anb1 g308(.dina(new_n381_), .dinb(G16), .dout(new_n382_));
  anb2 g309(.dina(new_n381_), .dinb(G16), .dout(new_n383_));
  anb2 g310(.dina(new_n382_), .dinb(new_n383_), .dout(G483));
  anb1 g311(.dina(new_n330_), .dinb(new_n367_), .dout(new_n385_));
  and2 g312(.dina(new_n204_), .dinb(new_n385_), .dout(new_n386_));
  anb2 g313(.dina(new_n223_), .dinb(new_n204_), .dout(new_n387_));
  anb2 g314(.dina(new_n224_), .dinb(new_n387_), .dout(new_n388_));
  and2 g315(.dina(new_n147_), .dinb(new_n184_), .dout(new_n389_));
  anb1 g316(.dina(new_n388_), .dinb(new_n389_), .dout(new_n390_));
  anb1 g317(.dina(new_n386_), .dinb(new_n390_), .dout(new_n391_));
  anb1 g318(.dina(new_n300_), .dinb(new_n306_), .dout(new_n392_));
  anb2 g319(.dina(new_n391_), .dinb(new_n392_), .dout(new_n393_));
  anb1 g320(.dina(new_n147_), .dinb(new_n393_), .dout(new_n394_));
  anb1 g321(.dina(new_n394_), .dinb(G17), .dout(new_n395_));
  anb2 g322(.dina(new_n394_), .dinb(G17), .dout(new_n396_));
  anb2 g323(.dina(new_n395_), .dinb(new_n396_), .dout(G484));
  anb1 g324(.dina(new_n184_), .dinb(new_n393_), .dout(new_n398_));
  anb1 g325(.dina(new_n398_), .dinb(G18), .dout(new_n399_));
  anb2 g326(.dina(new_n398_), .dinb(G18), .dout(new_n400_));
  anb2 g327(.dina(new_n399_), .dinb(new_n400_), .dout(G485));
  anb1 g328(.dina(new_n223_), .dinb(new_n393_), .dout(new_n402_));
  anb1 g329(.dina(new_n402_), .dinb(G19), .dout(new_n403_));
  anb2 g330(.dina(new_n402_), .dinb(G19), .dout(new_n404_));
  anb2 g331(.dina(new_n403_), .dinb(new_n404_), .dout(G486));
  anb1 g332(.dina(new_n204_), .dinb(new_n393_), .dout(new_n406_));
  anb1 g333(.dina(new_n406_), .dinb(G20), .dout(new_n407_));
  anb2 g334(.dina(new_n406_), .dinb(G20), .dout(new_n408_));
  anb2 g335(.dina(new_n407_), .dinb(new_n408_), .dout(G487));
  anb1 g336(.dina(new_n252_), .dinb(new_n391_), .dout(new_n410_));
  anb2 g337(.dina(new_n301_), .dinb(new_n410_), .dout(new_n411_));
  anb1 g338(.dina(new_n147_), .dinb(new_n411_), .dout(new_n412_));
  anb1 g339(.dina(new_n412_), .dinb(G21), .dout(new_n413_));
  anb2 g340(.dina(new_n412_), .dinb(G21), .dout(new_n414_));
  anb2 g341(.dina(new_n413_), .dinb(new_n414_), .dout(G488));
  anb1 g342(.dina(new_n184_), .dinb(new_n411_), .dout(new_n416_));
  anb1 g343(.dina(new_n416_), .dinb(G22), .dout(new_n417_));
  anb2 g344(.dina(new_n416_), .dinb(G22), .dout(new_n418_));
  anb2 g345(.dina(new_n417_), .dinb(new_n418_), .dout(G489));
  anb1 g346(.dina(new_n223_), .dinb(new_n411_), .dout(new_n420_));
  anb1 g347(.dina(new_n420_), .dinb(G23), .dout(new_n421_));
  anb2 g348(.dina(new_n420_), .dinb(G23), .dout(new_n422_));
  anb2 g349(.dina(new_n421_), .dinb(new_n422_), .dout(G490));
  anb1 g350(.dina(new_n204_), .dinb(new_n411_), .dout(new_n424_));
  anb1 g351(.dina(new_n424_), .dinb(G24), .dout(new_n425_));
  anb2 g352(.dina(new_n424_), .dinb(G24), .dout(new_n426_));
  anb2 g353(.dina(new_n425_), .dinb(new_n426_), .dout(G491));
  anb1 g354(.dina(new_n302_), .dinb(new_n306_), .dout(new_n428_));
  anb2 g355(.dina(new_n391_), .dinb(new_n428_), .dout(new_n429_));
  anb1 g356(.dina(new_n147_), .dinb(new_n429_), .dout(new_n430_));
  anb1 g357(.dina(new_n430_), .dinb(G25), .dout(new_n431_));
  anb2 g358(.dina(new_n430_), .dinb(G25), .dout(new_n432_));
  anb2 g359(.dina(new_n431_), .dinb(new_n432_), .dout(G492));
  anb1 g360(.dina(new_n184_), .dinb(new_n429_), .dout(new_n434_));
  anb1 g361(.dina(new_n434_), .dinb(G26), .dout(new_n435_));
  anb2 g362(.dina(new_n434_), .dinb(G26), .dout(new_n436_));
  anb2 g363(.dina(new_n435_), .dinb(new_n436_), .dout(G493));
  anb1 g364(.dina(new_n223_), .dinb(new_n429_), .dout(new_n438_));
  anb1 g365(.dina(new_n438_), .dinb(G27), .dout(new_n439_));
  anb2 g366(.dina(new_n438_), .dinb(G27), .dout(new_n440_));
  anb2 g367(.dina(new_n439_), .dinb(new_n440_), .dout(G494));
  anb1 g368(.dina(new_n204_), .dinb(new_n429_), .dout(new_n442_));
  anb1 g369(.dina(new_n442_), .dinb(G28), .dout(new_n443_));
  anb2 g370(.dina(new_n442_), .dinb(G28), .dout(new_n444_));
  anb2 g371(.dina(new_n443_), .dinb(new_n444_), .dout(G495));
  anb2 g372(.dina(new_n303_), .dinb(new_n410_), .dout(new_n446_));
  anb1 g373(.dina(new_n147_), .dinb(new_n446_), .dout(new_n447_));
  anb1 g374(.dina(new_n447_), .dinb(G29), .dout(new_n448_));
  anb2 g375(.dina(new_n447_), .dinb(G29), .dout(new_n449_));
  anb2 g376(.dina(new_n448_), .dinb(new_n449_), .dout(G496));
  anb1 g377(.dina(new_n184_), .dinb(new_n446_), .dout(new_n451_));
  anb1 g378(.dina(new_n451_), .dinb(G30), .dout(new_n452_));
  anb2 g379(.dina(new_n451_), .dinb(G30), .dout(new_n453_));
  anb2 g380(.dina(new_n452_), .dinb(new_n453_), .dout(G497));
  anb1 g381(.dina(new_n223_), .dinb(new_n446_), .dout(new_n455_));
  anb1 g382(.dina(new_n455_), .dinb(G31), .dout(new_n456_));
  anb2 g383(.dina(new_n455_), .dinb(G31), .dout(new_n457_));
  anb2 g384(.dina(new_n456_), .dinb(new_n457_), .dout(G498));
  anb1 g385(.dina(new_n204_), .dinb(new_n446_), .dout(new_n459_));
  anb1 g386(.dina(new_n459_), .dinb(G32), .dout(new_n460_));
  anb2 g387(.dina(new_n459_), .dinb(G32), .dout(new_n461_));
  anb2 g388(.dina(new_n460_), .dinb(new_n461_), .dout(G499));
endmodule


