
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  n229_lo,
  n253_lo,
  n256_lo,
  n259_lo,
  n262_lo,
  n277_lo,
  n301_lo,
  n304_lo,
  n307_lo,
  n310_lo,
  n325_lo,
  n349_lo,
  n352_lo,
  n355_lo,
  n358_lo,
  n373_lo,
  n397_lo,
  n400_lo,
  n403_lo,
  n406_lo,
  n421_lo,
  n445_lo,
  n448_lo,
  n451_lo,
  n454_lo,
  n469_lo,
  n493_lo,
  n496_lo,
  n499_lo,
  n502_lo,
  n517_lo,
  n520_lo,
  n541_lo,
  n544_lo,
  n547_lo,
  n550_lo,
  n565_lo,
  n589_lo,
  n592_lo,
  n595_lo,
  n598_lo,
  n613_lo,
  n625_lo,
  n628_lo,
  n631_lo,
  n634_lo,
  n852_o2,
  n853_o2,
  n955_o2,
  n956_o2,
  n531_o2,
  n549_o2,
  n537_o2,
  n540_o2,
  n546_o2,
  n534_o2,
  n552_o2,
  n543_o2,
  n961_o2,
  n223_inv,
  n555_o2,
  n1009_o2,
  n1010_o2,
  n1011_o2,
  n1012_o2,
  lo026_buf_o2,
  lo074_buf_o2,
  lo090_buf_o2,
  lo122_buf_o2,
  n510_o2,
  n498_o2,
  n516_o2,
  n507_o2,
  lo106_buf_o2,
  n519_o2,
  n1029_o2,
  n1041_o2,
  n1043_o2,
  n1045_o2,
  n558_o2,
  n563_o2,
  lo094_buf_o2,
  lo102_buf_o2,
  n522_o2,
  n298_inv,
  n486_o2,
  n304_inv,
  n564_o2,
  n528_o2,
  n492_o2,
  n530_o2,
  n548_o2,
  n536_o2,
  n539_o2,
  lo025_buf_o2,
  lo073_buf_o2,
  lo089_buf_o2,
  lo121_buf_o2,
  n509_o2,
  n513_o2,
  n501_o2,
  n504_o2,
  n495_o2,
  n497_o2,
  n515_o2,
  n506_o2,
  lo010_buf_o2,
  lo042_buf_o2,
  lo058_buf_o2,
  lo138_buf_o2,
  lo014_buf_o2,
  lo022_buf_o2,
  lo030_buf_o2,
  lo038_buf_o2,
  lo046_buf_o2,
  lo054_buf_o2,
  lo126_buf_o2,
  lo134_buf_o2,
  lo093_buf_o2,
  lo101_buf_o2,
  lo002_buf_o2,
  lo006_buf_o2,
  lo062_buf_o2,
  lo070_buf_o2,
  lo078_buf_o2,
  lo086_buf_o2,
  lo110_buf_o2,
  lo118_buf_o2,
  n476_o2,
  n482_o2,
  n478_o2,
  n479_o2,
  G426,
  G427,
  G428,
  G429,
  G430,
  G431,
  G432,
  n856_li008_li008,
  n880_li016_li016,
  n883_li017_li017,
  n886_li018_li018,
  n889_li019_li019,
  n904_li024_li024,
  n928_li032_li032,
  n931_li033_li033,
  n934_li034_li034,
  n937_li035_li035,
  n952_li040_li040,
  n976_li048_li048,
  n979_li049_li049,
  n982_li050_li050,
  n985_li051_li051,
  n1000_li056_li056,
  n1024_li064_li064,
  n1027_li065_li065,
  n1030_li066_li066,
  n1033_li067_li067,
  n1048_li072_li072,
  n1072_li080_li080,
  n1075_li081_li081,
  n1078_li082_li082,
  n1081_li083_li083,
  n1096_li088_li088,
  n1120_li096_li096,
  n1123_li097_li097,
  n1126_li098_li098,
  n1129_li099_li099,
  n1144_li104_li104,
  n1147_li105_li105,
  n1168_li112_li112,
  n1171_li113_li113,
  n1174_li114_li114,
  n1177_li115_li115,
  n1192_li120_li120,
  n1216_li128_li128,
  n1219_li129_li129,
  n1222_li130_li130,
  n1225_li131_li131,
  n1240_li136_li136,
  n1252_li140_li140,
  n1255_li141_li141,
  n1258_li142_li142,
  n1261_li143_li143,
  n852_i2,
  n853_i2,
  n955_i2,
  n956_i2,
  n531_i2,
  n549_i2,
  n537_i2,
  n540_i2,
  n546_i2,
  n534_i2,
  n552_i2,
  n543_i2,
  n961_i2,
  n962_i2,
  n555_i2,
  n1009_i2,
  n1010_i2,
  n1011_i2,
  n1012_i2,
  lo026_buf_i2,
  lo074_buf_i2,
  lo090_buf_i2,
  lo122_buf_i2,
  n510_i2,
  n498_i2,
  n516_i2,
  n507_i2,
  lo106_buf_i2,
  n519_i2,
  n1029_i2,
  n1041_i2,
  n1043_i2,
  n1045_i2,
  n558_i2,
  n563_i2,
  lo094_buf_i2,
  lo102_buf_i2,
  n522_i2,
  n527_i2,
  n486_i2,
  n491_i2,
  n564_i2,
  n528_i2,
  n492_i2,
  n530_i2,
  n548_i2,
  n536_i2,
  n539_i2,
  lo025_buf_i2,
  lo073_buf_i2,
  lo089_buf_i2,
  lo121_buf_i2,
  n509_i2,
  n513_i2,
  n501_i2,
  n504_i2,
  n495_i2,
  n497_i2,
  n515_i2,
  n506_i2,
  lo010_buf_i2,
  lo042_buf_i2,
  lo058_buf_i2,
  lo138_buf_i2,
  lo014_buf_i2,
  lo022_buf_i2,
  lo030_buf_i2,
  lo038_buf_i2,
  lo046_buf_i2,
  lo054_buf_i2,
  lo126_buf_i2,
  lo134_buf_i2,
  lo093_buf_i2,
  lo101_buf_i2,
  lo002_buf_i2,
  lo006_buf_i2,
  lo062_buf_i2,
  lo070_buf_i2,
  lo078_buf_i2,
  lo086_buf_i2,
  lo110_buf_i2,
  lo118_buf_i2,
  n476_i2,
  n482_i2,
  n478_i2,
  n479_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input n229_lo;input n253_lo;input n256_lo;input n259_lo;input n262_lo;input n277_lo;input n301_lo;input n304_lo;input n307_lo;input n310_lo;input n325_lo;input n349_lo;input n352_lo;input n355_lo;input n358_lo;input n373_lo;input n397_lo;input n400_lo;input n403_lo;input n406_lo;input n421_lo;input n445_lo;input n448_lo;input n451_lo;input n454_lo;input n469_lo;input n493_lo;input n496_lo;input n499_lo;input n502_lo;input n517_lo;input n520_lo;input n541_lo;input n544_lo;input n547_lo;input n550_lo;input n565_lo;input n589_lo;input n592_lo;input n595_lo;input n598_lo;input n613_lo;input n625_lo;input n628_lo;input n631_lo;input n634_lo;input n852_o2;input n853_o2;input n955_o2;input n956_o2;input n531_o2;input n549_o2;input n537_o2;input n540_o2;input n546_o2;input n534_o2;input n552_o2;input n543_o2;input n961_o2;input n223_inv;input n555_o2;input n1009_o2;input n1010_o2;input n1011_o2;input n1012_o2;input lo026_buf_o2;input lo074_buf_o2;input lo090_buf_o2;input lo122_buf_o2;input n510_o2;input n498_o2;input n516_o2;input n507_o2;input lo106_buf_o2;input n519_o2;input n1029_o2;input n1041_o2;input n1043_o2;input n1045_o2;input n558_o2;input n563_o2;input lo094_buf_o2;input lo102_buf_o2;input n522_o2;input n298_inv;input n486_o2;input n304_inv;input n564_o2;input n528_o2;input n492_o2;input n530_o2;input n548_o2;input n536_o2;input n539_o2;input lo025_buf_o2;input lo073_buf_o2;input lo089_buf_o2;input lo121_buf_o2;input n509_o2;input n513_o2;input n501_o2;input n504_o2;input n495_o2;input n497_o2;input n515_o2;input n506_o2;input lo010_buf_o2;input lo042_buf_o2;input lo058_buf_o2;input lo138_buf_o2;input lo014_buf_o2;input lo022_buf_o2;input lo030_buf_o2;input lo038_buf_o2;input lo046_buf_o2;input lo054_buf_o2;input lo126_buf_o2;input lo134_buf_o2;input lo093_buf_o2;input lo101_buf_o2;input lo002_buf_o2;input lo006_buf_o2;input lo062_buf_o2;input lo070_buf_o2;input lo078_buf_o2;input lo086_buf_o2;input lo110_buf_o2;input lo118_buf_o2;input n476_o2;input n482_o2;input n478_o2;input n479_o2;
  output G426;output G427;output G428;output G429;output G430;output G431;output G432;output n856_li008_li008;output n880_li016_li016;output n883_li017_li017;output n886_li018_li018;output n889_li019_li019;output n904_li024_li024;output n928_li032_li032;output n931_li033_li033;output n934_li034_li034;output n937_li035_li035;output n952_li040_li040;output n976_li048_li048;output n979_li049_li049;output n982_li050_li050;output n985_li051_li051;output n1000_li056_li056;output n1024_li064_li064;output n1027_li065_li065;output n1030_li066_li066;output n1033_li067_li067;output n1048_li072_li072;output n1072_li080_li080;output n1075_li081_li081;output n1078_li082_li082;output n1081_li083_li083;output n1096_li088_li088;output n1120_li096_li096;output n1123_li097_li097;output n1126_li098_li098;output n1129_li099_li099;output n1144_li104_li104;output n1147_li105_li105;output n1168_li112_li112;output n1171_li113_li113;output n1174_li114_li114;output n1177_li115_li115;output n1192_li120_li120;output n1216_li128_li128;output n1219_li129_li129;output n1222_li130_li130;output n1225_li131_li131;output n1240_li136_li136;output n1252_li140_li140;output n1255_li141_li141;output n1258_li142_li142;output n1261_li143_li143;output n852_i2;output n853_i2;output n955_i2;output n956_i2;output n531_i2;output n549_i2;output n537_i2;output n540_i2;output n546_i2;output n534_i2;output n552_i2;output n543_i2;output n961_i2;output n962_i2;output n555_i2;output n1009_i2;output n1010_i2;output n1011_i2;output n1012_i2;output lo026_buf_i2;output lo074_buf_i2;output lo090_buf_i2;output lo122_buf_i2;output n510_i2;output n498_i2;output n516_i2;output n507_i2;output lo106_buf_i2;output n519_i2;output n1029_i2;output n1041_i2;output n1043_i2;output n1045_i2;output n558_i2;output n563_i2;output lo094_buf_i2;output lo102_buf_i2;output n522_i2;output n527_i2;output n486_i2;output n491_i2;output n564_i2;output n528_i2;output n492_i2;output n530_i2;output n548_i2;output n536_i2;output n539_i2;output lo025_buf_i2;output lo073_buf_i2;output lo089_buf_i2;output lo121_buf_i2;output n509_i2;output n513_i2;output n501_i2;output n504_i2;output n495_i2;output n497_i2;output n515_i2;output n506_i2;output lo010_buf_i2;output lo042_buf_i2;output lo058_buf_i2;output lo138_buf_i2;output lo014_buf_i2;output lo022_buf_i2;output lo030_buf_i2;output lo038_buf_i2;output lo046_buf_i2;output lo054_buf_i2;output lo126_buf_i2;output lo134_buf_i2;output lo093_buf_i2;output lo101_buf_i2;output lo002_buf_i2;output lo006_buf_i2;output lo062_buf_i2;output lo070_buf_i2;output lo078_buf_i2;output lo086_buf_i2;output lo110_buf_i2;output lo118_buf_i2;output n476_i2;output n482_i2;output n478_i2;output n479_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire n229_lo_p;
  wire n229_lo_n;
  wire n253_lo_p;
  wire n253_lo_n;
  wire n256_lo_p;
  wire n256_lo_n;
  wire n259_lo_p;
  wire n259_lo_n;
  wire n262_lo_p;
  wire n262_lo_n;
  wire n277_lo_p;
  wire n277_lo_n;
  wire n301_lo_p;
  wire n301_lo_n;
  wire n304_lo_p;
  wire n304_lo_n;
  wire n307_lo_p;
  wire n307_lo_n;
  wire n310_lo_p;
  wire n310_lo_n;
  wire n325_lo_p;
  wire n325_lo_n;
  wire n349_lo_p;
  wire n349_lo_n;
  wire n352_lo_p;
  wire n352_lo_n;
  wire n355_lo_p;
  wire n355_lo_n;
  wire n358_lo_p;
  wire n358_lo_n;
  wire n373_lo_p;
  wire n373_lo_n;
  wire n397_lo_p;
  wire n397_lo_n;
  wire n400_lo_p;
  wire n400_lo_n;
  wire n403_lo_p;
  wire n403_lo_n;
  wire n406_lo_p;
  wire n406_lo_n;
  wire n421_lo_p;
  wire n421_lo_n;
  wire n445_lo_p;
  wire n445_lo_n;
  wire n448_lo_p;
  wire n448_lo_n;
  wire n451_lo_p;
  wire n451_lo_n;
  wire n454_lo_p;
  wire n454_lo_n;
  wire n469_lo_p;
  wire n469_lo_n;
  wire n493_lo_p;
  wire n493_lo_n;
  wire n496_lo_p;
  wire n496_lo_n;
  wire n499_lo_p;
  wire n499_lo_n;
  wire n502_lo_p;
  wire n502_lo_n;
  wire n517_lo_p;
  wire n517_lo_n;
  wire n520_lo_p;
  wire n520_lo_n;
  wire n541_lo_p;
  wire n541_lo_n;
  wire n544_lo_p;
  wire n544_lo_n;
  wire n547_lo_p;
  wire n547_lo_n;
  wire n550_lo_p;
  wire n550_lo_n;
  wire n565_lo_p;
  wire n565_lo_n;
  wire n589_lo_p;
  wire n589_lo_n;
  wire n592_lo_p;
  wire n592_lo_n;
  wire n595_lo_p;
  wire n595_lo_n;
  wire n598_lo_p;
  wire n598_lo_n;
  wire n613_lo_p;
  wire n613_lo_n;
  wire n625_lo_p;
  wire n625_lo_n;
  wire n628_lo_p;
  wire n628_lo_n;
  wire n631_lo_p;
  wire n631_lo_n;
  wire n634_lo_p;
  wire n634_lo_n;
  wire n852_o2_p;
  wire n852_o2_n;
  wire n853_o2_p;
  wire n853_o2_n;
  wire n955_o2_p;
  wire n955_o2_n;
  wire n956_o2_p;
  wire n956_o2_n;
  wire n531_o2_p;
  wire n531_o2_n;
  wire n549_o2_p;
  wire n549_o2_n;
  wire n537_o2_p;
  wire n537_o2_n;
  wire n540_o2_p;
  wire n540_o2_n;
  wire n546_o2_p;
  wire n546_o2_n;
  wire n534_o2_p;
  wire n534_o2_n;
  wire n552_o2_p;
  wire n552_o2_n;
  wire n543_o2_p;
  wire n543_o2_n;
  wire n961_o2_p;
  wire n961_o2_n;
  wire n223_inv_p;
  wire n223_inv_n;
  wire n555_o2_p;
  wire n555_o2_n;
  wire n1009_o2_p;
  wire n1009_o2_n;
  wire n1010_o2_p;
  wire n1010_o2_n;
  wire n1011_o2_p;
  wire n1011_o2_n;
  wire n1012_o2_p;
  wire n1012_o2_n;
  wire lo026_buf_o2_p;
  wire lo026_buf_o2_n;
  wire lo074_buf_o2_p;
  wire lo074_buf_o2_n;
  wire lo090_buf_o2_p;
  wire lo090_buf_o2_n;
  wire lo122_buf_o2_p;
  wire lo122_buf_o2_n;
  wire n510_o2_p;
  wire n510_o2_n;
  wire n498_o2_p;
  wire n498_o2_n;
  wire n516_o2_p;
  wire n516_o2_n;
  wire n507_o2_p;
  wire n507_o2_n;
  wire lo106_buf_o2_p;
  wire lo106_buf_o2_n;
  wire n519_o2_p;
  wire n519_o2_n;
  wire n1029_o2_p;
  wire n1029_o2_n;
  wire n1041_o2_p;
  wire n1041_o2_n;
  wire n1043_o2_p;
  wire n1043_o2_n;
  wire n1045_o2_p;
  wire n1045_o2_n;
  wire n558_o2_p;
  wire n558_o2_n;
  wire n563_o2_p;
  wire n563_o2_n;
  wire lo094_buf_o2_p;
  wire lo094_buf_o2_n;
  wire lo102_buf_o2_p;
  wire lo102_buf_o2_n;
  wire n522_o2_p;
  wire n522_o2_n;
  wire n298_inv_p;
  wire n298_inv_n;
  wire n486_o2_p;
  wire n486_o2_n;
  wire n304_inv_p;
  wire n304_inv_n;
  wire n564_o2_p;
  wire n564_o2_n;
  wire n528_o2_p;
  wire n528_o2_n;
  wire n492_o2_p;
  wire n492_o2_n;
  wire n530_o2_p;
  wire n530_o2_n;
  wire n548_o2_p;
  wire n548_o2_n;
  wire n536_o2_p;
  wire n536_o2_n;
  wire n539_o2_p;
  wire n539_o2_n;
  wire lo025_buf_o2_p;
  wire lo025_buf_o2_n;
  wire lo073_buf_o2_p;
  wire lo073_buf_o2_n;
  wire lo089_buf_o2_p;
  wire lo089_buf_o2_n;
  wire lo121_buf_o2_p;
  wire lo121_buf_o2_n;
  wire n509_o2_p;
  wire n509_o2_n;
  wire n513_o2_p;
  wire n513_o2_n;
  wire n501_o2_p;
  wire n501_o2_n;
  wire n504_o2_p;
  wire n504_o2_n;
  wire n495_o2_p;
  wire n495_o2_n;
  wire n497_o2_p;
  wire n497_o2_n;
  wire n515_o2_p;
  wire n515_o2_n;
  wire n506_o2_p;
  wire n506_o2_n;
  wire lo010_buf_o2_p;
  wire lo010_buf_o2_n;
  wire lo042_buf_o2_p;
  wire lo042_buf_o2_n;
  wire lo058_buf_o2_p;
  wire lo058_buf_o2_n;
  wire lo138_buf_o2_p;
  wire lo138_buf_o2_n;
  wire lo014_buf_o2_p;
  wire lo014_buf_o2_n;
  wire lo022_buf_o2_p;
  wire lo022_buf_o2_n;
  wire lo030_buf_o2_p;
  wire lo030_buf_o2_n;
  wire lo038_buf_o2_p;
  wire lo038_buf_o2_n;
  wire lo046_buf_o2_p;
  wire lo046_buf_o2_n;
  wire lo054_buf_o2_p;
  wire lo054_buf_o2_n;
  wire lo126_buf_o2_p;
  wire lo126_buf_o2_n;
  wire lo134_buf_o2_p;
  wire lo134_buf_o2_n;
  wire lo093_buf_o2_p;
  wire lo093_buf_o2_n;
  wire lo101_buf_o2_p;
  wire lo101_buf_o2_n;
  wire lo002_buf_o2_p;
  wire lo002_buf_o2_n;
  wire lo006_buf_o2_p;
  wire lo006_buf_o2_n;
  wire lo062_buf_o2_p;
  wire lo062_buf_o2_n;
  wire lo070_buf_o2_p;
  wire lo070_buf_o2_n;
  wire lo078_buf_o2_p;
  wire lo078_buf_o2_n;
  wire lo086_buf_o2_p;
  wire lo086_buf_o2_n;
  wire lo110_buf_o2_p;
  wire lo110_buf_o2_n;
  wire lo118_buf_o2_p;
  wire lo118_buf_o2_n;
  wire n476_o2_p;
  wire n476_o2_n;
  wire n482_o2_p;
  wire n482_o2_n;
  wire n478_o2_p;
  wire n478_o2_n;
  wire n479_o2_p;
  wire n479_o2_n;
  wire g169_p;
  wire g169_n;
  wire g170_p;
  wire g170_n;
  wire g171_p;
  wire g171_n;
  wire g172_p;
  wire g172_n;
  wire g173_p;
  wire g173_n;
  wire g174_p;
  wire g174_n;
  wire g175_p;
  wire g175_n;
  wire g176_p;
  wire g176_n;
  wire g177_p;
  wire g177_n;
  wire g178_p;
  wire g178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire n564_o2_n_spl_;
  wire n564_o2_n_spl_0;
  wire n564_o2_n_spl_00;
  wire n564_o2_n_spl_1;
  wire n564_o2_p_spl_;
  wire n564_o2_p_spl_0;
  wire n564_o2_p_spl_00;
  wire n564_o2_p_spl_01;
  wire n564_o2_p_spl_1;
  wire n564_o2_p_spl_10;
  wire n564_o2_p_spl_11;
  wire g175_n_spl_;
  wire g177_n_spl_;
  wire g180_n_spl_;
  wire g186_n_spl_;
  wire g186_p_spl_;
  wire g188_p_spl_;
  wire g191_n_spl_;
  wire g193_n_spl_;
  wire g195_p_spl_;
  wire g193_p_spl_;
  wire g200_p_spl_;
  wire n528_o2_p_spl_;
  wire n528_o2_p_spl_0;
  wire n528_o2_p_spl_00;
  wire n528_o2_p_spl_1;
  wire n547_lo_p_spl_;
  wire g222_n_spl_;
  wire n595_lo_p_spl_;
  wire g220_n_spl_;
  wire n307_lo_p_spl_;
  wire g214_n_spl_;
  wire n451_lo_p_spl_;
  wire g216_n_spl_;
  wire n499_lo_p_spl_;
  wire g218_n_spl_;
  wire n259_lo_p_spl_;
  wire g209_n_spl_;
  wire n631_lo_p_spl_;
  wire g212_n_spl_;
  wire n403_lo_p_spl_;
  wire g211_n_spl_;
  wire n355_lo_p_spl_;
  wire g210_n_spl_;
  wire n520_lo_p_spl_;
  wire g228_n_spl_;
  wire lo121_buf_o2_p_spl_;
  wire g226_n_spl_;
  wire lo025_buf_o2_p_spl_;
  wire g223_n_spl_;
  wire lo073_buf_o2_p_spl_;
  wire g224_n_spl_;
  wire lo089_buf_o2_p_spl_;
  wire g225_n_spl_;
  wire lo101_buf_o2_p_spl_;
  wire lo118_buf_o2_p_spl_;
  wire lo070_buf_o2_p_spl_;
  wire lo086_buf_o2_p_spl_;
  wire g233_p_spl_;
  wire g244_p_spl_;
  wire g249_p_spl_;
  wire g260_p_spl_;
  wire g265_n_spl_;
  wire g272_n_spl_;
  wire g274_p_spl_;
  wire g274_p_spl_0;
  wire g274_p_spl_00;
  wire g274_p_spl_1;
  wire g275_n_spl_;
  wire g275_n_spl_0;
  wire g275_n_spl_00;
  wire g275_n_spl_000;
  wire g275_n_spl_01;
  wire g275_n_spl_1;
  wire g275_n_spl_10;
  wire g275_n_spl_11;
  wire G6_p_spl_;
  wire G10_p_spl_;
  wire G14_p_spl_;
  wire G34_p_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    n229_lo_p,
    n229_lo
  );


  not

  (
    n229_lo_n,
    n229_lo
  );


  buf

  (
    n253_lo_p,
    n253_lo
  );


  not

  (
    n253_lo_n,
    n253_lo
  );


  buf

  (
    n256_lo_p,
    n256_lo
  );


  not

  (
    n256_lo_n,
    n256_lo
  );


  buf

  (
    n259_lo_p,
    n259_lo
  );


  not

  (
    n259_lo_n,
    n259_lo
  );


  buf

  (
    n262_lo_p,
    n262_lo
  );


  not

  (
    n262_lo_n,
    n262_lo
  );


  buf

  (
    n277_lo_p,
    n277_lo
  );


  not

  (
    n277_lo_n,
    n277_lo
  );


  buf

  (
    n301_lo_p,
    n301_lo
  );


  not

  (
    n301_lo_n,
    n301_lo
  );


  buf

  (
    n304_lo_p,
    n304_lo
  );


  not

  (
    n304_lo_n,
    n304_lo
  );


  buf

  (
    n307_lo_p,
    n307_lo
  );


  not

  (
    n307_lo_n,
    n307_lo
  );


  buf

  (
    n310_lo_p,
    n310_lo
  );


  not

  (
    n310_lo_n,
    n310_lo
  );


  buf

  (
    n325_lo_p,
    n325_lo
  );


  not

  (
    n325_lo_n,
    n325_lo
  );


  buf

  (
    n349_lo_p,
    n349_lo
  );


  not

  (
    n349_lo_n,
    n349_lo
  );


  buf

  (
    n352_lo_p,
    n352_lo
  );


  not

  (
    n352_lo_n,
    n352_lo
  );


  buf

  (
    n355_lo_p,
    n355_lo
  );


  not

  (
    n355_lo_n,
    n355_lo
  );


  buf

  (
    n358_lo_p,
    n358_lo
  );


  not

  (
    n358_lo_n,
    n358_lo
  );


  buf

  (
    n373_lo_p,
    n373_lo
  );


  not

  (
    n373_lo_n,
    n373_lo
  );


  buf

  (
    n397_lo_p,
    n397_lo
  );


  not

  (
    n397_lo_n,
    n397_lo
  );


  buf

  (
    n400_lo_p,
    n400_lo
  );


  not

  (
    n400_lo_n,
    n400_lo
  );


  buf

  (
    n403_lo_p,
    n403_lo
  );


  not

  (
    n403_lo_n,
    n403_lo
  );


  buf

  (
    n406_lo_p,
    n406_lo
  );


  not

  (
    n406_lo_n,
    n406_lo
  );


  buf

  (
    n421_lo_p,
    n421_lo
  );


  not

  (
    n421_lo_n,
    n421_lo
  );


  buf

  (
    n445_lo_p,
    n445_lo
  );


  not

  (
    n445_lo_n,
    n445_lo
  );


  buf

  (
    n448_lo_p,
    n448_lo
  );


  not

  (
    n448_lo_n,
    n448_lo
  );


  buf

  (
    n451_lo_p,
    n451_lo
  );


  not

  (
    n451_lo_n,
    n451_lo
  );


  buf

  (
    n454_lo_p,
    n454_lo
  );


  not

  (
    n454_lo_n,
    n454_lo
  );


  buf

  (
    n469_lo_p,
    n469_lo
  );


  not

  (
    n469_lo_n,
    n469_lo
  );


  buf

  (
    n493_lo_p,
    n493_lo
  );


  not

  (
    n493_lo_n,
    n493_lo
  );


  buf

  (
    n496_lo_p,
    n496_lo
  );


  not

  (
    n496_lo_n,
    n496_lo
  );


  buf

  (
    n499_lo_p,
    n499_lo
  );


  not

  (
    n499_lo_n,
    n499_lo
  );


  buf

  (
    n502_lo_p,
    n502_lo
  );


  not

  (
    n502_lo_n,
    n502_lo
  );


  buf

  (
    n517_lo_p,
    n517_lo
  );


  not

  (
    n517_lo_n,
    n517_lo
  );


  buf

  (
    n520_lo_p,
    n520_lo
  );


  not

  (
    n520_lo_n,
    n520_lo
  );


  buf

  (
    n541_lo_p,
    n541_lo
  );


  not

  (
    n541_lo_n,
    n541_lo
  );


  buf

  (
    n544_lo_p,
    n544_lo
  );


  not

  (
    n544_lo_n,
    n544_lo
  );


  buf

  (
    n547_lo_p,
    n547_lo
  );


  not

  (
    n547_lo_n,
    n547_lo
  );


  buf

  (
    n550_lo_p,
    n550_lo
  );


  not

  (
    n550_lo_n,
    n550_lo
  );


  buf

  (
    n565_lo_p,
    n565_lo
  );


  not

  (
    n565_lo_n,
    n565_lo
  );


  buf

  (
    n589_lo_p,
    n589_lo
  );


  not

  (
    n589_lo_n,
    n589_lo
  );


  buf

  (
    n592_lo_p,
    n592_lo
  );


  not

  (
    n592_lo_n,
    n592_lo
  );


  buf

  (
    n595_lo_p,
    n595_lo
  );


  not

  (
    n595_lo_n,
    n595_lo
  );


  buf

  (
    n598_lo_p,
    n598_lo
  );


  not

  (
    n598_lo_n,
    n598_lo
  );


  buf

  (
    n613_lo_p,
    n613_lo
  );


  not

  (
    n613_lo_n,
    n613_lo
  );


  buf

  (
    n625_lo_p,
    n625_lo
  );


  not

  (
    n625_lo_n,
    n625_lo
  );


  buf

  (
    n628_lo_p,
    n628_lo
  );


  not

  (
    n628_lo_n,
    n628_lo
  );


  buf

  (
    n631_lo_p,
    n631_lo
  );


  not

  (
    n631_lo_n,
    n631_lo
  );


  buf

  (
    n634_lo_p,
    n634_lo
  );


  not

  (
    n634_lo_n,
    n634_lo
  );


  buf

  (
    n852_o2_p,
    n852_o2
  );


  not

  (
    n852_o2_n,
    n852_o2
  );


  buf

  (
    n853_o2_p,
    n853_o2
  );


  not

  (
    n853_o2_n,
    n853_o2
  );


  buf

  (
    n955_o2_p,
    n955_o2
  );


  not

  (
    n955_o2_n,
    n955_o2
  );


  buf

  (
    n956_o2_p,
    n956_o2
  );


  not

  (
    n956_o2_n,
    n956_o2
  );


  buf

  (
    n531_o2_p,
    n531_o2
  );


  not

  (
    n531_o2_n,
    n531_o2
  );


  buf

  (
    n549_o2_p,
    n549_o2
  );


  not

  (
    n549_o2_n,
    n549_o2
  );


  buf

  (
    n537_o2_p,
    n537_o2
  );


  not

  (
    n537_o2_n,
    n537_o2
  );


  buf

  (
    n540_o2_p,
    n540_o2
  );


  not

  (
    n540_o2_n,
    n540_o2
  );


  buf

  (
    n546_o2_p,
    n546_o2
  );


  not

  (
    n546_o2_n,
    n546_o2
  );


  buf

  (
    n534_o2_p,
    n534_o2
  );


  not

  (
    n534_o2_n,
    n534_o2
  );


  buf

  (
    n552_o2_p,
    n552_o2
  );


  not

  (
    n552_o2_n,
    n552_o2
  );


  buf

  (
    n543_o2_p,
    n543_o2
  );


  not

  (
    n543_o2_n,
    n543_o2
  );


  buf

  (
    n961_o2_p,
    n961_o2
  );


  not

  (
    n961_o2_n,
    n961_o2
  );


  buf

  (
    n223_inv_p,
    n223_inv
  );


  not

  (
    n223_inv_n,
    n223_inv
  );


  buf

  (
    n555_o2_p,
    n555_o2
  );


  not

  (
    n555_o2_n,
    n555_o2
  );


  buf

  (
    n1009_o2_p,
    n1009_o2
  );


  not

  (
    n1009_o2_n,
    n1009_o2
  );


  buf

  (
    n1010_o2_p,
    n1010_o2
  );


  not

  (
    n1010_o2_n,
    n1010_o2
  );


  buf

  (
    n1011_o2_p,
    n1011_o2
  );


  not

  (
    n1011_o2_n,
    n1011_o2
  );


  buf

  (
    n1012_o2_p,
    n1012_o2
  );


  not

  (
    n1012_o2_n,
    n1012_o2
  );


  buf

  (
    lo026_buf_o2_p,
    lo026_buf_o2
  );


  not

  (
    lo026_buf_o2_n,
    lo026_buf_o2
  );


  buf

  (
    lo074_buf_o2_p,
    lo074_buf_o2
  );


  not

  (
    lo074_buf_o2_n,
    lo074_buf_o2
  );


  buf

  (
    lo090_buf_o2_p,
    lo090_buf_o2
  );


  not

  (
    lo090_buf_o2_n,
    lo090_buf_o2
  );


  buf

  (
    lo122_buf_o2_p,
    lo122_buf_o2
  );


  not

  (
    lo122_buf_o2_n,
    lo122_buf_o2
  );


  buf

  (
    n510_o2_p,
    n510_o2
  );


  not

  (
    n510_o2_n,
    n510_o2
  );


  buf

  (
    n498_o2_p,
    n498_o2
  );


  not

  (
    n498_o2_n,
    n498_o2
  );


  buf

  (
    n516_o2_p,
    n516_o2
  );


  not

  (
    n516_o2_n,
    n516_o2
  );


  buf

  (
    n507_o2_p,
    n507_o2
  );


  not

  (
    n507_o2_n,
    n507_o2
  );


  buf

  (
    lo106_buf_o2_p,
    lo106_buf_o2
  );


  not

  (
    lo106_buf_o2_n,
    lo106_buf_o2
  );


  buf

  (
    n519_o2_p,
    n519_o2
  );


  not

  (
    n519_o2_n,
    n519_o2
  );


  buf

  (
    n1029_o2_p,
    n1029_o2
  );


  not

  (
    n1029_o2_n,
    n1029_o2
  );


  buf

  (
    n1041_o2_p,
    n1041_o2
  );


  not

  (
    n1041_o2_n,
    n1041_o2
  );


  buf

  (
    n1043_o2_p,
    n1043_o2
  );


  not

  (
    n1043_o2_n,
    n1043_o2
  );


  buf

  (
    n1045_o2_p,
    n1045_o2
  );


  not

  (
    n1045_o2_n,
    n1045_o2
  );


  buf

  (
    n558_o2_p,
    n558_o2
  );


  not

  (
    n558_o2_n,
    n558_o2
  );


  buf

  (
    n563_o2_p,
    n563_o2
  );


  not

  (
    n563_o2_n,
    n563_o2
  );


  buf

  (
    lo094_buf_o2_p,
    lo094_buf_o2
  );


  not

  (
    lo094_buf_o2_n,
    lo094_buf_o2
  );


  buf

  (
    lo102_buf_o2_p,
    lo102_buf_o2
  );


  not

  (
    lo102_buf_o2_n,
    lo102_buf_o2
  );


  buf

  (
    n522_o2_p,
    n522_o2
  );


  not

  (
    n522_o2_n,
    n522_o2
  );


  buf

  (
    n298_inv_p,
    n298_inv
  );


  not

  (
    n298_inv_n,
    n298_inv
  );


  buf

  (
    n486_o2_p,
    n486_o2
  );


  not

  (
    n486_o2_n,
    n486_o2
  );


  buf

  (
    n304_inv_p,
    n304_inv
  );


  not

  (
    n304_inv_n,
    n304_inv
  );


  buf

  (
    n564_o2_p,
    n564_o2
  );


  not

  (
    n564_o2_n,
    n564_o2
  );


  buf

  (
    n528_o2_p,
    n528_o2
  );


  not

  (
    n528_o2_n,
    n528_o2
  );


  buf

  (
    n492_o2_p,
    n492_o2
  );


  not

  (
    n492_o2_n,
    n492_o2
  );


  buf

  (
    n530_o2_p,
    n530_o2
  );


  not

  (
    n530_o2_n,
    n530_o2
  );


  buf

  (
    n548_o2_p,
    n548_o2
  );


  not

  (
    n548_o2_n,
    n548_o2
  );


  buf

  (
    n536_o2_p,
    n536_o2
  );


  not

  (
    n536_o2_n,
    n536_o2
  );


  buf

  (
    n539_o2_p,
    n539_o2
  );


  not

  (
    n539_o2_n,
    n539_o2
  );


  buf

  (
    lo025_buf_o2_p,
    lo025_buf_o2
  );


  not

  (
    lo025_buf_o2_n,
    lo025_buf_o2
  );


  buf

  (
    lo073_buf_o2_p,
    lo073_buf_o2
  );


  not

  (
    lo073_buf_o2_n,
    lo073_buf_o2
  );


  buf

  (
    lo089_buf_o2_p,
    lo089_buf_o2
  );


  not

  (
    lo089_buf_o2_n,
    lo089_buf_o2
  );


  buf

  (
    lo121_buf_o2_p,
    lo121_buf_o2
  );


  not

  (
    lo121_buf_o2_n,
    lo121_buf_o2
  );


  buf

  (
    n509_o2_p,
    n509_o2
  );


  not

  (
    n509_o2_n,
    n509_o2
  );


  buf

  (
    n513_o2_p,
    n513_o2
  );


  not

  (
    n513_o2_n,
    n513_o2
  );


  buf

  (
    n501_o2_p,
    n501_o2
  );


  not

  (
    n501_o2_n,
    n501_o2
  );


  buf

  (
    n504_o2_p,
    n504_o2
  );


  not

  (
    n504_o2_n,
    n504_o2
  );


  buf

  (
    n495_o2_p,
    n495_o2
  );


  not

  (
    n495_o2_n,
    n495_o2
  );


  buf

  (
    n497_o2_p,
    n497_o2
  );


  not

  (
    n497_o2_n,
    n497_o2
  );


  buf

  (
    n515_o2_p,
    n515_o2
  );


  not

  (
    n515_o2_n,
    n515_o2
  );


  buf

  (
    n506_o2_p,
    n506_o2
  );


  not

  (
    n506_o2_n,
    n506_o2
  );


  buf

  (
    lo010_buf_o2_p,
    lo010_buf_o2
  );


  not

  (
    lo010_buf_o2_n,
    lo010_buf_o2
  );


  buf

  (
    lo042_buf_o2_p,
    lo042_buf_o2
  );


  not

  (
    lo042_buf_o2_n,
    lo042_buf_o2
  );


  buf

  (
    lo058_buf_o2_p,
    lo058_buf_o2
  );


  not

  (
    lo058_buf_o2_n,
    lo058_buf_o2
  );


  buf

  (
    lo138_buf_o2_p,
    lo138_buf_o2
  );


  not

  (
    lo138_buf_o2_n,
    lo138_buf_o2
  );


  buf

  (
    lo014_buf_o2_p,
    lo014_buf_o2
  );


  not

  (
    lo014_buf_o2_n,
    lo014_buf_o2
  );


  buf

  (
    lo022_buf_o2_p,
    lo022_buf_o2
  );


  not

  (
    lo022_buf_o2_n,
    lo022_buf_o2
  );


  buf

  (
    lo030_buf_o2_p,
    lo030_buf_o2
  );


  not

  (
    lo030_buf_o2_n,
    lo030_buf_o2
  );


  buf

  (
    lo038_buf_o2_p,
    lo038_buf_o2
  );


  not

  (
    lo038_buf_o2_n,
    lo038_buf_o2
  );


  buf

  (
    lo046_buf_o2_p,
    lo046_buf_o2
  );


  not

  (
    lo046_buf_o2_n,
    lo046_buf_o2
  );


  buf

  (
    lo054_buf_o2_p,
    lo054_buf_o2
  );


  not

  (
    lo054_buf_o2_n,
    lo054_buf_o2
  );


  buf

  (
    lo126_buf_o2_p,
    lo126_buf_o2
  );


  not

  (
    lo126_buf_o2_n,
    lo126_buf_o2
  );


  buf

  (
    lo134_buf_o2_p,
    lo134_buf_o2
  );


  not

  (
    lo134_buf_o2_n,
    lo134_buf_o2
  );


  buf

  (
    lo093_buf_o2_p,
    lo093_buf_o2
  );


  not

  (
    lo093_buf_o2_n,
    lo093_buf_o2
  );


  buf

  (
    lo101_buf_o2_p,
    lo101_buf_o2
  );


  not

  (
    lo101_buf_o2_n,
    lo101_buf_o2
  );


  buf

  (
    lo002_buf_o2_p,
    lo002_buf_o2
  );


  not

  (
    lo002_buf_o2_n,
    lo002_buf_o2
  );


  buf

  (
    lo006_buf_o2_p,
    lo006_buf_o2
  );


  not

  (
    lo006_buf_o2_n,
    lo006_buf_o2
  );


  buf

  (
    lo062_buf_o2_p,
    lo062_buf_o2
  );


  not

  (
    lo062_buf_o2_n,
    lo062_buf_o2
  );


  buf

  (
    lo070_buf_o2_p,
    lo070_buf_o2
  );


  not

  (
    lo070_buf_o2_n,
    lo070_buf_o2
  );


  buf

  (
    lo078_buf_o2_p,
    lo078_buf_o2
  );


  not

  (
    lo078_buf_o2_n,
    lo078_buf_o2
  );


  buf

  (
    lo086_buf_o2_p,
    lo086_buf_o2
  );


  not

  (
    lo086_buf_o2_n,
    lo086_buf_o2
  );


  buf

  (
    lo110_buf_o2_p,
    lo110_buf_o2
  );


  not

  (
    lo110_buf_o2_n,
    lo110_buf_o2
  );


  buf

  (
    lo118_buf_o2_p,
    lo118_buf_o2
  );


  not

  (
    lo118_buf_o2_n,
    lo118_buf_o2
  );


  buf

  (
    n476_o2_p,
    n476_o2
  );


  not

  (
    n476_o2_n,
    n476_o2
  );


  buf

  (
    n482_o2_p,
    n482_o2
  );


  not

  (
    n482_o2_n,
    n482_o2
  );


  buf

  (
    n478_o2_p,
    n478_o2
  );


  not

  (
    n478_o2_n,
    n478_o2
  );


  buf

  (
    n479_o2_p,
    n479_o2
  );


  not

  (
    n479_o2_n,
    n479_o2
  );


  or

  (
    g169_n,
    n852_o2_p,
    n853_o2_p
  );


  or

  (
    g170_n,
    n955_o2_p,
    n956_o2_p
  );


  or

  (
    g171_n,
    n558_o2_p,
    n563_o2_p
  );


  or

  (
    g172_n,
    n262_lo_n,
    n564_o2_n_spl_00
  );


  and

  (
    g173_p,
    n531_o2_p,
    g172_n
  );


  and

  (
    g174_p,
    n598_lo_p,
    n564_o2_p_spl_00
  );


  or

  (
    g175_n,
    n543_o2_n,
    g174_p
  );


  and

  (
    g176_p,
    n550_lo_p,
    n564_o2_p_spl_00
  );


  or

  (
    g176_n,
    n550_lo_n,
    n564_o2_n_spl_00
  );


  and

  (
    g177_p,
    n555_o2_p,
    g176_n
  );


  or

  (
    g177_n,
    n555_o2_n,
    g176_p
  );


  and

  (
    g178_p,
    g175_n_spl_,
    g177_n_spl_
  );


  and

  (
    g179_p,
    n502_lo_p,
    n564_o2_p_spl_01
  );


  or

  (
    g180_n,
    n552_o2_n,
    g179_p
  );


  and

  (
    g181_p,
    n634_lo_p,
    n564_o2_p_spl_01
  );


  or

  (
    g182_n,
    n540_o2_n,
    g181_p
  );


  and

  (
    g183_p,
    g180_n_spl_,
    g182_n
  );


  and

  (
    g184_p,
    g178_p,
    g183_p
  );


  and

  (
    g185_p,
    n358_lo_p,
    n564_o2_p_spl_10
  );


  or

  (
    g185_n,
    n358_lo_n,
    n564_o2_n_spl_0
  );


  and

  (
    g186_p,
    n549_o2_p,
    g185_n
  );


  or

  (
    g186_n,
    n549_o2_n,
    g185_p
  );


  and

  (
    g187_p,
    n454_lo_p,
    n564_o2_p_spl_10
  );


  or

  (
    g187_n,
    n454_lo_n,
    n564_o2_n_spl_1
  );


  and

  (
    g188_p,
    n534_o2_p,
    g187_n
  );


  or

  (
    g188_n,
    n534_o2_n,
    g187_p
  );


  and

  (
    g189_p,
    g186_n_spl_,
    g188_n
  );


  or

  (
    g189_n,
    g186_p_spl_,
    g188_p_spl_
  );


  and

  (
    g190_p,
    n310_lo_p,
    n564_o2_p_spl_11
  );


  or

  (
    g191_n,
    n546_o2_n,
    g190_p
  );


  and

  (
    g192_p,
    n406_lo_p,
    n564_o2_p_spl_11
  );


  or

  (
    g192_n,
    n406_lo_n,
    n564_o2_n_spl_1
  );


  and

  (
    g193_p,
    n537_o2_p,
    g192_n
  );


  or

  (
    g193_n,
    n537_o2_n,
    g192_p
  );


  and

  (
    g194_p,
    g191_n_spl_,
    g193_n_spl_
  );


  and

  (
    g195_p,
    g189_p,
    g194_p
  );


  and

  (
    g196_p,
    g184_p,
    g195_p_spl_
  );


  or

  (
    g197_n,
    g173_p,
    g196_p
  );


  or

  (
    g198_n,
    g180_n_spl_,
    g193_p_spl_
  );


  or

  (
    g199_n,
    g189_n,
    g198_n
  );


  and

  (
    g200_p,
    g191_n_spl_,
    g199_n
  );


  or

  (
    g201_n,
    g188_p_spl_,
    g193_p_spl_
  );


  or

  (
    g202_n,
    g177_n_spl_,
    g201_n
  );


  and

  (
    g203_p,
    g186_n_spl_,
    g202_n
  );


  and

  (
    g204_p,
    g200_p_spl_,
    g203_p
  );


  or

  (
    g205_n,
    g175_n_spl_,
    g177_p
  );


  and

  (
    g206_p,
    g193_n_spl_,
    g205_n
  );


  or

  (
    g207_n,
    g186_p_spl_,
    g206_p
  );


  and

  (
    g208_p,
    g200_p_spl_,
    g207_n
  );


  or

  (
    g209_n,
    n1012_o2_n,
    n530_o2_p
  );


  or

  (
    g210_n,
    n1009_o2_n,
    n548_o2_p
  );


  or

  (
    g211_n,
    n1010_o2_n,
    n536_o2_p
  );


  or

  (
    g212_n,
    n1011_o2_n,
    n539_o2_p
  );


  and

  (
    g213_p,
    lo026_buf_o2_p,
    n528_o2_p_spl_00
  );


  or

  (
    g214_n,
    n510_o2_n,
    g213_p
  );


  and

  (
    g215_p,
    lo074_buf_o2_p,
    n528_o2_p_spl_00
  );


  or

  (
    g216_n,
    n498_o2_n,
    g215_p
  );


  and

  (
    g217_p,
    lo090_buf_o2_p,
    n528_o2_p_spl_0
  );


  or

  (
    g218_n,
    n516_o2_n,
    g217_p
  );


  and

  (
    g219_p,
    lo122_buf_o2_p,
    n528_o2_p_spl_1
  );


  or

  (
    g220_n,
    n507_o2_n,
    g219_p
  );


  and

  (
    g221_p,
    lo106_buf_o2_p,
    n528_o2_p_spl_1
  );


  or

  (
    g222_n,
    n519_o2_n,
    g221_p
  );


  or

  (
    g223_n,
    n1029_o2_n,
    n509_o2_p
  );


  or

  (
    g224_n,
    n1041_o2_n,
    n497_o2_p
  );


  or

  (
    g225_n,
    n1043_o2_n,
    n515_o2_p
  );


  or

  (
    g226_n,
    n1045_o2_n,
    n506_o2_p
  );


  and

  (
    g227_p,
    lo094_buf_o2_p,
    n492_o2_p
  );


  or

  (
    g228_n,
    lo102_buf_o2_n,
    g227_p
  );


  or

  (
    g229_n,
    n547_lo_p_spl_,
    g222_n_spl_
  );


  or

  (
    g230_n,
    n595_lo_p_spl_,
    g220_n_spl_
  );


  or

  (
    g231_n,
    n307_lo_p_spl_,
    g214_n_spl_
  );


  and

  (
    g232_p,
    g230_n,
    g231_n
  );


  and

  (
    g233_p,
    g229_n,
    g232_p
  );


  or

  (
    g234_n,
    n451_lo_p_spl_,
    g216_n_spl_
  );


  or

  (
    g235_n,
    n499_lo_p_spl_,
    g218_n_spl_
  );


  and

  (
    g236_p,
    g234_n,
    g235_n
  );


  or

  (
    g237_n,
    n259_lo_p_spl_,
    g209_n_spl_
  );


  or

  (
    g238_n,
    n631_lo_p_spl_,
    g212_n_spl_
  );


  and

  (
    g239_p,
    g237_n,
    g238_n
  );


  or

  (
    g240_n,
    n403_lo_p_spl_,
    g211_n_spl_
  );


  or

  (
    g241_n,
    n355_lo_p_spl_,
    g210_n_spl_
  );


  and

  (
    g242_p,
    g240_n,
    g241_n
  );


  and

  (
    g243_p,
    g239_p,
    g242_p
  );


  and

  (
    g244_p,
    g236_p,
    g243_p
  );


  or

  (
    g245_n,
    n520_lo_p_spl_,
    g228_n_spl_
  );


  or

  (
    g246_n,
    lo121_buf_o2_p_spl_,
    g226_n_spl_
  );


  or

  (
    g247_n,
    lo025_buf_o2_p_spl_,
    g223_n_spl_
  );


  and

  (
    g248_p,
    g246_n,
    g247_n
  );


  and

  (
    g249_p,
    g245_n,
    g248_p
  );


  or

  (
    g250_n,
    lo073_buf_o2_p_spl_,
    g224_n_spl_
  );


  or

  (
    g251_n,
    lo089_buf_o2_p_spl_,
    g225_n_spl_
  );


  and

  (
    g252_p,
    g250_n,
    g251_n
  );


  or

  (
    g253_n,
    n495_o2_n,
    lo010_buf_o2_p
  );


  or

  (
    g254_n,
    n504_o2_n,
    lo138_buf_o2_p
  );


  and

  (
    g255_p,
    g253_n,
    g254_n
  );


  or

  (
    g256_n,
    n501_o2_n,
    lo058_buf_o2_p
  );


  or

  (
    g257_n,
    n513_o2_n,
    lo042_buf_o2_p
  );


  and

  (
    g258_p,
    g256_n,
    g257_n
  );


  and

  (
    g259_p,
    g255_p,
    g258_p
  );


  and

  (
    g260_p,
    g252_p,
    g259_p
  );


  and

  (
    g261_p,
    lo093_buf_o2_n,
    lo101_buf_o2_p_spl_
  );


  and

  (
    g262_p,
    lo110_buf_o2_n,
    lo118_buf_o2_p_spl_
  );


  and

  (
    g263_p,
    lo002_buf_o2_n,
    lo006_buf_o2_p
  );


  or

  (
    g264_n,
    g262_p,
    g263_p
  );


  or

  (
    g265_n,
    g261_p,
    g264_n
  );


  and

  (
    g266_p,
    lo062_buf_o2_n,
    lo070_buf_o2_p_spl_
  );


  and

  (
    g267_p,
    lo078_buf_o2_n,
    lo086_buf_o2_p_spl_
  );


  or

  (
    g268_n,
    g266_p,
    g267_p
  );


  or

  (
    g269_n,
    n476_o2_p,
    n479_o2_p
  );


  or

  (
    g270_n,
    n482_o2_p,
    n478_o2_p
  );


  or

  (
    g271_n,
    g269_n,
    g270_n
  );


  or

  (
    g272_n,
    g268_n,
    g271_n
  );


  and

  (
    g273_p,
    g233_p_spl_,
    g244_p_spl_
  );


  and

  (
    g274_p,
    g249_p_spl_,
    g260_p_spl_
  );


  or

  (
    g275_n,
    g265_n_spl_,
    g272_n_spl_
  );


  or

  (
    g276_n,
    lo010_buf_o2_n,
    g274_p_spl_00
  );


  or

  (
    g277_n,
    lo042_buf_o2_n,
    g274_p_spl_00
  );


  or

  (
    g278_n,
    lo058_buf_o2_n,
    g274_p_spl_0
  );


  or

  (
    g279_n,
    lo138_buf_o2_n,
    g274_p_spl_1
  );


  and

  (
    g280_p,
    lo014_buf_o2_p,
    g275_n_spl_000
  );


  and

  (
    g281_p,
    lo030_buf_o2_p,
    g275_n_spl_000
  );


  or

  (
    g282_n,
    lo038_buf_o2_n,
    g281_p
  );


  and

  (
    g283_p,
    lo046_buf_o2_p,
    g275_n_spl_00
  );


  or

  (
    g284_n,
    lo054_buf_o2_n,
    g283_p
  );


  and

  (
    g285_p,
    lo126_buf_o2_p,
    g275_n_spl_01
  );


  or

  (
    g286_n,
    lo134_buf_o2_n,
    g285_p
  );


  and

  (
    g287_p,
    lo002_buf_o2_p,
    g275_n_spl_01
  );


  or

  (
    g288_n,
    lo006_buf_o2_n,
    g287_p
  );


  and

  (
    g289_p,
    lo062_buf_o2_p,
    g275_n_spl_10
  );


  and

  (
    g290_p,
    lo078_buf_o2_p,
    g275_n_spl_10
  );


  and

  (
    g291_p,
    lo110_buf_o2_p,
    g275_n_spl_11
  );


  and

  (
    g292_p,
    G4_n,
    G6_p_spl_
  );


  and

  (
    g293_p,
    G8_n,
    G10_p_spl_
  );


  and

  (
    g294_p,
    G12_n,
    G14_p_spl_
  );


  and

  (
    g295_p,
    G32_n,
    G34_p_spl_
  );


  buf

  (
    G426,
    g169_n
  );


  buf

  (
    G427,
    g170_n
  );


  buf

  (
    G428,
    g171_n
  );


  not

  (
    G429,
    g197_n
  );


  not

  (
    G430,
    g195_p_spl_
  );


  not

  (
    G431,
    g204_p
  );


  not

  (
    G432,
    g208_p
  );


  buf

  (
    n856_li008_li008,
    G3_p
  );


  buf

  (
    n880_li016_li016,
    G5_p
  );


  buf

  (
    n883_li017_li017,
    n253_lo_p
  );


  buf

  (
    n886_li018_li018,
    n256_lo_p
  );


  buf

  (
    n889_li019_li019,
    n259_lo_p_spl_
  );


  buf

  (
    n904_li024_li024,
    G7_p
  );


  buf

  (
    n928_li032_li032,
    G9_p
  );


  buf

  (
    n931_li033_li033,
    n301_lo_p
  );


  buf

  (
    n934_li034_li034,
    n304_lo_p
  );


  buf

  (
    n937_li035_li035,
    n307_lo_p_spl_
  );


  buf

  (
    n952_li040_li040,
    G11_p
  );


  buf

  (
    n976_li048_li048,
    G13_p
  );


  buf

  (
    n979_li049_li049,
    n349_lo_p
  );


  buf

  (
    n982_li050_li050,
    n352_lo_p
  );


  buf

  (
    n985_li051_li051,
    n355_lo_p_spl_
  );


  buf

  (
    n1000_li056_li056,
    G15_p
  );


  buf

  (
    n1024_li064_li064,
    G17_p
  );


  buf

  (
    n1027_li065_li065,
    n397_lo_p
  );


  buf

  (
    n1030_li066_li066,
    n400_lo_p
  );


  buf

  (
    n1033_li067_li067,
    n403_lo_p_spl_
  );


  buf

  (
    n1048_li072_li072,
    G19_p
  );


  buf

  (
    n1072_li080_li080,
    G21_p
  );


  buf

  (
    n1075_li081_li081,
    n445_lo_p
  );


  buf

  (
    n1078_li082_li082,
    n448_lo_p
  );


  buf

  (
    n1081_li083_li083,
    n451_lo_p_spl_
  );


  buf

  (
    n1096_li088_li088,
    G23_p
  );


  buf

  (
    n1120_li096_li096,
    G25_p
  );


  buf

  (
    n1123_li097_li097,
    n493_lo_p
  );


  buf

  (
    n1126_li098_li098,
    n496_lo_p
  );


  buf

  (
    n1129_li099_li099,
    n499_lo_p_spl_
  );


  buf

  (
    n1144_li104_li104,
    G27_p
  );


  buf

  (
    n1147_li105_li105,
    n517_lo_p
  );


  buf

  (
    n1168_li112_li112,
    G29_p
  );


  buf

  (
    n1171_li113_li113,
    n541_lo_p
  );


  buf

  (
    n1174_li114_li114,
    n544_lo_p
  );


  buf

  (
    n1177_li115_li115,
    n547_lo_p_spl_
  );


  buf

  (
    n1192_li120_li120,
    G31_p
  );


  buf

  (
    n1216_li128_li128,
    G33_p
  );


  buf

  (
    n1219_li129_li129,
    n589_lo_p
  );


  buf

  (
    n1222_li130_li130,
    n592_lo_p
  );


  buf

  (
    n1225_li131_li131,
    n595_lo_p_spl_
  );


  buf

  (
    n1240_li136_li136,
    G35_p
  );


  buf

  (
    n1252_li140_li140,
    G36_p
  );


  buf

  (
    n1255_li141_li141,
    n625_lo_p
  );


  buf

  (
    n1258_li142_li142,
    n628_lo_p
  );


  buf

  (
    n1261_li143_li143,
    n631_lo_p_spl_
  );


  buf

  (
    n852_i2,
    n961_o2_p
  );


  buf

  (
    n853_i2,
    n223_inv_p
  );


  buf

  (
    n955_i2,
    n522_o2_p
  );


  buf

  (
    n956_i2,
    n298_inv_p
  );


  not

  (
    n531_i2,
    g209_n_spl_
  );


  not

  (
    n549_i2,
    g210_n_spl_
  );


  not

  (
    n537_i2,
    g211_n_spl_
  );


  not

  (
    n540_i2,
    g212_n_spl_
  );


  not

  (
    n546_i2,
    g214_n_spl_
  );


  not

  (
    n534_i2,
    g216_n_spl_
  );


  not

  (
    n552_i2,
    g218_n_spl_
  );


  not

  (
    n543_i2,
    g220_n_spl_
  );


  buf

  (
    n961_i2,
    n486_o2_p
  );


  buf

  (
    n962_i2,
    n304_inv_p
  );


  not

  (
    n555_i2,
    g222_n_spl_
  );


  buf

  (
    n1009_i2,
    n513_o2_p
  );


  buf

  (
    n1010_i2,
    n501_o2_p
  );


  buf

  (
    n1011_i2,
    n504_o2_p
  );


  buf

  (
    n1012_i2,
    n495_o2_p
  );


  buf

  (
    lo026_buf_i2,
    lo025_buf_o2_p_spl_
  );


  buf

  (
    lo074_buf_i2,
    lo073_buf_o2_p_spl_
  );


  buf

  (
    lo090_buf_i2,
    lo089_buf_o2_p_spl_
  );


  buf

  (
    lo122_buf_i2,
    lo121_buf_o2_p_spl_
  );


  not

  (
    n510_i2,
    g223_n_spl_
  );


  not

  (
    n498_i2,
    g224_n_spl_
  );


  not

  (
    n516_i2,
    g225_n_spl_
  );


  not

  (
    n507_i2,
    g226_n_spl_
  );


  buf

  (
    lo106_buf_i2,
    n520_lo_p_spl_
  );


  not

  (
    n519_i2,
    g228_n_spl_
  );


  buf

  (
    n1029_i2,
    lo022_buf_o2_p
  );


  buf

  (
    n1041_i2,
    lo070_buf_o2_p_spl_
  );


  buf

  (
    n1043_i2,
    lo086_buf_o2_p_spl_
  );


  buf

  (
    n1045_i2,
    lo118_buf_o2_p_spl_
  );


  not

  (
    n558_i2,
    g233_p_spl_
  );


  not

  (
    n563_i2,
    g244_p_spl_
  );


  buf

  (
    lo094_buf_i2,
    lo093_buf_o2_p
  );


  buf

  (
    lo102_buf_i2,
    lo101_buf_o2_p_spl_
  );


  not

  (
    n522_i2,
    g249_p_spl_
  );


  not

  (
    n527_i2,
    g260_p_spl_
  );


  buf

  (
    n486_i2,
    g265_n_spl_
  );


  buf

  (
    n491_i2,
    g272_n_spl_
  );


  not

  (
    n564_i2,
    g273_p
  );


  not

  (
    n528_i2,
    g274_p_spl_1
  );


  buf

  (
    n492_i2,
    g275_n_spl_11
  );


  not

  (
    n530_i2,
    g276_n
  );


  not

  (
    n548_i2,
    g277_n
  );


  not

  (
    n536_i2,
    g278_n
  );


  not

  (
    n539_i2,
    g279_n
  );


  buf

  (
    lo025_buf_i2,
    n277_lo_p
  );


  buf

  (
    lo073_buf_i2,
    n421_lo_p
  );


  buf

  (
    lo089_buf_i2,
    n469_lo_p
  );


  buf

  (
    lo121_buf_i2,
    n565_lo_p
  );


  buf

  (
    n509_i2,
    g280_p
  );


  not

  (
    n513_i2,
    g282_n
  );


  not

  (
    n501_i2,
    g284_n
  );


  not

  (
    n504_i2,
    g286_n
  );


  not

  (
    n495_i2,
    g288_n
  );


  buf

  (
    n497_i2,
    g289_p
  );


  buf

  (
    n515_i2,
    g290_p
  );


  buf

  (
    n506_i2,
    g291_p
  );


  buf

  (
    lo010_buf_i2,
    n229_lo_p
  );


  buf

  (
    lo042_buf_i2,
    n325_lo_p
  );


  buf

  (
    lo058_buf_i2,
    n373_lo_p
  );


  buf

  (
    lo138_buf_i2,
    n613_lo_p
  );


  buf

  (
    lo014_buf_i2,
    G4_p
  );


  buf

  (
    lo022_buf_i2,
    G6_p_spl_
  );


  buf

  (
    lo030_buf_i2,
    G8_p
  );


  buf

  (
    lo038_buf_i2,
    G10_p_spl_
  );


  buf

  (
    lo046_buf_i2,
    G12_p
  );


  buf

  (
    lo054_buf_i2,
    G14_p_spl_
  );


  buf

  (
    lo126_buf_i2,
    G32_p
  );


  buf

  (
    lo134_buf_i2,
    G34_p_spl_
  );


  buf

  (
    lo093_buf_i2,
    G24_p
  );


  buf

  (
    lo101_buf_i2,
    G26_p
  );


  buf

  (
    lo002_buf_i2,
    G1_p
  );


  buf

  (
    lo006_buf_i2,
    G2_p
  );


  buf

  (
    lo062_buf_i2,
    G16_p
  );


  buf

  (
    lo070_buf_i2,
    G18_p
  );


  buf

  (
    lo078_buf_i2,
    G20_p
  );


  buf

  (
    lo086_buf_i2,
    G22_p
  );


  buf

  (
    lo110_buf_i2,
    G28_p
  );


  buf

  (
    lo118_buf_i2,
    G30_p
  );


  buf

  (
    n476_i2,
    g292_p
  );


  buf

  (
    n482_i2,
    g293_p
  );


  buf

  (
    n478_i2,
    g294_p
  );


  buf

  (
    n479_i2,
    g295_p
  );


  buf

  (
    n564_o2_n_spl_,
    n564_o2_n
  );


  buf

  (
    n564_o2_n_spl_0,
    n564_o2_n_spl_
  );


  buf

  (
    n564_o2_n_spl_00,
    n564_o2_n_spl_0
  );


  buf

  (
    n564_o2_n_spl_1,
    n564_o2_n_spl_
  );


  buf

  (
    n564_o2_p_spl_,
    n564_o2_p
  );


  buf

  (
    n564_o2_p_spl_0,
    n564_o2_p_spl_
  );


  buf

  (
    n564_o2_p_spl_00,
    n564_o2_p_spl_0
  );


  buf

  (
    n564_o2_p_spl_01,
    n564_o2_p_spl_0
  );


  buf

  (
    n564_o2_p_spl_1,
    n564_o2_p_spl_
  );


  buf

  (
    n564_o2_p_spl_10,
    n564_o2_p_spl_1
  );


  buf

  (
    n564_o2_p_spl_11,
    n564_o2_p_spl_1
  );


  buf

  (
    g175_n_spl_,
    g175_n
  );


  buf

  (
    g177_n_spl_,
    g177_n
  );


  buf

  (
    g180_n_spl_,
    g180_n
  );


  buf

  (
    g186_n_spl_,
    g186_n
  );


  buf

  (
    g186_p_spl_,
    g186_p
  );


  buf

  (
    g188_p_spl_,
    g188_p
  );


  buf

  (
    g191_n_spl_,
    g191_n
  );


  buf

  (
    g193_n_spl_,
    g193_n
  );


  buf

  (
    g195_p_spl_,
    g195_p
  );


  buf

  (
    g193_p_spl_,
    g193_p
  );


  buf

  (
    g200_p_spl_,
    g200_p
  );


  buf

  (
    n528_o2_p_spl_,
    n528_o2_p
  );


  buf

  (
    n528_o2_p_spl_0,
    n528_o2_p_spl_
  );


  buf

  (
    n528_o2_p_spl_00,
    n528_o2_p_spl_0
  );


  buf

  (
    n528_o2_p_spl_1,
    n528_o2_p_spl_
  );


  buf

  (
    n547_lo_p_spl_,
    n547_lo_p
  );


  buf

  (
    g222_n_spl_,
    g222_n
  );


  buf

  (
    n595_lo_p_spl_,
    n595_lo_p
  );


  buf

  (
    g220_n_spl_,
    g220_n
  );


  buf

  (
    n307_lo_p_spl_,
    n307_lo_p
  );


  buf

  (
    g214_n_spl_,
    g214_n
  );


  buf

  (
    n451_lo_p_spl_,
    n451_lo_p
  );


  buf

  (
    g216_n_spl_,
    g216_n
  );


  buf

  (
    n499_lo_p_spl_,
    n499_lo_p
  );


  buf

  (
    g218_n_spl_,
    g218_n
  );


  buf

  (
    n259_lo_p_spl_,
    n259_lo_p
  );


  buf

  (
    g209_n_spl_,
    g209_n
  );


  buf

  (
    n631_lo_p_spl_,
    n631_lo_p
  );


  buf

  (
    g212_n_spl_,
    g212_n
  );


  buf

  (
    n403_lo_p_spl_,
    n403_lo_p
  );


  buf

  (
    g211_n_spl_,
    g211_n
  );


  buf

  (
    n355_lo_p_spl_,
    n355_lo_p
  );


  buf

  (
    g210_n_spl_,
    g210_n
  );


  buf

  (
    n520_lo_p_spl_,
    n520_lo_p
  );


  buf

  (
    g228_n_spl_,
    g228_n
  );


  buf

  (
    lo121_buf_o2_p_spl_,
    lo121_buf_o2_p
  );


  buf

  (
    g226_n_spl_,
    g226_n
  );


  buf

  (
    lo025_buf_o2_p_spl_,
    lo025_buf_o2_p
  );


  buf

  (
    g223_n_spl_,
    g223_n
  );


  buf

  (
    lo073_buf_o2_p_spl_,
    lo073_buf_o2_p
  );


  buf

  (
    g224_n_spl_,
    g224_n
  );


  buf

  (
    lo089_buf_o2_p_spl_,
    lo089_buf_o2_p
  );


  buf

  (
    g225_n_spl_,
    g225_n
  );


  buf

  (
    lo101_buf_o2_p_spl_,
    lo101_buf_o2_p
  );


  buf

  (
    lo118_buf_o2_p_spl_,
    lo118_buf_o2_p
  );


  buf

  (
    lo070_buf_o2_p_spl_,
    lo070_buf_o2_p
  );


  buf

  (
    lo086_buf_o2_p_spl_,
    lo086_buf_o2_p
  );


  buf

  (
    g233_p_spl_,
    g233_p
  );


  buf

  (
    g244_p_spl_,
    g244_p
  );


  buf

  (
    g249_p_spl_,
    g249_p
  );


  buf

  (
    g260_p_spl_,
    g260_p
  );


  buf

  (
    g265_n_spl_,
    g265_n
  );


  buf

  (
    g272_n_spl_,
    g272_n
  );


  buf

  (
    g274_p_spl_,
    g274_p
  );


  buf

  (
    g274_p_spl_0,
    g274_p_spl_
  );


  buf

  (
    g274_p_spl_00,
    g274_p_spl_0
  );


  buf

  (
    g274_p_spl_1,
    g274_p_spl_
  );


  buf

  (
    g275_n_spl_,
    g275_n
  );


  buf

  (
    g275_n_spl_0,
    g275_n_spl_
  );


  buf

  (
    g275_n_spl_00,
    g275_n_spl_0
  );


  buf

  (
    g275_n_spl_000,
    g275_n_spl_00
  );


  buf

  (
    g275_n_spl_01,
    g275_n_spl_0
  );


  buf

  (
    g275_n_spl_1,
    g275_n_spl_
  );


  buf

  (
    g275_n_spl_10,
    g275_n_spl_1
  );


  buf

  (
    g275_n_spl_11,
    g275_n_spl_1
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G34_p_spl_,
    G34_p
  );


endmodule
