
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  n286_lo,
  n298_lo,
  n310_lo,
  n322_lo,
  n334_lo,
  n346_lo,
  n358_lo,
  n370_lo,
  n382_lo,
  n394_lo,
  n406_lo,
  n418_lo,
  n430_lo,
  n442_lo,
  n454_lo,
  n466_lo,
  n478_lo,
  n490_lo,
  n502_lo,
  n514_lo,
  n526_lo,
  n538_lo,
  n550_lo,
  n562_lo,
  n574_lo,
  n586_lo,
  n598_lo,
  n610_lo,
  n622_lo,
  n634_lo,
  n646_lo,
  n658_lo,
  n661_lo,
  n673_lo,
  n685_lo,
  n697_lo,
  n709_lo,
  n721_lo,
  n733_lo,
  n745_lo,
  n757_lo,
  n1248_o2,
  n1249_o2,
  n1250_o2,
  n1251_o2,
  n1252_o2,
  n1253_o2,
  n1254_o2,
  n1255_o2,
  n1207_o2,
  n1208_o2,
  n1209_o2,
  n1210_o2,
  n1211_o2,
  n1212_o2,
  n1213_o2,
  n1214_o2,
  n1215_o2,
  n1216_o2,
  n1217_o2,
  n1218_o2,
  n1219_o2,
  n1220_o2,
  n1221_o2,
  n1222_o2,
  n1223_o2,
  n1224_o2,
  n1225_o2,
  n1226_o2,
  n1227_o2,
  n1228_o2,
  n1229_o2,
  n1230_o2,
  n1231_o2,
  n1232_o2,
  n1233_o2,
  n1234_o2,
  n1235_o2,
  n1236_o2,
  n1237_o2,
  n1238_o2,
  G374_o2,
  G376_o2,
  G370_o2,
  G372_o2,
  G373_o2,
  G377_o2,
  G371_o2,
  G375_o2,
  G354_o2,
  G356_o2,
  G350_o2,
  G352_o2,
  G353_o2,
  G357_o2,
  G351_o2,
  G355_o2,
  G386_o2,
  G391_o2,
  n283_lo_buf_o2,
  n295_lo_buf_o2,
  n307_lo_buf_o2,
  n319_lo_buf_o2,
  n331_lo_buf_o2,
  n343_lo_buf_o2,
  n355_lo_buf_o2,
  n367_lo_buf_o2,
  n379_lo_buf_o2,
  n391_lo_buf_o2,
  n403_lo_buf_o2,
  n415_lo_buf_o2,
  n427_lo_buf_o2,
  n439_lo_buf_o2,
  n451_lo_buf_o2,
  n463_lo_buf_o2,
  n475_lo_buf_o2,
  n487_lo_buf_o2,
  n499_lo_buf_o2,
  n511_lo_buf_o2,
  n523_lo_buf_o2,
  n535_lo_buf_o2,
  n547_lo_buf_o2,
  n559_lo_buf_o2,
  n571_lo_buf_o2,
  n583_lo_buf_o2,
  n595_lo_buf_o2,
  n607_lo_buf_o2,
  n619_lo_buf_o2,
  n631_lo_buf_o2,
  n643_lo_buf_o2,
  n655_lo_buf_o2,
  G234_o2,
  G247_o2,
  G260_o2,
  G273_o2,
  G286_o2,
  G299_o2,
  G312_o2,
  G325_o2,
  n667_lo_buf_o2,
  n679_lo_buf_o2,
  n691_lo_buf_o2,
  n703_lo_buf_o2,
  n715_lo_buf_o2,
  n727_lo_buf_o2,
  n739_lo_buf_o2,
  n751_lo_buf_o2,
  n763_lo_buf_o2,
  G186_o2,
  G189_o2,
  G192_o2,
  G195_o2,
  G198_o2,
  G201_o2,
  G204_o2,
  G207_o2,
  n280_lo_buf_o2,
  n292_lo_buf_o2,
  n304_lo_buf_o2,
  n316_lo_buf_o2,
  n328_lo_buf_o2,
  n340_lo_buf_o2,
  n352_lo_buf_o2,
  n364_lo_buf_o2,
  n376_lo_buf_o2,
  n388_lo_buf_o2,
  n400_lo_buf_o2,
  n412_lo_buf_o2,
  n424_lo_buf_o2,
  n436_lo_buf_o2,
  n448_lo_buf_o2,
  n460_lo_buf_o2,
  n472_lo_buf_o2,
  n484_lo_buf_o2,
  n496_lo_buf_o2,
  n508_lo_buf_o2,
  n520_lo_buf_o2,
  n532_lo_buf_o2,
  n544_lo_buf_o2,
  n556_lo_buf_o2,
  n568_lo_buf_o2,
  n580_lo_buf_o2,
  n592_lo_buf_o2,
  n604_lo_buf_o2,
  n616_lo_buf_o2,
  n628_lo_buf_o2,
  n640_lo_buf_o2,
  n652_lo_buf_o2,
  G468,
  G469,
  G470,
  G471,
  G472,
  G473,
  G474,
  G475,
  G476,
  G477,
  G478,
  G479,
  G480,
  G481,
  G482,
  G483,
  G484,
  G485,
  G486,
  G487,
  G488,
  G489,
  G490,
  G491,
  G492,
  G493,
  G494,
  G495,
  G496,
  G497,
  G498,
  G499,
  n286_li,
  n298_li,
  n310_li,
  n322_li,
  n334_li,
  n346_li,
  n358_li,
  n370_li,
  n382_li,
  n394_li,
  n406_li,
  n418_li,
  n430_li,
  n442_li,
  n454_li,
  n466_li,
  n478_li,
  n490_li,
  n502_li,
  n514_li,
  n526_li,
  n538_li,
  n550_li,
  n562_li,
  n574_li,
  n586_li,
  n598_li,
  n610_li,
  n622_li,
  n634_li,
  n646_li,
  n658_li,
  n661_li,
  n673_li,
  n685_li,
  n697_li,
  n709_li,
  n721_li,
  n733_li,
  n745_li,
  n757_li,
  n1248_i2,
  n1249_i2,
  n1250_i2,
  n1251_i2,
  n1252_i2,
  n1253_i2,
  n1254_i2,
  n1255_i2,
  n1207_i2,
  n1208_i2,
  n1209_i2,
  n1210_i2,
  n1211_i2,
  n1212_i2,
  n1213_i2,
  n1214_i2,
  n1215_i2,
  n1216_i2,
  n1217_i2,
  n1218_i2,
  n1219_i2,
  n1220_i2,
  n1221_i2,
  n1222_i2,
  n1223_i2,
  n1224_i2,
  n1225_i2,
  n1226_i2,
  n1227_i2,
  n1228_i2,
  n1229_i2,
  n1230_i2,
  n1231_i2,
  n1232_i2,
  n1233_i2,
  n1234_i2,
  n1235_i2,
  n1236_i2,
  n1237_i2,
  n1238_i2,
  G374_i2,
  G376_i2,
  G370_i2,
  G372_i2,
  G373_i2,
  G377_i2,
  G371_i2,
  G375_i2,
  G354_i2,
  G356_i2,
  G350_i2,
  G352_i2,
  G353_i2,
  G357_i2,
  G351_i2,
  G355_i2,
  G386_i2,
  G391_i2,
  n283_lo_buf_i2,
  n295_lo_buf_i2,
  n307_lo_buf_i2,
  n319_lo_buf_i2,
  n331_lo_buf_i2,
  n343_lo_buf_i2,
  n355_lo_buf_i2,
  n367_lo_buf_i2,
  n379_lo_buf_i2,
  n391_lo_buf_i2,
  n403_lo_buf_i2,
  n415_lo_buf_i2,
  n427_lo_buf_i2,
  n439_lo_buf_i2,
  n451_lo_buf_i2,
  n463_lo_buf_i2,
  n475_lo_buf_i2,
  n487_lo_buf_i2,
  n499_lo_buf_i2,
  n511_lo_buf_i2,
  n523_lo_buf_i2,
  n535_lo_buf_i2,
  n547_lo_buf_i2,
  n559_lo_buf_i2,
  n571_lo_buf_i2,
  n583_lo_buf_i2,
  n595_lo_buf_i2,
  n607_lo_buf_i2,
  n619_lo_buf_i2,
  n631_lo_buf_i2,
  n643_lo_buf_i2,
  n655_lo_buf_i2,
  G234_i2,
  G247_i2,
  G260_i2,
  G273_i2,
  G286_i2,
  G299_i2,
  G312_i2,
  G325_i2,
  n667_lo_buf_i2,
  n679_lo_buf_i2,
  n691_lo_buf_i2,
  n703_lo_buf_i2,
  n715_lo_buf_i2,
  n727_lo_buf_i2,
  n739_lo_buf_i2,
  n751_lo_buf_i2,
  n763_lo_buf_i2,
  G186_i2,
  G189_i2,
  G192_i2,
  G195_i2,
  G198_i2,
  G201_i2,
  G204_i2,
  G207_i2,
  n280_lo_buf_i2,
  n292_lo_buf_i2,
  n304_lo_buf_i2,
  n316_lo_buf_i2,
  n328_lo_buf_i2,
  n340_lo_buf_i2,
  n352_lo_buf_i2,
  n364_lo_buf_i2,
  n376_lo_buf_i2,
  n388_lo_buf_i2,
  n400_lo_buf_i2,
  n412_lo_buf_i2,
  n424_lo_buf_i2,
  n436_lo_buf_i2,
  n448_lo_buf_i2,
  n460_lo_buf_i2,
  n472_lo_buf_i2,
  n484_lo_buf_i2,
  n496_lo_buf_i2,
  n508_lo_buf_i2,
  n520_lo_buf_i2,
  n532_lo_buf_i2,
  n544_lo_buf_i2,
  n556_lo_buf_i2,
  n568_lo_buf_i2,
  n580_lo_buf_i2,
  n592_lo_buf_i2,
  n604_lo_buf_i2,
  n616_lo_buf_i2,
  n628_lo_buf_i2,
  n640_lo_buf_i2,
  n652_lo_buf_i2
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;input n286_lo;input n298_lo;input n310_lo;input n322_lo;input n334_lo;input n346_lo;input n358_lo;input n370_lo;input n382_lo;input n394_lo;input n406_lo;input n418_lo;input n430_lo;input n442_lo;input n454_lo;input n466_lo;input n478_lo;input n490_lo;input n502_lo;input n514_lo;input n526_lo;input n538_lo;input n550_lo;input n562_lo;input n574_lo;input n586_lo;input n598_lo;input n610_lo;input n622_lo;input n634_lo;input n646_lo;input n658_lo;input n661_lo;input n673_lo;input n685_lo;input n697_lo;input n709_lo;input n721_lo;input n733_lo;input n745_lo;input n757_lo;input n1248_o2;input n1249_o2;input n1250_o2;input n1251_o2;input n1252_o2;input n1253_o2;input n1254_o2;input n1255_o2;input n1207_o2;input n1208_o2;input n1209_o2;input n1210_o2;input n1211_o2;input n1212_o2;input n1213_o2;input n1214_o2;input n1215_o2;input n1216_o2;input n1217_o2;input n1218_o2;input n1219_o2;input n1220_o2;input n1221_o2;input n1222_o2;input n1223_o2;input n1224_o2;input n1225_o2;input n1226_o2;input n1227_o2;input n1228_o2;input n1229_o2;input n1230_o2;input n1231_o2;input n1232_o2;input n1233_o2;input n1234_o2;input n1235_o2;input n1236_o2;input n1237_o2;input n1238_o2;input G374_o2;input G376_o2;input G370_o2;input G372_o2;input G373_o2;input G377_o2;input G371_o2;input G375_o2;input G354_o2;input G356_o2;input G350_o2;input G352_o2;input G353_o2;input G357_o2;input G351_o2;input G355_o2;input G386_o2;input G391_o2;input n283_lo_buf_o2;input n295_lo_buf_o2;input n307_lo_buf_o2;input n319_lo_buf_o2;input n331_lo_buf_o2;input n343_lo_buf_o2;input n355_lo_buf_o2;input n367_lo_buf_o2;input n379_lo_buf_o2;input n391_lo_buf_o2;input n403_lo_buf_o2;input n415_lo_buf_o2;input n427_lo_buf_o2;input n439_lo_buf_o2;input n451_lo_buf_o2;input n463_lo_buf_o2;input n475_lo_buf_o2;input n487_lo_buf_o2;input n499_lo_buf_o2;input n511_lo_buf_o2;input n523_lo_buf_o2;input n535_lo_buf_o2;input n547_lo_buf_o2;input n559_lo_buf_o2;input n571_lo_buf_o2;input n583_lo_buf_o2;input n595_lo_buf_o2;input n607_lo_buf_o2;input n619_lo_buf_o2;input n631_lo_buf_o2;input n643_lo_buf_o2;input n655_lo_buf_o2;input G234_o2;input G247_o2;input G260_o2;input G273_o2;input G286_o2;input G299_o2;input G312_o2;input G325_o2;input n667_lo_buf_o2;input n679_lo_buf_o2;input n691_lo_buf_o2;input n703_lo_buf_o2;input n715_lo_buf_o2;input n727_lo_buf_o2;input n739_lo_buf_o2;input n751_lo_buf_o2;input n763_lo_buf_o2;input G186_o2;input G189_o2;input G192_o2;input G195_o2;input G198_o2;input G201_o2;input G204_o2;input G207_o2;input n280_lo_buf_o2;input n292_lo_buf_o2;input n304_lo_buf_o2;input n316_lo_buf_o2;input n328_lo_buf_o2;input n340_lo_buf_o2;input n352_lo_buf_o2;input n364_lo_buf_o2;input n376_lo_buf_o2;input n388_lo_buf_o2;input n400_lo_buf_o2;input n412_lo_buf_o2;input n424_lo_buf_o2;input n436_lo_buf_o2;input n448_lo_buf_o2;input n460_lo_buf_o2;input n472_lo_buf_o2;input n484_lo_buf_o2;input n496_lo_buf_o2;input n508_lo_buf_o2;input n520_lo_buf_o2;input n532_lo_buf_o2;input n544_lo_buf_o2;input n556_lo_buf_o2;input n568_lo_buf_o2;input n580_lo_buf_o2;input n592_lo_buf_o2;input n604_lo_buf_o2;input n616_lo_buf_o2;input n628_lo_buf_o2;input n640_lo_buf_o2;input n652_lo_buf_o2;
  output G468;output G469;output G470;output G471;output G472;output G473;output G474;output G475;output G476;output G477;output G478;output G479;output G480;output G481;output G482;output G483;output G484;output G485;output G486;output G487;output G488;output G489;output G490;output G491;output G492;output G493;output G494;output G495;output G496;output G497;output G498;output G499;output n286_li;output n298_li;output n310_li;output n322_li;output n334_li;output n346_li;output n358_li;output n370_li;output n382_li;output n394_li;output n406_li;output n418_li;output n430_li;output n442_li;output n454_li;output n466_li;output n478_li;output n490_li;output n502_li;output n514_li;output n526_li;output n538_li;output n550_li;output n562_li;output n574_li;output n586_li;output n598_li;output n610_li;output n622_li;output n634_li;output n646_li;output n658_li;output n661_li;output n673_li;output n685_li;output n697_li;output n709_li;output n721_li;output n733_li;output n745_li;output n757_li;output n1248_i2;output n1249_i2;output n1250_i2;output n1251_i2;output n1252_i2;output n1253_i2;output n1254_i2;output n1255_i2;output n1207_i2;output n1208_i2;output n1209_i2;output n1210_i2;output n1211_i2;output n1212_i2;output n1213_i2;output n1214_i2;output n1215_i2;output n1216_i2;output n1217_i2;output n1218_i2;output n1219_i2;output n1220_i2;output n1221_i2;output n1222_i2;output n1223_i2;output n1224_i2;output n1225_i2;output n1226_i2;output n1227_i2;output n1228_i2;output n1229_i2;output n1230_i2;output n1231_i2;output n1232_i2;output n1233_i2;output n1234_i2;output n1235_i2;output n1236_i2;output n1237_i2;output n1238_i2;output G374_i2;output G376_i2;output G370_i2;output G372_i2;output G373_i2;output G377_i2;output G371_i2;output G375_i2;output G354_i2;output G356_i2;output G350_i2;output G352_i2;output G353_i2;output G357_i2;output G351_i2;output G355_i2;output G386_i2;output G391_i2;output n283_lo_buf_i2;output n295_lo_buf_i2;output n307_lo_buf_i2;output n319_lo_buf_i2;output n331_lo_buf_i2;output n343_lo_buf_i2;output n355_lo_buf_i2;output n367_lo_buf_i2;output n379_lo_buf_i2;output n391_lo_buf_i2;output n403_lo_buf_i2;output n415_lo_buf_i2;output n427_lo_buf_i2;output n439_lo_buf_i2;output n451_lo_buf_i2;output n463_lo_buf_i2;output n475_lo_buf_i2;output n487_lo_buf_i2;output n499_lo_buf_i2;output n511_lo_buf_i2;output n523_lo_buf_i2;output n535_lo_buf_i2;output n547_lo_buf_i2;output n559_lo_buf_i2;output n571_lo_buf_i2;output n583_lo_buf_i2;output n595_lo_buf_i2;output n607_lo_buf_i2;output n619_lo_buf_i2;output n631_lo_buf_i2;output n643_lo_buf_i2;output n655_lo_buf_i2;output G234_i2;output G247_i2;output G260_i2;output G273_i2;output G286_i2;output G299_i2;output G312_i2;output G325_i2;output n667_lo_buf_i2;output n679_lo_buf_i2;output n691_lo_buf_i2;output n703_lo_buf_i2;output n715_lo_buf_i2;output n727_lo_buf_i2;output n739_lo_buf_i2;output n751_lo_buf_i2;output n763_lo_buf_i2;output G186_i2;output G189_i2;output G192_i2;output G195_i2;output G198_i2;output G201_i2;output G204_i2;output G207_i2;output n280_lo_buf_i2;output n292_lo_buf_i2;output n304_lo_buf_i2;output n316_lo_buf_i2;output n328_lo_buf_i2;output n340_lo_buf_i2;output n352_lo_buf_i2;output n364_lo_buf_i2;output n376_lo_buf_i2;output n388_lo_buf_i2;output n400_lo_buf_i2;output n412_lo_buf_i2;output n424_lo_buf_i2;output n436_lo_buf_i2;output n448_lo_buf_i2;output n460_lo_buf_i2;output n472_lo_buf_i2;output n484_lo_buf_i2;output n496_lo_buf_i2;output n508_lo_buf_i2;output n520_lo_buf_i2;output n532_lo_buf_i2;output n544_lo_buf_i2;output n556_lo_buf_i2;output n568_lo_buf_i2;output n580_lo_buf_i2;output n592_lo_buf_i2;output n604_lo_buf_i2;output n616_lo_buf_i2;output n628_lo_buf_i2;output n640_lo_buf_i2;output n652_lo_buf_i2;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire G33_p;
  wire G33_n;
  wire G34_p;
  wire G34_n;
  wire G35_p;
  wire G35_n;
  wire G36_p;
  wire G36_n;
  wire G37_p;
  wire G37_n;
  wire G38_p;
  wire G38_n;
  wire G39_p;
  wire G39_n;
  wire G40_p;
  wire G40_n;
  wire G41_p;
  wire G41_n;
  wire n286_lo_p;
  wire n286_lo_n;
  wire n298_lo_p;
  wire n298_lo_n;
  wire n310_lo_p;
  wire n310_lo_n;
  wire n322_lo_p;
  wire n322_lo_n;
  wire n334_lo_p;
  wire n334_lo_n;
  wire n346_lo_p;
  wire n346_lo_n;
  wire n358_lo_p;
  wire n358_lo_n;
  wire n370_lo_p;
  wire n370_lo_n;
  wire n382_lo_p;
  wire n382_lo_n;
  wire n394_lo_p;
  wire n394_lo_n;
  wire n406_lo_p;
  wire n406_lo_n;
  wire n418_lo_p;
  wire n418_lo_n;
  wire n430_lo_p;
  wire n430_lo_n;
  wire n442_lo_p;
  wire n442_lo_n;
  wire n454_lo_p;
  wire n454_lo_n;
  wire n466_lo_p;
  wire n466_lo_n;
  wire n478_lo_p;
  wire n478_lo_n;
  wire n490_lo_p;
  wire n490_lo_n;
  wire n502_lo_p;
  wire n502_lo_n;
  wire n514_lo_p;
  wire n514_lo_n;
  wire n526_lo_p;
  wire n526_lo_n;
  wire n538_lo_p;
  wire n538_lo_n;
  wire n550_lo_p;
  wire n550_lo_n;
  wire n562_lo_p;
  wire n562_lo_n;
  wire n574_lo_p;
  wire n574_lo_n;
  wire n586_lo_p;
  wire n586_lo_n;
  wire n598_lo_p;
  wire n598_lo_n;
  wire n610_lo_p;
  wire n610_lo_n;
  wire n622_lo_p;
  wire n622_lo_n;
  wire n634_lo_p;
  wire n634_lo_n;
  wire n646_lo_p;
  wire n646_lo_n;
  wire n658_lo_p;
  wire n658_lo_n;
  wire n661_lo_p;
  wire n661_lo_n;
  wire n673_lo_p;
  wire n673_lo_n;
  wire n685_lo_p;
  wire n685_lo_n;
  wire n697_lo_p;
  wire n697_lo_n;
  wire n709_lo_p;
  wire n709_lo_n;
  wire n721_lo_p;
  wire n721_lo_n;
  wire n733_lo_p;
  wire n733_lo_n;
  wire n745_lo_p;
  wire n745_lo_n;
  wire n757_lo_p;
  wire n757_lo_n;
  wire n1248_o2_p;
  wire n1248_o2_n;
  wire n1249_o2_p;
  wire n1249_o2_n;
  wire n1250_o2_p;
  wire n1250_o2_n;
  wire n1251_o2_p;
  wire n1251_o2_n;
  wire n1252_o2_p;
  wire n1252_o2_n;
  wire n1253_o2_p;
  wire n1253_o2_n;
  wire n1254_o2_p;
  wire n1254_o2_n;
  wire n1255_o2_p;
  wire n1255_o2_n;
  wire n1207_o2_p;
  wire n1207_o2_n;
  wire n1208_o2_p;
  wire n1208_o2_n;
  wire n1209_o2_p;
  wire n1209_o2_n;
  wire n1210_o2_p;
  wire n1210_o2_n;
  wire n1211_o2_p;
  wire n1211_o2_n;
  wire n1212_o2_p;
  wire n1212_o2_n;
  wire n1213_o2_p;
  wire n1213_o2_n;
  wire n1214_o2_p;
  wire n1214_o2_n;
  wire n1215_o2_p;
  wire n1215_o2_n;
  wire n1216_o2_p;
  wire n1216_o2_n;
  wire n1217_o2_p;
  wire n1217_o2_n;
  wire n1218_o2_p;
  wire n1218_o2_n;
  wire n1219_o2_p;
  wire n1219_o2_n;
  wire n1220_o2_p;
  wire n1220_o2_n;
  wire n1221_o2_p;
  wire n1221_o2_n;
  wire n1222_o2_p;
  wire n1222_o2_n;
  wire n1223_o2_p;
  wire n1223_o2_n;
  wire n1224_o2_p;
  wire n1224_o2_n;
  wire n1225_o2_p;
  wire n1225_o2_n;
  wire n1226_o2_p;
  wire n1226_o2_n;
  wire n1227_o2_p;
  wire n1227_o2_n;
  wire n1228_o2_p;
  wire n1228_o2_n;
  wire n1229_o2_p;
  wire n1229_o2_n;
  wire n1230_o2_p;
  wire n1230_o2_n;
  wire n1231_o2_p;
  wire n1231_o2_n;
  wire n1232_o2_p;
  wire n1232_o2_n;
  wire n1233_o2_p;
  wire n1233_o2_n;
  wire n1234_o2_p;
  wire n1234_o2_n;
  wire n1235_o2_p;
  wire n1235_o2_n;
  wire n1236_o2_p;
  wire n1236_o2_n;
  wire n1237_o2_p;
  wire n1237_o2_n;
  wire n1238_o2_p;
  wire n1238_o2_n;
  wire G374_o2_p;
  wire G374_o2_n;
  wire G376_o2_p;
  wire G376_o2_n;
  wire G370_o2_p;
  wire G370_o2_n;
  wire G372_o2_p;
  wire G372_o2_n;
  wire G373_o2_p;
  wire G373_o2_n;
  wire G377_o2_p;
  wire G377_o2_n;
  wire G371_o2_p;
  wire G371_o2_n;
  wire G375_o2_p;
  wire G375_o2_n;
  wire G354_o2_p;
  wire G354_o2_n;
  wire G356_o2_p;
  wire G356_o2_n;
  wire G350_o2_p;
  wire G350_o2_n;
  wire G352_o2_p;
  wire G352_o2_n;
  wire G353_o2_p;
  wire G353_o2_n;
  wire G357_o2_p;
  wire G357_o2_n;
  wire G351_o2_p;
  wire G351_o2_n;
  wire G355_o2_p;
  wire G355_o2_n;
  wire G386_o2_p;
  wire G386_o2_n;
  wire G391_o2_p;
  wire G391_o2_n;
  wire n283_lo_buf_o2_p;
  wire n283_lo_buf_o2_n;
  wire n295_lo_buf_o2_p;
  wire n295_lo_buf_o2_n;
  wire n307_lo_buf_o2_p;
  wire n307_lo_buf_o2_n;
  wire n319_lo_buf_o2_p;
  wire n319_lo_buf_o2_n;
  wire n331_lo_buf_o2_p;
  wire n331_lo_buf_o2_n;
  wire n343_lo_buf_o2_p;
  wire n343_lo_buf_o2_n;
  wire n355_lo_buf_o2_p;
  wire n355_lo_buf_o2_n;
  wire n367_lo_buf_o2_p;
  wire n367_lo_buf_o2_n;
  wire n379_lo_buf_o2_p;
  wire n379_lo_buf_o2_n;
  wire n391_lo_buf_o2_p;
  wire n391_lo_buf_o2_n;
  wire n403_lo_buf_o2_p;
  wire n403_lo_buf_o2_n;
  wire n415_lo_buf_o2_p;
  wire n415_lo_buf_o2_n;
  wire n427_lo_buf_o2_p;
  wire n427_lo_buf_o2_n;
  wire n439_lo_buf_o2_p;
  wire n439_lo_buf_o2_n;
  wire n451_lo_buf_o2_p;
  wire n451_lo_buf_o2_n;
  wire n463_lo_buf_o2_p;
  wire n463_lo_buf_o2_n;
  wire n475_lo_buf_o2_p;
  wire n475_lo_buf_o2_n;
  wire n487_lo_buf_o2_p;
  wire n487_lo_buf_o2_n;
  wire n499_lo_buf_o2_p;
  wire n499_lo_buf_o2_n;
  wire n511_lo_buf_o2_p;
  wire n511_lo_buf_o2_n;
  wire n523_lo_buf_o2_p;
  wire n523_lo_buf_o2_n;
  wire n535_lo_buf_o2_p;
  wire n535_lo_buf_o2_n;
  wire n547_lo_buf_o2_p;
  wire n547_lo_buf_o2_n;
  wire n559_lo_buf_o2_p;
  wire n559_lo_buf_o2_n;
  wire n571_lo_buf_o2_p;
  wire n571_lo_buf_o2_n;
  wire n583_lo_buf_o2_p;
  wire n583_lo_buf_o2_n;
  wire n595_lo_buf_o2_p;
  wire n595_lo_buf_o2_n;
  wire n607_lo_buf_o2_p;
  wire n607_lo_buf_o2_n;
  wire n619_lo_buf_o2_p;
  wire n619_lo_buf_o2_n;
  wire n631_lo_buf_o2_p;
  wire n631_lo_buf_o2_n;
  wire n643_lo_buf_o2_p;
  wire n643_lo_buf_o2_n;
  wire n655_lo_buf_o2_p;
  wire n655_lo_buf_o2_n;
  wire G234_o2_p;
  wire G234_o2_n;
  wire G247_o2_p;
  wire G247_o2_n;
  wire G260_o2_p;
  wire G260_o2_n;
  wire G273_o2_p;
  wire G273_o2_n;
  wire G286_o2_p;
  wire G286_o2_n;
  wire G299_o2_p;
  wire G299_o2_n;
  wire G312_o2_p;
  wire G312_o2_n;
  wire G325_o2_p;
  wire G325_o2_n;
  wire n667_lo_buf_o2_p;
  wire n667_lo_buf_o2_n;
  wire n679_lo_buf_o2_p;
  wire n679_lo_buf_o2_n;
  wire n691_lo_buf_o2_p;
  wire n691_lo_buf_o2_n;
  wire n703_lo_buf_o2_p;
  wire n703_lo_buf_o2_n;
  wire n715_lo_buf_o2_p;
  wire n715_lo_buf_o2_n;
  wire n727_lo_buf_o2_p;
  wire n727_lo_buf_o2_n;
  wire n739_lo_buf_o2_p;
  wire n739_lo_buf_o2_n;
  wire n751_lo_buf_o2_p;
  wire n751_lo_buf_o2_n;
  wire n763_lo_buf_o2_p;
  wire n763_lo_buf_o2_n;
  wire G186_o2_p;
  wire G186_o2_n;
  wire G189_o2_p;
  wire G189_o2_n;
  wire G192_o2_p;
  wire G192_o2_n;
  wire G195_o2_p;
  wire G195_o2_n;
  wire G198_o2_p;
  wire G198_o2_n;
  wire G201_o2_p;
  wire G201_o2_n;
  wire G204_o2_p;
  wire G204_o2_n;
  wire G207_o2_p;
  wire G207_o2_n;
  wire n280_lo_buf_o2_p;
  wire n280_lo_buf_o2_n;
  wire n292_lo_buf_o2_p;
  wire n292_lo_buf_o2_n;
  wire n304_lo_buf_o2_p;
  wire n304_lo_buf_o2_n;
  wire n316_lo_buf_o2_p;
  wire n316_lo_buf_o2_n;
  wire n328_lo_buf_o2_p;
  wire n328_lo_buf_o2_n;
  wire n340_lo_buf_o2_p;
  wire n340_lo_buf_o2_n;
  wire n352_lo_buf_o2_p;
  wire n352_lo_buf_o2_n;
  wire n364_lo_buf_o2_p;
  wire n364_lo_buf_o2_n;
  wire n376_lo_buf_o2_p;
  wire n376_lo_buf_o2_n;
  wire n388_lo_buf_o2_p;
  wire n388_lo_buf_o2_n;
  wire n400_lo_buf_o2_p;
  wire n400_lo_buf_o2_n;
  wire n412_lo_buf_o2_p;
  wire n412_lo_buf_o2_n;
  wire n424_lo_buf_o2_p;
  wire n424_lo_buf_o2_n;
  wire n436_lo_buf_o2_p;
  wire n436_lo_buf_o2_n;
  wire n448_lo_buf_o2_p;
  wire n448_lo_buf_o2_n;
  wire n460_lo_buf_o2_p;
  wire n460_lo_buf_o2_n;
  wire n472_lo_buf_o2_p;
  wire n472_lo_buf_o2_n;
  wire n484_lo_buf_o2_p;
  wire n484_lo_buf_o2_n;
  wire n496_lo_buf_o2_p;
  wire n496_lo_buf_o2_n;
  wire n508_lo_buf_o2_p;
  wire n508_lo_buf_o2_n;
  wire n520_lo_buf_o2_p;
  wire n520_lo_buf_o2_n;
  wire n532_lo_buf_o2_p;
  wire n532_lo_buf_o2_n;
  wire n544_lo_buf_o2_p;
  wire n544_lo_buf_o2_n;
  wire n556_lo_buf_o2_p;
  wire n556_lo_buf_o2_n;
  wire n568_lo_buf_o2_p;
  wire n568_lo_buf_o2_n;
  wire n580_lo_buf_o2_p;
  wire n580_lo_buf_o2_n;
  wire n592_lo_buf_o2_p;
  wire n592_lo_buf_o2_n;
  wire n604_lo_buf_o2_p;
  wire n604_lo_buf_o2_n;
  wire n616_lo_buf_o2_p;
  wire n616_lo_buf_o2_n;
  wire n628_lo_buf_o2_p;
  wire n628_lo_buf_o2_n;
  wire n640_lo_buf_o2_p;
  wire n640_lo_buf_o2_n;
  wire n652_lo_buf_o2_p;
  wire n652_lo_buf_o2_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire n1252_o2_p_spl_;
  wire n1252_o2_p_spl_0;
  wire n1252_o2_p_spl_00;
  wire n1252_o2_p_spl_01;
  wire n1252_o2_p_spl_1;
  wire n1252_o2_n_spl_;
  wire n1252_o2_n_spl_0;
  wire n1252_o2_n_spl_00;
  wire n1252_o2_n_spl_01;
  wire n1252_o2_n_spl_1;
  wire n1254_o2_p_spl_;
  wire n1254_o2_p_spl_0;
  wire n1254_o2_p_spl_00;
  wire n1254_o2_p_spl_01;
  wire n1254_o2_p_spl_1;
  wire n1254_o2_n_spl_;
  wire n1254_o2_n_spl_0;
  wire n1254_o2_n_spl_00;
  wire n1254_o2_n_spl_01;
  wire n1254_o2_n_spl_1;
  wire G386_o2_p_spl_;
  wire G386_o2_p_spl_0;
  wire G386_o2_p_spl_1;
  wire G386_o2_n_spl_;
  wire G386_o2_n_spl_0;
  wire G386_o2_n_spl_1;
  wire g233_p_spl_;
  wire g233_p_spl_0;
  wire g233_p_spl_1;
  wire n1248_o2_p_spl_;
  wire n1248_o2_p_spl_0;
  wire n1248_o2_p_spl_00;
  wire n1248_o2_p_spl_01;
  wire n1248_o2_p_spl_1;
  wire g233_n_spl_;
  wire g233_n_spl_0;
  wire g233_n_spl_1;
  wire n1248_o2_n_spl_;
  wire n1248_o2_n_spl_0;
  wire n1248_o2_n_spl_00;
  wire n1248_o2_n_spl_01;
  wire n1248_o2_n_spl_1;
  wire n1249_o2_p_spl_;
  wire n1249_o2_p_spl_0;
  wire n1249_o2_p_spl_00;
  wire n1249_o2_p_spl_01;
  wire n1249_o2_p_spl_1;
  wire n1249_o2_n_spl_;
  wire n1249_o2_n_spl_0;
  wire n1249_o2_n_spl_00;
  wire n1249_o2_n_spl_01;
  wire n1249_o2_n_spl_1;
  wire n1250_o2_p_spl_;
  wire n1250_o2_p_spl_0;
  wire n1250_o2_p_spl_00;
  wire n1250_o2_p_spl_01;
  wire n1250_o2_p_spl_1;
  wire n1250_o2_n_spl_;
  wire n1250_o2_n_spl_0;
  wire n1250_o2_n_spl_00;
  wire n1250_o2_n_spl_01;
  wire n1250_o2_n_spl_1;
  wire n1251_o2_p_spl_;
  wire n1251_o2_p_spl_0;
  wire n1251_o2_p_spl_00;
  wire n1251_o2_p_spl_01;
  wire n1251_o2_p_spl_1;
  wire n1251_o2_n_spl_;
  wire n1251_o2_n_spl_0;
  wire n1251_o2_n_spl_00;
  wire n1251_o2_n_spl_01;
  wire n1251_o2_n_spl_1;
  wire n1255_o2_p_spl_;
  wire n1255_o2_p_spl_0;
  wire n1255_o2_p_spl_00;
  wire n1255_o2_p_spl_01;
  wire n1255_o2_p_spl_1;
  wire n1255_o2_n_spl_;
  wire n1255_o2_n_spl_0;
  wire n1255_o2_n_spl_00;
  wire n1255_o2_n_spl_01;
  wire n1255_o2_n_spl_1;
  wire g253_p_spl_;
  wire g253_p_spl_0;
  wire g253_p_spl_1;
  wire g253_n_spl_;
  wire g253_n_spl_0;
  wire g253_n_spl_1;
  wire n1253_o2_p_spl_;
  wire n1253_o2_p_spl_0;
  wire n1253_o2_p_spl_00;
  wire n1253_o2_p_spl_01;
  wire n1253_o2_p_spl_1;
  wire n1253_o2_n_spl_;
  wire n1253_o2_n_spl_0;
  wire n1253_o2_n_spl_00;
  wire n1253_o2_n_spl_01;
  wire n1253_o2_n_spl_1;
  wire g273_p_spl_;
  wire g273_p_spl_0;
  wire g273_p_spl_1;
  wire g273_n_spl_;
  wire g273_n_spl_0;
  wire g273_n_spl_1;
  wire g293_p_spl_;
  wire g293_p_spl_0;
  wire g293_p_spl_1;
  wire g293_n_spl_;
  wire g293_n_spl_0;
  wire g293_n_spl_1;
  wire G391_o2_p_spl_;
  wire G391_o2_p_spl_0;
  wire G391_o2_p_spl_1;
  wire G391_o2_n_spl_;
  wire G391_o2_n_spl_0;
  wire G391_o2_n_spl_1;
  wire g313_p_spl_;
  wire g313_p_spl_0;
  wire g313_p_spl_1;
  wire g313_n_spl_;
  wire g313_n_spl_0;
  wire g313_n_spl_1;
  wire g333_p_spl_;
  wire g333_p_spl_0;
  wire g333_p_spl_1;
  wire g333_n_spl_;
  wire g333_n_spl_0;
  wire g333_n_spl_1;
  wire g353_p_spl_;
  wire g353_p_spl_0;
  wire g353_p_spl_1;
  wire g353_n_spl_;
  wire g353_n_spl_0;
  wire g353_n_spl_1;
  wire g373_p_spl_;
  wire g373_p_spl_0;
  wire g373_p_spl_1;
  wire g373_n_spl_;
  wire g373_n_spl_0;
  wire g373_n_spl_1;
  wire G247_o2_p_spl_;
  wire G234_o2_p_spl_;
  wire g390_n_spl_;
  wire G260_o2_p_spl_;
  wire G260_o2_p_spl_0;
  wire G273_o2_n_spl_;
  wire G273_o2_n_spl_0;
  wire G273_o2_n_spl_1;
  wire G260_o2_n_spl_;
  wire G260_o2_n_spl_0;
  wire G260_o2_n_spl_1;
  wire G273_o2_p_spl_;
  wire G273_o2_p_spl_0;
  wire G247_o2_n_spl_;
  wire G247_o2_n_spl_0;
  wire G247_o2_n_spl_1;
  wire G234_o2_n_spl_;
  wire G234_o2_n_spl_0;
  wire G234_o2_n_spl_1;
  wire G299_o2_p_spl_;
  wire G286_o2_p_spl_;
  wire g404_n_spl_;
  wire G312_o2_p_spl_;
  wire G312_o2_p_spl_0;
  wire G325_o2_n_spl_;
  wire G325_o2_n_spl_0;
  wire G325_o2_n_spl_1;
  wire G312_o2_n_spl_;
  wire G312_o2_n_spl_0;
  wire G312_o2_n_spl_1;
  wire G325_o2_p_spl_;
  wire G325_o2_p_spl_0;
  wire G299_o2_n_spl_;
  wire G299_o2_n_spl_0;
  wire G299_o2_n_spl_1;
  wire G286_o2_n_spl_;
  wire G286_o2_n_spl_0;
  wire G286_o2_n_spl_1;
  wire n331_lo_buf_o2_p_spl_;
  wire n283_lo_buf_o2_n_spl_;
  wire n283_lo_buf_o2_n_spl_0;
  wire n331_lo_buf_o2_n_spl_;
  wire n331_lo_buf_o2_n_spl_0;
  wire n283_lo_buf_o2_p_spl_;
  wire n427_lo_buf_o2_p_spl_;
  wire n379_lo_buf_o2_n_spl_;
  wire n379_lo_buf_o2_n_spl_0;
  wire n427_lo_buf_o2_n_spl_;
  wire n427_lo_buf_o2_n_spl_0;
  wire n379_lo_buf_o2_p_spl_;
  wire g423_n_spl_;
  wire g420_p_spl_;
  wire g423_p_spl_;
  wire g420_n_spl_;
  wire n763_lo_buf_o2_p_spl_;
  wire n763_lo_buf_o2_p_spl_0;
  wire n763_lo_buf_o2_p_spl_00;
  wire n763_lo_buf_o2_p_spl_01;
  wire n763_lo_buf_o2_p_spl_1;
  wire n763_lo_buf_o2_p_spl_10;
  wire n763_lo_buf_o2_p_spl_11;
  wire n763_lo_buf_o2_n_spl_;
  wire n763_lo_buf_o2_n_spl_0;
  wire n763_lo_buf_o2_n_spl_00;
  wire n763_lo_buf_o2_n_spl_01;
  wire n763_lo_buf_o2_n_spl_1;
  wire n763_lo_buf_o2_n_spl_10;
  wire n763_lo_buf_o2_n_spl_11;
  wire G201_o2_p_spl_;
  wire G201_o2_p_spl_0;
  wire G201_o2_p_spl_1;
  wire G198_o2_n_spl_;
  wire G198_o2_n_spl_0;
  wire G198_o2_n_spl_1;
  wire G201_o2_n_spl_;
  wire G201_o2_n_spl_0;
  wire G201_o2_n_spl_1;
  wire G198_o2_p_spl_;
  wire G198_o2_p_spl_0;
  wire G198_o2_p_spl_1;
  wire g430_n_spl_;
  wire g427_n_spl_;
  wire g430_p_spl_;
  wire g427_p_spl_;
  wire n343_lo_buf_o2_p_spl_;
  wire n295_lo_buf_o2_n_spl_;
  wire n295_lo_buf_o2_n_spl_0;
  wire n343_lo_buf_o2_n_spl_;
  wire n343_lo_buf_o2_n_spl_0;
  wire n295_lo_buf_o2_p_spl_;
  wire n439_lo_buf_o2_p_spl_;
  wire n391_lo_buf_o2_n_spl_;
  wire n391_lo_buf_o2_n_spl_0;
  wire n439_lo_buf_o2_n_spl_;
  wire n439_lo_buf_o2_n_spl_0;
  wire n391_lo_buf_o2_p_spl_;
  wire g442_n_spl_;
  wire g439_p_spl_;
  wire g442_p_spl_;
  wire g439_n_spl_;
  wire G207_o2_p_spl_;
  wire G207_o2_p_spl_0;
  wire G207_o2_p_spl_1;
  wire G204_o2_n_spl_;
  wire G204_o2_n_spl_0;
  wire G204_o2_n_spl_1;
  wire G207_o2_n_spl_;
  wire G207_o2_n_spl_0;
  wire G207_o2_n_spl_1;
  wire G204_o2_p_spl_;
  wire G204_o2_p_spl_0;
  wire G204_o2_p_spl_1;
  wire g449_n_spl_;
  wire g446_n_spl_;
  wire g449_p_spl_;
  wire g446_p_spl_;
  wire n355_lo_buf_o2_p_spl_;
  wire n307_lo_buf_o2_n_spl_;
  wire n307_lo_buf_o2_n_spl_0;
  wire n355_lo_buf_o2_n_spl_;
  wire n355_lo_buf_o2_n_spl_0;
  wire n307_lo_buf_o2_p_spl_;
  wire n451_lo_buf_o2_p_spl_;
  wire n403_lo_buf_o2_n_spl_;
  wire n403_lo_buf_o2_n_spl_0;
  wire n451_lo_buf_o2_n_spl_;
  wire n451_lo_buf_o2_n_spl_0;
  wire n403_lo_buf_o2_p_spl_;
  wire g461_n_spl_;
  wire g458_p_spl_;
  wire g461_p_spl_;
  wire g458_n_spl_;
  wire g468_n_spl_;
  wire g465_n_spl_;
  wire g468_p_spl_;
  wire g465_p_spl_;
  wire n367_lo_buf_o2_p_spl_;
  wire n319_lo_buf_o2_n_spl_;
  wire n319_lo_buf_o2_n_spl_0;
  wire n367_lo_buf_o2_n_spl_;
  wire n367_lo_buf_o2_n_spl_0;
  wire n319_lo_buf_o2_p_spl_;
  wire n463_lo_buf_o2_p_spl_;
  wire n415_lo_buf_o2_n_spl_;
  wire n415_lo_buf_o2_n_spl_0;
  wire n463_lo_buf_o2_n_spl_;
  wire n463_lo_buf_o2_n_spl_0;
  wire n415_lo_buf_o2_p_spl_;
  wire g480_n_spl_;
  wire g477_p_spl_;
  wire g480_p_spl_;
  wire g477_n_spl_;
  wire g487_n_spl_;
  wire g484_n_spl_;
  wire g487_p_spl_;
  wire g484_p_spl_;
  wire n523_lo_buf_o2_p_spl_;
  wire n475_lo_buf_o2_n_spl_;
  wire n475_lo_buf_o2_n_spl_0;
  wire n523_lo_buf_o2_n_spl_;
  wire n523_lo_buf_o2_n_spl_0;
  wire n475_lo_buf_o2_p_spl_;
  wire n619_lo_buf_o2_p_spl_;
  wire n571_lo_buf_o2_n_spl_;
  wire n571_lo_buf_o2_n_spl_0;
  wire n619_lo_buf_o2_n_spl_;
  wire n619_lo_buf_o2_n_spl_0;
  wire n571_lo_buf_o2_p_spl_;
  wire g499_n_spl_;
  wire g496_p_spl_;
  wire g499_p_spl_;
  wire g496_n_spl_;
  wire G189_o2_p_spl_;
  wire G189_o2_p_spl_0;
  wire G189_o2_p_spl_1;
  wire G186_o2_n_spl_;
  wire G186_o2_n_spl_0;
  wire G186_o2_n_spl_1;
  wire G189_o2_n_spl_;
  wire G189_o2_n_spl_0;
  wire G189_o2_n_spl_1;
  wire G186_o2_p_spl_;
  wire G186_o2_p_spl_0;
  wire G186_o2_p_spl_1;
  wire g506_n_spl_;
  wire g503_n_spl_;
  wire g506_p_spl_;
  wire g503_p_spl_;
  wire n535_lo_buf_o2_p_spl_;
  wire n487_lo_buf_o2_n_spl_;
  wire n487_lo_buf_o2_n_spl_0;
  wire n535_lo_buf_o2_n_spl_;
  wire n535_lo_buf_o2_n_spl_0;
  wire n487_lo_buf_o2_p_spl_;
  wire n631_lo_buf_o2_p_spl_;
  wire n583_lo_buf_o2_n_spl_;
  wire n583_lo_buf_o2_n_spl_0;
  wire n631_lo_buf_o2_n_spl_;
  wire n631_lo_buf_o2_n_spl_0;
  wire n583_lo_buf_o2_p_spl_;
  wire g518_n_spl_;
  wire g515_p_spl_;
  wire g518_p_spl_;
  wire g515_n_spl_;
  wire G195_o2_p_spl_;
  wire G195_o2_p_spl_0;
  wire G195_o2_p_spl_1;
  wire G192_o2_n_spl_;
  wire G192_o2_n_spl_0;
  wire G192_o2_n_spl_1;
  wire G195_o2_n_spl_;
  wire G195_o2_n_spl_0;
  wire G195_o2_n_spl_1;
  wire G192_o2_p_spl_;
  wire G192_o2_p_spl_0;
  wire G192_o2_p_spl_1;
  wire g525_n_spl_;
  wire g522_n_spl_;
  wire g525_p_spl_;
  wire g522_p_spl_;
  wire n547_lo_buf_o2_p_spl_;
  wire n499_lo_buf_o2_n_spl_;
  wire n499_lo_buf_o2_n_spl_0;
  wire n547_lo_buf_o2_n_spl_;
  wire n547_lo_buf_o2_n_spl_0;
  wire n499_lo_buf_o2_p_spl_;
  wire n643_lo_buf_o2_p_spl_;
  wire n595_lo_buf_o2_n_spl_;
  wire n595_lo_buf_o2_n_spl_0;
  wire n643_lo_buf_o2_n_spl_;
  wire n643_lo_buf_o2_n_spl_0;
  wire n595_lo_buf_o2_p_spl_;
  wire g537_n_spl_;
  wire g534_p_spl_;
  wire g537_p_spl_;
  wire g534_n_spl_;
  wire g544_n_spl_;
  wire g541_n_spl_;
  wire g544_p_spl_;
  wire g541_p_spl_;
  wire n559_lo_buf_o2_p_spl_;
  wire n511_lo_buf_o2_n_spl_;
  wire n511_lo_buf_o2_n_spl_0;
  wire n559_lo_buf_o2_n_spl_;
  wire n559_lo_buf_o2_n_spl_0;
  wire n511_lo_buf_o2_p_spl_;
  wire n655_lo_buf_o2_p_spl_;
  wire n607_lo_buf_o2_n_spl_;
  wire n607_lo_buf_o2_n_spl_0;
  wire n655_lo_buf_o2_n_spl_;
  wire n655_lo_buf_o2_n_spl_0;
  wire n607_lo_buf_o2_p_spl_;
  wire g556_n_spl_;
  wire g553_p_spl_;
  wire g556_p_spl_;
  wire g553_n_spl_;
  wire g563_n_spl_;
  wire g560_n_spl_;
  wire g563_p_spl_;
  wire g560_p_spl_;
  wire n292_lo_buf_o2_p_spl_;
  wire n280_lo_buf_o2_n_spl_;
  wire n280_lo_buf_o2_n_spl_0;
  wire n292_lo_buf_o2_n_spl_;
  wire n292_lo_buf_o2_n_spl_0;
  wire n280_lo_buf_o2_p_spl_;
  wire n316_lo_buf_o2_p_spl_;
  wire n304_lo_buf_o2_n_spl_;
  wire n304_lo_buf_o2_n_spl_0;
  wire n316_lo_buf_o2_n_spl_;
  wire n316_lo_buf_o2_n_spl_0;
  wire n304_lo_buf_o2_p_spl_;
  wire n340_lo_buf_o2_p_spl_;
  wire n328_lo_buf_o2_n_spl_;
  wire n328_lo_buf_o2_n_spl_0;
  wire n340_lo_buf_o2_n_spl_;
  wire n340_lo_buf_o2_n_spl_0;
  wire n328_lo_buf_o2_p_spl_;
  wire n364_lo_buf_o2_p_spl_;
  wire n352_lo_buf_o2_n_spl_;
  wire n352_lo_buf_o2_n_spl_0;
  wire n364_lo_buf_o2_n_spl_;
  wire n364_lo_buf_o2_n_spl_0;
  wire n352_lo_buf_o2_p_spl_;
  wire n388_lo_buf_o2_p_spl_;
  wire n376_lo_buf_o2_n_spl_;
  wire n376_lo_buf_o2_n_spl_0;
  wire n388_lo_buf_o2_n_spl_;
  wire n388_lo_buf_o2_n_spl_0;
  wire n376_lo_buf_o2_p_spl_;
  wire n412_lo_buf_o2_p_spl_;
  wire n400_lo_buf_o2_n_spl_;
  wire n400_lo_buf_o2_n_spl_0;
  wire n412_lo_buf_o2_n_spl_;
  wire n412_lo_buf_o2_n_spl_0;
  wire n400_lo_buf_o2_p_spl_;
  wire n436_lo_buf_o2_p_spl_;
  wire n424_lo_buf_o2_n_spl_;
  wire n424_lo_buf_o2_n_spl_0;
  wire n436_lo_buf_o2_n_spl_;
  wire n436_lo_buf_o2_n_spl_0;
  wire n424_lo_buf_o2_p_spl_;
  wire n460_lo_buf_o2_p_spl_;
  wire n448_lo_buf_o2_n_spl_;
  wire n448_lo_buf_o2_n_spl_0;
  wire n460_lo_buf_o2_n_spl_;
  wire n460_lo_buf_o2_n_spl_0;
  wire n448_lo_buf_o2_p_spl_;
  wire n484_lo_buf_o2_p_spl_;
  wire n472_lo_buf_o2_n_spl_;
  wire n472_lo_buf_o2_n_spl_0;
  wire n484_lo_buf_o2_n_spl_;
  wire n484_lo_buf_o2_n_spl_0;
  wire n472_lo_buf_o2_p_spl_;
  wire n508_lo_buf_o2_p_spl_;
  wire n496_lo_buf_o2_n_spl_;
  wire n496_lo_buf_o2_n_spl_0;
  wire n508_lo_buf_o2_n_spl_;
  wire n508_lo_buf_o2_n_spl_0;
  wire n496_lo_buf_o2_p_spl_;
  wire n532_lo_buf_o2_p_spl_;
  wire n520_lo_buf_o2_n_spl_;
  wire n520_lo_buf_o2_n_spl_0;
  wire n532_lo_buf_o2_n_spl_;
  wire n532_lo_buf_o2_n_spl_0;
  wire n520_lo_buf_o2_p_spl_;
  wire n556_lo_buf_o2_p_spl_;
  wire n544_lo_buf_o2_n_spl_;
  wire n544_lo_buf_o2_n_spl_0;
  wire n556_lo_buf_o2_n_spl_;
  wire n556_lo_buf_o2_n_spl_0;
  wire n544_lo_buf_o2_p_spl_;
  wire n580_lo_buf_o2_p_spl_;
  wire n568_lo_buf_o2_n_spl_;
  wire n568_lo_buf_o2_n_spl_0;
  wire n580_lo_buf_o2_n_spl_;
  wire n580_lo_buf_o2_n_spl_0;
  wire n568_lo_buf_o2_p_spl_;
  wire n604_lo_buf_o2_p_spl_;
  wire n592_lo_buf_o2_n_spl_;
  wire n592_lo_buf_o2_n_spl_0;
  wire n604_lo_buf_o2_n_spl_;
  wire n604_lo_buf_o2_n_spl_0;
  wire n592_lo_buf_o2_p_spl_;
  wire n628_lo_buf_o2_p_spl_;
  wire n616_lo_buf_o2_n_spl_;
  wire n616_lo_buf_o2_n_spl_0;
  wire n628_lo_buf_o2_n_spl_;
  wire n628_lo_buf_o2_n_spl_0;
  wire n616_lo_buf_o2_p_spl_;
  wire n652_lo_buf_o2_p_spl_;
  wire n640_lo_buf_o2_n_spl_;
  wire n640_lo_buf_o2_n_spl_0;
  wire n652_lo_buf_o2_n_spl_;
  wire n652_lo_buf_o2_n_spl_0;
  wire n640_lo_buf_o2_p_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  buf

  (
    G33_p,
    G33
  );


  not

  (
    G33_n,
    G33
  );


  buf

  (
    G34_p,
    G34
  );


  not

  (
    G34_n,
    G34
  );


  buf

  (
    G35_p,
    G35
  );


  not

  (
    G35_n,
    G35
  );


  buf

  (
    G36_p,
    G36
  );


  not

  (
    G36_n,
    G36
  );


  buf

  (
    G37_p,
    G37
  );


  not

  (
    G37_n,
    G37
  );


  buf

  (
    G38_p,
    G38
  );


  not

  (
    G38_n,
    G38
  );


  buf

  (
    G39_p,
    G39
  );


  not

  (
    G39_n,
    G39
  );


  buf

  (
    G40_p,
    G40
  );


  not

  (
    G40_n,
    G40
  );


  buf

  (
    G41_p,
    G41
  );


  not

  (
    G41_n,
    G41
  );


  buf

  (
    n286_lo_p,
    n286_lo
  );


  not

  (
    n286_lo_n,
    n286_lo
  );


  buf

  (
    n298_lo_p,
    n298_lo
  );


  not

  (
    n298_lo_n,
    n298_lo
  );


  buf

  (
    n310_lo_p,
    n310_lo
  );


  not

  (
    n310_lo_n,
    n310_lo
  );


  buf

  (
    n322_lo_p,
    n322_lo
  );


  not

  (
    n322_lo_n,
    n322_lo
  );


  buf

  (
    n334_lo_p,
    n334_lo
  );


  not

  (
    n334_lo_n,
    n334_lo
  );


  buf

  (
    n346_lo_p,
    n346_lo
  );


  not

  (
    n346_lo_n,
    n346_lo
  );


  buf

  (
    n358_lo_p,
    n358_lo
  );


  not

  (
    n358_lo_n,
    n358_lo
  );


  buf

  (
    n370_lo_p,
    n370_lo
  );


  not

  (
    n370_lo_n,
    n370_lo
  );


  buf

  (
    n382_lo_p,
    n382_lo
  );


  not

  (
    n382_lo_n,
    n382_lo
  );


  buf

  (
    n394_lo_p,
    n394_lo
  );


  not

  (
    n394_lo_n,
    n394_lo
  );


  buf

  (
    n406_lo_p,
    n406_lo
  );


  not

  (
    n406_lo_n,
    n406_lo
  );


  buf

  (
    n418_lo_p,
    n418_lo
  );


  not

  (
    n418_lo_n,
    n418_lo
  );


  buf

  (
    n430_lo_p,
    n430_lo
  );


  not

  (
    n430_lo_n,
    n430_lo
  );


  buf

  (
    n442_lo_p,
    n442_lo
  );


  not

  (
    n442_lo_n,
    n442_lo
  );


  buf

  (
    n454_lo_p,
    n454_lo
  );


  not

  (
    n454_lo_n,
    n454_lo
  );


  buf

  (
    n466_lo_p,
    n466_lo
  );


  not

  (
    n466_lo_n,
    n466_lo
  );


  buf

  (
    n478_lo_p,
    n478_lo
  );


  not

  (
    n478_lo_n,
    n478_lo
  );


  buf

  (
    n490_lo_p,
    n490_lo
  );


  not

  (
    n490_lo_n,
    n490_lo
  );


  buf

  (
    n502_lo_p,
    n502_lo
  );


  not

  (
    n502_lo_n,
    n502_lo
  );


  buf

  (
    n514_lo_p,
    n514_lo
  );


  not

  (
    n514_lo_n,
    n514_lo
  );


  buf

  (
    n526_lo_p,
    n526_lo
  );


  not

  (
    n526_lo_n,
    n526_lo
  );


  buf

  (
    n538_lo_p,
    n538_lo
  );


  not

  (
    n538_lo_n,
    n538_lo
  );


  buf

  (
    n550_lo_p,
    n550_lo
  );


  not

  (
    n550_lo_n,
    n550_lo
  );


  buf

  (
    n562_lo_p,
    n562_lo
  );


  not

  (
    n562_lo_n,
    n562_lo
  );


  buf

  (
    n574_lo_p,
    n574_lo
  );


  not

  (
    n574_lo_n,
    n574_lo
  );


  buf

  (
    n586_lo_p,
    n586_lo
  );


  not

  (
    n586_lo_n,
    n586_lo
  );


  buf

  (
    n598_lo_p,
    n598_lo
  );


  not

  (
    n598_lo_n,
    n598_lo
  );


  buf

  (
    n610_lo_p,
    n610_lo
  );


  not

  (
    n610_lo_n,
    n610_lo
  );


  buf

  (
    n622_lo_p,
    n622_lo
  );


  not

  (
    n622_lo_n,
    n622_lo
  );


  buf

  (
    n634_lo_p,
    n634_lo
  );


  not

  (
    n634_lo_n,
    n634_lo
  );


  buf

  (
    n646_lo_p,
    n646_lo
  );


  not

  (
    n646_lo_n,
    n646_lo
  );


  buf

  (
    n658_lo_p,
    n658_lo
  );


  not

  (
    n658_lo_n,
    n658_lo
  );


  buf

  (
    n661_lo_p,
    n661_lo
  );


  not

  (
    n661_lo_n,
    n661_lo
  );


  buf

  (
    n673_lo_p,
    n673_lo
  );


  not

  (
    n673_lo_n,
    n673_lo
  );


  buf

  (
    n685_lo_p,
    n685_lo
  );


  not

  (
    n685_lo_n,
    n685_lo
  );


  buf

  (
    n697_lo_p,
    n697_lo
  );


  not

  (
    n697_lo_n,
    n697_lo
  );


  buf

  (
    n709_lo_p,
    n709_lo
  );


  not

  (
    n709_lo_n,
    n709_lo
  );


  buf

  (
    n721_lo_p,
    n721_lo
  );


  not

  (
    n721_lo_n,
    n721_lo
  );


  buf

  (
    n733_lo_p,
    n733_lo
  );


  not

  (
    n733_lo_n,
    n733_lo
  );


  buf

  (
    n745_lo_p,
    n745_lo
  );


  not

  (
    n745_lo_n,
    n745_lo
  );


  buf

  (
    n757_lo_p,
    n757_lo
  );


  not

  (
    n757_lo_n,
    n757_lo
  );


  buf

  (
    n1248_o2_p,
    n1248_o2
  );


  not

  (
    n1248_o2_n,
    n1248_o2
  );


  buf

  (
    n1249_o2_p,
    n1249_o2
  );


  not

  (
    n1249_o2_n,
    n1249_o2
  );


  buf

  (
    n1250_o2_p,
    n1250_o2
  );


  not

  (
    n1250_o2_n,
    n1250_o2
  );


  buf

  (
    n1251_o2_p,
    n1251_o2
  );


  not

  (
    n1251_o2_n,
    n1251_o2
  );


  buf

  (
    n1252_o2_p,
    n1252_o2
  );


  not

  (
    n1252_o2_n,
    n1252_o2
  );


  buf

  (
    n1253_o2_p,
    n1253_o2
  );


  not

  (
    n1253_o2_n,
    n1253_o2
  );


  buf

  (
    n1254_o2_p,
    n1254_o2
  );


  not

  (
    n1254_o2_n,
    n1254_o2
  );


  buf

  (
    n1255_o2_p,
    n1255_o2
  );


  not

  (
    n1255_o2_n,
    n1255_o2
  );


  buf

  (
    n1207_o2_p,
    n1207_o2
  );


  not

  (
    n1207_o2_n,
    n1207_o2
  );


  buf

  (
    n1208_o2_p,
    n1208_o2
  );


  not

  (
    n1208_o2_n,
    n1208_o2
  );


  buf

  (
    n1209_o2_p,
    n1209_o2
  );


  not

  (
    n1209_o2_n,
    n1209_o2
  );


  buf

  (
    n1210_o2_p,
    n1210_o2
  );


  not

  (
    n1210_o2_n,
    n1210_o2
  );


  buf

  (
    n1211_o2_p,
    n1211_o2
  );


  not

  (
    n1211_o2_n,
    n1211_o2
  );


  buf

  (
    n1212_o2_p,
    n1212_o2
  );


  not

  (
    n1212_o2_n,
    n1212_o2
  );


  buf

  (
    n1213_o2_p,
    n1213_o2
  );


  not

  (
    n1213_o2_n,
    n1213_o2
  );


  buf

  (
    n1214_o2_p,
    n1214_o2
  );


  not

  (
    n1214_o2_n,
    n1214_o2
  );


  buf

  (
    n1215_o2_p,
    n1215_o2
  );


  not

  (
    n1215_o2_n,
    n1215_o2
  );


  buf

  (
    n1216_o2_p,
    n1216_o2
  );


  not

  (
    n1216_o2_n,
    n1216_o2
  );


  buf

  (
    n1217_o2_p,
    n1217_o2
  );


  not

  (
    n1217_o2_n,
    n1217_o2
  );


  buf

  (
    n1218_o2_p,
    n1218_o2
  );


  not

  (
    n1218_o2_n,
    n1218_o2
  );


  buf

  (
    n1219_o2_p,
    n1219_o2
  );


  not

  (
    n1219_o2_n,
    n1219_o2
  );


  buf

  (
    n1220_o2_p,
    n1220_o2
  );


  not

  (
    n1220_o2_n,
    n1220_o2
  );


  buf

  (
    n1221_o2_p,
    n1221_o2
  );


  not

  (
    n1221_o2_n,
    n1221_o2
  );


  buf

  (
    n1222_o2_p,
    n1222_o2
  );


  not

  (
    n1222_o2_n,
    n1222_o2
  );


  buf

  (
    n1223_o2_p,
    n1223_o2
  );


  not

  (
    n1223_o2_n,
    n1223_o2
  );


  buf

  (
    n1224_o2_p,
    n1224_o2
  );


  not

  (
    n1224_o2_n,
    n1224_o2
  );


  buf

  (
    n1225_o2_p,
    n1225_o2
  );


  not

  (
    n1225_o2_n,
    n1225_o2
  );


  buf

  (
    n1226_o2_p,
    n1226_o2
  );


  not

  (
    n1226_o2_n,
    n1226_o2
  );


  buf

  (
    n1227_o2_p,
    n1227_o2
  );


  not

  (
    n1227_o2_n,
    n1227_o2
  );


  buf

  (
    n1228_o2_p,
    n1228_o2
  );


  not

  (
    n1228_o2_n,
    n1228_o2
  );


  buf

  (
    n1229_o2_p,
    n1229_o2
  );


  not

  (
    n1229_o2_n,
    n1229_o2
  );


  buf

  (
    n1230_o2_p,
    n1230_o2
  );


  not

  (
    n1230_o2_n,
    n1230_o2
  );


  buf

  (
    n1231_o2_p,
    n1231_o2
  );


  not

  (
    n1231_o2_n,
    n1231_o2
  );


  buf

  (
    n1232_o2_p,
    n1232_o2
  );


  not

  (
    n1232_o2_n,
    n1232_o2
  );


  buf

  (
    n1233_o2_p,
    n1233_o2
  );


  not

  (
    n1233_o2_n,
    n1233_o2
  );


  buf

  (
    n1234_o2_p,
    n1234_o2
  );


  not

  (
    n1234_o2_n,
    n1234_o2
  );


  buf

  (
    n1235_o2_p,
    n1235_o2
  );


  not

  (
    n1235_o2_n,
    n1235_o2
  );


  buf

  (
    n1236_o2_p,
    n1236_o2
  );


  not

  (
    n1236_o2_n,
    n1236_o2
  );


  buf

  (
    n1237_o2_p,
    n1237_o2
  );


  not

  (
    n1237_o2_n,
    n1237_o2
  );


  buf

  (
    n1238_o2_p,
    n1238_o2
  );


  not

  (
    n1238_o2_n,
    n1238_o2
  );


  buf

  (
    G374_o2_p,
    G374_o2
  );


  not

  (
    G374_o2_n,
    G374_o2
  );


  buf

  (
    G376_o2_p,
    G376_o2
  );


  not

  (
    G376_o2_n,
    G376_o2
  );


  buf

  (
    G370_o2_p,
    G370_o2
  );


  not

  (
    G370_o2_n,
    G370_o2
  );


  buf

  (
    G372_o2_p,
    G372_o2
  );


  not

  (
    G372_o2_n,
    G372_o2
  );


  buf

  (
    G373_o2_p,
    G373_o2
  );


  not

  (
    G373_o2_n,
    G373_o2
  );


  buf

  (
    G377_o2_p,
    G377_o2
  );


  not

  (
    G377_o2_n,
    G377_o2
  );


  buf

  (
    G371_o2_p,
    G371_o2
  );


  not

  (
    G371_o2_n,
    G371_o2
  );


  buf

  (
    G375_o2_p,
    G375_o2
  );


  not

  (
    G375_o2_n,
    G375_o2
  );


  buf

  (
    G354_o2_p,
    G354_o2
  );


  not

  (
    G354_o2_n,
    G354_o2
  );


  buf

  (
    G356_o2_p,
    G356_o2
  );


  not

  (
    G356_o2_n,
    G356_o2
  );


  buf

  (
    G350_o2_p,
    G350_o2
  );


  not

  (
    G350_o2_n,
    G350_o2
  );


  buf

  (
    G352_o2_p,
    G352_o2
  );


  not

  (
    G352_o2_n,
    G352_o2
  );


  buf

  (
    G353_o2_p,
    G353_o2
  );


  not

  (
    G353_o2_n,
    G353_o2
  );


  buf

  (
    G357_o2_p,
    G357_o2
  );


  not

  (
    G357_o2_n,
    G357_o2
  );


  buf

  (
    G351_o2_p,
    G351_o2
  );


  not

  (
    G351_o2_n,
    G351_o2
  );


  buf

  (
    G355_o2_p,
    G355_o2
  );


  not

  (
    G355_o2_n,
    G355_o2
  );


  buf

  (
    G386_o2_p,
    G386_o2
  );


  not

  (
    G386_o2_n,
    G386_o2
  );


  buf

  (
    G391_o2_p,
    G391_o2
  );


  not

  (
    G391_o2_n,
    G391_o2
  );


  buf

  (
    n283_lo_buf_o2_p,
    n283_lo_buf_o2
  );


  not

  (
    n283_lo_buf_o2_n,
    n283_lo_buf_o2
  );


  buf

  (
    n295_lo_buf_o2_p,
    n295_lo_buf_o2
  );


  not

  (
    n295_lo_buf_o2_n,
    n295_lo_buf_o2
  );


  buf

  (
    n307_lo_buf_o2_p,
    n307_lo_buf_o2
  );


  not

  (
    n307_lo_buf_o2_n,
    n307_lo_buf_o2
  );


  buf

  (
    n319_lo_buf_o2_p,
    n319_lo_buf_o2
  );


  not

  (
    n319_lo_buf_o2_n,
    n319_lo_buf_o2
  );


  buf

  (
    n331_lo_buf_o2_p,
    n331_lo_buf_o2
  );


  not

  (
    n331_lo_buf_o2_n,
    n331_lo_buf_o2
  );


  buf

  (
    n343_lo_buf_o2_p,
    n343_lo_buf_o2
  );


  not

  (
    n343_lo_buf_o2_n,
    n343_lo_buf_o2
  );


  buf

  (
    n355_lo_buf_o2_p,
    n355_lo_buf_o2
  );


  not

  (
    n355_lo_buf_o2_n,
    n355_lo_buf_o2
  );


  buf

  (
    n367_lo_buf_o2_p,
    n367_lo_buf_o2
  );


  not

  (
    n367_lo_buf_o2_n,
    n367_lo_buf_o2
  );


  buf

  (
    n379_lo_buf_o2_p,
    n379_lo_buf_o2
  );


  not

  (
    n379_lo_buf_o2_n,
    n379_lo_buf_o2
  );


  buf

  (
    n391_lo_buf_o2_p,
    n391_lo_buf_o2
  );


  not

  (
    n391_lo_buf_o2_n,
    n391_lo_buf_o2
  );


  buf

  (
    n403_lo_buf_o2_p,
    n403_lo_buf_o2
  );


  not

  (
    n403_lo_buf_o2_n,
    n403_lo_buf_o2
  );


  buf

  (
    n415_lo_buf_o2_p,
    n415_lo_buf_o2
  );


  not

  (
    n415_lo_buf_o2_n,
    n415_lo_buf_o2
  );


  buf

  (
    n427_lo_buf_o2_p,
    n427_lo_buf_o2
  );


  not

  (
    n427_lo_buf_o2_n,
    n427_lo_buf_o2
  );


  buf

  (
    n439_lo_buf_o2_p,
    n439_lo_buf_o2
  );


  not

  (
    n439_lo_buf_o2_n,
    n439_lo_buf_o2
  );


  buf

  (
    n451_lo_buf_o2_p,
    n451_lo_buf_o2
  );


  not

  (
    n451_lo_buf_o2_n,
    n451_lo_buf_o2
  );


  buf

  (
    n463_lo_buf_o2_p,
    n463_lo_buf_o2
  );


  not

  (
    n463_lo_buf_o2_n,
    n463_lo_buf_o2
  );


  buf

  (
    n475_lo_buf_o2_p,
    n475_lo_buf_o2
  );


  not

  (
    n475_lo_buf_o2_n,
    n475_lo_buf_o2
  );


  buf

  (
    n487_lo_buf_o2_p,
    n487_lo_buf_o2
  );


  not

  (
    n487_lo_buf_o2_n,
    n487_lo_buf_o2
  );


  buf

  (
    n499_lo_buf_o2_p,
    n499_lo_buf_o2
  );


  not

  (
    n499_lo_buf_o2_n,
    n499_lo_buf_o2
  );


  buf

  (
    n511_lo_buf_o2_p,
    n511_lo_buf_o2
  );


  not

  (
    n511_lo_buf_o2_n,
    n511_lo_buf_o2
  );


  buf

  (
    n523_lo_buf_o2_p,
    n523_lo_buf_o2
  );


  not

  (
    n523_lo_buf_o2_n,
    n523_lo_buf_o2
  );


  buf

  (
    n535_lo_buf_o2_p,
    n535_lo_buf_o2
  );


  not

  (
    n535_lo_buf_o2_n,
    n535_lo_buf_o2
  );


  buf

  (
    n547_lo_buf_o2_p,
    n547_lo_buf_o2
  );


  not

  (
    n547_lo_buf_o2_n,
    n547_lo_buf_o2
  );


  buf

  (
    n559_lo_buf_o2_p,
    n559_lo_buf_o2
  );


  not

  (
    n559_lo_buf_o2_n,
    n559_lo_buf_o2
  );


  buf

  (
    n571_lo_buf_o2_p,
    n571_lo_buf_o2
  );


  not

  (
    n571_lo_buf_o2_n,
    n571_lo_buf_o2
  );


  buf

  (
    n583_lo_buf_o2_p,
    n583_lo_buf_o2
  );


  not

  (
    n583_lo_buf_o2_n,
    n583_lo_buf_o2
  );


  buf

  (
    n595_lo_buf_o2_p,
    n595_lo_buf_o2
  );


  not

  (
    n595_lo_buf_o2_n,
    n595_lo_buf_o2
  );


  buf

  (
    n607_lo_buf_o2_p,
    n607_lo_buf_o2
  );


  not

  (
    n607_lo_buf_o2_n,
    n607_lo_buf_o2
  );


  buf

  (
    n619_lo_buf_o2_p,
    n619_lo_buf_o2
  );


  not

  (
    n619_lo_buf_o2_n,
    n619_lo_buf_o2
  );


  buf

  (
    n631_lo_buf_o2_p,
    n631_lo_buf_o2
  );


  not

  (
    n631_lo_buf_o2_n,
    n631_lo_buf_o2
  );


  buf

  (
    n643_lo_buf_o2_p,
    n643_lo_buf_o2
  );


  not

  (
    n643_lo_buf_o2_n,
    n643_lo_buf_o2
  );


  buf

  (
    n655_lo_buf_o2_p,
    n655_lo_buf_o2
  );


  not

  (
    n655_lo_buf_o2_n,
    n655_lo_buf_o2
  );


  buf

  (
    G234_o2_p,
    G234_o2
  );


  not

  (
    G234_o2_n,
    G234_o2
  );


  buf

  (
    G247_o2_p,
    G247_o2
  );


  not

  (
    G247_o2_n,
    G247_o2
  );


  buf

  (
    G260_o2_p,
    G260_o2
  );


  not

  (
    G260_o2_n,
    G260_o2
  );


  buf

  (
    G273_o2_p,
    G273_o2
  );


  not

  (
    G273_o2_n,
    G273_o2
  );


  buf

  (
    G286_o2_p,
    G286_o2
  );


  not

  (
    G286_o2_n,
    G286_o2
  );


  buf

  (
    G299_o2_p,
    G299_o2
  );


  not

  (
    G299_o2_n,
    G299_o2
  );


  buf

  (
    G312_o2_p,
    G312_o2
  );


  not

  (
    G312_o2_n,
    G312_o2
  );


  buf

  (
    G325_o2_p,
    G325_o2
  );


  not

  (
    G325_o2_n,
    G325_o2
  );


  buf

  (
    n667_lo_buf_o2_p,
    n667_lo_buf_o2
  );


  not

  (
    n667_lo_buf_o2_n,
    n667_lo_buf_o2
  );


  buf

  (
    n679_lo_buf_o2_p,
    n679_lo_buf_o2
  );


  not

  (
    n679_lo_buf_o2_n,
    n679_lo_buf_o2
  );


  buf

  (
    n691_lo_buf_o2_p,
    n691_lo_buf_o2
  );


  not

  (
    n691_lo_buf_o2_n,
    n691_lo_buf_o2
  );


  buf

  (
    n703_lo_buf_o2_p,
    n703_lo_buf_o2
  );


  not

  (
    n703_lo_buf_o2_n,
    n703_lo_buf_o2
  );


  buf

  (
    n715_lo_buf_o2_p,
    n715_lo_buf_o2
  );


  not

  (
    n715_lo_buf_o2_n,
    n715_lo_buf_o2
  );


  buf

  (
    n727_lo_buf_o2_p,
    n727_lo_buf_o2
  );


  not

  (
    n727_lo_buf_o2_n,
    n727_lo_buf_o2
  );


  buf

  (
    n739_lo_buf_o2_p,
    n739_lo_buf_o2
  );


  not

  (
    n739_lo_buf_o2_n,
    n739_lo_buf_o2
  );


  buf

  (
    n751_lo_buf_o2_p,
    n751_lo_buf_o2
  );


  not

  (
    n751_lo_buf_o2_n,
    n751_lo_buf_o2
  );


  buf

  (
    n763_lo_buf_o2_p,
    n763_lo_buf_o2
  );


  not

  (
    n763_lo_buf_o2_n,
    n763_lo_buf_o2
  );


  buf

  (
    G186_o2_p,
    G186_o2
  );


  not

  (
    G186_o2_n,
    G186_o2
  );


  buf

  (
    G189_o2_p,
    G189_o2
  );


  not

  (
    G189_o2_n,
    G189_o2
  );


  buf

  (
    G192_o2_p,
    G192_o2
  );


  not

  (
    G192_o2_n,
    G192_o2
  );


  buf

  (
    G195_o2_p,
    G195_o2
  );


  not

  (
    G195_o2_n,
    G195_o2
  );


  buf

  (
    G198_o2_p,
    G198_o2
  );


  not

  (
    G198_o2_n,
    G198_o2
  );


  buf

  (
    G201_o2_p,
    G201_o2
  );


  not

  (
    G201_o2_n,
    G201_o2
  );


  buf

  (
    G204_o2_p,
    G204_o2
  );


  not

  (
    G204_o2_n,
    G204_o2
  );


  buf

  (
    G207_o2_p,
    G207_o2
  );


  not

  (
    G207_o2_n,
    G207_o2
  );


  buf

  (
    n280_lo_buf_o2_p,
    n280_lo_buf_o2
  );


  not

  (
    n280_lo_buf_o2_n,
    n280_lo_buf_o2
  );


  buf

  (
    n292_lo_buf_o2_p,
    n292_lo_buf_o2
  );


  not

  (
    n292_lo_buf_o2_n,
    n292_lo_buf_o2
  );


  buf

  (
    n304_lo_buf_o2_p,
    n304_lo_buf_o2
  );


  not

  (
    n304_lo_buf_o2_n,
    n304_lo_buf_o2
  );


  buf

  (
    n316_lo_buf_o2_p,
    n316_lo_buf_o2
  );


  not

  (
    n316_lo_buf_o2_n,
    n316_lo_buf_o2
  );


  buf

  (
    n328_lo_buf_o2_p,
    n328_lo_buf_o2
  );


  not

  (
    n328_lo_buf_o2_n,
    n328_lo_buf_o2
  );


  buf

  (
    n340_lo_buf_o2_p,
    n340_lo_buf_o2
  );


  not

  (
    n340_lo_buf_o2_n,
    n340_lo_buf_o2
  );


  buf

  (
    n352_lo_buf_o2_p,
    n352_lo_buf_o2
  );


  not

  (
    n352_lo_buf_o2_n,
    n352_lo_buf_o2
  );


  buf

  (
    n364_lo_buf_o2_p,
    n364_lo_buf_o2
  );


  not

  (
    n364_lo_buf_o2_n,
    n364_lo_buf_o2
  );


  buf

  (
    n376_lo_buf_o2_p,
    n376_lo_buf_o2
  );


  not

  (
    n376_lo_buf_o2_n,
    n376_lo_buf_o2
  );


  buf

  (
    n388_lo_buf_o2_p,
    n388_lo_buf_o2
  );


  not

  (
    n388_lo_buf_o2_n,
    n388_lo_buf_o2
  );


  buf

  (
    n400_lo_buf_o2_p,
    n400_lo_buf_o2
  );


  not

  (
    n400_lo_buf_o2_n,
    n400_lo_buf_o2
  );


  buf

  (
    n412_lo_buf_o2_p,
    n412_lo_buf_o2
  );


  not

  (
    n412_lo_buf_o2_n,
    n412_lo_buf_o2
  );


  buf

  (
    n424_lo_buf_o2_p,
    n424_lo_buf_o2
  );


  not

  (
    n424_lo_buf_o2_n,
    n424_lo_buf_o2
  );


  buf

  (
    n436_lo_buf_o2_p,
    n436_lo_buf_o2
  );


  not

  (
    n436_lo_buf_o2_n,
    n436_lo_buf_o2
  );


  buf

  (
    n448_lo_buf_o2_p,
    n448_lo_buf_o2
  );


  not

  (
    n448_lo_buf_o2_n,
    n448_lo_buf_o2
  );


  buf

  (
    n460_lo_buf_o2_p,
    n460_lo_buf_o2
  );


  not

  (
    n460_lo_buf_o2_n,
    n460_lo_buf_o2
  );


  buf

  (
    n472_lo_buf_o2_p,
    n472_lo_buf_o2
  );


  not

  (
    n472_lo_buf_o2_n,
    n472_lo_buf_o2
  );


  buf

  (
    n484_lo_buf_o2_p,
    n484_lo_buf_o2
  );


  not

  (
    n484_lo_buf_o2_n,
    n484_lo_buf_o2
  );


  buf

  (
    n496_lo_buf_o2_p,
    n496_lo_buf_o2
  );


  not

  (
    n496_lo_buf_o2_n,
    n496_lo_buf_o2
  );


  buf

  (
    n508_lo_buf_o2_p,
    n508_lo_buf_o2
  );


  not

  (
    n508_lo_buf_o2_n,
    n508_lo_buf_o2
  );


  buf

  (
    n520_lo_buf_o2_p,
    n520_lo_buf_o2
  );


  not

  (
    n520_lo_buf_o2_n,
    n520_lo_buf_o2
  );


  buf

  (
    n532_lo_buf_o2_p,
    n532_lo_buf_o2
  );


  not

  (
    n532_lo_buf_o2_n,
    n532_lo_buf_o2
  );


  buf

  (
    n544_lo_buf_o2_p,
    n544_lo_buf_o2
  );


  not

  (
    n544_lo_buf_o2_n,
    n544_lo_buf_o2
  );


  buf

  (
    n556_lo_buf_o2_p,
    n556_lo_buf_o2
  );


  not

  (
    n556_lo_buf_o2_n,
    n556_lo_buf_o2
  );


  buf

  (
    n568_lo_buf_o2_p,
    n568_lo_buf_o2
  );


  not

  (
    n568_lo_buf_o2_n,
    n568_lo_buf_o2
  );


  buf

  (
    n580_lo_buf_o2_p,
    n580_lo_buf_o2
  );


  not

  (
    n580_lo_buf_o2_n,
    n580_lo_buf_o2
  );


  buf

  (
    n592_lo_buf_o2_p,
    n592_lo_buf_o2
  );


  not

  (
    n592_lo_buf_o2_n,
    n592_lo_buf_o2
  );


  buf

  (
    n604_lo_buf_o2_p,
    n604_lo_buf_o2
  );


  not

  (
    n604_lo_buf_o2_n,
    n604_lo_buf_o2
  );


  buf

  (
    n616_lo_buf_o2_p,
    n616_lo_buf_o2
  );


  not

  (
    n616_lo_buf_o2_n,
    n616_lo_buf_o2
  );


  buf

  (
    n628_lo_buf_o2_p,
    n628_lo_buf_o2
  );


  not

  (
    n628_lo_buf_o2_n,
    n628_lo_buf_o2
  );


  buf

  (
    n640_lo_buf_o2_p,
    n640_lo_buf_o2
  );


  not

  (
    n640_lo_buf_o2_n,
    n640_lo_buf_o2
  );


  buf

  (
    n652_lo_buf_o2_p,
    n652_lo_buf_o2
  );


  not

  (
    n652_lo_buf_o2_n,
    n652_lo_buf_o2
  );


  and

  (
    g230_p,
    G350_o2_n,
    n1252_o2_p_spl_00
  );


  or

  (
    g230_n,
    G350_o2_p,
    n1252_o2_n_spl_00
  );


  and

  (
    g231_p,
    g230_p,
    n1254_o2_p_spl_00
  );


  or

  (
    g231_n,
    g230_n,
    n1254_o2_n_spl_00
  );


  and

  (
    g232_p,
    g231_p,
    G351_o2_n
  );


  or

  (
    g232_n,
    g231_n,
    G351_o2_p
  );


  and

  (
    g233_p,
    g232_p,
    G386_o2_p_spl_0
  );


  or

  (
    g233_n,
    g232_n,
    G386_o2_n_spl_0
  );


  and

  (
    g234_p,
    g233_p_spl_0,
    n1248_o2_p_spl_00
  );


  or

  (
    g234_n,
    g233_n_spl_0,
    n1248_o2_n_spl_00
  );


  or

  (
    g235_n,
    g234_n,
    n286_lo_p
  );


  or

  (
    g236_n,
    g234_p,
    n286_lo_n
  );


  and

  (
    g237_p,
    g236_n,
    g235_n
  );


  and

  (
    g238_p,
    g233_p_spl_0,
    n1249_o2_p_spl_00
  );


  or

  (
    g238_n,
    g233_n_spl_0,
    n1249_o2_n_spl_00
  );


  or

  (
    g239_n,
    g238_n,
    n298_lo_p
  );


  or

  (
    g240_n,
    g238_p,
    n298_lo_n
  );


  and

  (
    g241_p,
    g240_n,
    g239_n
  );


  and

  (
    g242_p,
    g233_p_spl_1,
    n1250_o2_p_spl_00
  );


  or

  (
    g242_n,
    g233_n_spl_1,
    n1250_o2_n_spl_00
  );


  or

  (
    g243_n,
    g242_n,
    n310_lo_p
  );


  or

  (
    g244_n,
    g242_p,
    n310_lo_n
  );


  and

  (
    g245_p,
    g244_n,
    g243_n
  );


  and

  (
    g246_p,
    g233_p_spl_1,
    n1251_o2_p_spl_00
  );


  or

  (
    g246_n,
    g233_n_spl_1,
    n1251_o2_n_spl_00
  );


  or

  (
    g247_n,
    g246_n,
    n322_lo_p
  );


  or

  (
    g248_n,
    g246_p,
    n322_lo_n
  );


  and

  (
    g249_p,
    g248_n,
    g247_n
  );


  and

  (
    g250_p,
    G352_o2_n,
    n1252_o2_p_spl_00
  );


  or

  (
    g250_n,
    G352_o2_p,
    n1252_o2_n_spl_00
  );


  and

  (
    g251_p,
    g250_p,
    G353_o2_n
  );


  or

  (
    g251_n,
    g250_n,
    G353_o2_p
  );


  and

  (
    g252_p,
    g251_p,
    n1255_o2_p_spl_00
  );


  or

  (
    g252_n,
    g251_n,
    n1255_o2_n_spl_00
  );


  and

  (
    g253_p,
    g252_p,
    G386_o2_p_spl_0
  );


  or

  (
    g253_n,
    g252_n,
    G386_o2_n_spl_0
  );


  and

  (
    g254_p,
    g253_p_spl_0,
    n1248_o2_p_spl_00
  );


  or

  (
    g254_n,
    g253_n_spl_0,
    n1248_o2_n_spl_00
  );


  or

  (
    g255_n,
    g254_n,
    n334_lo_p
  );


  or

  (
    g256_n,
    g254_p,
    n334_lo_n
  );


  and

  (
    g257_p,
    g256_n,
    g255_n
  );


  and

  (
    g258_p,
    g253_p_spl_0,
    n1249_o2_p_spl_00
  );


  or

  (
    g258_n,
    g253_n_spl_0,
    n1249_o2_n_spl_00
  );


  or

  (
    g259_n,
    g258_n,
    n346_lo_p
  );


  or

  (
    g260_n,
    g258_p,
    n346_lo_n
  );


  and

  (
    g261_p,
    g260_n,
    g259_n
  );


  and

  (
    g262_p,
    g253_p_spl_1,
    n1250_o2_p_spl_00
  );


  or

  (
    g262_n,
    g253_n_spl_1,
    n1250_o2_n_spl_00
  );


  or

  (
    g263_n,
    g262_n,
    n358_lo_p
  );


  or

  (
    g264_n,
    g262_p,
    n358_lo_n
  );


  and

  (
    g265_p,
    g264_n,
    g263_n
  );


  and

  (
    g266_p,
    g253_p_spl_1,
    n1251_o2_p_spl_00
  );


  or

  (
    g266_n,
    g253_n_spl_1,
    n1251_o2_n_spl_00
  );


  or

  (
    g267_n,
    g266_n,
    n370_lo_p
  );


  or

  (
    g268_n,
    g266_p,
    n370_lo_n
  );


  and

  (
    g269_p,
    g268_n,
    g267_n
  );


  and

  (
    g270_p,
    G354_o2_n,
    n1253_o2_p_spl_00
  );


  or

  (
    g270_n,
    G354_o2_p,
    n1253_o2_n_spl_00
  );


  and

  (
    g271_p,
    g270_p,
    n1254_o2_p_spl_00
  );


  or

  (
    g271_n,
    g270_n,
    n1254_o2_n_spl_00
  );


  and

  (
    g272_p,
    g271_p,
    G355_o2_n
  );


  or

  (
    g272_n,
    g271_n,
    G355_o2_p
  );


  and

  (
    g273_p,
    g272_p,
    G386_o2_p_spl_1
  );


  or

  (
    g273_n,
    g272_n,
    G386_o2_n_spl_1
  );


  and

  (
    g274_p,
    g273_p_spl_0,
    n1248_o2_p_spl_01
  );


  or

  (
    g274_n,
    g273_n_spl_0,
    n1248_o2_n_spl_01
  );


  or

  (
    g275_n,
    g274_n,
    n382_lo_p
  );


  or

  (
    g276_n,
    g274_p,
    n382_lo_n
  );


  and

  (
    g277_p,
    g276_n,
    g275_n
  );


  and

  (
    g278_p,
    g273_p_spl_0,
    n1249_o2_p_spl_01
  );


  or

  (
    g278_n,
    g273_n_spl_0,
    n1249_o2_n_spl_01
  );


  or

  (
    g279_n,
    g278_n,
    n394_lo_p
  );


  or

  (
    g280_n,
    g278_p,
    n394_lo_n
  );


  and

  (
    g281_p,
    g280_n,
    g279_n
  );


  and

  (
    g282_p,
    g273_p_spl_1,
    n1250_o2_p_spl_01
  );


  or

  (
    g282_n,
    g273_n_spl_1,
    n1250_o2_n_spl_01
  );


  or

  (
    g283_n,
    g282_n,
    n406_lo_p
  );


  or

  (
    g284_n,
    g282_p,
    n406_lo_n
  );


  and

  (
    g285_p,
    g284_n,
    g283_n
  );


  and

  (
    g286_p,
    g273_p_spl_1,
    n1251_o2_p_spl_01
  );


  or

  (
    g286_n,
    g273_n_spl_1,
    n1251_o2_n_spl_01
  );


  or

  (
    g287_n,
    g286_n,
    n418_lo_p
  );


  or

  (
    g288_n,
    g286_p,
    n418_lo_n
  );


  and

  (
    g289_p,
    g288_n,
    g287_n
  );


  and

  (
    g290_p,
    G356_o2_n,
    n1253_o2_p_spl_00
  );


  or

  (
    g290_n,
    G356_o2_p,
    n1253_o2_n_spl_00
  );


  and

  (
    g291_p,
    g290_p,
    G357_o2_n
  );


  or

  (
    g291_n,
    g290_n,
    G357_o2_p
  );


  and

  (
    g292_p,
    g291_p,
    n1255_o2_p_spl_00
  );


  or

  (
    g292_n,
    g291_n,
    n1255_o2_n_spl_00
  );


  and

  (
    g293_p,
    g292_p,
    G386_o2_p_spl_1
  );


  or

  (
    g293_n,
    g292_n,
    G386_o2_n_spl_1
  );


  and

  (
    g294_p,
    g293_p_spl_0,
    n1248_o2_p_spl_01
  );


  or

  (
    g294_n,
    g293_n_spl_0,
    n1248_o2_n_spl_01
  );


  or

  (
    g295_n,
    g294_n,
    n430_lo_p
  );


  or

  (
    g296_n,
    g294_p,
    n430_lo_n
  );


  and

  (
    g297_p,
    g296_n,
    g295_n
  );


  and

  (
    g298_p,
    g293_p_spl_0,
    n1249_o2_p_spl_01
  );


  or

  (
    g298_n,
    g293_n_spl_0,
    n1249_o2_n_spl_01
  );


  or

  (
    g299_n,
    g298_n,
    n442_lo_p
  );


  or

  (
    g300_n,
    g298_p,
    n442_lo_n
  );


  and

  (
    g301_p,
    g300_n,
    g299_n
  );


  and

  (
    g302_p,
    g293_p_spl_1,
    n1250_o2_p_spl_01
  );


  or

  (
    g302_n,
    g293_n_spl_1,
    n1250_o2_n_spl_01
  );


  or

  (
    g303_n,
    g302_n,
    n454_lo_p
  );


  or

  (
    g304_n,
    g302_p,
    n454_lo_n
  );


  and

  (
    g305_p,
    g304_n,
    g303_n
  );


  and

  (
    g306_p,
    g293_p_spl_1,
    n1251_o2_p_spl_01
  );


  or

  (
    g306_n,
    g293_n_spl_1,
    n1251_o2_n_spl_01
  );


  or

  (
    g307_n,
    g306_n,
    n466_lo_p
  );


  or

  (
    g308_n,
    g306_p,
    n466_lo_n
  );


  and

  (
    g309_p,
    g308_n,
    g307_n
  );


  and

  (
    g310_p,
    G370_o2_n,
    n1248_o2_p_spl_1
  );


  or

  (
    g310_n,
    G370_o2_p,
    n1248_o2_n_spl_1
  );


  and

  (
    g311_p,
    g310_p,
    n1250_o2_p_spl_1
  );


  or

  (
    g311_n,
    g310_n,
    n1250_o2_n_spl_1
  );


  and

  (
    g312_p,
    g311_p,
    G371_o2_n
  );


  or

  (
    g312_n,
    g311_n,
    G371_o2_p
  );


  and

  (
    g313_p,
    g312_p,
    G391_o2_p_spl_0
  );


  or

  (
    g313_n,
    g312_n,
    G391_o2_n_spl_0
  );


  and

  (
    g314_p,
    g313_p_spl_0,
    n1252_o2_p_spl_01
  );


  or

  (
    g314_n,
    g313_n_spl_0,
    n1252_o2_n_spl_01
  );


  or

  (
    g315_n,
    g314_n,
    n478_lo_p
  );


  or

  (
    g316_n,
    g314_p,
    n478_lo_n
  );


  and

  (
    g317_p,
    g316_n,
    g315_n
  );


  and

  (
    g318_p,
    g313_p_spl_0,
    n1253_o2_p_spl_01
  );


  or

  (
    g318_n,
    g313_n_spl_0,
    n1253_o2_n_spl_01
  );


  or

  (
    g319_n,
    g318_n,
    n490_lo_p
  );


  or

  (
    g320_n,
    g318_p,
    n490_lo_n
  );


  and

  (
    g321_p,
    g320_n,
    g319_n
  );


  and

  (
    g322_p,
    g313_p_spl_1,
    n1254_o2_p_spl_01
  );


  or

  (
    g322_n,
    g313_n_spl_1,
    n1254_o2_n_spl_01
  );


  or

  (
    g323_n,
    g322_n,
    n502_lo_p
  );


  or

  (
    g324_n,
    g322_p,
    n502_lo_n
  );


  and

  (
    g325_p,
    g324_n,
    g323_n
  );


  and

  (
    g326_p,
    g313_p_spl_1,
    n1255_o2_p_spl_01
  );


  or

  (
    g326_n,
    g313_n_spl_1,
    n1255_o2_n_spl_01
  );


  or

  (
    g327_n,
    g326_n,
    n514_lo_p
  );


  or

  (
    g328_n,
    g326_p,
    n514_lo_n
  );


  and

  (
    g329_p,
    g328_n,
    g327_n
  );


  and

  (
    g330_p,
    G372_o2_n,
    n1248_o2_p_spl_1
  );


  or

  (
    g330_n,
    G372_o2_p,
    n1248_o2_n_spl_1
  );


  and

  (
    g331_p,
    g330_p,
    G373_o2_n
  );


  or

  (
    g331_n,
    g330_n,
    G373_o2_p
  );


  and

  (
    g332_p,
    g331_p,
    n1251_o2_p_spl_1
  );


  or

  (
    g332_n,
    g331_n,
    n1251_o2_n_spl_1
  );


  and

  (
    g333_p,
    g332_p,
    G391_o2_p_spl_0
  );


  or

  (
    g333_n,
    g332_n,
    G391_o2_n_spl_0
  );


  and

  (
    g334_p,
    g333_p_spl_0,
    n1252_o2_p_spl_01
  );


  or

  (
    g334_n,
    g333_n_spl_0,
    n1252_o2_n_spl_01
  );


  or

  (
    g335_n,
    g334_n,
    n526_lo_p
  );


  or

  (
    g336_n,
    g334_p,
    n526_lo_n
  );


  and

  (
    g337_p,
    g336_n,
    g335_n
  );


  and

  (
    g338_p,
    g333_p_spl_0,
    n1253_o2_p_spl_01
  );


  or

  (
    g338_n,
    g333_n_spl_0,
    n1253_o2_n_spl_01
  );


  or

  (
    g339_n,
    g338_n,
    n538_lo_p
  );


  or

  (
    g340_n,
    g338_p,
    n538_lo_n
  );


  and

  (
    g341_p,
    g340_n,
    g339_n
  );


  and

  (
    g342_p,
    g333_p_spl_1,
    n1254_o2_p_spl_01
  );


  or

  (
    g342_n,
    g333_n_spl_1,
    n1254_o2_n_spl_01
  );


  or

  (
    g343_n,
    g342_n,
    n550_lo_p
  );


  or

  (
    g344_n,
    g342_p,
    n550_lo_n
  );


  and

  (
    g345_p,
    g344_n,
    g343_n
  );


  and

  (
    g346_p,
    g333_p_spl_1,
    n1255_o2_p_spl_01
  );


  or

  (
    g346_n,
    g333_n_spl_1,
    n1255_o2_n_spl_01
  );


  or

  (
    g347_n,
    g346_n,
    n562_lo_p
  );


  or

  (
    g348_n,
    g346_p,
    n562_lo_n
  );


  and

  (
    g349_p,
    g348_n,
    g347_n
  );


  and

  (
    g350_p,
    G374_o2_n,
    n1249_o2_p_spl_1
  );


  or

  (
    g350_n,
    G374_o2_p,
    n1249_o2_n_spl_1
  );


  and

  (
    g351_p,
    g350_p,
    n1250_o2_p_spl_1
  );


  or

  (
    g351_n,
    g350_n,
    n1250_o2_n_spl_1
  );


  and

  (
    g352_p,
    g351_p,
    G375_o2_n
  );


  or

  (
    g352_n,
    g351_n,
    G375_o2_p
  );


  and

  (
    g353_p,
    g352_p,
    G391_o2_p_spl_1
  );


  or

  (
    g353_n,
    g352_n,
    G391_o2_n_spl_1
  );


  and

  (
    g354_p,
    g353_p_spl_0,
    n1252_o2_p_spl_1
  );


  or

  (
    g354_n,
    g353_n_spl_0,
    n1252_o2_n_spl_1
  );


  or

  (
    g355_n,
    g354_n,
    n574_lo_p
  );


  or

  (
    g356_n,
    g354_p,
    n574_lo_n
  );


  and

  (
    g357_p,
    g356_n,
    g355_n
  );


  and

  (
    g358_p,
    g353_p_spl_0,
    n1253_o2_p_spl_1
  );


  or

  (
    g358_n,
    g353_n_spl_0,
    n1253_o2_n_spl_1
  );


  or

  (
    g359_n,
    g358_n,
    n586_lo_p
  );


  or

  (
    g360_n,
    g358_p,
    n586_lo_n
  );


  and

  (
    g361_p,
    g360_n,
    g359_n
  );


  and

  (
    g362_p,
    g353_p_spl_1,
    n1254_o2_p_spl_1
  );


  or

  (
    g362_n,
    g353_n_spl_1,
    n1254_o2_n_spl_1
  );


  or

  (
    g363_n,
    g362_n,
    n598_lo_p
  );


  or

  (
    g364_n,
    g362_p,
    n598_lo_n
  );


  and

  (
    g365_p,
    g364_n,
    g363_n
  );


  and

  (
    g366_p,
    g353_p_spl_1,
    n1255_o2_p_spl_1
  );


  or

  (
    g366_n,
    g353_n_spl_1,
    n1255_o2_n_spl_1
  );


  or

  (
    g367_n,
    g366_n,
    n610_lo_p
  );


  or

  (
    g368_n,
    g366_p,
    n610_lo_n
  );


  and

  (
    g369_p,
    g368_n,
    g367_n
  );


  and

  (
    g370_p,
    G376_o2_n,
    n1249_o2_p_spl_1
  );


  or

  (
    g370_n,
    G376_o2_p,
    n1249_o2_n_spl_1
  );


  and

  (
    g371_p,
    g370_p,
    G377_o2_n
  );


  or

  (
    g371_n,
    g370_n,
    G377_o2_p
  );


  and

  (
    g372_p,
    g371_p,
    n1251_o2_p_spl_1
  );


  or

  (
    g372_n,
    g371_n,
    n1251_o2_n_spl_1
  );


  and

  (
    g373_p,
    g372_p,
    G391_o2_p_spl_1
  );


  or

  (
    g373_n,
    g372_n,
    G391_o2_n_spl_1
  );


  and

  (
    g374_p,
    g373_p_spl_0,
    n1252_o2_p_spl_1
  );


  or

  (
    g374_n,
    g373_n_spl_0,
    n1252_o2_n_spl_1
  );


  or

  (
    g375_n,
    g374_n,
    n622_lo_p
  );


  or

  (
    g376_n,
    g374_p,
    n622_lo_n
  );


  and

  (
    g377_p,
    g376_n,
    g375_n
  );


  and

  (
    g378_p,
    g373_p_spl_0,
    n1253_o2_p_spl_1
  );


  or

  (
    g378_n,
    g373_n_spl_0,
    n1253_o2_n_spl_1
  );


  or

  (
    g379_n,
    g378_n,
    n634_lo_p
  );


  or

  (
    g380_n,
    g378_p,
    n634_lo_n
  );


  and

  (
    g381_p,
    g380_n,
    g379_n
  );


  and

  (
    g382_p,
    g373_p_spl_1,
    n1254_o2_p_spl_1
  );


  or

  (
    g382_n,
    g373_n_spl_1,
    n1254_o2_n_spl_1
  );


  or

  (
    g383_n,
    g382_n,
    n646_lo_p
  );


  or

  (
    g384_n,
    g382_p,
    n646_lo_n
  );


  and

  (
    g385_p,
    g384_n,
    g383_n
  );


  and

  (
    g386_p,
    g373_p_spl_1,
    n1255_o2_p_spl_1
  );


  or

  (
    g386_n,
    g373_n_spl_1,
    n1255_o2_n_spl_1
  );


  or

  (
    g387_n,
    g386_n,
    n658_lo_p
  );


  or

  (
    g388_n,
    g386_p,
    n658_lo_n
  );


  and

  (
    g389_p,
    g388_n,
    g387_n
  );


  or

  (
    g390_n,
    G247_o2_p_spl_,
    G234_o2_p_spl_
  );


  or

  (
    g391_n,
    g390_n_spl_,
    G260_o2_p_spl_0
  );


  or

  (
    g392_n,
    g391_n,
    G273_o2_n_spl_0
  );


  or

  (
    g393_n,
    g390_n_spl_,
    G260_o2_n_spl_0
  );


  or

  (
    g394_n,
    g393_n,
    G273_o2_p_spl_0
  );


  or

  (
    g395_n,
    G247_o2_n_spl_0,
    G234_o2_p_spl_
  );


  or

  (
    g396_n,
    g395_n,
    G260_o2_p_spl_0
  );


  or

  (
    g397_n,
    g396_n,
    G273_o2_p_spl_0
  );


  or

  (
    g398_n,
    G247_o2_p_spl_,
    G234_o2_n_spl_0
  );


  or

  (
    g399_n,
    g398_n,
    G260_o2_p_spl_
  );


  or

  (
    g400_n,
    g399_n,
    G273_o2_p_spl_
  );


  and

  (
    g401_p,
    g394_n,
    g392_n
  );


  and

  (
    g402_p,
    g401_p,
    g397_n
  );


  and

  (
    g403_p,
    g402_p,
    g400_n
  );


  or

  (
    g404_n,
    G299_o2_p_spl_,
    G286_o2_p_spl_
  );


  or

  (
    g405_n,
    g404_n_spl_,
    G312_o2_p_spl_0
  );


  or

  (
    g406_n,
    g405_n,
    G325_o2_n_spl_0
  );


  or

  (
    g407_n,
    g404_n_spl_,
    G312_o2_n_spl_0
  );


  or

  (
    g408_n,
    g407_n,
    G325_o2_p_spl_0
  );


  or

  (
    g409_n,
    G299_o2_n_spl_0,
    G286_o2_p_spl_
  );


  or

  (
    g410_n,
    g409_n,
    G312_o2_p_spl_0
  );


  or

  (
    g411_n,
    g410_n,
    G325_o2_p_spl_0
  );


  or

  (
    g412_n,
    G299_o2_p_spl_,
    G286_o2_n_spl_0
  );


  or

  (
    g413_n,
    g412_n,
    G312_o2_p_spl_
  );


  or

  (
    g414_n,
    g413_n,
    G325_o2_p_spl_
  );


  and

  (
    g415_p,
    g408_n,
    g406_n
  );


  and

  (
    g416_p,
    g415_p,
    g411_n
  );


  and

  (
    g417_p,
    g416_p,
    g414_n
  );


  and

  (
    g418_p,
    n331_lo_buf_o2_p_spl_,
    n283_lo_buf_o2_n_spl_0
  );


  or

  (
    g418_n,
    n331_lo_buf_o2_n_spl_0,
    n283_lo_buf_o2_p_spl_
  );


  and

  (
    g419_p,
    n331_lo_buf_o2_n_spl_0,
    n283_lo_buf_o2_p_spl_
  );


  or

  (
    g419_n,
    n331_lo_buf_o2_p_spl_,
    n283_lo_buf_o2_n_spl_0
  );


  and

  (
    g420_p,
    g419_n,
    g418_n
  );


  or

  (
    g420_n,
    g419_p,
    g418_p
  );


  and

  (
    g421_p,
    n427_lo_buf_o2_p_spl_,
    n379_lo_buf_o2_n_spl_0
  );


  or

  (
    g421_n,
    n427_lo_buf_o2_n_spl_0,
    n379_lo_buf_o2_p_spl_
  );


  and

  (
    g422_p,
    n427_lo_buf_o2_n_spl_0,
    n379_lo_buf_o2_p_spl_
  );


  or

  (
    g422_n,
    n427_lo_buf_o2_p_spl_,
    n379_lo_buf_o2_n_spl_0
  );


  and

  (
    g423_p,
    g422_n,
    g421_n
  );


  or

  (
    g423_n,
    g422_p,
    g421_p
  );


  and

  (
    g424_p,
    g423_n_spl_,
    g420_p_spl_
  );


  or

  (
    g424_n,
    g423_p_spl_,
    g420_n_spl_
  );


  and

  (
    g425_p,
    g423_p_spl_,
    g420_n_spl_
  );


  or

  (
    g425_n,
    g423_n_spl_,
    g420_p_spl_
  );


  and

  (
    g426_p,
    g425_n,
    g424_n
  );


  or

  (
    g426_n,
    g425_p,
    g424_p
  );


  and

  (
    g427_p,
    n763_lo_buf_o2_p_spl_00,
    n667_lo_buf_o2_p
  );


  or

  (
    g427_n,
    n763_lo_buf_o2_n_spl_00,
    n667_lo_buf_o2_n
  );


  and

  (
    g428_p,
    G201_o2_p_spl_0,
    G198_o2_n_spl_0
  );


  or

  (
    g428_n,
    G201_o2_n_spl_0,
    G198_o2_p_spl_0
  );


  and

  (
    g429_p,
    G201_o2_n_spl_0,
    G198_o2_p_spl_0
  );


  or

  (
    g429_n,
    G201_o2_p_spl_0,
    G198_o2_n_spl_0
  );


  and

  (
    g430_p,
    g429_n,
    g428_n
  );


  or

  (
    g430_n,
    g429_p,
    g428_p
  );


  and

  (
    g431_p,
    g430_n_spl_,
    g427_n_spl_
  );


  or

  (
    g431_n,
    g430_p_spl_,
    g427_p_spl_
  );


  and

  (
    g432_p,
    g430_p_spl_,
    g427_p_spl_
  );


  or

  (
    g432_n,
    g430_n_spl_,
    g427_n_spl_
  );


  and

  (
    g433_p,
    g432_n,
    g431_n
  );


  or

  (
    g433_n,
    g432_p,
    g431_p
  );


  or

  (
    g434_n,
    g433_p,
    g426_n
  );


  or

  (
    g435_n,
    g433_n,
    g426_p
  );


  and

  (
    g436_p,
    g435_n,
    g434_n
  );


  and

  (
    g437_p,
    n343_lo_buf_o2_p_spl_,
    n295_lo_buf_o2_n_spl_0
  );


  or

  (
    g437_n,
    n343_lo_buf_o2_n_spl_0,
    n295_lo_buf_o2_p_spl_
  );


  and

  (
    g438_p,
    n343_lo_buf_o2_n_spl_0,
    n295_lo_buf_o2_p_spl_
  );


  or

  (
    g438_n,
    n343_lo_buf_o2_p_spl_,
    n295_lo_buf_o2_n_spl_0
  );


  and

  (
    g439_p,
    g438_n,
    g437_n
  );


  or

  (
    g439_n,
    g438_p,
    g437_p
  );


  and

  (
    g440_p,
    n439_lo_buf_o2_p_spl_,
    n391_lo_buf_o2_n_spl_0
  );


  or

  (
    g440_n,
    n439_lo_buf_o2_n_spl_0,
    n391_lo_buf_o2_p_spl_
  );


  and

  (
    g441_p,
    n439_lo_buf_o2_n_spl_0,
    n391_lo_buf_o2_p_spl_
  );


  or

  (
    g441_n,
    n439_lo_buf_o2_p_spl_,
    n391_lo_buf_o2_n_spl_0
  );


  and

  (
    g442_p,
    g441_n,
    g440_n
  );


  or

  (
    g442_n,
    g441_p,
    g440_p
  );


  and

  (
    g443_p,
    g442_n_spl_,
    g439_p_spl_
  );


  or

  (
    g443_n,
    g442_p_spl_,
    g439_n_spl_
  );


  and

  (
    g444_p,
    g442_p_spl_,
    g439_n_spl_
  );


  or

  (
    g444_n,
    g442_n_spl_,
    g439_p_spl_
  );


  and

  (
    g445_p,
    g444_n,
    g443_n
  );


  or

  (
    g445_n,
    g444_p,
    g443_p
  );


  and

  (
    g446_p,
    n763_lo_buf_o2_p_spl_00,
    n679_lo_buf_o2_p
  );


  or

  (
    g446_n,
    n763_lo_buf_o2_n_spl_00,
    n679_lo_buf_o2_n
  );


  and

  (
    g447_p,
    G207_o2_p_spl_0,
    G204_o2_n_spl_0
  );


  or

  (
    g447_n,
    G207_o2_n_spl_0,
    G204_o2_p_spl_0
  );


  and

  (
    g448_p,
    G207_o2_n_spl_0,
    G204_o2_p_spl_0
  );


  or

  (
    g448_n,
    G207_o2_p_spl_0,
    G204_o2_n_spl_0
  );


  and

  (
    g449_p,
    g448_n,
    g447_n
  );


  or

  (
    g449_n,
    g448_p,
    g447_p
  );


  and

  (
    g450_p,
    g449_n_spl_,
    g446_n_spl_
  );


  or

  (
    g450_n,
    g449_p_spl_,
    g446_p_spl_
  );


  and

  (
    g451_p,
    g449_p_spl_,
    g446_p_spl_
  );


  or

  (
    g451_n,
    g449_n_spl_,
    g446_n_spl_
  );


  and

  (
    g452_p,
    g451_n,
    g450_n
  );


  or

  (
    g452_n,
    g451_p,
    g450_p
  );


  or

  (
    g453_n,
    g452_p,
    g445_n
  );


  or

  (
    g454_n,
    g452_n,
    g445_p
  );


  and

  (
    g455_p,
    g454_n,
    g453_n
  );


  and

  (
    g456_p,
    n355_lo_buf_o2_p_spl_,
    n307_lo_buf_o2_n_spl_0
  );


  or

  (
    g456_n,
    n355_lo_buf_o2_n_spl_0,
    n307_lo_buf_o2_p_spl_
  );


  and

  (
    g457_p,
    n355_lo_buf_o2_n_spl_0,
    n307_lo_buf_o2_p_spl_
  );


  or

  (
    g457_n,
    n355_lo_buf_o2_p_spl_,
    n307_lo_buf_o2_n_spl_0
  );


  and

  (
    g458_p,
    g457_n,
    g456_n
  );


  or

  (
    g458_n,
    g457_p,
    g456_p
  );


  and

  (
    g459_p,
    n451_lo_buf_o2_p_spl_,
    n403_lo_buf_o2_n_spl_0
  );


  or

  (
    g459_n,
    n451_lo_buf_o2_n_spl_0,
    n403_lo_buf_o2_p_spl_
  );


  and

  (
    g460_p,
    n451_lo_buf_o2_n_spl_0,
    n403_lo_buf_o2_p_spl_
  );


  or

  (
    g460_n,
    n451_lo_buf_o2_p_spl_,
    n403_lo_buf_o2_n_spl_0
  );


  and

  (
    g461_p,
    g460_n,
    g459_n
  );


  or

  (
    g461_n,
    g460_p,
    g459_p
  );


  and

  (
    g462_p,
    g461_n_spl_,
    g458_p_spl_
  );


  or

  (
    g462_n,
    g461_p_spl_,
    g458_n_spl_
  );


  and

  (
    g463_p,
    g461_p_spl_,
    g458_n_spl_
  );


  or

  (
    g463_n,
    g461_n_spl_,
    g458_p_spl_
  );


  and

  (
    g464_p,
    g463_n,
    g462_n
  );


  or

  (
    g464_n,
    g463_p,
    g462_p
  );


  and

  (
    g465_p,
    n763_lo_buf_o2_p_spl_01,
    n691_lo_buf_o2_p
  );


  or

  (
    g465_n,
    n763_lo_buf_o2_n_spl_01,
    n691_lo_buf_o2_n
  );


  and

  (
    g466_p,
    G204_o2_p_spl_1,
    G198_o2_n_spl_1
  );


  or

  (
    g466_n,
    G204_o2_n_spl_1,
    G198_o2_p_spl_1
  );


  and

  (
    g467_p,
    G204_o2_n_spl_1,
    G198_o2_p_spl_1
  );


  or

  (
    g467_n,
    G204_o2_p_spl_1,
    G198_o2_n_spl_1
  );


  and

  (
    g468_p,
    g467_n,
    g466_n
  );


  or

  (
    g468_n,
    g467_p,
    g466_p
  );


  and

  (
    g469_p,
    g468_n_spl_,
    g465_n_spl_
  );


  or

  (
    g469_n,
    g468_p_spl_,
    g465_p_spl_
  );


  and

  (
    g470_p,
    g468_p_spl_,
    g465_p_spl_
  );


  or

  (
    g470_n,
    g468_n_spl_,
    g465_n_spl_
  );


  and

  (
    g471_p,
    g470_n,
    g469_n
  );


  or

  (
    g471_n,
    g470_p,
    g469_p
  );


  or

  (
    g472_n,
    g471_p,
    g464_n
  );


  or

  (
    g473_n,
    g471_n,
    g464_p
  );


  and

  (
    g474_p,
    g473_n,
    g472_n
  );


  and

  (
    g475_p,
    n367_lo_buf_o2_p_spl_,
    n319_lo_buf_o2_n_spl_0
  );


  or

  (
    g475_n,
    n367_lo_buf_o2_n_spl_0,
    n319_lo_buf_o2_p_spl_
  );


  and

  (
    g476_p,
    n367_lo_buf_o2_n_spl_0,
    n319_lo_buf_o2_p_spl_
  );


  or

  (
    g476_n,
    n367_lo_buf_o2_p_spl_,
    n319_lo_buf_o2_n_spl_0
  );


  and

  (
    g477_p,
    g476_n,
    g475_n
  );


  or

  (
    g477_n,
    g476_p,
    g475_p
  );


  and

  (
    g478_p,
    n463_lo_buf_o2_p_spl_,
    n415_lo_buf_o2_n_spl_0
  );


  or

  (
    g478_n,
    n463_lo_buf_o2_n_spl_0,
    n415_lo_buf_o2_p_spl_
  );


  and

  (
    g479_p,
    n463_lo_buf_o2_n_spl_0,
    n415_lo_buf_o2_p_spl_
  );


  or

  (
    g479_n,
    n463_lo_buf_o2_p_spl_,
    n415_lo_buf_o2_n_spl_0
  );


  and

  (
    g480_p,
    g479_n,
    g478_n
  );


  or

  (
    g480_n,
    g479_p,
    g478_p
  );


  and

  (
    g481_p,
    g480_n_spl_,
    g477_p_spl_
  );


  or

  (
    g481_n,
    g480_p_spl_,
    g477_n_spl_
  );


  and

  (
    g482_p,
    g480_p_spl_,
    g477_n_spl_
  );


  or

  (
    g482_n,
    g480_n_spl_,
    g477_p_spl_
  );


  and

  (
    g483_p,
    g482_n,
    g481_n
  );


  or

  (
    g483_n,
    g482_p,
    g481_p
  );


  and

  (
    g484_p,
    n763_lo_buf_o2_p_spl_01,
    n703_lo_buf_o2_p
  );


  or

  (
    g484_n,
    n763_lo_buf_o2_n_spl_01,
    n703_lo_buf_o2_n
  );


  and

  (
    g485_p,
    G207_o2_p_spl_1,
    G201_o2_n_spl_1
  );


  or

  (
    g485_n,
    G207_o2_n_spl_1,
    G201_o2_p_spl_1
  );


  and

  (
    g486_p,
    G207_o2_n_spl_1,
    G201_o2_p_spl_1
  );


  or

  (
    g486_n,
    G207_o2_p_spl_1,
    G201_o2_n_spl_1
  );


  and

  (
    g487_p,
    g486_n,
    g485_n
  );


  or

  (
    g487_n,
    g486_p,
    g485_p
  );


  and

  (
    g488_p,
    g487_n_spl_,
    g484_n_spl_
  );


  or

  (
    g488_n,
    g487_p_spl_,
    g484_p_spl_
  );


  and

  (
    g489_p,
    g487_p_spl_,
    g484_p_spl_
  );


  or

  (
    g489_n,
    g487_n_spl_,
    g484_n_spl_
  );


  and

  (
    g490_p,
    g489_n,
    g488_n
  );


  or

  (
    g490_n,
    g489_p,
    g488_p
  );


  or

  (
    g491_n,
    g490_p,
    g483_n
  );


  or

  (
    g492_n,
    g490_n,
    g483_p
  );


  and

  (
    g493_p,
    g492_n,
    g491_n
  );


  and

  (
    g494_p,
    n523_lo_buf_o2_p_spl_,
    n475_lo_buf_o2_n_spl_0
  );


  or

  (
    g494_n,
    n523_lo_buf_o2_n_spl_0,
    n475_lo_buf_o2_p_spl_
  );


  and

  (
    g495_p,
    n523_lo_buf_o2_n_spl_0,
    n475_lo_buf_o2_p_spl_
  );


  or

  (
    g495_n,
    n523_lo_buf_o2_p_spl_,
    n475_lo_buf_o2_n_spl_0
  );


  and

  (
    g496_p,
    g495_n,
    g494_n
  );


  or

  (
    g496_n,
    g495_p,
    g494_p
  );


  and

  (
    g497_p,
    n619_lo_buf_o2_p_spl_,
    n571_lo_buf_o2_n_spl_0
  );


  or

  (
    g497_n,
    n619_lo_buf_o2_n_spl_0,
    n571_lo_buf_o2_p_spl_
  );


  and

  (
    g498_p,
    n619_lo_buf_o2_n_spl_0,
    n571_lo_buf_o2_p_spl_
  );


  or

  (
    g498_n,
    n619_lo_buf_o2_p_spl_,
    n571_lo_buf_o2_n_spl_0
  );


  and

  (
    g499_p,
    g498_n,
    g497_n
  );


  or

  (
    g499_n,
    g498_p,
    g497_p
  );


  and

  (
    g500_p,
    g499_n_spl_,
    g496_p_spl_
  );


  or

  (
    g500_n,
    g499_p_spl_,
    g496_n_spl_
  );


  and

  (
    g501_p,
    g499_p_spl_,
    g496_n_spl_
  );


  or

  (
    g501_n,
    g499_n_spl_,
    g496_p_spl_
  );


  and

  (
    g502_p,
    g501_n,
    g500_n
  );


  or

  (
    g502_n,
    g501_p,
    g500_p
  );


  and

  (
    g503_p,
    n763_lo_buf_o2_p_spl_10,
    n715_lo_buf_o2_p
  );


  or

  (
    g503_n,
    n763_lo_buf_o2_n_spl_10,
    n715_lo_buf_o2_n
  );


  and

  (
    g504_p,
    G189_o2_p_spl_0,
    G186_o2_n_spl_0
  );


  or

  (
    g504_n,
    G189_o2_n_spl_0,
    G186_o2_p_spl_0
  );


  and

  (
    g505_p,
    G189_o2_n_spl_0,
    G186_o2_p_spl_0
  );


  or

  (
    g505_n,
    G189_o2_p_spl_0,
    G186_o2_n_spl_0
  );


  and

  (
    g506_p,
    g505_n,
    g504_n
  );


  or

  (
    g506_n,
    g505_p,
    g504_p
  );


  and

  (
    g507_p,
    g506_n_spl_,
    g503_n_spl_
  );


  or

  (
    g507_n,
    g506_p_spl_,
    g503_p_spl_
  );


  and

  (
    g508_p,
    g506_p_spl_,
    g503_p_spl_
  );


  or

  (
    g508_n,
    g506_n_spl_,
    g503_n_spl_
  );


  and

  (
    g509_p,
    g508_n,
    g507_n
  );


  or

  (
    g509_n,
    g508_p,
    g507_p
  );


  or

  (
    g510_n,
    g509_p,
    g502_n
  );


  or

  (
    g511_n,
    g509_n,
    g502_p
  );


  and

  (
    g512_p,
    g511_n,
    g510_n
  );


  and

  (
    g513_p,
    n535_lo_buf_o2_p_spl_,
    n487_lo_buf_o2_n_spl_0
  );


  or

  (
    g513_n,
    n535_lo_buf_o2_n_spl_0,
    n487_lo_buf_o2_p_spl_
  );


  and

  (
    g514_p,
    n535_lo_buf_o2_n_spl_0,
    n487_lo_buf_o2_p_spl_
  );


  or

  (
    g514_n,
    n535_lo_buf_o2_p_spl_,
    n487_lo_buf_o2_n_spl_0
  );


  and

  (
    g515_p,
    g514_n,
    g513_n
  );


  or

  (
    g515_n,
    g514_p,
    g513_p
  );


  and

  (
    g516_p,
    n631_lo_buf_o2_p_spl_,
    n583_lo_buf_o2_n_spl_0
  );


  or

  (
    g516_n,
    n631_lo_buf_o2_n_spl_0,
    n583_lo_buf_o2_p_spl_
  );


  and

  (
    g517_p,
    n631_lo_buf_o2_n_spl_0,
    n583_lo_buf_o2_p_spl_
  );


  or

  (
    g517_n,
    n631_lo_buf_o2_p_spl_,
    n583_lo_buf_o2_n_spl_0
  );


  and

  (
    g518_p,
    g517_n,
    g516_n
  );


  or

  (
    g518_n,
    g517_p,
    g516_p
  );


  and

  (
    g519_p,
    g518_n_spl_,
    g515_p_spl_
  );


  or

  (
    g519_n,
    g518_p_spl_,
    g515_n_spl_
  );


  and

  (
    g520_p,
    g518_p_spl_,
    g515_n_spl_
  );


  or

  (
    g520_n,
    g518_n_spl_,
    g515_p_spl_
  );


  and

  (
    g521_p,
    g520_n,
    g519_n
  );


  or

  (
    g521_n,
    g520_p,
    g519_p
  );


  and

  (
    g522_p,
    n763_lo_buf_o2_p_spl_10,
    n727_lo_buf_o2_p
  );


  or

  (
    g522_n,
    n763_lo_buf_o2_n_spl_10,
    n727_lo_buf_o2_n
  );


  and

  (
    g523_p,
    G195_o2_p_spl_0,
    G192_o2_n_spl_0
  );


  or

  (
    g523_n,
    G195_o2_n_spl_0,
    G192_o2_p_spl_0
  );


  and

  (
    g524_p,
    G195_o2_n_spl_0,
    G192_o2_p_spl_0
  );


  or

  (
    g524_n,
    G195_o2_p_spl_0,
    G192_o2_n_spl_0
  );


  and

  (
    g525_p,
    g524_n,
    g523_n
  );


  or

  (
    g525_n,
    g524_p,
    g523_p
  );


  and

  (
    g526_p,
    g525_n_spl_,
    g522_n_spl_
  );


  or

  (
    g526_n,
    g525_p_spl_,
    g522_p_spl_
  );


  and

  (
    g527_p,
    g525_p_spl_,
    g522_p_spl_
  );


  or

  (
    g527_n,
    g525_n_spl_,
    g522_n_spl_
  );


  and

  (
    g528_p,
    g527_n,
    g526_n
  );


  or

  (
    g528_n,
    g527_p,
    g526_p
  );


  or

  (
    g529_n,
    g528_p,
    g521_n
  );


  or

  (
    g530_n,
    g528_n,
    g521_p
  );


  and

  (
    g531_p,
    g530_n,
    g529_n
  );


  and

  (
    g532_p,
    n547_lo_buf_o2_p_spl_,
    n499_lo_buf_o2_n_spl_0
  );


  or

  (
    g532_n,
    n547_lo_buf_o2_n_spl_0,
    n499_lo_buf_o2_p_spl_
  );


  and

  (
    g533_p,
    n547_lo_buf_o2_n_spl_0,
    n499_lo_buf_o2_p_spl_
  );


  or

  (
    g533_n,
    n547_lo_buf_o2_p_spl_,
    n499_lo_buf_o2_n_spl_0
  );


  and

  (
    g534_p,
    g533_n,
    g532_n
  );


  or

  (
    g534_n,
    g533_p,
    g532_p
  );


  and

  (
    g535_p,
    n643_lo_buf_o2_p_spl_,
    n595_lo_buf_o2_n_spl_0
  );


  or

  (
    g535_n,
    n643_lo_buf_o2_n_spl_0,
    n595_lo_buf_o2_p_spl_
  );


  and

  (
    g536_p,
    n643_lo_buf_o2_n_spl_0,
    n595_lo_buf_o2_p_spl_
  );


  or

  (
    g536_n,
    n643_lo_buf_o2_p_spl_,
    n595_lo_buf_o2_n_spl_0
  );


  and

  (
    g537_p,
    g536_n,
    g535_n
  );


  or

  (
    g537_n,
    g536_p,
    g535_p
  );


  and

  (
    g538_p,
    g537_n_spl_,
    g534_p_spl_
  );


  or

  (
    g538_n,
    g537_p_spl_,
    g534_n_spl_
  );


  and

  (
    g539_p,
    g537_p_spl_,
    g534_n_spl_
  );


  or

  (
    g539_n,
    g537_n_spl_,
    g534_p_spl_
  );


  and

  (
    g540_p,
    g539_n,
    g538_n
  );


  or

  (
    g540_n,
    g539_p,
    g538_p
  );


  and

  (
    g541_p,
    n763_lo_buf_o2_p_spl_11,
    n739_lo_buf_o2_p
  );


  or

  (
    g541_n,
    n763_lo_buf_o2_n_spl_11,
    n739_lo_buf_o2_n
  );


  and

  (
    g542_p,
    G192_o2_p_spl_1,
    G186_o2_n_spl_1
  );


  or

  (
    g542_n,
    G192_o2_n_spl_1,
    G186_o2_p_spl_1
  );


  and

  (
    g543_p,
    G192_o2_n_spl_1,
    G186_o2_p_spl_1
  );


  or

  (
    g543_n,
    G192_o2_p_spl_1,
    G186_o2_n_spl_1
  );


  and

  (
    g544_p,
    g543_n,
    g542_n
  );


  or

  (
    g544_n,
    g543_p,
    g542_p
  );


  and

  (
    g545_p,
    g544_n_spl_,
    g541_n_spl_
  );


  or

  (
    g545_n,
    g544_p_spl_,
    g541_p_spl_
  );


  and

  (
    g546_p,
    g544_p_spl_,
    g541_p_spl_
  );


  or

  (
    g546_n,
    g544_n_spl_,
    g541_n_spl_
  );


  and

  (
    g547_p,
    g546_n,
    g545_n
  );


  or

  (
    g547_n,
    g546_p,
    g545_p
  );


  or

  (
    g548_n,
    g547_p,
    g540_n
  );


  or

  (
    g549_n,
    g547_n,
    g540_p
  );


  and

  (
    g550_p,
    g549_n,
    g548_n
  );


  and

  (
    g551_p,
    n559_lo_buf_o2_p_spl_,
    n511_lo_buf_o2_n_spl_0
  );


  or

  (
    g551_n,
    n559_lo_buf_o2_n_spl_0,
    n511_lo_buf_o2_p_spl_
  );


  and

  (
    g552_p,
    n559_lo_buf_o2_n_spl_0,
    n511_lo_buf_o2_p_spl_
  );


  or

  (
    g552_n,
    n559_lo_buf_o2_p_spl_,
    n511_lo_buf_o2_n_spl_0
  );


  and

  (
    g553_p,
    g552_n,
    g551_n
  );


  or

  (
    g553_n,
    g552_p,
    g551_p
  );


  and

  (
    g554_p,
    n655_lo_buf_o2_p_spl_,
    n607_lo_buf_o2_n_spl_0
  );


  or

  (
    g554_n,
    n655_lo_buf_o2_n_spl_0,
    n607_lo_buf_o2_p_spl_
  );


  and

  (
    g555_p,
    n655_lo_buf_o2_n_spl_0,
    n607_lo_buf_o2_p_spl_
  );


  or

  (
    g555_n,
    n655_lo_buf_o2_p_spl_,
    n607_lo_buf_o2_n_spl_0
  );


  and

  (
    g556_p,
    g555_n,
    g554_n
  );


  or

  (
    g556_n,
    g555_p,
    g554_p
  );


  and

  (
    g557_p,
    g556_n_spl_,
    g553_p_spl_
  );


  or

  (
    g557_n,
    g556_p_spl_,
    g553_n_spl_
  );


  and

  (
    g558_p,
    g556_p_spl_,
    g553_n_spl_
  );


  or

  (
    g558_n,
    g556_n_spl_,
    g553_p_spl_
  );


  and

  (
    g559_p,
    g558_n,
    g557_n
  );


  or

  (
    g559_n,
    g558_p,
    g557_p
  );


  and

  (
    g560_p,
    n763_lo_buf_o2_p_spl_11,
    n751_lo_buf_o2_p
  );


  or

  (
    g560_n,
    n763_lo_buf_o2_n_spl_11,
    n751_lo_buf_o2_n
  );


  and

  (
    g561_p,
    G195_o2_p_spl_1,
    G189_o2_n_spl_1
  );


  or

  (
    g561_n,
    G195_o2_n_spl_1,
    G189_o2_p_spl_1
  );


  and

  (
    g562_p,
    G195_o2_n_spl_1,
    G189_o2_p_spl_1
  );


  or

  (
    g562_n,
    G195_o2_p_spl_1,
    G189_o2_n_spl_1
  );


  and

  (
    g563_p,
    g562_n,
    g561_n
  );


  or

  (
    g563_n,
    g562_p,
    g561_p
  );


  and

  (
    g564_p,
    g563_n_spl_,
    g560_n_spl_
  );


  or

  (
    g564_n,
    g563_p_spl_,
    g560_p_spl_
  );


  and

  (
    g565_p,
    g563_p_spl_,
    g560_p_spl_
  );


  or

  (
    g565_n,
    g563_n_spl_,
    g560_n_spl_
  );


  and

  (
    g566_p,
    g565_n,
    g564_n
  );


  or

  (
    g566_n,
    g565_p,
    g564_p
  );


  or

  (
    g567_n,
    g566_p,
    g559_n
  );


  or

  (
    g568_n,
    g566_n,
    g559_p
  );


  and

  (
    g569_p,
    g568_n,
    g567_n
  );


  and

  (
    g570_p,
    n292_lo_buf_o2_p_spl_,
    n280_lo_buf_o2_n_spl_0
  );


  or

  (
    g570_n,
    n292_lo_buf_o2_n_spl_0,
    n280_lo_buf_o2_p_spl_
  );


  and

  (
    g571_p,
    n292_lo_buf_o2_n_spl_0,
    n280_lo_buf_o2_p_spl_
  );


  or

  (
    g571_n,
    n292_lo_buf_o2_p_spl_,
    n280_lo_buf_o2_n_spl_0
  );


  and

  (
    g572_p,
    g571_n,
    g570_n
  );


  or

  (
    g572_n,
    g571_p,
    g570_p
  );


  and

  (
    g573_p,
    n316_lo_buf_o2_p_spl_,
    n304_lo_buf_o2_n_spl_0
  );


  or

  (
    g573_n,
    n316_lo_buf_o2_n_spl_0,
    n304_lo_buf_o2_p_spl_
  );


  and

  (
    g574_p,
    n316_lo_buf_o2_n_spl_0,
    n304_lo_buf_o2_p_spl_
  );


  or

  (
    g574_n,
    n316_lo_buf_o2_p_spl_,
    n304_lo_buf_o2_n_spl_0
  );


  and

  (
    g575_p,
    g574_n,
    g573_n
  );


  or

  (
    g575_n,
    g574_p,
    g573_p
  );


  or

  (
    g576_n,
    g575_p,
    g572_n
  );


  or

  (
    g577_n,
    g575_n,
    g572_p
  );


  and

  (
    g578_p,
    g577_n,
    g576_n
  );


  and

  (
    g579_p,
    n340_lo_buf_o2_p_spl_,
    n328_lo_buf_o2_n_spl_0
  );


  or

  (
    g579_n,
    n340_lo_buf_o2_n_spl_0,
    n328_lo_buf_o2_p_spl_
  );


  and

  (
    g580_p,
    n340_lo_buf_o2_n_spl_0,
    n328_lo_buf_o2_p_spl_
  );


  or

  (
    g580_n,
    n340_lo_buf_o2_p_spl_,
    n328_lo_buf_o2_n_spl_0
  );


  and

  (
    g581_p,
    g580_n,
    g579_n
  );


  or

  (
    g581_n,
    g580_p,
    g579_p
  );


  and

  (
    g582_p,
    n364_lo_buf_o2_p_spl_,
    n352_lo_buf_o2_n_spl_0
  );


  or

  (
    g582_n,
    n364_lo_buf_o2_n_spl_0,
    n352_lo_buf_o2_p_spl_
  );


  and

  (
    g583_p,
    n364_lo_buf_o2_n_spl_0,
    n352_lo_buf_o2_p_spl_
  );


  or

  (
    g583_n,
    n364_lo_buf_o2_p_spl_,
    n352_lo_buf_o2_n_spl_0
  );


  and

  (
    g584_p,
    g583_n,
    g582_n
  );


  or

  (
    g584_n,
    g583_p,
    g582_p
  );


  or

  (
    g585_n,
    g584_p,
    g581_n
  );


  or

  (
    g586_n,
    g584_n,
    g581_p
  );


  and

  (
    g587_p,
    g586_n,
    g585_n
  );


  and

  (
    g588_p,
    n388_lo_buf_o2_p_spl_,
    n376_lo_buf_o2_n_spl_0
  );


  or

  (
    g588_n,
    n388_lo_buf_o2_n_spl_0,
    n376_lo_buf_o2_p_spl_
  );


  and

  (
    g589_p,
    n388_lo_buf_o2_n_spl_0,
    n376_lo_buf_o2_p_spl_
  );


  or

  (
    g589_n,
    n388_lo_buf_o2_p_spl_,
    n376_lo_buf_o2_n_spl_0
  );


  and

  (
    g590_p,
    g589_n,
    g588_n
  );


  or

  (
    g590_n,
    g589_p,
    g588_p
  );


  and

  (
    g591_p,
    n412_lo_buf_o2_p_spl_,
    n400_lo_buf_o2_n_spl_0
  );


  or

  (
    g591_n,
    n412_lo_buf_o2_n_spl_0,
    n400_lo_buf_o2_p_spl_
  );


  and

  (
    g592_p,
    n412_lo_buf_o2_n_spl_0,
    n400_lo_buf_o2_p_spl_
  );


  or

  (
    g592_n,
    n412_lo_buf_o2_p_spl_,
    n400_lo_buf_o2_n_spl_0
  );


  and

  (
    g593_p,
    g592_n,
    g591_n
  );


  or

  (
    g593_n,
    g592_p,
    g591_p
  );


  or

  (
    g594_n,
    g593_p,
    g590_n
  );


  or

  (
    g595_n,
    g593_n,
    g590_p
  );


  and

  (
    g596_p,
    g595_n,
    g594_n
  );


  and

  (
    g597_p,
    n436_lo_buf_o2_p_spl_,
    n424_lo_buf_o2_n_spl_0
  );


  or

  (
    g597_n,
    n436_lo_buf_o2_n_spl_0,
    n424_lo_buf_o2_p_spl_
  );


  and

  (
    g598_p,
    n436_lo_buf_o2_n_spl_0,
    n424_lo_buf_o2_p_spl_
  );


  or

  (
    g598_n,
    n436_lo_buf_o2_p_spl_,
    n424_lo_buf_o2_n_spl_0
  );


  and

  (
    g599_p,
    g598_n,
    g597_n
  );


  or

  (
    g599_n,
    g598_p,
    g597_p
  );


  and

  (
    g600_p,
    n460_lo_buf_o2_p_spl_,
    n448_lo_buf_o2_n_spl_0
  );


  or

  (
    g600_n,
    n460_lo_buf_o2_n_spl_0,
    n448_lo_buf_o2_p_spl_
  );


  and

  (
    g601_p,
    n460_lo_buf_o2_n_spl_0,
    n448_lo_buf_o2_p_spl_
  );


  or

  (
    g601_n,
    n460_lo_buf_o2_p_spl_,
    n448_lo_buf_o2_n_spl_0
  );


  and

  (
    g602_p,
    g601_n,
    g600_n
  );


  or

  (
    g602_n,
    g601_p,
    g600_p
  );


  or

  (
    g603_n,
    g602_p,
    g599_n
  );


  or

  (
    g604_n,
    g602_n,
    g599_p
  );


  and

  (
    g605_p,
    g604_n,
    g603_n
  );


  and

  (
    g606_p,
    n484_lo_buf_o2_p_spl_,
    n472_lo_buf_o2_n_spl_0
  );


  or

  (
    g606_n,
    n484_lo_buf_o2_n_spl_0,
    n472_lo_buf_o2_p_spl_
  );


  and

  (
    g607_p,
    n484_lo_buf_o2_n_spl_0,
    n472_lo_buf_o2_p_spl_
  );


  or

  (
    g607_n,
    n484_lo_buf_o2_p_spl_,
    n472_lo_buf_o2_n_spl_0
  );


  and

  (
    g608_p,
    g607_n,
    g606_n
  );


  or

  (
    g608_n,
    g607_p,
    g606_p
  );


  and

  (
    g609_p,
    n508_lo_buf_o2_p_spl_,
    n496_lo_buf_o2_n_spl_0
  );


  or

  (
    g609_n,
    n508_lo_buf_o2_n_spl_0,
    n496_lo_buf_o2_p_spl_
  );


  and

  (
    g610_p,
    n508_lo_buf_o2_n_spl_0,
    n496_lo_buf_o2_p_spl_
  );


  or

  (
    g610_n,
    n508_lo_buf_o2_p_spl_,
    n496_lo_buf_o2_n_spl_0
  );


  and

  (
    g611_p,
    g610_n,
    g609_n
  );


  or

  (
    g611_n,
    g610_p,
    g609_p
  );


  or

  (
    g612_n,
    g611_p,
    g608_n
  );


  or

  (
    g613_n,
    g611_n,
    g608_p
  );


  and

  (
    g614_p,
    g613_n,
    g612_n
  );


  and

  (
    g615_p,
    n532_lo_buf_o2_p_spl_,
    n520_lo_buf_o2_n_spl_0
  );


  or

  (
    g615_n,
    n532_lo_buf_o2_n_spl_0,
    n520_lo_buf_o2_p_spl_
  );


  and

  (
    g616_p,
    n532_lo_buf_o2_n_spl_0,
    n520_lo_buf_o2_p_spl_
  );


  or

  (
    g616_n,
    n532_lo_buf_o2_p_spl_,
    n520_lo_buf_o2_n_spl_0
  );


  and

  (
    g617_p,
    g616_n,
    g615_n
  );


  or

  (
    g617_n,
    g616_p,
    g615_p
  );


  and

  (
    g618_p,
    n556_lo_buf_o2_p_spl_,
    n544_lo_buf_o2_n_spl_0
  );


  or

  (
    g618_n,
    n556_lo_buf_o2_n_spl_0,
    n544_lo_buf_o2_p_spl_
  );


  and

  (
    g619_p,
    n556_lo_buf_o2_n_spl_0,
    n544_lo_buf_o2_p_spl_
  );


  or

  (
    g619_n,
    n556_lo_buf_o2_p_spl_,
    n544_lo_buf_o2_n_spl_0
  );


  and

  (
    g620_p,
    g619_n,
    g618_n
  );


  or

  (
    g620_n,
    g619_p,
    g618_p
  );


  or

  (
    g621_n,
    g620_p,
    g617_n
  );


  or

  (
    g622_n,
    g620_n,
    g617_p
  );


  and

  (
    g623_p,
    g622_n,
    g621_n
  );


  and

  (
    g624_p,
    n580_lo_buf_o2_p_spl_,
    n568_lo_buf_o2_n_spl_0
  );


  or

  (
    g624_n,
    n580_lo_buf_o2_n_spl_0,
    n568_lo_buf_o2_p_spl_
  );


  and

  (
    g625_p,
    n580_lo_buf_o2_n_spl_0,
    n568_lo_buf_o2_p_spl_
  );


  or

  (
    g625_n,
    n580_lo_buf_o2_p_spl_,
    n568_lo_buf_o2_n_spl_0
  );


  and

  (
    g626_p,
    g625_n,
    g624_n
  );


  or

  (
    g626_n,
    g625_p,
    g624_p
  );


  and

  (
    g627_p,
    n604_lo_buf_o2_p_spl_,
    n592_lo_buf_o2_n_spl_0
  );


  or

  (
    g627_n,
    n604_lo_buf_o2_n_spl_0,
    n592_lo_buf_o2_p_spl_
  );


  and

  (
    g628_p,
    n604_lo_buf_o2_n_spl_0,
    n592_lo_buf_o2_p_spl_
  );


  or

  (
    g628_n,
    n604_lo_buf_o2_p_spl_,
    n592_lo_buf_o2_n_spl_0
  );


  and

  (
    g629_p,
    g628_n,
    g627_n
  );


  or

  (
    g629_n,
    g628_p,
    g627_p
  );


  or

  (
    g630_n,
    g629_p,
    g626_n
  );


  or

  (
    g631_n,
    g629_n,
    g626_p
  );


  and

  (
    g632_p,
    g631_n,
    g630_n
  );


  and

  (
    g633_p,
    n628_lo_buf_o2_p_spl_,
    n616_lo_buf_o2_n_spl_0
  );


  or

  (
    g633_n,
    n628_lo_buf_o2_n_spl_0,
    n616_lo_buf_o2_p_spl_
  );


  and

  (
    g634_p,
    n628_lo_buf_o2_n_spl_0,
    n616_lo_buf_o2_p_spl_
  );


  or

  (
    g634_n,
    n628_lo_buf_o2_p_spl_,
    n616_lo_buf_o2_n_spl_0
  );


  and

  (
    g635_p,
    g634_n,
    g633_n
  );


  or

  (
    g635_n,
    g634_p,
    g633_p
  );


  and

  (
    g636_p,
    n652_lo_buf_o2_p_spl_,
    n640_lo_buf_o2_n_spl_0
  );


  or

  (
    g636_n,
    n652_lo_buf_o2_n_spl_0,
    n640_lo_buf_o2_p_spl_
  );


  and

  (
    g637_p,
    n652_lo_buf_o2_n_spl_0,
    n640_lo_buf_o2_p_spl_
  );


  or

  (
    g637_n,
    n652_lo_buf_o2_p_spl_,
    n640_lo_buf_o2_n_spl_0
  );


  and

  (
    g638_p,
    g637_n,
    g636_n
  );


  or

  (
    g638_n,
    g637_p,
    g636_p
  );


  or

  (
    g639_n,
    g638_p,
    g635_n
  );


  or

  (
    g640_n,
    g638_n,
    g635_p
  );


  and

  (
    g641_p,
    g640_n,
    g639_n
  );


  not

  (
    G468,
    g237_p
  );


  not

  (
    G469,
    g241_p
  );


  not

  (
    G470,
    g245_p
  );


  not

  (
    G471,
    g249_p
  );


  not

  (
    G472,
    g257_p
  );


  not

  (
    G473,
    g261_p
  );


  not

  (
    G474,
    g265_p
  );


  not

  (
    G475,
    g269_p
  );


  not

  (
    G476,
    g277_p
  );


  not

  (
    G477,
    g281_p
  );


  not

  (
    G478,
    g285_p
  );


  not

  (
    G479,
    g289_p
  );


  not

  (
    G480,
    g297_p
  );


  not

  (
    G481,
    g301_p
  );


  not

  (
    G482,
    g305_p
  );


  not

  (
    G483,
    g309_p
  );


  not

  (
    G484,
    g317_p
  );


  not

  (
    G485,
    g321_p
  );


  not

  (
    G486,
    g325_p
  );


  not

  (
    G487,
    g329_p
  );


  not

  (
    G488,
    g337_p
  );


  not

  (
    G489,
    g341_p
  );


  not

  (
    G490,
    g345_p
  );


  not

  (
    G491,
    g349_p
  );


  not

  (
    G492,
    g357_p
  );


  not

  (
    G493,
    g361_p
  );


  not

  (
    G494,
    g365_p
  );


  not

  (
    G495,
    g369_p
  );


  not

  (
    G496,
    g377_p
  );


  not

  (
    G497,
    g381_p
  );


  not

  (
    G498,
    g385_p
  );


  not

  (
    G499,
    g389_p
  );


  not

  (
    n286_li,
    n1207_o2_n
  );


  not

  (
    n298_li,
    n1208_o2_n
  );


  not

  (
    n310_li,
    n1209_o2_n
  );


  not

  (
    n322_li,
    n1210_o2_n
  );


  not

  (
    n334_li,
    n1211_o2_n
  );


  not

  (
    n346_li,
    n1212_o2_n
  );


  not

  (
    n358_li,
    n1213_o2_n
  );


  not

  (
    n370_li,
    n1214_o2_n
  );


  not

  (
    n382_li,
    n1215_o2_n
  );


  not

  (
    n394_li,
    n1216_o2_n
  );


  not

  (
    n406_li,
    n1217_o2_n
  );


  not

  (
    n418_li,
    n1218_o2_n
  );


  not

  (
    n430_li,
    n1219_o2_n
  );


  not

  (
    n442_li,
    n1220_o2_n
  );


  not

  (
    n454_li,
    n1221_o2_n
  );


  not

  (
    n466_li,
    n1222_o2_n
  );


  not

  (
    n478_li,
    n1223_o2_n
  );


  not

  (
    n490_li,
    n1224_o2_n
  );


  not

  (
    n502_li,
    n1225_o2_n
  );


  not

  (
    n514_li,
    n1226_o2_n
  );


  not

  (
    n526_li,
    n1227_o2_n
  );


  not

  (
    n538_li,
    n1228_o2_n
  );


  not

  (
    n550_li,
    n1229_o2_n
  );


  not

  (
    n562_li,
    n1230_o2_n
  );


  not

  (
    n574_li,
    n1231_o2_n
  );


  not

  (
    n586_li,
    n1232_o2_n
  );


  not

  (
    n598_li,
    n1233_o2_n
  );


  not

  (
    n610_li,
    n1234_o2_n
  );


  not

  (
    n622_li,
    n1235_o2_n
  );


  not

  (
    n634_li,
    n1236_o2_n
  );


  not

  (
    n646_li,
    n1237_o2_n
  );


  not

  (
    n658_li,
    n1238_o2_n
  );


  not

  (
    n661_li,
    G33_n
  );


  not

  (
    n673_li,
    G34_n
  );


  not

  (
    n685_li,
    G35_n
  );


  not

  (
    n697_li,
    G36_n
  );


  not

  (
    n709_li,
    G37_n
  );


  not

  (
    n721_li,
    G38_n
  );


  not

  (
    n733_li,
    G39_n
  );


  not

  (
    n745_li,
    G40_n
  );


  not

  (
    n757_li,
    G41_n
  );


  not

  (
    n1248_i2,
    G234_o2_n_spl_0
  );


  not

  (
    n1249_i2,
    G247_o2_n_spl_0
  );


  not

  (
    n1250_i2,
    G260_o2_n_spl_0
  );


  not

  (
    n1251_i2,
    G273_o2_n_spl_0
  );


  not

  (
    n1252_i2,
    G286_o2_n_spl_0
  );


  not

  (
    n1253_i2,
    G299_o2_n_spl_0
  );


  not

  (
    n1254_i2,
    G312_o2_n_spl_0
  );


  not

  (
    n1255_i2,
    G325_o2_n_spl_0
  );


  not

  (
    n1207_i2,
    n283_lo_buf_o2_n_spl_
  );


  not

  (
    n1208_i2,
    n295_lo_buf_o2_n_spl_
  );


  not

  (
    n1209_i2,
    n307_lo_buf_o2_n_spl_
  );


  not

  (
    n1210_i2,
    n319_lo_buf_o2_n_spl_
  );


  not

  (
    n1211_i2,
    n331_lo_buf_o2_n_spl_
  );


  not

  (
    n1212_i2,
    n343_lo_buf_o2_n_spl_
  );


  not

  (
    n1213_i2,
    n355_lo_buf_o2_n_spl_
  );


  not

  (
    n1214_i2,
    n367_lo_buf_o2_n_spl_
  );


  not

  (
    n1215_i2,
    n379_lo_buf_o2_n_spl_
  );


  not

  (
    n1216_i2,
    n391_lo_buf_o2_n_spl_
  );


  not

  (
    n1217_i2,
    n403_lo_buf_o2_n_spl_
  );


  not

  (
    n1218_i2,
    n415_lo_buf_o2_n_spl_
  );


  not

  (
    n1219_i2,
    n427_lo_buf_o2_n_spl_
  );


  not

  (
    n1220_i2,
    n439_lo_buf_o2_n_spl_
  );


  not

  (
    n1221_i2,
    n451_lo_buf_o2_n_spl_
  );


  not

  (
    n1222_i2,
    n463_lo_buf_o2_n_spl_
  );


  not

  (
    n1223_i2,
    n475_lo_buf_o2_n_spl_
  );


  not

  (
    n1224_i2,
    n487_lo_buf_o2_n_spl_
  );


  not

  (
    n1225_i2,
    n499_lo_buf_o2_n_spl_
  );


  not

  (
    n1226_i2,
    n511_lo_buf_o2_n_spl_
  );


  not

  (
    n1227_i2,
    n523_lo_buf_o2_n_spl_
  );


  not

  (
    n1228_i2,
    n535_lo_buf_o2_n_spl_
  );


  not

  (
    n1229_i2,
    n547_lo_buf_o2_n_spl_
  );


  not

  (
    n1230_i2,
    n559_lo_buf_o2_n_spl_
  );


  not

  (
    n1231_i2,
    n571_lo_buf_o2_n_spl_
  );


  not

  (
    n1232_i2,
    n583_lo_buf_o2_n_spl_
  );


  not

  (
    n1233_i2,
    n595_lo_buf_o2_n_spl_
  );


  not

  (
    n1234_i2,
    n607_lo_buf_o2_n_spl_
  );


  not

  (
    n1235_i2,
    n619_lo_buf_o2_n_spl_
  );


  not

  (
    n1236_i2,
    n631_lo_buf_o2_n_spl_
  );


  not

  (
    n1237_i2,
    n643_lo_buf_o2_n_spl_
  );


  not

  (
    n1238_i2,
    n655_lo_buf_o2_n_spl_
  );


  not

  (
    G374_i2,
    G234_o2_n_spl_1
  );


  not

  (
    G376_i2,
    G234_o2_n_spl_1
  );


  not

  (
    G370_i2,
    G247_o2_n_spl_1
  );


  not

  (
    G372_i2,
    G247_o2_n_spl_1
  );


  not

  (
    G373_i2,
    G260_o2_n_spl_1
  );


  not

  (
    G377_i2,
    G260_o2_n_spl_1
  );


  not

  (
    G371_i2,
    G273_o2_n_spl_1
  );


  not

  (
    G375_i2,
    G273_o2_n_spl_1
  );


  not

  (
    G354_i2,
    G286_o2_n_spl_1
  );


  not

  (
    G356_i2,
    G286_o2_n_spl_1
  );


  not

  (
    G350_i2,
    G299_o2_n_spl_1
  );


  not

  (
    G352_i2,
    G299_o2_n_spl_1
  );


  not

  (
    G353_i2,
    G312_o2_n_spl_1
  );


  not

  (
    G357_i2,
    G312_o2_n_spl_1
  );


  not

  (
    G351_i2,
    G325_o2_n_spl_1
  );


  not

  (
    G355_i2,
    G325_o2_n_spl_1
  );


  not

  (
    G386_i2,
    g403_p
  );


  not

  (
    G391_i2,
    g417_p
  );


  not

  (
    n283_lo_buf_i2,
    n280_lo_buf_o2_n_spl_
  );


  not

  (
    n295_lo_buf_i2,
    n292_lo_buf_o2_n_spl_
  );


  not

  (
    n307_lo_buf_i2,
    n304_lo_buf_o2_n_spl_
  );


  not

  (
    n319_lo_buf_i2,
    n316_lo_buf_o2_n_spl_
  );


  not

  (
    n331_lo_buf_i2,
    n328_lo_buf_o2_n_spl_
  );


  not

  (
    n343_lo_buf_i2,
    n340_lo_buf_o2_n_spl_
  );


  not

  (
    n355_lo_buf_i2,
    n352_lo_buf_o2_n_spl_
  );


  not

  (
    n367_lo_buf_i2,
    n364_lo_buf_o2_n_spl_
  );


  not

  (
    n379_lo_buf_i2,
    n376_lo_buf_o2_n_spl_
  );


  not

  (
    n391_lo_buf_i2,
    n388_lo_buf_o2_n_spl_
  );


  not

  (
    n403_lo_buf_i2,
    n400_lo_buf_o2_n_spl_
  );


  not

  (
    n415_lo_buf_i2,
    n412_lo_buf_o2_n_spl_
  );


  not

  (
    n427_lo_buf_i2,
    n424_lo_buf_o2_n_spl_
  );


  not

  (
    n439_lo_buf_i2,
    n436_lo_buf_o2_n_spl_
  );


  not

  (
    n451_lo_buf_i2,
    n448_lo_buf_o2_n_spl_
  );


  not

  (
    n463_lo_buf_i2,
    n460_lo_buf_o2_n_spl_
  );


  not

  (
    n475_lo_buf_i2,
    n472_lo_buf_o2_n_spl_
  );


  not

  (
    n487_lo_buf_i2,
    n484_lo_buf_o2_n_spl_
  );


  not

  (
    n499_lo_buf_i2,
    n496_lo_buf_o2_n_spl_
  );


  not

  (
    n511_lo_buf_i2,
    n508_lo_buf_o2_n_spl_
  );


  not

  (
    n523_lo_buf_i2,
    n520_lo_buf_o2_n_spl_
  );


  not

  (
    n535_lo_buf_i2,
    n532_lo_buf_o2_n_spl_
  );


  not

  (
    n547_lo_buf_i2,
    n544_lo_buf_o2_n_spl_
  );


  not

  (
    n559_lo_buf_i2,
    n556_lo_buf_o2_n_spl_
  );


  not

  (
    n571_lo_buf_i2,
    n568_lo_buf_o2_n_spl_
  );


  not

  (
    n583_lo_buf_i2,
    n580_lo_buf_o2_n_spl_
  );


  not

  (
    n595_lo_buf_i2,
    n592_lo_buf_o2_n_spl_
  );


  not

  (
    n607_lo_buf_i2,
    n604_lo_buf_o2_n_spl_
  );


  not

  (
    n619_lo_buf_i2,
    n616_lo_buf_o2_n_spl_
  );


  not

  (
    n631_lo_buf_i2,
    n628_lo_buf_o2_n_spl_
  );


  not

  (
    n643_lo_buf_i2,
    n640_lo_buf_o2_n_spl_
  );


  not

  (
    n655_lo_buf_i2,
    n652_lo_buf_o2_n_spl_
  );


  not

  (
    G234_i2,
    g436_p
  );


  not

  (
    G247_i2,
    g455_p
  );


  not

  (
    G260_i2,
    g474_p
  );


  not

  (
    G273_i2,
    g493_p
  );


  not

  (
    G286_i2,
    g512_p
  );


  not

  (
    G299_i2,
    g531_p
  );


  not

  (
    G312_i2,
    g550_p
  );


  not

  (
    G325_i2,
    g569_p
  );


  not

  (
    n667_lo_buf_i2,
    n661_lo_n
  );


  not

  (
    n679_lo_buf_i2,
    n673_lo_n
  );


  not

  (
    n691_lo_buf_i2,
    n685_lo_n
  );


  not

  (
    n703_lo_buf_i2,
    n697_lo_n
  );


  not

  (
    n715_lo_buf_i2,
    n709_lo_n
  );


  not

  (
    n727_lo_buf_i2,
    n721_lo_n
  );


  not

  (
    n739_lo_buf_i2,
    n733_lo_n
  );


  not

  (
    n751_lo_buf_i2,
    n745_lo_n
  );


  not

  (
    n763_lo_buf_i2,
    n757_lo_n
  );


  not

  (
    G186_i2,
    g578_p
  );


  not

  (
    G189_i2,
    g587_p
  );


  not

  (
    G192_i2,
    g596_p
  );


  not

  (
    G195_i2,
    g605_p
  );


  not

  (
    G198_i2,
    g614_p
  );


  not

  (
    G201_i2,
    g623_p
  );


  not

  (
    G204_i2,
    g632_p
  );


  not

  (
    G207_i2,
    g641_p
  );


  not

  (
    n280_lo_buf_i2,
    G1_n
  );


  not

  (
    n292_lo_buf_i2,
    G2_n
  );


  not

  (
    n304_lo_buf_i2,
    G3_n
  );


  not

  (
    n316_lo_buf_i2,
    G4_n
  );


  not

  (
    n328_lo_buf_i2,
    G5_n
  );


  not

  (
    n340_lo_buf_i2,
    G6_n
  );


  not

  (
    n352_lo_buf_i2,
    G7_n
  );


  not

  (
    n364_lo_buf_i2,
    G8_n
  );


  not

  (
    n376_lo_buf_i2,
    G9_n
  );


  not

  (
    n388_lo_buf_i2,
    G10_n
  );


  not

  (
    n400_lo_buf_i2,
    G11_n
  );


  not

  (
    n412_lo_buf_i2,
    G12_n
  );


  not

  (
    n424_lo_buf_i2,
    G13_n
  );


  not

  (
    n436_lo_buf_i2,
    G14_n
  );


  not

  (
    n448_lo_buf_i2,
    G15_n
  );


  not

  (
    n460_lo_buf_i2,
    G16_n
  );


  not

  (
    n472_lo_buf_i2,
    G17_n
  );


  not

  (
    n484_lo_buf_i2,
    G18_n
  );


  not

  (
    n496_lo_buf_i2,
    G19_n
  );


  not

  (
    n508_lo_buf_i2,
    G20_n
  );


  not

  (
    n520_lo_buf_i2,
    G21_n
  );


  not

  (
    n532_lo_buf_i2,
    G22_n
  );


  not

  (
    n544_lo_buf_i2,
    G23_n
  );


  not

  (
    n556_lo_buf_i2,
    G24_n
  );


  not

  (
    n568_lo_buf_i2,
    G25_n
  );


  not

  (
    n580_lo_buf_i2,
    G26_n
  );


  not

  (
    n592_lo_buf_i2,
    G27_n
  );


  not

  (
    n604_lo_buf_i2,
    G28_n
  );


  not

  (
    n616_lo_buf_i2,
    G29_n
  );


  not

  (
    n628_lo_buf_i2,
    G30_n
  );


  not

  (
    n640_lo_buf_i2,
    G31_n
  );


  not

  (
    n652_lo_buf_i2,
    G32_n
  );


  buf

  (
    n1252_o2_p_spl_,
    n1252_o2_p
  );


  buf

  (
    n1252_o2_p_spl_0,
    n1252_o2_p_spl_
  );


  buf

  (
    n1252_o2_p_spl_00,
    n1252_o2_p_spl_0
  );


  buf

  (
    n1252_o2_p_spl_01,
    n1252_o2_p_spl_0
  );


  buf

  (
    n1252_o2_p_spl_1,
    n1252_o2_p_spl_
  );


  buf

  (
    n1252_o2_n_spl_,
    n1252_o2_n
  );


  buf

  (
    n1252_o2_n_spl_0,
    n1252_o2_n_spl_
  );


  buf

  (
    n1252_o2_n_spl_00,
    n1252_o2_n_spl_0
  );


  buf

  (
    n1252_o2_n_spl_01,
    n1252_o2_n_spl_0
  );


  buf

  (
    n1252_o2_n_spl_1,
    n1252_o2_n_spl_
  );


  buf

  (
    n1254_o2_p_spl_,
    n1254_o2_p
  );


  buf

  (
    n1254_o2_p_spl_0,
    n1254_o2_p_spl_
  );


  buf

  (
    n1254_o2_p_spl_00,
    n1254_o2_p_spl_0
  );


  buf

  (
    n1254_o2_p_spl_01,
    n1254_o2_p_spl_0
  );


  buf

  (
    n1254_o2_p_spl_1,
    n1254_o2_p_spl_
  );


  buf

  (
    n1254_o2_n_spl_,
    n1254_o2_n
  );


  buf

  (
    n1254_o2_n_spl_0,
    n1254_o2_n_spl_
  );


  buf

  (
    n1254_o2_n_spl_00,
    n1254_o2_n_spl_0
  );


  buf

  (
    n1254_o2_n_spl_01,
    n1254_o2_n_spl_0
  );


  buf

  (
    n1254_o2_n_spl_1,
    n1254_o2_n_spl_
  );


  buf

  (
    G386_o2_p_spl_,
    G386_o2_p
  );


  buf

  (
    G386_o2_p_spl_0,
    G386_o2_p_spl_
  );


  buf

  (
    G386_o2_p_spl_1,
    G386_o2_p_spl_
  );


  buf

  (
    G386_o2_n_spl_,
    G386_o2_n
  );


  buf

  (
    G386_o2_n_spl_0,
    G386_o2_n_spl_
  );


  buf

  (
    G386_o2_n_spl_1,
    G386_o2_n_spl_
  );


  buf

  (
    g233_p_spl_,
    g233_p
  );


  buf

  (
    g233_p_spl_0,
    g233_p_spl_
  );


  buf

  (
    g233_p_spl_1,
    g233_p_spl_
  );


  buf

  (
    n1248_o2_p_spl_,
    n1248_o2_p
  );


  buf

  (
    n1248_o2_p_spl_0,
    n1248_o2_p_spl_
  );


  buf

  (
    n1248_o2_p_spl_00,
    n1248_o2_p_spl_0
  );


  buf

  (
    n1248_o2_p_spl_01,
    n1248_o2_p_spl_0
  );


  buf

  (
    n1248_o2_p_spl_1,
    n1248_o2_p_spl_
  );


  buf

  (
    g233_n_spl_,
    g233_n
  );


  buf

  (
    g233_n_spl_0,
    g233_n_spl_
  );


  buf

  (
    g233_n_spl_1,
    g233_n_spl_
  );


  buf

  (
    n1248_o2_n_spl_,
    n1248_o2_n
  );


  buf

  (
    n1248_o2_n_spl_0,
    n1248_o2_n_spl_
  );


  buf

  (
    n1248_o2_n_spl_00,
    n1248_o2_n_spl_0
  );


  buf

  (
    n1248_o2_n_spl_01,
    n1248_o2_n_spl_0
  );


  buf

  (
    n1248_o2_n_spl_1,
    n1248_o2_n_spl_
  );


  buf

  (
    n1249_o2_p_spl_,
    n1249_o2_p
  );


  buf

  (
    n1249_o2_p_spl_0,
    n1249_o2_p_spl_
  );


  buf

  (
    n1249_o2_p_spl_00,
    n1249_o2_p_spl_0
  );


  buf

  (
    n1249_o2_p_spl_01,
    n1249_o2_p_spl_0
  );


  buf

  (
    n1249_o2_p_spl_1,
    n1249_o2_p_spl_
  );


  buf

  (
    n1249_o2_n_spl_,
    n1249_o2_n
  );


  buf

  (
    n1249_o2_n_spl_0,
    n1249_o2_n_spl_
  );


  buf

  (
    n1249_o2_n_spl_00,
    n1249_o2_n_spl_0
  );


  buf

  (
    n1249_o2_n_spl_01,
    n1249_o2_n_spl_0
  );


  buf

  (
    n1249_o2_n_spl_1,
    n1249_o2_n_spl_
  );


  buf

  (
    n1250_o2_p_spl_,
    n1250_o2_p
  );


  buf

  (
    n1250_o2_p_spl_0,
    n1250_o2_p_spl_
  );


  buf

  (
    n1250_o2_p_spl_00,
    n1250_o2_p_spl_0
  );


  buf

  (
    n1250_o2_p_spl_01,
    n1250_o2_p_spl_0
  );


  buf

  (
    n1250_o2_p_spl_1,
    n1250_o2_p_spl_
  );


  buf

  (
    n1250_o2_n_spl_,
    n1250_o2_n
  );


  buf

  (
    n1250_o2_n_spl_0,
    n1250_o2_n_spl_
  );


  buf

  (
    n1250_o2_n_spl_00,
    n1250_o2_n_spl_0
  );


  buf

  (
    n1250_o2_n_spl_01,
    n1250_o2_n_spl_0
  );


  buf

  (
    n1250_o2_n_spl_1,
    n1250_o2_n_spl_
  );


  buf

  (
    n1251_o2_p_spl_,
    n1251_o2_p
  );


  buf

  (
    n1251_o2_p_spl_0,
    n1251_o2_p_spl_
  );


  buf

  (
    n1251_o2_p_spl_00,
    n1251_o2_p_spl_0
  );


  buf

  (
    n1251_o2_p_spl_01,
    n1251_o2_p_spl_0
  );


  buf

  (
    n1251_o2_p_spl_1,
    n1251_o2_p_spl_
  );


  buf

  (
    n1251_o2_n_spl_,
    n1251_o2_n
  );


  buf

  (
    n1251_o2_n_spl_0,
    n1251_o2_n_spl_
  );


  buf

  (
    n1251_o2_n_spl_00,
    n1251_o2_n_spl_0
  );


  buf

  (
    n1251_o2_n_spl_01,
    n1251_o2_n_spl_0
  );


  buf

  (
    n1251_o2_n_spl_1,
    n1251_o2_n_spl_
  );


  buf

  (
    n1255_o2_p_spl_,
    n1255_o2_p
  );


  buf

  (
    n1255_o2_p_spl_0,
    n1255_o2_p_spl_
  );


  buf

  (
    n1255_o2_p_spl_00,
    n1255_o2_p_spl_0
  );


  buf

  (
    n1255_o2_p_spl_01,
    n1255_o2_p_spl_0
  );


  buf

  (
    n1255_o2_p_spl_1,
    n1255_o2_p_spl_
  );


  buf

  (
    n1255_o2_n_spl_,
    n1255_o2_n
  );


  buf

  (
    n1255_o2_n_spl_0,
    n1255_o2_n_spl_
  );


  buf

  (
    n1255_o2_n_spl_00,
    n1255_o2_n_spl_0
  );


  buf

  (
    n1255_o2_n_spl_01,
    n1255_o2_n_spl_0
  );


  buf

  (
    n1255_o2_n_spl_1,
    n1255_o2_n_spl_
  );


  buf

  (
    g253_p_spl_,
    g253_p
  );


  buf

  (
    g253_p_spl_0,
    g253_p_spl_
  );


  buf

  (
    g253_p_spl_1,
    g253_p_spl_
  );


  buf

  (
    g253_n_spl_,
    g253_n
  );


  buf

  (
    g253_n_spl_0,
    g253_n_spl_
  );


  buf

  (
    g253_n_spl_1,
    g253_n_spl_
  );


  buf

  (
    n1253_o2_p_spl_,
    n1253_o2_p
  );


  buf

  (
    n1253_o2_p_spl_0,
    n1253_o2_p_spl_
  );


  buf

  (
    n1253_o2_p_spl_00,
    n1253_o2_p_spl_0
  );


  buf

  (
    n1253_o2_p_spl_01,
    n1253_o2_p_spl_0
  );


  buf

  (
    n1253_o2_p_spl_1,
    n1253_o2_p_spl_
  );


  buf

  (
    n1253_o2_n_spl_,
    n1253_o2_n
  );


  buf

  (
    n1253_o2_n_spl_0,
    n1253_o2_n_spl_
  );


  buf

  (
    n1253_o2_n_spl_00,
    n1253_o2_n_spl_0
  );


  buf

  (
    n1253_o2_n_spl_01,
    n1253_o2_n_spl_0
  );


  buf

  (
    n1253_o2_n_spl_1,
    n1253_o2_n_spl_
  );


  buf

  (
    g273_p_spl_,
    g273_p
  );


  buf

  (
    g273_p_spl_0,
    g273_p_spl_
  );


  buf

  (
    g273_p_spl_1,
    g273_p_spl_
  );


  buf

  (
    g273_n_spl_,
    g273_n
  );


  buf

  (
    g273_n_spl_0,
    g273_n_spl_
  );


  buf

  (
    g273_n_spl_1,
    g273_n_spl_
  );


  buf

  (
    g293_p_spl_,
    g293_p
  );


  buf

  (
    g293_p_spl_0,
    g293_p_spl_
  );


  buf

  (
    g293_p_spl_1,
    g293_p_spl_
  );


  buf

  (
    g293_n_spl_,
    g293_n
  );


  buf

  (
    g293_n_spl_0,
    g293_n_spl_
  );


  buf

  (
    g293_n_spl_1,
    g293_n_spl_
  );


  buf

  (
    G391_o2_p_spl_,
    G391_o2_p
  );


  buf

  (
    G391_o2_p_spl_0,
    G391_o2_p_spl_
  );


  buf

  (
    G391_o2_p_spl_1,
    G391_o2_p_spl_
  );


  buf

  (
    G391_o2_n_spl_,
    G391_o2_n
  );


  buf

  (
    G391_o2_n_spl_0,
    G391_o2_n_spl_
  );


  buf

  (
    G391_o2_n_spl_1,
    G391_o2_n_spl_
  );


  buf

  (
    g313_p_spl_,
    g313_p
  );


  buf

  (
    g313_p_spl_0,
    g313_p_spl_
  );


  buf

  (
    g313_p_spl_1,
    g313_p_spl_
  );


  buf

  (
    g313_n_spl_,
    g313_n
  );


  buf

  (
    g313_n_spl_0,
    g313_n_spl_
  );


  buf

  (
    g313_n_spl_1,
    g313_n_spl_
  );


  buf

  (
    g333_p_spl_,
    g333_p
  );


  buf

  (
    g333_p_spl_0,
    g333_p_spl_
  );


  buf

  (
    g333_p_spl_1,
    g333_p_spl_
  );


  buf

  (
    g333_n_spl_,
    g333_n
  );


  buf

  (
    g333_n_spl_0,
    g333_n_spl_
  );


  buf

  (
    g333_n_spl_1,
    g333_n_spl_
  );


  buf

  (
    g353_p_spl_,
    g353_p
  );


  buf

  (
    g353_p_spl_0,
    g353_p_spl_
  );


  buf

  (
    g353_p_spl_1,
    g353_p_spl_
  );


  buf

  (
    g353_n_spl_,
    g353_n
  );


  buf

  (
    g353_n_spl_0,
    g353_n_spl_
  );


  buf

  (
    g353_n_spl_1,
    g353_n_spl_
  );


  buf

  (
    g373_p_spl_,
    g373_p
  );


  buf

  (
    g373_p_spl_0,
    g373_p_spl_
  );


  buf

  (
    g373_p_spl_1,
    g373_p_spl_
  );


  buf

  (
    g373_n_spl_,
    g373_n
  );


  buf

  (
    g373_n_spl_0,
    g373_n_spl_
  );


  buf

  (
    g373_n_spl_1,
    g373_n_spl_
  );


  buf

  (
    G247_o2_p_spl_,
    G247_o2_p
  );


  buf

  (
    G234_o2_p_spl_,
    G234_o2_p
  );


  buf

  (
    g390_n_spl_,
    g390_n
  );


  buf

  (
    G260_o2_p_spl_,
    G260_o2_p
  );


  buf

  (
    G260_o2_p_spl_0,
    G260_o2_p_spl_
  );


  buf

  (
    G273_o2_n_spl_,
    G273_o2_n
  );


  buf

  (
    G273_o2_n_spl_0,
    G273_o2_n_spl_
  );


  buf

  (
    G273_o2_n_spl_1,
    G273_o2_n_spl_
  );


  buf

  (
    G260_o2_n_spl_,
    G260_o2_n
  );


  buf

  (
    G260_o2_n_spl_0,
    G260_o2_n_spl_
  );


  buf

  (
    G260_o2_n_spl_1,
    G260_o2_n_spl_
  );


  buf

  (
    G273_o2_p_spl_,
    G273_o2_p
  );


  buf

  (
    G273_o2_p_spl_0,
    G273_o2_p_spl_
  );


  buf

  (
    G247_o2_n_spl_,
    G247_o2_n
  );


  buf

  (
    G247_o2_n_spl_0,
    G247_o2_n_spl_
  );


  buf

  (
    G247_o2_n_spl_1,
    G247_o2_n_spl_
  );


  buf

  (
    G234_o2_n_spl_,
    G234_o2_n
  );


  buf

  (
    G234_o2_n_spl_0,
    G234_o2_n_spl_
  );


  buf

  (
    G234_o2_n_spl_1,
    G234_o2_n_spl_
  );


  buf

  (
    G299_o2_p_spl_,
    G299_o2_p
  );


  buf

  (
    G286_o2_p_spl_,
    G286_o2_p
  );


  buf

  (
    g404_n_spl_,
    g404_n
  );


  buf

  (
    G312_o2_p_spl_,
    G312_o2_p
  );


  buf

  (
    G312_o2_p_spl_0,
    G312_o2_p_spl_
  );


  buf

  (
    G325_o2_n_spl_,
    G325_o2_n
  );


  buf

  (
    G325_o2_n_spl_0,
    G325_o2_n_spl_
  );


  buf

  (
    G325_o2_n_spl_1,
    G325_o2_n_spl_
  );


  buf

  (
    G312_o2_n_spl_,
    G312_o2_n
  );


  buf

  (
    G312_o2_n_spl_0,
    G312_o2_n_spl_
  );


  buf

  (
    G312_o2_n_spl_1,
    G312_o2_n_spl_
  );


  buf

  (
    G325_o2_p_spl_,
    G325_o2_p
  );


  buf

  (
    G325_o2_p_spl_0,
    G325_o2_p_spl_
  );


  buf

  (
    G299_o2_n_spl_,
    G299_o2_n
  );


  buf

  (
    G299_o2_n_spl_0,
    G299_o2_n_spl_
  );


  buf

  (
    G299_o2_n_spl_1,
    G299_o2_n_spl_
  );


  buf

  (
    G286_o2_n_spl_,
    G286_o2_n
  );


  buf

  (
    G286_o2_n_spl_0,
    G286_o2_n_spl_
  );


  buf

  (
    G286_o2_n_spl_1,
    G286_o2_n_spl_
  );


  buf

  (
    n331_lo_buf_o2_p_spl_,
    n331_lo_buf_o2_p
  );


  buf

  (
    n283_lo_buf_o2_n_spl_,
    n283_lo_buf_o2_n
  );


  buf

  (
    n283_lo_buf_o2_n_spl_0,
    n283_lo_buf_o2_n_spl_
  );


  buf

  (
    n331_lo_buf_o2_n_spl_,
    n331_lo_buf_o2_n
  );


  buf

  (
    n331_lo_buf_o2_n_spl_0,
    n331_lo_buf_o2_n_spl_
  );


  buf

  (
    n283_lo_buf_o2_p_spl_,
    n283_lo_buf_o2_p
  );


  buf

  (
    n427_lo_buf_o2_p_spl_,
    n427_lo_buf_o2_p
  );


  buf

  (
    n379_lo_buf_o2_n_spl_,
    n379_lo_buf_o2_n
  );


  buf

  (
    n379_lo_buf_o2_n_spl_0,
    n379_lo_buf_o2_n_spl_
  );


  buf

  (
    n427_lo_buf_o2_n_spl_,
    n427_lo_buf_o2_n
  );


  buf

  (
    n427_lo_buf_o2_n_spl_0,
    n427_lo_buf_o2_n_spl_
  );


  buf

  (
    n379_lo_buf_o2_p_spl_,
    n379_lo_buf_o2_p
  );


  buf

  (
    g423_n_spl_,
    g423_n
  );


  buf

  (
    g420_p_spl_,
    g420_p
  );


  buf

  (
    g423_p_spl_,
    g423_p
  );


  buf

  (
    g420_n_spl_,
    g420_n
  );


  buf

  (
    n763_lo_buf_o2_p_spl_,
    n763_lo_buf_o2_p
  );


  buf

  (
    n763_lo_buf_o2_p_spl_0,
    n763_lo_buf_o2_p_spl_
  );


  buf

  (
    n763_lo_buf_o2_p_spl_00,
    n763_lo_buf_o2_p_spl_0
  );


  buf

  (
    n763_lo_buf_o2_p_spl_01,
    n763_lo_buf_o2_p_spl_0
  );


  buf

  (
    n763_lo_buf_o2_p_spl_1,
    n763_lo_buf_o2_p_spl_
  );


  buf

  (
    n763_lo_buf_o2_p_spl_10,
    n763_lo_buf_o2_p_spl_1
  );


  buf

  (
    n763_lo_buf_o2_p_spl_11,
    n763_lo_buf_o2_p_spl_1
  );


  buf

  (
    n763_lo_buf_o2_n_spl_,
    n763_lo_buf_o2_n
  );


  buf

  (
    n763_lo_buf_o2_n_spl_0,
    n763_lo_buf_o2_n_spl_
  );


  buf

  (
    n763_lo_buf_o2_n_spl_00,
    n763_lo_buf_o2_n_spl_0
  );


  buf

  (
    n763_lo_buf_o2_n_spl_01,
    n763_lo_buf_o2_n_spl_0
  );


  buf

  (
    n763_lo_buf_o2_n_spl_1,
    n763_lo_buf_o2_n_spl_
  );


  buf

  (
    n763_lo_buf_o2_n_spl_10,
    n763_lo_buf_o2_n_spl_1
  );


  buf

  (
    n763_lo_buf_o2_n_spl_11,
    n763_lo_buf_o2_n_spl_1
  );


  buf

  (
    G201_o2_p_spl_,
    G201_o2_p
  );


  buf

  (
    G201_o2_p_spl_0,
    G201_o2_p_spl_
  );


  buf

  (
    G201_o2_p_spl_1,
    G201_o2_p_spl_
  );


  buf

  (
    G198_o2_n_spl_,
    G198_o2_n
  );


  buf

  (
    G198_o2_n_spl_0,
    G198_o2_n_spl_
  );


  buf

  (
    G198_o2_n_spl_1,
    G198_o2_n_spl_
  );


  buf

  (
    G201_o2_n_spl_,
    G201_o2_n
  );


  buf

  (
    G201_o2_n_spl_0,
    G201_o2_n_spl_
  );


  buf

  (
    G201_o2_n_spl_1,
    G201_o2_n_spl_
  );


  buf

  (
    G198_o2_p_spl_,
    G198_o2_p
  );


  buf

  (
    G198_o2_p_spl_0,
    G198_o2_p_spl_
  );


  buf

  (
    G198_o2_p_spl_1,
    G198_o2_p_spl_
  );


  buf

  (
    g430_n_spl_,
    g430_n
  );


  buf

  (
    g427_n_spl_,
    g427_n
  );


  buf

  (
    g430_p_spl_,
    g430_p
  );


  buf

  (
    g427_p_spl_,
    g427_p
  );


  buf

  (
    n343_lo_buf_o2_p_spl_,
    n343_lo_buf_o2_p
  );


  buf

  (
    n295_lo_buf_o2_n_spl_,
    n295_lo_buf_o2_n
  );


  buf

  (
    n295_lo_buf_o2_n_spl_0,
    n295_lo_buf_o2_n_spl_
  );


  buf

  (
    n343_lo_buf_o2_n_spl_,
    n343_lo_buf_o2_n
  );


  buf

  (
    n343_lo_buf_o2_n_spl_0,
    n343_lo_buf_o2_n_spl_
  );


  buf

  (
    n295_lo_buf_o2_p_spl_,
    n295_lo_buf_o2_p
  );


  buf

  (
    n439_lo_buf_o2_p_spl_,
    n439_lo_buf_o2_p
  );


  buf

  (
    n391_lo_buf_o2_n_spl_,
    n391_lo_buf_o2_n
  );


  buf

  (
    n391_lo_buf_o2_n_spl_0,
    n391_lo_buf_o2_n_spl_
  );


  buf

  (
    n439_lo_buf_o2_n_spl_,
    n439_lo_buf_o2_n
  );


  buf

  (
    n439_lo_buf_o2_n_spl_0,
    n439_lo_buf_o2_n_spl_
  );


  buf

  (
    n391_lo_buf_o2_p_spl_,
    n391_lo_buf_o2_p
  );


  buf

  (
    g442_n_spl_,
    g442_n
  );


  buf

  (
    g439_p_spl_,
    g439_p
  );


  buf

  (
    g442_p_spl_,
    g442_p
  );


  buf

  (
    g439_n_spl_,
    g439_n
  );


  buf

  (
    G207_o2_p_spl_,
    G207_o2_p
  );


  buf

  (
    G207_o2_p_spl_0,
    G207_o2_p_spl_
  );


  buf

  (
    G207_o2_p_spl_1,
    G207_o2_p_spl_
  );


  buf

  (
    G204_o2_n_spl_,
    G204_o2_n
  );


  buf

  (
    G204_o2_n_spl_0,
    G204_o2_n_spl_
  );


  buf

  (
    G204_o2_n_spl_1,
    G204_o2_n_spl_
  );


  buf

  (
    G207_o2_n_spl_,
    G207_o2_n
  );


  buf

  (
    G207_o2_n_spl_0,
    G207_o2_n_spl_
  );


  buf

  (
    G207_o2_n_spl_1,
    G207_o2_n_spl_
  );


  buf

  (
    G204_o2_p_spl_,
    G204_o2_p
  );


  buf

  (
    G204_o2_p_spl_0,
    G204_o2_p_spl_
  );


  buf

  (
    G204_o2_p_spl_1,
    G204_o2_p_spl_
  );


  buf

  (
    g449_n_spl_,
    g449_n
  );


  buf

  (
    g446_n_spl_,
    g446_n
  );


  buf

  (
    g449_p_spl_,
    g449_p
  );


  buf

  (
    g446_p_spl_,
    g446_p
  );


  buf

  (
    n355_lo_buf_o2_p_spl_,
    n355_lo_buf_o2_p
  );


  buf

  (
    n307_lo_buf_o2_n_spl_,
    n307_lo_buf_o2_n
  );


  buf

  (
    n307_lo_buf_o2_n_spl_0,
    n307_lo_buf_o2_n_spl_
  );


  buf

  (
    n355_lo_buf_o2_n_spl_,
    n355_lo_buf_o2_n
  );


  buf

  (
    n355_lo_buf_o2_n_spl_0,
    n355_lo_buf_o2_n_spl_
  );


  buf

  (
    n307_lo_buf_o2_p_spl_,
    n307_lo_buf_o2_p
  );


  buf

  (
    n451_lo_buf_o2_p_spl_,
    n451_lo_buf_o2_p
  );


  buf

  (
    n403_lo_buf_o2_n_spl_,
    n403_lo_buf_o2_n
  );


  buf

  (
    n403_lo_buf_o2_n_spl_0,
    n403_lo_buf_o2_n_spl_
  );


  buf

  (
    n451_lo_buf_o2_n_spl_,
    n451_lo_buf_o2_n
  );


  buf

  (
    n451_lo_buf_o2_n_spl_0,
    n451_lo_buf_o2_n_spl_
  );


  buf

  (
    n403_lo_buf_o2_p_spl_,
    n403_lo_buf_o2_p
  );


  buf

  (
    g461_n_spl_,
    g461_n
  );


  buf

  (
    g458_p_spl_,
    g458_p
  );


  buf

  (
    g461_p_spl_,
    g461_p
  );


  buf

  (
    g458_n_spl_,
    g458_n
  );


  buf

  (
    g468_n_spl_,
    g468_n
  );


  buf

  (
    g465_n_spl_,
    g465_n
  );


  buf

  (
    g468_p_spl_,
    g468_p
  );


  buf

  (
    g465_p_spl_,
    g465_p
  );


  buf

  (
    n367_lo_buf_o2_p_spl_,
    n367_lo_buf_o2_p
  );


  buf

  (
    n319_lo_buf_o2_n_spl_,
    n319_lo_buf_o2_n
  );


  buf

  (
    n319_lo_buf_o2_n_spl_0,
    n319_lo_buf_o2_n_spl_
  );


  buf

  (
    n367_lo_buf_o2_n_spl_,
    n367_lo_buf_o2_n
  );


  buf

  (
    n367_lo_buf_o2_n_spl_0,
    n367_lo_buf_o2_n_spl_
  );


  buf

  (
    n319_lo_buf_o2_p_spl_,
    n319_lo_buf_o2_p
  );


  buf

  (
    n463_lo_buf_o2_p_spl_,
    n463_lo_buf_o2_p
  );


  buf

  (
    n415_lo_buf_o2_n_spl_,
    n415_lo_buf_o2_n
  );


  buf

  (
    n415_lo_buf_o2_n_spl_0,
    n415_lo_buf_o2_n_spl_
  );


  buf

  (
    n463_lo_buf_o2_n_spl_,
    n463_lo_buf_o2_n
  );


  buf

  (
    n463_lo_buf_o2_n_spl_0,
    n463_lo_buf_o2_n_spl_
  );


  buf

  (
    n415_lo_buf_o2_p_spl_,
    n415_lo_buf_o2_p
  );


  buf

  (
    g480_n_spl_,
    g480_n
  );


  buf

  (
    g477_p_spl_,
    g477_p
  );


  buf

  (
    g480_p_spl_,
    g480_p
  );


  buf

  (
    g477_n_spl_,
    g477_n
  );


  buf

  (
    g487_n_spl_,
    g487_n
  );


  buf

  (
    g484_n_spl_,
    g484_n
  );


  buf

  (
    g487_p_spl_,
    g487_p
  );


  buf

  (
    g484_p_spl_,
    g484_p
  );


  buf

  (
    n523_lo_buf_o2_p_spl_,
    n523_lo_buf_o2_p
  );


  buf

  (
    n475_lo_buf_o2_n_spl_,
    n475_lo_buf_o2_n
  );


  buf

  (
    n475_lo_buf_o2_n_spl_0,
    n475_lo_buf_o2_n_spl_
  );


  buf

  (
    n523_lo_buf_o2_n_spl_,
    n523_lo_buf_o2_n
  );


  buf

  (
    n523_lo_buf_o2_n_spl_0,
    n523_lo_buf_o2_n_spl_
  );


  buf

  (
    n475_lo_buf_o2_p_spl_,
    n475_lo_buf_o2_p
  );


  buf

  (
    n619_lo_buf_o2_p_spl_,
    n619_lo_buf_o2_p
  );


  buf

  (
    n571_lo_buf_o2_n_spl_,
    n571_lo_buf_o2_n
  );


  buf

  (
    n571_lo_buf_o2_n_spl_0,
    n571_lo_buf_o2_n_spl_
  );


  buf

  (
    n619_lo_buf_o2_n_spl_,
    n619_lo_buf_o2_n
  );


  buf

  (
    n619_lo_buf_o2_n_spl_0,
    n619_lo_buf_o2_n_spl_
  );


  buf

  (
    n571_lo_buf_o2_p_spl_,
    n571_lo_buf_o2_p
  );


  buf

  (
    g499_n_spl_,
    g499_n
  );


  buf

  (
    g496_p_spl_,
    g496_p
  );


  buf

  (
    g499_p_spl_,
    g499_p
  );


  buf

  (
    g496_n_spl_,
    g496_n
  );


  buf

  (
    G189_o2_p_spl_,
    G189_o2_p
  );


  buf

  (
    G189_o2_p_spl_0,
    G189_o2_p_spl_
  );


  buf

  (
    G189_o2_p_spl_1,
    G189_o2_p_spl_
  );


  buf

  (
    G186_o2_n_spl_,
    G186_o2_n
  );


  buf

  (
    G186_o2_n_spl_0,
    G186_o2_n_spl_
  );


  buf

  (
    G186_o2_n_spl_1,
    G186_o2_n_spl_
  );


  buf

  (
    G189_o2_n_spl_,
    G189_o2_n
  );


  buf

  (
    G189_o2_n_spl_0,
    G189_o2_n_spl_
  );


  buf

  (
    G189_o2_n_spl_1,
    G189_o2_n_spl_
  );


  buf

  (
    G186_o2_p_spl_,
    G186_o2_p
  );


  buf

  (
    G186_o2_p_spl_0,
    G186_o2_p_spl_
  );


  buf

  (
    G186_o2_p_spl_1,
    G186_o2_p_spl_
  );


  buf

  (
    g506_n_spl_,
    g506_n
  );


  buf

  (
    g503_n_spl_,
    g503_n
  );


  buf

  (
    g506_p_spl_,
    g506_p
  );


  buf

  (
    g503_p_spl_,
    g503_p
  );


  buf

  (
    n535_lo_buf_o2_p_spl_,
    n535_lo_buf_o2_p
  );


  buf

  (
    n487_lo_buf_o2_n_spl_,
    n487_lo_buf_o2_n
  );


  buf

  (
    n487_lo_buf_o2_n_spl_0,
    n487_lo_buf_o2_n_spl_
  );


  buf

  (
    n535_lo_buf_o2_n_spl_,
    n535_lo_buf_o2_n
  );


  buf

  (
    n535_lo_buf_o2_n_spl_0,
    n535_lo_buf_o2_n_spl_
  );


  buf

  (
    n487_lo_buf_o2_p_spl_,
    n487_lo_buf_o2_p
  );


  buf

  (
    n631_lo_buf_o2_p_spl_,
    n631_lo_buf_o2_p
  );


  buf

  (
    n583_lo_buf_o2_n_spl_,
    n583_lo_buf_o2_n
  );


  buf

  (
    n583_lo_buf_o2_n_spl_0,
    n583_lo_buf_o2_n_spl_
  );


  buf

  (
    n631_lo_buf_o2_n_spl_,
    n631_lo_buf_o2_n
  );


  buf

  (
    n631_lo_buf_o2_n_spl_0,
    n631_lo_buf_o2_n_spl_
  );


  buf

  (
    n583_lo_buf_o2_p_spl_,
    n583_lo_buf_o2_p
  );


  buf

  (
    g518_n_spl_,
    g518_n
  );


  buf

  (
    g515_p_spl_,
    g515_p
  );


  buf

  (
    g518_p_spl_,
    g518_p
  );


  buf

  (
    g515_n_spl_,
    g515_n
  );


  buf

  (
    G195_o2_p_spl_,
    G195_o2_p
  );


  buf

  (
    G195_o2_p_spl_0,
    G195_o2_p_spl_
  );


  buf

  (
    G195_o2_p_spl_1,
    G195_o2_p_spl_
  );


  buf

  (
    G192_o2_n_spl_,
    G192_o2_n
  );


  buf

  (
    G192_o2_n_spl_0,
    G192_o2_n_spl_
  );


  buf

  (
    G192_o2_n_spl_1,
    G192_o2_n_spl_
  );


  buf

  (
    G195_o2_n_spl_,
    G195_o2_n
  );


  buf

  (
    G195_o2_n_spl_0,
    G195_o2_n_spl_
  );


  buf

  (
    G195_o2_n_spl_1,
    G195_o2_n_spl_
  );


  buf

  (
    G192_o2_p_spl_,
    G192_o2_p
  );


  buf

  (
    G192_o2_p_spl_0,
    G192_o2_p_spl_
  );


  buf

  (
    G192_o2_p_spl_1,
    G192_o2_p_spl_
  );


  buf

  (
    g525_n_spl_,
    g525_n
  );


  buf

  (
    g522_n_spl_,
    g522_n
  );


  buf

  (
    g525_p_spl_,
    g525_p
  );


  buf

  (
    g522_p_spl_,
    g522_p
  );


  buf

  (
    n547_lo_buf_o2_p_spl_,
    n547_lo_buf_o2_p
  );


  buf

  (
    n499_lo_buf_o2_n_spl_,
    n499_lo_buf_o2_n
  );


  buf

  (
    n499_lo_buf_o2_n_spl_0,
    n499_lo_buf_o2_n_spl_
  );


  buf

  (
    n547_lo_buf_o2_n_spl_,
    n547_lo_buf_o2_n
  );


  buf

  (
    n547_lo_buf_o2_n_spl_0,
    n547_lo_buf_o2_n_spl_
  );


  buf

  (
    n499_lo_buf_o2_p_spl_,
    n499_lo_buf_o2_p
  );


  buf

  (
    n643_lo_buf_o2_p_spl_,
    n643_lo_buf_o2_p
  );


  buf

  (
    n595_lo_buf_o2_n_spl_,
    n595_lo_buf_o2_n
  );


  buf

  (
    n595_lo_buf_o2_n_spl_0,
    n595_lo_buf_o2_n_spl_
  );


  buf

  (
    n643_lo_buf_o2_n_spl_,
    n643_lo_buf_o2_n
  );


  buf

  (
    n643_lo_buf_o2_n_spl_0,
    n643_lo_buf_o2_n_spl_
  );


  buf

  (
    n595_lo_buf_o2_p_spl_,
    n595_lo_buf_o2_p
  );


  buf

  (
    g537_n_spl_,
    g537_n
  );


  buf

  (
    g534_p_spl_,
    g534_p
  );


  buf

  (
    g537_p_spl_,
    g537_p
  );


  buf

  (
    g534_n_spl_,
    g534_n
  );


  buf

  (
    g544_n_spl_,
    g544_n
  );


  buf

  (
    g541_n_spl_,
    g541_n
  );


  buf

  (
    g544_p_spl_,
    g544_p
  );


  buf

  (
    g541_p_spl_,
    g541_p
  );


  buf

  (
    n559_lo_buf_o2_p_spl_,
    n559_lo_buf_o2_p
  );


  buf

  (
    n511_lo_buf_o2_n_spl_,
    n511_lo_buf_o2_n
  );


  buf

  (
    n511_lo_buf_o2_n_spl_0,
    n511_lo_buf_o2_n_spl_
  );


  buf

  (
    n559_lo_buf_o2_n_spl_,
    n559_lo_buf_o2_n
  );


  buf

  (
    n559_lo_buf_o2_n_spl_0,
    n559_lo_buf_o2_n_spl_
  );


  buf

  (
    n511_lo_buf_o2_p_spl_,
    n511_lo_buf_o2_p
  );


  buf

  (
    n655_lo_buf_o2_p_spl_,
    n655_lo_buf_o2_p
  );


  buf

  (
    n607_lo_buf_o2_n_spl_,
    n607_lo_buf_o2_n
  );


  buf

  (
    n607_lo_buf_o2_n_spl_0,
    n607_lo_buf_o2_n_spl_
  );


  buf

  (
    n655_lo_buf_o2_n_spl_,
    n655_lo_buf_o2_n
  );


  buf

  (
    n655_lo_buf_o2_n_spl_0,
    n655_lo_buf_o2_n_spl_
  );


  buf

  (
    n607_lo_buf_o2_p_spl_,
    n607_lo_buf_o2_p
  );


  buf

  (
    g556_n_spl_,
    g556_n
  );


  buf

  (
    g553_p_spl_,
    g553_p
  );


  buf

  (
    g556_p_spl_,
    g556_p
  );


  buf

  (
    g553_n_spl_,
    g553_n
  );


  buf

  (
    g563_n_spl_,
    g563_n
  );


  buf

  (
    g560_n_spl_,
    g560_n
  );


  buf

  (
    g563_p_spl_,
    g563_p
  );


  buf

  (
    g560_p_spl_,
    g560_p
  );


  buf

  (
    n292_lo_buf_o2_p_spl_,
    n292_lo_buf_o2_p
  );


  buf

  (
    n280_lo_buf_o2_n_spl_,
    n280_lo_buf_o2_n
  );


  buf

  (
    n280_lo_buf_o2_n_spl_0,
    n280_lo_buf_o2_n_spl_
  );


  buf

  (
    n292_lo_buf_o2_n_spl_,
    n292_lo_buf_o2_n
  );


  buf

  (
    n292_lo_buf_o2_n_spl_0,
    n292_lo_buf_o2_n_spl_
  );


  buf

  (
    n280_lo_buf_o2_p_spl_,
    n280_lo_buf_o2_p
  );


  buf

  (
    n316_lo_buf_o2_p_spl_,
    n316_lo_buf_o2_p
  );


  buf

  (
    n304_lo_buf_o2_n_spl_,
    n304_lo_buf_o2_n
  );


  buf

  (
    n304_lo_buf_o2_n_spl_0,
    n304_lo_buf_o2_n_spl_
  );


  buf

  (
    n316_lo_buf_o2_n_spl_,
    n316_lo_buf_o2_n
  );


  buf

  (
    n316_lo_buf_o2_n_spl_0,
    n316_lo_buf_o2_n_spl_
  );


  buf

  (
    n304_lo_buf_o2_p_spl_,
    n304_lo_buf_o2_p
  );


  buf

  (
    n340_lo_buf_o2_p_spl_,
    n340_lo_buf_o2_p
  );


  buf

  (
    n328_lo_buf_o2_n_spl_,
    n328_lo_buf_o2_n
  );


  buf

  (
    n328_lo_buf_o2_n_spl_0,
    n328_lo_buf_o2_n_spl_
  );


  buf

  (
    n340_lo_buf_o2_n_spl_,
    n340_lo_buf_o2_n
  );


  buf

  (
    n340_lo_buf_o2_n_spl_0,
    n340_lo_buf_o2_n_spl_
  );


  buf

  (
    n328_lo_buf_o2_p_spl_,
    n328_lo_buf_o2_p
  );


  buf

  (
    n364_lo_buf_o2_p_spl_,
    n364_lo_buf_o2_p
  );


  buf

  (
    n352_lo_buf_o2_n_spl_,
    n352_lo_buf_o2_n
  );


  buf

  (
    n352_lo_buf_o2_n_spl_0,
    n352_lo_buf_o2_n_spl_
  );


  buf

  (
    n364_lo_buf_o2_n_spl_,
    n364_lo_buf_o2_n
  );


  buf

  (
    n364_lo_buf_o2_n_spl_0,
    n364_lo_buf_o2_n_spl_
  );


  buf

  (
    n352_lo_buf_o2_p_spl_,
    n352_lo_buf_o2_p
  );


  buf

  (
    n388_lo_buf_o2_p_spl_,
    n388_lo_buf_o2_p
  );


  buf

  (
    n376_lo_buf_o2_n_spl_,
    n376_lo_buf_o2_n
  );


  buf

  (
    n376_lo_buf_o2_n_spl_0,
    n376_lo_buf_o2_n_spl_
  );


  buf

  (
    n388_lo_buf_o2_n_spl_,
    n388_lo_buf_o2_n
  );


  buf

  (
    n388_lo_buf_o2_n_spl_0,
    n388_lo_buf_o2_n_spl_
  );


  buf

  (
    n376_lo_buf_o2_p_spl_,
    n376_lo_buf_o2_p
  );


  buf

  (
    n412_lo_buf_o2_p_spl_,
    n412_lo_buf_o2_p
  );


  buf

  (
    n400_lo_buf_o2_n_spl_,
    n400_lo_buf_o2_n
  );


  buf

  (
    n400_lo_buf_o2_n_spl_0,
    n400_lo_buf_o2_n_spl_
  );


  buf

  (
    n412_lo_buf_o2_n_spl_,
    n412_lo_buf_o2_n
  );


  buf

  (
    n412_lo_buf_o2_n_spl_0,
    n412_lo_buf_o2_n_spl_
  );


  buf

  (
    n400_lo_buf_o2_p_spl_,
    n400_lo_buf_o2_p
  );


  buf

  (
    n436_lo_buf_o2_p_spl_,
    n436_lo_buf_o2_p
  );


  buf

  (
    n424_lo_buf_o2_n_spl_,
    n424_lo_buf_o2_n
  );


  buf

  (
    n424_lo_buf_o2_n_spl_0,
    n424_lo_buf_o2_n_spl_
  );


  buf

  (
    n436_lo_buf_o2_n_spl_,
    n436_lo_buf_o2_n
  );


  buf

  (
    n436_lo_buf_o2_n_spl_0,
    n436_lo_buf_o2_n_spl_
  );


  buf

  (
    n424_lo_buf_o2_p_spl_,
    n424_lo_buf_o2_p
  );


  buf

  (
    n460_lo_buf_o2_p_spl_,
    n460_lo_buf_o2_p
  );


  buf

  (
    n448_lo_buf_o2_n_spl_,
    n448_lo_buf_o2_n
  );


  buf

  (
    n448_lo_buf_o2_n_spl_0,
    n448_lo_buf_o2_n_spl_
  );


  buf

  (
    n460_lo_buf_o2_n_spl_,
    n460_lo_buf_o2_n
  );


  buf

  (
    n460_lo_buf_o2_n_spl_0,
    n460_lo_buf_o2_n_spl_
  );


  buf

  (
    n448_lo_buf_o2_p_spl_,
    n448_lo_buf_o2_p
  );


  buf

  (
    n484_lo_buf_o2_p_spl_,
    n484_lo_buf_o2_p
  );


  buf

  (
    n472_lo_buf_o2_n_spl_,
    n472_lo_buf_o2_n
  );


  buf

  (
    n472_lo_buf_o2_n_spl_0,
    n472_lo_buf_o2_n_spl_
  );


  buf

  (
    n484_lo_buf_o2_n_spl_,
    n484_lo_buf_o2_n
  );


  buf

  (
    n484_lo_buf_o2_n_spl_0,
    n484_lo_buf_o2_n_spl_
  );


  buf

  (
    n472_lo_buf_o2_p_spl_,
    n472_lo_buf_o2_p
  );


  buf

  (
    n508_lo_buf_o2_p_spl_,
    n508_lo_buf_o2_p
  );


  buf

  (
    n496_lo_buf_o2_n_spl_,
    n496_lo_buf_o2_n
  );


  buf

  (
    n496_lo_buf_o2_n_spl_0,
    n496_lo_buf_o2_n_spl_
  );


  buf

  (
    n508_lo_buf_o2_n_spl_,
    n508_lo_buf_o2_n
  );


  buf

  (
    n508_lo_buf_o2_n_spl_0,
    n508_lo_buf_o2_n_spl_
  );


  buf

  (
    n496_lo_buf_o2_p_spl_,
    n496_lo_buf_o2_p
  );


  buf

  (
    n532_lo_buf_o2_p_spl_,
    n532_lo_buf_o2_p
  );


  buf

  (
    n520_lo_buf_o2_n_spl_,
    n520_lo_buf_o2_n
  );


  buf

  (
    n520_lo_buf_o2_n_spl_0,
    n520_lo_buf_o2_n_spl_
  );


  buf

  (
    n532_lo_buf_o2_n_spl_,
    n532_lo_buf_o2_n
  );


  buf

  (
    n532_lo_buf_o2_n_spl_0,
    n532_lo_buf_o2_n_spl_
  );


  buf

  (
    n520_lo_buf_o2_p_spl_,
    n520_lo_buf_o2_p
  );


  buf

  (
    n556_lo_buf_o2_p_spl_,
    n556_lo_buf_o2_p
  );


  buf

  (
    n544_lo_buf_o2_n_spl_,
    n544_lo_buf_o2_n
  );


  buf

  (
    n544_lo_buf_o2_n_spl_0,
    n544_lo_buf_o2_n_spl_
  );


  buf

  (
    n556_lo_buf_o2_n_spl_,
    n556_lo_buf_o2_n
  );


  buf

  (
    n556_lo_buf_o2_n_spl_0,
    n556_lo_buf_o2_n_spl_
  );


  buf

  (
    n544_lo_buf_o2_p_spl_,
    n544_lo_buf_o2_p
  );


  buf

  (
    n580_lo_buf_o2_p_spl_,
    n580_lo_buf_o2_p
  );


  buf

  (
    n568_lo_buf_o2_n_spl_,
    n568_lo_buf_o2_n
  );


  buf

  (
    n568_lo_buf_o2_n_spl_0,
    n568_lo_buf_o2_n_spl_
  );


  buf

  (
    n580_lo_buf_o2_n_spl_,
    n580_lo_buf_o2_n
  );


  buf

  (
    n580_lo_buf_o2_n_spl_0,
    n580_lo_buf_o2_n_spl_
  );


  buf

  (
    n568_lo_buf_o2_p_spl_,
    n568_lo_buf_o2_p
  );


  buf

  (
    n604_lo_buf_o2_p_spl_,
    n604_lo_buf_o2_p
  );


  buf

  (
    n592_lo_buf_o2_n_spl_,
    n592_lo_buf_o2_n
  );


  buf

  (
    n592_lo_buf_o2_n_spl_0,
    n592_lo_buf_o2_n_spl_
  );


  buf

  (
    n604_lo_buf_o2_n_spl_,
    n604_lo_buf_o2_n
  );


  buf

  (
    n604_lo_buf_o2_n_spl_0,
    n604_lo_buf_o2_n_spl_
  );


  buf

  (
    n592_lo_buf_o2_p_spl_,
    n592_lo_buf_o2_p
  );


  buf

  (
    n628_lo_buf_o2_p_spl_,
    n628_lo_buf_o2_p
  );


  buf

  (
    n616_lo_buf_o2_n_spl_,
    n616_lo_buf_o2_n
  );


  buf

  (
    n616_lo_buf_o2_n_spl_0,
    n616_lo_buf_o2_n_spl_
  );


  buf

  (
    n628_lo_buf_o2_n_spl_,
    n628_lo_buf_o2_n
  );


  buf

  (
    n628_lo_buf_o2_n_spl_0,
    n628_lo_buf_o2_n_spl_
  );


  buf

  (
    n616_lo_buf_o2_p_spl_,
    n616_lo_buf_o2_p
  );


  buf

  (
    n652_lo_buf_o2_p_spl_,
    n652_lo_buf_o2_p
  );


  buf

  (
    n640_lo_buf_o2_n_spl_,
    n640_lo_buf_o2_n
  );


  buf

  (
    n640_lo_buf_o2_n_spl_0,
    n640_lo_buf_o2_n_spl_
  );


  buf

  (
    n652_lo_buf_o2_n_spl_,
    n652_lo_buf_o2_n
  );


  buf

  (
    n652_lo_buf_o2_n_spl_0,
    n652_lo_buf_o2_n_spl_
  );


  buf

  (
    n640_lo_buf_o2_p_spl_,
    n640_lo_buf_o2_p
  );


endmodule
