// Benchmark "mymod" written by ABC on Sun Oct 29 23:44:46 2023

module mymod (  
    G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
    G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
    G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44,
    G45, G46, G47, G48, G49, G50,
    G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528,
    G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538,
    G3539, G3540  );
  
  input  G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14,
    G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42,
    G43, G44, G45, G46, G47, G48, G49, G50;
  output G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528,
    G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538,
    G3539, G3540;
  reg n1752_lo, n1776_lo, n1824_lo, n1836_lo, n1848_lo, n1860_lo, n1872_lo,
    n1884_lo, n1896_lo, n1908_lo, n1911_lo, n1914_lo, n1923_lo, n1926_lo,
    n1935_lo, n1938_lo, n1947_lo, n1950_lo, n1959_lo, n1962_lo, n1971_lo,
    n1974_lo, n1983_lo, n1995_lo, n2055_lo, n2064_lo, n2067_lo, n2079_lo,
    n2100_lo, n2112_lo, n2124_lo, n2136_lo, n2148_lo, n2160_lo, n2172_lo,
    n2184_lo, n2235_lo, n2238_lo, n2247_lo, n2250_lo, n2259_lo, n2262_lo,
    n2271_lo, n2274_lo, n2283_lo, n2286_lo, n2289_lo, n2295_lo, n2298_lo,
    n2304_lo, n2307_lo, n2316_lo, n2331_lo, n2334_lo, n2337_lo, n2340_lo,
    n2071_o2, n2080_o2, n2137_o2, n2368_o2, n2383_o2, n2405_o2, n2471_o2,
    n2617_o2, n2765_o2, n2775_o2, n2829_o2, n2579_o2, n2580_o2, n2618_o2,
    n2619_o2, n2620_o2, n2621_o2, n2622_o2, n2623_o2, n2624_o2, n2625_o2,
    n2626_o2, n2627_o2, n3029_o2, n3035_o2, n2643_o2, n2644_o2, n2645_o2,
    n327_inv, n2658_o2, n2659_o2, n2674_o2, n2675_o2, n2676_o2, n3119_o2,
    n3153_o2, n351_inv, n2729_o2, n2730_o2, n2731_o2, n698_o2, n366_inv,
    n2757_o2, n2758_o2, n1000_o2, n1160_o2, n1153_o2, n2793_o2, n2794_o2,
    n2795_o2, n1001_o2, n2859_o2, n744_o2, n402_inv, n2926_o2, n408_inv,
    n2966_o2, n2967_o2, n2947_o2, n1010_o2, n2976_o2, n3069_o2, n3028_o2,
    n3081_o2, n3082_o2, n3142_o2, n3214_o2, n2992_o2, n2993_o2, n870_o2,
    n3086_o2, n3087_o2, n3088_o2, n3089_o2, n3090_o2, n3091_o2, n3092_o2,
    n3093_o2, n3094_o2, n3095_o2, n483_inv, n3170_o2, n3171_o2, n3172_o2,
    n3179_o2, n498_inv, n3193_o2, n3211_o2, n3212_o2, n3213_o2, n513_inv,
    n1125_o2, n1081_o2, n1139_o2, n3245_o2, n3246_o2, n3247_o2,
    lo074_buf_o2, lo078_buf_o2, lo186_buf_o2, lo118_buf_o2, lo146_buf_o2,
    n1038_o2, n1044_o2, n555_inv, n558_inv, lo026_buf_o2, lo030_buf_o2,
    lo090_buf_o2, lo094_buf_o2, lo098_buf_o2, lo102_buf_o2, lo066_buf_o2,
    lo070_buf_o2, n1202_o2, n1003_o2, n1031_o2, n1034_o2, n1040_o2,
    n1046_o2, n1380_o2, n1425_o2, n697_o2, n1143_o2, n673_o2, n789_o2,
    n786_o2, n1047_o2, n1036_o2, n1307_o2, n1035_o2, n1297_o2, n1099_o2,
    n1128_o2, n645_inv, n826_o2, n853_o2, n654_inv, n700_o2, n884_o2,
    lo082_buf_o2, lo086_buf_o2, n801_o2, n840_o2, n675_inv, lo002_buf_o2,
    lo010_buf_o2, lo166_buf_o2, lo170_buf_o2, n1426_o2, n1082_o2, n1310_o2,
    n1015_o2, n1206_o2, n1262_o2, n1456_o2, n1244_o2, n1280_o2, n1290_o2,
    n1012_o2, n1074_o2, n1112_o2, n1212_o2, n1454_o2, n1182_o2, n1220_o2,
    n701_o2, n744_inv, n1282_o2, n1144_o2, n1278_o2, n1459_o2, n1324_o2,
    n1288_o2, n1271_o2, n1132_o2, n1231_o2, n1462_o2, n1482_o2, n994_o2,
    n998_o2, lo106_buf_o2, n769_o2, n814_o2, n841_o2, n867_o2,
    lo006_buf_o2, lo014_buf_o2, lo022_buf_o2, lo042_buf_o2, lo046_buf_o2,
    lo050_buf_o2, lo054_buf_o2, lo130_buf_o2, lo134_buf_o2, lo154_buf_o2,
    lo174_buf_o2, lo178_buf_o2, n1007_o2, n1294_o2, n1084_o2, n1399_o2,
    n1311_o2, n1392_o2, n1102_o2, n1041_o2, n1298_o2, n738_o2, n1214_o2,
    n1222_o2, n1155_o2, n1147_o2, n1393_o2, n999_o2, n1306_o2, n1312_o2,
    n1382_o2, n1383_o2, n1152_o2, n1334_o2, n1335_o2, n906_inv, n773_o2,
    lo190_buf_o2, n1368_o2, n1362_o2, n1406_o2, n1403_o2, n741_o2,
    n1407_o2, n1395_o2, n1359_o2, n1159_o2, n1221_o2, n945_inv, n989_o2,
    n881_o2, n1340_o2, n1341_o2, n906_o2, n1388_o2, n791_o2, n1372_o2,
    n815_o2, n868_o2, lo018_buf_o2, lo138_buf_o2, lo158_buf_o2, n780_o2,
    n728_o2, n993_inv, n929_o2, n955_o2, n938_o2, n1117_o2, n1121_o2,
    n965_o2, n752_o2, n753_o2, n760_o2, n770_o2, n923_o2, n947_o2, n897_o2,
    n919_o2, n895_o2, n917_o2, n751_o2, n774_o2, lo126_buf_o2,
    lo142_buf_o2, lo162_buf_o2, n1059_inv, n792_o2, n869_o2, n1068_inv,
    lo024_buf_o2, lo028_buf_o2, lo088_buf_o2, lo092_buf_o2, lo096_buf_o2,
    lo100_buf_o2, n763_o2, n754_o2, n755_o2, n822_o2, n849_o2, n777_o2,
    n778_o2, n820_o2, n846_o2, n806_o2, n771_o2, n854_o2, n828_o2,
    lo117_buf_o2, lo145_buf_o2, n762_o2, n805_o2, n859_o2, n833_o2,
    lo034_buf_o2, lo038_buf_o2, lo122_buf_o2, lo150_buf_o2;
  wire new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n807_, new_n809_,
    new_n811_, new_n813_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n825_, new_n827_, new_n829_,
    new_n831_, new_n833_, new_n835_, new_n837_, new_n839_, new_n841_,
    new_n843_, new_n845_, new_n847_, new_n849_, new_n851_, new_n853_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n871_, new_n872_, new_n873_, new_n875_, new_n877_, new_n879_,
    new_n881_, new_n883_, new_n885_, new_n887_, new_n889_, new_n891_,
    new_n893_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n919_, new_n921_, new_n923_,
    new_n925_, new_n927_, new_n929_, new_n931_, new_n933_, new_n935_,
    new_n937_, new_n938_, new_n939_, new_n941_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n949_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n969_, new_n970_, new_n971_,
    new_n973_, new_n975_, new_n977_, new_n979_, new_n981_, new_n983_,
    new_n985_, new_n988_, new_n989_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1001_, new_n1003_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1012_, new_n1014_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1021_, new_n1023_, new_n1025_, new_n1026_,
    new_n1027_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1049_, new_n1051_, new_n1052_, new_n1053_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1068_, new_n1069_, new_n1071_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1079_,
    new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1087_,
    new_n1088_, new_n1090_, new_n1091_, new_n1093_, new_n1095_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1115_, new_n1116_, new_n1117_,
    new_n1119_, new_n1121_, new_n1123_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1139_, new_n1140_, new_n1141_,
    new_n1143_, new_n1144_, new_n1145_, new_n1147_, new_n1149_, new_n1150_,
    new_n1151_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1163_, new_n1165_,
    new_n1167_, new_n1169_, new_n1171_, new_n1173_, new_n1174_, new_n1175_,
    new_n1177_, new_n1180_, new_n1181_, new_n1183_, new_n1185_, new_n1187_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1194_, new_n1195_,
    new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1201_, new_n1202_,
    new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1209_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1217_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1225_,
    new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_,
    new_n1233_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1249_, new_n1251_, new_n1254_, new_n1255_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1263_, new_n1265_,
    new_n1267_, new_n1269_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1277_, new_n1279_, new_n1281_, new_n1283_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1316_, new_n1317_, new_n1318_, new_n1319_,
    new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1338_, new_n1339_, new_n1341_, new_n1343_, new_n1344_, new_n1345_,
    new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1371_, new_n1372_,
    new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1379_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1397_, new_n1398_, new_n1399_,
    new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1406_,
    new_n1408_, new_n1410_, new_n1411_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1420_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_,
    new_n1430_, new_n1431_, new_n1433_, new_n1434_, new_n1435_, new_n1437_,
    new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1451_,
    new_n1452_, new_n1453_, new_n1456_, new_n1458_, new_n1460_, new_n1462_,
    new_n1463_, new_n1464_, new_n1466_, new_n1467_, new_n1469_, new_n1471_,
    new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1489_, new_n1490_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1503_, new_n1504_,
    new_n1505_, new_n1507_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1523_, new_n1524_, new_n1525_,
    new_n1526_, new_n1527_, new_n1529_, new_n1530_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1551_,
    new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_,
    new_n1565_, new_n1566_, new_n1567_, new_n1569_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_,
    new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_,
    new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_,
    new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_,
    new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_,
    new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_,
    new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_,
    new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_,
    new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_,
    new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_,
    new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_,
    new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_,
    new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2094_,
    new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_,
    new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_,
    new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_,
    new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_,
    new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_,
    new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_,
    new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_,
    new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_,
    new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_,
    new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_,
    new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_,
    new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_,
    new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_,
    new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_,
    new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_,
    new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_,
    new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_,
    new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_,
    new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_,
    new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_,
    new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_,
    new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_,
    new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_,
    new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_,
    new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_,
    new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_,
    new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_,
    new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_,
    new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_,
    new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_,
    new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_,
    new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_,
    new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_,
    new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_,
    new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_,
    new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_,
    new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_,
    new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_,
    new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_,
    new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_,
    new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_,
    new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_,
    new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_,
    new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_,
    new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_,
    new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_,
    new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_,
    new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_,
    new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_,
    new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_,
    new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_,
    new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_,
    new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_,
    new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_,
    new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_,
    new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_,
    new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_,
    new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_,
    new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_,
    new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_,
    new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_,
    new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_,
    new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_,
    new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_,
    new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_,
    new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_,
    new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_,
    new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_,
    new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_,
    new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_,
    new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_,
    new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_,
    new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_,
    new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_,
    new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_,
    new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_,
    new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_,
    new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_,
    new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_,
    new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_,
    new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_,
    new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_,
    new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_,
    new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_,
    new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_,
    new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_,
    new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_,
    new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_,
    new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_,
    new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_,
    new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_,
    new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_,
    new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_,
    new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_,
    new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_,
    new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_,
    new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_,
    new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_,
    new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_,
    new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_,
    new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_,
    new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_,
    new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_,
    new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_,
    new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_,
    new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_,
    new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_,
    new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_,
    new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_,
    new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_,
    new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_,
    new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_,
    new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_,
    new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_,
    new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_,
    new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_,
    new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_,
    new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_,
    new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_,
    new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_,
    new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_,
    new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_,
    new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_,
    new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_,
    new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_,
    new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_,
    new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_,
    new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_,
    new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_,
    new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_,
    new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_,
    new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_,
    new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_,
    new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_,
    new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_,
    new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_,
    new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_,
    new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_,
    new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_,
    new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_,
    new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_,
    new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_,
    new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_,
    new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_,
    new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_,
    new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_,
    new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_,
    new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_,
    new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_,
    new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_,
    new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_,
    new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_,
    new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_,
    new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_,
    new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_,
    new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_,
    new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_,
    new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_,
    new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_,
    new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_,
    new_n3870_, n4070_li003_li003, n4094_li011_li011, n4142_li027_li027,
    n4154_li031_li031, n4166_li035_li035, n4178_li039_li039,
    n4190_li043_li043, n4202_li047_li047, n4214_li051_li051,
    n4226_li055_li055, n4229_li056_li056, n4232_li057_li057,
    n4241_li060_li060, n4244_li061_li061, n4253_li064_li064,
    n4256_li065_li065, n4265_li068_li068, n4268_li069_li069,
    n4277_li072_li072, n4280_li073_li073, n4289_li076_li076,
    n4292_li077_li077, n4301_li080_li080, n4313_li084_li084,
    n4373_li104_li104, n4382_li107_li107, n4385_li108_li108,
    n4397_li112_li112, n4418_li119_li119, n4430_li123_li123,
    n4442_li127_li127, n4454_li131_li131, n4466_li135_li135,
    n4478_li139_li139, n4490_li143_li143, n4502_li147_li147,
    n4553_li164_li164, n4556_li165_li165, n4565_li168_li168,
    n4568_li169_li169, n4577_li172_li172, n4580_li173_li173,
    n4589_li176_li176, n4592_li177_li177, n4601_li180_li180,
    n4604_li181_li181, n4607_li182_li182, n4613_li184_li184,
    n4616_li185_li185, n4622_li187_li187, n4625_li188_li188,
    n4634_li191_li191, n4649_li196_li196, n4652_li197_li197,
    n4655_li198_li198, n4658_li199_li199, n2071_i2, n2080_i2, n2137_i2,
    n2368_i2, n2383_i2, n2405_i2, n2471_i2, n2617_i2, n2765_i2, n2775_i2,
    n2829_i2, n2579_i2, n2580_i2, n2618_i2, n2619_i2, n2620_i2, n2621_i2,
    n2622_i2, n2623_i2, n2624_i2, n2625_i2, n2626_i2, n2627_i2, n3029_i2,
    n3035_i2, n2643_i2, n2644_i2, n2645_i2, n2640_i2, n2658_i2, n2659_i2,
    n2674_i2, n2675_i2, n2676_i2, n3119_i2, n3153_i2, n2681_i2, n2729_i2,
    n2730_i2, n2731_i2, n698_i2, n677_i2, n2757_i2, n2758_i2, n1000_i2,
    n1160_i2, n1153_i2, n2793_i2, n2794_i2, n2795_i2, n1001_i2, n2859_i2,
    n744_i2, n2908_i2, n2926_i2, n2928_i2, n2966_i2, n2967_i2, n2947_i2,
    n1010_i2, n2976_i2, n3069_i2, n3028_i2, n3081_i2, n3082_i2, n3142_i2,
    n3214_i2, n2992_i2, n2993_i2, n870_i2, n3086_i2, n3087_i2, n3088_i2,
    n3089_i2, n3090_i2, n3091_i2, n3092_i2, n3093_i2, n3094_i2, n3095_i2,
    n3136_i2, n3170_i2, n3171_i2, n3172_i2, n3179_i2, n3180_i2, n3193_i2,
    n3211_i2, n3212_i2, n3213_i2, n3219_i2, n1125_i2, n1081_i2, n1139_i2,
    n3245_i2, n3246_i2, n3247_i2, lo074_buf_i2, lo078_buf_i2, lo186_buf_i2,
    lo118_buf_i2, lo146_buf_i2, n1038_i2, n1044_i2, n980_i2, n1145_i2,
    lo026_buf_i2, lo030_buf_i2, lo090_buf_i2, lo094_buf_i2, lo098_buf_i2,
    lo102_buf_i2, lo066_buf_i2, lo070_buf_i2, n1202_i2, n1003_i2, n1031_i2,
    n1034_i2, n1040_i2, n1046_i2, n1380_i2, n1425_i2, n697_i2, n1143_i2,
    n673_i2, n789_i2, n786_i2, n1047_i2, n1036_i2, n1307_i2, n1035_i2,
    n1297_i2, n1099_i2, n1128_i2, n674_i2, n826_i2, n853_i2, n951_i2,
    n700_i2, n884_i2, lo082_buf_i2, lo086_buf_i2, n801_i2, n840_i2,
    n866_i2, lo002_buf_i2, lo010_buf_i2, lo166_buf_i2, lo170_buf_i2,
    n1426_i2, n1082_i2, n1310_i2, n1015_i2, n1206_i2, n1262_i2, n1456_i2,
    n1244_i2, n1280_i2, n1290_i2, n1012_i2, n1074_i2, n1112_i2, n1212_i2,
    n1454_i2, n1182_i2, n1220_i2, n701_i2, n973_i2, n1282_i2, n1144_i2,
    n1278_i2, n1459_i2, n1324_i2, n1288_i2, n1271_i2, n1132_i2, n1231_i2,
    n1462_i2, n1482_i2, n994_i2, n998_i2, lo106_buf_i2, n769_i2, n814_i2,
    n841_i2, n867_i2, lo006_buf_i2, lo014_buf_i2, lo022_buf_i2,
    lo042_buf_i2, lo046_buf_i2, lo050_buf_i2, lo054_buf_i2, lo130_buf_i2,
    lo134_buf_i2, lo154_buf_i2, lo174_buf_i2, lo178_buf_i2, n1007_i2,
    n1294_i2, n1084_i2, n1399_i2, n1311_i2, n1392_i2, n1102_i2, n1041_i2,
    n1298_i2, n738_i2, n1214_i2, n1222_i2, n1155_i2, n1147_i2, n1393_i2,
    n999_i2, n1306_i2, n1312_i2, n1382_i2, n1383_i2, n1152_i2, n1334_i2,
    n1335_i2, n695_i2, n773_i2, lo190_buf_i2, n1368_i2, n1362_i2, n1406_i2,
    n1403_i2, n741_i2, n1407_i2, n1395_i2, n1359_i2, n1159_i2, n1221_i2,
    n987_i2, n989_i2, n881_i2, n1340_i2, n1341_i2, n906_i2, n1388_i2,
    n791_i2, n1372_i2, n815_i2, n868_i2, lo018_buf_i2, lo138_buf_i2,
    lo158_buf_i2, n780_i2, n728_i2, n676_i2, n929_i2, n955_i2, n938_i2,
    n1117_i2, n1121_i2, n965_i2, n752_i2, n753_i2, n760_i2, n770_i2,
    n923_i2, n947_i2, n897_i2, n919_i2, n895_i2, n917_i2, n751_i2, n774_i2,
    lo126_buf_i2, lo142_buf_i2, lo162_buf_i2, n990_i2, n792_i2, n869_i2,
    n848_i2, lo024_buf_i2, lo028_buf_i2, lo088_buf_i2, lo092_buf_i2,
    lo096_buf_i2, lo100_buf_i2, n763_i2, n754_i2, n755_i2, n822_i2,
    n849_i2, n777_i2, n778_i2, n820_i2, n846_i2, n806_i2, n771_i2, n854_i2,
    n828_i2, lo117_buf_i2, lo145_buf_i2, n762_i2, n805_i2, n859_i2,
    n833_i2, lo034_buf_i2, lo038_buf_i2, lo122_buf_i2, lo150_buf_i2;
  assign new_n795_ = G1;
  assign new_n796_ = ~G1;
  assign new_n797_ = G2;
  assign new_n798_ = ~G2;
  assign new_n799_ = G3;
  assign new_n800_ = ~G3;
  assign new_n801_ = G4;
  assign new_n802_ = ~G4;
  assign new_n803_ = G5;
  assign new_n805_ = G6;
  assign new_n807_ = G7;
  assign new_n809_ = G8;
  assign new_n811_ = G9;
  assign new_n813_ = G10;
  assign new_n815_ = G11;
  assign new_n817_ = G12;
  assign new_n818_ = ~G12;
  assign new_n819_ = G13;
  assign new_n820_ = ~G13;
  assign new_n821_ = G14;
  assign new_n823_ = G15;
  assign new_n825_ = G16;
  assign new_n827_ = G17;
  assign new_n829_ = G18;
  assign new_n831_ = G19;
  assign new_n833_ = G20;
  assign new_n835_ = G21;
  assign new_n837_ = G22;
  assign new_n839_ = G23;
  assign new_n841_ = G24;
  assign new_n843_ = G25;
  assign new_n845_ = G26;
  assign new_n847_ = G27;
  assign new_n849_ = G28;
  assign new_n851_ = G29;
  assign new_n853_ = G30;
  assign new_n855_ = G31;
  assign new_n857_ = G32;
  assign new_n858_ = ~G32;
  assign new_n859_ = G33;
  assign new_n860_ = ~G33;
  assign new_n861_ = G34;
  assign new_n862_ = ~G34;
  assign new_n863_ = G35;
  assign new_n865_ = G36;
  assign new_n866_ = ~G36;
  assign new_n867_ = G37;
  assign new_n869_ = G38;
  assign new_n871_ = G39;
  assign new_n872_ = ~G39;
  assign new_n873_ = G40;
  assign new_n875_ = G41;
  assign new_n877_ = G42;
  assign new_n879_ = G43;
  assign new_n881_ = G44;
  assign new_n883_ = G45;
  assign new_n885_ = G46;
  assign new_n887_ = G47;
  assign new_n889_ = G48;
  assign new_n891_ = G49;
  assign new_n893_ = G50;
  assign new_n896_ = ~n1752_lo;
  assign new_n897_ = n1776_lo;
  assign new_n898_ = ~n1776_lo;
  assign new_n899_ = n1824_lo;
  assign new_n900_ = ~n1824_lo;
  assign new_n901_ = n1836_lo;
  assign new_n903_ = n1848_lo;
  assign new_n904_ = ~n1848_lo;
  assign new_n905_ = n1860_lo;
  assign new_n906_ = ~n1860_lo;
  assign new_n907_ = n1872_lo;
  assign new_n908_ = ~n1872_lo;
  assign new_n909_ = n1884_lo;
  assign new_n910_ = ~n1884_lo;
  assign new_n911_ = n1896_lo;
  assign new_n912_ = ~n1896_lo;
  assign new_n913_ = n1908_lo;
  assign new_n914_ = ~n1908_lo;
  assign new_n915_ = n1911_lo;
  assign new_n917_ = n1914_lo;
  assign new_n919_ = n1923_lo;
  assign new_n921_ = n1926_lo;
  assign new_n923_ = n1935_lo;
  assign new_n925_ = n1938_lo;
  assign new_n927_ = n1947_lo;
  assign new_n929_ = n1950_lo;
  assign new_n931_ = n1959_lo;
  assign new_n933_ = n1962_lo;
  assign new_n935_ = n1971_lo;
  assign new_n937_ = n1974_lo;
  assign new_n938_ = ~n1974_lo;
  assign new_n939_ = n1983_lo;
  assign new_n941_ = n1995_lo;
  assign new_n943_ = n2055_lo;
  assign new_n944_ = ~n2055_lo;
  assign new_n945_ = n2064_lo;
  assign new_n946_ = ~n2064_lo;
  assign new_n947_ = n2067_lo;
  assign new_n949_ = n2079_lo;
  assign new_n951_ = n2100_lo;
  assign new_n952_ = ~n2100_lo;
  assign new_n953_ = n2112_lo;
  assign new_n954_ = ~n2112_lo;
  assign new_n955_ = n2124_lo;
  assign new_n956_ = ~n2124_lo;
  assign new_n957_ = n2136_lo;
  assign new_n958_ = ~n2136_lo;
  assign new_n959_ = n2148_lo;
  assign new_n960_ = ~n2148_lo;
  assign new_n961_ = n2160_lo;
  assign new_n962_ = ~n2160_lo;
  assign new_n963_ = n2172_lo;
  assign new_n964_ = ~n2172_lo;
  assign new_n965_ = n2184_lo;
  assign new_n966_ = ~n2184_lo;
  assign new_n967_ = n2235_lo;
  assign new_n969_ = n2238_lo;
  assign new_n970_ = ~n2238_lo;
  assign new_n971_ = n2247_lo;
  assign new_n973_ = n2250_lo;
  assign new_n975_ = n2259_lo;
  assign new_n977_ = n2262_lo;
  assign new_n979_ = n2271_lo;
  assign new_n981_ = n2274_lo;
  assign new_n983_ = n2283_lo;
  assign new_n985_ = n2286_lo;
  assign new_n988_ = ~n2289_lo;
  assign new_n989_ = n2295_lo;
  assign new_n991_ = n2298_lo;
  assign new_n992_ = ~n2298_lo;
  assign new_n993_ = n2304_lo;
  assign new_n994_ = ~n2304_lo;
  assign new_n995_ = n2307_lo;
  assign new_n996_ = ~n2307_lo;
  assign new_n997_ = n2316_lo;
  assign new_n998_ = ~n2316_lo;
  assign new_n999_ = n2331_lo;
  assign new_n1001_ = n2334_lo;
  assign new_n1003_ = n2337_lo;
  assign new_n1005_ = n2340_lo;
  assign new_n1006_ = ~n2340_lo;
  assign new_n1007_ = n2071_o2;
  assign new_n1008_ = ~n2071_o2;
  assign new_n1009_ = n2080_o2;
  assign new_n1010_ = ~n2080_o2;
  assign new_n1012_ = ~n2137_o2;
  assign new_n1014_ = ~n2368_o2;
  assign new_n1016_ = ~n2383_o2;
  assign new_n1017_ = n2405_o2;
  assign new_n1018_ = ~n2405_o2;
  assign new_n1019_ = n2471_o2;
  assign new_n1021_ = n2617_o2;
  assign new_n1023_ = n2765_o2;
  assign new_n1025_ = n2775_o2;
  assign new_n1026_ = ~n2775_o2;
  assign new_n1027_ = n2829_o2;
  assign new_n1029_ = n2579_o2;
  assign new_n1030_ = ~n2579_o2;
  assign new_n1031_ = n2580_o2;
  assign new_n1032_ = ~n2580_o2;
  assign new_n1033_ = n2618_o2;
  assign new_n1035_ = n2619_o2;
  assign new_n1036_ = ~n2619_o2;
  assign new_n1037_ = n2620_o2;
  assign new_n1038_ = ~n2620_o2;
  assign new_n1039_ = n2621_o2;
  assign new_n1040_ = ~n2621_o2;
  assign new_n1041_ = n2622_o2;
  assign new_n1042_ = ~n2622_o2;
  assign new_n1043_ = n2623_o2;
  assign new_n1044_ = ~n2623_o2;
  assign new_n1045_ = n2624_o2;
  assign new_n1046_ = ~n2624_o2;
  assign new_n1047_ = n2625_o2;
  assign new_n1049_ = n2626_o2;
  assign new_n1051_ = n2627_o2;
  assign new_n1052_ = ~n2627_o2;
  assign new_n1053_ = n3029_o2;
  assign new_n1055_ = n3035_o2;
  assign new_n1056_ = ~n3035_o2;
  assign new_n1057_ = n2643_o2;
  assign new_n1058_ = ~n2643_o2;
  assign new_n1059_ = n2644_o2;
  assign new_n1061_ = n2645_o2;
  assign new_n1062_ = ~n2645_o2;
  assign new_n1063_ = n327_inv;
  assign new_n1064_ = ~n327_inv;
  assign new_n1065_ = n2658_o2;
  assign new_n1068_ = ~n2659_o2;
  assign new_n1069_ = n2674_o2;
  assign new_n1071_ = n2675_o2;
  assign new_n1073_ = n2676_o2;
  assign new_n1074_ = ~n2676_o2;
  assign new_n1075_ = n3119_o2;
  assign new_n1076_ = ~n3119_o2;
  assign new_n1077_ = n3153_o2;
  assign new_n1079_ = n351_inv;
  assign new_n1081_ = n2729_o2;
  assign new_n1082_ = ~n2729_o2;
  assign new_n1083_ = n2730_o2;
  assign new_n1084_ = ~n2730_o2;
  assign new_n1085_ = n2731_o2;
  assign new_n1087_ = n698_o2;
  assign new_n1088_ = ~n698_o2;
  assign new_n1090_ = ~n366_inv;
  assign new_n1091_ = n2757_o2;
  assign new_n1093_ = n2758_o2;
  assign new_n1095_ = n1000_o2;
  assign new_n1097_ = n1160_o2;
  assign new_n1098_ = ~n1160_o2;
  assign new_n1099_ = n1153_o2;
  assign new_n1100_ = ~n1153_o2;
  assign new_n1101_ = n2793_o2;
  assign new_n1102_ = ~n2793_o2;
  assign new_n1103_ = n2794_o2;
  assign new_n1104_ = ~n2794_o2;
  assign new_n1105_ = n2795_o2;
  assign new_n1106_ = ~n2795_o2;
  assign new_n1107_ = n1001_o2;
  assign new_n1108_ = ~n1001_o2;
  assign new_n1110_ = ~n2859_o2;
  assign new_n1111_ = n744_o2;
  assign new_n1112_ = ~n744_o2;
  assign new_n1113_ = n402_inv;
  assign new_n1115_ = n2926_o2;
  assign new_n1116_ = ~n2926_o2;
  assign new_n1117_ = n408_inv;
  assign new_n1119_ = n2966_o2;
  assign new_n1121_ = n2967_o2;
  assign new_n1123_ = n2947_o2;
  assign new_n1125_ = n1010_o2;
  assign new_n1126_ = ~n1010_o2;
  assign new_n1127_ = n2976_o2;
  assign new_n1128_ = ~n2976_o2;
  assign new_n1129_ = n3069_o2;
  assign new_n1131_ = n3028_o2;
  assign new_n1132_ = ~n3028_o2;
  assign new_n1133_ = n3081_o2;
  assign new_n1134_ = ~n3081_o2;
  assign new_n1135_ = n3082_o2;
  assign new_n1136_ = ~n3082_o2;
  assign new_n1137_ = n3142_o2;
  assign new_n1139_ = n3214_o2;
  assign new_n1140_ = ~n3214_o2;
  assign new_n1141_ = n2992_o2;
  assign new_n1143_ = n2993_o2;
  assign new_n1144_ = ~n2993_o2;
  assign new_n1145_ = n870_o2;
  assign new_n1147_ = n3086_o2;
  assign new_n1149_ = n3087_o2;
  assign new_n1150_ = ~n3087_o2;
  assign new_n1151_ = n3088_o2;
  assign new_n1153_ = n3089_o2;
  assign new_n1154_ = ~n3089_o2;
  assign new_n1155_ = n3090_o2;
  assign new_n1156_ = ~n3090_o2;
  assign new_n1157_ = n3091_o2;
  assign new_n1158_ = ~n3091_o2;
  assign new_n1159_ = n3092_o2;
  assign new_n1160_ = ~n3092_o2;
  assign new_n1161_ = n3093_o2;
  assign new_n1163_ = n3094_o2;
  assign new_n1165_ = n3095_o2;
  assign new_n1167_ = n483_inv;
  assign new_n1169_ = n3170_o2;
  assign new_n1171_ = n3171_o2;
  assign new_n1173_ = n3172_o2;
  assign new_n1174_ = ~n3172_o2;
  assign new_n1175_ = n3179_o2;
  assign new_n1177_ = n498_inv;
  assign new_n1180_ = ~n3193_o2;
  assign new_n1181_ = n3211_o2;
  assign new_n1183_ = n3212_o2;
  assign new_n1185_ = n3213_o2;
  assign new_n1187_ = n513_inv;
  assign new_n1189_ = n1125_o2;
  assign new_n1190_ = ~n1125_o2;
  assign new_n1191_ = n1081_o2;
  assign new_n1192_ = ~n1081_o2;
  assign new_n1194_ = ~n1139_o2;
  assign new_n1195_ = n3245_o2;
  assign new_n1196_ = ~n3245_o2;
  assign new_n1197_ = n3246_o2;
  assign new_n1198_ = ~n3246_o2;
  assign new_n1199_ = n3247_o2;
  assign new_n1201_ = lo074_buf_o2;
  assign new_n1202_ = ~lo074_buf_o2;
  assign new_n1203_ = lo078_buf_o2;
  assign new_n1204_ = ~lo078_buf_o2;
  assign new_n1205_ = lo186_buf_o2;
  assign new_n1206_ = ~lo186_buf_o2;
  assign new_n1207_ = lo118_buf_o2;
  assign new_n1209_ = lo146_buf_o2;
  assign new_n1211_ = n1038_o2;
  assign new_n1212_ = ~n1038_o2;
  assign new_n1213_ = n1044_o2;
  assign new_n1214_ = ~n1044_o2;
  assign new_n1215_ = n555_inv;
  assign new_n1217_ = n558_inv;
  assign new_n1219_ = lo026_buf_o2;
  assign new_n1220_ = ~lo026_buf_o2;
  assign new_n1221_ = lo030_buf_o2;
  assign new_n1222_ = ~lo030_buf_o2;
  assign new_n1223_ = lo090_buf_o2;
  assign new_n1225_ = lo094_buf_o2;
  assign new_n1226_ = ~lo094_buf_o2;
  assign new_n1227_ = lo098_buf_o2;
  assign new_n1228_ = ~lo098_buf_o2;
  assign new_n1229_ = lo102_buf_o2;
  assign new_n1230_ = ~lo102_buf_o2;
  assign new_n1231_ = lo066_buf_o2;
  assign new_n1233_ = lo070_buf_o2;
  assign new_n1236_ = ~n1202_o2;
  assign new_n1237_ = n1003_o2;
  assign new_n1238_ = ~n1003_o2;
  assign new_n1239_ = n1031_o2;
  assign new_n1240_ = ~n1031_o2;
  assign new_n1241_ = n1034_o2;
  assign new_n1242_ = ~n1034_o2;
  assign new_n1243_ = n1040_o2;
  assign new_n1244_ = ~n1040_o2;
  assign new_n1245_ = n1046_o2;
  assign new_n1246_ = ~n1046_o2;
  assign new_n1247_ = n1380_o2;
  assign new_n1249_ = n1425_o2;
  assign new_n1251_ = n697_o2;
  assign new_n1254_ = ~n1143_o2;
  assign new_n1255_ = n673_o2;
  assign new_n1257_ = n789_o2;
  assign new_n1258_ = ~n789_o2;
  assign new_n1259_ = n786_o2;
  assign new_n1260_ = ~n786_o2;
  assign new_n1261_ = n1047_o2;
  assign new_n1263_ = n1036_o2;
  assign new_n1265_ = n1307_o2;
  assign new_n1267_ = n1035_o2;
  assign new_n1269_ = n1297_o2;
  assign new_n1272_ = ~n1099_o2;
  assign new_n1273_ = n1128_o2;
  assign new_n1274_ = ~n1128_o2;
  assign new_n1275_ = n645_inv;
  assign new_n1277_ = n826_o2;
  assign new_n1279_ = n853_o2;
  assign new_n1281_ = n654_inv;
  assign new_n1283_ = n700_o2;
  assign new_n1285_ = n884_o2;
  assign new_n1286_ = ~n884_o2;
  assign new_n1287_ = lo082_buf_o2;
  assign new_n1288_ = ~lo082_buf_o2;
  assign new_n1289_ = lo086_buf_o2;
  assign new_n1290_ = ~lo086_buf_o2;
  assign new_n1291_ = n801_o2;
  assign new_n1292_ = ~n801_o2;
  assign new_n1293_ = n840_o2;
  assign new_n1294_ = ~n840_o2;
  assign new_n1295_ = n675_inv;
  assign new_n1296_ = ~n675_inv;
  assign new_n1297_ = lo002_buf_o2;
  assign new_n1298_ = ~lo002_buf_o2;
  assign new_n1299_ = lo010_buf_o2;
  assign new_n1300_ = ~lo010_buf_o2;
  assign new_n1301_ = lo166_buf_o2;
  assign new_n1302_ = ~lo166_buf_o2;
  assign new_n1303_ = lo170_buf_o2;
  assign new_n1304_ = ~lo170_buf_o2;
  assign new_n1305_ = n1426_o2;
  assign new_n1306_ = ~n1426_o2;
  assign new_n1307_ = n1082_o2;
  assign new_n1308_ = ~n1082_o2;
  assign new_n1310_ = ~n1310_o2;
  assign new_n1311_ = n1015_o2;
  assign new_n1312_ = ~n1015_o2;
  assign new_n1313_ = n1206_o2;
  assign new_n1316_ = ~n1262_o2;
  assign new_n1317_ = n1456_o2;
  assign new_n1318_ = ~n1456_o2;
  assign new_n1319_ = n1244_o2;
  assign new_n1320_ = ~n1244_o2;
  assign new_n1321_ = n1280_o2;
  assign new_n1322_ = ~n1280_o2;
  assign new_n1323_ = n1290_o2;
  assign new_n1324_ = ~n1290_o2;
  assign new_n1325_ = n1012_o2;
  assign new_n1326_ = ~n1012_o2;
  assign new_n1327_ = n1074_o2;
  assign new_n1328_ = ~n1074_o2;
  assign new_n1329_ = n1112_o2;
  assign new_n1330_ = ~n1112_o2;
  assign new_n1331_ = n1212_o2;
  assign new_n1332_ = ~n1212_o2;
  assign new_n1333_ = n1454_o2;
  assign new_n1334_ = ~n1454_o2;
  assign new_n1335_ = n1182_o2;
  assign new_n1336_ = ~n1182_o2;
  assign new_n1337_ = n1220_o2;
  assign new_n1338_ = ~n1220_o2;
  assign new_n1339_ = n701_o2;
  assign new_n1341_ = n744_inv;
  assign new_n1343_ = n1282_o2;
  assign new_n1344_ = ~n1282_o2;
  assign new_n1345_ = n1144_o2;
  assign new_n1347_ = n1278_o2;
  assign new_n1348_ = ~n1278_o2;
  assign new_n1349_ = n1459_o2;
  assign new_n1350_ = ~n1459_o2;
  assign new_n1351_ = n1324_o2;
  assign new_n1352_ = ~n1324_o2;
  assign new_n1353_ = n1288_o2;
  assign new_n1354_ = ~n1288_o2;
  assign new_n1356_ = ~n1271_o2;
  assign new_n1357_ = n1132_o2;
  assign new_n1358_ = ~n1132_o2;
  assign new_n1359_ = n1231_o2;
  assign new_n1360_ = ~n1231_o2;
  assign new_n1361_ = n1462_o2;
  assign new_n1362_ = ~n1462_o2;
  assign new_n1363_ = n1482_o2;
  assign new_n1364_ = ~n1482_o2;
  assign new_n1365_ = n994_o2;
  assign new_n1366_ = ~n994_o2;
  assign new_n1367_ = n998_o2;
  assign new_n1368_ = ~n998_o2;
  assign new_n1369_ = lo106_buf_o2;
  assign new_n1371_ = n769_o2;
  assign new_n1372_ = ~n769_o2;
  assign new_n1373_ = n814_o2;
  assign new_n1374_ = ~n814_o2;
  assign new_n1375_ = n841_o2;
  assign new_n1376_ = ~n841_o2;
  assign new_n1377_ = n867_o2;
  assign new_n1379_ = lo006_buf_o2;
  assign new_n1381_ = lo014_buf_o2;
  assign new_n1382_ = ~lo014_buf_o2;
  assign new_n1383_ = lo022_buf_o2;
  assign new_n1384_ = ~lo022_buf_o2;
  assign new_n1385_ = lo042_buf_o2;
  assign new_n1386_ = ~lo042_buf_o2;
  assign new_n1387_ = lo046_buf_o2;
  assign new_n1388_ = ~lo046_buf_o2;
  assign new_n1389_ = lo050_buf_o2;
  assign new_n1390_ = ~lo050_buf_o2;
  assign new_n1391_ = lo054_buf_o2;
  assign new_n1392_ = ~lo054_buf_o2;
  assign new_n1393_ = lo130_buf_o2;
  assign new_n1394_ = ~lo130_buf_o2;
  assign new_n1395_ = lo134_buf_o2;
  assign new_n1397_ = lo154_buf_o2;
  assign new_n1398_ = ~lo154_buf_o2;
  assign new_n1399_ = lo174_buf_o2;
  assign new_n1400_ = ~lo174_buf_o2;
  assign new_n1401_ = lo178_buf_o2;
  assign new_n1402_ = ~lo178_buf_o2;
  assign new_n1403_ = n1007_o2;
  assign new_n1404_ = ~n1007_o2;
  assign new_n1406_ = ~n1294_o2;
  assign new_n1408_ = ~n1084_o2;
  assign new_n1410_ = ~n1399_o2;
  assign new_n1411_ = n1311_o2;
  assign new_n1414_ = ~n1392_o2;
  assign new_n1415_ = n1102_o2;
  assign new_n1416_ = ~n1102_o2;
  assign new_n1417_ = n1041_o2;
  assign new_n1418_ = ~n1041_o2;
  assign new_n1420_ = ~n1298_o2;
  assign new_n1421_ = n738_o2;
  assign new_n1422_ = ~n738_o2;
  assign new_n1423_ = n1214_o2;
  assign new_n1424_ = ~n1214_o2;
  assign new_n1425_ = n1222_o2;
  assign new_n1426_ = ~n1222_o2;
  assign new_n1427_ = n1155_o2;
  assign new_n1428_ = ~n1155_o2;
  assign new_n1429_ = n1147_o2;
  assign new_n1430_ = ~n1147_o2;
  assign new_n1431_ = n1393_o2;
  assign new_n1433_ = n999_o2;
  assign new_n1434_ = ~n999_o2;
  assign new_n1435_ = n1306_o2;
  assign new_n1437_ = n1312_o2;
  assign new_n1439_ = n1382_o2;
  assign new_n1440_ = ~n1382_o2;
  assign new_n1441_ = n1383_o2;
  assign new_n1442_ = ~n1383_o2;
  assign new_n1443_ = n1152_o2;
  assign new_n1444_ = ~n1152_o2;
  assign new_n1445_ = n1334_o2;
  assign new_n1446_ = ~n1334_o2;
  assign new_n1447_ = n1335_o2;
  assign new_n1448_ = ~n1335_o2;
  assign new_n1449_ = n906_inv;
  assign new_n1451_ = n773_o2;
  assign new_n1452_ = ~n773_o2;
  assign new_n1453_ = lo190_buf_o2;
  assign new_n1456_ = ~n1368_o2;
  assign new_n1458_ = ~n1362_o2;
  assign new_n1460_ = ~n1406_o2;
  assign new_n1462_ = ~n1403_o2;
  assign new_n1463_ = n741_o2;
  assign new_n1464_ = ~n741_o2;
  assign new_n1466_ = ~n1407_o2;
  assign new_n1467_ = n1395_o2;
  assign new_n1469_ = n1359_o2;
  assign new_n1471_ = n1159_o2;
  assign new_n1472_ = ~n1159_o2;
  assign new_n1473_ = n1221_o2;
  assign new_n1474_ = ~n1221_o2;
  assign new_n1475_ = n945_inv;
  assign new_n1476_ = ~n945_inv;
  assign new_n1477_ = n989_o2;
  assign new_n1478_ = ~n989_o2;
  assign new_n1479_ = n881_o2;
  assign new_n1480_ = ~n881_o2;
  assign new_n1481_ = n1340_o2;
  assign new_n1482_ = ~n1340_o2;
  assign new_n1483_ = n1341_o2;
  assign new_n1484_ = ~n1341_o2;
  assign new_n1485_ = n906_o2;
  assign new_n1486_ = ~n906_o2;
  assign new_n1487_ = n1388_o2;
  assign new_n1489_ = n791_o2;
  assign new_n1490_ = ~n791_o2;
  assign new_n1492_ = ~n1372_o2;
  assign new_n1493_ = n815_o2;
  assign new_n1494_ = ~n815_o2;
  assign new_n1495_ = n868_o2;
  assign new_n1496_ = ~n868_o2;
  assign new_n1497_ = lo018_buf_o2;
  assign new_n1498_ = ~lo018_buf_o2;
  assign new_n1499_ = lo138_buf_o2;
  assign new_n1500_ = ~lo138_buf_o2;
  assign new_n1501_ = lo158_buf_o2;
  assign new_n1503_ = n780_o2;
  assign new_n1504_ = ~n780_o2;
  assign new_n1505_ = n728_o2;
  assign new_n1507_ = n993_inv;
  assign new_n1509_ = n929_o2;
  assign new_n1510_ = ~n929_o2;
  assign new_n1511_ = n955_o2;
  assign new_n1512_ = ~n955_o2;
  assign new_n1513_ = n938_o2;
  assign new_n1514_ = ~n938_o2;
  assign new_n1515_ = n1117_o2;
  assign new_n1516_ = ~n1117_o2;
  assign new_n1517_ = n1121_o2;
  assign new_n1518_ = ~n1121_o2;
  assign new_n1519_ = n965_o2;
  assign new_n1520_ = ~n965_o2;
  assign new_n1521_ = n752_o2;
  assign new_n1523_ = n753_o2;
  assign new_n1524_ = ~n753_o2;
  assign new_n1525_ = n760_o2;
  assign new_n1526_ = ~n760_o2;
  assign new_n1527_ = n770_o2;
  assign new_n1529_ = n923_o2;
  assign new_n1530_ = ~n923_o2;
  assign new_n1531_ = n947_o2;
  assign new_n1532_ = ~n947_o2;
  assign new_n1533_ = n897_o2;
  assign new_n1534_ = ~n897_o2;
  assign new_n1535_ = n919_o2;
  assign new_n1536_ = ~n919_o2;
  assign new_n1537_ = n895_o2;
  assign new_n1538_ = ~n895_o2;
  assign new_n1539_ = n917_o2;
  assign new_n1540_ = ~n917_o2;
  assign new_n1541_ = n751_o2;
  assign new_n1542_ = ~n751_o2;
  assign new_n1543_ = n774_o2;
  assign new_n1544_ = ~n774_o2;
  assign new_n1545_ = lo126_buf_o2;
  assign new_n1546_ = ~lo126_buf_o2;
  assign new_n1547_ = lo142_buf_o2;
  assign new_n1548_ = ~lo142_buf_o2;
  assign new_n1549_ = lo162_buf_o2;
  assign new_n1551_ = n1059_inv;
  assign new_n1552_ = ~n1059_inv;
  assign new_n1553_ = n792_o2;
  assign new_n1554_ = ~n792_o2;
  assign new_n1555_ = n869_o2;
  assign new_n1556_ = ~n869_o2;
  assign new_n1557_ = n1068_inv;
  assign new_n1559_ = lo024_buf_o2;
  assign new_n1560_ = ~lo024_buf_o2;
  assign new_n1561_ = lo028_buf_o2;
  assign new_n1562_ = ~lo028_buf_o2;
  assign new_n1563_ = lo088_buf_o2;
  assign new_n1564_ = ~lo088_buf_o2;
  assign new_n1565_ = lo092_buf_o2;
  assign new_n1566_ = ~lo092_buf_o2;
  assign new_n1567_ = lo096_buf_o2;
  assign new_n1569_ = lo100_buf_o2;
  assign new_n1571_ = n763_o2;
  assign new_n1572_ = ~n763_o2;
  assign new_n1573_ = n754_o2;
  assign new_n1574_ = ~n754_o2;
  assign new_n1575_ = n755_o2;
  assign new_n1576_ = ~n755_o2;
  assign new_n1577_ = n822_o2;
  assign new_n1578_ = ~n822_o2;
  assign new_n1579_ = n849_o2;
  assign new_n1580_ = ~n849_o2;
  assign new_n1581_ = n777_o2;
  assign new_n1582_ = ~n777_o2;
  assign new_n1583_ = n778_o2;
  assign new_n1584_ = ~n778_o2;
  assign new_n1585_ = n820_o2;
  assign new_n1586_ = ~n820_o2;
  assign new_n1587_ = n846_o2;
  assign new_n1588_ = ~n846_o2;
  assign new_n1589_ = n806_o2;
  assign new_n1590_ = ~n806_o2;
  assign new_n1591_ = n771_o2;
  assign new_n1592_ = ~n771_o2;
  assign new_n1593_ = n854_o2;
  assign new_n1594_ = ~n854_o2;
  assign new_n1595_ = n828_o2;
  assign new_n1596_ = ~n828_o2;
  assign new_n1597_ = lo117_buf_o2;
  assign new_n1598_ = ~lo117_buf_o2;
  assign new_n1599_ = lo145_buf_o2;
  assign new_n1600_ = ~lo145_buf_o2;
  assign new_n1601_ = n762_o2;
  assign new_n1602_ = ~n762_o2;
  assign new_n1603_ = n805_o2;
  assign new_n1604_ = ~n805_o2;
  assign new_n1605_ = n859_o2;
  assign new_n1606_ = ~n859_o2;
  assign new_n1607_ = n833_o2;
  assign new_n1608_ = ~n833_o2;
  assign new_n1609_ = lo034_buf_o2;
  assign new_n1610_ = ~lo034_buf_o2;
  assign new_n1611_ = lo038_buf_o2;
  assign new_n1612_ = ~lo038_buf_o2;
  assign new_n1613_ = lo122_buf_o2;
  assign new_n1614_ = ~lo122_buf_o2;
  assign new_n1615_ = lo150_buf_o2;
  assign new_n1616_ = ~lo150_buf_o2;
  assign new_n1617_ = new_n1014_ & new_n3063_;
  assign new_n1618_ = new_n3064_ & new_n3065_;
  assign new_n1619_ = new_n3067_ | new_n3069_;
  assign new_n1620_ = new_n3071_ | new_n903_;
  assign new_n1621_ = new_n1620_ & new_n1619_;
  assign new_n1622_ = new_n3073_ | new_n3074_;
  assign new_n1623_ = new_n3076_ | new_n905_;
  assign new_n1624_ = new_n1623_ & new_n1622_;
  assign new_n1625_ = new_n1624_ & new_n1621_;
  assign new_n1626_ = new_n3078_ | new_n3080_;
  assign new_n1627_ = new_n3082_ | new_n901_;
  assign new_n1628_ = new_n1627_ & new_n1626_;
  assign new_n1629_ = new_n3084_ | new_n3086_;
  assign new_n1630_ = new_n3088_ | new_n3091_;
  assign new_n1631_ = new_n1630_ & new_n1629_;
  assign new_n1632_ = new_n1631_ & new_n1628_;
  assign new_n1633_ = new_n1632_ & new_n1625_;
  assign new_n1634_ = new_n1633_ | new_n1618_;
  assign new_n1635_ = new_n1007_ & new_n3064_;
  assign new_n1636_ = new_n1008_ | new_n897_;
  assign new_n1637_ = new_n3092_ | new_n1088_;
  assign new_n1638_ = new_n3088_ & new_n3084_;
  assign new_n1639_ = new_n1638_ | new_n3067_;
  assign new_n1640_ = new_n1639_ | new_n1019_;
  assign new_n1641_ = new_n1640_ & new_n1637_;
  assign new_n1642_ = new_n1641_ & new_n1634_;
  assign new_n1643_ = new_n3078_ & new_n3093_;
  assign new_n1644_ = new_n3094_ | new_n3089_;
  assign new_n1645_ = new_n3094_ & new_n3089_;
  assign new_n1646_ = new_n3077_ | new_n3093_;
  assign new_n1647_ = new_n1646_ & new_n1644_;
  assign new_n1648_ = new_n1645_ | new_n1643_;
  assign new_n1649_ = new_n3085_ & new_n3095_;
  assign new_n1650_ = new_n3096_ | new_n3068_;
  assign new_n1651_ = new_n3096_ & new_n3068_;
  assign new_n1652_ = new_n3085_ | new_n3095_;
  assign new_n1653_ = new_n1652_ & new_n1650_;
  assign new_n1654_ = new_n1651_ | new_n1649_;
  assign new_n1655_ = new_n3097_ & new_n3098_;
  assign new_n1656_ = new_n3099_ | new_n3100_;
  assign new_n1657_ = new_n3099_ & new_n3100_;
  assign new_n1658_ = new_n3097_ | new_n3098_;
  assign new_n1659_ = new_n1658_ & new_n1656_;
  assign new_n1660_ = new_n1657_ | new_n1655_;
  assign new_n1661_ = new_n3076_ & new_n3101_;
  assign new_n1662_ = new_n3102_ | new_n3071_;
  assign new_n1663_ = new_n3102_ & new_n3070_;
  assign new_n1664_ = new_n3075_ | new_n3101_;
  assign new_n1665_ = new_n1664_ & new_n1662_;
  assign new_n1666_ = new_n1663_ | new_n1661_;
  assign new_n1667_ = new_n3082_ & new_n3103_;
  assign new_n1668_ = new_n3104_ | new_n3073_;
  assign new_n1669_ = new_n3104_ & new_n3072_;
  assign new_n1670_ = new_n3081_ | new_n3103_;
  assign new_n1671_ = new_n1670_ & new_n1668_;
  assign new_n1672_ = new_n1669_ | new_n1667_;
  assign new_n1673_ = new_n3105_ & new_n3106_;
  assign new_n1674_ = new_n3107_ | new_n3108_;
  assign new_n1675_ = new_n3107_ & new_n3108_;
  assign new_n1676_ = new_n3105_ | new_n3106_;
  assign new_n1677_ = new_n1676_ & new_n1674_;
  assign new_n1678_ = new_n1675_ | new_n1673_;
  assign new_n1679_ = new_n1677_ | new_n1659_;
  assign new_n1680_ = new_n1678_ | new_n1660_;
  assign new_n1681_ = new_n1680_ & new_n1679_;
  assign new_n1682_ = new_n3086_ & new_n3069_;
  assign new_n1683_ = new_n910_ | new_n908_;
  assign new_n1684_ = new_n1683_ & new_n1009_;
  assign new_n1685_ = new_n1682_ | new_n1010_;
  assign new_n1686_ = new_n3110_ & new_n3091_;
  assign new_n1687_ = new_n3080_ | new_n3111_;
  assign new_n1688_ = new_n3079_ & new_n3111_;
  assign new_n1689_ = new_n3110_ | new_n3090_;
  assign new_n1690_ = new_n1689_ & new_n1687_;
  assign new_n1691_ = new_n1688_ | new_n1686_;
  assign new_n1692_ = new_n3112_ & new_n3113_;
  assign new_n1693_ = new_n3114_ | new_n3115_;
  assign new_n1694_ = new_n3114_ & new_n3115_;
  assign new_n1695_ = new_n3112_ | new_n3113_;
  assign new_n1696_ = new_n1695_ & new_n1693_;
  assign new_n1697_ = new_n1694_ | new_n1692_;
  assign new_n1698_ = new_n1697_ & new_n1112_;
  assign new_n1699_ = new_n1696_ & new_n1111_;
  assign new_n1700_ = new_n1699_ | new_n1698_;
  assign new_n1701_ = new_n3116_ & new_n1021_;
  assign new_n1702_ = new_n3116_ & new_n1023_;
  assign new_n1703_ = new_n1702_ | new_n1077_;
  assign new_n1704_ = new_n3118_ & new_n1087_;
  assign new_n1705_ = new_n1027_ & new_n3065_;
  assign new_n1706_ = new_n1705_ | new_n1704_;
  assign new_n1707_ = new_n1326_ & new_n3119_;
  assign new_n1708_ = new_n1325_ | new_n3120_;
  assign new_n1709_ = new_n1327_ & new_n1312_;
  assign new_n1710_ = new_n1328_ | new_n1311_;
  assign new_n1711_ = new_n1710_ & new_n1708_;
  assign new_n1712_ = new_n1709_ | new_n1707_;
  assign new_n1713_ = new_n1329_ & new_n1308_;
  assign new_n1714_ = new_n1330_ | new_n1307_;
  assign new_n1715_ = new_n1357_ & new_n3119_;
  assign new_n1716_ = new_n1358_ | new_n3120_;
  assign new_n1717_ = new_n1716_ & new_n1714_;
  assign new_n1718_ = new_n1715_ | new_n1713_;
  assign new_n1719_ = new_n1055_ & new_n1025_;
  assign new_n1720_ = new_n1056_ | new_n1026_;
  assign new_n1721_ = new_n3121_ & new_n3122_;
  assign new_n1722_ = new_n3123_ | new_n3124_;
  assign new_n1723_ = new_n3123_ & new_n3124_;
  assign new_n1724_ = new_n3121_ | new_n3122_;
  assign new_n1725_ = new_n1724_ & new_n1722_;
  assign new_n1726_ = new_n1723_ | new_n1721_;
  assign new_n1727_ = new_n1726_ & new_n993_;
  assign new_n1728_ = new_n1725_ | new_n994_;
  assign new_n1729_ = new_n3125_ & new_n3126_;
  assign new_n1730_ = new_n3127_ | new_n3128_;
  assign new_n1731_ = new_n3127_ & new_n3128_;
  assign new_n1732_ = new_n3125_ | new_n3126_;
  assign new_n1733_ = new_n1732_ & new_n1730_;
  assign new_n1734_ = new_n1731_ | new_n1729_;
  assign new_n1735_ = new_n1733_ & new_n1727_;
  assign new_n1736_ = new_n1734_ & new_n1728_;
  assign new_n1737_ = new_n1736_ | new_n1735_;
  assign new_n1738_ = new_n3092_ & new_n1017_;
  assign new_n1739_ = new_n1738_ & new_n1737_;
  assign new_n1740_ = new_n1635_ & new_n3109_;
  assign new_n1741_ = new_n1740_ & new_n1012_;
  assign new_n1742_ = new_n1016_ & new_n3063_;
  assign new_n1743_ = new_n1742_ | new_n3074_;
  assign new_n1744_ = new_n904_ | new_n900_;
  assign new_n1745_ = new_n1744_ & new_n1018_;
  assign new_n1746_ = new_n1745_ & new_n1743_;
  assign new_n1747_ = new_n1746_ | new_n1741_;
  assign new_n1748_ = new_n1747_ | new_n1739_;
  assign new_n1749_ = new_n1336_ & new_n1331_;
  assign new_n1750_ = new_n1335_ | new_n1332_;
  assign new_n1751_ = new_n1359_ & new_n1320_;
  assign new_n1752_ = new_n1360_ | new_n1319_;
  assign new_n1753_ = new_n1752_ & new_n1750_;
  assign new_n1754_ = new_n1751_ | new_n1749_;
  assign new_n1755_ = new_n1343_ & new_n3118_;
  assign new_n1756_ = new_n1344_ | new_n3129_;
  assign new_n1757_ = new_n1348_ & new_n1322_;
  assign new_n1758_ = new_n1347_ | new_n1321_;
  assign new_n1759_ = new_n1757_ & new_n1756_;
  assign new_n1760_ = new_n1758_ | new_n1755_;
  assign new_n1761_ = new_n1353_ & new_n3117_;
  assign new_n1762_ = new_n1354_ | new_n3129_;
  assign new_n1763_ = new_n1352_ & new_n1324_;
  assign new_n1764_ = new_n1351_ | new_n1323_;
  assign new_n1765_ = new_n1763_ & new_n1762_;
  assign new_n1766_ = new_n1764_ | new_n1761_;
  assign new_n1767_ = new_n1333_ & new_n1306_;
  assign new_n1768_ = new_n1334_ | new_n1305_;
  assign new_n1769_ = new_n1349_ & new_n1318_;
  assign new_n1770_ = new_n1350_ | new_n1317_;
  assign new_n1771_ = new_n1770_ & new_n1768_;
  assign new_n1772_ = new_n1769_ | new_n1767_;
  assign new_n1773_ = new_n3130_ & new_n3131_;
  assign new_n1774_ = new_n3133_ | new_n3135_;
  assign new_n1775_ = new_n3136_ & new_n3137_;
  assign new_n1776_ = new_n3139_ | new_n3141_;
  assign new_n1777_ = new_n3142_ & new_n3143_;
  assign new_n1778_ = new_n3145_ | new_n3147_;
  assign new_n1779_ = new_n3148_ | new_n3149_;
  assign new_n1780_ = new_n1779_ | new_n3150_;
  assign new_n1781_ = new_n1780_ | new_n3152_;
  assign new_n1782_ = new_n997_ & new_n3153_;
  assign new_n1783_ = new_n998_ | new_n946_;
  assign new_n1784_ = new_n3154_ | new_n3152_;
  assign new_n1785_ = new_n1784_ & new_n3153_;
  assign new_n1786_ = new_n1785_ & new_n3155_;
  assign new_n1787_ = new_n3145_ & new_n3147_;
  assign new_n1788_ = new_n3142_ | new_n3143_;
  assign new_n1789_ = new_n1788_ & new_n3148_;
  assign new_n1790_ = new_n1787_ | new_n1777_;
  assign new_n1791_ = new_n3139_ & new_n3141_;
  assign new_n1792_ = new_n3136_ | new_n3137_;
  assign new_n1793_ = new_n1792_ & new_n3149_;
  assign new_n1794_ = new_n1791_ | new_n1775_;
  assign new_n1795_ = new_n3156_ & new_n3157_;
  assign new_n1796_ = new_n3158_ | new_n3159_;
  assign new_n1797_ = new_n3158_ & new_n3159_;
  assign new_n1798_ = new_n3156_ | new_n3157_;
  assign new_n1799_ = new_n1798_ & new_n1796_;
  assign new_n1800_ = new_n1797_ | new_n1795_;
  assign new_n1801_ = new_n3133_ & new_n3135_;
  assign new_n1802_ = new_n3130_ | new_n3131_;
  assign new_n1803_ = new_n1802_ & new_n3150_;
  assign new_n1804_ = new_n1801_ | new_n1773_;
  assign new_n1805_ = new_n1364_ & new_n3151_;
  assign new_n1806_ = new_n1363_ | new_n1362_;
  assign new_n1807_ = new_n3161_ & new_n3163_;
  assign new_n1808_ = new_n3165_ | new_n3167_;
  assign new_n1809_ = new_n3165_ & new_n3167_;
  assign new_n1810_ = new_n3161_ | new_n3163_;
  assign new_n1811_ = new_n1810_ & new_n1808_;
  assign new_n1812_ = new_n1809_ | new_n1807_;
  assign new_n1813_ = new_n1812_ & new_n3154_;
  assign new_n1814_ = new_n1811_ | new_n1782_;
  assign new_n1815_ = new_n3168_ & new_n3170_;
  assign new_n1816_ = new_n3172_ | new_n3174_;
  assign new_n1817_ = new_n3172_ & new_n3174_;
  assign new_n1818_ = new_n3168_ | new_n3170_;
  assign new_n1819_ = new_n1818_ & new_n1816_;
  assign new_n1820_ = new_n1817_ | new_n1815_;
  assign new_n1821_ = new_n1820_ & new_n3176_;
  assign new_n1822_ = new_n1819_ & new_n3177_;
  assign new_n1823_ = new_n1822_ | new_n1821_;
  assign new_n1824_ = new_n3162_ & new_n3175_;
  assign new_n1825_ = new_n3166_ | new_n3171_;
  assign new_n1826_ = new_n3166_ & new_n3171_;
  assign new_n1827_ = new_n3162_ | new_n3175_;
  assign new_n1828_ = new_n1827_ & new_n1825_;
  assign new_n1829_ = new_n1826_ | new_n1824_;
  assign new_n1830_ = new_n1828_ | new_n3177_;
  assign new_n1831_ = new_n1829_ | new_n3176_;
  assign new_n1832_ = new_n1831_ & new_n1830_;
  assign new_n1833_ = new_n1110_ | new_n3179_;
  assign new_n1834_ = new_n1068_ | new_n3181_;
  assign new_n1835_ = new_n1433_ & new_n3183_;
  assign new_n1836_ = new_n1434_ | new_n3184_;
  assign new_n1837_ = new_n1472_ & new_n1428_;
  assign new_n1838_ = new_n1471_ | new_n1427_;
  assign new_n1839_ = new_n1476_ & new_n1443_;
  assign new_n1840_ = new_n3185_ | new_n1444_;
  assign new_n1841_ = new_n3186_ & new_n1057_;
  assign new_n1842_ = new_n3188_ | new_n1058_;
  assign new_n1843_ = new_n1464_ & new_n1421_;
  assign new_n1844_ = new_n1463_ & new_n1422_;
  assign new_n1845_ = new_n1844_ | new_n1843_;
  assign new_n1846_ = new_n1404_ & new_n3189_;
  assign new_n1847_ = new_n3190_ | new_n3191_;
  assign new_n1848_ = new_n1847_ & new_n1030_;
  assign new_n1849_ = new_n1846_ | new_n3192_;
  assign new_n1850_ = new_n3193_ & new_n3195_;
  assign new_n1851_ = new_n3198_ | new_n3202_;
  assign new_n1852_ = new_n3204_ & new_n3205_;
  assign new_n1853_ = new_n3206_ | new_n3207_;
  assign new_n1854_ = new_n1518_ & new_n1516_;
  assign new_n1855_ = new_n1517_ | new_n1515_;
  assign new_n1856_ = new_n1854_ & new_n3211_;
  assign new_n1857_ = new_n1855_ | new_n3220_;
  assign new_n1858_ = new_n3228_ & new_n3220_;
  assign new_n1859_ = new_n1853_ | new_n3211_;
  assign new_n1860_ = new_n1859_ & new_n1857_;
  assign new_n1861_ = new_n1858_ | new_n1856_;
  assign new_n1862_ = new_n1537_ & new_n3230_;
  assign new_n1863_ = new_n1538_ | new_n3231_;
  assign new_n1864_ = new_n3221_ & new_n1479_;
  assign new_n1865_ = new_n3212_ | new_n1480_;
  assign new_n1866_ = new_n3232_ & new_n3234_;
  assign new_n1867_ = new_n3235_ | new_n3236_;
  assign new_n1868_ = new_n3235_ & new_n3236_;
  assign new_n1869_ = new_n3232_ | new_n3234_;
  assign new_n1870_ = new_n1869_ & new_n1867_;
  assign new_n1871_ = new_n1868_ | new_n1866_;
  assign new_n1872_ = new_n1539_ & new_n3238_;
  assign new_n1873_ = new_n1540_ | new_n3239_;
  assign new_n1874_ = new_n3221_ & new_n1485_;
  assign new_n1875_ = new_n3212_ | new_n1486_;
  assign new_n1876_ = new_n3240_ & new_n3242_;
  assign new_n1877_ = new_n3243_ | new_n3244_;
  assign new_n1878_ = new_n3243_ & new_n3244_;
  assign new_n1879_ = new_n3240_ | new_n3242_;
  assign new_n1880_ = new_n1879_ & new_n1877_;
  assign new_n1881_ = new_n1878_ | new_n1876_;
  assign new_n1882_ = new_n1225_ & new_n3247_;
  assign new_n1883_ = new_n1226_ | new_n3250_;
  assign new_n1884_ = new_n1227_ & new_n3247_;
  assign new_n1885_ = new_n1228_ | new_n3250_;
  assign new_n1886_ = new_n3253_ | new_n3256_;
  assign new_n1887_ = new_n1886_ | new_n3258_;
  assign new_n1888_ = new_n3253_ | new_n3260_;
  assign new_n1889_ = new_n1888_ | new_n3258_;
  assign new_n1890_ = new_n3204_ & new_n1489_;
  assign new_n1891_ = new_n3206_ | new_n3261_;
  assign new_n1892_ = new_n1495_ & new_n3262_;
  assign new_n1893_ = new_n1496_ | new_n1374_;
  assign new_n1894_ = new_n3263_ & new_n3264_;
  assign new_n1895_ = new_n1376_ | new_n1296_;
  assign new_n1896_ = new_n1895_ & new_n1294_;
  assign new_n1897_ = new_n1894_ | new_n1293_;
  assign new_n1898_ = new_n1896_ & new_n1893_;
  assign new_n1899_ = new_n1897_ | new_n1892_;
  assign new_n1900_ = new_n1898_ & new_n1891_;
  assign new_n1901_ = new_n1899_ | new_n1890_;
  assign new_n1902_ = new_n3266_ & new_n3268_;
  assign new_n1903_ = new_n1871_ | new_n1861_;
  assign new_n1904_ = new_n3269_ | new_n3271_;
  assign new_n1905_ = new_n3272_ & new_n3213_;
  assign new_n1906_ = new_n1900_ | new_n3223_;
  assign new_n1907_ = new_n3260_ & new_n3246_;
  assign new_n1908_ = new_n3256_ | new_n3249_;
  assign new_n1909_ = new_n3273_ & new_n3274_;
  assign new_n1910_ = new_n3275_ | new_n3259_;
  assign new_n1911_ = new_n3276_ & new_n3278_;
  assign new_n1912_ = new_n3280_ | new_n3254_;
  assign new_n1913_ = new_n3275_ & new_n3274_;
  assign new_n1914_ = new_n3273_ | new_n3259_;
  assign new_n1915_ = new_n3281_ & new_n3254_;
  assign new_n1916_ = new_n3282_ | new_n3278_;
  assign new_n1917_ = new_n3276_ & new_n3255_;
  assign new_n1918_ = new_n3280_ | new_n3279_;
  assign new_n1919_ = new_n3281_ & new_n3279_;
  assign new_n1920_ = new_n3282_ | new_n3255_;
  assign new_n1921_ = new_n1448_ & new_n3283_;
  assign new_n1922_ = new_n1447_ | new_n3284_;
  assign new_n1923_ = new_n1484_ & new_n1481_;
  assign new_n1924_ = new_n1483_ | new_n1482_;
  assign new_n1925_ = new_n3285_ & new_n3287_;
  assign new_n1926_ = new_n1430_ | new_n3290_;
  assign new_n1927_ = new_n1925_ & new_n1840_;
  assign new_n1928_ = new_n1926_ | new_n3292_;
  assign new_n1929_ = new_n3293_ & new_n3295_;
  assign new_n1930_ = new_n3296_ | new_n3297_;
  assign new_n1931_ = new_n3298_ & new_n1921_;
  assign new_n1932_ = new_n1929_ & new_n3300_;
  assign new_n1933_ = new_n1932_ | new_n1931_;
  assign new_n1934_ = new_n1933_ & new_n3202_;
  assign new_n1935_ = new_n3303_ | new_n1033_;
  assign new_n1936_ = new_n3308_ | new_n1254_;
  assign new_n1937_ = new_n1106_ & new_n3310_;
  assign new_n1938_ = new_n1105_ | new_n1032_;
  assign new_n1939_ = new_n1938_ & new_n3311_;
  assign new_n1940_ = new_n1937_ | new_n1064_;
  assign new_n1941_ = new_n1469_ | new_n1458_;
  assign new_n1942_ = new_n1492_ | new_n1456_;
  assign new_n1943_ = new_n1942_ & new_n1941_;
  assign new_n1944_ = new_n1943_ | new_n3314_;
  assign new_n1945_ = new_n1944_ & new_n3320_;
  assign new_n1946_ = new_n1945_ & new_n1936_;
  assign new_n1947_ = new_n3300_ & new_n3198_;
  assign new_n1948_ = new_n1947_ | new_n1946_;
  assign new_n1949_ = new_n1948_ | new_n1934_;
  assign new_n1950_ = new_n1442_ & new_n1439_;
  assign new_n1951_ = new_n1441_ | new_n1440_;
  assign new_n1952_ = new_n3325_ | new_n3308_;
  assign new_n1953_ = new_n1487_ | new_n1431_;
  assign new_n1954_ = new_n1467_ | new_n1414_;
  assign new_n1955_ = new_n1954_ | new_n1953_;
  assign new_n1956_ = new_n1462_ | new_n1410_;
  assign new_n1957_ = new_n1466_ | new_n1460_;
  assign new_n1958_ = new_n1957_ | new_n1956_;
  assign new_n1959_ = new_n1958_ & new_n1955_;
  assign new_n1960_ = new_n1959_ | new_n3314_;
  assign new_n1961_ = new_n1960_ & new_n3320_;
  assign new_n1962_ = new_n1961_ & new_n1952_;
  assign new_n1963_ = new_n3325_ & new_n3327_;
  assign new_n1964_ = new_n3328_ | new_n3329_;
  assign new_n1965_ = new_n3328_ & new_n3329_;
  assign new_n1966_ = new_n3324_ | new_n3327_;
  assign new_n1967_ = new_n1966_ & new_n1964_;
  assign new_n1968_ = new_n1965_ | new_n1963_;
  assign new_n1969_ = new_n1968_ & new_n3283_;
  assign new_n1970_ = new_n1967_ & new_n3284_;
  assign new_n1971_ = new_n1970_ | new_n1969_;
  assign new_n1972_ = new_n3295_ & new_n3299_;
  assign new_n1973_ = new_n1972_ | new_n3293_;
  assign new_n1974_ = new_n1973_ & new_n3203_;
  assign new_n1975_ = new_n1974_ | new_n3199_;
  assign new_n1976_ = new_n1975_ & new_n1971_;
  assign new_n1977_ = new_n1976_ | new_n1962_;
  assign new_n1978_ = new_n3332_ | new_n3335_;
  assign new_n1979_ = new_n3337_ & new_n1259_;
  assign new_n1980_ = new_n3338_ | new_n3339_;
  assign new_n1981_ = new_n1532_ & new_n1512_;
  assign new_n1982_ = new_n1531_ | new_n1511_;
  assign new_n1983_ = new_n3341_ & new_n1980_;
  assign new_n1984_ = new_n3343_ | new_n1979_;
  assign new_n1985_ = new_n3337_ & new_n3344_;
  assign new_n1986_ = new_n3338_ | new_n3345_;
  assign new_n1987_ = new_n1985_ & new_n3343_;
  assign new_n1988_ = new_n1986_ | new_n3341_;
  assign new_n1989_ = new_n3346_ & new_n1984_;
  assign new_n1990_ = new_n3347_ | new_n1983_;
  assign new_n1991_ = new_n3342_ & new_n1477_;
  assign new_n1992_ = new_n3340_ | new_n3349_;
  assign new_n1993_ = new_n3350_ & new_n3352_;
  assign new_n1994_ = new_n3353_ | new_n3354_;
  assign new_n1995_ = new_n3353_ & new_n3354_;
  assign new_n1996_ = new_n3350_ | new_n3352_;
  assign new_n1997_ = new_n1996_ & new_n1994_;
  assign new_n1998_ = new_n1995_ | new_n1993_;
  assign new_n1999_ = new_n3335_ | new_n3356_;
  assign new_n2000_ = new_n3358_ & new_n1564_;
  assign new_n2001_ = new_n3360_ | new_n3361_;
  assign new_n2002_ = new_n3362_ | new_n3363_;
  assign new_n2003_ = new_n3365_ & new_n3366_;
  assign new_n2004_ = new_n3368_ | new_n3369_;
  assign new_n2005_ = new_n3370_ | new_n1174_;
  assign new_n2006_ = new_n3372_ & new_n3374_;
  assign new_n2007_ = new_n3375_ | new_n3378_;
  assign new_n2008_ = new_n3381_ | new_n3383_;
  assign new_n2009_ = new_n3384_ & new_n3266_;
  assign new_n2010_ = new_n3385_ | new_n3332_;
  assign new_n2011_ = new_n3386_ & new_n1572_;
  assign new_n2012_ = new_n1601_ | new_n1571_;
  assign new_n2013_ = new_n3388_ & new_n3392_;
  assign new_n2014_ = new_n3395_ | new_n3398_;
  assign new_n2015_ = new_n3401_ & new_n3398_;
  assign new_n2016_ = new_n3405_ | new_n3392_;
  assign new_n2017_ = new_n2016_ & new_n2014_;
  assign new_n2018_ = new_n2015_ | new_n2013_;
  assign new_n2019_ = new_n3410_ & new_n3413_;
  assign new_n2020_ = new_n3331_ | new_n3416_;
  assign new_n2021_ = new_n1586_ & new_n1578_;
  assign new_n2022_ = new_n1585_ | new_n1577_;
  assign new_n2023_ = new_n2021_ & new_n2020_;
  assign new_n2024_ = new_n2022_ | new_n2019_;
  assign new_n2025_ = new_n2024_ & new_n3420_;
  assign new_n2026_ = new_n2023_ | new_n3427_;
  assign new_n2027_ = new_n2026_ & new_n2018_;
  assign new_n2028_ = new_n2025_ | new_n2017_;
  assign new_n2029_ = new_n3388_ & new_n3430_;
  assign new_n2030_ = new_n3395_ | new_n3433_;
  assign new_n2031_ = new_n3401_ & new_n3433_;
  assign new_n2032_ = new_n3405_ | new_n3430_;
  assign new_n2033_ = new_n2032_ & new_n2030_;
  assign new_n2034_ = new_n2031_ | new_n2029_;
  assign new_n2035_ = new_n3437_ & new_n3440_;
  assign new_n2036_ = new_n3442_ | new_n1575_;
  assign new_n2037_ = new_n1588_ & new_n1580_;
  assign new_n2038_ = new_n1587_ | new_n1579_;
  assign new_n2039_ = new_n2037_ & new_n2036_;
  assign new_n2040_ = new_n2038_ | new_n2035_;
  assign new_n2041_ = new_n2040_ & new_n3420_;
  assign new_n2042_ = new_n2039_ | new_n3427_;
  assign new_n2043_ = new_n2042_ & new_n2034_;
  assign new_n2044_ = new_n2041_ | new_n2033_;
  assign new_n2045_ = new_n3410_ | new_n3444_;
  assign new_n2046_ = new_n2045_ & new_n3446_;
  assign new_n2047_ = new_n3447_ | new_n3449_;
  assign new_n2048_ = new_n1615_ & new_n3453_;
  assign new_n2049_ = new_n1616_ | new_n3459_;
  assign new_n2050_ = new_n1498_ & new_n1384_;
  assign new_n2051_ = new_n3463_ | new_n3464_;
  assign new_n2052_ = new_n2051_ & new_n1298_;
  assign new_n2053_ = new_n2050_ | new_n3449_;
  assign new_n2054_ = new_n3466_ & new_n3468_;
  assign new_n2055_ = new_n3470_ | new_n3472_;
  assign new_n2056_ = new_n3419_ & new_n3475_;
  assign new_n2057_ = new_n3426_ | new_n3477_;
  assign new_n2058_ = new_n3478_ & new_n3402_;
  assign new_n2059_ = new_n3480_ | new_n3406_;
  assign new_n2060_ = new_n3481_ & new_n3483_;
  assign new_n2061_ = new_n2058_ | new_n3485_;
  assign new_n2062_ = new_n3413_ & new_n3399_;
  assign new_n2063_ = new_n3416_ | new_n3391_;
  assign new_n2064_ = new_n3487_ & new_n3489_;
  assign new_n2065_ = new_n3491_ | new_n3493_;
  assign new_n2066_ = new_n2065_ & new_n2063_;
  assign new_n2067_ = new_n2064_ | new_n2062_;
  assign new_n2068_ = new_n2067_ & new_n3421_;
  assign new_n2069_ = new_n2066_ | new_n3428_;
  assign new_n2070_ = new_n3396_ & new_n3485_;
  assign new_n2071_ = new_n3389_ | new_n3483_;
  assign new_n2072_ = new_n2071_ & new_n2069_;
  assign new_n2073_ = new_n2070_ | new_n2068_;
  assign new_n2074_ = new_n2072_ & new_n2061_;
  assign new_n2075_ = new_n2073_ | new_n2060_;
  assign new_n2076_ = new_n3468_ & new_n1452_;
  assign new_n2077_ = new_n3472_ | new_n1451_;
  assign new_n2078_ = new_n1608_ & new_n1596_;
  assign new_n2079_ = new_n1607_ | new_n1595_;
  assign new_n2080_ = new_n2079_ & new_n3453_;
  assign new_n2081_ = new_n2078_ | new_n3459_;
  assign new_n2082_ = new_n2081_ & new_n2077_;
  assign new_n2083_ = new_n2080_ | new_n2076_;
  assign new_n2084_ = new_n3494_ | new_n3496_;
  assign new_n2085_ = new_n2084_ | new_n2027_;
  assign new_n2086_ = new_n3467_ & new_n3499_;
  assign new_n2087_ = new_n3471_ | new_n3501_;
  assign new_n2088_ = new_n1606_ & new_n1594_;
  assign new_n2089_ = new_n1605_ | new_n1593_;
  assign new_n2090_ = new_n2089_ & new_n3454_;
  assign new_n2091_ = new_n2088_ | new_n3460_;
  assign new_n2092_ = new_n2091_ & new_n3503_;
  assign new_n2093_ = new_n2090_ | new_n3505_;
  assign new_n2094_ = new_n3506_ | new_n3496_;
  assign new_n2095_ = new_n2094_ | new_n2043_;
  assign new_n2096_ = new_n3309_ | new_n1194_;
  assign new_n2097_ = new_n3309_ | new_n3507_;
  assign new_n2098_ = new_n3508_ & new_n3510_;
  assign new_n2099_ = new_n3190_ | new_n3303_;
  assign new_n2100_ = new_n3512_ | new_n3514_;
  assign new_n2101_ = new_n3375_ | new_n3516_;
  assign new_n2102_ = new_n3518_ | new_n3378_;
  assign new_n2103_ = new_n3296_ & new_n3297_;
  assign new_n2104_ = new_n3514_ & new_n3287_;
  assign new_n2105_ = new_n3519_ | new_n3290_;
  assign new_n2106_ = new_n3184_ & new_n1337_;
  assign new_n2107_ = new_n3183_ | new_n1338_;
  assign new_n2108_ = new_n2107_ & new_n3520_;
  assign new_n2109_ = new_n2106_ | new_n3521_;
  assign new_n2110_ = new_n3522_ & new_n3523_;
  assign new_n2111_ = new_n3524_ | new_n3526_;
  assign new_n2112_ = new_n3524_ & new_n3526_;
  assign new_n2113_ = new_n3522_ | new_n3523_;
  assign new_n2114_ = new_n2113_ & new_n2111_;
  assign new_n2115_ = new_n2112_ | new_n2110_;
  assign new_n2116_ = new_n3527_ & new_n3528_;
  assign new_n2117_ = new_n3529_ | new_n3530_;
  assign new_n2118_ = new_n3529_ & new_n3530_;
  assign new_n2119_ = new_n3527_ | new_n3528_;
  assign new_n2120_ = new_n2119_ & new_n2117_;
  assign new_n2121_ = new_n2118_ | new_n2116_;
  assign new_n2122_ = new_n3520_ & new_n1426_;
  assign new_n2123_ = new_n3521_ | new_n1425_;
  assign new_n2124_ = new_n3531_ & new_n3532_;
  assign new_n2125_ = new_n3533_ | new_n3535_;
  assign new_n2126_ = new_n3536_ & new_n3538_;
  assign new_n2127_ = new_n3540_ | new_n3543_;
  assign new_n2128_ = new_n3540_ & new_n3543_;
  assign new_n2129_ = new_n3536_ | new_n3538_;
  assign new_n2130_ = new_n2129_ & new_n2127_;
  assign new_n2131_ = new_n2128_ | new_n2126_;
  assign new_n2132_ = new_n3545_ | new_n3546_;
  assign new_n2133_ = new_n2132_ & new_n3548_;
  assign new_n2134_ = new_n2133_ | new_n3195_;
  assign new_n2135_ = new_n2134_ & new_n3193_;
  assign new_n2136_ = new_n3551_ & new_n3199_;
  assign new_n2137_ = new_n3552_ & new_n3200_;
  assign new_n2138_ = new_n3519_ & new_n3291_;
  assign new_n2139_ = new_n2138_ | new_n3525_;
  assign new_n2140_ = new_n3186_ & new_n3304_;
  assign new_n2141_ = new_n3188_ | new_n3555_;
  assign new_n2142_ = new_n2140_ | new_n3560_;
  assign new_n2143_ = new_n3562_ & new_n3191_;
  assign new_n2144_ = new_n3563_ & new_n3189_;
  assign new_n2145_ = new_n2141_ | new_n3564_;
  assign new_n2146_ = new_n2145_ | new_n2144_;
  assign new_n2147_ = new_n2146_ | new_n2143_;
  assign new_n2148_ = new_n2147_ & new_n2142_;
  assign new_n2149_ = new_n2148_ | new_n3565_;
  assign new_n2150_ = new_n3568_ | new_n988_;
  assign new_n2151_ = new_n1400_ | new_n3571_;
  assign new_n2152_ = new_n1304_ | new_n3574_;
  assign new_n2153_ = new_n2152_ & new_n2151_;
  assign new_n2154_ = new_n2153_ & new_n2150_;
  assign new_n2155_ = new_n3574_ | new_n1052_;
  assign new_n2156_ = new_n1302_ | new_n3568_;
  assign new_n2157_ = new_n2156_ & new_n2155_;
  assign new_n2158_ = new_n3577_ | new_n3578_;
  assign new_n2159_ = new_n2158_ & new_n3555_;
  assign new_n2160_ = new_n1402_ | new_n3580_;
  assign new_n2161_ = new_n3583_ | new_n3584_;
  assign new_n2162_ = new_n2161_ & new_n2160_;
  assign new_n2163_ = new_n2162_ & new_n2159_;
  assign new_n2164_ = new_n2163_ & new_n3585_;
  assign new_n2165_ = new_n2164_ & new_n2154_;
  assign new_n2166_ = new_n3571_ | new_n3587_;
  assign new_n2167_ = new_n2166_ & new_n1267_;
  assign new_n2168_ = new_n3583_ | new_n3588_;
  assign new_n2169_ = new_n3589_ & new_n1263_;
  assign new_n2170_ = new_n2169_ & new_n2167_;
  assign new_n2171_ = new_n1417_ | new_n3567_;
  assign new_n2172_ = new_n2171_ & new_n3304_;
  assign new_n2173_ = new_n3580_ | new_n3179_;
  assign new_n2174_ = new_n2173_ & new_n1261_;
  assign new_n2175_ = new_n2174_ & new_n2172_;
  assign new_n2176_ = new_n2175_ & new_n2170_;
  assign new_n2177_ = new_n2176_ | new_n3315_;
  assign new_n2178_ = new_n2177_ | new_n2165_;
  assign new_n2179_ = new_n2178_ & new_n2149_;
  assign new_n2180_ = new_n2179_ | new_n3590_;
  assign new_n2181_ = new_n3569_ | new_n3591_;
  assign new_n2182_ = new_n3575_ | new_n3592_;
  assign new_n2183_ = new_n3581_ | new_n3578_;
  assign new_n2184_ = new_n2183_ & new_n2182_;
  assign new_n2185_ = new_n2184_ & new_n2181_;
  assign new_n2186_ = new_n3589_ & new_n3556_;
  assign new_n2187_ = new_n3577_ | new_n3593_;
  assign new_n2188_ = new_n3572_ | new_n3584_;
  assign new_n2189_ = new_n2188_ & new_n2187_;
  assign new_n2190_ = new_n2189_ & new_n2186_;
  assign new_n2191_ = new_n2190_ & new_n3585_;
  assign new_n2192_ = new_n2191_ & new_n2185_;
  assign new_n2193_ = new_n3582_ | new_n3587_;
  assign new_n2194_ = new_n3581_ | new_n1202_;
  assign new_n2195_ = new_n3572_ | new_n1204_;
  assign new_n2196_ = new_n2195_ & new_n2194_;
  assign new_n2197_ = new_n2196_ & new_n2193_;
  assign new_n2198_ = new_n1272_ | new_n3569_;
  assign new_n2199_ = new_n2198_ & new_n3306_;
  assign new_n2200_ = new_n3576_ | new_n3180_;
  assign new_n2201_ = new_n1415_ | new_n3575_;
  assign new_n2202_ = new_n2201_ & new_n2200_;
  assign new_n2203_ = new_n2202_ & new_n2199_;
  assign new_n2204_ = new_n2203_ & new_n2197_;
  assign new_n2205_ = new_n2204_ | new_n2192_;
  assign new_n2206_ = new_n2205_ & new_n3565_;
  assign new_n2207_ = new_n2206_ | new_n3590_;
  assign new_n2208_ = new_n3596_ & new_n3598_;
  assign new_n2209_ = new_n1301_ & new_n3601_;
  assign new_n2210_ = new_n3605_ | new_n3607_;
  assign new_n2211_ = new_n2210_ & new_n3612_;
  assign new_n2212_ = new_n2211_ | new_n2209_;
  assign new_n2213_ = new_n2212_ | new_n2208_;
  assign new_n2214_ = new_n3618_ | new_n3619_;
  assign new_n2215_ = new_n2214_ & new_n3622_;
  assign new_n2216_ = new_n2215_ | new_n3306_;
  assign new_n2217_ = new_n3627_ & new_n3560_;
  assign new_n2218_ = new_n3633_ & new_n3637_;
  assign new_n2219_ = new_n2218_ | new_n2217_;
  assign new_n2220_ = new_n2219_ | new_n2216_;
  assign new_n2221_ = new_n2220_ | new_n2213_;
  assign new_n2222_ = new_n3633_ & new_n3639_;
  assign new_n2223_ = new_n3601_ & new_n1203_;
  assign new_n2224_ = new_n1418_ & new_n3622_;
  assign new_n2225_ = new_n2224_ | new_n2223_;
  assign new_n2226_ = new_n2225_ | new_n2222_;
  assign new_n2227_ = new_n3612_ & new_n1236_;
  assign new_n2228_ = new_n2227_ | new_n3556_;
  assign new_n2229_ = new_n3627_ & new_n1104_;
  assign new_n2230_ = new_n2229_ | new_n1313_;
  assign new_n2231_ = new_n2230_ | new_n2228_;
  assign new_n2232_ = new_n2231_ | new_n2226_;
  assign new_n2233_ = new_n2232_ & new_n2221_;
  assign new_n2234_ = new_n2233_ | new_n3315_;
  assign new_n2235_ = new_n2234_ & new_n3321_;
  assign new_n2236_ = new_n3611_ & new_n3598_;
  assign new_n2237_ = new_n3634_ & new_n3607_;
  assign new_n2238_ = new_n2237_ | new_n2236_;
  assign new_n2239_ = new_n3602_ & new_n3618_;
  assign new_n2240_ = new_n1084_ | new_n3561_;
  assign new_n2241_ = new_n2240_ & new_n3623_;
  assign new_n2242_ = new_n2241_ | new_n2239_;
  assign new_n2243_ = new_n2242_ | new_n2238_;
  assign new_n2244_ = new_n3613_ & new_n3637_;
  assign new_n2245_ = new_n2244_ | new_n3305_;
  assign new_n2246_ = new_n3596_ & new_n3181_;
  assign new_n2247_ = new_n3628_ & new_n3619_;
  assign new_n2248_ = new_n2247_ | new_n3640_;
  assign new_n2249_ = new_n2248_ | new_n3641_;
  assign new_n2250_ = new_n2249_ | new_n2243_;
  assign new_n2251_ = new_n1231_ | new_n3639_;
  assign new_n2252_ = new_n2251_ & new_n3613_;
  assign new_n2253_ = new_n3628_ & new_n3643_;
  assign new_n2254_ = new_n3644_ & new_n3623_;
  assign new_n2255_ = new_n2254_ | new_n2253_;
  assign new_n2256_ = new_n2255_ | new_n2252_;
  assign new_n2257_ = new_n3595_ & new_n3645_;
  assign new_n2258_ = new_n3634_ & new_n1201_;
  assign new_n2259_ = new_n2258_ | new_n2257_;
  assign new_n2260_ = new_n1233_ & new_n3602_;
  assign new_n2261_ = new_n2260_ | new_n3558_;
  assign new_n2262_ = new_n2261_ | new_n2259_;
  assign new_n2263_ = new_n2262_ | new_n2256_;
  assign new_n2264_ = new_n2263_ & new_n2250_;
  assign new_n2265_ = new_n2264_ | new_n3317_;
  assign new_n2266_ = new_n2265_ & new_n3321_;
  assign new_n2267_ = new_n3646_ & new_n1115_;
  assign new_n2268_ = new_n3647_ | new_n1116_;
  assign new_n2269_ = new_n3648_ & new_n3649_;
  assign new_n2270_ = new_n3650_ | new_n3651_;
  assign new_n2271_ = new_n3650_ & new_n3651_;
  assign new_n2272_ = new_n3648_ | new_n3649_;
  assign new_n2273_ = new_n2272_ & new_n2270_;
  assign new_n2274_ = new_n2271_ | new_n2269_;
  assign new_n2275_ = new_n3653_ | new_n3512_;
  assign new_n2276_ = new_n3223_ | new_n3261_;
  assign new_n2277_ = new_n3654_ | new_n3475_;
  assign new_n2278_ = new_n1530_ & new_n1510_;
  assign new_n2279_ = new_n1529_ | new_n1509_;
  assign new_n2280_ = new_n1514_ & new_n1286_;
  assign new_n2281_ = new_n1513_ | new_n1285_;
  assign new_n2282_ = new_n3655_ | new_n3339_;
  assign new_n2283_ = new_n2282_ & new_n3657_;
  assign new_n2284_ = new_n2279_ & new_n3344_;
  assign new_n2285_ = new_n3657_ | new_n3345_;
  assign new_n2286_ = new_n2284_ & new_n2280_;
  assign new_n2287_ = new_n2285_ | new_n3655_;
  assign new_n2288_ = new_n2286_ | new_n2283_;
  assign new_n2289_ = new_n3659_ | new_n3351_;
  assign new_n2290_ = new_n3661_ | new_n3241_;
  assign new_n2291_ = new_n3662_ | new_n3233_;
  assign new_n2292_ = new_n3551_ | new_n3664_;
  assign new_n2293_ = new_n3550_ & new_n3664_;
  assign new_n2294_ = new_n3546_ | new_n3548_;
  assign new_n2295_ = new_n3665_ & new_n2292_;
  assign new_n2296_ = new_n3666_ | new_n3668_;
  assign new_n2297_ = new_n3513_ | new_n3182_;
  assign new_n2298_ = new_n3669_ & new_n3604_;
  assign new_n2299_ = new_n3597_ & new_n3608_;
  assign new_n2300_ = new_n2299_ | new_n2298_;
  assign new_n2301_ = new_n1408_ & new_n3624_;
  assign new_n2302_ = new_n3605_ & new_n3636_;
  assign new_n2303_ = new_n2302_ | new_n2301_;
  assign new_n2304_ = new_n2303_ | new_n2300_;
  assign new_n2305_ = new_n3630_ & new_n3617_;
  assign new_n2306_ = new_n1401_ & new_n3615_;
  assign new_n2307_ = new_n2306_ | new_n2305_;
  assign new_n2308_ = new_n2307_ | new_n3641_;
  assign new_n2309_ = new_n2308_ | new_n2304_;
  assign new_n2310_ = new_n3604_ & new_n3643_;
  assign new_n2311_ = new_n1416_ & new_n3615_;
  assign new_n2312_ = new_n2311_ | new_n2310_;
  assign new_n2313_ = new_n2312_ | new_n1316_;
  assign new_n2314_ = new_n3636_ & new_n3645_;
  assign new_n2315_ = new_n2314_ | new_n3640_;
  assign new_n2316_ = new_n1356_ | new_n3558_;
  assign new_n2317_ = new_n2316_ | new_n2315_;
  assign new_n2318_ = new_n2317_ | new_n2313_;
  assign new_n2319_ = new_n2318_ & new_n2309_;
  assign new_n2320_ = new_n2319_ | new_n3317_;
  assign new_n2321_ = new_n2320_ & new_n3323_;
  assign new_n2322_ = new_n2321_ & new_n2297_;
  assign new_n2323_ = new_n3294_ & new_n3200_;
  assign new_n2324_ = new_n3298_ & new_n3203_;
  assign new_n2325_ = new_n2324_ | new_n2323_;
  assign new_n2326_ = new_n3542_ | new_n3513_;
  assign new_n2327_ = new_n3630_ & new_n1082_;
  assign new_n2328_ = new_n3603_ & new_n3638_;
  assign new_n2329_ = new_n3635_ & new_n3642_;
  assign new_n2330_ = new_n2329_ | new_n2328_;
  assign new_n2331_ = new_n2330_ | new_n2327_;
  assign new_n2332_ = new_n3644_ & new_n3616_;
  assign new_n2333_ = new_n2332_ | new_n3557_;
  assign new_n2334_ = new_n1406_ & new_n3624_;
  assign new_n2335_ = new_n2334_ | new_n1269_;
  assign new_n2336_ = new_n2335_ | new_n2333_;
  assign new_n2337_ = new_n2336_ | new_n2331_;
  assign new_n2338_ = new_n3629_ & new_n3608_;
  assign new_n2339_ = new_n3669_ & new_n3616_;
  assign new_n2340_ = new_n3597_ & new_n3561_;
  assign new_n2341_ = new_n2340_ | new_n2339_;
  assign new_n2342_ = new_n2341_ | new_n2338_;
  assign new_n2343_ = new_n1435_ | new_n1265_;
  assign new_n2344_ = new_n1437_ | new_n1411_;
  assign new_n2345_ = new_n2344_ | new_n2343_;
  assign new_n2346_ = new_n2345_ | new_n1310_;
  assign new_n2347_ = new_n2346_ | new_n2342_;
  assign new_n2348_ = new_n2347_ & new_n2337_;
  assign new_n2349_ = new_n2348_ | new_n3316_;
  assign new_n2350_ = new_n2349_ & new_n3323_;
  assign new_n2351_ = new_n2350_ & new_n2326_;
  assign new_n2352_ = new_n3665_ & new_n3545_;
  assign new_n2353_ = new_n2293_ & new_n3552_;
  assign new_n2354_ = new_n2353_ | new_n2352_;
  assign new_n2355_ = new_n3671_ & new_n3672_;
  assign new_n2356_ = new_n2355_ | new_n3368_;
  assign new_n2357_ = new_n3288_ & new_n1190_;
  assign new_n2358_ = new_n3291_ | new_n1189_;
  assign new_n2359_ = new_n3549_ & new_n3507_;
  assign new_n2360_ = new_n3663_ | new_n1191_;
  assign new_n2361_ = new_n2360_ & new_n1274_;
  assign new_n2362_ = new_n2359_ | new_n1273_;
  assign new_n2363_ = new_n2361_ & new_n2357_;
  assign new_n2364_ = new_n2362_ & new_n2358_;
  assign new_n2365_ = new_n2364_ | new_n2363_;
  assign new_n2366_ = new_n3544_ & new_n3535_;
  assign new_n2367_ = new_n3539_ | new_n3532_;
  assign new_n2368_ = new_n3647_ & new_n1127_;
  assign new_n2369_ = new_n3646_ | new_n1128_;
  assign new_n2370_ = new_n3531_ & new_n3544_;
  assign new_n2371_ = new_n3533_ | new_n3539_;
  assign new_n2372_ = new_n2371_ & new_n2369_;
  assign new_n2373_ = new_n2370_ | new_n2368_;
  assign new_n2374_ = new_n3673_ & new_n3653_;
  assign new_n2375_ = new_n3674_ | new_n3675_;
  assign new_n2376_ = new_n3674_ & new_n3675_;
  assign new_n2377_ = new_n3673_ | new_n3652_;
  assign new_n2378_ = new_n2377_ & new_n2375_;
  assign new_n2379_ = new_n2376_ | new_n2374_;
  assign new_n2380_ = new_n2379_ & new_n2367_;
  assign new_n2381_ = new_n2378_ & new_n2366_;
  assign new_n2382_ = new_n2381_ | new_n2380_;
  assign new_n2383_ = new_n3677_ | new_n3679_;
  assign new_n2384_ = new_n3677_ & new_n3679_;
  assign new_n2385_ = new_n3224_ & new_n1291_;
  assign new_n2386_ = new_n3213_ | new_n1292_;
  assign new_n2387_ = new_n2386_ & new_n1494_;
  assign new_n2388_ = new_n2385_ & new_n1493_;
  assign new_n2389_ = new_n2388_ | new_n2387_;
  assign new_n2390_ = new_n3224_ & new_n1371_;
  assign new_n2391_ = new_n3215_ | new_n1372_;
  assign new_n2392_ = new_n2391_ & new_n3207_;
  assign new_n2393_ = new_n2390_ & new_n3205_;
  assign new_n2394_ = new_n2393_ | new_n2392_;
  assign new_n2395_ = new_n3414_ & new_n3434_;
  assign new_n2396_ = new_n3415_ | new_n3431_;
  assign new_n2397_ = new_n3487_ & new_n3680_;
  assign new_n2398_ = new_n3491_ | new_n1398_;
  assign new_n2399_ = new_n2398_ & new_n2396_;
  assign new_n2400_ = new_n2397_ | new_n2395_;
  assign new_n2401_ = new_n2400_ & new_n3421_;
  assign new_n2402_ = new_n2399_ | new_n3428_;
  assign new_n2403_ = new_n3402_ & new_n3493_;
  assign new_n2404_ = new_n3406_ | new_n3489_;
  assign new_n2405_ = new_n3478_ & new_n3490_;
  assign new_n2406_ = new_n3480_ | new_n3492_;
  assign new_n2407_ = new_n2405_ & new_n3389_;
  assign new_n2408_ = new_n2406_ | new_n3396_;
  assign new_n2409_ = new_n2408_ & new_n2404_;
  assign new_n2410_ = new_n2407_ | new_n2403_;
  assign new_n2411_ = new_n2410_ & new_n2402_;
  assign new_n2412_ = new_n2409_ | new_n2401_;
  assign new_n2413_ = new_n3681_ & new_n3501_;
  assign new_n2414_ = new_n1548_ | new_n3499_;
  assign new_n2415_ = new_n1604_ & new_n1590_;
  assign new_n2416_ = new_n1603_ | new_n1589_;
  assign new_n2417_ = new_n2415_ & new_n2414_;
  assign new_n2418_ = new_n2416_ | new_n2413_;
  assign new_n2419_ = new_n2418_ & new_n3454_;
  assign new_n2420_ = new_n2417_ | new_n3460_;
  assign new_n2421_ = new_n2420_ & new_n3503_;
  assign new_n2422_ = new_n2419_ | new_n3505_;
  assign new_n2423_ = new_n3682_ | new_n3497_;
  assign new_n2424_ = new_n2423_ | new_n2074_;
  assign new_n2425_ = new_n3683_ & new_n3686_;
  assign new_n2426_ = new_n2425_ | new_n3690_;
  assign new_n2427_ = new_n2426_ & new_n3691_;
  assign new_n2428_ = new_n3692_ & new_n3686_;
  assign new_n2429_ = new_n2428_ | new_n3693_;
  assign new_n2430_ = new_n2429_ & new_n3694_;
  assign new_n2431_ = new_n3695_ | new_n3248_;
  assign new_n2432_ = new_n3696_ & new_n3697_;
  assign new_n2433_ = new_n3698_ & new_n970_;
  assign new_n2434_ = new_n3701_ & new_n3704_;
  assign new_n2435_ = new_n3372_ & new_n3705_;
  assign new_n2436_ = new_n3708_ & new_n3712_;
  assign new_n2437_ = new_n2436_ | new_n1180_;
  assign new_n2438_ = new_n1288_ & new_n3516_;
  assign new_n2439_ = new_n1290_ & new_n3377_;
  assign new_n2440_ = new_n3671_ & new_n938_;
  assign new_n2441_ = new_n1222_ | new_n3269_;
  assign new_n2442_ = new_n2441_ & new_n1255_;
  assign new_n2443_ = new_n3226_ & new_n1279_;
  assign new_n2444_ = new_n3215_ & new_n3262_;
  assign new_n2445_ = new_n3216_ & new_n3231_;
  assign new_n2446_ = new_n3226_ | new_n3230_;
  assign new_n2447_ = new_n3714_ | new_n3715_;
  assign new_n2448_ = new_n3717_ & new_n3268_;
  assign new_n2449_ = new_n3701_ & new_n3718_;
  assign new_n2450_ = new_n3719_ | new_n3720_;
  assign new_n2451_ = new_n3702_ & new_n3721_;
  assign new_n2452_ = new_n3708_ & new_n3722_;
  assign new_n2453_ = new_n3656_ | new_n3349_;
  assign new_n2454_ = new_n3723_ & new_n3659_;
  assign new_n2455_ = new_n3723_ | new_n3660_;
  assign new_n2456_ = new_n3717_ & new_n3384_;
  assign new_n2457_ = new_n3724_ & new_n3725_;
  assign new_n2458_ = new_n1903_ | new_n3720_;
  assign new_n2459_ = new_n2458_ | new_n3668_;
  assign new_n2460_ = new_n3216_ & new_n3239_;
  assign new_n2461_ = new_n3227_ | new_n3238_;
  assign new_n2462_ = new_n2446_ & new_n3727_;
  assign new_n2463_ = new_n3714_ | new_n3667_;
  assign new_n2464_ = new_n2463_ & new_n2461_;
  assign new_n2465_ = new_n2462_ | new_n3728_;
  assign new_n2466_ = new_n2464_ & new_n3730_;
  assign new_n2467_ = new_n2465_ & new_n3666_;
  assign new_n2468_ = new_n2467_ | new_n2466_;
  assign new_n2469_ = new_n3731_ | new_n3733_;
  assign new_n2470_ = new_n3731_ & new_n3733_;
  assign new_n2471_ = new_n3734_ | new_n3736_;
  assign new_n2472_ = new_n3737_ | new_n3736_;
  assign new_n2473_ = new_n3738_ & new_n3739_;
  assign new_n2474_ = new_n2473_ & new_n3740_;
  assign new_n2475_ = new_n3365_ & new_n3742_;
  assign new_n2476_ = new_n3373_ & new_n3743_;
  assign new_n2477_ = new_n2476_ | new_n2475_;
  assign new_n2478_ = new_n3745_ | new_n3718_;
  assign new_n2479_ = new_n2478_ & new_n3747_;
  assign new_n2480_ = new_n2479_ | new_n3510_;
  assign new_n2481_ = new_n2480_ | new_n2477_;
  assign new_n2482_ = new_n3749_ & new_n1150_;
  assign new_n2483_ = new_n2482_ & new_n3750_;
  assign new_n2484_ = new_n3709_ & new_n1158_;
  assign new_n2485_ = new_n3752_ | new_n3366_;
  assign new_n2486_ = new_n2485_ & new_n3747_;
  assign new_n2487_ = new_n2486_ | new_n2484_;
  assign new_n2488_ = new_n3379_ | new_n3517_;
  assign new_n2489_ = new_n1198_ | new_n3374_;
  assign new_n2490_ = new_n2489_ & new_n2488_;
  assign new_n2491_ = new_n3753_ & new_n3754_;
  assign new_n2492_ = new_n3271_ | new_n917_;
  assign new_n2493_ = new_n2492_ & new_n3748_;
  assign new_n2494_ = new_n3756_ & new_n3742_;
  assign new_n2495_ = new_n2494_ | new_n2493_;
  assign new_n2496_ = new_n3756_ & new_n3381_;
  assign new_n2497_ = new_n3702_ & new_n3712_;
  assign new_n2498_ = new_n3709_ & new_n3383_;
  assign new_n2499_ = new_n2498_ | new_n2497_;
  assign new_n2500_ = new_n2499_ | new_n2496_;
  assign new_n2501_ = new_n3728_ & new_n3730_;
  assign new_n2502_ = new_n3347_ & new_n3348_;
  assign new_n2503_ = new_n2502_ | new_n2501_;
  assign new_n2504_ = new_n3757_ & new_n3758_;
  assign new_n2505_ = new_n3662_ | new_n3229_;
  assign new_n2506_ = new_n3661_ | new_n3237_;
  assign new_n2507_ = new_n3660_ | new_n3346_;
  assign new_n2508_ = new_n2507_ & new_n2287_;
  assign new_n2509_ = new_n2508_ & new_n2506_;
  assign new_n2510_ = new_n2509_ & new_n2505_;
  assign new_n2511_ = new_n3759_ | new_n944_;
  assign new_n2512_ = new_n3414_ & new_n3444_;
  assign new_n2513_ = new_n3761_ & new_n3399_;
  assign new_n2514_ = new_n2513_ | new_n2512_;
  assign new_n2515_ = new_n2514_ & new_n3423_;
  assign new_n2516_ = new_n3437_ | new_n3408_;
  assign new_n2517_ = new_n3479_ | new_n3442_;
  assign new_n2518_ = new_n3477_ | new_n3450_;
  assign new_n2519_ = new_n2518_ & new_n3386_;
  assign new_n2520_ = new_n3763_ | new_n2517_;
  assign new_n2521_ = new_n2520_ & new_n2516_;
  assign new_n2522_ = new_n2521_ | new_n2515_;
  assign new_n2523_ = new_n3713_ | new_n3765_;
  assign new_n2524_ = new_n2457_ | new_n3727_;
  assign new_n2525_ = new_n2524_ & new_n3732_;
  assign new_n2526_ = new_n3766_ | new_n3767_;
  assign new_n2527_ = new_n3766_ & new_n3767_;
  assign new_n2528_ = new_n3481_ & new_n3411_;
  assign new_n2529_ = new_n3440_ & new_n3356_;
  assign new_n2530_ = new_n3436_ & new_n3486_;
  assign new_n2531_ = new_n2530_ | new_n2529_;
  assign new_n2532_ = new_n2531_ & new_n3423_;
  assign new_n2533_ = new_n3763_ & new_n3333_;
  assign new_n2534_ = new_n2533_ | new_n2532_;
  assign new_n2535_ = new_n2534_ | new_n2528_;
  assign new_n2536_ = new_n3364_ & new_n3745_;
  assign new_n2537_ = new_n3768_ & new_n3373_;
  assign new_n2538_ = new_n2537_ | new_n2536_;
  assign new_n2539_ = new_n3769_ & new_n3500_;
  assign new_n2540_ = new_n1600_ | new_n3498_;
  assign new_n2541_ = new_n1584_ & new_n1581_;
  assign new_n2542_ = new_n1583_ | new_n1582_;
  assign new_n2543_ = new_n3771_ & new_n3772_;
  assign new_n2544_ = new_n3774_ | new_n1500_;
  assign new_n2545_ = new_n2544_ & new_n2542_;
  assign new_n2546_ = new_n2543_ | new_n2541_;
  assign new_n2547_ = new_n2545_ & new_n2540_;
  assign new_n2548_ = new_n2546_ | new_n2539_;
  assign new_n2549_ = new_n2548_ & new_n3456_;
  assign new_n2550_ = new_n2547_ | new_n3462_;
  assign new_n2551_ = new_n2550_ & new_n3502_;
  assign new_n2552_ = new_n2549_ | new_n3504_;
  assign new_n2553_ = new_n3775_ | new_n3497_;
  assign new_n2554_ = new_n2553_ | new_n2411_;
  assign new_n2555_ = new_n3748_ & new_n1156_;
  assign new_n2556_ = new_n2555_ | new_n3776_;
  assign new_n2557_ = new_n3703_ & new_n3752_;
  assign new_n2558_ = new_n3710_ & new_n3704_;
  assign new_n2559_ = new_n2558_ | new_n2557_;
  assign new_n2560_ = new_n2559_ | new_n3777_;
  assign new_n2561_ = new_n2560_ | new_n2556_;
  assign new_n2562_ = new_n3778_ & new_n3687_;
  assign new_n2563_ = new_n2562_ | new_n3779_;
  assign new_n2564_ = new_n2563_ & new_n3780_;
  assign new_n2565_ = new_n3781_ & new_n3782_;
  assign new_n2566_ = new_n891_ | new_n3786_;
  assign new_n2567_ = new_n3793_ | new_n3795_;
  assign new_n2568_ = new_n3797_ | new_n3793_;
  assign new_n2569_ = new_n3441_ & new_n3798_;
  assign new_n2570_ = new_n3445_ & new_n3761_;
  assign new_n2571_ = new_n3799_ & new_n3474_;
  assign new_n2572_ = new_n2571_ | new_n2570_;
  assign new_n2573_ = new_n2572_ | new_n2569_;
  assign new_n2574_ = new_n2573_ & new_n3424_;
  assign new_n2575_ = new_n3441_ & new_n3800_;
  assign new_n2576_ = new_n3411_ & new_n3760_;
  assign new_n2577_ = new_n3801_ & new_n3476_;
  assign new_n2578_ = new_n2577_ | new_n2576_;
  assign new_n2579_ = new_n2578_ | new_n2575_;
  assign new_n2580_ = new_n2579_ & new_n3424_;
  assign new_n2581_ = new_n3470_ & new_n3803_;
  assign new_n2582_ = new_n3438_ | new_n3806_;
  assign new_n2583_ = new_n3809_ | new_n3811_;
  assign new_n2584_ = new_n2583_ & new_n2582_;
  assign new_n2585_ = new_n3771_ & new_n947_;
  assign new_n2586_ = new_n2585_ | new_n2584_;
  assign new_n2587_ = new_n2586_ | new_n2581_;
  assign new_n2588_ = new_n2587_ & new_n3456_;
  assign new_n2589_ = new_n3812_ | new_n3778_;
  assign new_n2590_ = new_n3692_ | new_n3683_;
  assign new_n2591_ = new_n2590_ | new_n2589_;
  assign new_n2592_ = new_n2591_ & new_n3360_;
  assign new_n2593_ = new_n3775_ | new_n3682_;
  assign new_n2594_ = new_n3506_ | new_n3494_;
  assign new_n2595_ = new_n2594_ | new_n2593_;
  assign new_n2596_ = new_n2595_ & new_n3358_;
  assign new_n2597_ = new_n3469_ & new_n3813_;
  assign new_n2598_ = new_n3393_ | new_n3806_;
  assign new_n2599_ = new_n3803_ | new_n3809_;
  assign new_n2600_ = new_n2599_ & new_n2598_;
  assign new_n2601_ = new_n3770_ & new_n3811_;
  assign new_n2602_ = new_n2601_ | new_n2600_;
  assign new_n2603_ = new_n2602_ | new_n2597_;
  assign new_n2604_ = new_n2603_ & new_n3455_;
  assign new_n2605_ = new_n2604_ | new_n3814_;
  assign new_n2606_ = new_n3817_ | new_n3821_;
  assign new_n2607_ = new_n3823_ | new_n3824_;
  assign new_n2608_ = new_n3826_ & new_n3786_;
  assign new_n2609_ = new_n3764_ | new_n1560_;
  assign new_n2610_ = new_n3357_ | new_n3408_;
  assign new_n2611_ = new_n2610_ & new_n2609_;
  assign new_n2612_ = new_n3764_ | new_n3445_;
  assign new_n2613_ = new_n3336_ | new_n3407_;
  assign new_n2614_ = new_n2613_ & new_n2612_;
  assign new_n2615_ = new_n3466_ | new_n1394_;
  assign new_n2616_ = new_n3482_ & new_n3810_;
  assign new_n2617_ = new_n3827_ & new_n3805_;
  assign new_n2618_ = new_n2617_ | new_n2616_;
  assign new_n2619_ = new_n3828_ | new_n3774_;
  assign new_n2620_ = new_n2619_ & new_n2618_;
  assign new_n2621_ = new_n2620_ & new_n2615_;
  assign new_n2622_ = new_n2621_ | new_n3462_;
  assign new_n2623_ = new_n2622_ & new_n3829_;
  assign new_n2624_ = new_n3830_ & new_n3832_;
  assign new_n2625_ = new_n2624_ & new_n3834_;
  assign new_n2626_ = new_n3465_ | new_n3827_;
  assign new_n2627_ = new_n3434_ & new_n3810_;
  assign new_n2628_ = new_n3828_ & new_n3807_;
  assign new_n2629_ = new_n2628_ | new_n2627_;
  assign new_n2630_ = new_n1598_ | new_n3773_;
  assign new_n2631_ = new_n2630_ & new_n2629_;
  assign new_n2632_ = new_n2631_ & new_n2626_;
  assign new_n2633_ = new_n2632_ | new_n3461_;
  assign new_n2634_ = new_n2633_ & new_n3829_;
  assign new_n2635_ = new_n3835_ & new_n3832_;
  assign new_n2636_ = new_n2635_ & new_n3837_;
  assign new_n2637_ = new_n3830_ & new_n3687_;
  assign new_n2638_ = new_n2637_ | new_n3834_;
  assign new_n2639_ = new_n3835_ & new_n3689_;
  assign new_n2640_ = new_n2639_ | new_n3837_;
  assign new_n2641_ = new_n3734_ | new_n3839_;
  assign new_n2642_ = new_n3824_ | new_n3839_;
  assign new_n2643_ = new_n2642_ | new_n3817_;
  assign new_n2644_ = new_n2643_ & new_n3840_;
  assign new_n2645_ = new_n3842_ | new_n3826_;
  assign new_n2646_ = new_n3843_ | new_n996_;
  assign new_n2647_ = new_n3812_ & new_n3689_;
  assign new_n2648_ = new_n2647_ | new_n3844_;
  assign new_n2649_ = new_n2648_ & new_n3845_;
  assign new_n2650_ = new_n3846_ & new_n3847_;
  assign new_n2651_ = new_n3848_ | new_n818_;
  assign new_n2652_ = new_n2651_ & new_n3849_;
  assign new_n2653_ = new_n3787_ & new_n3838_;
  assign new_n2654_ = new_n3787_ | new_n3821_;
  assign new_n2655_ = new_n3850_ | new_n3797_;
  assign new_n2656_ = new_n2655_ & new_n3820_;
  assign new_n2657_ = new_n3851_ & new_n3822_;
  assign new_n2658_ = new_n3852_ | new_n3788_;
  assign new_n2659_ = new_n866_ & new_n3788_;
  assign new_n2660_ = new_n3854_ | new_n3794_;
  assign new_n2661_ = new_n3854_ | new_n3848_;
  assign new_n2662_ = new_n3857_ | new_n3859_;
  assign new_n2663_ = new_n3840_ | new_n3860_;
  assign new_n2664_ = new_n3861_ & new_n3863_;
  assign new_n2665_ = new_n3857_ | new_n858_;
  assign new_n2666_ = new_n3864_ & new_n3865_;
  assign new_n2667_ = new_n3866_ | new_n3790_;
  assign new_n2668_ = new_n3863_ | new_n3816_;
  assign new_n2669_ = new_n2668_ & new_n2667_;
  assign new_n2670_ = new_n872_ & new_n3818_;
  assign new_n2671_ = new_n3859_ & new_n3790_;
  assign new_n2672_ = new_n2671_ | new_n2670_;
  assign new_n2673_ = new_n3858_ | new_n860_;
  assign new_n2674_ = new_n2673_ & new_n2672_;
  assign new_n2675_ = new_n3867_ & new_n3791_;
  assign new_n2676_ = new_n3868_ & new_n3818_;
  assign new_n2677_ = new_n2676_ | new_n2675_;
  assign new_n2678_ = new_n3842_ & new_n3869_;
  assign new_n2679_ = new_n2678_ | new_n2677_;
  assign G3519 = new_n1617_;
  assign G3520 = new_n1090_;
  assign G3521 = new_n1642_;
  assign G3522 = new_n1681_;
  assign G3523 = new_n1700_;
  assign G3524 = new_n1701_;
  assign G3525 = new_n1703_;
  assign G3526 = new_n1095_;
  assign G3527 = new_n1706_;
  assign G3528 = new_n3146_;
  assign G3529 = new_n3134_;
  assign G3530 = new_n1748_;
  assign G3531 = new_n3140_;
  assign G3532 = new_n3144_;
  assign G3533 = new_n3138_;
  assign G3534 = new_n1247_;
  assign G3535 = new_n1249_;
  assign G3536 = new_n3132_;
  assign G3537 = new_n3155_;
  assign G3538 = ~new_n1786_;
  assign G3539 = new_n1823_;
  assign G3540 = new_n1832_;
  assign n4070_li003_li003 = new_n3192_;
  assign n4094_li011_li011 = new_n3310_;
  assign n4142_li027_li027 = new_n3180_;
  assign n4154_li031_li031 = new_n3586_;
  assign n4166_li035_li035 = new_n1081_;
  assign n4178_li039_li039 = new_n1083_;
  assign n4190_li043_li043 = new_n3592_;
  assign n4202_li047_li047 = new_n3588_;
  assign n4214_li051_li051 = new_n3593_;
  assign n4226_li055_li055 = new_n3591_;
  assign n4229_li056_li056 = new_n823_;
  assign n4232_li057_li057 = new_n915_;
  assign n4241_li060_li060 = new_n825_;
  assign n4244_li061_li061 = new_n919_;
  assign n4253_li064_li064 = new_n827_;
  assign n4256_li065_li065 = new_n923_;
  assign n4265_li068_li068 = new_n829_;
  assign n4268_li069_li069 = new_n927_;
  assign n4277_li072_li072 = new_n831_;
  assign n4280_li073_li073 = new_n931_;
  assign n4289_li076_li076 = new_n833_;
  assign n4292_li077_li077 = new_n935_;
  assign n4301_li080_li080 = new_n835_;
  assign n4313_li084_li084 = new_n837_;
  assign n4373_li104_li104 = new_n847_;
  assign n4382_li107_li107 = new_n1129_;
  assign n4385_li108_li108 = new_n849_;
  assign n4397_li112_li112 = new_n851_;
  assign n4418_li119_li119 = new_n1091_;
  assign n4430_li123_li123 = new_n1085_;
  assign n4442_li127_li127 = new_n1069_;
  assign n4454_li131_li131 = new_n1047_;
  assign n4466_li135_li135 = new_n1049_;
  assign n4478_li139_li139 = new_n1059_;
  assign n4490_li143_li143 = new_n1071_;
  assign n4502_li147_li147 = new_n1093_;
  assign n4553_li164_li164 = new_n877_;
  assign n4556_li165_li165 = new_n967_;
  assign n4565_li168_li168 = new_n879_;
  assign n4568_li169_li169 = new_n971_;
  assign n4577_li172_li172 = new_n881_;
  assign n4580_li173_li173 = new_n975_;
  assign n4589_li176_li176 = new_n883_;
  assign n4592_li177_li177 = new_n979_;
  assign n4601_li180_li180 = new_n885_;
  assign n4604_li181_li181 = new_n983_;
  assign n4607_li182_li182 = new_n985_;
  assign n4613_li184_li184 = new_n887_;
  assign n4616_li185_li185 = new_n989_;
  assign n4622_li187_li187 = new_n3288_;
  assign n4625_li188_li188 = new_n889_;
  assign n4634_li191_li191 = new_n1137_;
  assign n4649_li196_li196 = new_n893_;
  assign n4652_li197_li197 = new_n999_;
  assign n4655_li198_li198 = new_n1001_;
  assign n4658_li199_li199 = new_n1003_;
  assign n2071_i2 = new_n3311_;
  assign n2080_i2 = new_n1065_;
  assign n2137_i2 = new_n1079_;
  assign n2368_i2 = new_n1113_;
  assign n2383_i2 = new_n1117_;
  assign n2405_i2 = new_n1123_;
  assign n2471_i2 = new_n3187_;
  assign n2617_i2 = new_n1145_;
  assign n2765_i2 = new_n1215_;
  assign n2775_i2 = new_n1217_;
  assign n2829_i2 = new_n3549_;
  assign n2579_i2 = new_n1141_;
  assign n2580_i2 = new_n3248_;
  assign n2618_i2 = new_n3695_;
  assign n2619_i2 = new_n3509_;
  assign n2620_i2 = new_n1151_;
  assign n2621_i2 = new_n3697_;
  assign n2622_i2 = new_n3672_;
  assign n2623_i2 = new_n3369_;
  assign n2624_i2 = new_n3698_;
  assign n2625_i2 = new_n1161_;
  assign n2626_i2 = new_n1163_;
  assign n2627_i2 = new_n3751_;
  assign n3029_i2 = new_n1341_;
  assign n3035_i2 = new_n1345_;
  assign n2643_i2 = new_n3749_;
  assign n2644_i2 = new_n1171_;
  assign n2645_i2 = new_n1173_;
  assign n2640_i2 = new_n1167_;
  assign n2658_i2 = new_n1175_;
  assign n2659_i2 = new_n1177_;
  assign n2674_i2 = new_n1181_;
  assign n2675_i2 = new_n1183_;
  assign n2676_i2 = new_n3705_;
  assign n3119_i2 = new_n3285_;
  assign n3153_i2 = new_n3185_;
  assign n2681_i2 = new_n1187_;
  assign n2729_i2 = new_n3517_;
  assign n2730_i2 = new_n3379_;
  assign n2731_i2 = new_n1199_;
  assign n698_i2 = ~new_n3563_;
  assign n677_i2 = ~new_n3564_;
  assign n2757_i2 = new_n1207_;
  assign n2758_i2 = new_n1209_;
  assign n1000_i2 = new_n3534_;
  assign n1160_i2 = new_n3326_;
  assign n1153_i2 = new_n3292_;
  assign n2793_i2 = new_n3696_;
  assign n2794_i2 = new_n3670_;
  assign n2795_i2 = new_n1223_;
  assign n1001_i2 = new_n3194_;
  assign n2859_i2 = new_n1251_;
  assign n744_i2 = new_n3562_;
  assign n2908_i2 = new_n1275_;
  assign n2926_i2 = new_n1277_;
  assign n2928_i2 = new_n1281_;
  assign n2966_i2 = new_n3741_;
  assign n2967_i2 = new_n3380_;
  assign n2947_i2 = new_n1283_;
  assign n1010_i2 = new_n3322_;
  assign n2976_i2 = new_n3264_;
  assign n3069_i2 = new_n1369_;
  assign n3028_i2 = new_n1339_;
  assign n3081_i2 = new_n3263_;
  assign n3082_i2 = new_n1377_;
  assign n3142_i2 = new_n1453_;
  assign n3214_i2 = new_n3227_;
  assign n2992_i2 = new_n3450_;
  assign n2993_i2 = new_n3476_;
  assign n870_i2 = new_n3228_;
  assign n3086_i2 = new_n3447_;
  assign n3087_i2 = new_n3807_;
  assign n3088_i2 = new_n3464_;
  assign n3089_i2 = new_n3393_;
  assign n3090_i2 = new_n3431_;
  assign n3091_i2 = new_n3484_;
  assign n3092_i2 = new_n3490_;
  assign n3093_i2 = new_n1393_;
  assign n3094_i2 = new_n1395_;
  assign n3095_i2 = new_n3680_;
  assign n3136_i2 = new_n1449_;
  assign n3170_i2 = new_n3463_;
  assign n3171_i2 = new_n3772_;
  assign n3172_i2 = new_n1501_;
  assign n3179_i2 = new_n1505_;
  assign n3180_i2 = new_n1507_;
  assign n3193_i2 = new_n1527_;
  assign n3211_i2 = new_n1545_;
  assign n3212_i2 = new_n3681_;
  assign n3213_i2 = new_n1549_;
  assign n3219_i2 = new_n1557_;
  assign n1125_i2 = new_n3267_;
  assign n1081_i2 = new_n3265_;
  assign n1139_i2 = new_n3726_;
  assign n3245_i2 = new_n3333_;
  assign n3246_i2 = new_n3438_;
  assign n3247_i2 = new_n3813_;
  assign lo074_buf_i2 = new_n3270_;
  assign lo078_buf_i2 = new_n3744_;
  assign lo186_buf_i2 = new_n3725_;
  assign lo118_buf_i2 = new_n3802_;
  assign lo146_buf_i2 = new_n3769_;
  assign n1038_i2 = ~new_n3703_;
  assign n1044_i2 = new_n3710_;
  assign n980_i2 = new_n3272_;
  assign n1145_i2 = new_n3724_;
  assign lo026_buf_i2 = new_n3357_;
  assign lo030_buf_i2 = new_n3336_;
  assign lo090_buf_i2 = new_n3361_;
  assign lo094_buf_i2 = new_n3359_;
  assign lo098_buf_i2 = new_n3363_;
  assign lo102_buf_i2 = new_n3362_;
  assign lo066_buf_i2 = new_n3711_;
  assign lo070_buf_i2 = new_n3382_;
  assign n1202_i2 = ~new_n3743_;
  assign n1003_i2 = new_n1905_;
  assign n1031_i2 = new_n3755_;
  assign n1034_i2 = new_n3367_;
  assign n1040_i2 = new_n3370_;
  assign n1046_i2 = new_n3518_;
  assign n1380_i2 = new_n3678_;
  assign n1425_i2 = new_n3676_;
  assign n697_i2 = new_n3446_;
  assign n1143_i2 = new_n3729_;
  assign n673_i2 = new_n3385_;
  assign n789_i2 = new_n3831_;
  assign n786_i2 = new_n3688_;
  assign n1047_i2 = ~new_n3777_;
  assign n1036_i2 = new_n3508_;
  assign n1307_i2 = ~new_n3739_;
  assign n1035_i2 = ~new_n3776_;
  assign n1297_i2 = ~new_n3738_;
  assign n1099_i2 = new_n3768_;
  assign n1128_i2 = new_n3765_;
  assign n674_i2 = new_n3799_;
  assign n826_i2 = new_n3690_;
  assign n853_i2 = new_n3693_;
  assign n951_i2 = new_n3801_;
  assign n700_i2 = new_n3654_;
  assign n884_i2 = new_n3814_;
  assign lo082_buf_i2 = new_n3798_;
  assign lo086_buf_i2 = new_n3800_;
  assign n801_i2 = new_n3779_;
  assign n840_i2 = ~new_n3691_;
  assign n866_i2 = ~new_n3694_;
  assign lo002_buf_i2 = new_n3735_;
  assign lo010_buf_i2 = new_n3822_;
  assign lo166_buf_i2 = new_n3722_;
  assign lo170_buf_i2 = new_n3721_;
  assign n1426_i2 = ~new_n2096_;
  assign n1082_i2 = ~new_n2097_;
  assign n1310_i2 = new_n3740_;
  assign n1015_i2 = ~new_n2100_;
  assign n1206_i2 = ~new_n3750_;
  assign n1262_i2 = new_n3754_;
  assign n1456_i2 = new_n2103_;
  assign n1244_i2 = new_n2135_;
  assign n1280_i2 = new_n2136_;
  assign n1290_i2 = new_n2137_;
  assign n1012_i2 = new_n2139_;
  assign n1074_i2 = ~new_n2180_;
  assign n1112_i2 = ~new_n2207_;
  assign n1212_i2 = new_n2235_;
  assign n1454_i2 = new_n2266_;
  assign n1182_i2 = ~new_n2275_;
  assign n1220_i2 = ~new_n3758_;
  assign n701_i2 = new_n3759_;
  assign n973_i2 = ~new_n3716_;
  assign n1282_i2 = new_n2295_;
  assign n1144_i2 = ~new_n3715_;
  assign n1278_i2 = new_n2322_;
  assign n1459_i2 = new_n2325_;
  assign n1324_i2 = new_n2351_;
  assign n1288_i2 = new_n2354_;
  assign n1271_i2 = new_n3753_;
  assign n1132_i2 = new_n2365_;
  assign n1231_i2 = new_n2382_;
  assign n1462_i2 = new_n2383_;
  assign n1482_i2 = new_n2384_;
  assign n994_i2 = ~new_n3757_;
  assign n998_i2 = ~new_n3719_;
  assign lo106_buf_i2 = new_n943_;
  assign n769_i2 = new_n3844_;
  assign n814_i2 = ~new_n3780_;
  assign n841_i2 = new_n3782_;
  assign n867_i2 = new_n3781_;
  assign lo006_buf_i2 = new_n797_;
  assign lo014_buf_i2 = new_n3791_;
  assign lo022_buf_i2 = new_n3737_;
  assign lo042_buf_i2 = new_n3795_;
  assign lo046_buf_i2 = new_n3794_;
  assign lo050_buf_i2 = new_n3796_;
  assign lo054_buf_i2 = new_n3868_;
  assign lo130_buf_i2 = new_n3867_;
  assign lo134_buf_i2 = new_n3869_;
  assign lo154_buf_i2 = new_n871_;
  assign lo174_buf_i2 = new_n977_;
  assign lo178_buf_i2 = new_n981_;
  assign n1007_i2 = new_n2431_;
  assign n1294_i2 = new_n2432_;
  assign n1084_i2 = new_n2433_;
  assign n1399_i2 = ~new_n2434_;
  assign n1311_i2 = new_n2435_;
  assign n1392_i2 = ~new_n2437_;
  assign n1102_i2 = new_n2438_;
  assign n1041_i2 = new_n2439_;
  assign n1298_i2 = new_n2440_;
  assign n738_i2 = new_n2442_;
  assign n1214_i2 = new_n2443_;
  assign n1222_i2 = new_n2444_;
  assign n1155_i2 = ~new_n2447_;
  assign n1147_i2 = new_n2448_;
  assign n1393_i2 = new_n2449_;
  assign n999_i2 = ~new_n2450_;
  assign n1306_i2 = new_n2451_;
  assign n1312_i2 = new_n2452_;
  assign n1382_i2 = ~new_n2454_;
  assign n1383_i2 = ~new_n2455_;
  assign n1152_i2 = ~new_n2456_;
  assign n1334_i2 = ~new_n2469_;
  assign n1335_i2 = new_n2470_;
  assign n695_i2 = ~new_n3823_;
  assign n773_i2 = new_n3841_;
  assign lo190_buf_i2 = new_n995_;
  assign n1368_i2 = new_n2474_;
  assign n1362_i2 = ~new_n2481_;
  assign n1406_i2 = new_n2483_;
  assign n1403_i2 = ~new_n2487_;
  assign n741_i2 = new_n2490_;
  assign n1407_i2 = new_n2491_;
  assign n1395_i2 = new_n2495_;
  assign n1359_i2 = new_n2500_;
  assign n1159_i2 = new_n2503_;
  assign n1221_i2 = ~new_n2504_;
  assign n987_i2 = ~new_n2510_;
  assign n989_i2 = ~new_n3843_;
  assign n881_i2 = new_n3833_;
  assign n1340_i2 = new_n2526_;
  assign n1341_i2 = new_n2527_;
  assign n906_i2 = new_n3836_;
  assign n1388_i2 = new_n2538_;
  assign n791_i2 = ~new_n3845_;
  assign n1372_i2 = ~new_n2561_;
  assign n815_i2 = new_n3847_;
  assign n868_i2 = new_n3846_;
  assign lo018_buf_i2 = new_n3825_;
  assign lo138_buf_i2 = new_n3862_;
  assign lo158_buf_i2 = new_n3866_;
  assign n780_i2 = new_n3858_;
  assign n728_i2 = new_n3850_;
  assign n676_i2 = new_n3849_;
  assign n929_i2 = new_n2574_;
  assign n955_i2 = new_n2580_;
  assign n938_i2 = new_n2588_;
  assign n1117_i2 = new_n2592_;
  assign n1121_i2 = new_n2596_;
  assign n965_i2 = new_n2605_;
  assign n752_i2 = ~new_n3855_;
  assign n753_i2 = n752_i2;
  assign n760_i2 = ~new_n3865_;
  assign n770_i2 = new_n3860_;
  assign n923_i2 = new_n2611_;
  assign n947_i2 = new_n2614_;
  assign n897_i2 = new_n2625_;
  assign n919_i2 = new_n2636_;
  assign n895_i2 = new_n2638_;
  assign n917_i2 = new_n2640_;
  assign n751_i2 = ~new_n3864_;
  assign n774_i2 = new_n3861_;
  assign lo126_buf_i2 = new_n857_;
  assign lo142_buf_i2 = new_n865_;
  assign lo162_buf_i2 = new_n3852_;
  assign n990_i2 = ~new_n2646_;
  assign n792_i2 = new_n2649_;
  assign n869_i2 = new_n2650_;
  assign n848_i2 = new_n3851_;
  assign lo024_buf_i2 = new_n807_;
  assign lo028_buf_i2 = new_n809_;
  assign lo088_buf_i2 = new_n839_;
  assign lo092_buf_i2 = new_n841_;
  assign lo096_buf_i2 = new_n843_;
  assign lo100_buf_i2 = new_n845_;
  assign n763_i2 = new_n2653_;
  assign n754_i2 = new_n3870_;
  assign n755_i2 = n754_i2;
  assign n822_i2 = new_n2656_;
  assign n849_i2 = new_n2657_;
  assign n777_i2 = new_n2658_;
  assign n778_i2 = new_n2659_;
  assign n820_i2 = ~new_n2660_;
  assign n846_i2 = ~new_n2661_;
  assign n806_i2 = ~new_n2662_;
  assign n771_i2 = ~new_n2663_;
  assign n854_i2 = new_n2664_;
  assign n828_i2 = ~new_n2665_;
  assign lo117_buf_i2 = new_n853_;
  assign lo145_buf_i2 = new_n867_;
  assign n762_i2 = ~new_n2666_;
  assign n805_i2 = new_n2669_;
  assign n859_i2 = ~new_n2674_;
  assign n833_i2 = new_n2679_;
  assign lo034_buf_i2 = new_n811_;
  assign lo038_buf_i2 = new_n813_;
  assign lo122_buf_i2 = new_n855_;
  assign lo150_buf_i2 = new_n869_;
  assign new_n3063_ = new_n906_;
  assign new_n3064_ = new_n898_;
  assign new_n3065_ = new_n896_;
  assign new_n3066_ = new_n960_;
  assign new_n3067_ = new_n3066_;
  assign new_n3068_ = new_n3066_;
  assign new_n3069_ = new_n907_;
  assign new_n3070_ = new_n956_;
  assign new_n3071_ = new_n3070_;
  assign new_n3072_ = new_n952_;
  assign new_n3073_ = new_n3072_;
  assign new_n3074_ = new_n899_;
  assign new_n3075_ = new_n958_;
  assign new_n3076_ = new_n3075_;
  assign new_n3077_ = new_n966_;
  assign new_n3078_ = new_n3077_;
  assign new_n3079_ = new_n913_;
  assign new_n3080_ = new_n3079_;
  assign new_n3081_ = new_n954_;
  assign new_n3082_ = new_n3081_;
  assign new_n3083_ = new_n962_;
  assign new_n3084_ = new_n3083_;
  assign new_n3085_ = new_n3083_;
  assign new_n3086_ = new_n909_;
  assign new_n3087_ = new_n964_;
  assign new_n3088_ = new_n3087_;
  assign new_n3089_ = new_n3087_;
  assign new_n3090_ = new_n911_;
  assign new_n3091_ = new_n3090_;
  assign new_n3092_ = new_n1636_;
  assign new_n3093_ = new_n963_;
  assign new_n3094_ = new_n965_;
  assign new_n3095_ = new_n959_;
  assign new_n3096_ = new_n961_;
  assign new_n3097_ = new_n1653_;
  assign new_n3098_ = new_n1648_;
  assign new_n3099_ = new_n1654_;
  assign new_n3100_ = new_n1647_;
  assign new_n3101_ = new_n955_;
  assign new_n3102_ = new_n957_;
  assign new_n3103_ = new_n951_;
  assign new_n3104_ = new_n953_;
  assign new_n3105_ = new_n1672_;
  assign new_n3106_ = new_n1665_;
  assign new_n3107_ = new_n1671_;
  assign new_n3108_ = new_n1666_;
  assign new_n3109_ = new_n914_;
  assign new_n3110_ = new_n3109_;
  assign new_n3111_ = new_n912_;
  assign new_n3112_ = new_n1690_;
  assign new_n3113_ = new_n1684_;
  assign new_n3114_ = new_n1691_;
  assign new_n3115_ = new_n1685_;
  assign new_n3116_ = new_n1053_;
  assign new_n3117_ = new_n1108_;
  assign new_n3118_ = new_n3117_;
  assign new_n3119_ = new_n1126_;
  assign new_n3120_ = new_n1125_;
  assign new_n3121_ = new_n1720_;
  assign new_n3122_ = new_n1075_;
  assign new_n3123_ = new_n1719_;
  assign new_n3124_ = new_n1076_;
  assign new_n3125_ = new_n1099_;
  assign new_n3126_ = new_n1097_;
  assign new_n3127_ = new_n1100_;
  assign new_n3128_ = new_n1098_;
  assign new_n3129_ = new_n1107_;
  assign new_n3130_ = new_n1771_;
  assign new_n3131_ = new_n1717_;
  assign new_n3132_ = new_n1772_;
  assign new_n3133_ = new_n3132_;
  assign new_n3134_ = new_n1718_;
  assign new_n3135_ = new_n3134_;
  assign new_n3136_ = new_n1765_;
  assign new_n3137_ = new_n1753_;
  assign new_n3138_ = new_n1766_;
  assign new_n3139_ = new_n3138_;
  assign new_n3140_ = new_n1754_;
  assign new_n3141_ = new_n3140_;
  assign new_n3142_ = new_n1759_;
  assign new_n3143_ = new_n1711_;
  assign new_n3144_ = new_n1760_;
  assign new_n3145_ = new_n3144_;
  assign new_n3146_ = new_n1712_;
  assign new_n3147_ = new_n3146_;
  assign new_n3148_ = new_n1778_;
  assign new_n3149_ = new_n1776_;
  assign new_n3150_ = new_n1774_;
  assign new_n3151_ = new_n1361_;
  assign new_n3152_ = new_n3151_;
  assign new_n3153_ = new_n945_;
  assign new_n3154_ = new_n1783_;
  assign new_n3155_ = new_n1781_;
  assign new_n3156_ = new_n1794_;
  assign new_n3157_ = new_n1789_;
  assign new_n3158_ = new_n1793_;
  assign new_n3159_ = new_n1790_;
  assign new_n3160_ = new_n1806_;
  assign new_n3161_ = new_n3160_;
  assign new_n3162_ = new_n3160_;
  assign new_n3163_ = new_n1005_;
  assign new_n3164_ = new_n1805_;
  assign new_n3165_ = new_n3164_;
  assign new_n3166_ = new_n3164_;
  assign new_n3167_ = new_n1006_;
  assign new_n3168_ = new_n1813_;
  assign new_n3169_ = new_n1803_;
  assign new_n3170_ = new_n3169_;
  assign new_n3171_ = new_n3169_;
  assign new_n3172_ = new_n1814_;
  assign new_n3173_ = new_n1804_;
  assign new_n3174_ = new_n3173_;
  assign new_n3175_ = new_n3173_;
  assign new_n3176_ = new_n1800_;
  assign new_n3177_ = new_n1799_;
  assign new_n3178_ = new_n1101_;
  assign new_n3179_ = new_n3178_;
  assign new_n3180_ = new_n3178_;
  assign new_n3181_ = new_n1040_;
  assign new_n3182_ = new_n1366_;
  assign new_n3183_ = new_n3182_;
  assign new_n3184_ = new_n1365_;
  assign new_n3185_ = new_n1475_;
  assign new_n3186_ = new_n1132_;
  assign new_n3187_ = new_n1131_;
  assign new_n3188_ = new_n3187_;
  assign new_n3189_ = new_n1037_;
  assign new_n3190_ = new_n1403_;
  assign new_n3191_ = new_n1038_;
  assign new_n3192_ = new_n1029_;
  assign new_n3193_ = new_n1848_;
  assign new_n3194_ = new_n1841_;
  assign new_n3195_ = new_n3194_;
  assign new_n3196_ = new_n1849_;
  assign new_n3197_ = new_n3196_;
  assign new_n3198_ = new_n3197_;
  assign new_n3199_ = new_n3197_;
  assign new_n3200_ = new_n3196_;
  assign new_n3201_ = new_n1842_;
  assign new_n3202_ = new_n3201_;
  assign new_n3203_ = new_n3201_;
  assign new_n3204_ = new_n1555_;
  assign new_n3205_ = new_n1553_;
  assign new_n3206_ = new_n1556_;
  assign new_n3207_ = new_n1554_;
  assign new_n3208_ = new_n1552_;
  assign new_n3209_ = new_n3208_;
  assign new_n3210_ = new_n3209_;
  assign new_n3211_ = new_n3210_;
  assign new_n3212_ = new_n3210_;
  assign new_n3213_ = new_n3209_;
  assign new_n3214_ = new_n3208_;
  assign new_n3215_ = new_n3214_;
  assign new_n3216_ = new_n3214_;
  assign new_n3217_ = new_n1551_;
  assign new_n3218_ = new_n3217_;
  assign new_n3219_ = new_n3218_;
  assign new_n3220_ = new_n3219_;
  assign new_n3221_ = new_n3219_;
  assign new_n3222_ = new_n3218_;
  assign new_n3223_ = new_n3222_;
  assign new_n3224_ = new_n3222_;
  assign new_n3225_ = new_n3217_;
  assign new_n3226_ = new_n3225_;
  assign new_n3227_ = new_n3225_;
  assign new_n3228_ = new_n1852_;
  assign new_n3229_ = new_n1534_;
  assign new_n3230_ = new_n3229_;
  assign new_n3231_ = new_n1533_;
  assign new_n3232_ = new_n1865_;
  assign new_n3233_ = new_n1863_;
  assign new_n3234_ = new_n3233_;
  assign new_n3235_ = new_n1864_;
  assign new_n3236_ = new_n1862_;
  assign new_n3237_ = new_n1536_;
  assign new_n3238_ = new_n3237_;
  assign new_n3239_ = new_n1535_;
  assign new_n3240_ = new_n1875_;
  assign new_n3241_ = new_n1873_;
  assign new_n3242_ = new_n3241_;
  assign new_n3243_ = new_n1874_;
  assign new_n3244_ = new_n1872_;
  assign new_n3245_ = new_n1143_;
  assign new_n3246_ = new_n3245_;
  assign new_n3247_ = new_n3246_;
  assign new_n3248_ = new_n3245_;
  assign new_n3249_ = new_n1144_;
  assign new_n3250_ = new_n3249_;
  assign new_n3251_ = new_n1884_;
  assign new_n3252_ = new_n3251_;
  assign new_n3253_ = new_n3252_;
  assign new_n3254_ = new_n3252_;
  assign new_n3255_ = new_n3251_;
  assign new_n3256_ = new_n1230_;
  assign new_n3257_ = new_n1882_;
  assign new_n3258_ = new_n3257_;
  assign new_n3259_ = new_n3257_;
  assign new_n3260_ = new_n1229_;
  assign new_n3261_ = new_n1490_;
  assign new_n3262_ = new_n1373_;
  assign new_n3263_ = new_n1375_;
  assign new_n3264_ = new_n1295_;
  assign new_n3265_ = new_n1870_;
  assign new_n3266_ = new_n3265_;
  assign new_n3267_ = new_n1860_;
  assign new_n3268_ = new_n3267_;
  assign new_n3269_ = new_n1220_;
  assign new_n3270_ = new_n933_;
  assign new_n3271_ = new_n3270_;
  assign new_n3272_ = new_n1901_;
  assign new_n3273_ = new_n1908_;
  assign new_n3274_ = new_n1883_;
  assign new_n3275_ = new_n1907_;
  assign new_n3276_ = new_n1909_;
  assign new_n3277_ = new_n1885_;
  assign new_n3278_ = new_n3277_;
  assign new_n3279_ = new_n3277_;
  assign new_n3280_ = new_n1910_;
  assign new_n3281_ = new_n1913_;
  assign new_n3282_ = new_n1914_;
  assign new_n3283_ = new_n1446_;
  assign new_n3284_ = new_n1445_;
  assign new_n3285_ = new_n1429_;
  assign new_n3286_ = new_n1205_;
  assign new_n3287_ = new_n3286_;
  assign new_n3288_ = new_n3286_;
  assign new_n3289_ = new_n1206_;
  assign new_n3290_ = new_n3289_;
  assign new_n3291_ = new_n3289_;
  assign new_n3292_ = new_n1839_;
  assign new_n3293_ = new_n1928_;
  assign new_n3294_ = new_n1924_;
  assign new_n3295_ = new_n3294_;
  assign new_n3296_ = new_n1927_;
  assign new_n3297_ = new_n1923_;
  assign new_n3298_ = new_n1930_;
  assign new_n3299_ = new_n1922_;
  assign new_n3300_ = new_n3299_;
  assign new_n3301_ = new_n1036_;
  assign new_n3302_ = new_n3301_;
  assign new_n3303_ = new_n3302_;
  assign new_n3304_ = new_n3302_;
  assign new_n3305_ = new_n3301_;
  assign new_n3306_ = new_n3305_;
  assign new_n3307_ = new_n1935_;
  assign new_n3308_ = new_n3307_;
  assign new_n3309_ = new_n3307_;
  assign new_n3310_ = new_n1031_;
  assign new_n3311_ = new_n1063_;
  assign new_n3312_ = new_n1939_;
  assign new_n3313_ = new_n3312_;
  assign new_n3314_ = new_n3313_;
  assign new_n3315_ = new_n3313_;
  assign new_n3316_ = new_n3312_;
  assign new_n3317_ = new_n3316_;
  assign new_n3318_ = new_n1850_;
  assign new_n3319_ = new_n3318_;
  assign new_n3320_ = new_n3319_;
  assign new_n3321_ = new_n3319_;
  assign new_n3322_ = new_n3318_;
  assign new_n3323_ = new_n3322_;
  assign new_n3324_ = new_n1951_;
  assign new_n3325_ = new_n3324_;
  assign new_n3326_ = new_n1838_;
  assign new_n3327_ = new_n3326_;
  assign new_n3328_ = new_n1950_;
  assign new_n3329_ = new_n1837_;
  assign new_n3330_ = new_n1609_;
  assign new_n3331_ = new_n3330_;
  assign new_n3332_ = new_n3331_;
  assign new_n3333_ = new_n3330_;
  assign new_n3334_ = new_n1561_;
  assign new_n3335_ = new_n3334_;
  assign new_n3336_ = new_n3334_;
  assign new_n3337_ = new_n1520_;
  assign new_n3338_ = new_n1519_;
  assign new_n3339_ = new_n1260_;
  assign new_n3340_ = new_n1981_;
  assign new_n3341_ = new_n3340_;
  assign new_n3342_ = new_n1982_;
  assign new_n3343_ = new_n3342_;
  assign new_n3344_ = new_n1257_;
  assign new_n3345_ = new_n1258_;
  assign new_n3346_ = new_n1988_;
  assign new_n3347_ = new_n1987_;
  assign new_n3348_ = new_n1478_;
  assign new_n3349_ = new_n3348_;
  assign new_n3350_ = new_n1992_;
  assign new_n3351_ = new_n1990_;
  assign new_n3352_ = new_n3351_;
  assign new_n3353_ = new_n1991_;
  assign new_n3354_ = new_n1989_;
  assign new_n3355_ = new_n1559_;
  assign new_n3356_ = new_n3355_;
  assign new_n3357_ = new_n3355_;
  assign new_n3358_ = new_n1566_;
  assign new_n3359_ = new_n1565_;
  assign new_n3360_ = new_n3359_;
  assign new_n3361_ = new_n1563_;
  assign new_n3362_ = new_n1569_;
  assign new_n3363_ = new_n1567_;
  assign new_n3364_ = new_n1920_;
  assign new_n3365_ = new_n3364_;
  assign new_n3366_ = new_n1154_;
  assign new_n3367_ = new_n1915_;
  assign new_n3368_ = new_n3367_;
  assign new_n3369_ = new_n1157_;
  assign new_n3370_ = new_n1917_;
  assign new_n3371_ = new_n1916_;
  assign new_n3372_ = new_n3371_;
  assign new_n3373_ = new_n3371_;
  assign new_n3374_ = new_n1196_;
  assign new_n3375_ = new_n1911_;
  assign new_n3376_ = new_n1197_;
  assign new_n3377_ = new_n3376_;
  assign new_n3378_ = new_n3377_;
  assign new_n3379_ = new_n3376_;
  assign new_n3380_ = new_n1289_;
  assign new_n3381_ = new_n3380_;
  assign new_n3382_ = new_n929_;
  assign new_n3383_ = new_n3382_;
  assign new_n3384_ = new_n1906_;
  assign new_n3385_ = new_n1999_;
  assign new_n3386_ = new_n1602_;
  assign new_n3387_ = new_n2012_;
  assign new_n3388_ = new_n3387_;
  assign new_n3389_ = new_n3387_;
  assign new_n3390_ = new_n1385_;
  assign new_n3391_ = new_n3390_;
  assign new_n3392_ = new_n3391_;
  assign new_n3393_ = new_n3390_;
  assign new_n3394_ = new_n2011_;
  assign new_n3395_ = new_n3394_;
  assign new_n3396_ = new_n3394_;
  assign new_n3397_ = new_n1386_;
  assign new_n3398_ = new_n3397_;
  assign new_n3399_ = new_n3397_;
  assign new_n3400_ = new_n1526_;
  assign new_n3401_ = new_n3400_;
  assign new_n3402_ = new_n3400_;
  assign new_n3403_ = new_n1525_;
  assign new_n3404_ = new_n3403_;
  assign new_n3405_ = new_n3404_;
  assign new_n3406_ = new_n3404_;
  assign new_n3407_ = new_n3403_;
  assign new_n3408_ = new_n3407_;
  assign new_n3409_ = new_n1610_;
  assign new_n3410_ = new_n3409_;
  assign new_n3411_ = new_n3409_;
  assign new_n3412_ = new_n1574_;
  assign new_n3413_ = new_n3412_;
  assign new_n3414_ = new_n3412_;
  assign new_n3415_ = new_n1573_;
  assign new_n3416_ = new_n3415_;
  assign new_n3417_ = new_n1541_;
  assign new_n3418_ = new_n3417_;
  assign new_n3419_ = new_n3418_;
  assign new_n3420_ = new_n3419_;
  assign new_n3421_ = new_n3418_;
  assign new_n3422_ = new_n3417_;
  assign new_n3423_ = new_n3422_;
  assign new_n3424_ = new_n3422_;
  assign new_n3425_ = new_n1542_;
  assign new_n3426_ = new_n3425_;
  assign new_n3427_ = new_n3426_;
  assign new_n3428_ = new_n3425_;
  assign new_n3429_ = new_n1387_;
  assign new_n3430_ = new_n3429_;
  assign new_n3431_ = new_n3429_;
  assign new_n3432_ = new_n1388_;
  assign new_n3433_ = new_n3432_;
  assign new_n3434_ = new_n3432_;
  assign new_n3435_ = new_n1611_;
  assign new_n3436_ = new_n3435_;
  assign new_n3437_ = new_n3436_;
  assign new_n3438_ = new_n3435_;
  assign new_n3439_ = new_n1576_;
  assign new_n3440_ = new_n3439_;
  assign new_n3441_ = new_n3439_;
  assign new_n3442_ = new_n1612_;
  assign new_n3443_ = new_n1562_;
  assign new_n3444_ = new_n3443_;
  assign new_n3445_ = new_n3443_;
  assign new_n3446_ = new_n1978_;
  assign new_n3447_ = new_n1379_;
  assign new_n3448_ = new_n1297_;
  assign new_n3449_ = new_n3448_;
  assign new_n3450_ = new_n3448_;
  assign new_n3451_ = new_n1592_;
  assign new_n3452_ = new_n3451_;
  assign new_n3453_ = new_n3452_;
  assign new_n3454_ = new_n3452_;
  assign new_n3455_ = new_n3451_;
  assign new_n3456_ = new_n3455_;
  assign new_n3457_ = new_n1591_;
  assign new_n3458_ = new_n3457_;
  assign new_n3459_ = new_n3458_;
  assign new_n3460_ = new_n3458_;
  assign new_n3461_ = new_n3457_;
  assign new_n3462_ = new_n3461_;
  assign new_n3463_ = new_n1497_;
  assign new_n3464_ = new_n1383_;
  assign new_n3465_ = new_n2052_;
  assign new_n3466_ = new_n3465_;
  assign new_n3467_ = new_n2048_;
  assign new_n3468_ = new_n3467_;
  assign new_n3469_ = new_n2053_;
  assign new_n3470_ = new_n3469_;
  assign new_n3471_ = new_n2049_;
  assign new_n3472_ = new_n3471_;
  assign new_n3473_ = new_n1299_;
  assign new_n3474_ = new_n3473_;
  assign new_n3475_ = new_n3474_;
  assign new_n3476_ = new_n3473_;
  assign new_n3477_ = new_n1300_;
  assign new_n3478_ = new_n2057_;
  assign new_n3479_ = new_n2056_;
  assign new_n3480_ = new_n3479_;
  assign new_n3481_ = new_n2059_;
  assign new_n3482_ = new_n1390_;
  assign new_n3483_ = new_n3482_;
  assign new_n3484_ = new_n1389_;
  assign new_n3485_ = new_n3484_;
  assign new_n3486_ = new_n1523_;
  assign new_n3487_ = new_n3486_;
  assign new_n3488_ = new_n1391_;
  assign new_n3489_ = new_n3488_;
  assign new_n3490_ = new_n3488_;
  assign new_n3491_ = new_n1524_;
  assign new_n3492_ = new_n1392_;
  assign new_n3493_ = new_n3492_;
  assign new_n3494_ = new_n2083_;
  assign new_n3495_ = new_n2000_;
  assign new_n3496_ = new_n3495_;
  assign new_n3497_ = new_n3495_;
  assign new_n3498_ = new_n1544_;
  assign new_n3499_ = new_n3498_;
  assign new_n3500_ = new_n1543_;
  assign new_n3501_ = new_n3500_;
  assign new_n3502_ = new_n2087_;
  assign new_n3503_ = new_n3502_;
  assign new_n3504_ = new_n2086_;
  assign new_n3505_ = new_n3504_;
  assign new_n3506_ = new_n2093_;
  assign new_n3507_ = new_n1192_;
  assign new_n3508_ = new_n2004_;
  assign new_n3509_ = new_n1149_;
  assign new_n3510_ = new_n3509_;
  assign new_n3511_ = new_n2099_;
  assign new_n3512_ = new_n3511_;
  assign new_n3513_ = new_n3511_;
  assign new_n3514_ = new_n1368_;
  assign new_n3515_ = new_n1195_;
  assign new_n3516_ = new_n3515_;
  assign new_n3517_ = new_n3515_;
  assign new_n3518_ = new_n1919_;
  assign new_n3519_ = new_n1367_;
  assign new_n3520_ = new_n1473_;
  assign new_n3521_ = new_n1474_;
  assign new_n3522_ = new_n2109_;
  assign new_n3523_ = new_n2105_;
  assign new_n3524_ = new_n2108_;
  assign new_n3525_ = new_n2104_;
  assign new_n3526_ = new_n3525_;
  assign new_n3527_ = new_n1424_;
  assign new_n3528_ = new_n1136_;
  assign new_n3529_ = new_n1423_;
  assign new_n3530_ = new_n1135_;
  assign new_n3531_ = new_n2123_;
  assign new_n3532_ = new_n1836_;
  assign new_n3533_ = new_n2122_;
  assign new_n3534_ = new_n1835_;
  assign new_n3535_ = new_n3534_;
  assign new_n3536_ = new_n2124_;
  assign new_n3537_ = new_n2120_;
  assign new_n3538_ = new_n3537_;
  assign new_n3539_ = new_n3537_;
  assign new_n3540_ = new_n2125_;
  assign new_n3541_ = new_n2121_;
  assign new_n3542_ = new_n3541_;
  assign new_n3543_ = new_n3542_;
  assign new_n3544_ = new_n3541_;
  assign new_n3545_ = new_n2130_;
  assign new_n3546_ = new_n2114_;
  assign new_n3547_ = new_n1237_;
  assign new_n3548_ = new_n3547_;
  assign new_n3549_ = new_n3547_;
  assign new_n3550_ = new_n2115_;
  assign new_n3551_ = new_n3550_;
  assign new_n3552_ = new_n2131_;
  assign new_n3553_ = new_n1035_;
  assign new_n3554_ = new_n3553_;
  assign new_n3555_ = new_n3554_;
  assign new_n3556_ = new_n3554_;
  assign new_n3557_ = new_n3553_;
  assign new_n3558_ = new_n3557_;
  assign new_n3559_ = new_n1046_;
  assign new_n3560_ = new_n3559_;
  assign new_n3561_ = new_n3559_;
  assign new_n3562_ = new_n1845_;
  assign new_n3563_ = new_n1833_;
  assign new_n3564_ = new_n1834_;
  assign new_n3565_ = new_n1940_;
  assign new_n3566_ = new_n1243_;
  assign new_n3567_ = new_n3566_;
  assign new_n3568_ = new_n3567_;
  assign new_n3569_ = new_n3566_;
  assign new_n3570_ = new_n1214_;
  assign new_n3571_ = new_n3570_;
  assign new_n3572_ = new_n3570_;
  assign new_n3573_ = new_n1241_;
  assign new_n3574_ = new_n3573_;
  assign new_n3575_ = new_n3573_;
  assign new_n3576_ = new_n1245_;
  assign new_n3577_ = new_n3576_;
  assign new_n3578_ = new_n1074_;
  assign new_n3579_ = new_n1211_;
  assign new_n3580_ = new_n3579_;
  assign new_n3581_ = new_n3579_;
  assign new_n3582_ = new_n1240_;
  assign new_n3583_ = new_n3582_;
  assign new_n3584_ = new_n1062_;
  assign new_n3585_ = new_n2157_;
  assign new_n3586_ = new_n1103_;
  assign new_n3587_ = new_n3586_;
  assign new_n3588_ = new_n1041_;
  assign new_n3589_ = new_n2168_;
  assign new_n3590_ = new_n1851_;
  assign new_n3591_ = new_n1045_;
  assign new_n3592_ = new_n1039_;
  assign new_n3593_ = new_n1043_;
  assign new_n3594_ = new_n1239_;
  assign new_n3595_ = new_n3594_;
  assign new_n3596_ = new_n3595_;
  assign new_n3597_ = new_n3594_;
  assign new_n3598_ = new_n1044_;
  assign new_n3599_ = new_n1212_;
  assign new_n3600_ = new_n3599_;
  assign new_n3601_ = new_n3600_;
  assign new_n3602_ = new_n3600_;
  assign new_n3603_ = new_n3599_;
  assign new_n3604_ = new_n3603_;
  assign new_n3605_ = new_n1303_;
  assign new_n3606_ = new_n1051_;
  assign new_n3607_ = new_n3606_;
  assign new_n3608_ = new_n3606_;
  assign new_n3609_ = new_n1244_;
  assign new_n3610_ = new_n3609_;
  assign new_n3611_ = new_n3610_;
  assign new_n3612_ = new_n3611_;
  assign new_n3613_ = new_n3610_;
  assign new_n3614_ = new_n3609_;
  assign new_n3615_ = new_n3614_;
  assign new_n3616_ = new_n3614_;
  assign new_n3617_ = new_n1061_;
  assign new_n3618_ = new_n3617_;
  assign new_n3619_ = new_n1042_;
  assign new_n3620_ = new_n1242_;
  assign new_n3621_ = new_n3620_;
  assign new_n3622_ = new_n3621_;
  assign new_n3623_ = new_n3621_;
  assign new_n3624_ = new_n3620_;
  assign new_n3625_ = new_n1246_;
  assign new_n3626_ = new_n3625_;
  assign new_n3627_ = new_n3626_;
  assign new_n3628_ = new_n3626_;
  assign new_n3629_ = new_n3625_;
  assign new_n3630_ = new_n3629_;
  assign new_n3631_ = new_n1213_;
  assign new_n3632_ = new_n3631_;
  assign new_n3633_ = new_n3632_;
  assign new_n3634_ = new_n3632_;
  assign new_n3635_ = new_n3631_;
  assign new_n3636_ = new_n3635_;
  assign new_n3637_ = new_n1073_;
  assign new_n3638_ = new_n1119_;
  assign new_n3639_ = new_n3638_;
  assign new_n3640_ = new_n2246_;
  assign new_n3641_ = new_n2245_;
  assign new_n3642_ = new_n1121_;
  assign new_n3643_ = new_n3642_;
  assign new_n3644_ = new_n1420_;
  assign new_n3645_ = new_n1102_;
  assign new_n3646_ = new_n1139_;
  assign new_n3647_ = new_n1140_;
  assign new_n3648_ = new_n2268_;
  assign new_n3649_ = new_n1134_;
  assign new_n3650_ = new_n2267_;
  assign new_n3651_ = new_n1133_;
  assign new_n3652_ = new_n2274_;
  assign new_n3653_ = new_n3652_;
  assign new_n3654_ = new_n2047_;
  assign new_n3655_ = new_n2281_;
  assign new_n3656_ = new_n2278_;
  assign new_n3657_ = new_n3656_;
  assign new_n3658_ = new_n2288_;
  assign new_n3659_ = new_n3658_;
  assign new_n3660_ = new_n3658_;
  assign new_n3661_ = new_n2289_;
  assign new_n3662_ = new_n2290_;
  assign new_n3663_ = new_n1238_;
  assign new_n3664_ = new_n3663_;
  assign new_n3665_ = new_n2294_;
  assign new_n3666_ = new_n1998_;
  assign new_n3667_ = new_n1881_;
  assign new_n3668_ = new_n3667_;
  assign new_n3669_ = new_n1399_;
  assign new_n3670_ = new_n1221_;
  assign new_n3671_ = new_n3670_;
  assign new_n3672_ = new_n1155_;
  assign new_n3673_ = new_n2372_;
  assign new_n3674_ = new_n2373_;
  assign new_n3675_ = new_n2273_;
  assign new_n3676_ = new_n1977_;
  assign new_n3677_ = new_n3676_;
  assign new_n3678_ = new_n1949_;
  assign new_n3679_ = new_n3678_;
  assign new_n3680_ = new_n1397_;
  assign new_n3681_ = new_n1547_;
  assign new_n3682_ = new_n2422_;
  assign new_n3683_ = new_n2082_;
  assign new_n3684_ = new_n2002_;
  assign new_n3685_ = new_n3684_;
  assign new_n3686_ = new_n3685_;
  assign new_n3687_ = new_n3685_;
  assign new_n3688_ = new_n3684_;
  assign new_n3689_ = new_n3688_;
  assign new_n3690_ = new_n2028_;
  assign new_n3691_ = new_n2085_;
  assign new_n3692_ = new_n2092_;
  assign new_n3693_ = new_n2044_;
  assign new_n3694_ = new_n2095_;
  assign new_n3695_ = new_n1147_;
  assign new_n3696_ = new_n1219_;
  assign new_n3697_ = new_n1153_;
  assign new_n3698_ = new_n1159_;
  assign new_n3699_ = new_n1887_;
  assign new_n3700_ = new_n3699_;
  assign new_n3701_ = new_n3700_;
  assign new_n3702_ = new_n3700_;
  assign new_n3703_ = new_n3699_;
  assign new_n3704_ = new_n1160_;
  assign new_n3705_ = new_n1185_;
  assign new_n3706_ = new_n1889_;
  assign new_n3707_ = new_n3706_;
  assign new_n3708_ = new_n3707_;
  assign new_n3709_ = new_n3707_;
  assign new_n3710_ = new_n3706_;
  assign new_n3711_ = new_n925_;
  assign new_n3712_ = new_n3711_;
  assign new_n3713_ = new_n2445_;
  assign new_n3714_ = new_n3713_;
  assign new_n3715_ = new_n2296_;
  assign new_n3716_ = new_n2291_;
  assign new_n3717_ = new_n3716_;
  assign new_n3718_ = new_n921_;
  assign new_n3719_ = new_n2394_;
  assign new_n3720_ = new_n992_;
  assign new_n3721_ = new_n973_;
  assign new_n3722_ = new_n969_;
  assign new_n3723_ = new_n2453_;
  assign new_n3724_ = new_n1902_;
  assign new_n3725_ = new_n991_;
  assign new_n3726_ = new_n1880_;
  assign new_n3727_ = new_n3726_;
  assign new_n3728_ = new_n2460_;
  assign new_n3729_ = new_n1997_;
  assign new_n3730_ = new_n3729_;
  assign new_n3731_ = new_n2468_;
  assign new_n3732_ = new_n2459_;
  assign new_n3733_ = new_n3732_;
  assign new_n3734_ = new_n798_;
  assign new_n3735_ = new_n795_;
  assign new_n3736_ = new_n3735_;
  assign new_n3737_ = new_n805_;
  assign new_n3738_ = new_n2007_;
  assign new_n3739_ = new_n2005_;
  assign new_n3740_ = new_n2098_;
  assign new_n3741_ = new_n1287_;
  assign new_n3742_ = new_n3741_;
  assign new_n3743_ = new_n1904_;
  assign new_n3744_ = new_n937_;
  assign new_n3745_ = new_n3744_;
  assign new_n3746_ = new_n1918_;
  assign new_n3747_ = new_n3746_;
  assign new_n3748_ = new_n3746_;
  assign new_n3749_ = new_n1169_;
  assign new_n3750_ = new_n2101_;
  assign new_n3751_ = new_n1165_;
  assign new_n3752_ = new_n3751_;
  assign new_n3753_ = new_n2356_;
  assign new_n3754_ = new_n2102_;
  assign new_n3755_ = new_n1912_;
  assign new_n3756_ = new_n3755_;
  assign new_n3757_ = new_n2389_;
  assign new_n3758_ = new_n2276_;
  assign new_n3759_ = new_n2277_;
  assign new_n3760_ = new_n1521_;
  assign new_n3761_ = new_n3760_;
  assign new_n3762_ = new_n2519_;
  assign new_n3763_ = new_n3762_;
  assign new_n3764_ = new_n3762_;
  assign new_n3765_ = new_n2009_;
  assign new_n3766_ = new_n2525_;
  assign new_n3767_ = new_n2523_;
  assign new_n3768_ = new_n2008_;
  assign new_n3769_ = new_n1599_;
  assign new_n3770_ = new_n1504_;
  assign new_n3771_ = new_n3770_;
  assign new_n3772_ = new_n1499_;
  assign new_n3773_ = new_n1503_;
  assign new_n3774_ = new_n3773_;
  assign new_n3775_ = new_n2552_;
  assign new_n3776_ = new_n2006_;
  assign new_n3777_ = new_n2003_;
  assign new_n3778_ = new_n2421_;
  assign new_n3779_ = new_n2075_;
  assign new_n3780_ = new_n2424_;
  assign new_n3781_ = new_n2430_;
  assign new_n3782_ = new_n2427_;
  assign new_n3783_ = new_n801_;
  assign new_n3784_ = new_n3783_;
  assign new_n3785_ = new_n3784_;
  assign new_n3786_ = new_n3785_;
  assign new_n3787_ = new_n3785_;
  assign new_n3788_ = new_n3784_;
  assign new_n3789_ = new_n3783_;
  assign new_n3790_ = new_n3789_;
  assign new_n3791_ = new_n3789_;
  assign new_n3792_ = new_n817_;
  assign new_n3793_ = new_n3792_;
  assign new_n3794_ = new_n3792_;
  assign new_n3795_ = new_n815_;
  assign new_n3796_ = new_n819_;
  assign new_n3797_ = new_n3796_;
  assign new_n3798_ = new_n939_;
  assign new_n3799_ = new_n2010_;
  assign new_n3800_ = new_n941_;
  assign new_n3801_ = new_n2046_;
  assign new_n3802_ = new_n1597_;
  assign new_n3803_ = new_n3802_;
  assign new_n3804_ = new_n1381_;
  assign new_n3805_ = new_n3804_;
  assign new_n3806_ = new_n3805_;
  assign new_n3807_ = new_n3804_;
  assign new_n3808_ = new_n1382_;
  assign new_n3809_ = new_n3808_;
  assign new_n3810_ = new_n3808_;
  assign new_n3811_ = new_n949_;
  assign new_n3812_ = new_n2551_;
  assign new_n3813_ = new_n1613_;
  assign new_n3814_ = new_n2054_;
  assign new_n3815_ = new_n802_;
  assign new_n3816_ = new_n3815_;
  assign new_n3817_ = new_n3816_;
  assign new_n3818_ = new_n3815_;
  assign new_n3819_ = new_n799_;
  assign new_n3820_ = new_n3819_;
  assign new_n3821_ = new_n3820_;
  assign new_n3822_ = new_n3819_;
  assign new_n3823_ = new_n2471_;
  assign new_n3824_ = new_n800_;
  assign new_n3825_ = new_n803_;
  assign new_n3826_ = new_n3825_;
  assign new_n3827_ = new_n1546_;
  assign new_n3828_ = new_n1614_;
  assign new_n3829_ = new_n2055_;
  assign new_n3830_ = new_n2623_;
  assign new_n3831_ = new_n2001_;
  assign new_n3832_ = new_n3831_;
  assign new_n3833_ = new_n2522_;
  assign new_n3834_ = new_n3833_;
  assign new_n3835_ = new_n2634_;
  assign new_n3836_ = new_n2535_;
  assign new_n3837_ = new_n3836_;
  assign new_n3838_ = new_n796_;
  assign new_n3839_ = new_n3838_;
  assign new_n3840_ = new_n2641_;
  assign new_n3841_ = new_n2472_;
  assign new_n3842_ = new_n3841_;
  assign new_n3843_ = new_n2511_;
  assign new_n3844_ = new_n2412_;
  assign new_n3845_ = new_n2554_;
  assign new_n3846_ = new_n2565_;
  assign new_n3847_ = new_n2564_;
  assign new_n3848_ = new_n820_;
  assign new_n3849_ = new_n2568_;
  assign new_n3850_ = new_n2567_;
  assign new_n3851_ = new_n2652_;
  assign new_n3852_ = new_n875_;
  assign new_n3853_ = new_n2606_;
  assign new_n3854_ = new_n3853_;
  assign new_n3855_ = new_n3853_;
  assign new_n3856_ = new_n2566_;
  assign new_n3857_ = new_n3856_;
  assign new_n3858_ = new_n3856_;
  assign new_n3859_ = new_n862_;
  assign new_n3860_ = new_n2608_;
  assign new_n3861_ = new_n2645_;
  assign new_n3862_ = new_n863_;
  assign new_n3863_ = new_n3862_;
  assign new_n3864_ = new_n2644_;
  assign new_n3865_ = new_n2607_;
  assign new_n3866_ = new_n873_;
  assign new_n3867_ = new_n859_;
  assign new_n3868_ = new_n821_;
  assign new_n3869_ = new_n861_;
  assign new_n3870_ = new_n2654_;
  always @ (posedge clock) begin
    n1752_lo <= n4070_li003_li003;
    n1776_lo <= n4094_li011_li011;
    n1824_lo <= n4142_li027_li027;
    n1836_lo <= n4154_li031_li031;
    n1848_lo <= n4166_li035_li035;
    n1860_lo <= n4178_li039_li039;
    n1872_lo <= n4190_li043_li043;
    n1884_lo <= n4202_li047_li047;
    n1896_lo <= n4214_li051_li051;
    n1908_lo <= n4226_li055_li055;
    n1911_lo <= n4229_li056_li056;
    n1914_lo <= n4232_li057_li057;
    n1923_lo <= n4241_li060_li060;
    n1926_lo <= n4244_li061_li061;
    n1935_lo <= n4253_li064_li064;
    n1938_lo <= n4256_li065_li065;
    n1947_lo <= n4265_li068_li068;
    n1950_lo <= n4268_li069_li069;
    n1959_lo <= n4277_li072_li072;
    n1962_lo <= n4280_li073_li073;
    n1971_lo <= n4289_li076_li076;
    n1974_lo <= n4292_li077_li077;
    n1983_lo <= n4301_li080_li080;
    n1995_lo <= n4313_li084_li084;
    n2055_lo <= n4373_li104_li104;
    n2064_lo <= n4382_li107_li107;
    n2067_lo <= n4385_li108_li108;
    n2079_lo <= n4397_li112_li112;
    n2100_lo <= n4418_li119_li119;
    n2112_lo <= n4430_li123_li123;
    n2124_lo <= n4442_li127_li127;
    n2136_lo <= n4454_li131_li131;
    n2148_lo <= n4466_li135_li135;
    n2160_lo <= n4478_li139_li139;
    n2172_lo <= n4490_li143_li143;
    n2184_lo <= n4502_li147_li147;
    n2235_lo <= n4553_li164_li164;
    n2238_lo <= n4556_li165_li165;
    n2247_lo <= n4565_li168_li168;
    n2250_lo <= n4568_li169_li169;
    n2259_lo <= n4577_li172_li172;
    n2262_lo <= n4580_li173_li173;
    n2271_lo <= n4589_li176_li176;
    n2274_lo <= n4592_li177_li177;
    n2283_lo <= n4601_li180_li180;
    n2286_lo <= n4604_li181_li181;
    n2289_lo <= n4607_li182_li182;
    n2295_lo <= n4613_li184_li184;
    n2298_lo <= n4616_li185_li185;
    n2304_lo <= n4622_li187_li187;
    n2307_lo <= n4625_li188_li188;
    n2316_lo <= n4634_li191_li191;
    n2331_lo <= n4649_li196_li196;
    n2334_lo <= n4652_li197_li197;
    n2337_lo <= n4655_li198_li198;
    n2340_lo <= n4658_li199_li199;
    n2071_o2 <= n2071_i2;
    n2080_o2 <= n2080_i2;
    n2137_o2 <= n2137_i2;
    n2368_o2 <= n2368_i2;
    n2383_o2 <= n2383_i2;
    n2405_o2 <= n2405_i2;
    n2471_o2 <= n2471_i2;
    n2617_o2 <= n2617_i2;
    n2765_o2 <= n2765_i2;
    n2775_o2 <= n2775_i2;
    n2829_o2 <= n2829_i2;
    n2579_o2 <= n2579_i2;
    n2580_o2 <= n2580_i2;
    n2618_o2 <= n2618_i2;
    n2619_o2 <= n2619_i2;
    n2620_o2 <= n2620_i2;
    n2621_o2 <= n2621_i2;
    n2622_o2 <= n2622_i2;
    n2623_o2 <= n2623_i2;
    n2624_o2 <= n2624_i2;
    n2625_o2 <= n2625_i2;
    n2626_o2 <= n2626_i2;
    n2627_o2 <= n2627_i2;
    n3029_o2 <= n3029_i2;
    n3035_o2 <= n3035_i2;
    n2643_o2 <= n2643_i2;
    n2644_o2 <= n2644_i2;
    n2645_o2 <= n2645_i2;
    n327_inv <= n2640_i2;
    n2658_o2 <= n2658_i2;
    n2659_o2 <= n2659_i2;
    n2674_o2 <= n2674_i2;
    n2675_o2 <= n2675_i2;
    n2676_o2 <= n2676_i2;
    n3119_o2 <= n3119_i2;
    n3153_o2 <= n3153_i2;
    n351_inv <= n2681_i2;
    n2729_o2 <= n2729_i2;
    n2730_o2 <= n2730_i2;
    n2731_o2 <= n2731_i2;
    n698_o2 <= n698_i2;
    n366_inv <= n677_i2;
    n2757_o2 <= n2757_i2;
    n2758_o2 <= n2758_i2;
    n1000_o2 <= n1000_i2;
    n1160_o2 <= n1160_i2;
    n1153_o2 <= n1153_i2;
    n2793_o2 <= n2793_i2;
    n2794_o2 <= n2794_i2;
    n2795_o2 <= n2795_i2;
    n1001_o2 <= n1001_i2;
    n2859_o2 <= n2859_i2;
    n744_o2 <= n744_i2;
    n402_inv <= n2908_i2;
    n2926_o2 <= n2926_i2;
    n408_inv <= n2928_i2;
    n2966_o2 <= n2966_i2;
    n2967_o2 <= n2967_i2;
    n2947_o2 <= n2947_i2;
    n1010_o2 <= n1010_i2;
    n2976_o2 <= n2976_i2;
    n3069_o2 <= n3069_i2;
    n3028_o2 <= n3028_i2;
    n3081_o2 <= n3081_i2;
    n3082_o2 <= n3082_i2;
    n3142_o2 <= n3142_i2;
    n3214_o2 <= n3214_i2;
    n2992_o2 <= n2992_i2;
    n2993_o2 <= n2993_i2;
    n870_o2 <= n870_i2;
    n3086_o2 <= n3086_i2;
    n3087_o2 <= n3087_i2;
    n3088_o2 <= n3088_i2;
    n3089_o2 <= n3089_i2;
    n3090_o2 <= n3090_i2;
    n3091_o2 <= n3091_i2;
    n3092_o2 <= n3092_i2;
    n3093_o2 <= n3093_i2;
    n3094_o2 <= n3094_i2;
    n3095_o2 <= n3095_i2;
    n483_inv <= n3136_i2;
    n3170_o2 <= n3170_i2;
    n3171_o2 <= n3171_i2;
    n3172_o2 <= n3172_i2;
    n3179_o2 <= n3179_i2;
    n498_inv <= n3180_i2;
    n3193_o2 <= n3193_i2;
    n3211_o2 <= n3211_i2;
    n3212_o2 <= n3212_i2;
    n3213_o2 <= n3213_i2;
    n513_inv <= n3219_i2;
    n1125_o2 <= n1125_i2;
    n1081_o2 <= n1081_i2;
    n1139_o2 <= n1139_i2;
    n3245_o2 <= n3245_i2;
    n3246_o2 <= n3246_i2;
    n3247_o2 <= n3247_i2;
    lo074_buf_o2 <= lo074_buf_i2;
    lo078_buf_o2 <= lo078_buf_i2;
    lo186_buf_o2 <= lo186_buf_i2;
    lo118_buf_o2 <= lo118_buf_i2;
    lo146_buf_o2 <= lo146_buf_i2;
    n1038_o2 <= n1038_i2;
    n1044_o2 <= n1044_i2;
    n555_inv <= n980_i2;
    n558_inv <= n1145_i2;
    lo026_buf_o2 <= lo026_buf_i2;
    lo030_buf_o2 <= lo030_buf_i2;
    lo090_buf_o2 <= lo090_buf_i2;
    lo094_buf_o2 <= lo094_buf_i2;
    lo098_buf_o2 <= lo098_buf_i2;
    lo102_buf_o2 <= lo102_buf_i2;
    lo066_buf_o2 <= lo066_buf_i2;
    lo070_buf_o2 <= lo070_buf_i2;
    n1202_o2 <= n1202_i2;
    n1003_o2 <= n1003_i2;
    n1031_o2 <= n1031_i2;
    n1034_o2 <= n1034_i2;
    n1040_o2 <= n1040_i2;
    n1046_o2 <= n1046_i2;
    n1380_o2 <= n1380_i2;
    n1425_o2 <= n1425_i2;
    n697_o2 <= n697_i2;
    n1143_o2 <= n1143_i2;
    n673_o2 <= n673_i2;
    n789_o2 <= n789_i2;
    n786_o2 <= n786_i2;
    n1047_o2 <= n1047_i2;
    n1036_o2 <= n1036_i2;
    n1307_o2 <= n1307_i2;
    n1035_o2 <= n1035_i2;
    n1297_o2 <= n1297_i2;
    n1099_o2 <= n1099_i2;
    n1128_o2 <= n1128_i2;
    n645_inv <= n674_i2;
    n826_o2 <= n826_i2;
    n853_o2 <= n853_i2;
    n654_inv <= n951_i2;
    n700_o2 <= n700_i2;
    n884_o2 <= n884_i2;
    lo082_buf_o2 <= lo082_buf_i2;
    lo086_buf_o2 <= lo086_buf_i2;
    n801_o2 <= n801_i2;
    n840_o2 <= n840_i2;
    n675_inv <= n866_i2;
    lo002_buf_o2 <= lo002_buf_i2;
    lo010_buf_o2 <= lo010_buf_i2;
    lo166_buf_o2 <= lo166_buf_i2;
    lo170_buf_o2 <= lo170_buf_i2;
    n1426_o2 <= n1426_i2;
    n1082_o2 <= n1082_i2;
    n1310_o2 <= n1310_i2;
    n1015_o2 <= n1015_i2;
    n1206_o2 <= n1206_i2;
    n1262_o2 <= n1262_i2;
    n1456_o2 <= n1456_i2;
    n1244_o2 <= n1244_i2;
    n1280_o2 <= n1280_i2;
    n1290_o2 <= n1290_i2;
    n1012_o2 <= n1012_i2;
    n1074_o2 <= n1074_i2;
    n1112_o2 <= n1112_i2;
    n1212_o2 <= n1212_i2;
    n1454_o2 <= n1454_i2;
    n1182_o2 <= n1182_i2;
    n1220_o2 <= n1220_i2;
    n701_o2 <= n701_i2;
    n744_inv <= n973_i2;
    n1282_o2 <= n1282_i2;
    n1144_o2 <= n1144_i2;
    n1278_o2 <= n1278_i2;
    n1459_o2 <= n1459_i2;
    n1324_o2 <= n1324_i2;
    n1288_o2 <= n1288_i2;
    n1271_o2 <= n1271_i2;
    n1132_o2 <= n1132_i2;
    n1231_o2 <= n1231_i2;
    n1462_o2 <= n1462_i2;
    n1482_o2 <= n1482_i2;
    n994_o2 <= n994_i2;
    n998_o2 <= n998_i2;
    lo106_buf_o2 <= lo106_buf_i2;
    n769_o2 <= n769_i2;
    n814_o2 <= n814_i2;
    n841_o2 <= n841_i2;
    n867_o2 <= n867_i2;
    lo006_buf_o2 <= lo006_buf_i2;
    lo014_buf_o2 <= lo014_buf_i2;
    lo022_buf_o2 <= lo022_buf_i2;
    lo042_buf_o2 <= lo042_buf_i2;
    lo046_buf_o2 <= lo046_buf_i2;
    lo050_buf_o2 <= lo050_buf_i2;
    lo054_buf_o2 <= lo054_buf_i2;
    lo130_buf_o2 <= lo130_buf_i2;
    lo134_buf_o2 <= lo134_buf_i2;
    lo154_buf_o2 <= lo154_buf_i2;
    lo174_buf_o2 <= lo174_buf_i2;
    lo178_buf_o2 <= lo178_buf_i2;
    n1007_o2 <= n1007_i2;
    n1294_o2 <= n1294_i2;
    n1084_o2 <= n1084_i2;
    n1399_o2 <= n1399_i2;
    n1311_o2 <= n1311_i2;
    n1392_o2 <= n1392_i2;
    n1102_o2 <= n1102_i2;
    n1041_o2 <= n1041_i2;
    n1298_o2 <= n1298_i2;
    n738_o2 <= n738_i2;
    n1214_o2 <= n1214_i2;
    n1222_o2 <= n1222_i2;
    n1155_o2 <= n1155_i2;
    n1147_o2 <= n1147_i2;
    n1393_o2 <= n1393_i2;
    n999_o2 <= n999_i2;
    n1306_o2 <= n1306_i2;
    n1312_o2 <= n1312_i2;
    n1382_o2 <= n1382_i2;
    n1383_o2 <= n1383_i2;
    n1152_o2 <= n1152_i2;
    n1334_o2 <= n1334_i2;
    n1335_o2 <= n1335_i2;
    n906_inv <= n695_i2;
    n773_o2 <= n773_i2;
    lo190_buf_o2 <= lo190_buf_i2;
    n1368_o2 <= n1368_i2;
    n1362_o2 <= n1362_i2;
    n1406_o2 <= n1406_i2;
    n1403_o2 <= n1403_i2;
    n741_o2 <= n741_i2;
    n1407_o2 <= n1407_i2;
    n1395_o2 <= n1395_i2;
    n1359_o2 <= n1359_i2;
    n1159_o2 <= n1159_i2;
    n1221_o2 <= n1221_i2;
    n945_inv <= n987_i2;
    n989_o2 <= n989_i2;
    n881_o2 <= n881_i2;
    n1340_o2 <= n1340_i2;
    n1341_o2 <= n1341_i2;
    n906_o2 <= n906_i2;
    n1388_o2 <= n1388_i2;
    n791_o2 <= n791_i2;
    n1372_o2 <= n1372_i2;
    n815_o2 <= n815_i2;
    n868_o2 <= n868_i2;
    lo018_buf_o2 <= lo018_buf_i2;
    lo138_buf_o2 <= lo138_buf_i2;
    lo158_buf_o2 <= lo158_buf_i2;
    n780_o2 <= n780_i2;
    n728_o2 <= n728_i2;
    n993_inv <= n676_i2;
    n929_o2 <= n929_i2;
    n955_o2 <= n955_i2;
    n938_o2 <= n938_i2;
    n1117_o2 <= n1117_i2;
    n1121_o2 <= n1121_i2;
    n965_o2 <= n965_i2;
    n752_o2 <= n752_i2;
    n753_o2 <= n753_i2;
    n760_o2 <= n760_i2;
    n770_o2 <= n770_i2;
    n923_o2 <= n923_i2;
    n947_o2 <= n947_i2;
    n897_o2 <= n897_i2;
    n919_o2 <= n919_i2;
    n895_o2 <= n895_i2;
    n917_o2 <= n917_i2;
    n751_o2 <= n751_i2;
    n774_o2 <= n774_i2;
    lo126_buf_o2 <= lo126_buf_i2;
    lo142_buf_o2 <= lo142_buf_i2;
    lo162_buf_o2 <= lo162_buf_i2;
    n1059_inv <= n990_i2;
    n792_o2 <= n792_i2;
    n869_o2 <= n869_i2;
    n1068_inv <= n848_i2;
    lo024_buf_o2 <= lo024_buf_i2;
    lo028_buf_o2 <= lo028_buf_i2;
    lo088_buf_o2 <= lo088_buf_i2;
    lo092_buf_o2 <= lo092_buf_i2;
    lo096_buf_o2 <= lo096_buf_i2;
    lo100_buf_o2 <= lo100_buf_i2;
    n763_o2 <= n763_i2;
    n754_o2 <= n754_i2;
    n755_o2 <= n755_i2;
    n822_o2 <= n822_i2;
    n849_o2 <= n849_i2;
    n777_o2 <= n777_i2;
    n778_o2 <= n778_i2;
    n820_o2 <= n820_i2;
    n846_o2 <= n846_i2;
    n806_o2 <= n806_i2;
    n771_o2 <= n771_i2;
    n854_o2 <= n854_i2;
    n828_o2 <= n828_i2;
    lo117_buf_o2 <= lo117_buf_i2;
    lo145_buf_o2 <= lo145_buf_i2;
    n762_o2 <= n762_i2;
    n805_o2 <= n805_i2;
    n859_o2 <= n859_i2;
    n833_o2 <= n833_i2;
    lo034_buf_o2 <= lo034_buf_i2;
    lo038_buf_o2 <= lo038_buf_i2;
    lo122_buf_o2 <= lo122_buf_i2;
    lo150_buf_o2 <= lo150_buf_i2;
  end
  initial begin
    n1752_lo <= 1'b0;
    n1776_lo <= 1'b0;
    n1824_lo <= 1'b0;
    n1836_lo <= 1'b0;
    n1848_lo <= 1'b0;
    n1860_lo <= 1'b0;
    n1872_lo <= 1'b0;
    n1884_lo <= 1'b0;
    n1896_lo <= 1'b0;
    n1908_lo <= 1'b0;
    n1911_lo <= 1'b0;
    n1914_lo <= 1'b0;
    n1923_lo <= 1'b0;
    n1926_lo <= 1'b0;
    n1935_lo <= 1'b0;
    n1938_lo <= 1'b0;
    n1947_lo <= 1'b0;
    n1950_lo <= 1'b0;
    n1959_lo <= 1'b0;
    n1962_lo <= 1'b0;
    n1971_lo <= 1'b0;
    n1974_lo <= 1'b0;
    n1983_lo <= 1'b0;
    n1995_lo <= 1'b0;
    n2055_lo <= 1'b0;
    n2064_lo <= 1'b0;
    n2067_lo <= 1'b0;
    n2079_lo <= 1'b0;
    n2100_lo <= 1'b0;
    n2112_lo <= 1'b0;
    n2124_lo <= 1'b0;
    n2136_lo <= 1'b0;
    n2148_lo <= 1'b0;
    n2160_lo <= 1'b0;
    n2172_lo <= 1'b0;
    n2184_lo <= 1'b0;
    n2235_lo <= 1'b0;
    n2238_lo <= 1'b0;
    n2247_lo <= 1'b0;
    n2250_lo <= 1'b0;
    n2259_lo <= 1'b0;
    n2262_lo <= 1'b0;
    n2271_lo <= 1'b0;
    n2274_lo <= 1'b0;
    n2283_lo <= 1'b0;
    n2286_lo <= 1'b0;
    n2289_lo <= 1'b0;
    n2295_lo <= 1'b0;
    n2298_lo <= 1'b0;
    n2304_lo <= 1'b0;
    n2307_lo <= 1'b0;
    n2316_lo <= 1'b0;
    n2331_lo <= 1'b0;
    n2334_lo <= 1'b0;
    n2337_lo <= 1'b0;
    n2340_lo <= 1'b0;
    n2071_o2 <= 1'b0;
    n2080_o2 <= 1'b0;
    n2137_o2 <= 1'b0;
    n2368_o2 <= 1'b0;
    n2383_o2 <= 1'b0;
    n2405_o2 <= 1'b0;
    n2471_o2 <= 1'b0;
    n2617_o2 <= 1'b0;
    n2765_o2 <= 1'b0;
    n2775_o2 <= 1'b0;
    n2829_o2 <= 1'b0;
    n2579_o2 <= 1'b0;
    n2580_o2 <= 1'b0;
    n2618_o2 <= 1'b0;
    n2619_o2 <= 1'b0;
    n2620_o2 <= 1'b0;
    n2621_o2 <= 1'b0;
    n2622_o2 <= 1'b0;
    n2623_o2 <= 1'b0;
    n2624_o2 <= 1'b0;
    n2625_o2 <= 1'b0;
    n2626_o2 <= 1'b0;
    n2627_o2 <= 1'b0;
    n3029_o2 <= 1'b0;
    n3035_o2 <= 1'b0;
    n2643_o2 <= 1'b0;
    n2644_o2 <= 1'b0;
    n2645_o2 <= 1'b0;
    n327_inv <= 1'b0;
    n2658_o2 <= 1'b0;
    n2659_o2 <= 1'b0;
    n2674_o2 <= 1'b0;
    n2675_o2 <= 1'b0;
    n2676_o2 <= 1'b0;
    n3119_o2 <= 1'b0;
    n3153_o2 <= 1'b0;
    n351_inv <= 1'b0;
    n2729_o2 <= 1'b0;
    n2730_o2 <= 1'b0;
    n2731_o2 <= 1'b0;
    n698_o2 <= 1'b0;
    n366_inv <= 1'b0;
    n2757_o2 <= 1'b0;
    n2758_o2 <= 1'b0;
    n1000_o2 <= 1'b0;
    n1160_o2 <= 1'b0;
    n1153_o2 <= 1'b0;
    n2793_o2 <= 1'b0;
    n2794_o2 <= 1'b0;
    n2795_o2 <= 1'b0;
    n1001_o2 <= 1'b0;
    n2859_o2 <= 1'b0;
    n744_o2 <= 1'b0;
    n402_inv <= 1'b0;
    n2926_o2 <= 1'b0;
    n408_inv <= 1'b0;
    n2966_o2 <= 1'b0;
    n2967_o2 <= 1'b0;
    n2947_o2 <= 1'b0;
    n1010_o2 <= 1'b0;
    n2976_o2 <= 1'b0;
    n3069_o2 <= 1'b0;
    n3028_o2 <= 1'b0;
    n3081_o2 <= 1'b0;
    n3082_o2 <= 1'b0;
    n3142_o2 <= 1'b0;
    n3214_o2 <= 1'b0;
    n2992_o2 <= 1'b0;
    n2993_o2 <= 1'b0;
    n870_o2 <= 1'b0;
    n3086_o2 <= 1'b0;
    n3087_o2 <= 1'b0;
    n3088_o2 <= 1'b0;
    n3089_o2 <= 1'b0;
    n3090_o2 <= 1'b0;
    n3091_o2 <= 1'b0;
    n3092_o2 <= 1'b0;
    n3093_o2 <= 1'b0;
    n3094_o2 <= 1'b0;
    n3095_o2 <= 1'b0;
    n483_inv <= 1'b0;
    n3170_o2 <= 1'b0;
    n3171_o2 <= 1'b0;
    n3172_o2 <= 1'b0;
    n3179_o2 <= 1'b0;
    n498_inv <= 1'b0;
    n3193_o2 <= 1'b0;
    n3211_o2 <= 1'b0;
    n3212_o2 <= 1'b0;
    n3213_o2 <= 1'b0;
    n513_inv <= 1'b0;
    n1125_o2 <= 1'b0;
    n1081_o2 <= 1'b0;
    n1139_o2 <= 1'b0;
    n3245_o2 <= 1'b0;
    n3246_o2 <= 1'b0;
    n3247_o2 <= 1'b0;
    lo074_buf_o2 <= 1'b0;
    lo078_buf_o2 <= 1'b0;
    lo186_buf_o2 <= 1'b0;
    lo118_buf_o2 <= 1'b0;
    lo146_buf_o2 <= 1'b0;
    n1038_o2 <= 1'b0;
    n1044_o2 <= 1'b0;
    n555_inv <= 1'b0;
    n558_inv <= 1'b0;
    lo026_buf_o2 <= 1'b0;
    lo030_buf_o2 <= 1'b0;
    lo090_buf_o2 <= 1'b0;
    lo094_buf_o2 <= 1'b0;
    lo098_buf_o2 <= 1'b0;
    lo102_buf_o2 <= 1'b0;
    lo066_buf_o2 <= 1'b0;
    lo070_buf_o2 <= 1'b0;
    n1202_o2 <= 1'b0;
    n1003_o2 <= 1'b0;
    n1031_o2 <= 1'b0;
    n1034_o2 <= 1'b0;
    n1040_o2 <= 1'b0;
    n1046_o2 <= 1'b0;
    n1380_o2 <= 1'b0;
    n1425_o2 <= 1'b0;
    n697_o2 <= 1'b0;
    n1143_o2 <= 1'b0;
    n673_o2 <= 1'b0;
    n789_o2 <= 1'b0;
    n786_o2 <= 1'b0;
    n1047_o2 <= 1'b0;
    n1036_o2 <= 1'b0;
    n1307_o2 <= 1'b0;
    n1035_o2 <= 1'b0;
    n1297_o2 <= 1'b0;
    n1099_o2 <= 1'b0;
    n1128_o2 <= 1'b0;
    n645_inv <= 1'b0;
    n826_o2 <= 1'b0;
    n853_o2 <= 1'b0;
    n654_inv <= 1'b0;
    n700_o2 <= 1'b0;
    n884_o2 <= 1'b0;
    lo082_buf_o2 <= 1'b0;
    lo086_buf_o2 <= 1'b0;
    n801_o2 <= 1'b0;
    n840_o2 <= 1'b0;
    n675_inv <= 1'b0;
    lo002_buf_o2 <= 1'b0;
    lo010_buf_o2 <= 1'b0;
    lo166_buf_o2 <= 1'b0;
    lo170_buf_o2 <= 1'b0;
    n1426_o2 <= 1'b0;
    n1082_o2 <= 1'b0;
    n1310_o2 <= 1'b0;
    n1015_o2 <= 1'b0;
    n1206_o2 <= 1'b0;
    n1262_o2 <= 1'b0;
    n1456_o2 <= 1'b0;
    n1244_o2 <= 1'b0;
    n1280_o2 <= 1'b0;
    n1290_o2 <= 1'b0;
    n1012_o2 <= 1'b0;
    n1074_o2 <= 1'b0;
    n1112_o2 <= 1'b0;
    n1212_o2 <= 1'b0;
    n1454_o2 <= 1'b0;
    n1182_o2 <= 1'b0;
    n1220_o2 <= 1'b0;
    n701_o2 <= 1'b0;
    n744_inv <= 1'b0;
    n1282_o2 <= 1'b0;
    n1144_o2 <= 1'b0;
    n1278_o2 <= 1'b0;
    n1459_o2 <= 1'b0;
    n1324_o2 <= 1'b0;
    n1288_o2 <= 1'b0;
    n1271_o2 <= 1'b0;
    n1132_o2 <= 1'b0;
    n1231_o2 <= 1'b0;
    n1462_o2 <= 1'b0;
    n1482_o2 <= 1'b0;
    n994_o2 <= 1'b0;
    n998_o2 <= 1'b0;
    lo106_buf_o2 <= 1'b0;
    n769_o2 <= 1'b0;
    n814_o2 <= 1'b0;
    n841_o2 <= 1'b0;
    n867_o2 <= 1'b0;
    lo006_buf_o2 <= 1'b0;
    lo014_buf_o2 <= 1'b0;
    lo022_buf_o2 <= 1'b0;
    lo042_buf_o2 <= 1'b0;
    lo046_buf_o2 <= 1'b0;
    lo050_buf_o2 <= 1'b0;
    lo054_buf_o2 <= 1'b0;
    lo130_buf_o2 <= 1'b0;
    lo134_buf_o2 <= 1'b0;
    lo154_buf_o2 <= 1'b0;
    lo174_buf_o2 <= 1'b0;
    lo178_buf_o2 <= 1'b0;
    n1007_o2 <= 1'b0;
    n1294_o2 <= 1'b0;
    n1084_o2 <= 1'b0;
    n1399_o2 <= 1'b0;
    n1311_o2 <= 1'b0;
    n1392_o2 <= 1'b0;
    n1102_o2 <= 1'b0;
    n1041_o2 <= 1'b0;
    n1298_o2 <= 1'b0;
    n738_o2 <= 1'b0;
    n1214_o2 <= 1'b0;
    n1222_o2 <= 1'b0;
    n1155_o2 <= 1'b0;
    n1147_o2 <= 1'b0;
    n1393_o2 <= 1'b0;
    n999_o2 <= 1'b0;
    n1306_o2 <= 1'b0;
    n1312_o2 <= 1'b0;
    n1382_o2 <= 1'b0;
    n1383_o2 <= 1'b0;
    n1152_o2 <= 1'b0;
    n1334_o2 <= 1'b0;
    n1335_o2 <= 1'b0;
    n906_inv <= 1'b0;
    n773_o2 <= 1'b0;
    lo190_buf_o2 <= 1'b0;
    n1368_o2 <= 1'b0;
    n1362_o2 <= 1'b0;
    n1406_o2 <= 1'b0;
    n1403_o2 <= 1'b0;
    n741_o2 <= 1'b0;
    n1407_o2 <= 1'b0;
    n1395_o2 <= 1'b0;
    n1359_o2 <= 1'b0;
    n1159_o2 <= 1'b0;
    n1221_o2 <= 1'b0;
    n945_inv <= 1'b0;
    n989_o2 <= 1'b0;
    n881_o2 <= 1'b0;
    n1340_o2 <= 1'b0;
    n1341_o2 <= 1'b0;
    n906_o2 <= 1'b0;
    n1388_o2 <= 1'b0;
    n791_o2 <= 1'b0;
    n1372_o2 <= 1'b0;
    n815_o2 <= 1'b0;
    n868_o2 <= 1'b0;
    lo018_buf_o2 <= 1'b0;
    lo138_buf_o2 <= 1'b0;
    lo158_buf_o2 <= 1'b0;
    n780_o2 <= 1'b0;
    n728_o2 <= 1'b0;
    n993_inv <= 1'b0;
    n929_o2 <= 1'b0;
    n955_o2 <= 1'b0;
    n938_o2 <= 1'b0;
    n1117_o2 <= 1'b0;
    n1121_o2 <= 1'b0;
    n965_o2 <= 1'b0;
    n752_o2 <= 1'b0;
    n753_o2 <= 1'b0;
    n760_o2 <= 1'b0;
    n770_o2 <= 1'b0;
    n923_o2 <= 1'b0;
    n947_o2 <= 1'b0;
    n897_o2 <= 1'b0;
    n919_o2 <= 1'b0;
    n895_o2 <= 1'b0;
    n917_o2 <= 1'b0;
    n751_o2 <= 1'b0;
    n774_o2 <= 1'b0;
    lo126_buf_o2 <= 1'b0;
    lo142_buf_o2 <= 1'b0;
    lo162_buf_o2 <= 1'b0;
    n1059_inv <= 1'b0;
    n792_o2 <= 1'b0;
    n869_o2 <= 1'b0;
    n1068_inv <= 1'b0;
    lo024_buf_o2 <= 1'b0;
    lo028_buf_o2 <= 1'b0;
    lo088_buf_o2 <= 1'b0;
    lo092_buf_o2 <= 1'b0;
    lo096_buf_o2 <= 1'b0;
    lo100_buf_o2 <= 1'b0;
    n763_o2 <= 1'b0;
    n754_o2 <= 1'b0;
    n755_o2 <= 1'b0;
    n822_o2 <= 1'b0;
    n849_o2 <= 1'b0;
    n777_o2 <= 1'b0;
    n778_o2 <= 1'b0;
    n820_o2 <= 1'b0;
    n846_o2 <= 1'b0;
    n806_o2 <= 1'b0;
    n771_o2 <= 1'b0;
    n854_o2 <= 1'b0;
    n828_o2 <= 1'b0;
    lo117_buf_o2 <= 1'b0;
    lo145_buf_o2 <= 1'b0;
    n762_o2 <= 1'b0;
    n805_o2 <= 1'b0;
    n859_o2 <= 1'b0;
    n833_o2 <= 1'b0;
    lo034_buf_o2 <= 1'b0;
    lo038_buf_o2 <= 1'b0;
    lo122_buf_o2 <= 1'b0;
    lo150_buf_o2 <= 1'b0;
  end
endmodule


