
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G33,
  G34,
  G35,
  G36,
  G37,
  G38,
  G39,
  G40,
  G41,
  G1324,
  G1325,
  G1326,
  G1327,
  G1328,
  G1329,
  G1330,
  G1331,
  G1332,
  G1333,
  G1334,
  G1335,
  G1336,
  G1337,
  G1338,
  G1339,
  G1340,
  G1341,
  G1342,
  G1343,
  G1344,
  G1345,
  G1346,
  G1347,
  G1348,
  G1349,
  G1350,
  G1351,
  G1352,
  G1353,
  G1354,
  G1355
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;input G33;input G34;input G35;input G36;input G37;input G38;input G39;input G40;input G41;
  output G1324;output G1325;output G1326;output G1327;output G1328;output G1329;output G1330;output G1331;output G1332;output G1333;output G1334;output G1335;output G1336;output G1337;output G1338;output G1339;output G1340;output G1341;output G1342;output G1343;output G1344;output G1345;output G1346;output G1347;output G1348;output G1349;output G1350;output G1351;output G1352;output G1353;output G1354;output G1355;
  wire new_n74_;wire new_n75_;wire new_n76_;wire new_n77_;wire new_n78_;wire new_n79_;wire new_n80_;wire new_n81_;wire new_n82_;wire new_n83_;wire new_n84_;wire new_n85_;wire new_n86_;wire new_n87_;wire new_n88_;wire new_n89_;wire new_n90_;wire new_n91_;wire new_n92_;wire new_n93_;wire new_n94_;wire new_n95_;wire new_n96_;wire new_n97_;wire new_n98_;wire new_n99_;wire new_n100_;wire new_n101_;wire new_n102_;wire new_n103_;wire new_n104_;wire new_n105_;wire new_n106_;wire new_n107_;wire new_n108_;wire new_n109_;wire new_n110_;wire new_n111_;wire new_n112_;wire new_n113_;wire new_n114_;wire new_n115_;wire new_n116_;wire new_n117_;wire new_n118_;wire new_n119_;wire new_n120_;wire new_n121_;wire new_n122_;wire new_n123_;wire new_n124_;wire new_n125_;wire new_n126_;wire new_n127_;wire new_n128_;wire new_n129_;wire new_n130_;wire new_n131_;wire new_n132_;wire new_n133_;wire new_n134_;wire new_n135_;wire new_n136_;wire new_n137_;wire new_n138_;wire new_n139_;wire new_n140_;wire new_n141_;wire new_n142_;wire new_n143_;wire new_n144_;wire new_n145_;wire new_n146_;wire new_n147_;wire new_n148_;wire new_n149_;wire new_n150_;wire new_n151_;wire new_n152_;wire new_n153_;wire new_n154_;wire new_n155_;wire new_n156_;wire new_n157_;wire new_n158_;wire new_n159_;wire new_n160_;wire new_n161_;wire new_n162_;wire new_n163_;wire new_n164_;wire new_n165_;wire new_n166_;wire new_n167_;wire new_n168_;wire new_n169_;wire new_n170_;wire new_n171_;wire new_n172_;wire new_n173_;wire new_n174_;wire new_n175_;wire new_n176_;wire new_n177_;wire new_n178_;wire new_n179_;wire new_n180_;wire new_n181_;wire new_n182_;wire new_n183_;wire new_n184_;wire new_n185_;wire new_n186_;wire new_n187_;wire new_n188_;wire new_n189_;wire new_n190_;wire new_n191_;wire new_n192_;wire new_n193_;wire new_n194_;wire new_n195_;wire new_n196_;wire new_n197_;wire new_n198_;wire new_n199_;wire new_n200_;wire new_n201_;wire new_n202_;wire new_n203_;wire new_n204_;wire new_n205_;wire new_n206_;wire new_n207_;wire new_n208_;wire new_n209_;wire new_n210_;wire new_n211_;wire new_n212_;wire new_n213_;wire new_n214_;wire new_n215_;wire new_n216_;wire new_n217_;wire new_n218_;wire new_n219_;wire new_n220_;wire new_n221_;wire new_n222_;wire new_n223_;wire new_n224_;wire new_n225_;wire new_n226_;wire new_n227_;wire new_n228_;wire new_n229_;wire new_n230_;wire new_n231_;wire new_n232_;wire new_n233_;wire new_n234_;wire new_n235_;wire new_n236_;wire new_n237_;wire new_n238_;wire new_n239_;wire new_n240_;wire new_n241_;wire new_n242_;wire new_n243_;wire new_n244_;wire new_n245_;wire new_n246_;wire new_n247_;wire new_n248_;wire new_n249_;wire new_n250_;wire new_n251_;wire new_n252_;wire new_n253_;wire new_n254_;wire new_n255_;wire new_n256_;wire new_n257_;wire new_n258_;wire new_n259_;wire new_n260_;wire new_n261_;wire new_n262_;wire new_n263_;wire new_n264_;wire new_n265_;wire new_n266_;wire new_n267_;wire new_n268_;wire new_n269_;wire new_n270_;wire new_n271_;wire new_n272_;wire new_n273_;wire new_n274_;wire new_n275_;wire new_n276_;wire new_n277_;wire new_n278_;wire new_n279_;wire new_n280_;wire new_n281_;wire new_n282_;wire new_n283_;wire new_n284_;wire new_n285_;wire new_n286_;wire new_n287_;wire new_n288_;wire new_n289_;wire new_n290_;wire new_n291_;wire new_n292_;wire new_n293_;wire new_n294_;wire new_n295_;wire new_n296_;wire new_n297_;wire new_n298_;wire new_n299_;wire new_n300_;wire new_n301_;wire new_n302_;wire new_n303_;wire new_n304_;wire new_n305_;wire new_n306_;wire new_n307_;wire new_n308_;wire new_n309_;wire new_n310_;wire new_n311_;wire new_n312_;wire new_n313_;wire new_n314_;wire new_n315_;wire new_n316_;wire new_n318_;wire new_n319_;wire new_n320_;wire new_n322_;wire new_n323_;wire new_n324_;wire new_n326_;wire new_n327_;wire new_n328_;wire new_n330_;wire new_n331_;wire new_n332_;wire new_n333_;wire new_n334_;wire new_n335_;wire new_n337_;wire new_n338_;wire new_n339_;wire new_n341_;wire new_n342_;wire new_n343_;wire new_n345_;wire new_n346_;wire new_n347_;wire new_n349_;wire new_n350_;wire new_n351_;wire new_n352_;wire new_n353_;wire new_n355_;wire new_n356_;wire new_n357_;wire new_n359_;wire new_n360_;wire new_n361_;wire new_n363_;wire new_n364_;wire new_n365_;wire new_n367_;wire new_n368_;wire new_n369_;wire new_n370_;wire new_n371_;wire new_n373_;wire new_n374_;wire new_n375_;wire new_n377_;wire new_n378_;wire new_n379_;wire new_n381_;wire new_n382_;wire new_n383_;wire new_n385_;wire new_n386_;wire new_n387_;wire new_n388_;wire new_n389_;wire new_n390_;wire new_n391_;wire new_n392_;wire new_n393_;wire new_n394_;wire new_n395_;wire new_n396_;wire new_n398_;wire new_n399_;wire new_n400_;wire new_n402_;wire new_n403_;wire new_n404_;wire new_n406_;wire new_n407_;wire new_n408_;wire new_n410_;wire new_n411_;wire new_n412_;wire new_n413_;wire new_n414_;wire new_n416_;wire new_n417_;wire new_n418_;wire new_n420_;wire new_n421_;wire new_n422_;wire new_n424_;wire new_n425_;wire new_n426_;wire new_n428_;wire new_n429_;wire new_n430_;wire new_n431_;wire new_n432_;wire new_n434_;wire new_n435_;wire new_n436_;wire new_n438_;wire new_n439_;wire new_n440_;wire new_n442_;wire new_n443_;wire new_n444_;wire new_n446_;wire new_n447_;wire new_n448_;wire new_n449_;wire new_n451_;wire new_n452_;wire new_n453_;wire new_n455_;wire new_n456_;wire new_n457_;wire new_n459_;wire new_n460_;wire new_n461_;
  wire G13_spl_;
  wire G13_spl_0;
  wire G13_spl_00;
  wire G13_spl_01;
  wire G13_spl_1;
  wire G9_spl_;
  wire G9_spl_0;
  wire G9_spl_00;
  wire G9_spl_01;
  wire G9_spl_1;
  wire G1_spl_;
  wire G1_spl_0;
  wire G1_spl_00;
  wire G1_spl_01;
  wire G1_spl_1;
  wire G5_spl_;
  wire G5_spl_0;
  wire G5_spl_00;
  wire G5_spl_01;
  wire G5_spl_1;
  wire new_n76__spl_;
  wire new_n79__spl_;
  wire G41_spl_;
  wire G41_spl_0;
  wire G41_spl_00;
  wire G41_spl_01;
  wire G41_spl_1;
  wire G41_spl_10;
  wire G41_spl_11;
  wire new_n82__spl_;
  wire new_n83__spl_;
  wire G20_spl_;
  wire G20_spl_0;
  wire G20_spl_00;
  wire G20_spl_01;
  wire G20_spl_1;
  wire G19_spl_;
  wire G19_spl_0;
  wire G19_spl_00;
  wire G19_spl_01;
  wire G19_spl_1;
  wire G17_spl_;
  wire G17_spl_0;
  wire G17_spl_00;
  wire G17_spl_01;
  wire G17_spl_1;
  wire G18_spl_;
  wire G18_spl_0;
  wire G18_spl_00;
  wire G18_spl_01;
  wire G18_spl_1;
  wire new_n89__spl_;
  wire new_n92__spl_;
  wire G24_spl_;
  wire G24_spl_0;
  wire G24_spl_00;
  wire G24_spl_01;
  wire G24_spl_1;
  wire G23_spl_;
  wire G23_spl_0;
  wire G23_spl_00;
  wire G23_spl_01;
  wire G23_spl_1;
  wire G21_spl_;
  wire G21_spl_0;
  wire G21_spl_00;
  wire G21_spl_01;
  wire G21_spl_1;
  wire G22_spl_;
  wire G22_spl_0;
  wire G22_spl_00;
  wire G22_spl_01;
  wire G22_spl_1;
  wire new_n98__spl_;
  wire new_n101__spl_;
  wire new_n95__spl_;
  wire new_n95__spl_0;
  wire new_n95__spl_1;
  wire new_n104__spl_;
  wire new_n104__spl_0;
  wire new_n104__spl_1;
  wire new_n86__spl_;
  wire new_n107__spl_;
  wire G29_spl_;
  wire G29_spl_0;
  wire G29_spl_00;
  wire G29_spl_01;
  wire G29_spl_1;
  wire G25_spl_;
  wire G25_spl_0;
  wire G25_spl_00;
  wire G25_spl_01;
  wire G25_spl_1;
  wire new_n113__spl_;
  wire new_n116__spl_;
  wire new_n119__spl_;
  wire new_n120__spl_;
  wire G8_spl_;
  wire G8_spl_0;
  wire G8_spl_00;
  wire G8_spl_01;
  wire G8_spl_1;
  wire G7_spl_;
  wire G7_spl_0;
  wire G7_spl_00;
  wire G7_spl_01;
  wire G7_spl_1;
  wire G6_spl_;
  wire G6_spl_0;
  wire G6_spl_00;
  wire G6_spl_01;
  wire G6_spl_1;
  wire new_n126__spl_;
  wire new_n129__spl_;
  wire G4_spl_;
  wire G4_spl_0;
  wire G4_spl_00;
  wire G4_spl_01;
  wire G4_spl_1;
  wire G3_spl_;
  wire G3_spl_0;
  wire G3_spl_00;
  wire G3_spl_01;
  wire G3_spl_1;
  wire G2_spl_;
  wire G2_spl_0;
  wire G2_spl_00;
  wire G2_spl_01;
  wire G2_spl_1;
  wire new_n135__spl_;
  wire new_n138__spl_;
  wire new_n132__spl_;
  wire new_n132__spl_0;
  wire new_n132__spl_1;
  wire new_n141__spl_;
  wire new_n141__spl_0;
  wire new_n141__spl_1;
  wire new_n123__spl_;
  wire new_n144__spl_;
  wire G30_spl_;
  wire G30_spl_0;
  wire G30_spl_00;
  wire G30_spl_01;
  wire G30_spl_1;
  wire G26_spl_;
  wire G26_spl_0;
  wire G26_spl_00;
  wire G26_spl_01;
  wire G26_spl_1;
  wire new_n150__spl_;
  wire new_n153__spl_;
  wire new_n156__spl_;
  wire new_n157__spl_;
  wire G16_spl_;
  wire G16_spl_0;
  wire G16_spl_00;
  wire G16_spl_01;
  wire G16_spl_1;
  wire G15_spl_;
  wire G15_spl_0;
  wire G15_spl_00;
  wire G15_spl_01;
  wire G15_spl_1;
  wire G14_spl_;
  wire G14_spl_0;
  wire G14_spl_00;
  wire G14_spl_01;
  wire G14_spl_1;
  wire new_n163__spl_;
  wire new_n166__spl_;
  wire G12_spl_;
  wire G12_spl_0;
  wire G12_spl_00;
  wire G12_spl_01;
  wire G12_spl_1;
  wire G11_spl_;
  wire G11_spl_0;
  wire G11_spl_00;
  wire G11_spl_01;
  wire G11_spl_1;
  wire G10_spl_;
  wire G10_spl_0;
  wire G10_spl_00;
  wire G10_spl_01;
  wire G10_spl_1;
  wire new_n172__spl_;
  wire new_n175__spl_;
  wire new_n169__spl_;
  wire new_n169__spl_0;
  wire new_n169__spl_1;
  wire new_n178__spl_;
  wire new_n178__spl_0;
  wire new_n178__spl_1;
  wire new_n160__spl_;
  wire new_n181__spl_;
  wire new_n184__spl_;
  wire new_n184__spl_0;
  wire new_n184__spl_00;
  wire new_n184__spl_01;
  wire new_n184__spl_1;
  wire new_n184__spl_10;
  wire new_n147__spl_;
  wire new_n147__spl_0;
  wire new_n147__spl_00;
  wire new_n147__spl_01;
  wire new_n147__spl_1;
  wire new_n147__spl_10;
  wire G32_spl_;
  wire G32_spl_0;
  wire G32_spl_00;
  wire G32_spl_01;
  wire G32_spl_1;
  wire G28_spl_;
  wire G28_spl_0;
  wire G28_spl_00;
  wire G28_spl_01;
  wire G28_spl_1;
  wire new_n188__spl_;
  wire new_n191__spl_;
  wire new_n194__spl_;
  wire new_n195__spl_;
  wire new_n198__spl_;
  wire new_n201__spl_;
  wire G31_spl_;
  wire G31_spl_0;
  wire G31_spl_00;
  wire G31_spl_01;
  wire G31_spl_1;
  wire G27_spl_;
  wire G27_spl_0;
  wire G27_spl_00;
  wire G27_spl_01;
  wire G27_spl_1;
  wire new_n207__spl_;
  wire new_n210__spl_;
  wire new_n213__spl_;
  wire new_n214__spl_;
  wire new_n217__spl_;
  wire new_n220__spl_;
  wire new_n223__spl_;
  wire new_n223__spl_0;
  wire new_n223__spl_00;
  wire new_n223__spl_01;
  wire new_n223__spl_1;
  wire new_n223__spl_10;
  wire new_n223__spl_11;
  wire new_n204__spl_;
  wire new_n204__spl_0;
  wire new_n204__spl_00;
  wire new_n204__spl_01;
  wire new_n204__spl_1;
  wire new_n204__spl_10;
  wire new_n204__spl_11;
  wire new_n227__spl_;
  wire new_n230__spl_;
  wire new_n233__spl_;
  wire new_n234__spl_;
  wire new_n240__spl_;
  wire new_n243__spl_;
  wire new_n246__spl_;
  wire new_n246__spl_0;
  wire new_n246__spl_1;
  wire new_n237__spl_;
  wire new_n249__spl_;
  wire new_n255__spl_;
  wire new_n258__spl_;
  wire new_n261__spl_;
  wire new_n262__spl_;
  wire new_n268__spl_;
  wire new_n271__spl_;
  wire new_n274__spl_;
  wire new_n274__spl_0;
  wire new_n274__spl_1;
  wire new_n265__spl_;
  wire new_n277__spl_;
  wire new_n283__spl_;
  wire new_n286__spl_;
  wire new_n289__spl_;
  wire new_n290__spl_;
  wire new_n293__spl_;
  wire new_n296__spl_;
  wire new_n110__spl_;
  wire new_n110__spl_0;
  wire new_n110__spl_00;
  wire new_n110__spl_01;
  wire new_n110__spl_1;
  wire new_n110__spl_10;
  wire new_n299__spl_;
  wire new_n299__spl_0;
  wire new_n299__spl_00;
  wire new_n299__spl_01;
  wire new_n299__spl_1;
  wire new_n299__spl_10;
  wire new_n280__spl_;
  wire new_n280__spl_0;
  wire new_n280__spl_00;
  wire new_n280__spl_01;
  wire new_n280__spl_1;
  wire new_n280__spl_10;
  wire new_n280__spl_11;
  wire new_n300__spl_;
  wire new_n302__spl_;
  wire new_n301__spl_;
  wire new_n303__spl_;
  wire new_n252__spl_;
  wire new_n252__spl_0;
  wire new_n252__spl_00;
  wire new_n252__spl_01;
  wire new_n252__spl_1;
  wire new_n252__spl_10;
  wire new_n252__spl_11;
  wire new_n306__spl_;
  wire new_n306__spl_0;
  wire new_n224__spl_;
  wire new_n311__spl_;
  wire new_n185__spl_;
  wire new_n312__spl_;
  wire new_n313__spl_;
  wire new_n313__spl_0;
  wire new_n313__spl_1;
  wire new_n314__spl_;
  wire new_n318__spl_;
  wire new_n322__spl_;
  wire new_n326__spl_;
  wire new_n330__spl_;
  wire new_n331__spl_;
  wire new_n332__spl_;
  wire new_n332__spl_0;
  wire new_n332__spl_1;
  wire new_n333__spl_;
  wire new_n337__spl_;
  wire new_n341__spl_;
  wire new_n345__spl_;
  wire new_n349__spl_;
  wire new_n350__spl_;
  wire new_n350__spl_0;
  wire new_n350__spl_1;
  wire new_n351__spl_;
  wire new_n355__spl_;
  wire new_n359__spl_;
  wire new_n363__spl_;
  wire new_n367__spl_;
  wire new_n368__spl_;
  wire new_n368__spl_0;
  wire new_n368__spl_1;
  wire new_n369__spl_;
  wire new_n373__spl_;
  wire new_n377__spl_;
  wire new_n381__spl_;
  wire new_n391__spl_;
  wire new_n391__spl_0;
  wire new_n393__spl_;
  wire new_n393__spl_0;
  wire new_n393__spl_1;
  wire new_n394__spl_;
  wire new_n398__spl_;
  wire new_n402__spl_;
  wire new_n406__spl_;
  wire new_n410__spl_;
  wire new_n411__spl_;
  wire new_n411__spl_0;
  wire new_n411__spl_1;
  wire new_n412__spl_;
  wire new_n416__spl_;
  wire new_n420__spl_;
  wire new_n424__spl_;
  wire new_n429__spl_;
  wire new_n429__spl_0;
  wire new_n429__spl_1;
  wire new_n430__spl_;
  wire new_n434__spl_;
  wire new_n438__spl_;
  wire new_n442__spl_;
  wire new_n446__spl_;
  wire new_n446__spl_0;
  wire new_n446__spl_1;
  wire new_n447__spl_;
  wire new_n451__spl_;
  wire new_n455__spl_;
  wire new_n459__spl_;

  anb2
  g000
  (
    .dina(G13_spl_00),
    .dinb(G9_spl_00),
    .dout(new_n74_)
  );


  anb1
  g001
  (
    .dina(G13_spl_00),
    .dinb(G9_spl_00),
    .dout(new_n75_)
  );


  anb1
  g002
  (
    .dina(new_n74_),
    .dinb(new_n75_),
    .dout(new_n76_)
  );


  nor1
  g003
  (
    .dina(G1_spl_00),
    .dinb(G5_spl_00),
    .dout(new_n77_)
  );


  nor2
  g004
  (
    .dina(G1_spl_00),
    .dinb(G5_spl_00),
    .dout(new_n78_)
  );


  anb2
  g005
  (
    .dina(new_n77_),
    .dinb(new_n78_),
    .dout(new_n79_)
  );


  anb1
  g006
  (
    .dina(new_n76__spl_),
    .dinb(new_n79__spl_),
    .dout(new_n80_)
  );


  anb2
  g007
  (
    .dina(new_n76__spl_),
    .dinb(new_n79__spl_),
    .dout(new_n81_)
  );


  anb2
  g008
  (
    .dina(new_n80_),
    .dinb(new_n81_),
    .dout(new_n82_)
  );


  nor2
  g009
  (
    .dina(G33),
    .dinb(G41_spl_00),
    .dout(new_n83_)
  );


  anb1
  g010
  (
    .dina(new_n82__spl_),
    .dinb(new_n83__spl_),
    .dout(new_n84_)
  );


  anb2
  g011
  (
    .dina(new_n82__spl_),
    .dinb(new_n83__spl_),
    .dout(new_n85_)
  );


  anb2
  g012
  (
    .dina(new_n84_),
    .dinb(new_n85_),
    .dout(new_n86_)
  );


  anb2
  g013
  (
    .dina(G20_spl_00),
    .dinb(G19_spl_00),
    .dout(new_n87_)
  );


  anb1
  g014
  (
    .dina(G20_spl_00),
    .dinb(G19_spl_00),
    .dout(new_n88_)
  );


  anb1
  g015
  (
    .dina(new_n87_),
    .dinb(new_n88_),
    .dout(new_n89_)
  );


  nor1
  g016
  (
    .dina(G17_spl_00),
    .dinb(G18_spl_00),
    .dout(new_n90_)
  );


  nor2
  g017
  (
    .dina(G17_spl_00),
    .dinb(G18_spl_00),
    .dout(new_n91_)
  );


  anb2
  g018
  (
    .dina(new_n90_),
    .dinb(new_n91_),
    .dout(new_n92_)
  );


  anb1
  g019
  (
    .dina(new_n89__spl_),
    .dinb(new_n92__spl_),
    .dout(new_n93_)
  );


  anb2
  g020
  (
    .dina(new_n89__spl_),
    .dinb(new_n92__spl_),
    .dout(new_n94_)
  );


  anb2
  g021
  (
    .dina(new_n93_),
    .dinb(new_n94_),
    .dout(new_n95_)
  );


  anb2
  g022
  (
    .dina(G24_spl_00),
    .dinb(G23_spl_00),
    .dout(new_n96_)
  );


  anb1
  g023
  (
    .dina(G24_spl_00),
    .dinb(G23_spl_00),
    .dout(new_n97_)
  );


  anb1
  g024
  (
    .dina(new_n96_),
    .dinb(new_n97_),
    .dout(new_n98_)
  );


  nor1
  g025
  (
    .dina(G21_spl_00),
    .dinb(G22_spl_00),
    .dout(new_n99_)
  );


  nor2
  g026
  (
    .dina(G21_spl_00),
    .dinb(G22_spl_00),
    .dout(new_n100_)
  );


  anb2
  g027
  (
    .dina(new_n99_),
    .dinb(new_n100_),
    .dout(new_n101_)
  );


  anb1
  g028
  (
    .dina(new_n98__spl_),
    .dinb(new_n101__spl_),
    .dout(new_n102_)
  );


  anb2
  g029
  (
    .dina(new_n98__spl_),
    .dinb(new_n101__spl_),
    .dout(new_n103_)
  );


  anb2
  g030
  (
    .dina(new_n102_),
    .dinb(new_n103_),
    .dout(new_n104_)
  );


  anb2
  g031
  (
    .dina(new_n95__spl_0),
    .dinb(new_n104__spl_0),
    .dout(new_n105_)
  );


  anb1
  g032
  (
    .dina(new_n95__spl_0),
    .dinb(new_n104__spl_0),
    .dout(new_n106_)
  );


  anb1
  g033
  (
    .dina(new_n105_),
    .dinb(new_n106_),
    .dout(new_n107_)
  );


  anb1
  g034
  (
    .dina(new_n86__spl_),
    .dinb(new_n107__spl_),
    .dout(new_n108_)
  );


  anb2
  g035
  (
    .dina(new_n86__spl_),
    .dinb(new_n107__spl_),
    .dout(new_n109_)
  );


  anb2
  g036
  (
    .dina(new_n108_),
    .dinb(new_n109_),
    .dout(new_n110_)
  );


  anb2
  g037
  (
    .dina(G29_spl_00),
    .dinb(G25_spl_00),
    .dout(new_n111_)
  );


  anb1
  g038
  (
    .dina(G29_spl_00),
    .dinb(G25_spl_00),
    .dout(new_n112_)
  );


  anb1
  g039
  (
    .dina(new_n111_),
    .dinb(new_n112_),
    .dout(new_n113_)
  );


  nor1
  g040
  (
    .dina(G17_spl_01),
    .dinb(G21_spl_01),
    .dout(new_n114_)
  );


  nor2
  g041
  (
    .dina(G17_spl_01),
    .dinb(G21_spl_01),
    .dout(new_n115_)
  );


  anb2
  g042
  (
    .dina(new_n114_),
    .dinb(new_n115_),
    .dout(new_n116_)
  );


  anb1
  g043
  (
    .dina(new_n113__spl_),
    .dinb(new_n116__spl_),
    .dout(new_n117_)
  );


  anb2
  g044
  (
    .dina(new_n113__spl_),
    .dinb(new_n116__spl_),
    .dout(new_n118_)
  );


  anb2
  g045
  (
    .dina(new_n117_),
    .dinb(new_n118_),
    .dout(new_n119_)
  );


  nor2
  g046
  (
    .dina(G37),
    .dinb(G41_spl_00),
    .dout(new_n120_)
  );


  anb1
  g047
  (
    .dina(new_n119__spl_),
    .dinb(new_n120__spl_),
    .dout(new_n121_)
  );


  anb2
  g048
  (
    .dina(new_n119__spl_),
    .dinb(new_n120__spl_),
    .dout(new_n122_)
  );


  anb2
  g049
  (
    .dina(new_n121_),
    .dinb(new_n122_),
    .dout(new_n123_)
  );


  anb2
  g050
  (
    .dina(G8_spl_00),
    .dinb(G7_spl_00),
    .dout(new_n124_)
  );


  anb1
  g051
  (
    .dina(G8_spl_00),
    .dinb(G7_spl_00),
    .dout(new_n125_)
  );


  anb1
  g052
  (
    .dina(new_n124_),
    .dinb(new_n125_),
    .dout(new_n126_)
  );


  nor1
  g053
  (
    .dina(G5_spl_01),
    .dinb(G6_spl_00),
    .dout(new_n127_)
  );


  nor2
  g054
  (
    .dina(G5_spl_01),
    .dinb(G6_spl_00),
    .dout(new_n128_)
  );


  anb2
  g055
  (
    .dina(new_n127_),
    .dinb(new_n128_),
    .dout(new_n129_)
  );


  anb1
  g056
  (
    .dina(new_n126__spl_),
    .dinb(new_n129__spl_),
    .dout(new_n130_)
  );


  anb2
  g057
  (
    .dina(new_n126__spl_),
    .dinb(new_n129__spl_),
    .dout(new_n131_)
  );


  anb2
  g058
  (
    .dina(new_n130_),
    .dinb(new_n131_),
    .dout(new_n132_)
  );


  anb2
  g059
  (
    .dina(G4_spl_00),
    .dinb(G3_spl_00),
    .dout(new_n133_)
  );


  anb1
  g060
  (
    .dina(G4_spl_00),
    .dinb(G3_spl_00),
    .dout(new_n134_)
  );


  anb1
  g061
  (
    .dina(new_n133_),
    .dinb(new_n134_),
    .dout(new_n135_)
  );


  nor1
  g062
  (
    .dina(G1_spl_01),
    .dinb(G2_spl_00),
    .dout(new_n136_)
  );


  nor2
  g063
  (
    .dina(G1_spl_01),
    .dinb(G2_spl_00),
    .dout(new_n137_)
  );


  anb2
  g064
  (
    .dina(new_n136_),
    .dinb(new_n137_),
    .dout(new_n138_)
  );


  anb1
  g065
  (
    .dina(new_n135__spl_),
    .dinb(new_n138__spl_),
    .dout(new_n139_)
  );


  anb2
  g066
  (
    .dina(new_n135__spl_),
    .dinb(new_n138__spl_),
    .dout(new_n140_)
  );


  anb2
  g067
  (
    .dina(new_n139_),
    .dinb(new_n140_),
    .dout(new_n141_)
  );


  anb2
  g068
  (
    .dina(new_n132__spl_0),
    .dinb(new_n141__spl_0),
    .dout(new_n142_)
  );


  anb1
  g069
  (
    .dina(new_n132__spl_0),
    .dinb(new_n141__spl_0),
    .dout(new_n143_)
  );


  anb1
  g070
  (
    .dina(new_n142_),
    .dinb(new_n143_),
    .dout(new_n144_)
  );


  anb1
  g071
  (
    .dina(new_n123__spl_),
    .dinb(new_n144__spl_),
    .dout(new_n145_)
  );


  anb2
  g072
  (
    .dina(new_n123__spl_),
    .dinb(new_n144__spl_),
    .dout(new_n146_)
  );


  anb2
  g073
  (
    .dina(new_n145_),
    .dinb(new_n146_),
    .dout(new_n147_)
  );


  anb2
  g074
  (
    .dina(G30_spl_00),
    .dinb(G26_spl_00),
    .dout(new_n148_)
  );


  anb1
  g075
  (
    .dina(G30_spl_00),
    .dinb(G26_spl_00),
    .dout(new_n149_)
  );


  anb1
  g076
  (
    .dina(new_n148_),
    .dinb(new_n149_),
    .dout(new_n150_)
  );


  nor1
  g077
  (
    .dina(G18_spl_01),
    .dinb(G22_spl_01),
    .dout(new_n151_)
  );


  nor2
  g078
  (
    .dina(G18_spl_01),
    .dinb(G22_spl_01),
    .dout(new_n152_)
  );


  anb2
  g079
  (
    .dina(new_n151_),
    .dinb(new_n152_),
    .dout(new_n153_)
  );


  anb1
  g080
  (
    .dina(new_n150__spl_),
    .dinb(new_n153__spl_),
    .dout(new_n154_)
  );


  anb2
  g081
  (
    .dina(new_n150__spl_),
    .dinb(new_n153__spl_),
    .dout(new_n155_)
  );


  anb2
  g082
  (
    .dina(new_n154_),
    .dinb(new_n155_),
    .dout(new_n156_)
  );


  nor2
  g083
  (
    .dina(G38),
    .dinb(G41_spl_01),
    .dout(new_n157_)
  );


  anb1
  g084
  (
    .dina(new_n156__spl_),
    .dinb(new_n157__spl_),
    .dout(new_n158_)
  );


  anb2
  g085
  (
    .dina(new_n156__spl_),
    .dinb(new_n157__spl_),
    .dout(new_n159_)
  );


  anb2
  g086
  (
    .dina(new_n158_),
    .dinb(new_n159_),
    .dout(new_n160_)
  );


  anb2
  g087
  (
    .dina(G16_spl_00),
    .dinb(G15_spl_00),
    .dout(new_n161_)
  );


  anb1
  g088
  (
    .dina(G16_spl_00),
    .dinb(G15_spl_00),
    .dout(new_n162_)
  );


  anb1
  g089
  (
    .dina(new_n161_),
    .dinb(new_n162_),
    .dout(new_n163_)
  );


  nor1
  g090
  (
    .dina(G13_spl_01),
    .dinb(G14_spl_00),
    .dout(new_n164_)
  );


  nor2
  g091
  (
    .dina(G13_spl_01),
    .dinb(G14_spl_00),
    .dout(new_n165_)
  );


  anb2
  g092
  (
    .dina(new_n164_),
    .dinb(new_n165_),
    .dout(new_n166_)
  );


  anb1
  g093
  (
    .dina(new_n163__spl_),
    .dinb(new_n166__spl_),
    .dout(new_n167_)
  );


  anb2
  g094
  (
    .dina(new_n163__spl_),
    .dinb(new_n166__spl_),
    .dout(new_n168_)
  );


  anb2
  g095
  (
    .dina(new_n167_),
    .dinb(new_n168_),
    .dout(new_n169_)
  );


  anb2
  g096
  (
    .dina(G12_spl_00),
    .dinb(G11_spl_00),
    .dout(new_n170_)
  );


  anb1
  g097
  (
    .dina(G12_spl_00),
    .dinb(G11_spl_00),
    .dout(new_n171_)
  );


  anb1
  g098
  (
    .dina(new_n170_),
    .dinb(new_n171_),
    .dout(new_n172_)
  );


  nor1
  g099
  (
    .dina(G9_spl_01),
    .dinb(G10_spl_00),
    .dout(new_n173_)
  );


  nor2
  g100
  (
    .dina(G9_spl_01),
    .dinb(G10_spl_00),
    .dout(new_n174_)
  );


  anb2
  g101
  (
    .dina(new_n173_),
    .dinb(new_n174_),
    .dout(new_n175_)
  );


  anb1
  g102
  (
    .dina(new_n172__spl_),
    .dinb(new_n175__spl_),
    .dout(new_n176_)
  );


  anb2
  g103
  (
    .dina(new_n172__spl_),
    .dinb(new_n175__spl_),
    .dout(new_n177_)
  );


  anb2
  g104
  (
    .dina(new_n176_),
    .dinb(new_n177_),
    .dout(new_n178_)
  );


  anb2
  g105
  (
    .dina(new_n169__spl_0),
    .dinb(new_n178__spl_0),
    .dout(new_n179_)
  );


  anb1
  g106
  (
    .dina(new_n169__spl_0),
    .dinb(new_n178__spl_0),
    .dout(new_n180_)
  );


  anb1
  g107
  (
    .dina(new_n179_),
    .dinb(new_n180_),
    .dout(new_n181_)
  );


  anb1
  g108
  (
    .dina(new_n160__spl_),
    .dinb(new_n181__spl_),
    .dout(new_n182_)
  );


  anb2
  g109
  (
    .dina(new_n160__spl_),
    .dinb(new_n181__spl_),
    .dout(new_n183_)
  );


  anb2
  g110
  (
    .dina(new_n182_),
    .dinb(new_n183_),
    .dout(new_n184_)
  );


  anb2
  g111
  (
    .dina(new_n184__spl_00),
    .dinb(new_n147__spl_00),
    .dout(new_n185_)
  );


  anb2
  g112
  (
    .dina(G32_spl_00),
    .dinb(G28_spl_00),
    .dout(new_n186_)
  );


  anb1
  g113
  (
    .dina(G32_spl_00),
    .dinb(G28_spl_00),
    .dout(new_n187_)
  );


  anb1
  g114
  (
    .dina(new_n186_),
    .dinb(new_n187_),
    .dout(new_n188_)
  );


  nor1
  g115
  (
    .dina(G20_spl_01),
    .dinb(G24_spl_01),
    .dout(new_n189_)
  );


  nor2
  g116
  (
    .dina(G20_spl_01),
    .dinb(G24_spl_01),
    .dout(new_n190_)
  );


  anb2
  g117
  (
    .dina(new_n189_),
    .dinb(new_n190_),
    .dout(new_n191_)
  );


  anb1
  g118
  (
    .dina(new_n188__spl_),
    .dinb(new_n191__spl_),
    .dout(new_n192_)
  );


  anb2
  g119
  (
    .dina(new_n188__spl_),
    .dinb(new_n191__spl_),
    .dout(new_n193_)
  );


  anb2
  g120
  (
    .dina(new_n192_),
    .dinb(new_n193_),
    .dout(new_n194_)
  );


  nor2
  g121
  (
    .dina(G40),
    .dinb(G41_spl_01),
    .dout(new_n195_)
  );


  anb1
  g122
  (
    .dina(new_n194__spl_),
    .dinb(new_n195__spl_),
    .dout(new_n196_)
  );


  anb2
  g123
  (
    .dina(new_n194__spl_),
    .dinb(new_n195__spl_),
    .dout(new_n197_)
  );


  anb2
  g124
  (
    .dina(new_n196_),
    .dinb(new_n197_),
    .dout(new_n198_)
  );


  anb2
  g125
  (
    .dina(new_n132__spl_1),
    .dinb(new_n169__spl_1),
    .dout(new_n199_)
  );


  anb1
  g126
  (
    .dina(new_n132__spl_1),
    .dinb(new_n169__spl_1),
    .dout(new_n200_)
  );


  anb1
  g127
  (
    .dina(new_n199_),
    .dinb(new_n200_),
    .dout(new_n201_)
  );


  anb1
  g128
  (
    .dina(new_n198__spl_),
    .dinb(new_n201__spl_),
    .dout(new_n202_)
  );


  anb2
  g129
  (
    .dina(new_n198__spl_),
    .dinb(new_n201__spl_),
    .dout(new_n203_)
  );


  anb2
  g130
  (
    .dina(new_n202_),
    .dinb(new_n203_),
    .dout(new_n204_)
  );


  anb2
  g131
  (
    .dina(G31_spl_00),
    .dinb(G27_spl_00),
    .dout(new_n205_)
  );


  anb1
  g132
  (
    .dina(G31_spl_00),
    .dinb(G27_spl_00),
    .dout(new_n206_)
  );


  anb1
  g133
  (
    .dina(new_n205_),
    .dinb(new_n206_),
    .dout(new_n207_)
  );


  nor1
  g134
  (
    .dina(G19_spl_01),
    .dinb(G23_spl_01),
    .dout(new_n208_)
  );


  nor2
  g135
  (
    .dina(G19_spl_01),
    .dinb(G23_spl_01),
    .dout(new_n209_)
  );


  anb2
  g136
  (
    .dina(new_n208_),
    .dinb(new_n209_),
    .dout(new_n210_)
  );


  anb1
  g137
  (
    .dina(new_n207__spl_),
    .dinb(new_n210__spl_),
    .dout(new_n211_)
  );


  anb2
  g138
  (
    .dina(new_n207__spl_),
    .dinb(new_n210__spl_),
    .dout(new_n212_)
  );


  anb2
  g139
  (
    .dina(new_n211_),
    .dinb(new_n212_),
    .dout(new_n213_)
  );


  nor2
  g140
  (
    .dina(G39),
    .dinb(G41_spl_10),
    .dout(new_n214_)
  );


  anb1
  g141
  (
    .dina(new_n213__spl_),
    .dinb(new_n214__spl_),
    .dout(new_n215_)
  );


  anb2
  g142
  (
    .dina(new_n213__spl_),
    .dinb(new_n214__spl_),
    .dout(new_n216_)
  );


  anb2
  g143
  (
    .dina(new_n215_),
    .dinb(new_n216_),
    .dout(new_n217_)
  );


  anb2
  g144
  (
    .dina(new_n141__spl_1),
    .dinb(new_n178__spl_1),
    .dout(new_n218_)
  );


  anb1
  g145
  (
    .dina(new_n141__spl_1),
    .dinb(new_n178__spl_1),
    .dout(new_n219_)
  );


  anb1
  g146
  (
    .dina(new_n218_),
    .dinb(new_n219_),
    .dout(new_n220_)
  );


  anb1
  g147
  (
    .dina(new_n217__spl_),
    .dinb(new_n220__spl_),
    .dout(new_n221_)
  );


  anb2
  g148
  (
    .dina(new_n217__spl_),
    .dinb(new_n220__spl_),
    .dout(new_n222_)
  );


  anb2
  g149
  (
    .dina(new_n221_),
    .dinb(new_n222_),
    .dout(new_n223_)
  );


  anb1
  g150
  (
    .dina(new_n223__spl_00),
    .dinb(new_n204__spl_00),
    .dout(new_n224_)
  );


  anb2
  g151
  (
    .dina(G16_spl_01),
    .dinb(G12_spl_01),
    .dout(new_n225_)
  );


  anb1
  g152
  (
    .dina(G16_spl_01),
    .dinb(G12_spl_01),
    .dout(new_n226_)
  );


  anb1
  g153
  (
    .dina(new_n225_),
    .dinb(new_n226_),
    .dout(new_n227_)
  );


  nor1
  g154
  (
    .dina(G4_spl_01),
    .dinb(G8_spl_01),
    .dout(new_n228_)
  );


  nor2
  g155
  (
    .dina(G4_spl_01),
    .dinb(G8_spl_01),
    .dout(new_n229_)
  );


  anb2
  g156
  (
    .dina(new_n228_),
    .dinb(new_n229_),
    .dout(new_n230_)
  );


  anb1
  g157
  (
    .dina(new_n227__spl_),
    .dinb(new_n230__spl_),
    .dout(new_n231_)
  );


  anb2
  g158
  (
    .dina(new_n227__spl_),
    .dinb(new_n230__spl_),
    .dout(new_n232_)
  );


  anb2
  g159
  (
    .dina(new_n231_),
    .dinb(new_n232_),
    .dout(new_n233_)
  );


  nor2
  g160
  (
    .dina(G36),
    .dinb(G41_spl_10),
    .dout(new_n234_)
  );


  anb1
  g161
  (
    .dina(new_n233__spl_),
    .dinb(new_n234__spl_),
    .dout(new_n235_)
  );


  anb2
  g162
  (
    .dina(new_n233__spl_),
    .dinb(new_n234__spl_),
    .dout(new_n236_)
  );


  anb2
  g163
  (
    .dina(new_n235_),
    .dinb(new_n236_),
    .dout(new_n237_)
  );


  anb2
  g164
  (
    .dina(G32_spl_01),
    .dinb(G31_spl_01),
    .dout(new_n238_)
  );


  anb1
  g165
  (
    .dina(G32_spl_01),
    .dinb(G31_spl_01),
    .dout(new_n239_)
  );


  anb1
  g166
  (
    .dina(new_n238_),
    .dinb(new_n239_),
    .dout(new_n240_)
  );


  nor1
  g167
  (
    .dina(G29_spl_01),
    .dinb(G30_spl_01),
    .dout(new_n241_)
  );


  nor2
  g168
  (
    .dina(G29_spl_01),
    .dinb(G30_spl_01),
    .dout(new_n242_)
  );


  anb2
  g169
  (
    .dina(new_n241_),
    .dinb(new_n242_),
    .dout(new_n243_)
  );


  anb1
  g170
  (
    .dina(new_n240__spl_),
    .dinb(new_n243__spl_),
    .dout(new_n244_)
  );


  anb2
  g171
  (
    .dina(new_n240__spl_),
    .dinb(new_n243__spl_),
    .dout(new_n245_)
  );


  anb2
  g172
  (
    .dina(new_n244_),
    .dinb(new_n245_),
    .dout(new_n246_)
  );


  anb2
  g173
  (
    .dina(new_n104__spl_1),
    .dinb(new_n246__spl_0),
    .dout(new_n247_)
  );


  anb1
  g174
  (
    .dina(new_n104__spl_1),
    .dinb(new_n246__spl_0),
    .dout(new_n248_)
  );


  anb1
  g175
  (
    .dina(new_n247_),
    .dinb(new_n248_),
    .dout(new_n249_)
  );


  anb1
  g176
  (
    .dina(new_n237__spl_),
    .dinb(new_n249__spl_),
    .dout(new_n250_)
  );


  anb2
  g177
  (
    .dina(new_n237__spl_),
    .dinb(new_n249__spl_),
    .dout(new_n251_)
  );


  anb2
  g178
  (
    .dina(new_n250_),
    .dinb(new_n251_),
    .dout(new_n252_)
  );


  anb2
  g179
  (
    .dina(G15_spl_01),
    .dinb(G11_spl_01),
    .dout(new_n253_)
  );


  anb1
  g180
  (
    .dina(G15_spl_01),
    .dinb(G11_spl_01),
    .dout(new_n254_)
  );


  anb1
  g181
  (
    .dina(new_n253_),
    .dinb(new_n254_),
    .dout(new_n255_)
  );


  nor1
  g182
  (
    .dina(G3_spl_01),
    .dinb(G7_spl_01),
    .dout(new_n256_)
  );


  nor2
  g183
  (
    .dina(G3_spl_01),
    .dinb(G7_spl_01),
    .dout(new_n257_)
  );


  anb2
  g184
  (
    .dina(new_n256_),
    .dinb(new_n257_),
    .dout(new_n258_)
  );


  anb1
  g185
  (
    .dina(new_n255__spl_),
    .dinb(new_n258__spl_),
    .dout(new_n259_)
  );


  anb2
  g186
  (
    .dina(new_n255__spl_),
    .dinb(new_n258__spl_),
    .dout(new_n260_)
  );


  anb2
  g187
  (
    .dina(new_n259_),
    .dinb(new_n260_),
    .dout(new_n261_)
  );


  nor2
  g188
  (
    .dina(G35),
    .dinb(G41_spl_11),
    .dout(new_n262_)
  );


  anb1
  g189
  (
    .dina(new_n261__spl_),
    .dinb(new_n262__spl_),
    .dout(new_n263_)
  );


  anb2
  g190
  (
    .dina(new_n261__spl_),
    .dinb(new_n262__spl_),
    .dout(new_n264_)
  );


  anb2
  g191
  (
    .dina(new_n263_),
    .dinb(new_n264_),
    .dout(new_n265_)
  );


  anb2
  g192
  (
    .dina(G28_spl_01),
    .dinb(G27_spl_01),
    .dout(new_n266_)
  );


  anb1
  g193
  (
    .dina(G28_spl_01),
    .dinb(G27_spl_01),
    .dout(new_n267_)
  );


  anb1
  g194
  (
    .dina(new_n266_),
    .dinb(new_n267_),
    .dout(new_n268_)
  );


  nor1
  g195
  (
    .dina(G25_spl_01),
    .dinb(G26_spl_01),
    .dout(new_n269_)
  );


  nor2
  g196
  (
    .dina(G25_spl_01),
    .dinb(G26_spl_01),
    .dout(new_n270_)
  );


  anb2
  g197
  (
    .dina(new_n269_),
    .dinb(new_n270_),
    .dout(new_n271_)
  );


  anb1
  g198
  (
    .dina(new_n268__spl_),
    .dinb(new_n271__spl_),
    .dout(new_n272_)
  );


  anb2
  g199
  (
    .dina(new_n268__spl_),
    .dinb(new_n271__spl_),
    .dout(new_n273_)
  );


  anb2
  g200
  (
    .dina(new_n272_),
    .dinb(new_n273_),
    .dout(new_n274_)
  );


  anb2
  g201
  (
    .dina(new_n95__spl_1),
    .dinb(new_n274__spl_0),
    .dout(new_n275_)
  );


  anb1
  g202
  (
    .dina(new_n95__spl_1),
    .dinb(new_n274__spl_0),
    .dout(new_n276_)
  );


  anb1
  g203
  (
    .dina(new_n275_),
    .dinb(new_n276_),
    .dout(new_n277_)
  );


  anb1
  g204
  (
    .dina(new_n265__spl_),
    .dinb(new_n277__spl_),
    .dout(new_n278_)
  );


  anb2
  g205
  (
    .dina(new_n265__spl_),
    .dinb(new_n277__spl_),
    .dout(new_n279_)
  );


  anb2
  g206
  (
    .dina(new_n278_),
    .dinb(new_n279_),
    .dout(new_n280_)
  );


  anb2
  g207
  (
    .dina(G14_spl_01),
    .dinb(G10_spl_01),
    .dout(new_n281_)
  );


  anb1
  g208
  (
    .dina(G14_spl_01),
    .dinb(G10_spl_01),
    .dout(new_n282_)
  );


  anb1
  g209
  (
    .dina(new_n281_),
    .dinb(new_n282_),
    .dout(new_n283_)
  );


  nor1
  g210
  (
    .dina(G2_spl_01),
    .dinb(G6_spl_01),
    .dout(new_n284_)
  );


  nor2
  g211
  (
    .dina(G2_spl_01),
    .dinb(G6_spl_01),
    .dout(new_n285_)
  );


  anb2
  g212
  (
    .dina(new_n284_),
    .dinb(new_n285_),
    .dout(new_n286_)
  );


  anb1
  g213
  (
    .dina(new_n283__spl_),
    .dinb(new_n286__spl_),
    .dout(new_n287_)
  );


  anb2
  g214
  (
    .dina(new_n283__spl_),
    .dinb(new_n286__spl_),
    .dout(new_n288_)
  );


  anb2
  g215
  (
    .dina(new_n287_),
    .dinb(new_n288_),
    .dout(new_n289_)
  );


  nor2
  g216
  (
    .dina(G34),
    .dinb(G41_spl_11),
    .dout(new_n290_)
  );


  anb1
  g217
  (
    .dina(new_n289__spl_),
    .dinb(new_n290__spl_),
    .dout(new_n291_)
  );


  anb2
  g218
  (
    .dina(new_n289__spl_),
    .dinb(new_n290__spl_),
    .dout(new_n292_)
  );


  anb2
  g219
  (
    .dina(new_n291_),
    .dinb(new_n292_),
    .dout(new_n293_)
  );


  anb2
  g220
  (
    .dina(new_n246__spl_1),
    .dinb(new_n274__spl_1),
    .dout(new_n294_)
  );


  anb1
  g221
  (
    .dina(new_n246__spl_1),
    .dinb(new_n274__spl_1),
    .dout(new_n295_)
  );


  anb1
  g222
  (
    .dina(new_n294_),
    .dinb(new_n295_),
    .dout(new_n296_)
  );


  anb1
  g223
  (
    .dina(new_n293__spl_),
    .dinb(new_n296__spl_),
    .dout(new_n297_)
  );


  anb2
  g224
  (
    .dina(new_n293__spl_),
    .dinb(new_n296__spl_),
    .dout(new_n298_)
  );


  anb2
  g225
  (
    .dina(new_n297_),
    .dinb(new_n298_),
    .dout(new_n299_)
  );


  anb1
  g226
  (
    .dina(new_n110__spl_00),
    .dinb(new_n299__spl_00),
    .dout(new_n300_)
  );


  anb2
  g227
  (
    .dina(new_n280__spl_00),
    .dinb(new_n300__spl_),
    .dout(new_n301_)
  );


  anb1
  g228
  (
    .dina(new_n299__spl_00),
    .dinb(new_n110__spl_00),
    .dout(new_n302_)
  );


  anb2
  g229
  (
    .dina(new_n280__spl_00),
    .dinb(new_n302__spl_),
    .dout(new_n303_)
  );


  nor2
  g230
  (
    .dina(new_n301__spl_),
    .dinb(new_n303__spl_),
    .dout(new_n304_)
  );


  anb2
  g231
  (
    .dina(new_n252__spl_00),
    .dinb(new_n304_),
    .dout(new_n305_)
  );


  anb2
  g232
  (
    .dina(new_n252__spl_00),
    .dinb(new_n280__spl_01),
    .dout(new_n306_)
  );


  anb1
  g233
  (
    .dina(new_n252__spl_01),
    .dinb(new_n280__spl_01),
    .dout(new_n307_)
  );


  nab2
  g234
  (
    .dina(new_n306__spl_0),
    .dinb(new_n307_),
    .dout(new_n308_)
  );


  and2
  g235
  (
    .dina(new_n110__spl_01),
    .dinb(new_n299__spl_01),
    .dout(new_n309_)
  );


  anb1
  g236
  (
    .dina(new_n308_),
    .dinb(new_n309_),
    .dout(new_n310_)
  );


  anb1
  g237
  (
    .dina(new_n305_),
    .dinb(new_n310_),
    .dout(new_n311_)
  );


  anb1
  g238
  (
    .dina(new_n224__spl_),
    .dinb(new_n311__spl_),
    .dout(new_n312_)
  );


  anb2
  g239
  (
    .dina(new_n185__spl_),
    .dinb(new_n312__spl_),
    .dout(new_n313_)
  );


  anb1
  g240
  (
    .dina(new_n110__spl_01),
    .dinb(new_n313__spl_0),
    .dout(new_n314_)
  );


  anb2
  g241
  (
    .dina(new_n314__spl_),
    .dinb(G1_spl_1),
    .dout(new_n315_)
  );


  anb1
  g242
  (
    .dina(new_n314__spl_),
    .dinb(G1_spl_1),
    .dout(new_n316_)
  );


  anb1
  g243
  (
    .dina(new_n315_),
    .dinb(new_n316_),
    .dout(G1324)
  );


  anb1
  g244
  (
    .dina(new_n299__spl_01),
    .dinb(new_n313__spl_0),
    .dout(new_n318_)
  );


  anb2
  g245
  (
    .dina(new_n318__spl_),
    .dinb(G2_spl_1),
    .dout(new_n319_)
  );


  anb1
  g246
  (
    .dina(new_n318__spl_),
    .dinb(G2_spl_1),
    .dout(new_n320_)
  );


  anb1
  g247
  (
    .dina(new_n319_),
    .dinb(new_n320_),
    .dout(G1325)
  );


  anb1
  g248
  (
    .dina(new_n280__spl_10),
    .dinb(new_n313__spl_1),
    .dout(new_n322_)
  );


  anb2
  g249
  (
    .dina(new_n322__spl_),
    .dinb(G3_spl_1),
    .dout(new_n323_)
  );


  anb1
  g250
  (
    .dina(new_n322__spl_),
    .dinb(G3_spl_1),
    .dout(new_n324_)
  );


  anb1
  g251
  (
    .dina(new_n323_),
    .dinb(new_n324_),
    .dout(G1326)
  );


  anb1
  g252
  (
    .dina(new_n252__spl_01),
    .dinb(new_n313__spl_1),
    .dout(new_n326_)
  );


  anb2
  g253
  (
    .dina(new_n326__spl_),
    .dinb(G4_spl_1),
    .dout(new_n327_)
  );


  anb1
  g254
  (
    .dina(new_n326__spl_),
    .dinb(G4_spl_1),
    .dout(new_n328_)
  );


  anb1
  g255
  (
    .dina(new_n327_),
    .dinb(new_n328_),
    .dout(G1327)
  );


  and2
  g256
  (
    .dina(new_n185__spl_),
    .dinb(new_n223__spl_00),
    .dout(new_n330_)
  );


  anb1
  g257
  (
    .dina(new_n204__spl_00),
    .dinb(new_n311__spl_),
    .dout(new_n331_)
  );


  anb2
  g258
  (
    .dina(new_n330__spl_),
    .dinb(new_n331__spl_),
    .dout(new_n332_)
  );


  anb1
  g259
  (
    .dina(new_n110__spl_10),
    .dinb(new_n332__spl_0),
    .dout(new_n333_)
  );


  anb2
  g260
  (
    .dina(new_n333__spl_),
    .dinb(G5_spl_1),
    .dout(new_n334_)
  );


  anb1
  g261
  (
    .dina(new_n333__spl_),
    .dinb(G5_spl_1),
    .dout(new_n335_)
  );


  anb1
  g262
  (
    .dina(new_n334_),
    .dinb(new_n335_),
    .dout(G1328)
  );


  anb1
  g263
  (
    .dina(new_n299__spl_10),
    .dinb(new_n332__spl_0),
    .dout(new_n337_)
  );


  anb2
  g264
  (
    .dina(new_n337__spl_),
    .dinb(G6_spl_1),
    .dout(new_n338_)
  );


  anb1
  g265
  (
    .dina(new_n337__spl_),
    .dinb(G6_spl_1),
    .dout(new_n339_)
  );


  anb1
  g266
  (
    .dina(new_n338_),
    .dinb(new_n339_),
    .dout(G1329)
  );


  anb1
  g267
  (
    .dina(new_n280__spl_10),
    .dinb(new_n332__spl_1),
    .dout(new_n341_)
  );


  anb2
  g268
  (
    .dina(new_n341__spl_),
    .dinb(G7_spl_1),
    .dout(new_n342_)
  );


  anb1
  g269
  (
    .dina(new_n341__spl_),
    .dinb(G7_spl_1),
    .dout(new_n343_)
  );


  anb1
  g270
  (
    .dina(new_n342_),
    .dinb(new_n343_),
    .dout(G1330)
  );


  anb1
  g271
  (
    .dina(new_n252__spl_10),
    .dinb(new_n332__spl_1),
    .dout(new_n345_)
  );


  anb2
  g272
  (
    .dina(new_n345__spl_),
    .dinb(G8_spl_1),
    .dout(new_n346_)
  );


  anb1
  g273
  (
    .dina(new_n345__spl_),
    .dinb(G8_spl_1),
    .dout(new_n347_)
  );


  anb1
  g274
  (
    .dina(new_n346_),
    .dinb(new_n347_),
    .dout(G1331)
  );


  anb1
  g275
  (
    .dina(new_n184__spl_00),
    .dinb(new_n147__spl_00),
    .dout(new_n349_)
  );


  nor2
  g276
  (
    .dina(new_n312__spl_),
    .dinb(new_n349__spl_),
    .dout(new_n350_)
  );


  anb1
  g277
  (
    .dina(new_n110__spl_10),
    .dinb(new_n350__spl_0),
    .dout(new_n351_)
  );


  anb2
  g278
  (
    .dina(new_n351__spl_),
    .dinb(G9_spl_1),
    .dout(new_n352_)
  );


  anb1
  g279
  (
    .dina(new_n351__spl_),
    .dinb(G9_spl_1),
    .dout(new_n353_)
  );


  anb1
  g280
  (
    .dina(new_n352_),
    .dinb(new_n353_),
    .dout(G1332)
  );


  anb1
  g281
  (
    .dina(new_n299__spl_10),
    .dinb(new_n350__spl_0),
    .dout(new_n355_)
  );


  anb2
  g282
  (
    .dina(new_n355__spl_),
    .dinb(G10_spl_1),
    .dout(new_n356_)
  );


  anb1
  g283
  (
    .dina(new_n355__spl_),
    .dinb(G10_spl_1),
    .dout(new_n357_)
  );


  anb1
  g284
  (
    .dina(new_n356_),
    .dinb(new_n357_),
    .dout(G1333)
  );


  anb1
  g285
  (
    .dina(new_n280__spl_11),
    .dinb(new_n350__spl_1),
    .dout(new_n359_)
  );


  anb2
  g286
  (
    .dina(new_n359__spl_),
    .dinb(G11_spl_1),
    .dout(new_n360_)
  );


  anb1
  g287
  (
    .dina(new_n359__spl_),
    .dinb(G11_spl_1),
    .dout(new_n361_)
  );


  anb1
  g288
  (
    .dina(new_n360_),
    .dinb(new_n361_),
    .dout(G1334)
  );


  anb1
  g289
  (
    .dina(new_n252__spl_10),
    .dinb(new_n350__spl_1),
    .dout(new_n363_)
  );


  anb2
  g290
  (
    .dina(new_n363__spl_),
    .dinb(G12_spl_1),
    .dout(new_n364_)
  );


  anb1
  g291
  (
    .dina(new_n363__spl_),
    .dinb(G12_spl_1),
    .dout(new_n365_)
  );


  anb1
  g292
  (
    .dina(new_n364_),
    .dinb(new_n365_),
    .dout(G1335)
  );


  nab1
  g293
  (
    .dina(new_n223__spl_01),
    .dinb(new_n349__spl_),
    .dout(new_n367_)
  );


  nor2
  g294
  (
    .dina(new_n331__spl_),
    .dinb(new_n367__spl_),
    .dout(new_n368_)
  );


  anb1
  g295
  (
    .dina(new_n110__spl_1),
    .dinb(new_n368__spl_0),
    .dout(new_n369_)
  );


  anb2
  g296
  (
    .dina(new_n369__spl_),
    .dinb(G13_spl_1),
    .dout(new_n370_)
  );


  anb1
  g297
  (
    .dina(new_n369__spl_),
    .dinb(G13_spl_1),
    .dout(new_n371_)
  );


  anb1
  g298
  (
    .dina(new_n370_),
    .dinb(new_n371_),
    .dout(G1336)
  );


  anb1
  g299
  (
    .dina(new_n299__spl_1),
    .dinb(new_n368__spl_0),
    .dout(new_n373_)
  );


  anb2
  g300
  (
    .dina(new_n373__spl_),
    .dinb(G14_spl_1),
    .dout(new_n374_)
  );


  anb1
  g301
  (
    .dina(new_n373__spl_),
    .dinb(G14_spl_1),
    .dout(new_n375_)
  );


  anb1
  g302
  (
    .dina(new_n374_),
    .dinb(new_n375_),
    .dout(G1337)
  );


  anb1
  g303
  (
    .dina(new_n280__spl_11),
    .dinb(new_n368__spl_1),
    .dout(new_n377_)
  );


  anb2
  g304
  (
    .dina(new_n377__spl_),
    .dinb(G15_spl_1),
    .dout(new_n378_)
  );


  anb1
  g305
  (
    .dina(new_n377__spl_),
    .dinb(G15_spl_1),
    .dout(new_n379_)
  );


  anb1
  g306
  (
    .dina(new_n378_),
    .dinb(new_n379_),
    .dout(G1338)
  );


  anb1
  g307
  (
    .dina(new_n252__spl_11),
    .dinb(new_n368__spl_1),
    .dout(new_n381_)
  );


  anb2
  g308
  (
    .dina(new_n381__spl_),
    .dinb(G16_spl_1),
    .dout(new_n382_)
  );


  anb1
  g309
  (
    .dina(new_n381__spl_),
    .dinb(G16_spl_1),
    .dout(new_n383_)
  );


  anb1
  g310
  (
    .dina(new_n382_),
    .dinb(new_n383_),
    .dout(G1339)
  );


  anb1
  g311
  (
    .dina(new_n330__spl_),
    .dinb(new_n367__spl_),
    .dout(new_n385_)
  );


  and2
  g312
  (
    .dina(new_n204__spl_01),
    .dinb(new_n385_),
    .dout(new_n386_)
  );


  anb2
  g313
  (
    .dina(new_n223__spl_01),
    .dinb(new_n204__spl_01),
    .dout(new_n387_)
  );


  anb2
  g314
  (
    .dina(new_n224__spl_),
    .dinb(new_n387_),
    .dout(new_n388_)
  );


  and2
  g315
  (
    .dina(new_n147__spl_01),
    .dinb(new_n184__spl_01),
    .dout(new_n389_)
  );


  anb1
  g316
  (
    .dina(new_n388_),
    .dinb(new_n389_),
    .dout(new_n390_)
  );


  anb1
  g317
  (
    .dina(new_n386_),
    .dinb(new_n390_),
    .dout(new_n391_)
  );


  anb1
  g318
  (
    .dina(new_n300__spl_),
    .dinb(new_n306__spl_0),
    .dout(new_n392_)
  );


  anb2
  g319
  (
    .dina(new_n391__spl_0),
    .dinb(new_n392_),
    .dout(new_n393_)
  );


  anb1
  g320
  (
    .dina(new_n147__spl_01),
    .dinb(new_n393__spl_0),
    .dout(new_n394_)
  );


  anb2
  g321
  (
    .dina(new_n394__spl_),
    .dinb(G17_spl_1),
    .dout(new_n395_)
  );


  anb1
  g322
  (
    .dina(new_n394__spl_),
    .dinb(G17_spl_1),
    .dout(new_n396_)
  );


  anb1
  g323
  (
    .dina(new_n395_),
    .dinb(new_n396_),
    .dout(G1340)
  );


  anb1
  g324
  (
    .dina(new_n184__spl_01),
    .dinb(new_n393__spl_0),
    .dout(new_n398_)
  );


  anb2
  g325
  (
    .dina(new_n398__spl_),
    .dinb(G18_spl_1),
    .dout(new_n399_)
  );


  anb1
  g326
  (
    .dina(new_n398__spl_),
    .dinb(G18_spl_1),
    .dout(new_n400_)
  );


  anb1
  g327
  (
    .dina(new_n399_),
    .dinb(new_n400_),
    .dout(G1341)
  );


  anb1
  g328
  (
    .dina(new_n223__spl_10),
    .dinb(new_n393__spl_1),
    .dout(new_n402_)
  );


  anb2
  g329
  (
    .dina(new_n402__spl_),
    .dinb(G19_spl_1),
    .dout(new_n403_)
  );


  anb1
  g330
  (
    .dina(new_n402__spl_),
    .dinb(G19_spl_1),
    .dout(new_n404_)
  );


  anb1
  g331
  (
    .dina(new_n403_),
    .dinb(new_n404_),
    .dout(G1342)
  );


  anb1
  g332
  (
    .dina(new_n204__spl_10),
    .dinb(new_n393__spl_1),
    .dout(new_n406_)
  );


  anb2
  g333
  (
    .dina(new_n406__spl_),
    .dinb(G20_spl_1),
    .dout(new_n407_)
  );


  anb1
  g334
  (
    .dina(new_n406__spl_),
    .dinb(G20_spl_1),
    .dout(new_n408_)
  );


  anb1
  g335
  (
    .dina(new_n407_),
    .dinb(new_n408_),
    .dout(G1343)
  );


  anb1
  g336
  (
    .dina(new_n252__spl_11),
    .dinb(new_n391__spl_0),
    .dout(new_n410_)
  );


  anb2
  g337
  (
    .dina(new_n301__spl_),
    .dinb(new_n410__spl_),
    .dout(new_n411_)
  );


  anb1
  g338
  (
    .dina(new_n147__spl_10),
    .dinb(new_n411__spl_0),
    .dout(new_n412_)
  );


  anb2
  g339
  (
    .dina(new_n412__spl_),
    .dinb(G21_spl_1),
    .dout(new_n413_)
  );


  anb1
  g340
  (
    .dina(new_n412__spl_),
    .dinb(G21_spl_1),
    .dout(new_n414_)
  );


  anb1
  g341
  (
    .dina(new_n413_),
    .dinb(new_n414_),
    .dout(G1344)
  );


  anb1
  g342
  (
    .dina(new_n184__spl_10),
    .dinb(new_n411__spl_0),
    .dout(new_n416_)
  );


  anb2
  g343
  (
    .dina(new_n416__spl_),
    .dinb(G22_spl_1),
    .dout(new_n417_)
  );


  anb1
  g344
  (
    .dina(new_n416__spl_),
    .dinb(G22_spl_1),
    .dout(new_n418_)
  );


  anb1
  g345
  (
    .dina(new_n417_),
    .dinb(new_n418_),
    .dout(G1345)
  );


  anb1
  g346
  (
    .dina(new_n223__spl_10),
    .dinb(new_n411__spl_1),
    .dout(new_n420_)
  );


  anb2
  g347
  (
    .dina(new_n420__spl_),
    .dinb(G23_spl_1),
    .dout(new_n421_)
  );


  anb1
  g348
  (
    .dina(new_n420__spl_),
    .dinb(G23_spl_1),
    .dout(new_n422_)
  );


  anb1
  g349
  (
    .dina(new_n421_),
    .dinb(new_n422_),
    .dout(G1346)
  );


  anb1
  g350
  (
    .dina(new_n204__spl_10),
    .dinb(new_n411__spl_1),
    .dout(new_n424_)
  );


  anb2
  g351
  (
    .dina(new_n424__spl_),
    .dinb(G24_spl_1),
    .dout(new_n425_)
  );


  anb1
  g352
  (
    .dina(new_n424__spl_),
    .dinb(G24_spl_1),
    .dout(new_n426_)
  );


  anb1
  g353
  (
    .dina(new_n425_),
    .dinb(new_n426_),
    .dout(G1347)
  );


  anb1
  g354
  (
    .dina(new_n302__spl_),
    .dinb(new_n306__spl_),
    .dout(new_n428_)
  );


  anb2
  g355
  (
    .dina(new_n391__spl_),
    .dinb(new_n428_),
    .dout(new_n429_)
  );


  anb1
  g356
  (
    .dina(new_n147__spl_10),
    .dinb(new_n429__spl_0),
    .dout(new_n430_)
  );


  anb2
  g357
  (
    .dina(new_n430__spl_),
    .dinb(G25_spl_1),
    .dout(new_n431_)
  );


  anb1
  g358
  (
    .dina(new_n430__spl_),
    .dinb(G25_spl_1),
    .dout(new_n432_)
  );


  anb1
  g359
  (
    .dina(new_n431_),
    .dinb(new_n432_),
    .dout(G1348)
  );


  anb1
  g360
  (
    .dina(new_n184__spl_10),
    .dinb(new_n429__spl_0),
    .dout(new_n434_)
  );


  anb2
  g361
  (
    .dina(new_n434__spl_),
    .dinb(G26_spl_1),
    .dout(new_n435_)
  );


  anb1
  g362
  (
    .dina(new_n434__spl_),
    .dinb(G26_spl_1),
    .dout(new_n436_)
  );


  anb1
  g363
  (
    .dina(new_n435_),
    .dinb(new_n436_),
    .dout(G1349)
  );


  anb1
  g364
  (
    .dina(new_n223__spl_11),
    .dinb(new_n429__spl_1),
    .dout(new_n438_)
  );


  anb2
  g365
  (
    .dina(new_n438__spl_),
    .dinb(G27_spl_1),
    .dout(new_n439_)
  );


  anb1
  g366
  (
    .dina(new_n438__spl_),
    .dinb(G27_spl_1),
    .dout(new_n440_)
  );


  anb1
  g367
  (
    .dina(new_n439_),
    .dinb(new_n440_),
    .dout(G1350)
  );


  anb1
  g368
  (
    .dina(new_n204__spl_11),
    .dinb(new_n429__spl_1),
    .dout(new_n442_)
  );


  anb2
  g369
  (
    .dina(new_n442__spl_),
    .dinb(G28_spl_1),
    .dout(new_n443_)
  );


  anb1
  g370
  (
    .dina(new_n442__spl_),
    .dinb(G28_spl_1),
    .dout(new_n444_)
  );


  anb1
  g371
  (
    .dina(new_n443_),
    .dinb(new_n444_),
    .dout(G1351)
  );


  anb2
  g372
  (
    .dina(new_n303__spl_),
    .dinb(new_n410__spl_),
    .dout(new_n446_)
  );


  anb1
  g373
  (
    .dina(new_n147__spl_1),
    .dinb(new_n446__spl_0),
    .dout(new_n447_)
  );


  anb2
  g374
  (
    .dina(new_n447__spl_),
    .dinb(G29_spl_1),
    .dout(new_n448_)
  );


  anb1
  g375
  (
    .dina(new_n447__spl_),
    .dinb(G29_spl_1),
    .dout(new_n449_)
  );


  anb1
  g376
  (
    .dina(new_n448_),
    .dinb(new_n449_),
    .dout(G1352)
  );


  anb1
  g377
  (
    .dina(new_n184__spl_1),
    .dinb(new_n446__spl_0),
    .dout(new_n451_)
  );


  anb2
  g378
  (
    .dina(new_n451__spl_),
    .dinb(G30_spl_1),
    .dout(new_n452_)
  );


  anb1
  g379
  (
    .dina(new_n451__spl_),
    .dinb(G30_spl_1),
    .dout(new_n453_)
  );


  anb1
  g380
  (
    .dina(new_n452_),
    .dinb(new_n453_),
    .dout(G1353)
  );


  anb1
  g381
  (
    .dina(new_n223__spl_11),
    .dinb(new_n446__spl_1),
    .dout(new_n455_)
  );


  anb2
  g382
  (
    .dina(new_n455__spl_),
    .dinb(G31_spl_1),
    .dout(new_n456_)
  );


  anb1
  g383
  (
    .dina(new_n455__spl_),
    .dinb(G31_spl_1),
    .dout(new_n457_)
  );


  anb1
  g384
  (
    .dina(new_n456_),
    .dinb(new_n457_),
    .dout(G1354)
  );


  anb1
  g385
  (
    .dina(new_n204__spl_11),
    .dinb(new_n446__spl_1),
    .dout(new_n459_)
  );


  anb2
  g386
  (
    .dina(new_n459__spl_),
    .dinb(G32_spl_1),
    .dout(new_n460_)
  );


  anb1
  g387
  (
    .dina(new_n459__spl_),
    .dinb(G32_spl_1),
    .dout(new_n461_)
  );


  anb1
  g388
  (
    .dina(new_n460_),
    .dinb(new_n461_),
    .dout(G1355)
  );


  splt
  gG13
  (
    .dout(G13_spl_),
    .din(G13)
  );


  splt
  gG13_spl_
  (
    .dout(G13_spl_0),
    .din(G13_spl_)
  );


  splt
  gG13_spl_0
  (
    .dout(G13_spl_00),
    .din(G13_spl_0)
  );


  splt
  gG13_spl_0
  (
    .dout(G13_spl_01),
    .din(G13_spl_0)
  );


  splt
  gG13_spl_
  (
    .dout(G13_spl_1),
    .din(G13_spl_)
  );


  splt
  gG9
  (
    .dout(G9_spl_),
    .din(G9)
  );


  splt
  gG9_spl_
  (
    .dout(G9_spl_0),
    .din(G9_spl_)
  );


  splt
  gG9_spl_0
  (
    .dout(G9_spl_00),
    .din(G9_spl_0)
  );


  splt
  gG9_spl_0
  (
    .dout(G9_spl_01),
    .din(G9_spl_0)
  );


  splt
  gG9_spl_
  (
    .dout(G9_spl_1),
    .din(G9_spl_)
  );


  splt
  gG1
  (
    .dout(G1_spl_),
    .din(G1)
  );


  splt
  gG1_spl_
  (
    .dout(G1_spl_0),
    .din(G1_spl_)
  );


  splt
  gG1_spl_0
  (
    .dout(G1_spl_00),
    .din(G1_spl_0)
  );


  splt
  gG1_spl_0
  (
    .dout(G1_spl_01),
    .din(G1_spl_0)
  );


  splt
  gG1_spl_
  (
    .dout(G1_spl_1),
    .din(G1_spl_)
  );


  splt
  gG5
  (
    .dout(G5_spl_),
    .din(G5)
  );


  splt
  gG5_spl_
  (
    .dout(G5_spl_0),
    .din(G5_spl_)
  );


  splt
  gG5_spl_0
  (
    .dout(G5_spl_00),
    .din(G5_spl_0)
  );


  splt
  gG5_spl_0
  (
    .dout(G5_spl_01),
    .din(G5_spl_0)
  );


  splt
  gG5_spl_
  (
    .dout(G5_spl_1),
    .din(G5_spl_)
  );


  splt
  gnew_n76_
  (
    .dout(new_n76__spl_),
    .din(new_n76_)
  );


  splt
  gnew_n79_
  (
    .dout(new_n79__spl_),
    .din(new_n79_)
  );


  splt
  gG41
  (
    .dout(G41_spl_),
    .din(G41)
  );


  splt
  gG41_spl_
  (
    .dout(G41_spl_0),
    .din(G41_spl_)
  );


  splt
  gG41_spl_0
  (
    .dout(G41_spl_00),
    .din(G41_spl_0)
  );


  splt
  gG41_spl_0
  (
    .dout(G41_spl_01),
    .din(G41_spl_0)
  );


  splt
  gG41_spl_
  (
    .dout(G41_spl_1),
    .din(G41_spl_)
  );


  splt
  gG41_spl_1
  (
    .dout(G41_spl_10),
    .din(G41_spl_1)
  );


  splt
  gG41_spl_1
  (
    .dout(G41_spl_11),
    .din(G41_spl_1)
  );


  splt
  gnew_n82_
  (
    .dout(new_n82__spl_),
    .din(new_n82_)
  );


  splt
  gnew_n83_
  (
    .dout(new_n83__spl_),
    .din(new_n83_)
  );


  splt
  gG20
  (
    .dout(G20_spl_),
    .din(G20)
  );


  splt
  gG20_spl_
  (
    .dout(G20_spl_0),
    .din(G20_spl_)
  );


  splt
  gG20_spl_0
  (
    .dout(G20_spl_00),
    .din(G20_spl_0)
  );


  splt
  gG20_spl_0
  (
    .dout(G20_spl_01),
    .din(G20_spl_0)
  );


  splt
  gG20_spl_
  (
    .dout(G20_spl_1),
    .din(G20_spl_)
  );


  splt
  gG19
  (
    .dout(G19_spl_),
    .din(G19)
  );


  splt
  gG19_spl_
  (
    .dout(G19_spl_0),
    .din(G19_spl_)
  );


  splt
  gG19_spl_0
  (
    .dout(G19_spl_00),
    .din(G19_spl_0)
  );


  splt
  gG19_spl_0
  (
    .dout(G19_spl_01),
    .din(G19_spl_0)
  );


  splt
  gG19_spl_
  (
    .dout(G19_spl_1),
    .din(G19_spl_)
  );


  splt
  gG17
  (
    .dout(G17_spl_),
    .din(G17)
  );


  splt
  gG17_spl_
  (
    .dout(G17_spl_0),
    .din(G17_spl_)
  );


  splt
  gG17_spl_0
  (
    .dout(G17_spl_00),
    .din(G17_spl_0)
  );


  splt
  gG17_spl_0
  (
    .dout(G17_spl_01),
    .din(G17_spl_0)
  );


  splt
  gG17_spl_
  (
    .dout(G17_spl_1),
    .din(G17_spl_)
  );


  splt
  gG18
  (
    .dout(G18_spl_),
    .din(G18)
  );


  splt
  gG18_spl_
  (
    .dout(G18_spl_0),
    .din(G18_spl_)
  );


  splt
  gG18_spl_0
  (
    .dout(G18_spl_00),
    .din(G18_spl_0)
  );


  splt
  gG18_spl_0
  (
    .dout(G18_spl_01),
    .din(G18_spl_0)
  );


  splt
  gG18_spl_
  (
    .dout(G18_spl_1),
    .din(G18_spl_)
  );


  splt
  gnew_n89_
  (
    .dout(new_n89__spl_),
    .din(new_n89_)
  );


  splt
  gnew_n92_
  (
    .dout(new_n92__spl_),
    .din(new_n92_)
  );


  splt
  gG24
  (
    .dout(G24_spl_),
    .din(G24)
  );


  splt
  gG24_spl_
  (
    .dout(G24_spl_0),
    .din(G24_spl_)
  );


  splt
  gG24_spl_0
  (
    .dout(G24_spl_00),
    .din(G24_spl_0)
  );


  splt
  gG24_spl_0
  (
    .dout(G24_spl_01),
    .din(G24_spl_0)
  );


  splt
  gG24_spl_
  (
    .dout(G24_spl_1),
    .din(G24_spl_)
  );


  splt
  gG23
  (
    .dout(G23_spl_),
    .din(G23)
  );


  splt
  gG23_spl_
  (
    .dout(G23_spl_0),
    .din(G23_spl_)
  );


  splt
  gG23_spl_0
  (
    .dout(G23_spl_00),
    .din(G23_spl_0)
  );


  splt
  gG23_spl_0
  (
    .dout(G23_spl_01),
    .din(G23_spl_0)
  );


  splt
  gG23_spl_
  (
    .dout(G23_spl_1),
    .din(G23_spl_)
  );


  splt
  gG21
  (
    .dout(G21_spl_),
    .din(G21)
  );


  splt
  gG21_spl_
  (
    .dout(G21_spl_0),
    .din(G21_spl_)
  );


  splt
  gG21_spl_0
  (
    .dout(G21_spl_00),
    .din(G21_spl_0)
  );


  splt
  gG21_spl_0
  (
    .dout(G21_spl_01),
    .din(G21_spl_0)
  );


  splt
  gG21_spl_
  (
    .dout(G21_spl_1),
    .din(G21_spl_)
  );


  splt
  gG22
  (
    .dout(G22_spl_),
    .din(G22)
  );


  splt
  gG22_spl_
  (
    .dout(G22_spl_0),
    .din(G22_spl_)
  );


  splt
  gG22_spl_0
  (
    .dout(G22_spl_00),
    .din(G22_spl_0)
  );


  splt
  gG22_spl_0
  (
    .dout(G22_spl_01),
    .din(G22_spl_0)
  );


  splt
  gG22_spl_
  (
    .dout(G22_spl_1),
    .din(G22_spl_)
  );


  splt
  gnew_n98_
  (
    .dout(new_n98__spl_),
    .din(new_n98_)
  );


  splt
  gnew_n101_
  (
    .dout(new_n101__spl_),
    .din(new_n101_)
  );


  splt
  gnew_n95_
  (
    .dout(new_n95__spl_),
    .din(new_n95_)
  );


  splt
  gnew_n95__spl_
  (
    .dout(new_n95__spl_0),
    .din(new_n95__spl_)
  );


  splt
  gnew_n95__spl_
  (
    .dout(new_n95__spl_1),
    .din(new_n95__spl_)
  );


  splt
  gnew_n104_
  (
    .dout(new_n104__spl_),
    .din(new_n104_)
  );


  splt
  gnew_n104__spl_
  (
    .dout(new_n104__spl_0),
    .din(new_n104__spl_)
  );


  splt
  gnew_n104__spl_
  (
    .dout(new_n104__spl_1),
    .din(new_n104__spl_)
  );


  splt
  gnew_n86_
  (
    .dout(new_n86__spl_),
    .din(new_n86_)
  );


  splt
  gnew_n107_
  (
    .dout(new_n107__spl_),
    .din(new_n107_)
  );


  splt
  gG29
  (
    .dout(G29_spl_),
    .din(G29)
  );


  splt
  gG29_spl_
  (
    .dout(G29_spl_0),
    .din(G29_spl_)
  );


  splt
  gG29_spl_0
  (
    .dout(G29_spl_00),
    .din(G29_spl_0)
  );


  splt
  gG29_spl_0
  (
    .dout(G29_spl_01),
    .din(G29_spl_0)
  );


  splt
  gG29_spl_
  (
    .dout(G29_spl_1),
    .din(G29_spl_)
  );


  splt
  gG25
  (
    .dout(G25_spl_),
    .din(G25)
  );


  splt
  gG25_spl_
  (
    .dout(G25_spl_0),
    .din(G25_spl_)
  );


  splt
  gG25_spl_0
  (
    .dout(G25_spl_00),
    .din(G25_spl_0)
  );


  splt
  gG25_spl_0
  (
    .dout(G25_spl_01),
    .din(G25_spl_0)
  );


  splt
  gG25_spl_
  (
    .dout(G25_spl_1),
    .din(G25_spl_)
  );


  splt
  gnew_n113_
  (
    .dout(new_n113__spl_),
    .din(new_n113_)
  );


  splt
  gnew_n116_
  (
    .dout(new_n116__spl_),
    .din(new_n116_)
  );


  splt
  gnew_n119_
  (
    .dout(new_n119__spl_),
    .din(new_n119_)
  );


  splt
  gnew_n120_
  (
    .dout(new_n120__spl_),
    .din(new_n120_)
  );


  splt
  gG8
  (
    .dout(G8_spl_),
    .din(G8)
  );


  splt
  gG8_spl_
  (
    .dout(G8_spl_0),
    .din(G8_spl_)
  );


  splt
  gG8_spl_0
  (
    .dout(G8_spl_00),
    .din(G8_spl_0)
  );


  splt
  gG8_spl_0
  (
    .dout(G8_spl_01),
    .din(G8_spl_0)
  );


  splt
  gG8_spl_
  (
    .dout(G8_spl_1),
    .din(G8_spl_)
  );


  splt
  gG7
  (
    .dout(G7_spl_),
    .din(G7)
  );


  splt
  gG7_spl_
  (
    .dout(G7_spl_0),
    .din(G7_spl_)
  );


  splt
  gG7_spl_0
  (
    .dout(G7_spl_00),
    .din(G7_spl_0)
  );


  splt
  gG7_spl_0
  (
    .dout(G7_spl_01),
    .din(G7_spl_0)
  );


  splt
  gG7_spl_
  (
    .dout(G7_spl_1),
    .din(G7_spl_)
  );


  splt
  gG6
  (
    .dout(G6_spl_),
    .din(G6)
  );


  splt
  gG6_spl_
  (
    .dout(G6_spl_0),
    .din(G6_spl_)
  );


  splt
  gG6_spl_0
  (
    .dout(G6_spl_00),
    .din(G6_spl_0)
  );


  splt
  gG6_spl_0
  (
    .dout(G6_spl_01),
    .din(G6_spl_0)
  );


  splt
  gG6_spl_
  (
    .dout(G6_spl_1),
    .din(G6_spl_)
  );


  splt
  gnew_n126_
  (
    .dout(new_n126__spl_),
    .din(new_n126_)
  );


  splt
  gnew_n129_
  (
    .dout(new_n129__spl_),
    .din(new_n129_)
  );


  splt
  gG4
  (
    .dout(G4_spl_),
    .din(G4)
  );


  splt
  gG4_spl_
  (
    .dout(G4_spl_0),
    .din(G4_spl_)
  );


  splt
  gG4_spl_0
  (
    .dout(G4_spl_00),
    .din(G4_spl_0)
  );


  splt
  gG4_spl_0
  (
    .dout(G4_spl_01),
    .din(G4_spl_0)
  );


  splt
  gG4_spl_
  (
    .dout(G4_spl_1),
    .din(G4_spl_)
  );


  splt
  gG3
  (
    .dout(G3_spl_),
    .din(G3)
  );


  splt
  gG3_spl_
  (
    .dout(G3_spl_0),
    .din(G3_spl_)
  );


  splt
  gG3_spl_0
  (
    .dout(G3_spl_00),
    .din(G3_spl_0)
  );


  splt
  gG3_spl_0
  (
    .dout(G3_spl_01),
    .din(G3_spl_0)
  );


  splt
  gG3_spl_
  (
    .dout(G3_spl_1),
    .din(G3_spl_)
  );


  splt
  gG2
  (
    .dout(G2_spl_),
    .din(G2)
  );


  splt
  gG2_spl_
  (
    .dout(G2_spl_0),
    .din(G2_spl_)
  );


  splt
  gG2_spl_0
  (
    .dout(G2_spl_00),
    .din(G2_spl_0)
  );


  splt
  gG2_spl_0
  (
    .dout(G2_spl_01),
    .din(G2_spl_0)
  );


  splt
  gG2_spl_
  (
    .dout(G2_spl_1),
    .din(G2_spl_)
  );


  splt
  gnew_n135_
  (
    .dout(new_n135__spl_),
    .din(new_n135_)
  );


  splt
  gnew_n138_
  (
    .dout(new_n138__spl_),
    .din(new_n138_)
  );


  splt
  gnew_n132_
  (
    .dout(new_n132__spl_),
    .din(new_n132_)
  );


  splt
  gnew_n132__spl_
  (
    .dout(new_n132__spl_0),
    .din(new_n132__spl_)
  );


  splt
  gnew_n132__spl_
  (
    .dout(new_n132__spl_1),
    .din(new_n132__spl_)
  );


  splt
  gnew_n141_
  (
    .dout(new_n141__spl_),
    .din(new_n141_)
  );


  splt
  gnew_n141__spl_
  (
    .dout(new_n141__spl_0),
    .din(new_n141__spl_)
  );


  splt
  gnew_n141__spl_
  (
    .dout(new_n141__spl_1),
    .din(new_n141__spl_)
  );


  splt
  gnew_n123_
  (
    .dout(new_n123__spl_),
    .din(new_n123_)
  );


  splt
  gnew_n144_
  (
    .dout(new_n144__spl_),
    .din(new_n144_)
  );


  splt
  gG30
  (
    .dout(G30_spl_),
    .din(G30)
  );


  splt
  gG30_spl_
  (
    .dout(G30_spl_0),
    .din(G30_spl_)
  );


  splt
  gG30_spl_0
  (
    .dout(G30_spl_00),
    .din(G30_spl_0)
  );


  splt
  gG30_spl_0
  (
    .dout(G30_spl_01),
    .din(G30_spl_0)
  );


  splt
  gG30_spl_
  (
    .dout(G30_spl_1),
    .din(G30_spl_)
  );


  splt
  gG26
  (
    .dout(G26_spl_),
    .din(G26)
  );


  splt
  gG26_spl_
  (
    .dout(G26_spl_0),
    .din(G26_spl_)
  );


  splt
  gG26_spl_0
  (
    .dout(G26_spl_00),
    .din(G26_spl_0)
  );


  splt
  gG26_spl_0
  (
    .dout(G26_spl_01),
    .din(G26_spl_0)
  );


  splt
  gG26_spl_
  (
    .dout(G26_spl_1),
    .din(G26_spl_)
  );


  splt
  gnew_n150_
  (
    .dout(new_n150__spl_),
    .din(new_n150_)
  );


  splt
  gnew_n153_
  (
    .dout(new_n153__spl_),
    .din(new_n153_)
  );


  splt
  gnew_n156_
  (
    .dout(new_n156__spl_),
    .din(new_n156_)
  );


  splt
  gnew_n157_
  (
    .dout(new_n157__spl_),
    .din(new_n157_)
  );


  splt
  gG16
  (
    .dout(G16_spl_),
    .din(G16)
  );


  splt
  gG16_spl_
  (
    .dout(G16_spl_0),
    .din(G16_spl_)
  );


  splt
  gG16_spl_0
  (
    .dout(G16_spl_00),
    .din(G16_spl_0)
  );


  splt
  gG16_spl_0
  (
    .dout(G16_spl_01),
    .din(G16_spl_0)
  );


  splt
  gG16_spl_
  (
    .dout(G16_spl_1),
    .din(G16_spl_)
  );


  splt
  gG15
  (
    .dout(G15_spl_),
    .din(G15)
  );


  splt
  gG15_spl_
  (
    .dout(G15_spl_0),
    .din(G15_spl_)
  );


  splt
  gG15_spl_0
  (
    .dout(G15_spl_00),
    .din(G15_spl_0)
  );


  splt
  gG15_spl_0
  (
    .dout(G15_spl_01),
    .din(G15_spl_0)
  );


  splt
  gG15_spl_
  (
    .dout(G15_spl_1),
    .din(G15_spl_)
  );


  splt
  gG14
  (
    .dout(G14_spl_),
    .din(G14)
  );


  splt
  gG14_spl_
  (
    .dout(G14_spl_0),
    .din(G14_spl_)
  );


  splt
  gG14_spl_0
  (
    .dout(G14_spl_00),
    .din(G14_spl_0)
  );


  splt
  gG14_spl_0
  (
    .dout(G14_spl_01),
    .din(G14_spl_0)
  );


  splt
  gG14_spl_
  (
    .dout(G14_spl_1),
    .din(G14_spl_)
  );


  splt
  gnew_n163_
  (
    .dout(new_n163__spl_),
    .din(new_n163_)
  );


  splt
  gnew_n166_
  (
    .dout(new_n166__spl_),
    .din(new_n166_)
  );


  splt
  gG12
  (
    .dout(G12_spl_),
    .din(G12)
  );


  splt
  gG12_spl_
  (
    .dout(G12_spl_0),
    .din(G12_spl_)
  );


  splt
  gG12_spl_0
  (
    .dout(G12_spl_00),
    .din(G12_spl_0)
  );


  splt
  gG12_spl_0
  (
    .dout(G12_spl_01),
    .din(G12_spl_0)
  );


  splt
  gG12_spl_
  (
    .dout(G12_spl_1),
    .din(G12_spl_)
  );


  splt
  gG11
  (
    .dout(G11_spl_),
    .din(G11)
  );


  splt
  gG11_spl_
  (
    .dout(G11_spl_0),
    .din(G11_spl_)
  );


  splt
  gG11_spl_0
  (
    .dout(G11_spl_00),
    .din(G11_spl_0)
  );


  splt
  gG11_spl_0
  (
    .dout(G11_spl_01),
    .din(G11_spl_0)
  );


  splt
  gG11_spl_
  (
    .dout(G11_spl_1),
    .din(G11_spl_)
  );


  splt
  gG10
  (
    .dout(G10_spl_),
    .din(G10)
  );


  splt
  gG10_spl_
  (
    .dout(G10_spl_0),
    .din(G10_spl_)
  );


  splt
  gG10_spl_0
  (
    .dout(G10_spl_00),
    .din(G10_spl_0)
  );


  splt
  gG10_spl_0
  (
    .dout(G10_spl_01),
    .din(G10_spl_0)
  );


  splt
  gG10_spl_
  (
    .dout(G10_spl_1),
    .din(G10_spl_)
  );


  splt
  gnew_n172_
  (
    .dout(new_n172__spl_),
    .din(new_n172_)
  );


  splt
  gnew_n175_
  (
    .dout(new_n175__spl_),
    .din(new_n175_)
  );


  splt
  gnew_n169_
  (
    .dout(new_n169__spl_),
    .din(new_n169_)
  );


  splt
  gnew_n169__spl_
  (
    .dout(new_n169__spl_0),
    .din(new_n169__spl_)
  );


  splt
  gnew_n169__spl_
  (
    .dout(new_n169__spl_1),
    .din(new_n169__spl_)
  );


  splt
  gnew_n178_
  (
    .dout(new_n178__spl_),
    .din(new_n178_)
  );


  splt
  gnew_n178__spl_
  (
    .dout(new_n178__spl_0),
    .din(new_n178__spl_)
  );


  splt
  gnew_n178__spl_
  (
    .dout(new_n178__spl_1),
    .din(new_n178__spl_)
  );


  splt
  gnew_n160_
  (
    .dout(new_n160__spl_),
    .din(new_n160_)
  );


  splt
  gnew_n181_
  (
    .dout(new_n181__spl_),
    .din(new_n181_)
  );


  splt
  gnew_n184_
  (
    .dout(new_n184__spl_),
    .din(new_n184_)
  );


  splt
  gnew_n184__spl_
  (
    .dout(new_n184__spl_0),
    .din(new_n184__spl_)
  );


  splt
  gnew_n184__spl_0
  (
    .dout(new_n184__spl_00),
    .din(new_n184__spl_0)
  );


  splt
  gnew_n184__spl_0
  (
    .dout(new_n184__spl_01),
    .din(new_n184__spl_0)
  );


  splt
  gnew_n184__spl_
  (
    .dout(new_n184__spl_1),
    .din(new_n184__spl_)
  );


  splt
  gnew_n184__spl_1
  (
    .dout(new_n184__spl_10),
    .din(new_n184__spl_1)
  );


  splt
  gnew_n147_
  (
    .dout(new_n147__spl_),
    .din(new_n147_)
  );


  splt
  gnew_n147__spl_
  (
    .dout(new_n147__spl_0),
    .din(new_n147__spl_)
  );


  splt
  gnew_n147__spl_0
  (
    .dout(new_n147__spl_00),
    .din(new_n147__spl_0)
  );


  splt
  gnew_n147__spl_0
  (
    .dout(new_n147__spl_01),
    .din(new_n147__spl_0)
  );


  splt
  gnew_n147__spl_
  (
    .dout(new_n147__spl_1),
    .din(new_n147__spl_)
  );


  splt
  gnew_n147__spl_1
  (
    .dout(new_n147__spl_10),
    .din(new_n147__spl_1)
  );


  splt
  gG32
  (
    .dout(G32_spl_),
    .din(G32)
  );


  splt
  gG32_spl_
  (
    .dout(G32_spl_0),
    .din(G32_spl_)
  );


  splt
  gG32_spl_0
  (
    .dout(G32_spl_00),
    .din(G32_spl_0)
  );


  splt
  gG32_spl_0
  (
    .dout(G32_spl_01),
    .din(G32_spl_0)
  );


  splt
  gG32_spl_
  (
    .dout(G32_spl_1),
    .din(G32_spl_)
  );


  splt
  gG28
  (
    .dout(G28_spl_),
    .din(G28)
  );


  splt
  gG28_spl_
  (
    .dout(G28_spl_0),
    .din(G28_spl_)
  );


  splt
  gG28_spl_0
  (
    .dout(G28_spl_00),
    .din(G28_spl_0)
  );


  splt
  gG28_spl_0
  (
    .dout(G28_spl_01),
    .din(G28_spl_0)
  );


  splt
  gG28_spl_
  (
    .dout(G28_spl_1),
    .din(G28_spl_)
  );


  splt
  gnew_n188_
  (
    .dout(new_n188__spl_),
    .din(new_n188_)
  );


  splt
  gnew_n191_
  (
    .dout(new_n191__spl_),
    .din(new_n191_)
  );


  splt
  gnew_n194_
  (
    .dout(new_n194__spl_),
    .din(new_n194_)
  );


  splt
  gnew_n195_
  (
    .dout(new_n195__spl_),
    .din(new_n195_)
  );


  splt
  gnew_n198_
  (
    .dout(new_n198__spl_),
    .din(new_n198_)
  );


  splt
  gnew_n201_
  (
    .dout(new_n201__spl_),
    .din(new_n201_)
  );


  splt
  gG31
  (
    .dout(G31_spl_),
    .din(G31)
  );


  splt
  gG31_spl_
  (
    .dout(G31_spl_0),
    .din(G31_spl_)
  );


  splt
  gG31_spl_0
  (
    .dout(G31_spl_00),
    .din(G31_spl_0)
  );


  splt
  gG31_spl_0
  (
    .dout(G31_spl_01),
    .din(G31_spl_0)
  );


  splt
  gG31_spl_
  (
    .dout(G31_spl_1),
    .din(G31_spl_)
  );


  splt
  gG27
  (
    .dout(G27_spl_),
    .din(G27)
  );


  splt
  gG27_spl_
  (
    .dout(G27_spl_0),
    .din(G27_spl_)
  );


  splt
  gG27_spl_0
  (
    .dout(G27_spl_00),
    .din(G27_spl_0)
  );


  splt
  gG27_spl_0
  (
    .dout(G27_spl_01),
    .din(G27_spl_0)
  );


  splt
  gG27_spl_
  (
    .dout(G27_spl_1),
    .din(G27_spl_)
  );


  splt
  gnew_n207_
  (
    .dout(new_n207__spl_),
    .din(new_n207_)
  );


  splt
  gnew_n210_
  (
    .dout(new_n210__spl_),
    .din(new_n210_)
  );


  splt
  gnew_n213_
  (
    .dout(new_n213__spl_),
    .din(new_n213_)
  );


  splt
  gnew_n214_
  (
    .dout(new_n214__spl_),
    .din(new_n214_)
  );


  splt
  gnew_n217_
  (
    .dout(new_n217__spl_),
    .din(new_n217_)
  );


  splt
  gnew_n220_
  (
    .dout(new_n220__spl_),
    .din(new_n220_)
  );


  splt
  gnew_n223_
  (
    .dout(new_n223__spl_),
    .din(new_n223_)
  );


  splt
  gnew_n223__spl_
  (
    .dout(new_n223__spl_0),
    .din(new_n223__spl_)
  );


  splt
  gnew_n223__spl_0
  (
    .dout(new_n223__spl_00),
    .din(new_n223__spl_0)
  );


  splt
  gnew_n223__spl_0
  (
    .dout(new_n223__spl_01),
    .din(new_n223__spl_0)
  );


  splt
  gnew_n223__spl_
  (
    .dout(new_n223__spl_1),
    .din(new_n223__spl_)
  );


  splt
  gnew_n223__spl_1
  (
    .dout(new_n223__spl_10),
    .din(new_n223__spl_1)
  );


  splt
  gnew_n223__spl_1
  (
    .dout(new_n223__spl_11),
    .din(new_n223__spl_1)
  );


  splt
  gnew_n204_
  (
    .dout(new_n204__spl_),
    .din(new_n204_)
  );


  splt
  gnew_n204__spl_
  (
    .dout(new_n204__spl_0),
    .din(new_n204__spl_)
  );


  splt
  gnew_n204__spl_0
  (
    .dout(new_n204__spl_00),
    .din(new_n204__spl_0)
  );


  splt
  gnew_n204__spl_0
  (
    .dout(new_n204__spl_01),
    .din(new_n204__spl_0)
  );


  splt
  gnew_n204__spl_
  (
    .dout(new_n204__spl_1),
    .din(new_n204__spl_)
  );


  splt
  gnew_n204__spl_1
  (
    .dout(new_n204__spl_10),
    .din(new_n204__spl_1)
  );


  splt
  gnew_n204__spl_1
  (
    .dout(new_n204__spl_11),
    .din(new_n204__spl_1)
  );


  splt
  gnew_n227_
  (
    .dout(new_n227__spl_),
    .din(new_n227_)
  );


  splt
  gnew_n230_
  (
    .dout(new_n230__spl_),
    .din(new_n230_)
  );


  splt
  gnew_n233_
  (
    .dout(new_n233__spl_),
    .din(new_n233_)
  );


  splt
  gnew_n234_
  (
    .dout(new_n234__spl_),
    .din(new_n234_)
  );


  splt
  gnew_n240_
  (
    .dout(new_n240__spl_),
    .din(new_n240_)
  );


  splt
  gnew_n243_
  (
    .dout(new_n243__spl_),
    .din(new_n243_)
  );


  splt
  gnew_n246_
  (
    .dout(new_n246__spl_),
    .din(new_n246_)
  );


  splt
  gnew_n246__spl_
  (
    .dout(new_n246__spl_0),
    .din(new_n246__spl_)
  );


  splt
  gnew_n246__spl_
  (
    .dout(new_n246__spl_1),
    .din(new_n246__spl_)
  );


  splt
  gnew_n237_
  (
    .dout(new_n237__spl_),
    .din(new_n237_)
  );


  splt
  gnew_n249_
  (
    .dout(new_n249__spl_),
    .din(new_n249_)
  );


  splt
  gnew_n255_
  (
    .dout(new_n255__spl_),
    .din(new_n255_)
  );


  splt
  gnew_n258_
  (
    .dout(new_n258__spl_),
    .din(new_n258_)
  );


  splt
  gnew_n261_
  (
    .dout(new_n261__spl_),
    .din(new_n261_)
  );


  splt
  gnew_n262_
  (
    .dout(new_n262__spl_),
    .din(new_n262_)
  );


  splt
  gnew_n268_
  (
    .dout(new_n268__spl_),
    .din(new_n268_)
  );


  splt
  gnew_n271_
  (
    .dout(new_n271__spl_),
    .din(new_n271_)
  );


  splt
  gnew_n274_
  (
    .dout(new_n274__spl_),
    .din(new_n274_)
  );


  splt
  gnew_n274__spl_
  (
    .dout(new_n274__spl_0),
    .din(new_n274__spl_)
  );


  splt
  gnew_n274__spl_
  (
    .dout(new_n274__spl_1),
    .din(new_n274__spl_)
  );


  splt
  gnew_n265_
  (
    .dout(new_n265__spl_),
    .din(new_n265_)
  );


  splt
  gnew_n277_
  (
    .dout(new_n277__spl_),
    .din(new_n277_)
  );


  splt
  gnew_n283_
  (
    .dout(new_n283__spl_),
    .din(new_n283_)
  );


  splt
  gnew_n286_
  (
    .dout(new_n286__spl_),
    .din(new_n286_)
  );


  splt
  gnew_n289_
  (
    .dout(new_n289__spl_),
    .din(new_n289_)
  );


  splt
  gnew_n290_
  (
    .dout(new_n290__spl_),
    .din(new_n290_)
  );


  splt
  gnew_n293_
  (
    .dout(new_n293__spl_),
    .din(new_n293_)
  );


  splt
  gnew_n296_
  (
    .dout(new_n296__spl_),
    .din(new_n296_)
  );


  splt
  gnew_n110_
  (
    .dout(new_n110__spl_),
    .din(new_n110_)
  );


  splt
  gnew_n110__spl_
  (
    .dout(new_n110__spl_0),
    .din(new_n110__spl_)
  );


  splt
  gnew_n110__spl_0
  (
    .dout(new_n110__spl_00),
    .din(new_n110__spl_0)
  );


  splt
  gnew_n110__spl_0
  (
    .dout(new_n110__spl_01),
    .din(new_n110__spl_0)
  );


  splt
  gnew_n110__spl_
  (
    .dout(new_n110__spl_1),
    .din(new_n110__spl_)
  );


  splt
  gnew_n110__spl_1
  (
    .dout(new_n110__spl_10),
    .din(new_n110__spl_1)
  );


  splt
  gnew_n299_
  (
    .dout(new_n299__spl_),
    .din(new_n299_)
  );


  splt
  gnew_n299__spl_
  (
    .dout(new_n299__spl_0),
    .din(new_n299__spl_)
  );


  splt
  gnew_n299__spl_0
  (
    .dout(new_n299__spl_00),
    .din(new_n299__spl_0)
  );


  splt
  gnew_n299__spl_0
  (
    .dout(new_n299__spl_01),
    .din(new_n299__spl_0)
  );


  splt
  gnew_n299__spl_
  (
    .dout(new_n299__spl_1),
    .din(new_n299__spl_)
  );


  splt
  gnew_n299__spl_1
  (
    .dout(new_n299__spl_10),
    .din(new_n299__spl_1)
  );


  splt
  gnew_n280_
  (
    .dout(new_n280__spl_),
    .din(new_n280_)
  );


  splt
  gnew_n280__spl_
  (
    .dout(new_n280__spl_0),
    .din(new_n280__spl_)
  );


  splt
  gnew_n280__spl_0
  (
    .dout(new_n280__spl_00),
    .din(new_n280__spl_0)
  );


  splt
  gnew_n280__spl_0
  (
    .dout(new_n280__spl_01),
    .din(new_n280__spl_0)
  );


  splt
  gnew_n280__spl_
  (
    .dout(new_n280__spl_1),
    .din(new_n280__spl_)
  );


  splt
  gnew_n280__spl_1
  (
    .dout(new_n280__spl_10),
    .din(new_n280__spl_1)
  );


  splt
  gnew_n280__spl_1
  (
    .dout(new_n280__spl_11),
    .din(new_n280__spl_1)
  );


  splt
  gnew_n300_
  (
    .dout(new_n300__spl_),
    .din(new_n300_)
  );


  splt
  gnew_n302_
  (
    .dout(new_n302__spl_),
    .din(new_n302_)
  );


  splt
  gnew_n301_
  (
    .dout(new_n301__spl_),
    .din(new_n301_)
  );


  splt
  gnew_n303_
  (
    .dout(new_n303__spl_),
    .din(new_n303_)
  );


  splt
  gnew_n252_
  (
    .dout(new_n252__spl_),
    .din(new_n252_)
  );


  splt
  gnew_n252__spl_
  (
    .dout(new_n252__spl_0),
    .din(new_n252__spl_)
  );


  splt
  gnew_n252__spl_0
  (
    .dout(new_n252__spl_00),
    .din(new_n252__spl_0)
  );


  splt
  gnew_n252__spl_0
  (
    .dout(new_n252__spl_01),
    .din(new_n252__spl_0)
  );


  splt
  gnew_n252__spl_
  (
    .dout(new_n252__spl_1),
    .din(new_n252__spl_)
  );


  splt
  gnew_n252__spl_1
  (
    .dout(new_n252__spl_10),
    .din(new_n252__spl_1)
  );


  splt
  gnew_n252__spl_1
  (
    .dout(new_n252__spl_11),
    .din(new_n252__spl_1)
  );


  splt
  gnew_n306_
  (
    .dout(new_n306__spl_),
    .din(new_n306_)
  );


  splt
  gnew_n306__spl_
  (
    .dout(new_n306__spl_0),
    .din(new_n306__spl_)
  );


  splt
  gnew_n224_
  (
    .dout(new_n224__spl_),
    .din(new_n224_)
  );


  splt
  gnew_n311_
  (
    .dout(new_n311__spl_),
    .din(new_n311_)
  );


  splt
  gnew_n185_
  (
    .dout(new_n185__spl_),
    .din(new_n185_)
  );


  splt
  gnew_n312_
  (
    .dout(new_n312__spl_),
    .din(new_n312_)
  );


  splt
  gnew_n313_
  (
    .dout(new_n313__spl_),
    .din(new_n313_)
  );


  splt
  gnew_n313__spl_
  (
    .dout(new_n313__spl_0),
    .din(new_n313__spl_)
  );


  splt
  gnew_n313__spl_
  (
    .dout(new_n313__spl_1),
    .din(new_n313__spl_)
  );


  splt
  gnew_n314_
  (
    .dout(new_n314__spl_),
    .din(new_n314_)
  );


  splt
  gnew_n318_
  (
    .dout(new_n318__spl_),
    .din(new_n318_)
  );


  splt
  gnew_n322_
  (
    .dout(new_n322__spl_),
    .din(new_n322_)
  );


  splt
  gnew_n326_
  (
    .dout(new_n326__spl_),
    .din(new_n326_)
  );


  splt
  gnew_n330_
  (
    .dout(new_n330__spl_),
    .din(new_n330_)
  );


  splt
  gnew_n331_
  (
    .dout(new_n331__spl_),
    .din(new_n331_)
  );


  splt
  gnew_n332_
  (
    .dout(new_n332__spl_),
    .din(new_n332_)
  );


  splt
  gnew_n332__spl_
  (
    .dout(new_n332__spl_0),
    .din(new_n332__spl_)
  );


  splt
  gnew_n332__spl_
  (
    .dout(new_n332__spl_1),
    .din(new_n332__spl_)
  );


  splt
  gnew_n333_
  (
    .dout(new_n333__spl_),
    .din(new_n333_)
  );


  splt
  gnew_n337_
  (
    .dout(new_n337__spl_),
    .din(new_n337_)
  );


  splt
  gnew_n341_
  (
    .dout(new_n341__spl_),
    .din(new_n341_)
  );


  splt
  gnew_n345_
  (
    .dout(new_n345__spl_),
    .din(new_n345_)
  );


  splt
  gnew_n349_
  (
    .dout(new_n349__spl_),
    .din(new_n349_)
  );


  splt
  gnew_n350_
  (
    .dout(new_n350__spl_),
    .din(new_n350_)
  );


  splt
  gnew_n350__spl_
  (
    .dout(new_n350__spl_0),
    .din(new_n350__spl_)
  );


  splt
  gnew_n350__spl_
  (
    .dout(new_n350__spl_1),
    .din(new_n350__spl_)
  );


  splt
  gnew_n351_
  (
    .dout(new_n351__spl_),
    .din(new_n351_)
  );


  splt
  gnew_n355_
  (
    .dout(new_n355__spl_),
    .din(new_n355_)
  );


  splt
  gnew_n359_
  (
    .dout(new_n359__spl_),
    .din(new_n359_)
  );


  splt
  gnew_n363_
  (
    .dout(new_n363__spl_),
    .din(new_n363_)
  );


  splt
  gnew_n367_
  (
    .dout(new_n367__spl_),
    .din(new_n367_)
  );


  splt
  gnew_n368_
  (
    .dout(new_n368__spl_),
    .din(new_n368_)
  );


  splt
  gnew_n368__spl_
  (
    .dout(new_n368__spl_0),
    .din(new_n368__spl_)
  );


  splt
  gnew_n368__spl_
  (
    .dout(new_n368__spl_1),
    .din(new_n368__spl_)
  );


  splt
  gnew_n369_
  (
    .dout(new_n369__spl_),
    .din(new_n369_)
  );


  splt
  gnew_n373_
  (
    .dout(new_n373__spl_),
    .din(new_n373_)
  );


  splt
  gnew_n377_
  (
    .dout(new_n377__spl_),
    .din(new_n377_)
  );


  splt
  gnew_n381_
  (
    .dout(new_n381__spl_),
    .din(new_n381_)
  );


  splt
  gnew_n391_
  (
    .dout(new_n391__spl_),
    .din(new_n391_)
  );


  splt
  gnew_n391__spl_
  (
    .dout(new_n391__spl_0),
    .din(new_n391__spl_)
  );


  splt
  gnew_n393_
  (
    .dout(new_n393__spl_),
    .din(new_n393_)
  );


  splt
  gnew_n393__spl_
  (
    .dout(new_n393__spl_0),
    .din(new_n393__spl_)
  );


  splt
  gnew_n393__spl_
  (
    .dout(new_n393__spl_1),
    .din(new_n393__spl_)
  );


  splt
  gnew_n394_
  (
    .dout(new_n394__spl_),
    .din(new_n394_)
  );


  splt
  gnew_n398_
  (
    .dout(new_n398__spl_),
    .din(new_n398_)
  );


  splt
  gnew_n402_
  (
    .dout(new_n402__spl_),
    .din(new_n402_)
  );


  splt
  gnew_n406_
  (
    .dout(new_n406__spl_),
    .din(new_n406_)
  );


  splt
  gnew_n410_
  (
    .dout(new_n410__spl_),
    .din(new_n410_)
  );


  splt
  gnew_n411_
  (
    .dout(new_n411__spl_),
    .din(new_n411_)
  );


  splt
  gnew_n411__spl_
  (
    .dout(new_n411__spl_0),
    .din(new_n411__spl_)
  );


  splt
  gnew_n411__spl_
  (
    .dout(new_n411__spl_1),
    .din(new_n411__spl_)
  );


  splt
  gnew_n412_
  (
    .dout(new_n412__spl_),
    .din(new_n412_)
  );


  splt
  gnew_n416_
  (
    .dout(new_n416__spl_),
    .din(new_n416_)
  );


  splt
  gnew_n420_
  (
    .dout(new_n420__spl_),
    .din(new_n420_)
  );


  splt
  gnew_n424_
  (
    .dout(new_n424__spl_),
    .din(new_n424_)
  );


  splt
  gnew_n429_
  (
    .dout(new_n429__spl_),
    .din(new_n429_)
  );


  splt
  gnew_n429__spl_
  (
    .dout(new_n429__spl_0),
    .din(new_n429__spl_)
  );


  splt
  gnew_n429__spl_
  (
    .dout(new_n429__spl_1),
    .din(new_n429__spl_)
  );


  splt
  gnew_n430_
  (
    .dout(new_n430__spl_),
    .din(new_n430_)
  );


  splt
  gnew_n434_
  (
    .dout(new_n434__spl_),
    .din(new_n434_)
  );


  splt
  gnew_n438_
  (
    .dout(new_n438__spl_),
    .din(new_n438_)
  );


  splt
  gnew_n442_
  (
    .dout(new_n442__spl_),
    .din(new_n442_)
  );


  splt
  gnew_n446_
  (
    .dout(new_n446__spl_),
    .din(new_n446_)
  );


  splt
  gnew_n446__spl_
  (
    .dout(new_n446__spl_0),
    .din(new_n446__spl_)
  );


  splt
  gnew_n446__spl_
  (
    .dout(new_n446__spl_1),
    .din(new_n446__spl_)
  );


  splt
  gnew_n447_
  (
    .dout(new_n447__spl_),
    .din(new_n447_)
  );


  splt
  gnew_n451_
  (
    .dout(new_n451__spl_),
    .din(new_n451_)
  );


  splt
  gnew_n455_
  (
    .dout(new_n455__spl_),
    .din(new_n455_)
  );


  splt
  gnew_n459_
  (
    .dout(new_n459__spl_),
    .din(new_n459_)
  );


endmodule
