
module mymod
(
  G1,
  G2,
  G3,
  G4,
  G5,
  G6,
  G7,
  G8,
  G9,
  G10,
  G11,
  G12,
  G13,
  G14,
  G15,
  G16,
  G17,
  G18,
  G19,
  G20,
  G21,
  G22,
  G23,
  G24,
  G25,
  G26,
  G27,
  G28,
  G29,
  G30,
  G31,
  G32,
  G6257,
  G6258,
  G6259,
  G6260,
  G6261,
  G6262,
  G6263,
  G6264,
  G6265,
  G6266,
  G6267,
  G6268,
  G6269,
  G6270,
  G6271,
  G6272,
  G6273,
  G6274,
  G6275,
  G6276,
  G6277,
  G6278,
  G6279,
  G6280,
  G6281,
  G6282,
  G6283,
  G6284,
  G6285,
  G6286,
  G6287,
  G6288
);

  input G1;input G2;input G3;input G4;input G5;input G6;input G7;input G8;input G9;input G10;input G11;input G12;input G13;input G14;input G15;input G16;input G17;input G18;input G19;input G20;input G21;input G22;input G23;input G24;input G25;input G26;input G27;input G28;input G29;input G30;input G31;input G32;
  output G6257;output G6258;output G6259;output G6260;output G6261;output G6262;output G6263;output G6264;output G6265;output G6266;output G6267;output G6268;output G6269;output G6270;output G6271;output G6272;output G6273;output G6274;output G6275;output G6276;output G6277;output G6278;output G6279;output G6280;output G6281;output G6282;output G6283;output G6284;output G6285;output G6286;output G6287;output G6288;
  wire G1_p;
  wire G1_n;
  wire G2_p;
  wire G2_n;
  wire G3_p;
  wire G3_n;
  wire G4_p;
  wire G4_n;
  wire G5_p;
  wire G5_n;
  wire G6_p;
  wire G6_n;
  wire G7_p;
  wire G7_n;
  wire G8_p;
  wire G8_n;
  wire G9_p;
  wire G9_n;
  wire G10_p;
  wire G10_n;
  wire G11_p;
  wire G11_n;
  wire G12_p;
  wire G12_n;
  wire G13_p;
  wire G13_n;
  wire G14_p;
  wire G14_n;
  wire G15_p;
  wire G15_n;
  wire G16_p;
  wire G16_n;
  wire G17_p;
  wire G17_n;
  wire G18_p;
  wire G18_n;
  wire G19_p;
  wire G19_n;
  wire G20_p;
  wire G20_n;
  wire G21_p;
  wire G21_n;
  wire G22_p;
  wire G22_n;
  wire G23_p;
  wire G23_n;
  wire G24_p;
  wire G24_n;
  wire G25_p;
  wire G25_n;
  wire G26_p;
  wire G26_n;
  wire G27_p;
  wire G27_n;
  wire G28_p;
  wire G28_n;
  wire G29_p;
  wire G29_n;
  wire G30_p;
  wire G30_n;
  wire G31_p;
  wire G31_n;
  wire G32_p;
  wire G32_n;
  wire g33_p;
  wire g33_n;
  wire g34_p;
  wire g34_n;
  wire g35_p;
  wire g35_n;
  wire g36_p;
  wire g36_n;
  wire g37_p;
  wire g37_n;
  wire g38_p;
  wire g38_n;
  wire g39_p;
  wire g39_n;
  wire g40_p;
  wire g40_n;
  wire g41_p;
  wire g41_n;
  wire g42_p;
  wire g42_n;
  wire g43_p;
  wire g43_n;
  wire g44_p;
  wire g44_n;
  wire g45_p;
  wire g45_n;
  wire g46_p;
  wire g46_n;
  wire g47_p;
  wire g47_n;
  wire g48_p;
  wire g48_n;
  wire g49_p;
  wire g49_n;
  wire g50_p;
  wire g50_n;
  wire g51_p;
  wire g51_n;
  wire g52_p;
  wire g52_n;
  wire g53_p;
  wire g53_n;
  wire g54_p;
  wire g54_n;
  wire g55_p;
  wire g55_n;
  wire g56_p;
  wire g56_n;
  wire g57_p;
  wire g57_n;
  wire g58_p;
  wire g58_n;
  wire g59_p;
  wire g59_n;
  wire g60_p;
  wire g60_n;
  wire g61_p;
  wire g61_n;
  wire g62_p;
  wire g62_n;
  wire g63_p;
  wire g63_n;
  wire g64_p;
  wire g64_n;
  wire g65_p;
  wire g65_n;
  wire g66_p;
  wire g66_n;
  wire g67_p;
  wire g67_n;
  wire g68_p;
  wire g68_n;
  wire g69_p;
  wire g69_n;
  wire g70_p;
  wire g70_n;
  wire g71_p;
  wire g71_n;
  wire g72_p;
  wire g72_n;
  wire g73_p;
  wire g73_n;
  wire g74_p;
  wire g74_n;
  wire g75_p;
  wire g75_n;
  wire g76_p;
  wire g76_n;
  wire g77_p;
  wire g77_n;
  wire g78_p;
  wire g78_n;
  wire g79_p;
  wire g79_n;
  wire g80_p;
  wire g80_n;
  wire g81_p;
  wire g81_n;
  wire g82_p;
  wire g82_n;
  wire g83_p;
  wire g83_n;
  wire g84_p;
  wire g84_n;
  wire g85_p;
  wire g85_n;
  wire g86_p;
  wire g86_n;
  wire g87_p;
  wire g87_n;
  wire g88_p;
  wire g88_n;
  wire g89_p;
  wire g89_n;
  wire g90_p;
  wire g90_n;
  wire g91_p;
  wire g91_n;
  wire g92_p;
  wire g92_n;
  wire g93_p;
  wire g93_n;
  wire g94_p;
  wire g94_n;
  wire g95_p;
  wire g95_n;
  wire g96_p;
  wire g96_n;
  wire g97_p;
  wire g97_n;
  wire g98_p;
  wire g98_n;
  wire g99_p;
  wire g99_n;
  wire g100_p;
  wire g100_n;
  wire g101_p;
  wire g101_n;
  wire g102_p;
  wire g102_n;
  wire g103_p;
  wire g103_n;
  wire g104_p;
  wire g104_n;
  wire g105_p;
  wire g105_n;
  wire g106_p;
  wire g106_n;
  wire g107_p;
  wire g107_n;
  wire g108_p;
  wire g108_n;
  wire g109_p;
  wire g109_n;
  wire g110_p;
  wire g110_n;
  wire g111_p;
  wire g111_n;
  wire g112_p;
  wire g112_n;
  wire g113_p;
  wire g113_n;
  wire g114_p;
  wire g114_n;
  wire g115_p;
  wire g115_n;
  wire g116_p;
  wire g116_n;
  wire g117_p;
  wire g117_n;
  wire g118_p;
  wire g118_n;
  wire g119_p;
  wire g119_n;
  wire g120_p;
  wire g120_n;
  wire g121_p;
  wire g121_n;
  wire g122_p;
  wire g122_n;
  wire g123_p;
  wire g123_n;
  wire g124_p;
  wire g124_n;
  wire g125_p;
  wire g125_n;
  wire g126_p;
  wire g126_n;
  wire g127_p;
  wire g127_n;
  wire g128_p;
  wire g128_n;
  wire g129_p;
  wire g129_n;
  wire g130_p;
  wire g130_n;
  wire g131_p;
  wire g131_n;
  wire g132_p;
  wire g132_n;
  wire g133_p;
  wire g133_n;
  wire g134_p;
  wire g134_n;
  wire g135_p;
  wire g135_n;
  wire g136_p;
  wire g136_n;
  wire g137_p;
  wire g137_n;
  wire g138_p;
  wire g138_n;
  wire g139_p;
  wire g139_n;
  wire g140_p;
  wire g140_n;
  wire g141_p;
  wire g141_n;
  wire g142_p;
  wire g142_n;
  wire g143_p;
  wire g143_n;
  wire g144_p;
  wire g144_n;
  wire g145_p;
  wire g145_n;
  wire g146_p;
  wire g146_n;
  wire g147_p;
  wire g147_n;
  wire g148_p;
  wire g148_n;
  wire g149_p;
  wire g149_n;
  wire g150_p;
  wire g150_n;
  wire g151_p;
  wire g151_n;
  wire g152_p;
  wire g152_n;
  wire g153_p;
  wire g153_n;
  wire g154_p;
  wire g154_n;
  wire g155_p;
  wire g155_n;
  wire g156_p;
  wire g156_n;
  wire g157_p;
  wire g157_n;
  wire g158_p;
  wire g158_n;
  wire g159_p;
  wire g159_n;
  wire g160_p;
  wire g160_n;
  wire g161_p;
  wire g161_n;
  wire g162_p;
  wire g162_n;
  wire g163_p;
  wire g163_n;
  wire g164_p;
  wire g164_n;
  wire g165_p;
  wire g165_n;
  wire g166_p;
  wire g166_n;
  wire g167_p;
  wire g167_n;
  wire g168_p;
  wire g168_n;
  wire g169_p;
  wire g169_n;
  wire g170_p;
  wire g170_n;
  wire g171_p;
  wire g171_n;
  wire g172_p;
  wire g172_n;
  wire g173_p;
  wire g173_n;
  wire g174_p;
  wire g174_n;
  wire g175_p;
  wire g175_n;
  wire g176_p;
  wire g176_n;
  wire g177_p;
  wire g177_n;
  wire g178_p;
  wire g178_n;
  wire g179_p;
  wire g179_n;
  wire g180_p;
  wire g180_n;
  wire g181_p;
  wire g181_n;
  wire g182_p;
  wire g182_n;
  wire g183_p;
  wire g183_n;
  wire g184_p;
  wire g184_n;
  wire g185_p;
  wire g185_n;
  wire g186_p;
  wire g186_n;
  wire g187_p;
  wire g187_n;
  wire g188_p;
  wire g188_n;
  wire g189_p;
  wire g189_n;
  wire g190_p;
  wire g190_n;
  wire g191_p;
  wire g191_n;
  wire g192_p;
  wire g192_n;
  wire g193_p;
  wire g193_n;
  wire g194_p;
  wire g194_n;
  wire g195_p;
  wire g195_n;
  wire g196_p;
  wire g196_n;
  wire g197_p;
  wire g197_n;
  wire g198_p;
  wire g198_n;
  wire g199_p;
  wire g199_n;
  wire g200_p;
  wire g200_n;
  wire g201_p;
  wire g201_n;
  wire g202_p;
  wire g202_n;
  wire g203_p;
  wire g203_n;
  wire g204_p;
  wire g204_n;
  wire g205_p;
  wire g205_n;
  wire g206_p;
  wire g206_n;
  wire g207_p;
  wire g207_n;
  wire g208_p;
  wire g208_n;
  wire g209_p;
  wire g209_n;
  wire g210_p;
  wire g210_n;
  wire g211_p;
  wire g211_n;
  wire g212_p;
  wire g212_n;
  wire g213_p;
  wire g213_n;
  wire g214_p;
  wire g214_n;
  wire g215_p;
  wire g215_n;
  wire g216_p;
  wire g216_n;
  wire g217_p;
  wire g217_n;
  wire g218_p;
  wire g218_n;
  wire g219_p;
  wire g219_n;
  wire g220_p;
  wire g220_n;
  wire g221_p;
  wire g221_n;
  wire g222_p;
  wire g222_n;
  wire g223_p;
  wire g223_n;
  wire g224_p;
  wire g224_n;
  wire g225_p;
  wire g225_n;
  wire g226_p;
  wire g226_n;
  wire g227_p;
  wire g227_n;
  wire g228_p;
  wire g228_n;
  wire g229_p;
  wire g229_n;
  wire g230_p;
  wire g230_n;
  wire g231_p;
  wire g231_n;
  wire g232_p;
  wire g232_n;
  wire g233_p;
  wire g233_n;
  wire g234_p;
  wire g234_n;
  wire g235_p;
  wire g235_n;
  wire g236_p;
  wire g236_n;
  wire g237_p;
  wire g237_n;
  wire g238_p;
  wire g238_n;
  wire g239_p;
  wire g239_n;
  wire g240_p;
  wire g240_n;
  wire g241_p;
  wire g241_n;
  wire g242_p;
  wire g242_n;
  wire g243_p;
  wire g243_n;
  wire g244_p;
  wire g244_n;
  wire g245_p;
  wire g245_n;
  wire g246_p;
  wire g246_n;
  wire g247_p;
  wire g247_n;
  wire g248_p;
  wire g248_n;
  wire g249_p;
  wire g249_n;
  wire g250_p;
  wire g250_n;
  wire g251_p;
  wire g251_n;
  wire g252_p;
  wire g252_n;
  wire g253_p;
  wire g253_n;
  wire g254_p;
  wire g254_n;
  wire g255_p;
  wire g255_n;
  wire g256_p;
  wire g256_n;
  wire g257_p;
  wire g257_n;
  wire g258_p;
  wire g258_n;
  wire g259_p;
  wire g259_n;
  wire g260_p;
  wire g260_n;
  wire g261_p;
  wire g261_n;
  wire g262_p;
  wire g262_n;
  wire g263_p;
  wire g263_n;
  wire g264_p;
  wire g264_n;
  wire g265_p;
  wire g265_n;
  wire g266_p;
  wire g266_n;
  wire g267_p;
  wire g267_n;
  wire g268_p;
  wire g268_n;
  wire g269_p;
  wire g269_n;
  wire g270_p;
  wire g270_n;
  wire g271_p;
  wire g271_n;
  wire g272_p;
  wire g272_n;
  wire g273_p;
  wire g273_n;
  wire g274_p;
  wire g274_n;
  wire g275_p;
  wire g275_n;
  wire g276_p;
  wire g276_n;
  wire g277_p;
  wire g277_n;
  wire g278_p;
  wire g278_n;
  wire g279_p;
  wire g279_n;
  wire g280_p;
  wire g280_n;
  wire g281_p;
  wire g281_n;
  wire g282_p;
  wire g282_n;
  wire g283_p;
  wire g283_n;
  wire g284_p;
  wire g284_n;
  wire g285_p;
  wire g285_n;
  wire g286_p;
  wire g286_n;
  wire g287_p;
  wire g287_n;
  wire g288_p;
  wire g288_n;
  wire g289_p;
  wire g289_n;
  wire g290_p;
  wire g290_n;
  wire g291_p;
  wire g291_n;
  wire g292_p;
  wire g292_n;
  wire g293_p;
  wire g293_n;
  wire g294_p;
  wire g294_n;
  wire g295_p;
  wire g295_n;
  wire g296_p;
  wire g296_n;
  wire g297_p;
  wire g297_n;
  wire g298_p;
  wire g298_n;
  wire g299_p;
  wire g299_n;
  wire g300_p;
  wire g300_n;
  wire g301_p;
  wire g301_n;
  wire g302_p;
  wire g302_n;
  wire g303_p;
  wire g303_n;
  wire g304_p;
  wire g304_n;
  wire g305_p;
  wire g305_n;
  wire g306_p;
  wire g306_n;
  wire g307_p;
  wire g307_n;
  wire g308_p;
  wire g308_n;
  wire g309_p;
  wire g309_n;
  wire g310_p;
  wire g310_n;
  wire g311_p;
  wire g311_n;
  wire g312_p;
  wire g312_n;
  wire g313_p;
  wire g313_n;
  wire g314_p;
  wire g314_n;
  wire g315_p;
  wire g315_n;
  wire g316_p;
  wire g316_n;
  wire g317_p;
  wire g317_n;
  wire g318_p;
  wire g318_n;
  wire g319_p;
  wire g319_n;
  wire g320_p;
  wire g320_n;
  wire g321_p;
  wire g321_n;
  wire g322_p;
  wire g322_n;
  wire g323_p;
  wire g323_n;
  wire g324_p;
  wire g324_n;
  wire g325_p;
  wire g325_n;
  wire g326_p;
  wire g326_n;
  wire g327_p;
  wire g327_n;
  wire g328_p;
  wire g328_n;
  wire g329_p;
  wire g329_n;
  wire g330_p;
  wire g330_n;
  wire g331_p;
  wire g331_n;
  wire g332_p;
  wire g332_n;
  wire g333_p;
  wire g333_n;
  wire g334_p;
  wire g334_n;
  wire g335_p;
  wire g335_n;
  wire g336_p;
  wire g336_n;
  wire g337_p;
  wire g337_n;
  wire g338_p;
  wire g338_n;
  wire g339_p;
  wire g339_n;
  wire g340_p;
  wire g340_n;
  wire g341_p;
  wire g341_n;
  wire g342_p;
  wire g342_n;
  wire g343_p;
  wire g343_n;
  wire g344_p;
  wire g344_n;
  wire g345_p;
  wire g345_n;
  wire g346_p;
  wire g346_n;
  wire g347_p;
  wire g347_n;
  wire g348_p;
  wire g348_n;
  wire g349_p;
  wire g349_n;
  wire g350_p;
  wire g350_n;
  wire g351_p;
  wire g351_n;
  wire g352_p;
  wire g352_n;
  wire g353_p;
  wire g353_n;
  wire g354_p;
  wire g354_n;
  wire g355_p;
  wire g355_n;
  wire g356_p;
  wire g356_n;
  wire g357_p;
  wire g357_n;
  wire g358_p;
  wire g358_n;
  wire g359_p;
  wire g359_n;
  wire g360_p;
  wire g360_n;
  wire g361_p;
  wire g361_n;
  wire g362_p;
  wire g362_n;
  wire g363_p;
  wire g363_n;
  wire g364_p;
  wire g364_n;
  wire g365_p;
  wire g365_n;
  wire g366_p;
  wire g366_n;
  wire g367_p;
  wire g367_n;
  wire g368_p;
  wire g368_n;
  wire g369_p;
  wire g369_n;
  wire g370_p;
  wire g370_n;
  wire g371_p;
  wire g371_n;
  wire g372_p;
  wire g372_n;
  wire g373_p;
  wire g373_n;
  wire g374_p;
  wire g374_n;
  wire g375_p;
  wire g375_n;
  wire g376_p;
  wire g376_n;
  wire g377_p;
  wire g377_n;
  wire g378_p;
  wire g378_n;
  wire g379_p;
  wire g379_n;
  wire g380_p;
  wire g380_n;
  wire g381_p;
  wire g381_n;
  wire g382_p;
  wire g382_n;
  wire g383_p;
  wire g383_n;
  wire g384_p;
  wire g384_n;
  wire g385_p;
  wire g385_n;
  wire g386_p;
  wire g386_n;
  wire g387_p;
  wire g387_n;
  wire g388_p;
  wire g388_n;
  wire g389_p;
  wire g389_n;
  wire g390_p;
  wire g390_n;
  wire g391_p;
  wire g391_n;
  wire g392_p;
  wire g392_n;
  wire g393_p;
  wire g393_n;
  wire g394_p;
  wire g394_n;
  wire g395_p;
  wire g395_n;
  wire g396_p;
  wire g396_n;
  wire g397_p;
  wire g397_n;
  wire g398_p;
  wire g398_n;
  wire g399_p;
  wire g399_n;
  wire g400_p;
  wire g400_n;
  wire g401_p;
  wire g401_n;
  wire g402_p;
  wire g402_n;
  wire g403_p;
  wire g403_n;
  wire g404_p;
  wire g404_n;
  wire g405_p;
  wire g405_n;
  wire g406_p;
  wire g406_n;
  wire g407_p;
  wire g407_n;
  wire g408_p;
  wire g408_n;
  wire g409_p;
  wire g409_n;
  wire g410_p;
  wire g410_n;
  wire g411_p;
  wire g411_n;
  wire g412_p;
  wire g412_n;
  wire g413_p;
  wire g413_n;
  wire g414_p;
  wire g414_n;
  wire g415_p;
  wire g415_n;
  wire g416_p;
  wire g416_n;
  wire g417_p;
  wire g417_n;
  wire g418_p;
  wire g418_n;
  wire g419_p;
  wire g419_n;
  wire g420_p;
  wire g420_n;
  wire g421_p;
  wire g421_n;
  wire g422_p;
  wire g422_n;
  wire g423_p;
  wire g423_n;
  wire g424_p;
  wire g424_n;
  wire g425_p;
  wire g425_n;
  wire g426_p;
  wire g426_n;
  wire g427_p;
  wire g427_n;
  wire g428_p;
  wire g428_n;
  wire g429_p;
  wire g429_n;
  wire g430_p;
  wire g430_n;
  wire g431_p;
  wire g431_n;
  wire g432_p;
  wire g432_n;
  wire g433_p;
  wire g433_n;
  wire g434_p;
  wire g434_n;
  wire g435_p;
  wire g435_n;
  wire g436_p;
  wire g436_n;
  wire g437_p;
  wire g437_n;
  wire g438_p;
  wire g438_n;
  wire g439_p;
  wire g439_n;
  wire g440_p;
  wire g440_n;
  wire g441_p;
  wire g441_n;
  wire g442_p;
  wire g442_n;
  wire g443_p;
  wire g443_n;
  wire g444_p;
  wire g444_n;
  wire g445_p;
  wire g445_n;
  wire g446_p;
  wire g446_n;
  wire g447_p;
  wire g447_n;
  wire g448_p;
  wire g448_n;
  wire g449_p;
  wire g449_n;
  wire g450_p;
  wire g450_n;
  wire g451_p;
  wire g451_n;
  wire g452_p;
  wire g452_n;
  wire g453_p;
  wire g453_n;
  wire g454_p;
  wire g454_n;
  wire g455_p;
  wire g455_n;
  wire g456_p;
  wire g456_n;
  wire g457_p;
  wire g457_n;
  wire g458_p;
  wire g458_n;
  wire g459_p;
  wire g459_n;
  wire g460_p;
  wire g460_n;
  wire g461_p;
  wire g461_n;
  wire g462_p;
  wire g462_n;
  wire g463_p;
  wire g463_n;
  wire g464_p;
  wire g464_n;
  wire g465_p;
  wire g465_n;
  wire g466_p;
  wire g466_n;
  wire g467_p;
  wire g467_n;
  wire g468_p;
  wire g468_n;
  wire g469_p;
  wire g469_n;
  wire g470_p;
  wire g470_n;
  wire g471_p;
  wire g471_n;
  wire g472_p;
  wire g472_n;
  wire g473_p;
  wire g473_n;
  wire g474_p;
  wire g474_n;
  wire g475_p;
  wire g475_n;
  wire g476_p;
  wire g476_n;
  wire g477_p;
  wire g477_n;
  wire g478_p;
  wire g478_n;
  wire g479_p;
  wire g479_n;
  wire g480_p;
  wire g480_n;
  wire g481_p;
  wire g481_n;
  wire g482_p;
  wire g482_n;
  wire g483_p;
  wire g483_n;
  wire g484_p;
  wire g484_n;
  wire g485_p;
  wire g485_n;
  wire g486_p;
  wire g486_n;
  wire g487_p;
  wire g487_n;
  wire g488_p;
  wire g488_n;
  wire g489_p;
  wire g489_n;
  wire g490_p;
  wire g490_n;
  wire g491_p;
  wire g491_n;
  wire g492_p;
  wire g492_n;
  wire g493_p;
  wire g493_n;
  wire g494_p;
  wire g494_n;
  wire g495_p;
  wire g495_n;
  wire g496_p;
  wire g496_n;
  wire g497_p;
  wire g497_n;
  wire g498_p;
  wire g498_n;
  wire g499_p;
  wire g499_n;
  wire g500_p;
  wire g500_n;
  wire g501_p;
  wire g501_n;
  wire g502_p;
  wire g502_n;
  wire g503_p;
  wire g503_n;
  wire g504_p;
  wire g504_n;
  wire g505_p;
  wire g505_n;
  wire g506_p;
  wire g506_n;
  wire g507_p;
  wire g507_n;
  wire g508_p;
  wire g508_n;
  wire g509_p;
  wire g509_n;
  wire g510_p;
  wire g510_n;
  wire g511_p;
  wire g511_n;
  wire g512_p;
  wire g512_n;
  wire g513_p;
  wire g513_n;
  wire g514_p;
  wire g514_n;
  wire g515_p;
  wire g515_n;
  wire g516_p;
  wire g516_n;
  wire g517_p;
  wire g517_n;
  wire g518_p;
  wire g518_n;
  wire g519_p;
  wire g519_n;
  wire g520_p;
  wire g520_n;
  wire g521_p;
  wire g521_n;
  wire g522_p;
  wire g522_n;
  wire g523_p;
  wire g523_n;
  wire g524_p;
  wire g524_n;
  wire g525_p;
  wire g525_n;
  wire g526_p;
  wire g526_n;
  wire g527_p;
  wire g527_n;
  wire g528_p;
  wire g528_n;
  wire g529_p;
  wire g529_n;
  wire g530_p;
  wire g530_n;
  wire g531_p;
  wire g531_n;
  wire g532_p;
  wire g532_n;
  wire g533_p;
  wire g533_n;
  wire g534_p;
  wire g534_n;
  wire g535_p;
  wire g535_n;
  wire g536_p;
  wire g536_n;
  wire g537_p;
  wire g537_n;
  wire g538_p;
  wire g538_n;
  wire g539_p;
  wire g539_n;
  wire g540_p;
  wire g540_n;
  wire g541_p;
  wire g541_n;
  wire g542_p;
  wire g542_n;
  wire g543_p;
  wire g543_n;
  wire g544_p;
  wire g544_n;
  wire g545_p;
  wire g545_n;
  wire g546_p;
  wire g546_n;
  wire g547_p;
  wire g547_n;
  wire g548_p;
  wire g548_n;
  wire g549_p;
  wire g549_n;
  wire g550_p;
  wire g550_n;
  wire g551_p;
  wire g551_n;
  wire g552_p;
  wire g552_n;
  wire g553_p;
  wire g553_n;
  wire g554_p;
  wire g554_n;
  wire g555_p;
  wire g555_n;
  wire g556_p;
  wire g556_n;
  wire g557_p;
  wire g557_n;
  wire g558_p;
  wire g558_n;
  wire g559_p;
  wire g559_n;
  wire g560_p;
  wire g560_n;
  wire g561_p;
  wire g561_n;
  wire g562_p;
  wire g562_n;
  wire g563_p;
  wire g563_n;
  wire g564_p;
  wire g564_n;
  wire g565_p;
  wire g565_n;
  wire g566_p;
  wire g566_n;
  wire g567_p;
  wire g567_n;
  wire g568_p;
  wire g568_n;
  wire g569_p;
  wire g569_n;
  wire g570_p;
  wire g570_n;
  wire g571_p;
  wire g571_n;
  wire g572_p;
  wire g572_n;
  wire g573_p;
  wire g573_n;
  wire g574_p;
  wire g574_n;
  wire g575_p;
  wire g575_n;
  wire g576_p;
  wire g576_n;
  wire g577_p;
  wire g577_n;
  wire g578_p;
  wire g578_n;
  wire g579_p;
  wire g579_n;
  wire g580_p;
  wire g580_n;
  wire g581_p;
  wire g581_n;
  wire g582_p;
  wire g582_n;
  wire g583_p;
  wire g583_n;
  wire g584_p;
  wire g584_n;
  wire g585_p;
  wire g585_n;
  wire g586_p;
  wire g586_n;
  wire g587_p;
  wire g587_n;
  wire g588_p;
  wire g588_n;
  wire g589_p;
  wire g589_n;
  wire g590_p;
  wire g590_n;
  wire g591_p;
  wire g591_n;
  wire g592_p;
  wire g592_n;
  wire g593_p;
  wire g593_n;
  wire g594_p;
  wire g594_n;
  wire g595_p;
  wire g595_n;
  wire g596_p;
  wire g596_n;
  wire g597_p;
  wire g597_n;
  wire g598_p;
  wire g598_n;
  wire g599_p;
  wire g599_n;
  wire g600_p;
  wire g600_n;
  wire g601_p;
  wire g601_n;
  wire g602_p;
  wire g602_n;
  wire g603_p;
  wire g603_n;
  wire g604_p;
  wire g604_n;
  wire g605_p;
  wire g605_n;
  wire g606_p;
  wire g606_n;
  wire g607_p;
  wire g607_n;
  wire g608_p;
  wire g608_n;
  wire g609_p;
  wire g609_n;
  wire g610_p;
  wire g610_n;
  wire g611_p;
  wire g611_n;
  wire g612_p;
  wire g612_n;
  wire g613_p;
  wire g613_n;
  wire g614_p;
  wire g614_n;
  wire g615_p;
  wire g615_n;
  wire g616_p;
  wire g616_n;
  wire g617_p;
  wire g617_n;
  wire g618_p;
  wire g618_n;
  wire g619_p;
  wire g619_n;
  wire g620_p;
  wire g620_n;
  wire g621_p;
  wire g621_n;
  wire g622_p;
  wire g622_n;
  wire g623_p;
  wire g623_n;
  wire g624_p;
  wire g624_n;
  wire g625_p;
  wire g625_n;
  wire g626_p;
  wire g626_n;
  wire g627_p;
  wire g627_n;
  wire g628_p;
  wire g628_n;
  wire g629_p;
  wire g629_n;
  wire g630_p;
  wire g630_n;
  wire g631_p;
  wire g631_n;
  wire g632_p;
  wire g632_n;
  wire g633_p;
  wire g633_n;
  wire g634_p;
  wire g634_n;
  wire g635_p;
  wire g635_n;
  wire g636_p;
  wire g636_n;
  wire g637_p;
  wire g637_n;
  wire g638_p;
  wire g638_n;
  wire g639_p;
  wire g639_n;
  wire g640_p;
  wire g640_n;
  wire g641_p;
  wire g641_n;
  wire g642_p;
  wire g642_n;
  wire g643_p;
  wire g643_n;
  wire g644_p;
  wire g644_n;
  wire g645_p;
  wire g645_n;
  wire g646_p;
  wire g646_n;
  wire g647_p;
  wire g647_n;
  wire g648_p;
  wire g648_n;
  wire g649_p;
  wire g649_n;
  wire g650_p;
  wire g650_n;
  wire g651_p;
  wire g651_n;
  wire g652_p;
  wire g652_n;
  wire g653_p;
  wire g653_n;
  wire g654_p;
  wire g654_n;
  wire g655_p;
  wire g655_n;
  wire g656_p;
  wire g656_n;
  wire g657_p;
  wire g657_n;
  wire g658_p;
  wire g658_n;
  wire g659_p;
  wire g659_n;
  wire g660_p;
  wire g660_n;
  wire g661_p;
  wire g661_n;
  wire g662_p;
  wire g662_n;
  wire g663_p;
  wire g663_n;
  wire g664_p;
  wire g664_n;
  wire g665_p;
  wire g665_n;
  wire g666_p;
  wire g666_n;
  wire g667_p;
  wire g667_n;
  wire g668_p;
  wire g668_n;
  wire g669_p;
  wire g669_n;
  wire g670_p;
  wire g670_n;
  wire g671_p;
  wire g671_n;
  wire g672_p;
  wire g672_n;
  wire g673_p;
  wire g673_n;
  wire g674_p;
  wire g674_n;
  wire g675_p;
  wire g675_n;
  wire g676_p;
  wire g676_n;
  wire g677_p;
  wire g677_n;
  wire g678_p;
  wire g678_n;
  wire g679_p;
  wire g679_n;
  wire g680_p;
  wire g680_n;
  wire g681_p;
  wire g681_n;
  wire g682_p;
  wire g682_n;
  wire g683_p;
  wire g683_n;
  wire g684_p;
  wire g684_n;
  wire g685_p;
  wire g685_n;
  wire g686_p;
  wire g686_n;
  wire g687_p;
  wire g687_n;
  wire g688_p;
  wire g688_n;
  wire g689_p;
  wire g689_n;
  wire g690_p;
  wire g690_n;
  wire g691_p;
  wire g691_n;
  wire g692_p;
  wire g692_n;
  wire g693_p;
  wire g693_n;
  wire g694_p;
  wire g694_n;
  wire g695_p;
  wire g695_n;
  wire g696_p;
  wire g696_n;
  wire g697_p;
  wire g697_n;
  wire g698_p;
  wire g698_n;
  wire g699_p;
  wire g699_n;
  wire g700_p;
  wire g700_n;
  wire g701_p;
  wire g701_n;
  wire g702_p;
  wire g702_n;
  wire g703_p;
  wire g703_n;
  wire g704_p;
  wire g704_n;
  wire g705_p;
  wire g705_n;
  wire g706_p;
  wire g706_n;
  wire g707_p;
  wire g707_n;
  wire g708_p;
  wire g708_n;
  wire g709_p;
  wire g709_n;
  wire g710_p;
  wire g710_n;
  wire g711_p;
  wire g711_n;
  wire g712_p;
  wire g712_n;
  wire g713_p;
  wire g713_n;
  wire g714_p;
  wire g714_n;
  wire g715_p;
  wire g715_n;
  wire g716_p;
  wire g716_n;
  wire g717_p;
  wire g717_n;
  wire g718_p;
  wire g718_n;
  wire g719_p;
  wire g719_n;
  wire g720_p;
  wire g720_n;
  wire g721_p;
  wire g721_n;
  wire g722_p;
  wire g722_n;
  wire g723_p;
  wire g723_n;
  wire g724_p;
  wire g724_n;
  wire g725_p;
  wire g725_n;
  wire g726_p;
  wire g726_n;
  wire g727_p;
  wire g727_n;
  wire g728_p;
  wire g728_n;
  wire g729_p;
  wire g729_n;
  wire g730_p;
  wire g730_n;
  wire g731_p;
  wire g731_n;
  wire g732_p;
  wire g732_n;
  wire g733_p;
  wire g733_n;
  wire g734_p;
  wire g734_n;
  wire g735_p;
  wire g735_n;
  wire g736_p;
  wire g736_n;
  wire g737_p;
  wire g737_n;
  wire g738_p;
  wire g738_n;
  wire g739_p;
  wire g739_n;
  wire g740_p;
  wire g740_n;
  wire g741_p;
  wire g741_n;
  wire g742_p;
  wire g742_n;
  wire g743_p;
  wire g743_n;
  wire g744_p;
  wire g744_n;
  wire g745_p;
  wire g745_n;
  wire g746_p;
  wire g746_n;
  wire g747_p;
  wire g747_n;
  wire g748_p;
  wire g748_n;
  wire g749_p;
  wire g749_n;
  wire g750_p;
  wire g750_n;
  wire g751_p;
  wire g751_n;
  wire g752_p;
  wire g752_n;
  wire g753_p;
  wire g753_n;
  wire g754_p;
  wire g754_n;
  wire g755_p;
  wire g755_n;
  wire g756_p;
  wire g756_n;
  wire g757_p;
  wire g757_n;
  wire g758_p;
  wire g758_n;
  wire g759_p;
  wire g759_n;
  wire g760_p;
  wire g760_n;
  wire g761_p;
  wire g761_n;
  wire g762_p;
  wire g762_n;
  wire g763_p;
  wire g763_n;
  wire g764_p;
  wire g764_n;
  wire g765_p;
  wire g765_n;
  wire g766_p;
  wire g766_n;
  wire g767_p;
  wire g767_n;
  wire g768_p;
  wire g768_n;
  wire g769_p;
  wire g769_n;
  wire g770_p;
  wire g770_n;
  wire g771_p;
  wire g771_n;
  wire g772_p;
  wire g772_n;
  wire g773_p;
  wire g773_n;
  wire g774_p;
  wire g774_n;
  wire g775_p;
  wire g775_n;
  wire g776_p;
  wire g776_n;
  wire g777_p;
  wire g777_n;
  wire g778_p;
  wire g778_n;
  wire g779_p;
  wire g779_n;
  wire g780_p;
  wire g780_n;
  wire g781_p;
  wire g781_n;
  wire g782_p;
  wire g782_n;
  wire g783_p;
  wire g783_n;
  wire g784_p;
  wire g784_n;
  wire g785_p;
  wire g785_n;
  wire g786_p;
  wire g786_n;
  wire g787_p;
  wire g787_n;
  wire g788_p;
  wire g788_n;
  wire g789_p;
  wire g789_n;
  wire g790_p;
  wire g790_n;
  wire g791_p;
  wire g791_n;
  wire g792_p;
  wire g792_n;
  wire g793_p;
  wire g793_n;
  wire g794_p;
  wire g794_n;
  wire g795_p;
  wire g795_n;
  wire g796_p;
  wire g796_n;
  wire g797_p;
  wire g797_n;
  wire g798_p;
  wire g798_n;
  wire g799_p;
  wire g799_n;
  wire g800_p;
  wire g800_n;
  wire g801_p;
  wire g801_n;
  wire g802_p;
  wire g802_n;
  wire g803_p;
  wire g803_n;
  wire g804_p;
  wire g804_n;
  wire g805_p;
  wire g805_n;
  wire g806_p;
  wire g806_n;
  wire g807_p;
  wire g807_n;
  wire g808_p;
  wire g808_n;
  wire g809_p;
  wire g809_n;
  wire g810_p;
  wire g810_n;
  wire g811_p;
  wire g811_n;
  wire g812_p;
  wire g812_n;
  wire g813_p;
  wire g813_n;
  wire g814_p;
  wire g814_n;
  wire g815_p;
  wire g815_n;
  wire g816_p;
  wire g816_n;
  wire g817_p;
  wire g817_n;
  wire g818_p;
  wire g818_n;
  wire g819_p;
  wire g819_n;
  wire g820_p;
  wire g820_n;
  wire g821_p;
  wire g821_n;
  wire g822_p;
  wire g822_n;
  wire g823_p;
  wire g823_n;
  wire g824_p;
  wire g824_n;
  wire g825_p;
  wire g825_n;
  wire g826_p;
  wire g826_n;
  wire g827_p;
  wire g827_n;
  wire g828_p;
  wire g828_n;
  wire g829_p;
  wire g829_n;
  wire g830_p;
  wire g830_n;
  wire g831_p;
  wire g831_n;
  wire g832_p;
  wire g832_n;
  wire g833_p;
  wire g833_n;
  wire g834_p;
  wire g834_n;
  wire g835_p;
  wire g835_n;
  wire g836_p;
  wire g836_n;
  wire g837_p;
  wire g837_n;
  wire g838_p;
  wire g838_n;
  wire g839_p;
  wire g839_n;
  wire g840_p;
  wire g840_n;
  wire g841_p;
  wire g841_n;
  wire g842_p;
  wire g842_n;
  wire g843_p;
  wire g843_n;
  wire g844_p;
  wire g844_n;
  wire g845_p;
  wire g845_n;
  wire g846_p;
  wire g846_n;
  wire g847_p;
  wire g847_n;
  wire g848_p;
  wire g848_n;
  wire g849_p;
  wire g849_n;
  wire g850_p;
  wire g850_n;
  wire g851_p;
  wire g851_n;
  wire g852_p;
  wire g852_n;
  wire g853_p;
  wire g853_n;
  wire g854_p;
  wire g854_n;
  wire g855_p;
  wire g855_n;
  wire g856_p;
  wire g856_n;
  wire g857_p;
  wire g857_n;
  wire g858_p;
  wire g858_n;
  wire g859_p;
  wire g859_n;
  wire g860_p;
  wire g860_n;
  wire g861_p;
  wire g861_n;
  wire g862_p;
  wire g862_n;
  wire g863_p;
  wire g863_n;
  wire g864_p;
  wire g864_n;
  wire g865_p;
  wire g865_n;
  wire g866_p;
  wire g866_n;
  wire g867_p;
  wire g867_n;
  wire g868_p;
  wire g868_n;
  wire g869_p;
  wire g869_n;
  wire g870_p;
  wire g870_n;
  wire g871_p;
  wire g871_n;
  wire g872_p;
  wire g872_n;
  wire g873_p;
  wire g873_n;
  wire g874_p;
  wire g874_n;
  wire g875_p;
  wire g875_n;
  wire g876_p;
  wire g876_n;
  wire g877_p;
  wire g877_n;
  wire g878_p;
  wire g878_n;
  wire g879_p;
  wire g879_n;
  wire g880_p;
  wire g880_n;
  wire g881_p;
  wire g881_n;
  wire g882_p;
  wire g882_n;
  wire g883_p;
  wire g883_n;
  wire g884_p;
  wire g884_n;
  wire g885_p;
  wire g885_n;
  wire g886_p;
  wire g886_n;
  wire g887_p;
  wire g887_n;
  wire g888_p;
  wire g888_n;
  wire g889_p;
  wire g889_n;
  wire g890_p;
  wire g890_n;
  wire g891_p;
  wire g891_n;
  wire g892_p;
  wire g892_n;
  wire g893_p;
  wire g893_n;
  wire g894_p;
  wire g894_n;
  wire g895_p;
  wire g895_n;
  wire g896_p;
  wire g896_n;
  wire g897_p;
  wire g897_n;
  wire g898_p;
  wire g898_n;
  wire g899_p;
  wire g899_n;
  wire g900_p;
  wire g900_n;
  wire g901_p;
  wire g901_n;
  wire g902_p;
  wire g902_n;
  wire g903_p;
  wire g903_n;
  wire g904_p;
  wire g904_n;
  wire g905_p;
  wire g905_n;
  wire g906_p;
  wire g906_n;
  wire g907_p;
  wire g907_n;
  wire g908_p;
  wire g908_n;
  wire g909_p;
  wire g909_n;
  wire g910_p;
  wire g910_n;
  wire g911_p;
  wire g911_n;
  wire g912_p;
  wire g912_n;
  wire g913_p;
  wire g913_n;
  wire g914_p;
  wire g914_n;
  wire g915_p;
  wire g915_n;
  wire g916_p;
  wire g916_n;
  wire g917_p;
  wire g917_n;
  wire g918_p;
  wire g918_n;
  wire g919_p;
  wire g919_n;
  wire g920_p;
  wire g920_n;
  wire g921_p;
  wire g921_n;
  wire g922_p;
  wire g922_n;
  wire g923_p;
  wire g923_n;
  wire g924_p;
  wire g924_n;
  wire g925_p;
  wire g925_n;
  wire g926_p;
  wire g926_n;
  wire g927_p;
  wire g927_n;
  wire g928_p;
  wire g928_n;
  wire g929_p;
  wire g929_n;
  wire g930_p;
  wire g930_n;
  wire g931_p;
  wire g931_n;
  wire g932_p;
  wire g932_n;
  wire g933_p;
  wire g933_n;
  wire g934_p;
  wire g934_n;
  wire g935_p;
  wire g935_n;
  wire g936_p;
  wire g936_n;
  wire g937_p;
  wire g937_n;
  wire g938_p;
  wire g938_n;
  wire g939_p;
  wire g939_n;
  wire g940_p;
  wire g940_n;
  wire g941_p;
  wire g941_n;
  wire g942_p;
  wire g942_n;
  wire g943_p;
  wire g943_n;
  wire g944_p;
  wire g944_n;
  wire g945_p;
  wire g945_n;
  wire g946_p;
  wire g946_n;
  wire g947_p;
  wire g947_n;
  wire g948_p;
  wire g948_n;
  wire g949_p;
  wire g949_n;
  wire g950_p;
  wire g950_n;
  wire g951_p;
  wire g951_n;
  wire g952_p;
  wire g952_n;
  wire g953_p;
  wire g953_n;
  wire g954_p;
  wire g954_n;
  wire g955_p;
  wire g955_n;
  wire g956_p;
  wire g956_n;
  wire g957_p;
  wire g957_n;
  wire g958_p;
  wire g958_n;
  wire g959_p;
  wire g959_n;
  wire g960_p;
  wire g960_n;
  wire g961_p;
  wire g961_n;
  wire g962_p;
  wire g962_n;
  wire g963_p;
  wire g963_n;
  wire g964_p;
  wire g964_n;
  wire g965_p;
  wire g965_n;
  wire g966_p;
  wire g966_n;
  wire g967_p;
  wire g967_n;
  wire g968_p;
  wire g968_n;
  wire g969_p;
  wire g969_n;
  wire g970_p;
  wire g970_n;
  wire g971_p;
  wire g971_n;
  wire g972_p;
  wire g972_n;
  wire g973_p;
  wire g973_n;
  wire g974_p;
  wire g974_n;
  wire g975_p;
  wire g975_n;
  wire g976_p;
  wire g976_n;
  wire g977_p;
  wire g977_n;
  wire g978_p;
  wire g978_n;
  wire g979_p;
  wire g979_n;
  wire g980_p;
  wire g980_n;
  wire g981_p;
  wire g981_n;
  wire g982_p;
  wire g982_n;
  wire g983_p;
  wire g983_n;
  wire g984_p;
  wire g984_n;
  wire g985_p;
  wire g985_n;
  wire g986_p;
  wire g986_n;
  wire g987_p;
  wire g987_n;
  wire g988_p;
  wire g988_n;
  wire g989_p;
  wire g989_n;
  wire g990_p;
  wire g990_n;
  wire g991_p;
  wire g991_n;
  wire g992_p;
  wire g992_n;
  wire g993_p;
  wire g993_n;
  wire g994_p;
  wire g994_n;
  wire g995_p;
  wire g995_n;
  wire g996_p;
  wire g996_n;
  wire g997_p;
  wire g997_n;
  wire g998_p;
  wire g998_n;
  wire g999_p;
  wire g999_n;
  wire g1000_p;
  wire g1000_n;
  wire g1001_p;
  wire g1001_n;
  wire g1002_p;
  wire g1002_n;
  wire g1003_p;
  wire g1003_n;
  wire g1004_p;
  wire g1004_n;
  wire g1005_p;
  wire g1005_n;
  wire g1006_p;
  wire g1006_n;
  wire g1007_p;
  wire g1007_n;
  wire g1008_p;
  wire g1008_n;
  wire g1009_p;
  wire g1009_n;
  wire g1010_p;
  wire g1010_n;
  wire g1011_p;
  wire g1011_n;
  wire g1012_p;
  wire g1012_n;
  wire g1013_p;
  wire g1013_n;
  wire g1014_p;
  wire g1014_n;
  wire g1015_p;
  wire g1015_n;
  wire g1016_p;
  wire g1016_n;
  wire g1017_p;
  wire g1017_n;
  wire g1018_p;
  wire g1018_n;
  wire g1019_p;
  wire g1019_n;
  wire g1020_p;
  wire g1020_n;
  wire g1021_p;
  wire g1021_n;
  wire g1022_p;
  wire g1022_n;
  wire g1023_p;
  wire g1023_n;
  wire g1024_p;
  wire g1024_n;
  wire g1025_p;
  wire g1025_n;
  wire g1026_p;
  wire g1026_n;
  wire g1027_p;
  wire g1027_n;
  wire g1028_p;
  wire g1028_n;
  wire g1029_p;
  wire g1029_n;
  wire g1030_p;
  wire g1030_n;
  wire g1031_p;
  wire g1031_n;
  wire g1032_p;
  wire g1032_n;
  wire g1033_p;
  wire g1033_n;
  wire g1034_p;
  wire g1034_n;
  wire g1035_p;
  wire g1035_n;
  wire g1036_p;
  wire g1036_n;
  wire g1037_p;
  wire g1037_n;
  wire g1038_p;
  wire g1038_n;
  wire g1039_p;
  wire g1039_n;
  wire g1040_p;
  wire g1040_n;
  wire g1041_p;
  wire g1041_n;
  wire g1042_p;
  wire g1042_n;
  wire g1043_p;
  wire g1043_n;
  wire g1044_p;
  wire g1044_n;
  wire g1045_p;
  wire g1045_n;
  wire g1046_p;
  wire g1046_n;
  wire g1047_p;
  wire g1047_n;
  wire g1048_p;
  wire g1048_n;
  wire g1049_p;
  wire g1049_n;
  wire g1050_p;
  wire g1050_n;
  wire g1051_p;
  wire g1051_n;
  wire g1052_p;
  wire g1052_n;
  wire g1053_p;
  wire g1053_n;
  wire g1054_p;
  wire g1054_n;
  wire g1055_p;
  wire g1055_n;
  wire g1056_p;
  wire g1056_n;
  wire g1057_p;
  wire g1057_n;
  wire g1058_p;
  wire g1058_n;
  wire g1059_p;
  wire g1059_n;
  wire g1060_p;
  wire g1060_n;
  wire g1061_p;
  wire g1061_n;
  wire g1062_p;
  wire g1062_n;
  wire g1063_p;
  wire g1063_n;
  wire g1064_p;
  wire g1064_n;
  wire g1065_p;
  wire g1065_n;
  wire g1066_p;
  wire g1066_n;
  wire g1067_p;
  wire g1067_n;
  wire g1068_p;
  wire g1068_n;
  wire g1069_p;
  wire g1069_n;
  wire g1070_p;
  wire g1070_n;
  wire g1071_p;
  wire g1071_n;
  wire g1072_p;
  wire g1072_n;
  wire g1073_p;
  wire g1073_n;
  wire g1074_p;
  wire g1074_n;
  wire g1075_p;
  wire g1075_n;
  wire g1076_p;
  wire g1076_n;
  wire g1077_p;
  wire g1077_n;
  wire g1078_p;
  wire g1078_n;
  wire g1079_p;
  wire g1079_n;
  wire g1080_p;
  wire g1080_n;
  wire g1081_p;
  wire g1081_n;
  wire g1082_p;
  wire g1082_n;
  wire g1083_p;
  wire g1083_n;
  wire g1084_p;
  wire g1084_n;
  wire g1085_p;
  wire g1085_n;
  wire g1086_p;
  wire g1086_n;
  wire g1087_p;
  wire g1087_n;
  wire g1088_p;
  wire g1088_n;
  wire g1089_p;
  wire g1089_n;
  wire g1090_p;
  wire g1090_n;
  wire g1091_p;
  wire g1091_n;
  wire g1092_p;
  wire g1092_n;
  wire g1093_p;
  wire g1093_n;
  wire g1094_p;
  wire g1094_n;
  wire g1095_p;
  wire g1095_n;
  wire g1096_p;
  wire g1096_n;
  wire g1097_p;
  wire g1097_n;
  wire g1098_p;
  wire g1098_n;
  wire g1099_p;
  wire g1099_n;
  wire g1100_p;
  wire g1100_n;
  wire g1101_p;
  wire g1101_n;
  wire g1102_p;
  wire g1102_n;
  wire g1103_p;
  wire g1103_n;
  wire g1104_p;
  wire g1104_n;
  wire g1105_p;
  wire g1105_n;
  wire g1106_p;
  wire g1106_n;
  wire g1107_p;
  wire g1107_n;
  wire g1108_p;
  wire g1108_n;
  wire g1109_p;
  wire g1109_n;
  wire g1110_p;
  wire g1110_n;
  wire g1111_p;
  wire g1111_n;
  wire g1112_p;
  wire g1112_n;
  wire g1113_p;
  wire g1113_n;
  wire g1114_p;
  wire g1114_n;
  wire g1115_p;
  wire g1115_n;
  wire g1116_p;
  wire g1116_n;
  wire g1117_p;
  wire g1117_n;
  wire g1118_p;
  wire g1118_n;
  wire g1119_p;
  wire g1119_n;
  wire g1120_p;
  wire g1120_n;
  wire g1121_p;
  wire g1121_n;
  wire g1122_p;
  wire g1122_n;
  wire g1123_p;
  wire g1123_n;
  wire g1124_p;
  wire g1124_n;
  wire g1125_p;
  wire g1125_n;
  wire g1126_p;
  wire g1126_n;
  wire g1127_p;
  wire g1127_n;
  wire g1128_p;
  wire g1128_n;
  wire g1129_p;
  wire g1129_n;
  wire g1130_p;
  wire g1130_n;
  wire g1131_p;
  wire g1131_n;
  wire g1132_p;
  wire g1132_n;
  wire g1133_p;
  wire g1133_n;
  wire g1134_p;
  wire g1134_n;
  wire g1135_p;
  wire g1135_n;
  wire g1136_p;
  wire g1136_n;
  wire g1137_p;
  wire g1137_n;
  wire g1138_p;
  wire g1138_n;
  wire g1139_p;
  wire g1139_n;
  wire g1140_p;
  wire g1140_n;
  wire g1141_p;
  wire g1141_n;
  wire g1142_p;
  wire g1142_n;
  wire g1143_p;
  wire g1143_n;
  wire g1144_p;
  wire g1144_n;
  wire g1145_p;
  wire g1145_n;
  wire g1146_p;
  wire g1146_n;
  wire g1147_p;
  wire g1147_n;
  wire g1148_p;
  wire g1148_n;
  wire g1149_p;
  wire g1149_n;
  wire g1150_p;
  wire g1150_n;
  wire g1151_p;
  wire g1151_n;
  wire g1152_p;
  wire g1152_n;
  wire g1153_p;
  wire g1153_n;
  wire g1154_p;
  wire g1154_n;
  wire g1155_p;
  wire g1155_n;
  wire g1156_p;
  wire g1156_n;
  wire g1157_p;
  wire g1157_n;
  wire g1158_p;
  wire g1158_n;
  wire g1159_p;
  wire g1159_n;
  wire g1160_p;
  wire g1160_n;
  wire g1161_p;
  wire g1161_n;
  wire g1162_p;
  wire g1162_n;
  wire g1163_p;
  wire g1163_n;
  wire g1164_p;
  wire g1164_n;
  wire g1165_p;
  wire g1165_n;
  wire g1166_p;
  wire g1166_n;
  wire g1167_p;
  wire g1167_n;
  wire g1168_p;
  wire g1168_n;
  wire g1169_p;
  wire g1169_n;
  wire g1170_p;
  wire g1170_n;
  wire g1171_p;
  wire g1171_n;
  wire g1172_p;
  wire g1172_n;
  wire g1173_p;
  wire g1173_n;
  wire g1174_p;
  wire g1174_n;
  wire g1175_p;
  wire g1175_n;
  wire g1176_p;
  wire g1176_n;
  wire g1177_p;
  wire g1177_n;
  wire g1178_p;
  wire g1178_n;
  wire g1179_p;
  wire g1179_n;
  wire g1180_p;
  wire g1180_n;
  wire g1181_p;
  wire g1181_n;
  wire g1182_p;
  wire g1182_n;
  wire g1183_p;
  wire g1183_n;
  wire g1184_p;
  wire g1184_n;
  wire g1185_p;
  wire g1185_n;
  wire g1186_p;
  wire g1186_n;
  wire g1187_p;
  wire g1187_n;
  wire g1188_p;
  wire g1188_n;
  wire g1189_p;
  wire g1189_n;
  wire g1190_p;
  wire g1190_n;
  wire g1191_p;
  wire g1191_n;
  wire g1192_p;
  wire g1192_n;
  wire g1193_p;
  wire g1193_n;
  wire g1194_p;
  wire g1194_n;
  wire g1195_p;
  wire g1195_n;
  wire g1196_p;
  wire g1196_n;
  wire g1197_p;
  wire g1197_n;
  wire g1198_p;
  wire g1198_n;
  wire g1199_p;
  wire g1199_n;
  wire g1200_p;
  wire g1200_n;
  wire g1201_p;
  wire g1201_n;
  wire g1202_p;
  wire g1202_n;
  wire g1203_p;
  wire g1203_n;
  wire g1204_p;
  wire g1204_n;
  wire g1205_p;
  wire g1205_n;
  wire g1206_p;
  wire g1206_n;
  wire g1207_p;
  wire g1207_n;
  wire g1208_p;
  wire g1208_n;
  wire g1209_p;
  wire g1209_n;
  wire g1210_p;
  wire g1210_n;
  wire g1211_p;
  wire g1211_n;
  wire g1212_p;
  wire g1212_n;
  wire g1213_p;
  wire g1213_n;
  wire g1214_p;
  wire g1214_n;
  wire g1215_p;
  wire g1215_n;
  wire g1216_p;
  wire g1216_n;
  wire g1217_p;
  wire g1217_n;
  wire g1218_p;
  wire g1218_n;
  wire g1219_p;
  wire g1219_n;
  wire g1220_p;
  wire g1220_n;
  wire g1221_p;
  wire g1221_n;
  wire g1222_p;
  wire g1222_n;
  wire g1223_p;
  wire g1223_n;
  wire g1224_p;
  wire g1224_n;
  wire g1225_p;
  wire g1225_n;
  wire g1226_p;
  wire g1226_n;
  wire g1227_p;
  wire g1227_n;
  wire g1228_p;
  wire g1228_n;
  wire g1229_p;
  wire g1229_n;
  wire g1230_p;
  wire g1230_n;
  wire g1231_p;
  wire g1231_n;
  wire g1232_p;
  wire g1232_n;
  wire g1233_p;
  wire g1233_n;
  wire g1234_p;
  wire g1234_n;
  wire g1235_p;
  wire g1235_n;
  wire g1236_p;
  wire g1236_n;
  wire g1237_p;
  wire g1237_n;
  wire g1238_p;
  wire g1238_n;
  wire g1239_p;
  wire g1239_n;
  wire g1240_p;
  wire g1240_n;
  wire g1241_p;
  wire g1241_n;
  wire g1242_p;
  wire g1242_n;
  wire g1243_p;
  wire g1243_n;
  wire g1244_p;
  wire g1244_n;
  wire g1245_p;
  wire g1245_n;
  wire g1246_p;
  wire g1246_n;
  wire g1247_p;
  wire g1247_n;
  wire g1248_p;
  wire g1248_n;
  wire g1249_p;
  wire g1249_n;
  wire g1250_p;
  wire g1250_n;
  wire g1251_p;
  wire g1251_n;
  wire g1252_p;
  wire g1252_n;
  wire g1253_p;
  wire g1253_n;
  wire g1254_p;
  wire g1254_n;
  wire g1255_p;
  wire g1255_n;
  wire g1256_p;
  wire g1256_n;
  wire g1257_p;
  wire g1257_n;
  wire g1258_p;
  wire g1258_n;
  wire g1259_p;
  wire g1259_n;
  wire g1260_p;
  wire g1260_n;
  wire g1261_p;
  wire g1261_n;
  wire g1262_p;
  wire g1262_n;
  wire g1263_p;
  wire g1263_n;
  wire g1264_p;
  wire g1264_n;
  wire g1265_p;
  wire g1265_n;
  wire g1266_p;
  wire g1266_n;
  wire g1267_p;
  wire g1267_n;
  wire g1268_p;
  wire g1268_n;
  wire g1269_p;
  wire g1269_n;
  wire g1270_p;
  wire g1270_n;
  wire g1271_p;
  wire g1271_n;
  wire g1272_p;
  wire g1272_n;
  wire g1273_p;
  wire g1273_n;
  wire g1274_p;
  wire g1274_n;
  wire g1275_p;
  wire g1275_n;
  wire g1276_p;
  wire g1276_n;
  wire g1277_p;
  wire g1277_n;
  wire g1278_p;
  wire g1278_n;
  wire g1279_p;
  wire g1279_n;
  wire g1280_p;
  wire g1280_n;
  wire g1281_p;
  wire g1281_n;
  wire g1282_p;
  wire g1282_n;
  wire g1283_p;
  wire g1283_n;
  wire g1284_p;
  wire g1284_n;
  wire g1285_p;
  wire g1285_n;
  wire g1286_p;
  wire g1286_n;
  wire g1287_p;
  wire g1287_n;
  wire g1288_p;
  wire g1288_n;
  wire g1289_p;
  wire g1289_n;
  wire g1290_p;
  wire g1290_n;
  wire g1291_p;
  wire g1291_n;
  wire g1292_p;
  wire g1292_n;
  wire g1293_p;
  wire g1293_n;
  wire g1294_p;
  wire g1294_n;
  wire g1295_p;
  wire g1295_n;
  wire g1296_p;
  wire g1296_n;
  wire g1297_p;
  wire g1297_n;
  wire g1298_p;
  wire g1298_n;
  wire g1299_p;
  wire g1299_n;
  wire g1300_p;
  wire g1300_n;
  wire g1301_p;
  wire g1301_n;
  wire g1302_p;
  wire g1302_n;
  wire g1303_p;
  wire g1303_n;
  wire g1304_p;
  wire g1304_n;
  wire g1305_p;
  wire g1305_n;
  wire g1306_p;
  wire g1306_n;
  wire g1307_p;
  wire g1307_n;
  wire g1308_p;
  wire g1308_n;
  wire g1309_p;
  wire g1309_n;
  wire g1310_p;
  wire g1310_n;
  wire g1311_p;
  wire g1311_n;
  wire g1312_p;
  wire g1312_n;
  wire g1313_p;
  wire g1313_n;
  wire g1314_p;
  wire g1314_n;
  wire g1315_p;
  wire g1315_n;
  wire g1316_p;
  wire g1316_n;
  wire g1317_p;
  wire g1317_n;
  wire g1318_p;
  wire g1318_n;
  wire g1319_p;
  wire g1319_n;
  wire g1320_p;
  wire g1320_n;
  wire g1321_p;
  wire g1321_n;
  wire g1322_p;
  wire g1322_n;
  wire g1323_p;
  wire g1323_n;
  wire g1324_p;
  wire g1324_n;
  wire g1325_p;
  wire g1325_n;
  wire g1326_p;
  wire g1326_n;
  wire g1327_p;
  wire g1327_n;
  wire g1328_p;
  wire g1328_n;
  wire g1329_p;
  wire g1329_n;
  wire g1330_p;
  wire g1330_n;
  wire g1331_p;
  wire g1331_n;
  wire g1332_p;
  wire g1332_n;
  wire g1333_p;
  wire g1333_n;
  wire g1334_p;
  wire g1334_n;
  wire g1335_p;
  wire g1335_n;
  wire g1336_p;
  wire g1336_n;
  wire g1337_p;
  wire g1337_n;
  wire g1338_p;
  wire g1338_n;
  wire g1339_p;
  wire g1339_n;
  wire g1340_p;
  wire g1340_n;
  wire g1341_p;
  wire g1341_n;
  wire g1342_p;
  wire g1342_n;
  wire g1343_p;
  wire g1343_n;
  wire g1344_p;
  wire g1344_n;
  wire g1345_p;
  wire g1345_n;
  wire g1346_p;
  wire g1346_n;
  wire g1347_p;
  wire g1347_n;
  wire g1348_p;
  wire g1348_n;
  wire g1349_p;
  wire g1349_n;
  wire g1350_p;
  wire g1350_n;
  wire g1351_p;
  wire g1351_n;
  wire g1352_p;
  wire g1352_n;
  wire g1353_p;
  wire g1353_n;
  wire g1354_p;
  wire g1354_n;
  wire g1355_p;
  wire g1355_n;
  wire g1356_p;
  wire g1356_n;
  wire g1357_p;
  wire g1357_n;
  wire g1358_p;
  wire g1358_n;
  wire g1359_p;
  wire g1359_n;
  wire g1360_p;
  wire g1360_n;
  wire g1361_p;
  wire g1361_n;
  wire g1362_p;
  wire g1362_n;
  wire g1363_p;
  wire g1363_n;
  wire g1364_p;
  wire g1364_n;
  wire g1365_p;
  wire g1365_n;
  wire g1366_p;
  wire g1366_n;
  wire g1367_p;
  wire g1367_n;
  wire g1368_p;
  wire g1368_n;
  wire g1369_p;
  wire g1369_n;
  wire g1370_p;
  wire g1370_n;
  wire g1371_p;
  wire g1371_n;
  wire g1372_p;
  wire g1372_n;
  wire g1373_p;
  wire g1373_n;
  wire g1374_p;
  wire g1374_n;
  wire g1375_p;
  wire g1375_n;
  wire g1376_p;
  wire g1376_n;
  wire g1377_p;
  wire g1377_n;
  wire g1378_p;
  wire g1378_n;
  wire g1379_p;
  wire g1379_n;
  wire g1380_p;
  wire g1380_n;
  wire g1381_p;
  wire g1381_n;
  wire g1382_p;
  wire g1382_n;
  wire g1383_p;
  wire g1383_n;
  wire g1384_p;
  wire g1384_n;
  wire g1385_p;
  wire g1385_n;
  wire g1386_p;
  wire g1386_n;
  wire g1387_p;
  wire g1387_n;
  wire g1388_p;
  wire g1388_n;
  wire g1389_p;
  wire g1389_n;
  wire g1390_p;
  wire g1390_n;
  wire g1391_p;
  wire g1391_n;
  wire g1392_p;
  wire g1392_n;
  wire g1393_p;
  wire g1393_n;
  wire g1394_p;
  wire g1394_n;
  wire g1395_p;
  wire g1395_n;
  wire g1396_p;
  wire g1396_n;
  wire g1397_p;
  wire g1397_n;
  wire g1398_p;
  wire g1398_n;
  wire g1399_p;
  wire g1399_n;
  wire g1400_p;
  wire g1400_n;
  wire g1401_p;
  wire g1401_n;
  wire g1402_p;
  wire g1402_n;
  wire g1403_p;
  wire g1403_n;
  wire g1404_p;
  wire g1404_n;
  wire g1405_p;
  wire g1405_n;
  wire g1406_p;
  wire g1406_n;
  wire g1407_p;
  wire g1407_n;
  wire g1408_p;
  wire g1408_n;
  wire g1409_p;
  wire g1409_n;
  wire g1410_p;
  wire g1410_n;
  wire g1411_p;
  wire g1411_n;
  wire g1412_p;
  wire g1412_n;
  wire g1413_p;
  wire g1413_n;
  wire g1414_p;
  wire g1414_n;
  wire g1415_p;
  wire g1415_n;
  wire g1416_p;
  wire g1416_n;
  wire g1417_p;
  wire g1417_n;
  wire g1418_p;
  wire g1418_n;
  wire g1419_p;
  wire g1419_n;
  wire g1420_p;
  wire g1420_n;
  wire g1421_p;
  wire g1421_n;
  wire g1422_p;
  wire g1422_n;
  wire g1423_p;
  wire g1423_n;
  wire g1424_p;
  wire g1424_n;
  wire g1425_p;
  wire g1425_n;
  wire g1426_p;
  wire g1426_n;
  wire g1427_p;
  wire g1427_n;
  wire g1428_p;
  wire g1428_n;
  wire g1429_p;
  wire g1429_n;
  wire g1430_p;
  wire g1430_n;
  wire g1431_p;
  wire g1431_n;
  wire g1432_p;
  wire g1432_n;
  wire g1433_p;
  wire g1433_n;
  wire g1434_p;
  wire g1434_n;
  wire g1435_p;
  wire g1435_n;
  wire g1436_p;
  wire g1436_n;
  wire g1437_p;
  wire g1437_n;
  wire g1438_p;
  wire g1438_n;
  wire g1439_p;
  wire g1439_n;
  wire g1440_p;
  wire g1440_n;
  wire g1441_p;
  wire g1441_n;
  wire g1442_p;
  wire g1442_n;
  wire g1443_p;
  wire g1443_n;
  wire g1444_p;
  wire g1444_n;
  wire g1445_p;
  wire g1445_n;
  wire g1446_p;
  wire g1446_n;
  wire g1447_p;
  wire g1447_n;
  wire g1448_p;
  wire g1448_n;
  wire g1449_p;
  wire g1449_n;
  wire g1450_p;
  wire g1450_n;
  wire g1451_p;
  wire g1451_n;
  wire g1452_p;
  wire g1452_n;
  wire g1453_p;
  wire g1453_n;
  wire g1454_p;
  wire g1454_n;
  wire g1455_p;
  wire g1455_n;
  wire g1456_p;
  wire g1456_n;
  wire g1457_p;
  wire g1457_n;
  wire g1458_p;
  wire g1458_n;
  wire g1459_p;
  wire g1459_n;
  wire g1460_p;
  wire g1460_n;
  wire g1461_p;
  wire g1461_n;
  wire g1462_p;
  wire g1462_n;
  wire g1463_p;
  wire g1463_n;
  wire g1464_p;
  wire g1464_n;
  wire g1465_p;
  wire g1465_n;
  wire g1466_p;
  wire g1466_n;
  wire g1467_p;
  wire g1467_n;
  wire g1468_p;
  wire g1468_n;
  wire g1469_p;
  wire g1469_n;
  wire g1470_p;
  wire g1470_n;
  wire g1471_p;
  wire g1471_n;
  wire g1472_p;
  wire g1472_n;
  wire g1473_p;
  wire g1473_n;
  wire g1474_p;
  wire g1474_n;
  wire g1475_p;
  wire g1475_n;
  wire g1476_p;
  wire g1476_n;
  wire g1477_p;
  wire g1477_n;
  wire g1478_p;
  wire g1478_n;
  wire g1479_p;
  wire g1479_n;
  wire g1480_p;
  wire g1480_n;
  wire g1481_p;
  wire g1481_n;
  wire g1482_p;
  wire g1482_n;
  wire g1483_p;
  wire g1483_n;
  wire g1484_p;
  wire g1484_n;
  wire g1485_p;
  wire g1485_n;
  wire g1486_p;
  wire g1486_n;
  wire g1487_p;
  wire g1487_n;
  wire g1488_p;
  wire g1488_n;
  wire g1489_p;
  wire g1489_n;
  wire g1490_p;
  wire g1490_n;
  wire g1491_p;
  wire g1491_n;
  wire g1492_p;
  wire g1492_n;
  wire g1493_p;
  wire g1493_n;
  wire g1494_p;
  wire g1494_n;
  wire g1495_p;
  wire g1495_n;
  wire g1496_p;
  wire g1496_n;
  wire g1497_p;
  wire g1497_n;
  wire g1498_p;
  wire g1498_n;
  wire g1499_p;
  wire g1499_n;
  wire g1500_p;
  wire g1500_n;
  wire g1501_p;
  wire g1501_n;
  wire g1502_p;
  wire g1502_n;
  wire g1503_p;
  wire g1503_n;
  wire g1504_p;
  wire g1504_n;
  wire g1505_p;
  wire g1505_n;
  wire g1506_p;
  wire g1506_n;
  wire g1507_p;
  wire g1507_n;
  wire g1508_p;
  wire g1508_n;
  wire g1509_p;
  wire g1509_n;
  wire g1510_p;
  wire g1510_n;
  wire g1511_p;
  wire g1511_n;
  wire g1512_p;
  wire g1512_n;
  wire g1513_p;
  wire g1513_n;
  wire g1514_p;
  wire g1514_n;
  wire g1515_p;
  wire g1515_n;
  wire g1516_p;
  wire g1516_n;
  wire g1517_p;
  wire g1517_n;
  wire g1518_p;
  wire g1518_n;
  wire g1519_p;
  wire g1519_n;
  wire g1520_p;
  wire g1520_n;
  wire g1521_p;
  wire g1521_n;
  wire g1522_p;
  wire g1522_n;
  wire g1523_p;
  wire g1523_n;
  wire g1524_p;
  wire g1524_n;
  wire g1525_p;
  wire g1525_n;
  wire g1526_p;
  wire g1526_n;
  wire g1527_p;
  wire g1527_n;
  wire g1528_p;
  wire g1528_n;
  wire g1529_p;
  wire g1529_n;
  wire g1530_p;
  wire g1530_n;
  wire g1531_p;
  wire g1531_n;
  wire g1532_p;
  wire g1532_n;
  wire g1533_p;
  wire g1533_n;
  wire g1534_p;
  wire g1534_n;
  wire g1535_p;
  wire g1535_n;
  wire g1536_p;
  wire g1536_n;
  wire g1537_p;
  wire g1537_n;
  wire g1538_p;
  wire g1538_n;
  wire g1539_p;
  wire g1539_n;
  wire g1540_p;
  wire g1540_n;
  wire g1541_p;
  wire g1541_n;
  wire g1542_p;
  wire g1542_n;
  wire g1543_p;
  wire g1543_n;
  wire g1544_p;
  wire g1544_n;
  wire g1545_p;
  wire g1545_n;
  wire g1546_p;
  wire g1546_n;
  wire g1547_p;
  wire g1547_n;
  wire g1548_p;
  wire g1548_n;
  wire g1549_p;
  wire g1549_n;
  wire g1550_p;
  wire g1550_n;
  wire g1551_p;
  wire g1551_n;
  wire g1552_p;
  wire g1552_n;
  wire g1553_p;
  wire g1553_n;
  wire g1554_p;
  wire g1554_n;
  wire g1555_p;
  wire g1555_n;
  wire g1556_p;
  wire g1556_n;
  wire g1557_p;
  wire g1557_n;
  wire g1558_p;
  wire g1558_n;
  wire g1559_p;
  wire g1559_n;
  wire g1560_p;
  wire g1560_n;
  wire g1561_p;
  wire g1561_n;
  wire g1562_p;
  wire g1562_n;
  wire g1563_p;
  wire g1563_n;
  wire g1564_p;
  wire g1564_n;
  wire g1565_p;
  wire g1565_n;
  wire g1566_p;
  wire g1566_n;
  wire g1567_p;
  wire g1567_n;
  wire g1568_p;
  wire g1568_n;
  wire g1569_p;
  wire g1569_n;
  wire g1570_p;
  wire g1570_n;
  wire g1571_p;
  wire g1571_n;
  wire g1572_p;
  wire g1572_n;
  wire g1573_p;
  wire g1573_n;
  wire g1574_p;
  wire g1574_n;
  wire g1575_p;
  wire g1575_n;
  wire g1576_p;
  wire g1576_n;
  wire g1577_p;
  wire g1577_n;
  wire g1578_p;
  wire g1578_n;
  wire g1579_p;
  wire g1579_n;
  wire g1580_p;
  wire g1580_n;
  wire g1581_p;
  wire g1581_n;
  wire g1582_p;
  wire g1582_n;
  wire g1583_p;
  wire g1583_n;
  wire g1584_p;
  wire g1584_n;
  wire g1585_p;
  wire g1585_n;
  wire g1586_p;
  wire g1586_n;
  wire g1587_p;
  wire g1587_n;
  wire g1588_p;
  wire g1588_n;
  wire g1589_p;
  wire g1589_n;
  wire g1590_p;
  wire g1590_n;
  wire g1591_p;
  wire g1591_n;
  wire g1592_p;
  wire g1592_n;
  wire g1593_p;
  wire g1593_n;
  wire g1594_p;
  wire g1594_n;
  wire g1595_p;
  wire g1595_n;
  wire g1596_p;
  wire g1596_n;
  wire g1597_p;
  wire g1597_n;
  wire g1598_p;
  wire g1598_n;
  wire g1599_p;
  wire g1599_n;
  wire g1600_p;
  wire g1600_n;
  wire g1601_p;
  wire g1601_n;
  wire g1602_p;
  wire g1602_n;
  wire g1603_p;
  wire g1603_n;
  wire g1604_p;
  wire g1604_n;
  wire g1605_p;
  wire g1605_n;
  wire g1606_p;
  wire g1606_n;
  wire g1607_p;
  wire g1607_n;
  wire g1608_p;
  wire g1608_n;
  wire g1609_p;
  wire g1609_n;
  wire g1610_p;
  wire g1610_n;
  wire g1611_p;
  wire g1611_n;
  wire g1612_p;
  wire g1612_n;
  wire g1613_p;
  wire g1613_n;
  wire g1614_p;
  wire g1614_n;
  wire g1615_p;
  wire g1615_n;
  wire g1616_p;
  wire g1616_n;
  wire g1617_p;
  wire g1617_n;
  wire g1618_p;
  wire g1618_n;
  wire g1619_p;
  wire g1619_n;
  wire g1620_p;
  wire g1620_n;
  wire g1621_p;
  wire g1621_n;
  wire g1622_p;
  wire g1622_n;
  wire g1623_p;
  wire g1623_n;
  wire g1624_p;
  wire g1624_n;
  wire g1625_p;
  wire g1625_n;
  wire g1626_p;
  wire g1626_n;
  wire g1627_p;
  wire g1627_n;
  wire g1628_p;
  wire g1628_n;
  wire g1629_p;
  wire g1629_n;
  wire g1630_p;
  wire g1630_n;
  wire g1631_p;
  wire g1631_n;
  wire g1632_p;
  wire g1632_n;
  wire g1633_p;
  wire g1633_n;
  wire g1634_p;
  wire g1634_n;
  wire g1635_p;
  wire g1635_n;
  wire g1636_p;
  wire g1636_n;
  wire g1637_p;
  wire g1637_n;
  wire g1638_p;
  wire g1638_n;
  wire g1639_p;
  wire g1639_n;
  wire g1640_p;
  wire g1640_n;
  wire g1641_p;
  wire g1641_n;
  wire g1642_p;
  wire g1642_n;
  wire g1643_p;
  wire g1643_n;
  wire g1644_p;
  wire g1644_n;
  wire g1645_p;
  wire g1645_n;
  wire g1646_p;
  wire g1646_n;
  wire g1647_p;
  wire g1647_n;
  wire g1648_p;
  wire g1648_n;
  wire g1649_p;
  wire g1649_n;
  wire g1650_p;
  wire g1650_n;
  wire g1651_p;
  wire g1651_n;
  wire g1652_p;
  wire g1652_n;
  wire g1653_p;
  wire g1653_n;
  wire g1654_p;
  wire g1654_n;
  wire g1655_p;
  wire g1655_n;
  wire g1656_p;
  wire g1656_n;
  wire g1657_p;
  wire g1657_n;
  wire g1658_p;
  wire g1658_n;
  wire g1659_p;
  wire g1659_n;
  wire g1660_p;
  wire g1660_n;
  wire g1661_p;
  wire g1661_n;
  wire g1662_p;
  wire g1662_n;
  wire g1663_p;
  wire g1663_n;
  wire g1664_p;
  wire g1664_n;
  wire g1665_p;
  wire g1665_n;
  wire g1666_p;
  wire g1666_n;
  wire g1667_p;
  wire g1667_n;
  wire g1668_p;
  wire g1668_n;
  wire g1669_p;
  wire g1669_n;
  wire g1670_p;
  wire g1670_n;
  wire g1671_p;
  wire g1671_n;
  wire g1672_p;
  wire g1672_n;
  wire g1673_p;
  wire g1673_n;
  wire g1674_p;
  wire g1674_n;
  wire g1675_p;
  wire g1675_n;
  wire g1676_p;
  wire g1676_n;
  wire g1677_p;
  wire g1677_n;
  wire g1678_p;
  wire g1678_n;
  wire g1679_p;
  wire g1679_n;
  wire g1680_p;
  wire g1680_n;
  wire g1681_p;
  wire g1681_n;
  wire g1682_p;
  wire g1682_n;
  wire g1683_p;
  wire g1683_n;
  wire g1684_p;
  wire g1684_n;
  wire g1685_p;
  wire g1685_n;
  wire g1686_p;
  wire g1686_n;
  wire g1687_p;
  wire g1687_n;
  wire g1688_p;
  wire g1688_n;
  wire g1689_p;
  wire g1689_n;
  wire g1690_p;
  wire g1690_n;
  wire g1691_p;
  wire g1691_n;
  wire g1692_p;
  wire g1692_n;
  wire g1693_p;
  wire g1693_n;
  wire g1694_p;
  wire g1694_n;
  wire g1695_p;
  wire g1695_n;
  wire g1696_p;
  wire g1696_n;
  wire g1697_p;
  wire g1697_n;
  wire g1698_p;
  wire g1698_n;
  wire g1699_p;
  wire g1699_n;
  wire g1700_p;
  wire g1700_n;
  wire g1701_p;
  wire g1701_n;
  wire g1702_p;
  wire g1702_n;
  wire g1703_p;
  wire g1703_n;
  wire g1704_p;
  wire g1704_n;
  wire g1705_p;
  wire g1705_n;
  wire g1706_p;
  wire g1706_n;
  wire g1707_p;
  wire g1707_n;
  wire g1708_p;
  wire g1708_n;
  wire g1709_p;
  wire g1709_n;
  wire g1710_p;
  wire g1710_n;
  wire g1711_p;
  wire g1711_n;
  wire g1712_p;
  wire g1712_n;
  wire g1713_p;
  wire g1713_n;
  wire g1714_p;
  wire g1714_n;
  wire g1715_p;
  wire g1715_n;
  wire g1716_p;
  wire g1716_n;
  wire g1717_p;
  wire g1717_n;
  wire g1718_p;
  wire g1718_n;
  wire g1719_p;
  wire g1719_n;
  wire g1720_p;
  wire g1720_n;
  wire g1721_p;
  wire g1721_n;
  wire g1722_p;
  wire g1722_n;
  wire g1723_p;
  wire g1723_n;
  wire g1724_p;
  wire g1724_n;
  wire g1725_p;
  wire g1725_n;
  wire g1726_p;
  wire g1726_n;
  wire g1727_p;
  wire g1727_n;
  wire g1728_p;
  wire g1728_n;
  wire g1729_p;
  wire g1729_n;
  wire g1730_p;
  wire g1730_n;
  wire g1731_p;
  wire g1731_n;
  wire g1732_p;
  wire g1732_n;
  wire g1733_p;
  wire g1733_n;
  wire g1734_p;
  wire g1734_n;
  wire g1735_p;
  wire g1735_n;
  wire g1736_p;
  wire g1736_n;
  wire g1737_p;
  wire g1737_n;
  wire g1738_p;
  wire g1738_n;
  wire g1739_p;
  wire g1739_n;
  wire g1740_p;
  wire g1740_n;
  wire g1741_p;
  wire g1741_n;
  wire g1742_p;
  wire g1742_n;
  wire g1743_p;
  wire g1743_n;
  wire g1744_p;
  wire g1744_n;
  wire g1745_p;
  wire g1745_n;
  wire g1746_p;
  wire g1746_n;
  wire g1747_p;
  wire g1747_n;
  wire g1748_p;
  wire g1748_n;
  wire g1749_p;
  wire g1749_n;
  wire g1750_p;
  wire g1750_n;
  wire g1751_p;
  wire g1751_n;
  wire g1752_p;
  wire g1752_n;
  wire g1753_p;
  wire g1753_n;
  wire g1754_p;
  wire g1754_n;
  wire g1755_p;
  wire g1755_n;
  wire g1756_p;
  wire g1756_n;
  wire g1757_p;
  wire g1757_n;
  wire g1758_p;
  wire g1758_n;
  wire g1759_p;
  wire g1759_n;
  wire g1760_p;
  wire g1760_n;
  wire g1761_p;
  wire g1761_n;
  wire g1762_p;
  wire g1762_n;
  wire g1763_p;
  wire g1763_n;
  wire g1764_p;
  wire g1764_n;
  wire g1765_p;
  wire g1765_n;
  wire g1766_p;
  wire g1766_n;
  wire g1767_p;
  wire g1767_n;
  wire g1768_p;
  wire g1768_n;
  wire g1769_p;
  wire g1769_n;
  wire g1770_p;
  wire g1770_n;
  wire g1771_p;
  wire g1771_n;
  wire g1772_p;
  wire g1772_n;
  wire g1773_p;
  wire g1773_n;
  wire g1774_p;
  wire g1774_n;
  wire g1775_p;
  wire g1775_n;
  wire g1776_p;
  wire g1776_n;
  wire g1777_p;
  wire g1777_n;
  wire g1778_p;
  wire g1778_n;
  wire g1779_p;
  wire g1779_n;
  wire g1780_p;
  wire g1780_n;
  wire g1781_p;
  wire g1781_n;
  wire g1782_p;
  wire g1782_n;
  wire g1783_p;
  wire g1783_n;
  wire g1784_p;
  wire g1784_n;
  wire g1785_p;
  wire g1785_n;
  wire g1786_p;
  wire g1786_n;
  wire g1787_p;
  wire g1787_n;
  wire g1788_p;
  wire g1788_n;
  wire g1789_p;
  wire g1789_n;
  wire g1790_p;
  wire g1790_n;
  wire g1791_p;
  wire g1791_n;
  wire g1792_p;
  wire g1792_n;
  wire g1793_p;
  wire g1793_n;
  wire g1794_p;
  wire g1794_n;
  wire g1795_p;
  wire g1795_n;
  wire g1796_p;
  wire g1796_n;
  wire g1797_p;
  wire g1797_n;
  wire g1798_p;
  wire g1798_n;
  wire g1799_p;
  wire g1799_n;
  wire g1800_p;
  wire g1800_n;
  wire g1801_p;
  wire g1801_n;
  wire g1802_p;
  wire g1802_n;
  wire g1803_p;
  wire g1803_n;
  wire g1804_p;
  wire g1804_n;
  wire g1805_p;
  wire g1805_n;
  wire g1806_p;
  wire g1806_n;
  wire g1807_p;
  wire g1807_n;
  wire g1808_p;
  wire g1808_n;
  wire g1809_p;
  wire g1809_n;
  wire g1810_p;
  wire g1810_n;
  wire g1811_p;
  wire g1811_n;
  wire g1812_p;
  wire g1812_n;
  wire g1813_p;
  wire g1813_n;
  wire g1814_p;
  wire g1814_n;
  wire g1815_p;
  wire g1815_n;
  wire g1816_p;
  wire g1816_n;
  wire g1817_p;
  wire g1817_n;
  wire g1818_p;
  wire g1818_n;
  wire g1819_p;
  wire g1819_n;
  wire g1820_p;
  wire g1820_n;
  wire g1821_p;
  wire g1821_n;
  wire g1822_p;
  wire g1822_n;
  wire g1823_p;
  wire g1823_n;
  wire g1824_p;
  wire g1824_n;
  wire g1825_p;
  wire g1825_n;
  wire g1826_p;
  wire g1826_n;
  wire g1827_p;
  wire g1827_n;
  wire g1828_p;
  wire g1828_n;
  wire g1829_p;
  wire g1829_n;
  wire g1830_p;
  wire g1830_n;
  wire g1831_p;
  wire g1831_n;
  wire g1832_p;
  wire g1832_n;
  wire g1833_p;
  wire g1833_n;
  wire g1834_p;
  wire g1834_n;
  wire g1835_p;
  wire g1835_n;
  wire g1836_p;
  wire g1836_n;
  wire g1837_p;
  wire g1837_n;
  wire g1838_p;
  wire g1838_n;
  wire g1839_p;
  wire g1839_n;
  wire g1840_p;
  wire g1840_n;
  wire g1841_p;
  wire g1841_n;
  wire g1842_p;
  wire g1842_n;
  wire g1843_p;
  wire g1843_n;
  wire g1844_p;
  wire g1844_n;
  wire g1845_p;
  wire g1845_n;
  wire g1846_p;
  wire g1846_n;
  wire g1847_p;
  wire g1847_n;
  wire g1848_p;
  wire g1848_n;
  wire g1849_p;
  wire g1849_n;
  wire g1850_p;
  wire g1850_n;
  wire g1851_p;
  wire g1851_n;
  wire g1852_p;
  wire g1852_n;
  wire g1853_p;
  wire g1853_n;
  wire g1854_p;
  wire g1854_n;
  wire g1855_p;
  wire g1855_n;
  wire g1856_p;
  wire g1856_n;
  wire g1857_p;
  wire g1857_n;
  wire g1858_p;
  wire g1858_n;
  wire g1859_p;
  wire g1859_n;
  wire g1860_p;
  wire g1860_n;
  wire g1861_p;
  wire g1861_n;
  wire g1862_p;
  wire g1862_n;
  wire g1863_p;
  wire g1863_n;
  wire g1864_p;
  wire g1864_n;
  wire g1865_p;
  wire g1865_n;
  wire g1866_p;
  wire g1866_n;
  wire g1867_p;
  wire g1867_n;
  wire g1868_p;
  wire g1868_n;
  wire g1869_p;
  wire g1869_n;
  wire g1870_p;
  wire g1870_n;
  wire g1871_p;
  wire g1871_n;
  wire g1872_p;
  wire g1872_n;
  wire g1873_p;
  wire g1873_n;
  wire g1874_p;
  wire g1874_n;
  wire g1875_p;
  wire g1875_n;
  wire g1876_p;
  wire g1876_n;
  wire g1877_p;
  wire g1877_n;
  wire g1878_p;
  wire g1878_n;
  wire g1879_p;
  wire g1879_n;
  wire g1880_p;
  wire g1880_n;
  wire g1881_p;
  wire g1881_n;
  wire g1882_p;
  wire g1882_n;
  wire g1883_p;
  wire g1883_n;
  wire g1884_p;
  wire g1884_n;
  wire g1885_p;
  wire g1885_n;
  wire g1886_p;
  wire g1886_n;
  wire g1887_p;
  wire g1887_n;
  wire g1888_p;
  wire g1888_n;
  wire g1889_p;
  wire g1889_n;
  wire g1890_p;
  wire g1890_n;
  wire g1891_p;
  wire g1891_n;
  wire g1892_p;
  wire g1892_n;
  wire g1893_p;
  wire g1893_n;
  wire g1894_p;
  wire g1894_n;
  wire g1895_p;
  wire g1895_n;
  wire g1896_p;
  wire g1896_n;
  wire g1897_p;
  wire g1897_n;
  wire g1898_p;
  wire g1898_n;
  wire g1899_p;
  wire g1899_n;
  wire g1900_p;
  wire g1900_n;
  wire g1901_p;
  wire g1901_n;
  wire g1902_p;
  wire g1902_n;
  wire g1903_p;
  wire g1903_n;
  wire g1904_p;
  wire g1904_n;
  wire g1905_p;
  wire g1905_n;
  wire g1906_p;
  wire g1906_n;
  wire g1907_p;
  wire g1907_n;
  wire g1908_p;
  wire g1908_n;
  wire g1909_p;
  wire g1909_n;
  wire g1910_p;
  wire g1910_n;
  wire g1911_p;
  wire g1911_n;
  wire g1912_p;
  wire g1912_n;
  wire g1913_p;
  wire g1913_n;
  wire g1914_p;
  wire g1914_n;
  wire g1915_p;
  wire g1915_n;
  wire g1916_p;
  wire g1916_n;
  wire g1917_p;
  wire g1917_n;
  wire G17_p_spl_;
  wire G17_p_spl_0;
  wire G17_p_spl_00;
  wire G17_p_spl_000;
  wire G17_p_spl_001;
  wire G17_p_spl_01;
  wire G17_p_spl_010;
  wire G17_p_spl_011;
  wire G17_p_spl_1;
  wire G17_p_spl_10;
  wire G17_p_spl_100;
  wire G17_p_spl_101;
  wire G17_p_spl_11;
  wire G17_p_spl_110;
  wire G17_p_spl_111;
  wire G1_p_spl_;
  wire G1_p_spl_0;
  wire G1_p_spl_00;
  wire G1_p_spl_000;
  wire G1_p_spl_001;
  wire G1_p_spl_01;
  wire G1_p_spl_010;
  wire G1_p_spl_011;
  wire G1_p_spl_1;
  wire G1_p_spl_10;
  wire G1_p_spl_100;
  wire G1_p_spl_101;
  wire G1_p_spl_11;
  wire G1_p_spl_110;
  wire G1_p_spl_111;
  wire G2_p_spl_;
  wire G2_p_spl_0;
  wire G2_p_spl_00;
  wire G2_p_spl_000;
  wire G2_p_spl_001;
  wire G2_p_spl_01;
  wire G2_p_spl_010;
  wire G2_p_spl_011;
  wire G2_p_spl_1;
  wire G2_p_spl_10;
  wire G2_p_spl_100;
  wire G2_p_spl_101;
  wire G2_p_spl_11;
  wire G2_p_spl_110;
  wire G2_p_spl_111;
  wire G17_n_spl_;
  wire G17_n_spl_0;
  wire G17_n_spl_00;
  wire G17_n_spl_000;
  wire G17_n_spl_001;
  wire G17_n_spl_01;
  wire G17_n_spl_010;
  wire G17_n_spl_011;
  wire G17_n_spl_1;
  wire G17_n_spl_10;
  wire G17_n_spl_100;
  wire G17_n_spl_101;
  wire G17_n_spl_11;
  wire G17_n_spl_110;
  wire G2_n_spl_;
  wire G2_n_spl_0;
  wire G2_n_spl_00;
  wire G2_n_spl_000;
  wire G2_n_spl_001;
  wire G2_n_spl_01;
  wire G2_n_spl_010;
  wire G2_n_spl_011;
  wire G2_n_spl_1;
  wire G2_n_spl_10;
  wire G2_n_spl_100;
  wire G2_n_spl_101;
  wire G2_n_spl_11;
  wire G2_n_spl_110;
  wire G2_n_spl_111;
  wire G18_p_spl_;
  wire G18_p_spl_0;
  wire G18_p_spl_00;
  wire G18_p_spl_000;
  wire G18_p_spl_001;
  wire G18_p_spl_01;
  wire G18_p_spl_010;
  wire G18_p_spl_011;
  wire G18_p_spl_1;
  wire G18_p_spl_10;
  wire G18_p_spl_100;
  wire G18_p_spl_101;
  wire G18_p_spl_11;
  wire G18_p_spl_110;
  wire G18_p_spl_111;
  wire G18_n_spl_;
  wire G18_n_spl_0;
  wire G18_n_spl_00;
  wire G18_n_spl_000;
  wire G18_n_spl_001;
  wire G18_n_spl_01;
  wire G18_n_spl_010;
  wire G18_n_spl_011;
  wire G18_n_spl_1;
  wire G18_n_spl_10;
  wire G18_n_spl_100;
  wire G18_n_spl_101;
  wire G18_n_spl_11;
  wire G18_n_spl_110;
  wire G18_n_spl_111;
  wire G1_n_spl_;
  wire G1_n_spl_0;
  wire G1_n_spl_00;
  wire G1_n_spl_000;
  wire G1_n_spl_001;
  wire G1_n_spl_01;
  wire G1_n_spl_010;
  wire G1_n_spl_011;
  wire G1_n_spl_1;
  wire G1_n_spl_10;
  wire G1_n_spl_100;
  wire G1_n_spl_101;
  wire G1_n_spl_11;
  wire G1_n_spl_110;
  wire g34_p_spl_;
  wire g35_p_spl_;
  wire g34_n_spl_;
  wire g36_p_spl_;
  wire g37_n_spl_;
  wire g37_n_spl_0;
  wire G19_p_spl_;
  wire G19_p_spl_0;
  wire G19_p_spl_00;
  wire G19_p_spl_000;
  wire G19_p_spl_001;
  wire G19_p_spl_01;
  wire G19_p_spl_010;
  wire G19_p_spl_011;
  wire G19_p_spl_1;
  wire G19_p_spl_10;
  wire G19_p_spl_100;
  wire G19_p_spl_101;
  wire G19_p_spl_11;
  wire G19_p_spl_110;
  wire G19_p_spl_111;
  wire G19_n_spl_;
  wire G19_n_spl_0;
  wire G19_n_spl_00;
  wire G19_n_spl_000;
  wire G19_n_spl_001;
  wire G19_n_spl_01;
  wire G19_n_spl_010;
  wire G19_n_spl_011;
  wire G19_n_spl_1;
  wire G19_n_spl_10;
  wire G19_n_spl_100;
  wire G19_n_spl_101;
  wire G19_n_spl_11;
  wire G19_n_spl_110;
  wire G19_n_spl_111;
  wire G3_p_spl_;
  wire G3_p_spl_0;
  wire G3_p_spl_00;
  wire G3_p_spl_000;
  wire G3_p_spl_001;
  wire G3_p_spl_01;
  wire G3_p_spl_010;
  wire G3_p_spl_011;
  wire G3_p_spl_1;
  wire G3_p_spl_10;
  wire G3_p_spl_100;
  wire G3_p_spl_101;
  wire G3_p_spl_11;
  wire G3_p_spl_110;
  wire G3_p_spl_111;
  wire G3_n_spl_;
  wire G3_n_spl_0;
  wire G3_n_spl_00;
  wire G3_n_spl_000;
  wire G3_n_spl_001;
  wire G3_n_spl_01;
  wire G3_n_spl_010;
  wire G3_n_spl_011;
  wire G3_n_spl_1;
  wire G3_n_spl_10;
  wire G3_n_spl_100;
  wire G3_n_spl_101;
  wire G3_n_spl_11;
  wire G3_n_spl_110;
  wire G3_n_spl_111;
  wire g42_n_spl_;
  wire g41_p_spl_;
  wire g42_p_spl_;
  wire g41_n_spl_;
  wire g43_n_spl_;
  wire g43_p_spl_;
  wire g44_n_spl_;
  wire g44_n_spl_0;
  wire g44_p_spl_;
  wire g44_p_spl_0;
  wire g46_n_spl_;
  wire g46_p_spl_;
  wire g37_p_spl_;
  wire g47_n_spl_;
  wire g47_p_spl_;
  wire g49_n_spl_;
  wire g40_p_spl_;
  wire g50_p_spl_;
  wire G20_p_spl_;
  wire G20_p_spl_0;
  wire G20_p_spl_00;
  wire G20_p_spl_000;
  wire G20_p_spl_001;
  wire G20_p_spl_01;
  wire G20_p_spl_010;
  wire G20_p_spl_011;
  wire G20_p_spl_1;
  wire G20_p_spl_10;
  wire G20_p_spl_100;
  wire G20_p_spl_101;
  wire G20_p_spl_11;
  wire G20_p_spl_110;
  wire G20_p_spl_111;
  wire G20_n_spl_;
  wire G20_n_spl_0;
  wire G20_n_spl_00;
  wire G20_n_spl_000;
  wire G20_n_spl_001;
  wire G20_n_spl_01;
  wire G20_n_spl_010;
  wire G20_n_spl_011;
  wire G20_n_spl_1;
  wire G20_n_spl_10;
  wire G20_n_spl_100;
  wire G20_n_spl_101;
  wire G20_n_spl_11;
  wire G20_n_spl_110;
  wire G20_n_spl_111;
  wire G4_p_spl_;
  wire G4_p_spl_0;
  wire G4_p_spl_00;
  wire G4_p_spl_000;
  wire G4_p_spl_001;
  wire G4_p_spl_01;
  wire G4_p_spl_010;
  wire G4_p_spl_011;
  wire G4_p_spl_1;
  wire G4_p_spl_10;
  wire G4_p_spl_100;
  wire G4_p_spl_101;
  wire G4_p_spl_11;
  wire G4_p_spl_110;
  wire G4_p_spl_111;
  wire G4_n_spl_;
  wire G4_n_spl_0;
  wire G4_n_spl_00;
  wire G4_n_spl_000;
  wire G4_n_spl_001;
  wire G4_n_spl_01;
  wire G4_n_spl_010;
  wire G4_n_spl_011;
  wire G4_n_spl_1;
  wire G4_n_spl_10;
  wire G4_n_spl_100;
  wire G4_n_spl_101;
  wire G4_n_spl_11;
  wire G4_n_spl_110;
  wire G4_n_spl_111;
  wire g57_n_spl_;
  wire g56_p_spl_;
  wire g57_p_spl_;
  wire g56_n_spl_;
  wire g58_n_spl_;
  wire g58_p_spl_;
  wire g59_n_spl_;
  wire g59_n_spl_0;
  wire g59_p_spl_;
  wire g59_p_spl_0;
  wire g61_n_spl_;
  wire g61_p_spl_;
  wire g62_n_spl_;
  wire g62_p_spl_;
  wire g64_p_spl_;
  wire g55_n_spl_;
  wire g64_n_spl_;
  wire g55_p_spl_;
  wire g65_n_spl_;
  wire g65_p_spl_;
  wire g67_p_spl_;
  wire g54_n_spl_;
  wire g67_n_spl_;
  wire g54_p_spl_;
  wire g68_n_spl_;
  wire g68_p_spl_;
  wire g70_n_spl_;
  wire g53_p_spl_;
  wire g71_p_spl_;
  wire G21_p_spl_;
  wire G21_p_spl_0;
  wire G21_p_spl_00;
  wire G21_p_spl_000;
  wire G21_p_spl_001;
  wire G21_p_spl_01;
  wire G21_p_spl_010;
  wire G21_p_spl_011;
  wire G21_p_spl_1;
  wire G21_p_spl_10;
  wire G21_p_spl_100;
  wire G21_p_spl_101;
  wire G21_p_spl_11;
  wire G21_p_spl_110;
  wire G21_p_spl_111;
  wire G21_n_spl_;
  wire G21_n_spl_0;
  wire G21_n_spl_00;
  wire G21_n_spl_000;
  wire G21_n_spl_001;
  wire G21_n_spl_01;
  wire G21_n_spl_010;
  wire G21_n_spl_011;
  wire G21_n_spl_1;
  wire G21_n_spl_10;
  wire G21_n_spl_100;
  wire G21_n_spl_101;
  wire G21_n_spl_11;
  wire G21_n_spl_110;
  wire G21_n_spl_111;
  wire G5_p_spl_;
  wire G5_p_spl_0;
  wire G5_p_spl_00;
  wire G5_p_spl_000;
  wire G5_p_spl_001;
  wire G5_p_spl_01;
  wire G5_p_spl_010;
  wire G5_p_spl_011;
  wire G5_p_spl_1;
  wire G5_p_spl_10;
  wire G5_p_spl_100;
  wire G5_p_spl_101;
  wire G5_p_spl_11;
  wire G5_p_spl_110;
  wire G5_p_spl_111;
  wire G5_n_spl_;
  wire G5_n_spl_0;
  wire G5_n_spl_00;
  wire G5_n_spl_000;
  wire G5_n_spl_001;
  wire G5_n_spl_01;
  wire G5_n_spl_010;
  wire G5_n_spl_011;
  wire G5_n_spl_1;
  wire G5_n_spl_10;
  wire G5_n_spl_100;
  wire G5_n_spl_101;
  wire G5_n_spl_11;
  wire G5_n_spl_110;
  wire G5_n_spl_111;
  wire g80_n_spl_;
  wire g79_p_spl_;
  wire g80_p_spl_;
  wire g79_n_spl_;
  wire g81_n_spl_;
  wire g81_p_spl_;
  wire g82_n_spl_;
  wire g82_n_spl_0;
  wire g82_p_spl_;
  wire g82_p_spl_0;
  wire g84_n_spl_;
  wire g84_p_spl_;
  wire g85_n_spl_;
  wire g85_p_spl_;
  wire g87_p_spl_;
  wire g78_n_spl_;
  wire g87_n_spl_;
  wire g78_p_spl_;
  wire g88_n_spl_;
  wire g88_p_spl_;
  wire g90_p_spl_;
  wire g77_n_spl_;
  wire g90_n_spl_;
  wire g77_p_spl_;
  wire g91_n_spl_;
  wire g91_p_spl_;
  wire g93_p_spl_;
  wire g76_n_spl_;
  wire g93_n_spl_;
  wire g76_p_spl_;
  wire g94_n_spl_;
  wire g94_p_spl_;
  wire g96_p_spl_;
  wire g75_n_spl_;
  wire g96_n_spl_;
  wire g75_p_spl_;
  wire g97_n_spl_;
  wire g97_p_spl_;
  wire g99_n_spl_;
  wire g74_p_spl_;
  wire g100_p_spl_;
  wire G22_p_spl_;
  wire G22_p_spl_0;
  wire G22_p_spl_00;
  wire G22_p_spl_000;
  wire G22_p_spl_001;
  wire G22_p_spl_01;
  wire G22_p_spl_010;
  wire G22_p_spl_011;
  wire G22_p_spl_1;
  wire G22_p_spl_10;
  wire G22_p_spl_100;
  wire G22_p_spl_101;
  wire G22_p_spl_11;
  wire G22_p_spl_110;
  wire G22_p_spl_111;
  wire G22_n_spl_;
  wire G22_n_spl_0;
  wire G22_n_spl_00;
  wire G22_n_spl_000;
  wire G22_n_spl_001;
  wire G22_n_spl_01;
  wire G22_n_spl_010;
  wire G22_n_spl_011;
  wire G22_n_spl_1;
  wire G22_n_spl_10;
  wire G22_n_spl_100;
  wire G22_n_spl_101;
  wire G22_n_spl_11;
  wire G22_n_spl_110;
  wire G22_n_spl_111;
  wire G6_p_spl_;
  wire G6_p_spl_0;
  wire G6_p_spl_00;
  wire G6_p_spl_000;
  wire G6_p_spl_001;
  wire G6_p_spl_01;
  wire G6_p_spl_010;
  wire G6_p_spl_011;
  wire G6_p_spl_1;
  wire G6_p_spl_10;
  wire G6_p_spl_100;
  wire G6_p_spl_101;
  wire G6_p_spl_11;
  wire G6_p_spl_110;
  wire G6_p_spl_111;
  wire G6_n_spl_;
  wire G6_n_spl_0;
  wire G6_n_spl_00;
  wire G6_n_spl_000;
  wire G6_n_spl_001;
  wire G6_n_spl_01;
  wire G6_n_spl_010;
  wire G6_n_spl_011;
  wire G6_n_spl_1;
  wire G6_n_spl_10;
  wire G6_n_spl_100;
  wire G6_n_spl_101;
  wire G6_n_spl_11;
  wire G6_n_spl_110;
  wire G6_n_spl_111;
  wire g111_n_spl_;
  wire g110_p_spl_;
  wire g111_p_spl_;
  wire g110_n_spl_;
  wire g112_n_spl_;
  wire g112_p_spl_;
  wire g113_n_spl_;
  wire g113_n_spl_0;
  wire g113_p_spl_;
  wire g113_p_spl_0;
  wire g115_n_spl_;
  wire g115_p_spl_;
  wire g116_n_spl_;
  wire g116_p_spl_;
  wire g118_p_spl_;
  wire g109_n_spl_;
  wire g118_n_spl_;
  wire g109_p_spl_;
  wire g119_n_spl_;
  wire g119_p_spl_;
  wire g121_p_spl_;
  wire g108_n_spl_;
  wire g121_n_spl_;
  wire g108_p_spl_;
  wire g122_n_spl_;
  wire g122_p_spl_;
  wire g124_p_spl_;
  wire g107_n_spl_;
  wire g124_n_spl_;
  wire g107_p_spl_;
  wire g125_n_spl_;
  wire g125_p_spl_;
  wire g127_p_spl_;
  wire g106_n_spl_;
  wire g127_n_spl_;
  wire g106_p_spl_;
  wire g128_n_spl_;
  wire g128_p_spl_;
  wire g130_p_spl_;
  wire g105_n_spl_;
  wire g130_n_spl_;
  wire g105_p_spl_;
  wire g131_n_spl_;
  wire g131_p_spl_;
  wire g133_p_spl_;
  wire g104_n_spl_;
  wire g133_n_spl_;
  wire g104_p_spl_;
  wire g134_n_spl_;
  wire g134_p_spl_;
  wire g136_n_spl_;
  wire g103_p_spl_;
  wire g137_p_spl_;
  wire G23_p_spl_;
  wire G23_p_spl_0;
  wire G23_p_spl_00;
  wire G23_p_spl_000;
  wire G23_p_spl_001;
  wire G23_p_spl_01;
  wire G23_p_spl_010;
  wire G23_p_spl_011;
  wire G23_p_spl_1;
  wire G23_p_spl_10;
  wire G23_p_spl_100;
  wire G23_p_spl_101;
  wire G23_p_spl_11;
  wire G23_p_spl_110;
  wire G23_p_spl_111;
  wire G23_n_spl_;
  wire G23_n_spl_0;
  wire G23_n_spl_00;
  wire G23_n_spl_000;
  wire G23_n_spl_001;
  wire G23_n_spl_01;
  wire G23_n_spl_010;
  wire G23_n_spl_011;
  wire G23_n_spl_1;
  wire G23_n_spl_10;
  wire G23_n_spl_100;
  wire G23_n_spl_101;
  wire G23_n_spl_11;
  wire G23_n_spl_110;
  wire G23_n_spl_111;
  wire G7_p_spl_;
  wire G7_p_spl_0;
  wire G7_p_spl_00;
  wire G7_p_spl_000;
  wire G7_p_spl_001;
  wire G7_p_spl_01;
  wire G7_p_spl_010;
  wire G7_p_spl_011;
  wire G7_p_spl_1;
  wire G7_p_spl_10;
  wire G7_p_spl_100;
  wire G7_p_spl_101;
  wire G7_p_spl_11;
  wire G7_p_spl_110;
  wire G7_p_spl_111;
  wire G7_n_spl_;
  wire G7_n_spl_0;
  wire G7_n_spl_00;
  wire G7_n_spl_000;
  wire G7_n_spl_001;
  wire G7_n_spl_01;
  wire G7_n_spl_010;
  wire G7_n_spl_011;
  wire G7_n_spl_1;
  wire G7_n_spl_10;
  wire G7_n_spl_100;
  wire G7_n_spl_101;
  wire G7_n_spl_11;
  wire G7_n_spl_110;
  wire G7_n_spl_111;
  wire g150_n_spl_;
  wire g149_p_spl_;
  wire g150_p_spl_;
  wire g149_n_spl_;
  wire g151_n_spl_;
  wire g151_p_spl_;
  wire g152_n_spl_;
  wire g152_n_spl_0;
  wire g152_p_spl_;
  wire g152_p_spl_0;
  wire g154_n_spl_;
  wire g154_p_spl_;
  wire g155_n_spl_;
  wire g155_p_spl_;
  wire g157_p_spl_;
  wire g148_n_spl_;
  wire g157_n_spl_;
  wire g148_p_spl_;
  wire g158_n_spl_;
  wire g158_p_spl_;
  wire g160_p_spl_;
  wire g147_n_spl_;
  wire g160_n_spl_;
  wire g147_p_spl_;
  wire g161_n_spl_;
  wire g161_p_spl_;
  wire g163_p_spl_;
  wire g146_n_spl_;
  wire g163_n_spl_;
  wire g146_p_spl_;
  wire g164_n_spl_;
  wire g164_p_spl_;
  wire g166_p_spl_;
  wire g145_n_spl_;
  wire g166_n_spl_;
  wire g145_p_spl_;
  wire g167_n_spl_;
  wire g167_p_spl_;
  wire g169_p_spl_;
  wire g144_n_spl_;
  wire g169_n_spl_;
  wire g144_p_spl_;
  wire g170_n_spl_;
  wire g170_p_spl_;
  wire g172_p_spl_;
  wire g143_n_spl_;
  wire g172_n_spl_;
  wire g143_p_spl_;
  wire g173_n_spl_;
  wire g173_p_spl_;
  wire g175_p_spl_;
  wire g142_n_spl_;
  wire g175_n_spl_;
  wire g142_p_spl_;
  wire g176_n_spl_;
  wire g176_p_spl_;
  wire g178_p_spl_;
  wire g141_n_spl_;
  wire g178_n_spl_;
  wire g141_p_spl_;
  wire g179_n_spl_;
  wire g179_p_spl_;
  wire g181_n_spl_;
  wire g140_p_spl_;
  wire g182_p_spl_;
  wire G24_p_spl_;
  wire G24_p_spl_0;
  wire G24_p_spl_00;
  wire G24_p_spl_000;
  wire G24_p_spl_001;
  wire G24_p_spl_01;
  wire G24_p_spl_010;
  wire G24_p_spl_011;
  wire G24_p_spl_1;
  wire G24_p_spl_10;
  wire G24_p_spl_100;
  wire G24_p_spl_101;
  wire G24_p_spl_11;
  wire G24_p_spl_110;
  wire G24_p_spl_111;
  wire G24_n_spl_;
  wire G24_n_spl_0;
  wire G24_n_spl_00;
  wire G24_n_spl_000;
  wire G24_n_spl_001;
  wire G24_n_spl_01;
  wire G24_n_spl_010;
  wire G24_n_spl_011;
  wire G24_n_spl_1;
  wire G24_n_spl_10;
  wire G24_n_spl_100;
  wire G24_n_spl_101;
  wire G24_n_spl_11;
  wire G24_n_spl_110;
  wire G24_n_spl_111;
  wire G8_p_spl_;
  wire G8_p_spl_0;
  wire G8_p_spl_00;
  wire G8_p_spl_000;
  wire G8_p_spl_001;
  wire G8_p_spl_01;
  wire G8_p_spl_010;
  wire G8_p_spl_011;
  wire G8_p_spl_1;
  wire G8_p_spl_10;
  wire G8_p_spl_100;
  wire G8_p_spl_101;
  wire G8_p_spl_11;
  wire G8_p_spl_110;
  wire G8_p_spl_111;
  wire G8_n_spl_;
  wire G8_n_spl_0;
  wire G8_n_spl_00;
  wire G8_n_spl_000;
  wire G8_n_spl_001;
  wire G8_n_spl_01;
  wire G8_n_spl_010;
  wire G8_n_spl_011;
  wire G8_n_spl_1;
  wire G8_n_spl_10;
  wire G8_n_spl_100;
  wire G8_n_spl_101;
  wire G8_n_spl_11;
  wire G8_n_spl_110;
  wire G8_n_spl_111;
  wire g197_n_spl_;
  wire g196_p_spl_;
  wire g197_p_spl_;
  wire g196_n_spl_;
  wire g198_n_spl_;
  wire g198_p_spl_;
  wire g199_n_spl_;
  wire g199_n_spl_0;
  wire g199_p_spl_;
  wire g199_p_spl_0;
  wire g201_n_spl_;
  wire g201_p_spl_;
  wire g202_n_spl_;
  wire g202_p_spl_;
  wire g204_p_spl_;
  wire g195_n_spl_;
  wire g204_n_spl_;
  wire g195_p_spl_;
  wire g205_n_spl_;
  wire g205_p_spl_;
  wire g207_p_spl_;
  wire g194_n_spl_;
  wire g207_n_spl_;
  wire g194_p_spl_;
  wire g208_n_spl_;
  wire g208_p_spl_;
  wire g210_p_spl_;
  wire g193_n_spl_;
  wire g210_n_spl_;
  wire g193_p_spl_;
  wire g211_n_spl_;
  wire g211_p_spl_;
  wire g213_p_spl_;
  wire g192_n_spl_;
  wire g213_n_spl_;
  wire g192_p_spl_;
  wire g214_n_spl_;
  wire g214_p_spl_;
  wire g216_p_spl_;
  wire g191_n_spl_;
  wire g216_n_spl_;
  wire g191_p_spl_;
  wire g217_n_spl_;
  wire g217_p_spl_;
  wire g219_p_spl_;
  wire g190_n_spl_;
  wire g219_n_spl_;
  wire g190_p_spl_;
  wire g220_n_spl_;
  wire g220_p_spl_;
  wire g222_p_spl_;
  wire g189_n_spl_;
  wire g222_n_spl_;
  wire g189_p_spl_;
  wire g223_n_spl_;
  wire g223_p_spl_;
  wire g225_p_spl_;
  wire g188_n_spl_;
  wire g225_n_spl_;
  wire g188_p_spl_;
  wire g226_n_spl_;
  wire g226_p_spl_;
  wire g228_p_spl_;
  wire g187_n_spl_;
  wire g228_n_spl_;
  wire g187_p_spl_;
  wire g229_n_spl_;
  wire g229_p_spl_;
  wire g231_p_spl_;
  wire g186_n_spl_;
  wire g231_n_spl_;
  wire g186_p_spl_;
  wire g232_n_spl_;
  wire g232_p_spl_;
  wire g234_n_spl_;
  wire g185_p_spl_;
  wire g235_p_spl_;
  wire G25_p_spl_;
  wire G25_p_spl_0;
  wire G25_p_spl_00;
  wire G25_p_spl_000;
  wire G25_p_spl_001;
  wire G25_p_spl_01;
  wire G25_p_spl_010;
  wire G25_p_spl_011;
  wire G25_p_spl_1;
  wire G25_p_spl_10;
  wire G25_p_spl_100;
  wire G25_p_spl_101;
  wire G25_p_spl_11;
  wire G25_p_spl_110;
  wire G25_p_spl_111;
  wire G25_n_spl_;
  wire G25_n_spl_0;
  wire G25_n_spl_00;
  wire G25_n_spl_000;
  wire G25_n_spl_001;
  wire G25_n_spl_01;
  wire G25_n_spl_010;
  wire G25_n_spl_011;
  wire G25_n_spl_1;
  wire G25_n_spl_10;
  wire G25_n_spl_100;
  wire G25_n_spl_101;
  wire G25_n_spl_11;
  wire G25_n_spl_110;
  wire G25_n_spl_111;
  wire G9_p_spl_;
  wire G9_p_spl_0;
  wire G9_p_spl_00;
  wire G9_p_spl_000;
  wire G9_p_spl_001;
  wire G9_p_spl_01;
  wire G9_p_spl_010;
  wire G9_p_spl_011;
  wire G9_p_spl_1;
  wire G9_p_spl_10;
  wire G9_p_spl_100;
  wire G9_p_spl_101;
  wire G9_p_spl_11;
  wire G9_p_spl_110;
  wire G9_p_spl_111;
  wire G9_n_spl_;
  wire G9_n_spl_0;
  wire G9_n_spl_00;
  wire G9_n_spl_000;
  wire G9_n_spl_001;
  wire G9_n_spl_01;
  wire G9_n_spl_010;
  wire G9_n_spl_011;
  wire G9_n_spl_1;
  wire G9_n_spl_10;
  wire G9_n_spl_100;
  wire G9_n_spl_101;
  wire G9_n_spl_11;
  wire G9_n_spl_110;
  wire G9_n_spl_111;
  wire g252_n_spl_;
  wire g251_p_spl_;
  wire g252_p_spl_;
  wire g251_n_spl_;
  wire g253_n_spl_;
  wire g253_p_spl_;
  wire g254_n_spl_;
  wire g254_n_spl_0;
  wire g254_p_spl_;
  wire g254_p_spl_0;
  wire g256_n_spl_;
  wire g256_p_spl_;
  wire g257_n_spl_;
  wire g257_p_spl_;
  wire g259_p_spl_;
  wire g250_n_spl_;
  wire g259_n_spl_;
  wire g250_p_spl_;
  wire g260_n_spl_;
  wire g260_p_spl_;
  wire g262_p_spl_;
  wire g249_n_spl_;
  wire g262_n_spl_;
  wire g249_p_spl_;
  wire g263_n_spl_;
  wire g263_p_spl_;
  wire g265_p_spl_;
  wire g248_n_spl_;
  wire g265_n_spl_;
  wire g248_p_spl_;
  wire g266_n_spl_;
  wire g266_p_spl_;
  wire g268_p_spl_;
  wire g247_n_spl_;
  wire g268_n_spl_;
  wire g247_p_spl_;
  wire g269_n_spl_;
  wire g269_p_spl_;
  wire g271_p_spl_;
  wire g246_n_spl_;
  wire g271_n_spl_;
  wire g246_p_spl_;
  wire g272_n_spl_;
  wire g272_p_spl_;
  wire g274_p_spl_;
  wire g245_n_spl_;
  wire g274_n_spl_;
  wire g245_p_spl_;
  wire g275_n_spl_;
  wire g275_p_spl_;
  wire g277_p_spl_;
  wire g244_n_spl_;
  wire g277_n_spl_;
  wire g244_p_spl_;
  wire g278_n_spl_;
  wire g278_p_spl_;
  wire g280_p_spl_;
  wire g243_n_spl_;
  wire g280_n_spl_;
  wire g243_p_spl_;
  wire g281_n_spl_;
  wire g281_p_spl_;
  wire g283_p_spl_;
  wire g242_n_spl_;
  wire g283_n_spl_;
  wire g242_p_spl_;
  wire g284_n_spl_;
  wire g284_p_spl_;
  wire g286_p_spl_;
  wire g241_n_spl_;
  wire g286_n_spl_;
  wire g241_p_spl_;
  wire g287_n_spl_;
  wire g287_p_spl_;
  wire g289_p_spl_;
  wire g240_n_spl_;
  wire g289_n_spl_;
  wire g240_p_spl_;
  wire g290_n_spl_;
  wire g290_p_spl_;
  wire g292_p_spl_;
  wire g239_n_spl_;
  wire g292_n_spl_;
  wire g239_p_spl_;
  wire g293_n_spl_;
  wire g293_p_spl_;
  wire g295_n_spl_;
  wire g238_p_spl_;
  wire g296_p_spl_;
  wire G26_p_spl_;
  wire G26_p_spl_0;
  wire G26_p_spl_00;
  wire G26_p_spl_000;
  wire G26_p_spl_001;
  wire G26_p_spl_01;
  wire G26_p_spl_010;
  wire G26_p_spl_011;
  wire G26_p_spl_1;
  wire G26_p_spl_10;
  wire G26_p_spl_100;
  wire G26_p_spl_101;
  wire G26_p_spl_11;
  wire G26_p_spl_110;
  wire G26_p_spl_111;
  wire G26_n_spl_;
  wire G26_n_spl_0;
  wire G26_n_spl_00;
  wire G26_n_spl_000;
  wire G26_n_spl_001;
  wire G26_n_spl_01;
  wire G26_n_spl_010;
  wire G26_n_spl_011;
  wire G26_n_spl_1;
  wire G26_n_spl_10;
  wire G26_n_spl_100;
  wire G26_n_spl_101;
  wire G26_n_spl_11;
  wire G26_n_spl_110;
  wire G26_n_spl_111;
  wire G10_p_spl_;
  wire G10_p_spl_0;
  wire G10_p_spl_00;
  wire G10_p_spl_000;
  wire G10_p_spl_001;
  wire G10_p_spl_01;
  wire G10_p_spl_010;
  wire G10_p_spl_011;
  wire G10_p_spl_1;
  wire G10_p_spl_10;
  wire G10_p_spl_100;
  wire G10_p_spl_101;
  wire G10_p_spl_11;
  wire G10_p_spl_110;
  wire G10_p_spl_111;
  wire G10_n_spl_;
  wire G10_n_spl_0;
  wire G10_n_spl_00;
  wire G10_n_spl_000;
  wire G10_n_spl_001;
  wire G10_n_spl_01;
  wire G10_n_spl_010;
  wire G10_n_spl_011;
  wire G10_n_spl_1;
  wire G10_n_spl_10;
  wire G10_n_spl_100;
  wire G10_n_spl_101;
  wire G10_n_spl_11;
  wire G10_n_spl_110;
  wire G10_n_spl_111;
  wire g315_n_spl_;
  wire g314_p_spl_;
  wire g315_p_spl_;
  wire g314_n_spl_;
  wire g316_n_spl_;
  wire g316_p_spl_;
  wire g317_n_spl_;
  wire g317_n_spl_0;
  wire g317_p_spl_;
  wire g317_p_spl_0;
  wire g319_n_spl_;
  wire g319_p_spl_;
  wire g320_n_spl_;
  wire g320_p_spl_;
  wire g322_p_spl_;
  wire g313_n_spl_;
  wire g322_n_spl_;
  wire g313_p_spl_;
  wire g323_n_spl_;
  wire g323_p_spl_;
  wire g325_p_spl_;
  wire g312_n_spl_;
  wire g325_n_spl_;
  wire g312_p_spl_;
  wire g326_n_spl_;
  wire g326_p_spl_;
  wire g328_p_spl_;
  wire g311_n_spl_;
  wire g328_n_spl_;
  wire g311_p_spl_;
  wire g329_n_spl_;
  wire g329_p_spl_;
  wire g331_p_spl_;
  wire g310_n_spl_;
  wire g331_n_spl_;
  wire g310_p_spl_;
  wire g332_n_spl_;
  wire g332_p_spl_;
  wire g334_p_spl_;
  wire g309_n_spl_;
  wire g334_n_spl_;
  wire g309_p_spl_;
  wire g335_n_spl_;
  wire g335_p_spl_;
  wire g337_p_spl_;
  wire g308_n_spl_;
  wire g337_n_spl_;
  wire g308_p_spl_;
  wire g338_n_spl_;
  wire g338_p_spl_;
  wire g340_p_spl_;
  wire g307_n_spl_;
  wire g340_n_spl_;
  wire g307_p_spl_;
  wire g341_n_spl_;
  wire g341_p_spl_;
  wire g343_p_spl_;
  wire g306_n_spl_;
  wire g343_n_spl_;
  wire g306_p_spl_;
  wire g344_n_spl_;
  wire g344_p_spl_;
  wire g346_p_spl_;
  wire g305_n_spl_;
  wire g346_n_spl_;
  wire g305_p_spl_;
  wire g347_n_spl_;
  wire g347_p_spl_;
  wire g349_p_spl_;
  wire g304_n_spl_;
  wire g349_n_spl_;
  wire g304_p_spl_;
  wire g350_n_spl_;
  wire g350_p_spl_;
  wire g352_p_spl_;
  wire g303_n_spl_;
  wire g352_n_spl_;
  wire g303_p_spl_;
  wire g353_n_spl_;
  wire g353_p_spl_;
  wire g355_p_spl_;
  wire g302_n_spl_;
  wire g355_n_spl_;
  wire g302_p_spl_;
  wire g356_n_spl_;
  wire g356_p_spl_;
  wire g358_p_spl_;
  wire g301_n_spl_;
  wire g358_n_spl_;
  wire g301_p_spl_;
  wire g359_n_spl_;
  wire g359_p_spl_;
  wire g361_p_spl_;
  wire g300_n_spl_;
  wire g361_n_spl_;
  wire g300_p_spl_;
  wire g362_n_spl_;
  wire g362_p_spl_;
  wire g364_n_spl_;
  wire g299_p_spl_;
  wire g365_p_spl_;
  wire G27_p_spl_;
  wire G27_p_spl_0;
  wire G27_p_spl_00;
  wire G27_p_spl_000;
  wire G27_p_spl_001;
  wire G27_p_spl_01;
  wire G27_p_spl_010;
  wire G27_p_spl_011;
  wire G27_p_spl_1;
  wire G27_p_spl_10;
  wire G27_p_spl_100;
  wire G27_p_spl_101;
  wire G27_p_spl_11;
  wire G27_p_spl_110;
  wire G27_p_spl_111;
  wire G27_n_spl_;
  wire G27_n_spl_0;
  wire G27_n_spl_00;
  wire G27_n_spl_000;
  wire G27_n_spl_001;
  wire G27_n_spl_01;
  wire G27_n_spl_010;
  wire G27_n_spl_011;
  wire G27_n_spl_1;
  wire G27_n_spl_10;
  wire G27_n_spl_100;
  wire G27_n_spl_101;
  wire G27_n_spl_11;
  wire G27_n_spl_110;
  wire G27_n_spl_111;
  wire G11_p_spl_;
  wire G11_p_spl_0;
  wire G11_p_spl_00;
  wire G11_p_spl_000;
  wire G11_p_spl_001;
  wire G11_p_spl_01;
  wire G11_p_spl_010;
  wire G11_p_spl_011;
  wire G11_p_spl_1;
  wire G11_p_spl_10;
  wire G11_p_spl_100;
  wire G11_p_spl_101;
  wire G11_p_spl_11;
  wire G11_p_spl_110;
  wire G11_p_spl_111;
  wire G11_n_spl_;
  wire G11_n_spl_0;
  wire G11_n_spl_00;
  wire G11_n_spl_000;
  wire G11_n_spl_001;
  wire G11_n_spl_01;
  wire G11_n_spl_010;
  wire G11_n_spl_011;
  wire G11_n_spl_1;
  wire G11_n_spl_10;
  wire G11_n_spl_100;
  wire G11_n_spl_101;
  wire G11_n_spl_11;
  wire G11_n_spl_110;
  wire G11_n_spl_111;
  wire g386_n_spl_;
  wire g385_p_spl_;
  wire g386_p_spl_;
  wire g385_n_spl_;
  wire g387_n_spl_;
  wire g387_p_spl_;
  wire g388_n_spl_;
  wire g388_n_spl_0;
  wire g388_p_spl_;
  wire g388_p_spl_0;
  wire g390_n_spl_;
  wire g390_p_spl_;
  wire g391_n_spl_;
  wire g391_p_spl_;
  wire g393_p_spl_;
  wire g384_n_spl_;
  wire g393_n_spl_;
  wire g384_p_spl_;
  wire g394_n_spl_;
  wire g394_p_spl_;
  wire g396_p_spl_;
  wire g383_n_spl_;
  wire g396_n_spl_;
  wire g383_p_spl_;
  wire g397_n_spl_;
  wire g397_p_spl_;
  wire g399_p_spl_;
  wire g382_n_spl_;
  wire g399_n_spl_;
  wire g382_p_spl_;
  wire g400_n_spl_;
  wire g400_p_spl_;
  wire g402_p_spl_;
  wire g381_n_spl_;
  wire g402_n_spl_;
  wire g381_p_spl_;
  wire g403_n_spl_;
  wire g403_p_spl_;
  wire g405_p_spl_;
  wire g380_n_spl_;
  wire g405_n_spl_;
  wire g380_p_spl_;
  wire g406_n_spl_;
  wire g406_p_spl_;
  wire g408_p_spl_;
  wire g379_n_spl_;
  wire g408_n_spl_;
  wire g379_p_spl_;
  wire g409_n_spl_;
  wire g409_p_spl_;
  wire g411_p_spl_;
  wire g378_n_spl_;
  wire g411_n_spl_;
  wire g378_p_spl_;
  wire g412_n_spl_;
  wire g412_p_spl_;
  wire g414_p_spl_;
  wire g377_n_spl_;
  wire g414_n_spl_;
  wire g377_p_spl_;
  wire g415_n_spl_;
  wire g415_p_spl_;
  wire g417_p_spl_;
  wire g376_n_spl_;
  wire g417_n_spl_;
  wire g376_p_spl_;
  wire g418_n_spl_;
  wire g418_p_spl_;
  wire g420_p_spl_;
  wire g375_n_spl_;
  wire g420_n_spl_;
  wire g375_p_spl_;
  wire g421_n_spl_;
  wire g421_p_spl_;
  wire g423_p_spl_;
  wire g374_n_spl_;
  wire g423_n_spl_;
  wire g374_p_spl_;
  wire g424_n_spl_;
  wire g424_p_spl_;
  wire g426_p_spl_;
  wire g373_n_spl_;
  wire g426_n_spl_;
  wire g373_p_spl_;
  wire g427_n_spl_;
  wire g427_p_spl_;
  wire g429_p_spl_;
  wire g372_n_spl_;
  wire g429_n_spl_;
  wire g372_p_spl_;
  wire g430_n_spl_;
  wire g430_p_spl_;
  wire g432_p_spl_;
  wire g371_n_spl_;
  wire g432_n_spl_;
  wire g371_p_spl_;
  wire g433_n_spl_;
  wire g433_p_spl_;
  wire g435_p_spl_;
  wire g370_n_spl_;
  wire g435_n_spl_;
  wire g370_p_spl_;
  wire g436_n_spl_;
  wire g436_p_spl_;
  wire g438_p_spl_;
  wire g369_n_spl_;
  wire g438_n_spl_;
  wire g369_p_spl_;
  wire g439_n_spl_;
  wire g439_p_spl_;
  wire g441_n_spl_;
  wire g368_p_spl_;
  wire g442_p_spl_;
  wire G28_p_spl_;
  wire G28_p_spl_0;
  wire G28_p_spl_00;
  wire G28_p_spl_000;
  wire G28_p_spl_001;
  wire G28_p_spl_01;
  wire G28_p_spl_010;
  wire G28_p_spl_011;
  wire G28_p_spl_1;
  wire G28_p_spl_10;
  wire G28_p_spl_100;
  wire G28_p_spl_101;
  wire G28_p_spl_11;
  wire G28_p_spl_110;
  wire G28_p_spl_111;
  wire G28_n_spl_;
  wire G28_n_spl_0;
  wire G28_n_spl_00;
  wire G28_n_spl_000;
  wire G28_n_spl_001;
  wire G28_n_spl_01;
  wire G28_n_spl_010;
  wire G28_n_spl_011;
  wire G28_n_spl_1;
  wire G28_n_spl_10;
  wire G28_n_spl_100;
  wire G28_n_spl_101;
  wire G28_n_spl_11;
  wire G28_n_spl_110;
  wire G28_n_spl_111;
  wire G12_p_spl_;
  wire G12_p_spl_0;
  wire G12_p_spl_00;
  wire G12_p_spl_000;
  wire G12_p_spl_001;
  wire G12_p_spl_01;
  wire G12_p_spl_010;
  wire G12_p_spl_011;
  wire G12_p_spl_1;
  wire G12_p_spl_10;
  wire G12_p_spl_100;
  wire G12_p_spl_101;
  wire G12_p_spl_11;
  wire G12_p_spl_110;
  wire G12_p_spl_111;
  wire G12_n_spl_;
  wire G12_n_spl_0;
  wire G12_n_spl_00;
  wire G12_n_spl_000;
  wire G12_n_spl_001;
  wire G12_n_spl_01;
  wire G12_n_spl_010;
  wire G12_n_spl_011;
  wire G12_n_spl_1;
  wire G12_n_spl_10;
  wire G12_n_spl_100;
  wire G12_n_spl_101;
  wire G12_n_spl_11;
  wire G12_n_spl_110;
  wire G12_n_spl_111;
  wire g465_n_spl_;
  wire g464_p_spl_;
  wire g465_p_spl_;
  wire g464_n_spl_;
  wire g466_n_spl_;
  wire g466_p_spl_;
  wire g467_n_spl_;
  wire g467_n_spl_0;
  wire g467_p_spl_;
  wire g467_p_spl_0;
  wire g469_n_spl_;
  wire g469_p_spl_;
  wire g470_n_spl_;
  wire g470_p_spl_;
  wire g472_p_spl_;
  wire g463_n_spl_;
  wire g472_n_spl_;
  wire g463_p_spl_;
  wire g473_n_spl_;
  wire g473_p_spl_;
  wire g475_p_spl_;
  wire g462_n_spl_;
  wire g475_n_spl_;
  wire g462_p_spl_;
  wire g476_n_spl_;
  wire g476_p_spl_;
  wire g478_p_spl_;
  wire g461_n_spl_;
  wire g478_n_spl_;
  wire g461_p_spl_;
  wire g479_n_spl_;
  wire g479_p_spl_;
  wire g481_p_spl_;
  wire g460_n_spl_;
  wire g481_n_spl_;
  wire g460_p_spl_;
  wire g482_n_spl_;
  wire g482_p_spl_;
  wire g484_p_spl_;
  wire g459_n_spl_;
  wire g484_n_spl_;
  wire g459_p_spl_;
  wire g485_n_spl_;
  wire g485_p_spl_;
  wire g487_p_spl_;
  wire g458_n_spl_;
  wire g487_n_spl_;
  wire g458_p_spl_;
  wire g488_n_spl_;
  wire g488_p_spl_;
  wire g490_p_spl_;
  wire g457_n_spl_;
  wire g490_n_spl_;
  wire g457_p_spl_;
  wire g491_n_spl_;
  wire g491_p_spl_;
  wire g493_p_spl_;
  wire g456_n_spl_;
  wire g493_n_spl_;
  wire g456_p_spl_;
  wire g494_n_spl_;
  wire g494_p_spl_;
  wire g496_p_spl_;
  wire g455_n_spl_;
  wire g496_n_spl_;
  wire g455_p_spl_;
  wire g497_n_spl_;
  wire g497_p_spl_;
  wire g499_p_spl_;
  wire g454_n_spl_;
  wire g499_n_spl_;
  wire g454_p_spl_;
  wire g500_n_spl_;
  wire g500_p_spl_;
  wire g502_p_spl_;
  wire g453_n_spl_;
  wire g502_n_spl_;
  wire g453_p_spl_;
  wire g503_n_spl_;
  wire g503_p_spl_;
  wire g505_p_spl_;
  wire g452_n_spl_;
  wire g505_n_spl_;
  wire g452_p_spl_;
  wire g506_n_spl_;
  wire g506_p_spl_;
  wire g508_p_spl_;
  wire g451_n_spl_;
  wire g508_n_spl_;
  wire g451_p_spl_;
  wire g509_n_spl_;
  wire g509_p_spl_;
  wire g511_p_spl_;
  wire g450_n_spl_;
  wire g511_n_spl_;
  wire g450_p_spl_;
  wire g512_n_spl_;
  wire g512_p_spl_;
  wire g514_p_spl_;
  wire g449_n_spl_;
  wire g514_n_spl_;
  wire g449_p_spl_;
  wire g515_n_spl_;
  wire g515_p_spl_;
  wire g517_p_spl_;
  wire g448_n_spl_;
  wire g517_n_spl_;
  wire g448_p_spl_;
  wire g518_n_spl_;
  wire g518_p_spl_;
  wire g520_p_spl_;
  wire g447_n_spl_;
  wire g520_n_spl_;
  wire g447_p_spl_;
  wire g521_n_spl_;
  wire g521_p_spl_;
  wire g523_p_spl_;
  wire g446_n_spl_;
  wire g523_n_spl_;
  wire g446_p_spl_;
  wire g524_n_spl_;
  wire g524_p_spl_;
  wire g526_n_spl_;
  wire g445_p_spl_;
  wire g527_p_spl_;
  wire G29_p_spl_;
  wire G29_p_spl_0;
  wire G29_p_spl_00;
  wire G29_p_spl_000;
  wire G29_p_spl_001;
  wire G29_p_spl_01;
  wire G29_p_spl_010;
  wire G29_p_spl_011;
  wire G29_p_spl_1;
  wire G29_p_spl_10;
  wire G29_p_spl_100;
  wire G29_p_spl_101;
  wire G29_p_spl_11;
  wire G29_p_spl_110;
  wire G29_p_spl_111;
  wire G29_n_spl_;
  wire G29_n_spl_0;
  wire G29_n_spl_00;
  wire G29_n_spl_000;
  wire G29_n_spl_001;
  wire G29_n_spl_01;
  wire G29_n_spl_010;
  wire G29_n_spl_011;
  wire G29_n_spl_1;
  wire G29_n_spl_10;
  wire G29_n_spl_100;
  wire G29_n_spl_101;
  wire G29_n_spl_11;
  wire G29_n_spl_110;
  wire G29_n_spl_111;
  wire G13_p_spl_;
  wire G13_p_spl_0;
  wire G13_p_spl_00;
  wire G13_p_spl_000;
  wire G13_p_spl_001;
  wire G13_p_spl_01;
  wire G13_p_spl_010;
  wire G13_p_spl_011;
  wire G13_p_spl_1;
  wire G13_p_spl_10;
  wire G13_p_spl_100;
  wire G13_p_spl_101;
  wire G13_p_spl_11;
  wire G13_p_spl_110;
  wire G13_p_spl_111;
  wire G13_n_spl_;
  wire G13_n_spl_0;
  wire G13_n_spl_00;
  wire G13_n_spl_000;
  wire G13_n_spl_001;
  wire G13_n_spl_01;
  wire G13_n_spl_010;
  wire G13_n_spl_011;
  wire G13_n_spl_1;
  wire G13_n_spl_10;
  wire G13_n_spl_100;
  wire G13_n_spl_101;
  wire G13_n_spl_11;
  wire G13_n_spl_110;
  wire G13_n_spl_111;
  wire g552_n_spl_;
  wire g551_p_spl_;
  wire g552_p_spl_;
  wire g551_n_spl_;
  wire g553_n_spl_;
  wire g553_p_spl_;
  wire g554_n_spl_;
  wire g554_n_spl_0;
  wire g554_p_spl_;
  wire g554_p_spl_0;
  wire g556_n_spl_;
  wire g556_p_spl_;
  wire g557_n_spl_;
  wire g557_p_spl_;
  wire g559_p_spl_;
  wire g550_n_spl_;
  wire g559_n_spl_;
  wire g550_p_spl_;
  wire g560_n_spl_;
  wire g560_p_spl_;
  wire g562_p_spl_;
  wire g549_n_spl_;
  wire g562_n_spl_;
  wire g549_p_spl_;
  wire g563_n_spl_;
  wire g563_p_spl_;
  wire g565_p_spl_;
  wire g548_n_spl_;
  wire g565_n_spl_;
  wire g548_p_spl_;
  wire g566_n_spl_;
  wire g566_p_spl_;
  wire g568_p_spl_;
  wire g547_n_spl_;
  wire g568_n_spl_;
  wire g547_p_spl_;
  wire g569_n_spl_;
  wire g569_p_spl_;
  wire g571_p_spl_;
  wire g546_n_spl_;
  wire g571_n_spl_;
  wire g546_p_spl_;
  wire g572_n_spl_;
  wire g572_p_spl_;
  wire g574_p_spl_;
  wire g545_n_spl_;
  wire g574_n_spl_;
  wire g545_p_spl_;
  wire g575_n_spl_;
  wire g575_p_spl_;
  wire g577_p_spl_;
  wire g544_n_spl_;
  wire g577_n_spl_;
  wire g544_p_spl_;
  wire g578_n_spl_;
  wire g578_p_spl_;
  wire g580_p_spl_;
  wire g543_n_spl_;
  wire g580_n_spl_;
  wire g543_p_spl_;
  wire g581_n_spl_;
  wire g581_p_spl_;
  wire g583_p_spl_;
  wire g542_n_spl_;
  wire g583_n_spl_;
  wire g542_p_spl_;
  wire g584_n_spl_;
  wire g584_p_spl_;
  wire g586_p_spl_;
  wire g541_n_spl_;
  wire g586_n_spl_;
  wire g541_p_spl_;
  wire g587_n_spl_;
  wire g587_p_spl_;
  wire g589_p_spl_;
  wire g540_n_spl_;
  wire g589_n_spl_;
  wire g540_p_spl_;
  wire g590_n_spl_;
  wire g590_p_spl_;
  wire g592_p_spl_;
  wire g539_n_spl_;
  wire g592_n_spl_;
  wire g539_p_spl_;
  wire g593_n_spl_;
  wire g593_p_spl_;
  wire g595_p_spl_;
  wire g538_n_spl_;
  wire g595_n_spl_;
  wire g538_p_spl_;
  wire g596_n_spl_;
  wire g596_p_spl_;
  wire g598_p_spl_;
  wire g537_n_spl_;
  wire g598_n_spl_;
  wire g537_p_spl_;
  wire g599_n_spl_;
  wire g599_p_spl_;
  wire g601_p_spl_;
  wire g536_n_spl_;
  wire g601_n_spl_;
  wire g536_p_spl_;
  wire g602_n_spl_;
  wire g602_p_spl_;
  wire g604_p_spl_;
  wire g535_n_spl_;
  wire g604_n_spl_;
  wire g535_p_spl_;
  wire g605_n_spl_;
  wire g605_p_spl_;
  wire g607_p_spl_;
  wire g534_n_spl_;
  wire g607_n_spl_;
  wire g534_p_spl_;
  wire g608_n_spl_;
  wire g608_p_spl_;
  wire g610_p_spl_;
  wire g533_n_spl_;
  wire g610_n_spl_;
  wire g533_p_spl_;
  wire g611_n_spl_;
  wire g611_p_spl_;
  wire g613_p_spl_;
  wire g532_n_spl_;
  wire g613_n_spl_;
  wire g532_p_spl_;
  wire g614_n_spl_;
  wire g614_p_spl_;
  wire g616_p_spl_;
  wire g531_n_spl_;
  wire g616_n_spl_;
  wire g531_p_spl_;
  wire g617_n_spl_;
  wire g617_p_spl_;
  wire g619_n_spl_;
  wire g530_p_spl_;
  wire g620_p_spl_;
  wire G30_p_spl_;
  wire G30_p_spl_0;
  wire G30_p_spl_00;
  wire G30_p_spl_000;
  wire G30_p_spl_001;
  wire G30_p_spl_01;
  wire G30_p_spl_010;
  wire G30_p_spl_011;
  wire G30_p_spl_1;
  wire G30_p_spl_10;
  wire G30_p_spl_100;
  wire G30_p_spl_101;
  wire G30_p_spl_11;
  wire G30_p_spl_110;
  wire G30_p_spl_111;
  wire G30_n_spl_;
  wire G30_n_spl_0;
  wire G30_n_spl_00;
  wire G30_n_spl_000;
  wire G30_n_spl_001;
  wire G30_n_spl_01;
  wire G30_n_spl_010;
  wire G30_n_spl_011;
  wire G30_n_spl_1;
  wire G30_n_spl_10;
  wire G30_n_spl_100;
  wire G30_n_spl_101;
  wire G30_n_spl_11;
  wire G30_n_spl_110;
  wire G30_n_spl_111;
  wire G14_p_spl_;
  wire G14_p_spl_0;
  wire G14_p_spl_00;
  wire G14_p_spl_000;
  wire G14_p_spl_001;
  wire G14_p_spl_01;
  wire G14_p_spl_010;
  wire G14_p_spl_011;
  wire G14_p_spl_1;
  wire G14_p_spl_10;
  wire G14_p_spl_100;
  wire G14_p_spl_101;
  wire G14_p_spl_11;
  wire G14_p_spl_110;
  wire G14_p_spl_111;
  wire G14_n_spl_;
  wire G14_n_spl_0;
  wire G14_n_spl_00;
  wire G14_n_spl_000;
  wire G14_n_spl_001;
  wire G14_n_spl_01;
  wire G14_n_spl_010;
  wire G14_n_spl_011;
  wire G14_n_spl_1;
  wire G14_n_spl_10;
  wire G14_n_spl_100;
  wire G14_n_spl_101;
  wire G14_n_spl_11;
  wire G14_n_spl_110;
  wire G14_n_spl_111;
  wire g647_n_spl_;
  wire g646_p_spl_;
  wire g647_p_spl_;
  wire g646_n_spl_;
  wire g648_n_spl_;
  wire g648_p_spl_;
  wire g649_n_spl_;
  wire g649_n_spl_0;
  wire g649_p_spl_;
  wire g649_p_spl_0;
  wire g651_n_spl_;
  wire g651_p_spl_;
  wire g652_n_spl_;
  wire g652_p_spl_;
  wire g654_p_spl_;
  wire g645_n_spl_;
  wire g654_n_spl_;
  wire g645_p_spl_;
  wire g655_n_spl_;
  wire g655_p_spl_;
  wire g657_p_spl_;
  wire g644_n_spl_;
  wire g657_n_spl_;
  wire g644_p_spl_;
  wire g658_n_spl_;
  wire g658_p_spl_;
  wire g660_p_spl_;
  wire g643_n_spl_;
  wire g660_n_spl_;
  wire g643_p_spl_;
  wire g661_n_spl_;
  wire g661_p_spl_;
  wire g663_p_spl_;
  wire g642_n_spl_;
  wire g663_n_spl_;
  wire g642_p_spl_;
  wire g664_n_spl_;
  wire g664_p_spl_;
  wire g666_p_spl_;
  wire g641_n_spl_;
  wire g666_n_spl_;
  wire g641_p_spl_;
  wire g667_n_spl_;
  wire g667_p_spl_;
  wire g669_p_spl_;
  wire g640_n_spl_;
  wire g669_n_spl_;
  wire g640_p_spl_;
  wire g670_n_spl_;
  wire g670_p_spl_;
  wire g672_p_spl_;
  wire g639_n_spl_;
  wire g672_n_spl_;
  wire g639_p_spl_;
  wire g673_n_spl_;
  wire g673_p_spl_;
  wire g675_p_spl_;
  wire g638_n_spl_;
  wire g675_n_spl_;
  wire g638_p_spl_;
  wire g676_n_spl_;
  wire g676_p_spl_;
  wire g678_p_spl_;
  wire g637_n_spl_;
  wire g678_n_spl_;
  wire g637_p_spl_;
  wire g679_n_spl_;
  wire g679_p_spl_;
  wire g681_p_spl_;
  wire g636_n_spl_;
  wire g681_n_spl_;
  wire g636_p_spl_;
  wire g682_n_spl_;
  wire g682_p_spl_;
  wire g684_p_spl_;
  wire g635_n_spl_;
  wire g684_n_spl_;
  wire g635_p_spl_;
  wire g685_n_spl_;
  wire g685_p_spl_;
  wire g687_p_spl_;
  wire g634_n_spl_;
  wire g687_n_spl_;
  wire g634_p_spl_;
  wire g688_n_spl_;
  wire g688_p_spl_;
  wire g690_p_spl_;
  wire g633_n_spl_;
  wire g690_n_spl_;
  wire g633_p_spl_;
  wire g691_n_spl_;
  wire g691_p_spl_;
  wire g693_p_spl_;
  wire g632_n_spl_;
  wire g693_n_spl_;
  wire g632_p_spl_;
  wire g694_n_spl_;
  wire g694_p_spl_;
  wire g696_p_spl_;
  wire g631_n_spl_;
  wire g696_n_spl_;
  wire g631_p_spl_;
  wire g697_n_spl_;
  wire g697_p_spl_;
  wire g699_p_spl_;
  wire g630_n_spl_;
  wire g699_n_spl_;
  wire g630_p_spl_;
  wire g700_n_spl_;
  wire g700_p_spl_;
  wire g702_p_spl_;
  wire g629_n_spl_;
  wire g702_n_spl_;
  wire g629_p_spl_;
  wire g703_n_spl_;
  wire g703_p_spl_;
  wire g705_p_spl_;
  wire g628_n_spl_;
  wire g705_n_spl_;
  wire g628_p_spl_;
  wire g706_n_spl_;
  wire g706_p_spl_;
  wire g708_p_spl_;
  wire g627_n_spl_;
  wire g708_n_spl_;
  wire g627_p_spl_;
  wire g709_n_spl_;
  wire g709_p_spl_;
  wire g711_p_spl_;
  wire g626_n_spl_;
  wire g711_n_spl_;
  wire g626_p_spl_;
  wire g712_n_spl_;
  wire g712_p_spl_;
  wire g714_p_spl_;
  wire g625_n_spl_;
  wire g714_n_spl_;
  wire g625_p_spl_;
  wire g715_n_spl_;
  wire g715_p_spl_;
  wire g717_p_spl_;
  wire g624_n_spl_;
  wire g717_n_spl_;
  wire g624_p_spl_;
  wire g718_n_spl_;
  wire g718_p_spl_;
  wire g720_n_spl_;
  wire g623_p_spl_;
  wire g721_p_spl_;
  wire G31_p_spl_;
  wire G31_p_spl_0;
  wire G31_p_spl_00;
  wire G31_p_spl_000;
  wire G31_p_spl_001;
  wire G31_p_spl_01;
  wire G31_p_spl_010;
  wire G31_p_spl_011;
  wire G31_p_spl_1;
  wire G31_p_spl_10;
  wire G31_p_spl_100;
  wire G31_p_spl_101;
  wire G31_p_spl_11;
  wire G31_p_spl_110;
  wire G31_p_spl_111;
  wire G31_n_spl_;
  wire G31_n_spl_0;
  wire G31_n_spl_00;
  wire G31_n_spl_000;
  wire G31_n_spl_001;
  wire G31_n_spl_01;
  wire G31_n_spl_010;
  wire G31_n_spl_011;
  wire G31_n_spl_1;
  wire G31_n_spl_10;
  wire G31_n_spl_100;
  wire G31_n_spl_101;
  wire G31_n_spl_11;
  wire G31_n_spl_110;
  wire G31_n_spl_111;
  wire G15_p_spl_;
  wire G15_p_spl_0;
  wire G15_p_spl_00;
  wire G15_p_spl_000;
  wire G15_p_spl_001;
  wire G15_p_spl_01;
  wire G15_p_spl_010;
  wire G15_p_spl_011;
  wire G15_p_spl_1;
  wire G15_p_spl_10;
  wire G15_p_spl_100;
  wire G15_p_spl_101;
  wire G15_p_spl_11;
  wire G15_p_spl_110;
  wire G15_p_spl_111;
  wire G15_n_spl_;
  wire G15_n_spl_0;
  wire G15_n_spl_00;
  wire G15_n_spl_000;
  wire G15_n_spl_001;
  wire G15_n_spl_01;
  wire G15_n_spl_010;
  wire G15_n_spl_011;
  wire G15_n_spl_1;
  wire G15_n_spl_10;
  wire G15_n_spl_100;
  wire G15_n_spl_101;
  wire G15_n_spl_11;
  wire G15_n_spl_110;
  wire G15_n_spl_111;
  wire g750_n_spl_;
  wire g749_p_spl_;
  wire g750_p_spl_;
  wire g749_n_spl_;
  wire g751_n_spl_;
  wire g751_p_spl_;
  wire g752_n_spl_;
  wire g752_n_spl_0;
  wire g752_p_spl_;
  wire g752_p_spl_0;
  wire g754_n_spl_;
  wire g754_p_spl_;
  wire g755_n_spl_;
  wire g755_p_spl_;
  wire g757_p_spl_;
  wire g748_n_spl_;
  wire g757_n_spl_;
  wire g748_p_spl_;
  wire g758_n_spl_;
  wire g758_p_spl_;
  wire g760_p_spl_;
  wire g747_n_spl_;
  wire g760_n_spl_;
  wire g747_p_spl_;
  wire g761_n_spl_;
  wire g761_p_spl_;
  wire g763_p_spl_;
  wire g746_n_spl_;
  wire g763_n_spl_;
  wire g746_p_spl_;
  wire g764_n_spl_;
  wire g764_p_spl_;
  wire g766_p_spl_;
  wire g745_n_spl_;
  wire g766_n_spl_;
  wire g745_p_spl_;
  wire g767_n_spl_;
  wire g767_p_spl_;
  wire g769_p_spl_;
  wire g744_n_spl_;
  wire g769_n_spl_;
  wire g744_p_spl_;
  wire g770_n_spl_;
  wire g770_p_spl_;
  wire g772_p_spl_;
  wire g743_n_spl_;
  wire g772_n_spl_;
  wire g743_p_spl_;
  wire g773_n_spl_;
  wire g773_p_spl_;
  wire g775_p_spl_;
  wire g742_n_spl_;
  wire g775_n_spl_;
  wire g742_p_spl_;
  wire g776_n_spl_;
  wire g776_p_spl_;
  wire g778_p_spl_;
  wire g741_n_spl_;
  wire g778_n_spl_;
  wire g741_p_spl_;
  wire g779_n_spl_;
  wire g779_p_spl_;
  wire g781_p_spl_;
  wire g740_n_spl_;
  wire g781_n_spl_;
  wire g740_p_spl_;
  wire g782_n_spl_;
  wire g782_p_spl_;
  wire g784_p_spl_;
  wire g739_n_spl_;
  wire g784_n_spl_;
  wire g739_p_spl_;
  wire g785_n_spl_;
  wire g785_p_spl_;
  wire g787_p_spl_;
  wire g738_n_spl_;
  wire g787_n_spl_;
  wire g738_p_spl_;
  wire g788_n_spl_;
  wire g788_p_spl_;
  wire g790_p_spl_;
  wire g737_n_spl_;
  wire g790_n_spl_;
  wire g737_p_spl_;
  wire g791_n_spl_;
  wire g791_p_spl_;
  wire g793_p_spl_;
  wire g736_n_spl_;
  wire g793_n_spl_;
  wire g736_p_spl_;
  wire g794_n_spl_;
  wire g794_p_spl_;
  wire g796_p_spl_;
  wire g735_n_spl_;
  wire g796_n_spl_;
  wire g735_p_spl_;
  wire g797_n_spl_;
  wire g797_p_spl_;
  wire g799_p_spl_;
  wire g734_n_spl_;
  wire g799_n_spl_;
  wire g734_p_spl_;
  wire g800_n_spl_;
  wire g800_p_spl_;
  wire g802_p_spl_;
  wire g733_n_spl_;
  wire g802_n_spl_;
  wire g733_p_spl_;
  wire g803_n_spl_;
  wire g803_p_spl_;
  wire g805_p_spl_;
  wire g732_n_spl_;
  wire g805_n_spl_;
  wire g732_p_spl_;
  wire g806_n_spl_;
  wire g806_p_spl_;
  wire g808_p_spl_;
  wire g731_n_spl_;
  wire g808_n_spl_;
  wire g731_p_spl_;
  wire g809_n_spl_;
  wire g809_p_spl_;
  wire g811_p_spl_;
  wire g730_n_spl_;
  wire g811_n_spl_;
  wire g730_p_spl_;
  wire g812_n_spl_;
  wire g812_p_spl_;
  wire g814_p_spl_;
  wire g729_n_spl_;
  wire g814_n_spl_;
  wire g729_p_spl_;
  wire g815_n_spl_;
  wire g815_p_spl_;
  wire g817_p_spl_;
  wire g728_n_spl_;
  wire g817_n_spl_;
  wire g728_p_spl_;
  wire g818_n_spl_;
  wire g818_p_spl_;
  wire g820_p_spl_;
  wire g727_n_spl_;
  wire g820_n_spl_;
  wire g727_p_spl_;
  wire g821_n_spl_;
  wire g821_p_spl_;
  wire g823_p_spl_;
  wire g726_n_spl_;
  wire g823_n_spl_;
  wire g726_p_spl_;
  wire g824_n_spl_;
  wire g824_p_spl_;
  wire g826_p_spl_;
  wire g725_n_spl_;
  wire g826_n_spl_;
  wire g725_p_spl_;
  wire g827_n_spl_;
  wire g827_p_spl_;
  wire g829_n_spl_;
  wire g724_p_spl_;
  wire g830_p_spl_;
  wire G32_p_spl_;
  wire G32_p_spl_0;
  wire G32_p_spl_00;
  wire G32_p_spl_000;
  wire G32_p_spl_001;
  wire G32_p_spl_01;
  wire G32_p_spl_010;
  wire G32_p_spl_011;
  wire G32_p_spl_1;
  wire G32_p_spl_10;
  wire G32_p_spl_100;
  wire G32_p_spl_101;
  wire G32_p_spl_11;
  wire G32_p_spl_110;
  wire G32_p_spl_111;
  wire G32_n_spl_;
  wire G32_n_spl_0;
  wire G32_n_spl_00;
  wire G32_n_spl_000;
  wire G32_n_spl_001;
  wire G32_n_spl_01;
  wire G32_n_spl_010;
  wire G32_n_spl_011;
  wire G32_n_spl_1;
  wire G32_n_spl_10;
  wire G32_n_spl_100;
  wire G32_n_spl_101;
  wire G32_n_spl_11;
  wire G32_n_spl_110;
  wire G32_n_spl_111;
  wire G16_p_spl_;
  wire G16_p_spl_0;
  wire G16_p_spl_00;
  wire G16_p_spl_000;
  wire G16_p_spl_001;
  wire G16_p_spl_01;
  wire G16_p_spl_010;
  wire G16_p_spl_011;
  wire G16_p_spl_1;
  wire G16_p_spl_10;
  wire G16_p_spl_100;
  wire G16_p_spl_101;
  wire G16_p_spl_11;
  wire G16_p_spl_110;
  wire G16_p_spl_111;
  wire G16_n_spl_;
  wire G16_n_spl_0;
  wire G16_n_spl_00;
  wire G16_n_spl_000;
  wire G16_n_spl_001;
  wire G16_n_spl_01;
  wire G16_n_spl_010;
  wire G16_n_spl_011;
  wire G16_n_spl_1;
  wire G16_n_spl_10;
  wire G16_n_spl_100;
  wire G16_n_spl_101;
  wire G16_n_spl_11;
  wire G16_n_spl_110;
  wire G16_n_spl_111;
  wire g861_n_spl_;
  wire g860_p_spl_;
  wire g861_p_spl_;
  wire g860_n_spl_;
  wire g862_n_spl_;
  wire g862_p_spl_;
  wire g863_n_spl_;
  wire g863_p_spl_;
  wire g865_n_spl_;
  wire g865_p_spl_;
  wire g866_n_spl_;
  wire g866_p_spl_;
  wire g868_p_spl_;
  wire g859_n_spl_;
  wire g868_n_spl_;
  wire g859_p_spl_;
  wire g869_n_spl_;
  wire g869_p_spl_;
  wire g871_p_spl_;
  wire g858_n_spl_;
  wire g871_n_spl_;
  wire g858_p_spl_;
  wire g872_n_spl_;
  wire g872_p_spl_;
  wire g874_p_spl_;
  wire g857_n_spl_;
  wire g874_n_spl_;
  wire g857_p_spl_;
  wire g875_n_spl_;
  wire g875_p_spl_;
  wire g877_p_spl_;
  wire g856_n_spl_;
  wire g877_n_spl_;
  wire g856_p_spl_;
  wire g878_n_spl_;
  wire g878_p_spl_;
  wire g880_p_spl_;
  wire g855_n_spl_;
  wire g880_n_spl_;
  wire g855_p_spl_;
  wire g881_n_spl_;
  wire g881_p_spl_;
  wire g883_p_spl_;
  wire g854_n_spl_;
  wire g883_n_spl_;
  wire g854_p_spl_;
  wire g884_n_spl_;
  wire g884_p_spl_;
  wire g886_p_spl_;
  wire g853_n_spl_;
  wire g886_n_spl_;
  wire g853_p_spl_;
  wire g887_n_spl_;
  wire g887_p_spl_;
  wire g889_p_spl_;
  wire g852_n_spl_;
  wire g889_n_spl_;
  wire g852_p_spl_;
  wire g890_n_spl_;
  wire g890_p_spl_;
  wire g892_p_spl_;
  wire g851_n_spl_;
  wire g892_n_spl_;
  wire g851_p_spl_;
  wire g893_n_spl_;
  wire g893_p_spl_;
  wire g895_p_spl_;
  wire g850_n_spl_;
  wire g895_n_spl_;
  wire g850_p_spl_;
  wire g896_n_spl_;
  wire g896_p_spl_;
  wire g898_p_spl_;
  wire g849_n_spl_;
  wire g898_n_spl_;
  wire g849_p_spl_;
  wire g899_n_spl_;
  wire g899_p_spl_;
  wire g901_p_spl_;
  wire g848_n_spl_;
  wire g901_n_spl_;
  wire g848_p_spl_;
  wire g902_n_spl_;
  wire g902_p_spl_;
  wire g904_p_spl_;
  wire g847_n_spl_;
  wire g904_n_spl_;
  wire g847_p_spl_;
  wire g905_n_spl_;
  wire g905_p_spl_;
  wire g907_p_spl_;
  wire g846_n_spl_;
  wire g907_n_spl_;
  wire g846_p_spl_;
  wire g908_n_spl_;
  wire g908_p_spl_;
  wire g910_p_spl_;
  wire g845_n_spl_;
  wire g910_n_spl_;
  wire g845_p_spl_;
  wire g911_n_spl_;
  wire g911_p_spl_;
  wire g913_p_spl_;
  wire g844_n_spl_;
  wire g913_n_spl_;
  wire g844_p_spl_;
  wire g914_n_spl_;
  wire g914_p_spl_;
  wire g916_p_spl_;
  wire g843_n_spl_;
  wire g916_n_spl_;
  wire g843_p_spl_;
  wire g917_n_spl_;
  wire g917_p_spl_;
  wire g919_p_spl_;
  wire g842_n_spl_;
  wire g919_n_spl_;
  wire g842_p_spl_;
  wire g920_n_spl_;
  wire g920_p_spl_;
  wire g922_p_spl_;
  wire g841_n_spl_;
  wire g922_n_spl_;
  wire g841_p_spl_;
  wire g923_n_spl_;
  wire g923_p_spl_;
  wire g925_p_spl_;
  wire g840_n_spl_;
  wire g925_n_spl_;
  wire g840_p_spl_;
  wire g926_n_spl_;
  wire g926_p_spl_;
  wire g928_p_spl_;
  wire g839_n_spl_;
  wire g928_n_spl_;
  wire g839_p_spl_;
  wire g929_n_spl_;
  wire g929_p_spl_;
  wire g931_p_spl_;
  wire g838_n_spl_;
  wire g931_n_spl_;
  wire g838_p_spl_;
  wire g932_n_spl_;
  wire g932_p_spl_;
  wire g934_p_spl_;
  wire g837_n_spl_;
  wire g934_n_spl_;
  wire g837_p_spl_;
  wire g935_n_spl_;
  wire g935_p_spl_;
  wire g937_p_spl_;
  wire g836_n_spl_;
  wire g937_n_spl_;
  wire g836_p_spl_;
  wire g938_n_spl_;
  wire g938_p_spl_;
  wire g940_p_spl_;
  wire g835_n_spl_;
  wire g940_n_spl_;
  wire g835_p_spl_;
  wire g941_n_spl_;
  wire g941_p_spl_;
  wire g943_p_spl_;
  wire g834_n_spl_;
  wire g943_n_spl_;
  wire g834_p_spl_;
  wire g944_n_spl_;
  wire g944_p_spl_;
  wire g946_n_spl_;
  wire g833_p_spl_;
  wire g947_p_spl_;
  wire g977_p_spl_;
  wire g977_n_spl_;
  wire g979_n_spl_;
  wire g978_p_spl_;
  wire g979_p_spl_;
  wire g978_n_spl_;
  wire g980_n_spl_;
  wire g980_p_spl_;
  wire g982_p_spl_;
  wire g976_n_spl_;
  wire g982_n_spl_;
  wire g976_p_spl_;
  wire g983_n_spl_;
  wire g983_p_spl_;
  wire g985_p_spl_;
  wire g975_n_spl_;
  wire g985_n_spl_;
  wire g975_p_spl_;
  wire g986_n_spl_;
  wire g986_p_spl_;
  wire g988_p_spl_;
  wire g974_n_spl_;
  wire g988_n_spl_;
  wire g974_p_spl_;
  wire g989_n_spl_;
  wire g989_p_spl_;
  wire g991_p_spl_;
  wire g973_n_spl_;
  wire g991_n_spl_;
  wire g973_p_spl_;
  wire g992_n_spl_;
  wire g992_p_spl_;
  wire g994_p_spl_;
  wire g972_n_spl_;
  wire g994_n_spl_;
  wire g972_p_spl_;
  wire g995_n_spl_;
  wire g995_p_spl_;
  wire g997_p_spl_;
  wire g971_n_spl_;
  wire g997_n_spl_;
  wire g971_p_spl_;
  wire g998_n_spl_;
  wire g998_p_spl_;
  wire g1000_p_spl_;
  wire g970_n_spl_;
  wire g1000_n_spl_;
  wire g970_p_spl_;
  wire g1001_n_spl_;
  wire g1001_p_spl_;
  wire g1003_p_spl_;
  wire g969_n_spl_;
  wire g1003_n_spl_;
  wire g969_p_spl_;
  wire g1004_n_spl_;
  wire g1004_p_spl_;
  wire g1006_p_spl_;
  wire g968_n_spl_;
  wire g1006_n_spl_;
  wire g968_p_spl_;
  wire g1007_n_spl_;
  wire g1007_p_spl_;
  wire g1009_p_spl_;
  wire g967_n_spl_;
  wire g1009_n_spl_;
  wire g967_p_spl_;
  wire g1010_n_spl_;
  wire g1010_p_spl_;
  wire g1012_p_spl_;
  wire g966_n_spl_;
  wire g1012_n_spl_;
  wire g966_p_spl_;
  wire g1013_n_spl_;
  wire g1013_p_spl_;
  wire g1015_p_spl_;
  wire g965_n_spl_;
  wire g1015_n_spl_;
  wire g965_p_spl_;
  wire g1016_n_spl_;
  wire g1016_p_spl_;
  wire g1018_p_spl_;
  wire g964_n_spl_;
  wire g1018_n_spl_;
  wire g964_p_spl_;
  wire g1019_n_spl_;
  wire g1019_p_spl_;
  wire g1021_p_spl_;
  wire g963_n_spl_;
  wire g1021_n_spl_;
  wire g963_p_spl_;
  wire g1022_n_spl_;
  wire g1022_p_spl_;
  wire g1024_p_spl_;
  wire g962_n_spl_;
  wire g1024_n_spl_;
  wire g962_p_spl_;
  wire g1025_n_spl_;
  wire g1025_p_spl_;
  wire g1027_p_spl_;
  wire g961_n_spl_;
  wire g1027_n_spl_;
  wire g961_p_spl_;
  wire g1028_n_spl_;
  wire g1028_p_spl_;
  wire g1030_p_spl_;
  wire g960_n_spl_;
  wire g1030_n_spl_;
  wire g960_p_spl_;
  wire g1031_n_spl_;
  wire g1031_p_spl_;
  wire g1033_p_spl_;
  wire g959_n_spl_;
  wire g1033_n_spl_;
  wire g959_p_spl_;
  wire g1034_n_spl_;
  wire g1034_p_spl_;
  wire g1036_p_spl_;
  wire g958_n_spl_;
  wire g1036_n_spl_;
  wire g958_p_spl_;
  wire g1037_n_spl_;
  wire g1037_p_spl_;
  wire g1039_p_spl_;
  wire g957_n_spl_;
  wire g1039_n_spl_;
  wire g957_p_spl_;
  wire g1040_n_spl_;
  wire g1040_p_spl_;
  wire g1042_p_spl_;
  wire g956_n_spl_;
  wire g1042_n_spl_;
  wire g956_p_spl_;
  wire g1043_n_spl_;
  wire g1043_p_spl_;
  wire g1045_p_spl_;
  wire g955_n_spl_;
  wire g1045_n_spl_;
  wire g955_p_spl_;
  wire g1046_n_spl_;
  wire g1046_p_spl_;
  wire g1048_p_spl_;
  wire g954_n_spl_;
  wire g1048_n_spl_;
  wire g954_p_spl_;
  wire g1049_n_spl_;
  wire g1049_p_spl_;
  wire g1051_p_spl_;
  wire g953_n_spl_;
  wire g1051_n_spl_;
  wire g953_p_spl_;
  wire g1052_n_spl_;
  wire g1052_p_spl_;
  wire g1054_p_spl_;
  wire g952_n_spl_;
  wire g1054_n_spl_;
  wire g952_p_spl_;
  wire g1055_n_spl_;
  wire g1055_p_spl_;
  wire g1057_p_spl_;
  wire g951_n_spl_;
  wire g1057_n_spl_;
  wire g951_p_spl_;
  wire g1058_n_spl_;
  wire g1058_p_spl_;
  wire g1060_n_spl_;
  wire g950_p_spl_;
  wire g1062_n_spl_;
  wire g1091_n_spl_;
  wire g1090_n_spl_;
  wire g1091_p_spl_;
  wire g1090_p_spl_;
  wire g1092_n_spl_;
  wire g1092_p_spl_;
  wire g1094_p_spl_;
  wire g1089_n_spl_;
  wire g1094_n_spl_;
  wire g1089_p_spl_;
  wire g1095_n_spl_;
  wire g1095_p_spl_;
  wire g1097_p_spl_;
  wire g1088_n_spl_;
  wire g1097_n_spl_;
  wire g1088_p_spl_;
  wire g1098_n_spl_;
  wire g1098_p_spl_;
  wire g1100_p_spl_;
  wire g1087_n_spl_;
  wire g1100_n_spl_;
  wire g1087_p_spl_;
  wire g1101_n_spl_;
  wire g1101_p_spl_;
  wire g1103_p_spl_;
  wire g1086_n_spl_;
  wire g1103_n_spl_;
  wire g1086_p_spl_;
  wire g1104_n_spl_;
  wire g1104_p_spl_;
  wire g1106_p_spl_;
  wire g1085_n_spl_;
  wire g1106_n_spl_;
  wire g1085_p_spl_;
  wire g1107_n_spl_;
  wire g1107_p_spl_;
  wire g1109_p_spl_;
  wire g1084_n_spl_;
  wire g1109_n_spl_;
  wire g1084_p_spl_;
  wire g1110_n_spl_;
  wire g1110_p_spl_;
  wire g1112_p_spl_;
  wire g1083_n_spl_;
  wire g1112_n_spl_;
  wire g1083_p_spl_;
  wire g1113_n_spl_;
  wire g1113_p_spl_;
  wire g1115_p_spl_;
  wire g1082_n_spl_;
  wire g1115_n_spl_;
  wire g1082_p_spl_;
  wire g1116_n_spl_;
  wire g1116_p_spl_;
  wire g1118_p_spl_;
  wire g1081_n_spl_;
  wire g1118_n_spl_;
  wire g1081_p_spl_;
  wire g1119_n_spl_;
  wire g1119_p_spl_;
  wire g1121_p_spl_;
  wire g1080_n_spl_;
  wire g1121_n_spl_;
  wire g1080_p_spl_;
  wire g1122_n_spl_;
  wire g1122_p_spl_;
  wire g1124_p_spl_;
  wire g1079_n_spl_;
  wire g1124_n_spl_;
  wire g1079_p_spl_;
  wire g1125_n_spl_;
  wire g1125_p_spl_;
  wire g1127_p_spl_;
  wire g1078_n_spl_;
  wire g1127_n_spl_;
  wire g1078_p_spl_;
  wire g1128_n_spl_;
  wire g1128_p_spl_;
  wire g1130_p_spl_;
  wire g1077_n_spl_;
  wire g1130_n_spl_;
  wire g1077_p_spl_;
  wire g1131_n_spl_;
  wire g1131_p_spl_;
  wire g1133_p_spl_;
  wire g1076_n_spl_;
  wire g1133_n_spl_;
  wire g1076_p_spl_;
  wire g1134_n_spl_;
  wire g1134_p_spl_;
  wire g1136_p_spl_;
  wire g1075_n_spl_;
  wire g1136_n_spl_;
  wire g1075_p_spl_;
  wire g1137_n_spl_;
  wire g1137_p_spl_;
  wire g1139_p_spl_;
  wire g1074_n_spl_;
  wire g1139_n_spl_;
  wire g1074_p_spl_;
  wire g1140_n_spl_;
  wire g1140_p_spl_;
  wire g1142_p_spl_;
  wire g1073_n_spl_;
  wire g1142_n_spl_;
  wire g1073_p_spl_;
  wire g1143_n_spl_;
  wire g1143_p_spl_;
  wire g1145_p_spl_;
  wire g1072_n_spl_;
  wire g1145_n_spl_;
  wire g1072_p_spl_;
  wire g1146_n_spl_;
  wire g1146_p_spl_;
  wire g1148_p_spl_;
  wire g1071_n_spl_;
  wire g1148_n_spl_;
  wire g1071_p_spl_;
  wire g1149_n_spl_;
  wire g1149_p_spl_;
  wire g1151_p_spl_;
  wire g1070_n_spl_;
  wire g1151_n_spl_;
  wire g1070_p_spl_;
  wire g1152_n_spl_;
  wire g1152_p_spl_;
  wire g1154_p_spl_;
  wire g1069_n_spl_;
  wire g1154_n_spl_;
  wire g1069_p_spl_;
  wire g1155_n_spl_;
  wire g1155_p_spl_;
  wire g1157_p_spl_;
  wire g1068_n_spl_;
  wire g1157_n_spl_;
  wire g1068_p_spl_;
  wire g1158_n_spl_;
  wire g1158_p_spl_;
  wire g1160_p_spl_;
  wire g1067_n_spl_;
  wire g1160_n_spl_;
  wire g1067_p_spl_;
  wire g1161_n_spl_;
  wire g1161_p_spl_;
  wire g1163_p_spl_;
  wire g1066_n_spl_;
  wire g1163_n_spl_;
  wire g1066_p_spl_;
  wire g1164_n_spl_;
  wire g1164_p_spl_;
  wire g1166_p_spl_;
  wire g1065_n_spl_;
  wire g1166_n_spl_;
  wire g1065_p_spl_;
  wire g1167_n_spl_;
  wire g1167_p_spl_;
  wire g1169_p_spl_;
  wire g1064_n_spl_;
  wire g1169_n_spl_;
  wire g1064_p_spl_;
  wire g1170_n_spl_;
  wire g1170_p_spl_;
  wire g1172_n_spl_;
  wire g1062_p_spl_;
  wire g1173_p_spl_;
  wire g1202_n_spl_;
  wire g1201_n_spl_;
  wire g1202_p_spl_;
  wire g1201_p_spl_;
  wire g1203_n_spl_;
  wire g1203_p_spl_;
  wire g1205_p_spl_;
  wire g1200_n_spl_;
  wire g1205_n_spl_;
  wire g1200_p_spl_;
  wire g1206_n_spl_;
  wire g1206_p_spl_;
  wire g1208_p_spl_;
  wire g1199_n_spl_;
  wire g1208_n_spl_;
  wire g1199_p_spl_;
  wire g1209_n_spl_;
  wire g1209_p_spl_;
  wire g1211_p_spl_;
  wire g1198_n_spl_;
  wire g1211_n_spl_;
  wire g1198_p_spl_;
  wire g1212_n_spl_;
  wire g1212_p_spl_;
  wire g1214_p_spl_;
  wire g1197_n_spl_;
  wire g1214_n_spl_;
  wire g1197_p_spl_;
  wire g1215_n_spl_;
  wire g1215_p_spl_;
  wire g1217_p_spl_;
  wire g1196_n_spl_;
  wire g1217_n_spl_;
  wire g1196_p_spl_;
  wire g1218_n_spl_;
  wire g1218_p_spl_;
  wire g1220_p_spl_;
  wire g1195_n_spl_;
  wire g1220_n_spl_;
  wire g1195_p_spl_;
  wire g1221_n_spl_;
  wire g1221_p_spl_;
  wire g1223_p_spl_;
  wire g1194_n_spl_;
  wire g1223_n_spl_;
  wire g1194_p_spl_;
  wire g1224_n_spl_;
  wire g1224_p_spl_;
  wire g1226_p_spl_;
  wire g1193_n_spl_;
  wire g1226_n_spl_;
  wire g1193_p_spl_;
  wire g1227_n_spl_;
  wire g1227_p_spl_;
  wire g1229_p_spl_;
  wire g1192_n_spl_;
  wire g1229_n_spl_;
  wire g1192_p_spl_;
  wire g1230_n_spl_;
  wire g1230_p_spl_;
  wire g1232_p_spl_;
  wire g1191_n_spl_;
  wire g1232_n_spl_;
  wire g1191_p_spl_;
  wire g1233_n_spl_;
  wire g1233_p_spl_;
  wire g1235_p_spl_;
  wire g1190_n_spl_;
  wire g1235_n_spl_;
  wire g1190_p_spl_;
  wire g1236_n_spl_;
  wire g1236_p_spl_;
  wire g1238_p_spl_;
  wire g1189_n_spl_;
  wire g1238_n_spl_;
  wire g1189_p_spl_;
  wire g1239_n_spl_;
  wire g1239_p_spl_;
  wire g1241_p_spl_;
  wire g1188_n_spl_;
  wire g1241_n_spl_;
  wire g1188_p_spl_;
  wire g1242_n_spl_;
  wire g1242_p_spl_;
  wire g1244_p_spl_;
  wire g1187_n_spl_;
  wire g1244_n_spl_;
  wire g1187_p_spl_;
  wire g1245_n_spl_;
  wire g1245_p_spl_;
  wire g1247_p_spl_;
  wire g1186_n_spl_;
  wire g1247_n_spl_;
  wire g1186_p_spl_;
  wire g1248_n_spl_;
  wire g1248_p_spl_;
  wire g1250_p_spl_;
  wire g1185_n_spl_;
  wire g1250_n_spl_;
  wire g1185_p_spl_;
  wire g1251_n_spl_;
  wire g1251_p_spl_;
  wire g1253_p_spl_;
  wire g1184_n_spl_;
  wire g1253_n_spl_;
  wire g1184_p_spl_;
  wire g1254_n_spl_;
  wire g1254_p_spl_;
  wire g1256_p_spl_;
  wire g1183_n_spl_;
  wire g1256_n_spl_;
  wire g1183_p_spl_;
  wire g1257_n_spl_;
  wire g1257_p_spl_;
  wire g1259_p_spl_;
  wire g1182_n_spl_;
  wire g1259_n_spl_;
  wire g1182_p_spl_;
  wire g1260_n_spl_;
  wire g1260_p_spl_;
  wire g1262_p_spl_;
  wire g1181_n_spl_;
  wire g1262_n_spl_;
  wire g1181_p_spl_;
  wire g1263_n_spl_;
  wire g1263_p_spl_;
  wire g1265_p_spl_;
  wire g1180_n_spl_;
  wire g1265_n_spl_;
  wire g1180_p_spl_;
  wire g1266_n_spl_;
  wire g1266_p_spl_;
  wire g1268_p_spl_;
  wire g1179_n_spl_;
  wire g1268_n_spl_;
  wire g1179_p_spl_;
  wire g1269_n_spl_;
  wire g1269_p_spl_;
  wire g1271_p_spl_;
  wire g1178_n_spl_;
  wire g1271_n_spl_;
  wire g1178_p_spl_;
  wire g1272_n_spl_;
  wire g1272_p_spl_;
  wire g1274_p_spl_;
  wire g1177_n_spl_;
  wire g1274_n_spl_;
  wire g1177_p_spl_;
  wire g1275_n_spl_;
  wire g1275_p_spl_;
  wire g1277_n_spl_;
  wire g1176_p_spl_;
  wire g1278_p_spl_;
  wire g1305_n_spl_;
  wire g1304_n_spl_;
  wire g1305_p_spl_;
  wire g1304_p_spl_;
  wire g1306_n_spl_;
  wire g1306_p_spl_;
  wire g1308_p_spl_;
  wire g1303_n_spl_;
  wire g1308_n_spl_;
  wire g1303_p_spl_;
  wire g1309_n_spl_;
  wire g1309_p_spl_;
  wire g1311_p_spl_;
  wire g1302_n_spl_;
  wire g1311_n_spl_;
  wire g1302_p_spl_;
  wire g1312_n_spl_;
  wire g1312_p_spl_;
  wire g1314_p_spl_;
  wire g1301_n_spl_;
  wire g1314_n_spl_;
  wire g1301_p_spl_;
  wire g1315_n_spl_;
  wire g1315_p_spl_;
  wire g1317_p_spl_;
  wire g1300_n_spl_;
  wire g1317_n_spl_;
  wire g1300_p_spl_;
  wire g1318_n_spl_;
  wire g1318_p_spl_;
  wire g1320_p_spl_;
  wire g1299_n_spl_;
  wire g1320_n_spl_;
  wire g1299_p_spl_;
  wire g1321_n_spl_;
  wire g1321_p_spl_;
  wire g1323_p_spl_;
  wire g1298_n_spl_;
  wire g1323_n_spl_;
  wire g1298_p_spl_;
  wire g1324_n_spl_;
  wire g1324_p_spl_;
  wire g1326_p_spl_;
  wire g1297_n_spl_;
  wire g1326_n_spl_;
  wire g1297_p_spl_;
  wire g1327_n_spl_;
  wire g1327_p_spl_;
  wire g1329_p_spl_;
  wire g1296_n_spl_;
  wire g1329_n_spl_;
  wire g1296_p_spl_;
  wire g1330_n_spl_;
  wire g1330_p_spl_;
  wire g1332_p_spl_;
  wire g1295_n_spl_;
  wire g1332_n_spl_;
  wire g1295_p_spl_;
  wire g1333_n_spl_;
  wire g1333_p_spl_;
  wire g1335_p_spl_;
  wire g1294_n_spl_;
  wire g1335_n_spl_;
  wire g1294_p_spl_;
  wire g1336_n_spl_;
  wire g1336_p_spl_;
  wire g1338_p_spl_;
  wire g1293_n_spl_;
  wire g1338_n_spl_;
  wire g1293_p_spl_;
  wire g1339_n_spl_;
  wire g1339_p_spl_;
  wire g1341_p_spl_;
  wire g1292_n_spl_;
  wire g1341_n_spl_;
  wire g1292_p_spl_;
  wire g1342_n_spl_;
  wire g1342_p_spl_;
  wire g1344_p_spl_;
  wire g1291_n_spl_;
  wire g1344_n_spl_;
  wire g1291_p_spl_;
  wire g1345_n_spl_;
  wire g1345_p_spl_;
  wire g1347_p_spl_;
  wire g1290_n_spl_;
  wire g1347_n_spl_;
  wire g1290_p_spl_;
  wire g1348_n_spl_;
  wire g1348_p_spl_;
  wire g1350_p_spl_;
  wire g1289_n_spl_;
  wire g1350_n_spl_;
  wire g1289_p_spl_;
  wire g1351_n_spl_;
  wire g1351_p_spl_;
  wire g1353_p_spl_;
  wire g1288_n_spl_;
  wire g1353_n_spl_;
  wire g1288_p_spl_;
  wire g1354_n_spl_;
  wire g1354_p_spl_;
  wire g1356_p_spl_;
  wire g1287_n_spl_;
  wire g1356_n_spl_;
  wire g1287_p_spl_;
  wire g1357_n_spl_;
  wire g1357_p_spl_;
  wire g1359_p_spl_;
  wire g1286_n_spl_;
  wire g1359_n_spl_;
  wire g1286_p_spl_;
  wire g1360_n_spl_;
  wire g1360_p_spl_;
  wire g1362_p_spl_;
  wire g1285_n_spl_;
  wire g1362_n_spl_;
  wire g1285_p_spl_;
  wire g1363_n_spl_;
  wire g1363_p_spl_;
  wire g1365_p_spl_;
  wire g1284_n_spl_;
  wire g1365_n_spl_;
  wire g1284_p_spl_;
  wire g1366_n_spl_;
  wire g1366_p_spl_;
  wire g1368_p_spl_;
  wire g1283_n_spl_;
  wire g1368_n_spl_;
  wire g1283_p_spl_;
  wire g1369_n_spl_;
  wire g1369_p_spl_;
  wire g1371_p_spl_;
  wire g1282_n_spl_;
  wire g1371_n_spl_;
  wire g1282_p_spl_;
  wire g1372_n_spl_;
  wire g1372_p_spl_;
  wire g1374_n_spl_;
  wire g1281_p_spl_;
  wire g1375_p_spl_;
  wire g1400_n_spl_;
  wire g1399_n_spl_;
  wire g1400_p_spl_;
  wire g1399_p_spl_;
  wire g1401_n_spl_;
  wire g1401_p_spl_;
  wire g1403_p_spl_;
  wire g1398_n_spl_;
  wire g1403_n_spl_;
  wire g1398_p_spl_;
  wire g1404_n_spl_;
  wire g1404_p_spl_;
  wire g1406_p_spl_;
  wire g1397_n_spl_;
  wire g1406_n_spl_;
  wire g1397_p_spl_;
  wire g1407_n_spl_;
  wire g1407_p_spl_;
  wire g1409_p_spl_;
  wire g1396_n_spl_;
  wire g1409_n_spl_;
  wire g1396_p_spl_;
  wire g1410_n_spl_;
  wire g1410_p_spl_;
  wire g1412_p_spl_;
  wire g1395_n_spl_;
  wire g1412_n_spl_;
  wire g1395_p_spl_;
  wire g1413_n_spl_;
  wire g1413_p_spl_;
  wire g1415_p_spl_;
  wire g1394_n_spl_;
  wire g1415_n_spl_;
  wire g1394_p_spl_;
  wire g1416_n_spl_;
  wire g1416_p_spl_;
  wire g1418_p_spl_;
  wire g1393_n_spl_;
  wire g1418_n_spl_;
  wire g1393_p_spl_;
  wire g1419_n_spl_;
  wire g1419_p_spl_;
  wire g1421_p_spl_;
  wire g1392_n_spl_;
  wire g1421_n_spl_;
  wire g1392_p_spl_;
  wire g1422_n_spl_;
  wire g1422_p_spl_;
  wire g1424_p_spl_;
  wire g1391_n_spl_;
  wire g1424_n_spl_;
  wire g1391_p_spl_;
  wire g1425_n_spl_;
  wire g1425_p_spl_;
  wire g1427_p_spl_;
  wire g1390_n_spl_;
  wire g1427_n_spl_;
  wire g1390_p_spl_;
  wire g1428_n_spl_;
  wire g1428_p_spl_;
  wire g1430_p_spl_;
  wire g1389_n_spl_;
  wire g1430_n_spl_;
  wire g1389_p_spl_;
  wire g1431_n_spl_;
  wire g1431_p_spl_;
  wire g1433_p_spl_;
  wire g1388_n_spl_;
  wire g1433_n_spl_;
  wire g1388_p_spl_;
  wire g1434_n_spl_;
  wire g1434_p_spl_;
  wire g1436_p_spl_;
  wire g1387_n_spl_;
  wire g1436_n_spl_;
  wire g1387_p_spl_;
  wire g1437_n_spl_;
  wire g1437_p_spl_;
  wire g1439_p_spl_;
  wire g1386_n_spl_;
  wire g1439_n_spl_;
  wire g1386_p_spl_;
  wire g1440_n_spl_;
  wire g1440_p_spl_;
  wire g1442_p_spl_;
  wire g1385_n_spl_;
  wire g1442_n_spl_;
  wire g1385_p_spl_;
  wire g1443_n_spl_;
  wire g1443_p_spl_;
  wire g1445_p_spl_;
  wire g1384_n_spl_;
  wire g1445_n_spl_;
  wire g1384_p_spl_;
  wire g1446_n_spl_;
  wire g1446_p_spl_;
  wire g1448_p_spl_;
  wire g1383_n_spl_;
  wire g1448_n_spl_;
  wire g1383_p_spl_;
  wire g1449_n_spl_;
  wire g1449_p_spl_;
  wire g1451_p_spl_;
  wire g1382_n_spl_;
  wire g1451_n_spl_;
  wire g1382_p_spl_;
  wire g1452_n_spl_;
  wire g1452_p_spl_;
  wire g1454_p_spl_;
  wire g1381_n_spl_;
  wire g1454_n_spl_;
  wire g1381_p_spl_;
  wire g1455_n_spl_;
  wire g1455_p_spl_;
  wire g1457_p_spl_;
  wire g1380_n_spl_;
  wire g1457_n_spl_;
  wire g1380_p_spl_;
  wire g1458_n_spl_;
  wire g1458_p_spl_;
  wire g1460_p_spl_;
  wire g1379_n_spl_;
  wire g1460_n_spl_;
  wire g1379_p_spl_;
  wire g1461_n_spl_;
  wire g1461_p_spl_;
  wire g1463_n_spl_;
  wire g1378_p_spl_;
  wire g1464_p_spl_;
  wire g1487_n_spl_;
  wire g1486_n_spl_;
  wire g1487_p_spl_;
  wire g1486_p_spl_;
  wire g1488_n_spl_;
  wire g1488_p_spl_;
  wire g1490_p_spl_;
  wire g1485_n_spl_;
  wire g1490_n_spl_;
  wire g1485_p_spl_;
  wire g1491_n_spl_;
  wire g1491_p_spl_;
  wire g1493_p_spl_;
  wire g1484_n_spl_;
  wire g1493_n_spl_;
  wire g1484_p_spl_;
  wire g1494_n_spl_;
  wire g1494_p_spl_;
  wire g1496_p_spl_;
  wire g1483_n_spl_;
  wire g1496_n_spl_;
  wire g1483_p_spl_;
  wire g1497_n_spl_;
  wire g1497_p_spl_;
  wire g1499_p_spl_;
  wire g1482_n_spl_;
  wire g1499_n_spl_;
  wire g1482_p_spl_;
  wire g1500_n_spl_;
  wire g1500_p_spl_;
  wire g1502_p_spl_;
  wire g1481_n_spl_;
  wire g1502_n_spl_;
  wire g1481_p_spl_;
  wire g1503_n_spl_;
  wire g1503_p_spl_;
  wire g1505_p_spl_;
  wire g1480_n_spl_;
  wire g1505_n_spl_;
  wire g1480_p_spl_;
  wire g1506_n_spl_;
  wire g1506_p_spl_;
  wire g1508_p_spl_;
  wire g1479_n_spl_;
  wire g1508_n_spl_;
  wire g1479_p_spl_;
  wire g1509_n_spl_;
  wire g1509_p_spl_;
  wire g1511_p_spl_;
  wire g1478_n_spl_;
  wire g1511_n_spl_;
  wire g1478_p_spl_;
  wire g1512_n_spl_;
  wire g1512_p_spl_;
  wire g1514_p_spl_;
  wire g1477_n_spl_;
  wire g1514_n_spl_;
  wire g1477_p_spl_;
  wire g1515_n_spl_;
  wire g1515_p_spl_;
  wire g1517_p_spl_;
  wire g1476_n_spl_;
  wire g1517_n_spl_;
  wire g1476_p_spl_;
  wire g1518_n_spl_;
  wire g1518_p_spl_;
  wire g1520_p_spl_;
  wire g1475_n_spl_;
  wire g1520_n_spl_;
  wire g1475_p_spl_;
  wire g1521_n_spl_;
  wire g1521_p_spl_;
  wire g1523_p_spl_;
  wire g1474_n_spl_;
  wire g1523_n_spl_;
  wire g1474_p_spl_;
  wire g1524_n_spl_;
  wire g1524_p_spl_;
  wire g1526_p_spl_;
  wire g1473_n_spl_;
  wire g1526_n_spl_;
  wire g1473_p_spl_;
  wire g1527_n_spl_;
  wire g1527_p_spl_;
  wire g1529_p_spl_;
  wire g1472_n_spl_;
  wire g1529_n_spl_;
  wire g1472_p_spl_;
  wire g1530_n_spl_;
  wire g1530_p_spl_;
  wire g1532_p_spl_;
  wire g1471_n_spl_;
  wire g1532_n_spl_;
  wire g1471_p_spl_;
  wire g1533_n_spl_;
  wire g1533_p_spl_;
  wire g1535_p_spl_;
  wire g1470_n_spl_;
  wire g1535_n_spl_;
  wire g1470_p_spl_;
  wire g1536_n_spl_;
  wire g1536_p_spl_;
  wire g1538_p_spl_;
  wire g1469_n_spl_;
  wire g1538_n_spl_;
  wire g1469_p_spl_;
  wire g1539_n_spl_;
  wire g1539_p_spl_;
  wire g1541_p_spl_;
  wire g1468_n_spl_;
  wire g1541_n_spl_;
  wire g1468_p_spl_;
  wire g1542_n_spl_;
  wire g1542_p_spl_;
  wire g1544_n_spl_;
  wire g1467_p_spl_;
  wire g1545_p_spl_;
  wire g1566_n_spl_;
  wire g1565_n_spl_;
  wire g1566_p_spl_;
  wire g1565_p_spl_;
  wire g1567_n_spl_;
  wire g1567_p_spl_;
  wire g1569_p_spl_;
  wire g1564_n_spl_;
  wire g1569_n_spl_;
  wire g1564_p_spl_;
  wire g1570_n_spl_;
  wire g1570_p_spl_;
  wire g1572_p_spl_;
  wire g1563_n_spl_;
  wire g1572_n_spl_;
  wire g1563_p_spl_;
  wire g1573_n_spl_;
  wire g1573_p_spl_;
  wire g1575_p_spl_;
  wire g1562_n_spl_;
  wire g1575_n_spl_;
  wire g1562_p_spl_;
  wire g1576_n_spl_;
  wire g1576_p_spl_;
  wire g1578_p_spl_;
  wire g1561_n_spl_;
  wire g1578_n_spl_;
  wire g1561_p_spl_;
  wire g1579_n_spl_;
  wire g1579_p_spl_;
  wire g1581_p_spl_;
  wire g1560_n_spl_;
  wire g1581_n_spl_;
  wire g1560_p_spl_;
  wire g1582_n_spl_;
  wire g1582_p_spl_;
  wire g1584_p_spl_;
  wire g1559_n_spl_;
  wire g1584_n_spl_;
  wire g1559_p_spl_;
  wire g1585_n_spl_;
  wire g1585_p_spl_;
  wire g1587_p_spl_;
  wire g1558_n_spl_;
  wire g1587_n_spl_;
  wire g1558_p_spl_;
  wire g1588_n_spl_;
  wire g1588_p_spl_;
  wire g1590_p_spl_;
  wire g1557_n_spl_;
  wire g1590_n_spl_;
  wire g1557_p_spl_;
  wire g1591_n_spl_;
  wire g1591_p_spl_;
  wire g1593_p_spl_;
  wire g1556_n_spl_;
  wire g1593_n_spl_;
  wire g1556_p_spl_;
  wire g1594_n_spl_;
  wire g1594_p_spl_;
  wire g1596_p_spl_;
  wire g1555_n_spl_;
  wire g1596_n_spl_;
  wire g1555_p_spl_;
  wire g1597_n_spl_;
  wire g1597_p_spl_;
  wire g1599_p_spl_;
  wire g1554_n_spl_;
  wire g1599_n_spl_;
  wire g1554_p_spl_;
  wire g1600_n_spl_;
  wire g1600_p_spl_;
  wire g1602_p_spl_;
  wire g1553_n_spl_;
  wire g1602_n_spl_;
  wire g1553_p_spl_;
  wire g1603_n_spl_;
  wire g1603_p_spl_;
  wire g1605_p_spl_;
  wire g1552_n_spl_;
  wire g1605_n_spl_;
  wire g1552_p_spl_;
  wire g1606_n_spl_;
  wire g1606_p_spl_;
  wire g1608_p_spl_;
  wire g1551_n_spl_;
  wire g1608_n_spl_;
  wire g1551_p_spl_;
  wire g1609_n_spl_;
  wire g1609_p_spl_;
  wire g1611_p_spl_;
  wire g1550_n_spl_;
  wire g1611_n_spl_;
  wire g1550_p_spl_;
  wire g1612_n_spl_;
  wire g1612_p_spl_;
  wire g1614_p_spl_;
  wire g1549_n_spl_;
  wire g1614_n_spl_;
  wire g1549_p_spl_;
  wire g1615_n_spl_;
  wire g1615_p_spl_;
  wire g1617_n_spl_;
  wire g1548_p_spl_;
  wire g1618_p_spl_;
  wire g1637_n_spl_;
  wire g1636_n_spl_;
  wire g1637_p_spl_;
  wire g1636_p_spl_;
  wire g1638_n_spl_;
  wire g1638_p_spl_;
  wire g1640_p_spl_;
  wire g1635_n_spl_;
  wire g1640_n_spl_;
  wire g1635_p_spl_;
  wire g1641_n_spl_;
  wire g1641_p_spl_;
  wire g1643_p_spl_;
  wire g1634_n_spl_;
  wire g1643_n_spl_;
  wire g1634_p_spl_;
  wire g1644_n_spl_;
  wire g1644_p_spl_;
  wire g1646_p_spl_;
  wire g1633_n_spl_;
  wire g1646_n_spl_;
  wire g1633_p_spl_;
  wire g1647_n_spl_;
  wire g1647_p_spl_;
  wire g1649_p_spl_;
  wire g1632_n_spl_;
  wire g1649_n_spl_;
  wire g1632_p_spl_;
  wire g1650_n_spl_;
  wire g1650_p_spl_;
  wire g1652_p_spl_;
  wire g1631_n_spl_;
  wire g1652_n_spl_;
  wire g1631_p_spl_;
  wire g1653_n_spl_;
  wire g1653_p_spl_;
  wire g1655_p_spl_;
  wire g1630_n_spl_;
  wire g1655_n_spl_;
  wire g1630_p_spl_;
  wire g1656_n_spl_;
  wire g1656_p_spl_;
  wire g1658_p_spl_;
  wire g1629_n_spl_;
  wire g1658_n_spl_;
  wire g1629_p_spl_;
  wire g1659_n_spl_;
  wire g1659_p_spl_;
  wire g1661_p_spl_;
  wire g1628_n_spl_;
  wire g1661_n_spl_;
  wire g1628_p_spl_;
  wire g1662_n_spl_;
  wire g1662_p_spl_;
  wire g1664_p_spl_;
  wire g1627_n_spl_;
  wire g1664_n_spl_;
  wire g1627_p_spl_;
  wire g1665_n_spl_;
  wire g1665_p_spl_;
  wire g1667_p_spl_;
  wire g1626_n_spl_;
  wire g1667_n_spl_;
  wire g1626_p_spl_;
  wire g1668_n_spl_;
  wire g1668_p_spl_;
  wire g1670_p_spl_;
  wire g1625_n_spl_;
  wire g1670_n_spl_;
  wire g1625_p_spl_;
  wire g1671_n_spl_;
  wire g1671_p_spl_;
  wire g1673_p_spl_;
  wire g1624_n_spl_;
  wire g1673_n_spl_;
  wire g1624_p_spl_;
  wire g1674_n_spl_;
  wire g1674_p_spl_;
  wire g1676_p_spl_;
  wire g1623_n_spl_;
  wire g1676_n_spl_;
  wire g1623_p_spl_;
  wire g1677_n_spl_;
  wire g1677_p_spl_;
  wire g1679_p_spl_;
  wire g1622_n_spl_;
  wire g1679_n_spl_;
  wire g1622_p_spl_;
  wire g1680_n_spl_;
  wire g1680_p_spl_;
  wire g1682_n_spl_;
  wire g1621_p_spl_;
  wire g1683_p_spl_;
  wire g1700_n_spl_;
  wire g1699_n_spl_;
  wire g1700_p_spl_;
  wire g1699_p_spl_;
  wire g1701_n_spl_;
  wire g1701_p_spl_;
  wire g1703_p_spl_;
  wire g1698_n_spl_;
  wire g1703_n_spl_;
  wire g1698_p_spl_;
  wire g1704_n_spl_;
  wire g1704_p_spl_;
  wire g1706_p_spl_;
  wire g1697_n_spl_;
  wire g1706_n_spl_;
  wire g1697_p_spl_;
  wire g1707_n_spl_;
  wire g1707_p_spl_;
  wire g1709_p_spl_;
  wire g1696_n_spl_;
  wire g1709_n_spl_;
  wire g1696_p_spl_;
  wire g1710_n_spl_;
  wire g1710_p_spl_;
  wire g1712_p_spl_;
  wire g1695_n_spl_;
  wire g1712_n_spl_;
  wire g1695_p_spl_;
  wire g1713_n_spl_;
  wire g1713_p_spl_;
  wire g1715_p_spl_;
  wire g1694_n_spl_;
  wire g1715_n_spl_;
  wire g1694_p_spl_;
  wire g1716_n_spl_;
  wire g1716_p_spl_;
  wire g1718_p_spl_;
  wire g1693_n_spl_;
  wire g1718_n_spl_;
  wire g1693_p_spl_;
  wire g1719_n_spl_;
  wire g1719_p_spl_;
  wire g1721_p_spl_;
  wire g1692_n_spl_;
  wire g1721_n_spl_;
  wire g1692_p_spl_;
  wire g1722_n_spl_;
  wire g1722_p_spl_;
  wire g1724_p_spl_;
  wire g1691_n_spl_;
  wire g1724_n_spl_;
  wire g1691_p_spl_;
  wire g1725_n_spl_;
  wire g1725_p_spl_;
  wire g1727_p_spl_;
  wire g1690_n_spl_;
  wire g1727_n_spl_;
  wire g1690_p_spl_;
  wire g1728_n_spl_;
  wire g1728_p_spl_;
  wire g1730_p_spl_;
  wire g1689_n_spl_;
  wire g1730_n_spl_;
  wire g1689_p_spl_;
  wire g1731_n_spl_;
  wire g1731_p_spl_;
  wire g1733_p_spl_;
  wire g1688_n_spl_;
  wire g1733_n_spl_;
  wire g1688_p_spl_;
  wire g1734_n_spl_;
  wire g1734_p_spl_;
  wire g1736_p_spl_;
  wire g1687_n_spl_;
  wire g1736_n_spl_;
  wire g1687_p_spl_;
  wire g1737_n_spl_;
  wire g1737_p_spl_;
  wire g1739_n_spl_;
  wire g1686_p_spl_;
  wire g1740_p_spl_;
  wire g1755_n_spl_;
  wire g1754_n_spl_;
  wire g1755_p_spl_;
  wire g1754_p_spl_;
  wire g1756_n_spl_;
  wire g1756_p_spl_;
  wire g1758_p_spl_;
  wire g1753_n_spl_;
  wire g1758_n_spl_;
  wire g1753_p_spl_;
  wire g1759_n_spl_;
  wire g1759_p_spl_;
  wire g1761_p_spl_;
  wire g1752_n_spl_;
  wire g1761_n_spl_;
  wire g1752_p_spl_;
  wire g1762_n_spl_;
  wire g1762_p_spl_;
  wire g1764_p_spl_;
  wire g1751_n_spl_;
  wire g1764_n_spl_;
  wire g1751_p_spl_;
  wire g1765_n_spl_;
  wire g1765_p_spl_;
  wire g1767_p_spl_;
  wire g1750_n_spl_;
  wire g1767_n_spl_;
  wire g1750_p_spl_;
  wire g1768_n_spl_;
  wire g1768_p_spl_;
  wire g1770_p_spl_;
  wire g1749_n_spl_;
  wire g1770_n_spl_;
  wire g1749_p_spl_;
  wire g1771_n_spl_;
  wire g1771_p_spl_;
  wire g1773_p_spl_;
  wire g1748_n_spl_;
  wire g1773_n_spl_;
  wire g1748_p_spl_;
  wire g1774_n_spl_;
  wire g1774_p_spl_;
  wire g1776_p_spl_;
  wire g1747_n_spl_;
  wire g1776_n_spl_;
  wire g1747_p_spl_;
  wire g1777_n_spl_;
  wire g1777_p_spl_;
  wire g1779_p_spl_;
  wire g1746_n_spl_;
  wire g1779_n_spl_;
  wire g1746_p_spl_;
  wire g1780_n_spl_;
  wire g1780_p_spl_;
  wire g1782_p_spl_;
  wire g1745_n_spl_;
  wire g1782_n_spl_;
  wire g1745_p_spl_;
  wire g1783_n_spl_;
  wire g1783_p_spl_;
  wire g1785_p_spl_;
  wire g1744_n_spl_;
  wire g1785_n_spl_;
  wire g1744_p_spl_;
  wire g1786_n_spl_;
  wire g1786_p_spl_;
  wire g1788_n_spl_;
  wire g1743_p_spl_;
  wire g1789_p_spl_;
  wire g1802_n_spl_;
  wire g1801_n_spl_;
  wire g1802_p_spl_;
  wire g1801_p_spl_;
  wire g1803_n_spl_;
  wire g1803_p_spl_;
  wire g1805_p_spl_;
  wire g1800_n_spl_;
  wire g1805_n_spl_;
  wire g1800_p_spl_;
  wire g1806_n_spl_;
  wire g1806_p_spl_;
  wire g1808_p_spl_;
  wire g1799_n_spl_;
  wire g1808_n_spl_;
  wire g1799_p_spl_;
  wire g1809_n_spl_;
  wire g1809_p_spl_;
  wire g1811_p_spl_;
  wire g1798_n_spl_;
  wire g1811_n_spl_;
  wire g1798_p_spl_;
  wire g1812_n_spl_;
  wire g1812_p_spl_;
  wire g1814_p_spl_;
  wire g1797_n_spl_;
  wire g1814_n_spl_;
  wire g1797_p_spl_;
  wire g1815_n_spl_;
  wire g1815_p_spl_;
  wire g1817_p_spl_;
  wire g1796_n_spl_;
  wire g1817_n_spl_;
  wire g1796_p_spl_;
  wire g1818_n_spl_;
  wire g1818_p_spl_;
  wire g1820_p_spl_;
  wire g1795_n_spl_;
  wire g1820_n_spl_;
  wire g1795_p_spl_;
  wire g1821_n_spl_;
  wire g1821_p_spl_;
  wire g1823_p_spl_;
  wire g1794_n_spl_;
  wire g1823_n_spl_;
  wire g1794_p_spl_;
  wire g1824_n_spl_;
  wire g1824_p_spl_;
  wire g1826_p_spl_;
  wire g1793_n_spl_;
  wire g1826_n_spl_;
  wire g1793_p_spl_;
  wire g1827_n_spl_;
  wire g1827_p_spl_;
  wire g1829_n_spl_;
  wire g1792_p_spl_;
  wire g1830_p_spl_;
  wire g1841_n_spl_;
  wire g1840_n_spl_;
  wire g1841_p_spl_;
  wire g1840_p_spl_;
  wire g1842_n_spl_;
  wire g1842_p_spl_;
  wire g1844_p_spl_;
  wire g1839_n_spl_;
  wire g1844_n_spl_;
  wire g1839_p_spl_;
  wire g1845_n_spl_;
  wire g1845_p_spl_;
  wire g1847_p_spl_;
  wire g1838_n_spl_;
  wire g1847_n_spl_;
  wire g1838_p_spl_;
  wire g1848_n_spl_;
  wire g1848_p_spl_;
  wire g1850_p_spl_;
  wire g1837_n_spl_;
  wire g1850_n_spl_;
  wire g1837_p_spl_;
  wire g1851_n_spl_;
  wire g1851_p_spl_;
  wire g1853_p_spl_;
  wire g1836_n_spl_;
  wire g1853_n_spl_;
  wire g1836_p_spl_;
  wire g1854_n_spl_;
  wire g1854_p_spl_;
  wire g1856_p_spl_;
  wire g1835_n_spl_;
  wire g1856_n_spl_;
  wire g1835_p_spl_;
  wire g1857_n_spl_;
  wire g1857_p_spl_;
  wire g1859_p_spl_;
  wire g1834_n_spl_;
  wire g1859_n_spl_;
  wire g1834_p_spl_;
  wire g1860_n_spl_;
  wire g1860_p_spl_;
  wire g1862_n_spl_;
  wire g1833_p_spl_;
  wire g1863_p_spl_;
  wire g1872_n_spl_;
  wire g1871_n_spl_;
  wire g1872_p_spl_;
  wire g1871_p_spl_;
  wire g1873_n_spl_;
  wire g1873_p_spl_;
  wire g1875_p_spl_;
  wire g1870_n_spl_;
  wire g1875_n_spl_;
  wire g1870_p_spl_;
  wire g1876_n_spl_;
  wire g1876_p_spl_;
  wire g1878_p_spl_;
  wire g1869_n_spl_;
  wire g1878_n_spl_;
  wire g1869_p_spl_;
  wire g1879_n_spl_;
  wire g1879_p_spl_;
  wire g1881_p_spl_;
  wire g1868_n_spl_;
  wire g1881_n_spl_;
  wire g1868_p_spl_;
  wire g1882_n_spl_;
  wire g1882_p_spl_;
  wire g1884_p_spl_;
  wire g1867_n_spl_;
  wire g1884_n_spl_;
  wire g1867_p_spl_;
  wire g1885_n_spl_;
  wire g1885_p_spl_;
  wire g1887_n_spl_;
  wire g1866_p_spl_;
  wire g1888_p_spl_;
  wire g1895_n_spl_;
  wire g1894_n_spl_;
  wire g1895_p_spl_;
  wire g1894_p_spl_;
  wire g1896_n_spl_;
  wire g1896_p_spl_;
  wire g1898_p_spl_;
  wire g1893_n_spl_;
  wire g1898_n_spl_;
  wire g1893_p_spl_;
  wire g1899_n_spl_;
  wire g1899_p_spl_;
  wire g1901_p_spl_;
  wire g1892_n_spl_;
  wire g1901_n_spl_;
  wire g1892_p_spl_;
  wire g1902_n_spl_;
  wire g1902_p_spl_;
  wire g1904_n_spl_;
  wire g1891_p_spl_;
  wire g1905_p_spl_;
  wire g1909_n_spl_;
  wire g1908_n_spl_;
  wire g1909_p_spl_;
  wire g1908_p_spl_;
  wire g1910_n_spl_;
  wire g1914_n_spl_;

  buf

  (
    G1_p,
    G1
  );


  not

  (
    G1_n,
    G1
  );


  buf

  (
    G2_p,
    G2
  );


  not

  (
    G2_n,
    G2
  );


  buf

  (
    G3_p,
    G3
  );


  not

  (
    G3_n,
    G3
  );


  buf

  (
    G4_p,
    G4
  );


  not

  (
    G4_n,
    G4
  );


  buf

  (
    G5_p,
    G5
  );


  not

  (
    G5_n,
    G5
  );


  buf

  (
    G6_p,
    G6
  );


  not

  (
    G6_n,
    G6
  );


  buf

  (
    G7_p,
    G7
  );


  not

  (
    G7_n,
    G7
  );


  buf

  (
    G8_p,
    G8
  );


  not

  (
    G8_n,
    G8
  );


  buf

  (
    G9_p,
    G9
  );


  not

  (
    G9_n,
    G9
  );


  buf

  (
    G10_p,
    G10
  );


  not

  (
    G10_n,
    G10
  );


  buf

  (
    G11_p,
    G11
  );


  not

  (
    G11_n,
    G11
  );


  buf

  (
    G12_p,
    G12
  );


  not

  (
    G12_n,
    G12
  );


  buf

  (
    G13_p,
    G13
  );


  not

  (
    G13_n,
    G13
  );


  buf

  (
    G14_p,
    G14
  );


  not

  (
    G14_n,
    G14
  );


  buf

  (
    G15_p,
    G15
  );


  not

  (
    G15_n,
    G15
  );


  buf

  (
    G16_p,
    G16
  );


  not

  (
    G16_n,
    G16
  );


  buf

  (
    G17_p,
    G17
  );


  not

  (
    G17_n,
    G17
  );


  buf

  (
    G18_p,
    G18
  );


  not

  (
    G18_n,
    G18
  );


  buf

  (
    G19_p,
    G19
  );


  not

  (
    G19_n,
    G19
  );


  buf

  (
    G20_p,
    G20
  );


  not

  (
    G20_n,
    G20
  );


  buf

  (
    G21_p,
    G21
  );


  not

  (
    G21_n,
    G21
  );


  buf

  (
    G22_p,
    G22
  );


  not

  (
    G22_n,
    G22
  );


  buf

  (
    G23_p,
    G23
  );


  not

  (
    G23_n,
    G23
  );


  buf

  (
    G24_p,
    G24
  );


  not

  (
    G24_n,
    G24
  );


  buf

  (
    G25_p,
    G25
  );


  not

  (
    G25_n,
    G25
  );


  buf

  (
    G26_p,
    G26
  );


  not

  (
    G26_n,
    G26
  );


  buf

  (
    G27_p,
    G27
  );


  not

  (
    G27_n,
    G27
  );


  buf

  (
    G28_p,
    G28
  );


  not

  (
    G28_n,
    G28
  );


  buf

  (
    G29_p,
    G29
  );


  not

  (
    G29_n,
    G29
  );


  buf

  (
    G30_p,
    G30
  );


  not

  (
    G30_n,
    G30
  );


  buf

  (
    G31_p,
    G31
  );


  not

  (
    G31_n,
    G31
  );


  buf

  (
    G32_p,
    G32
  );


  not

  (
    G32_n,
    G32
  );


  and

  (
    g33_p,
    G17_p_spl_000,
    G1_p_spl_000
  );


  and

  (
    g34_p,
    G17_p_spl_000,
    G2_p_spl_000
  );


  or

  (
    g34_n,
    G17_n_spl_000,
    G2_n_spl_000
  );


  and

  (
    g35_p,
    G18_p_spl_000,
    G1_p_spl_000
  );


  or

  (
    g35_n,
    G18_n_spl_000,
    G1_n_spl_000
  );


  and

  (
    g36_p,
    g35_n,
    g34_p_spl_
  );


  or

  (
    g36_n,
    g35_p_spl_,
    g34_n_spl_
  );


  and

  (
    g37_p,
    g36_n,
    g34_p_spl_
  );


  or

  (
    g37_n,
    g36_p_spl_,
    g34_n_spl_
  );


  or

  (
    g38_n,
    g36_p_spl_,
    g35_p_spl_
  );


  and

  (
    g39_p,
    g38_n,
    g37_n_spl_0
  );


  and

  (
    g40_p,
    G19_p_spl_000,
    G1_p_spl_001
  );


  or

  (
    g40_n,
    G19_n_spl_000,
    G1_n_spl_000
  );


  and

  (
    g41_p,
    G17_p_spl_001,
    G3_p_spl_000
  );


  or

  (
    g41_n,
    G17_n_spl_000,
    G3_n_spl_000
  );


  and

  (
    g42_p,
    G18_p_spl_000,
    G2_p_spl_000
  );


  or

  (
    g42_n,
    G18_n_spl_000,
    G2_n_spl_000
  );


  and

  (
    g43_p,
    g42_n_spl_,
    g41_p_spl_
  );


  or

  (
    g43_n,
    g42_p_spl_,
    g41_n_spl_
  );


  and

  (
    g44_p,
    g43_n_spl_,
    g41_p_spl_
  );


  or

  (
    g44_n,
    g43_p_spl_,
    g41_n_spl_
  );


  and

  (
    g45_p,
    g43_n_spl_,
    g42_n_spl_
  );


  or

  (
    g45_n,
    g43_p_spl_,
    g42_p_spl_
  );


  and

  (
    g46_p,
    g45_n,
    g44_n_spl_0
  );


  or

  (
    g46_n,
    g45_p,
    g44_p_spl_0
  );


  and

  (
    g47_p,
    g46_n_spl_,
    g37_n_spl_0
  );


  or

  (
    g47_n,
    g46_p_spl_,
    g37_p_spl_
  );


  and

  (
    g48_p,
    g46_p_spl_,
    g37_p_spl_
  );


  or

  (
    g48_n,
    g46_n_spl_,
    g37_n_spl_
  );


  and

  (
    g49_p,
    g48_n,
    g47_n_spl_
  );


  or

  (
    g49_n,
    g48_p,
    g47_p_spl_
  );


  and

  (
    g50_p,
    g49_p,
    g40_n
  );


  or

  (
    g50_n,
    g49_n_spl_,
    g40_p_spl_
  );


  and

  (
    g51_p,
    g49_n_spl_,
    g40_p_spl_
  );


  or

  (
    g52_n,
    g51_p,
    g50_p_spl_
  );


  and

  (
    g53_p,
    G20_p_spl_000,
    G1_p_spl_001
  );


  or

  (
    g53_n,
    G20_n_spl_000,
    G1_n_spl_001
  );


  and

  (
    g54_p,
    g50_n,
    g47_n_spl_
  );


  or

  (
    g54_n,
    g50_p_spl_,
    g47_p_spl_
  );


  and

  (
    g55_p,
    G19_p_spl_000,
    G2_p_spl_001
  );


  or

  (
    g55_n,
    G19_n_spl_000,
    G2_n_spl_001
  );


  and

  (
    g56_p,
    G17_p_spl_001,
    G4_p_spl_000
  );


  or

  (
    g56_n,
    G17_n_spl_001,
    G4_n_spl_000
  );


  and

  (
    g57_p,
    G18_p_spl_001,
    G3_p_spl_000
  );


  or

  (
    g57_n,
    G18_n_spl_001,
    G3_n_spl_000
  );


  and

  (
    g58_p,
    g57_n_spl_,
    g56_p_spl_
  );


  or

  (
    g58_n,
    g57_p_spl_,
    g56_n_spl_
  );


  and

  (
    g59_p,
    g58_n_spl_,
    g56_p_spl_
  );


  or

  (
    g59_n,
    g58_p_spl_,
    g56_n_spl_
  );


  and

  (
    g60_p,
    g58_n_spl_,
    g57_n_spl_
  );


  or

  (
    g60_n,
    g58_p_spl_,
    g57_p_spl_
  );


  and

  (
    g61_p,
    g60_n,
    g59_n_spl_0
  );


  or

  (
    g61_n,
    g60_p,
    g59_p_spl_0
  );


  and

  (
    g62_p,
    g61_n_spl_,
    g44_n_spl_0
  );


  or

  (
    g62_n,
    g61_p_spl_,
    g44_p_spl_0
  );


  and

  (
    g63_p,
    g61_p_spl_,
    g44_p_spl_
  );


  or

  (
    g63_n,
    g61_n_spl_,
    g44_n_spl_
  );


  and

  (
    g64_p,
    g63_n,
    g62_n_spl_
  );


  or

  (
    g64_n,
    g63_p,
    g62_p_spl_
  );


  and

  (
    g65_p,
    g64_p_spl_,
    g55_n_spl_
  );


  or

  (
    g65_n,
    g64_n_spl_,
    g55_p_spl_
  );


  and

  (
    g66_p,
    g64_n_spl_,
    g55_p_spl_
  );


  or

  (
    g66_n,
    g64_p_spl_,
    g55_n_spl_
  );


  and

  (
    g67_p,
    g66_n,
    g65_n_spl_
  );


  or

  (
    g67_n,
    g66_p,
    g65_p_spl_
  );


  and

  (
    g68_p,
    g67_p_spl_,
    g54_n_spl_
  );


  or

  (
    g68_n,
    g67_n_spl_,
    g54_p_spl_
  );


  and

  (
    g69_p,
    g67_n_spl_,
    g54_p_spl_
  );


  or

  (
    g69_n,
    g67_p_spl_,
    g54_n_spl_
  );


  and

  (
    g70_p,
    g69_n,
    g68_n_spl_
  );


  or

  (
    g70_n,
    g69_p,
    g68_p_spl_
  );


  and

  (
    g71_p,
    g70_p,
    g53_n
  );


  or

  (
    g71_n,
    g70_n_spl_,
    g53_p_spl_
  );


  and

  (
    g72_p,
    g70_n_spl_,
    g53_p_spl_
  );


  or

  (
    g73_n,
    g72_p,
    g71_p_spl_
  );


  and

  (
    g74_p,
    G21_p_spl_000,
    G1_p_spl_010
  );


  or

  (
    g74_n,
    G21_n_spl_000,
    G1_n_spl_001
  );


  and

  (
    g75_p,
    g71_n,
    g68_n_spl_
  );


  or

  (
    g75_n,
    g71_p_spl_,
    g68_p_spl_
  );


  and

  (
    g76_p,
    G20_p_spl_000,
    G2_p_spl_001
  );


  or

  (
    g76_n,
    G20_n_spl_000,
    G2_n_spl_001
  );


  and

  (
    g77_p,
    g65_n_spl_,
    g62_n_spl_
  );


  or

  (
    g77_n,
    g65_p_spl_,
    g62_p_spl_
  );


  and

  (
    g78_p,
    G19_p_spl_001,
    G3_p_spl_001
  );


  or

  (
    g78_n,
    G19_n_spl_001,
    G3_n_spl_001
  );


  and

  (
    g79_p,
    G17_p_spl_010,
    G5_p_spl_000
  );


  or

  (
    g79_n,
    G17_n_spl_001,
    G5_n_spl_000
  );


  and

  (
    g80_p,
    G18_p_spl_001,
    G4_p_spl_000
  );


  or

  (
    g80_n,
    G18_n_spl_001,
    G4_n_spl_000
  );


  and

  (
    g81_p,
    g80_n_spl_,
    g79_p_spl_
  );


  or

  (
    g81_n,
    g80_p_spl_,
    g79_n_spl_
  );


  and

  (
    g82_p,
    g81_n_spl_,
    g79_p_spl_
  );


  or

  (
    g82_n,
    g81_p_spl_,
    g79_n_spl_
  );


  and

  (
    g83_p,
    g81_n_spl_,
    g80_n_spl_
  );


  or

  (
    g83_n,
    g81_p_spl_,
    g80_p_spl_
  );


  and

  (
    g84_p,
    g83_n,
    g82_n_spl_0
  );


  or

  (
    g84_n,
    g83_p,
    g82_p_spl_0
  );


  and

  (
    g85_p,
    g84_n_spl_,
    g59_n_spl_0
  );


  or

  (
    g85_n,
    g84_p_spl_,
    g59_p_spl_0
  );


  and

  (
    g86_p,
    g84_p_spl_,
    g59_p_spl_
  );


  or

  (
    g86_n,
    g84_n_spl_,
    g59_n_spl_
  );


  and

  (
    g87_p,
    g86_n,
    g85_n_spl_
  );


  or

  (
    g87_n,
    g86_p,
    g85_p_spl_
  );


  and

  (
    g88_p,
    g87_p_spl_,
    g78_n_spl_
  );


  or

  (
    g88_n,
    g87_n_spl_,
    g78_p_spl_
  );


  and

  (
    g89_p,
    g87_n_spl_,
    g78_p_spl_
  );


  or

  (
    g89_n,
    g87_p_spl_,
    g78_n_spl_
  );


  and

  (
    g90_p,
    g89_n,
    g88_n_spl_
  );


  or

  (
    g90_n,
    g89_p,
    g88_p_spl_
  );


  and

  (
    g91_p,
    g90_p_spl_,
    g77_n_spl_
  );


  or

  (
    g91_n,
    g90_n_spl_,
    g77_p_spl_
  );


  and

  (
    g92_p,
    g90_n_spl_,
    g77_p_spl_
  );


  or

  (
    g92_n,
    g90_p_spl_,
    g77_n_spl_
  );


  and

  (
    g93_p,
    g92_n,
    g91_n_spl_
  );


  or

  (
    g93_n,
    g92_p,
    g91_p_spl_
  );


  and

  (
    g94_p,
    g93_p_spl_,
    g76_n_spl_
  );


  or

  (
    g94_n,
    g93_n_spl_,
    g76_p_spl_
  );


  and

  (
    g95_p,
    g93_n_spl_,
    g76_p_spl_
  );


  or

  (
    g95_n,
    g93_p_spl_,
    g76_n_spl_
  );


  and

  (
    g96_p,
    g95_n,
    g94_n_spl_
  );


  or

  (
    g96_n,
    g95_p,
    g94_p_spl_
  );


  and

  (
    g97_p,
    g96_p_spl_,
    g75_n_spl_
  );


  or

  (
    g97_n,
    g96_n_spl_,
    g75_p_spl_
  );


  and

  (
    g98_p,
    g96_n_spl_,
    g75_p_spl_
  );


  or

  (
    g98_n,
    g96_p_spl_,
    g75_n_spl_
  );


  and

  (
    g99_p,
    g98_n,
    g97_n_spl_
  );


  or

  (
    g99_n,
    g98_p,
    g97_p_spl_
  );


  and

  (
    g100_p,
    g99_p,
    g74_n
  );


  or

  (
    g100_n,
    g99_n_spl_,
    g74_p_spl_
  );


  and

  (
    g101_p,
    g99_n_spl_,
    g74_p_spl_
  );


  or

  (
    g102_n,
    g101_p,
    g100_p_spl_
  );


  and

  (
    g103_p,
    G22_p_spl_000,
    G1_p_spl_010
  );


  or

  (
    g103_n,
    G22_n_spl_000,
    G1_n_spl_010
  );


  and

  (
    g104_p,
    g100_n,
    g97_n_spl_
  );


  or

  (
    g104_n,
    g100_p_spl_,
    g97_p_spl_
  );


  and

  (
    g105_p,
    G21_p_spl_000,
    G2_p_spl_010
  );


  or

  (
    g105_n,
    G21_n_spl_000,
    G2_n_spl_010
  );


  and

  (
    g106_p,
    g94_n_spl_,
    g91_n_spl_
  );


  or

  (
    g106_n,
    g94_p_spl_,
    g91_p_spl_
  );


  and

  (
    g107_p,
    G20_p_spl_001,
    G3_p_spl_001
  );


  or

  (
    g107_n,
    G20_n_spl_001,
    G3_n_spl_001
  );


  and

  (
    g108_p,
    g88_n_spl_,
    g85_n_spl_
  );


  or

  (
    g108_n,
    g88_p_spl_,
    g85_p_spl_
  );


  and

  (
    g109_p,
    G19_p_spl_001,
    G4_p_spl_001
  );


  or

  (
    g109_n,
    G19_n_spl_001,
    G4_n_spl_001
  );


  and

  (
    g110_p,
    G17_p_spl_010,
    G6_p_spl_000
  );


  or

  (
    g110_n,
    G17_n_spl_010,
    G6_n_spl_000
  );


  and

  (
    g111_p,
    G18_p_spl_010,
    G5_p_spl_000
  );


  or

  (
    g111_n,
    G18_n_spl_010,
    G5_n_spl_000
  );


  and

  (
    g112_p,
    g111_n_spl_,
    g110_p_spl_
  );


  or

  (
    g112_n,
    g111_p_spl_,
    g110_n_spl_
  );


  and

  (
    g113_p,
    g112_n_spl_,
    g110_p_spl_
  );


  or

  (
    g113_n,
    g112_p_spl_,
    g110_n_spl_
  );


  and

  (
    g114_p,
    g112_n_spl_,
    g111_n_spl_
  );


  or

  (
    g114_n,
    g112_p_spl_,
    g111_p_spl_
  );


  and

  (
    g115_p,
    g114_n,
    g113_n_spl_0
  );


  or

  (
    g115_n,
    g114_p,
    g113_p_spl_0
  );


  and

  (
    g116_p,
    g115_n_spl_,
    g82_n_spl_0
  );


  or

  (
    g116_n,
    g115_p_spl_,
    g82_p_spl_0
  );


  and

  (
    g117_p,
    g115_p_spl_,
    g82_p_spl_
  );


  or

  (
    g117_n,
    g115_n_spl_,
    g82_n_spl_
  );


  and

  (
    g118_p,
    g117_n,
    g116_n_spl_
  );


  or

  (
    g118_n,
    g117_p,
    g116_p_spl_
  );


  and

  (
    g119_p,
    g118_p_spl_,
    g109_n_spl_
  );


  or

  (
    g119_n,
    g118_n_spl_,
    g109_p_spl_
  );


  and

  (
    g120_p,
    g118_n_spl_,
    g109_p_spl_
  );


  or

  (
    g120_n,
    g118_p_spl_,
    g109_n_spl_
  );


  and

  (
    g121_p,
    g120_n,
    g119_n_spl_
  );


  or

  (
    g121_n,
    g120_p,
    g119_p_spl_
  );


  and

  (
    g122_p,
    g121_p_spl_,
    g108_n_spl_
  );


  or

  (
    g122_n,
    g121_n_spl_,
    g108_p_spl_
  );


  and

  (
    g123_p,
    g121_n_spl_,
    g108_p_spl_
  );


  or

  (
    g123_n,
    g121_p_spl_,
    g108_n_spl_
  );


  and

  (
    g124_p,
    g123_n,
    g122_n_spl_
  );


  or

  (
    g124_n,
    g123_p,
    g122_p_spl_
  );


  and

  (
    g125_p,
    g124_p_spl_,
    g107_n_spl_
  );


  or

  (
    g125_n,
    g124_n_spl_,
    g107_p_spl_
  );


  and

  (
    g126_p,
    g124_n_spl_,
    g107_p_spl_
  );


  or

  (
    g126_n,
    g124_p_spl_,
    g107_n_spl_
  );


  and

  (
    g127_p,
    g126_n,
    g125_n_spl_
  );


  or

  (
    g127_n,
    g126_p,
    g125_p_spl_
  );


  and

  (
    g128_p,
    g127_p_spl_,
    g106_n_spl_
  );


  or

  (
    g128_n,
    g127_n_spl_,
    g106_p_spl_
  );


  and

  (
    g129_p,
    g127_n_spl_,
    g106_p_spl_
  );


  or

  (
    g129_n,
    g127_p_spl_,
    g106_n_spl_
  );


  and

  (
    g130_p,
    g129_n,
    g128_n_spl_
  );


  or

  (
    g130_n,
    g129_p,
    g128_p_spl_
  );


  and

  (
    g131_p,
    g130_p_spl_,
    g105_n_spl_
  );


  or

  (
    g131_n,
    g130_n_spl_,
    g105_p_spl_
  );


  and

  (
    g132_p,
    g130_n_spl_,
    g105_p_spl_
  );


  or

  (
    g132_n,
    g130_p_spl_,
    g105_n_spl_
  );


  and

  (
    g133_p,
    g132_n,
    g131_n_spl_
  );


  or

  (
    g133_n,
    g132_p,
    g131_p_spl_
  );


  and

  (
    g134_p,
    g133_p_spl_,
    g104_n_spl_
  );


  or

  (
    g134_n,
    g133_n_spl_,
    g104_p_spl_
  );


  and

  (
    g135_p,
    g133_n_spl_,
    g104_p_spl_
  );


  or

  (
    g135_n,
    g133_p_spl_,
    g104_n_spl_
  );


  and

  (
    g136_p,
    g135_n,
    g134_n_spl_
  );


  or

  (
    g136_n,
    g135_p,
    g134_p_spl_
  );


  and

  (
    g137_p,
    g136_p,
    g103_n
  );


  or

  (
    g137_n,
    g136_n_spl_,
    g103_p_spl_
  );


  and

  (
    g138_p,
    g136_n_spl_,
    g103_p_spl_
  );


  or

  (
    g139_n,
    g138_p,
    g137_p_spl_
  );


  and

  (
    g140_p,
    G23_p_spl_000,
    G1_p_spl_011
  );


  or

  (
    g140_n,
    G23_n_spl_000,
    G1_n_spl_010
  );


  and

  (
    g141_p,
    g137_n,
    g134_n_spl_
  );


  or

  (
    g141_n,
    g137_p_spl_,
    g134_p_spl_
  );


  and

  (
    g142_p,
    G22_p_spl_000,
    G2_p_spl_010
  );


  or

  (
    g142_n,
    G22_n_spl_000,
    G2_n_spl_010
  );


  and

  (
    g143_p,
    g131_n_spl_,
    g128_n_spl_
  );


  or

  (
    g143_n,
    g131_p_spl_,
    g128_p_spl_
  );


  and

  (
    g144_p,
    G21_p_spl_001,
    G3_p_spl_010
  );


  or

  (
    g144_n,
    G21_n_spl_001,
    G3_n_spl_010
  );


  and

  (
    g145_p,
    g125_n_spl_,
    g122_n_spl_
  );


  or

  (
    g145_n,
    g125_p_spl_,
    g122_p_spl_
  );


  and

  (
    g146_p,
    G20_p_spl_001,
    G4_p_spl_001
  );


  or

  (
    g146_n,
    G20_n_spl_001,
    G4_n_spl_001
  );


  and

  (
    g147_p,
    g119_n_spl_,
    g116_n_spl_
  );


  or

  (
    g147_n,
    g119_p_spl_,
    g116_p_spl_
  );


  and

  (
    g148_p,
    G19_p_spl_010,
    G5_p_spl_001
  );


  or

  (
    g148_n,
    G19_n_spl_010,
    G5_n_spl_001
  );


  and

  (
    g149_p,
    G17_p_spl_011,
    G7_p_spl_000
  );


  or

  (
    g149_n,
    G17_n_spl_010,
    G7_n_spl_000
  );


  and

  (
    g150_p,
    G18_p_spl_010,
    G6_p_spl_000
  );


  or

  (
    g150_n,
    G18_n_spl_010,
    G6_n_spl_000
  );


  and

  (
    g151_p,
    g150_n_spl_,
    g149_p_spl_
  );


  or

  (
    g151_n,
    g150_p_spl_,
    g149_n_spl_
  );


  and

  (
    g152_p,
    g151_n_spl_,
    g149_p_spl_
  );


  or

  (
    g152_n,
    g151_p_spl_,
    g149_n_spl_
  );


  and

  (
    g153_p,
    g151_n_spl_,
    g150_n_spl_
  );


  or

  (
    g153_n,
    g151_p_spl_,
    g150_p_spl_
  );


  and

  (
    g154_p,
    g153_n,
    g152_n_spl_0
  );


  or

  (
    g154_n,
    g153_p,
    g152_p_spl_0
  );


  and

  (
    g155_p,
    g154_n_spl_,
    g113_n_spl_0
  );


  or

  (
    g155_n,
    g154_p_spl_,
    g113_p_spl_0
  );


  and

  (
    g156_p,
    g154_p_spl_,
    g113_p_spl_
  );


  or

  (
    g156_n,
    g154_n_spl_,
    g113_n_spl_
  );


  and

  (
    g157_p,
    g156_n,
    g155_n_spl_
  );


  or

  (
    g157_n,
    g156_p,
    g155_p_spl_
  );


  and

  (
    g158_p,
    g157_p_spl_,
    g148_n_spl_
  );


  or

  (
    g158_n,
    g157_n_spl_,
    g148_p_spl_
  );


  and

  (
    g159_p,
    g157_n_spl_,
    g148_p_spl_
  );


  or

  (
    g159_n,
    g157_p_spl_,
    g148_n_spl_
  );


  and

  (
    g160_p,
    g159_n,
    g158_n_spl_
  );


  or

  (
    g160_n,
    g159_p,
    g158_p_spl_
  );


  and

  (
    g161_p,
    g160_p_spl_,
    g147_n_spl_
  );


  or

  (
    g161_n,
    g160_n_spl_,
    g147_p_spl_
  );


  and

  (
    g162_p,
    g160_n_spl_,
    g147_p_spl_
  );


  or

  (
    g162_n,
    g160_p_spl_,
    g147_n_spl_
  );


  and

  (
    g163_p,
    g162_n,
    g161_n_spl_
  );


  or

  (
    g163_n,
    g162_p,
    g161_p_spl_
  );


  and

  (
    g164_p,
    g163_p_spl_,
    g146_n_spl_
  );


  or

  (
    g164_n,
    g163_n_spl_,
    g146_p_spl_
  );


  and

  (
    g165_p,
    g163_n_spl_,
    g146_p_spl_
  );


  or

  (
    g165_n,
    g163_p_spl_,
    g146_n_spl_
  );


  and

  (
    g166_p,
    g165_n,
    g164_n_spl_
  );


  or

  (
    g166_n,
    g165_p,
    g164_p_spl_
  );


  and

  (
    g167_p,
    g166_p_spl_,
    g145_n_spl_
  );


  or

  (
    g167_n,
    g166_n_spl_,
    g145_p_spl_
  );


  and

  (
    g168_p,
    g166_n_spl_,
    g145_p_spl_
  );


  or

  (
    g168_n,
    g166_p_spl_,
    g145_n_spl_
  );


  and

  (
    g169_p,
    g168_n,
    g167_n_spl_
  );


  or

  (
    g169_n,
    g168_p,
    g167_p_spl_
  );


  and

  (
    g170_p,
    g169_p_spl_,
    g144_n_spl_
  );


  or

  (
    g170_n,
    g169_n_spl_,
    g144_p_spl_
  );


  and

  (
    g171_p,
    g169_n_spl_,
    g144_p_spl_
  );


  or

  (
    g171_n,
    g169_p_spl_,
    g144_n_spl_
  );


  and

  (
    g172_p,
    g171_n,
    g170_n_spl_
  );


  or

  (
    g172_n,
    g171_p,
    g170_p_spl_
  );


  and

  (
    g173_p,
    g172_p_spl_,
    g143_n_spl_
  );


  or

  (
    g173_n,
    g172_n_spl_,
    g143_p_spl_
  );


  and

  (
    g174_p,
    g172_n_spl_,
    g143_p_spl_
  );


  or

  (
    g174_n,
    g172_p_spl_,
    g143_n_spl_
  );


  and

  (
    g175_p,
    g174_n,
    g173_n_spl_
  );


  or

  (
    g175_n,
    g174_p,
    g173_p_spl_
  );


  and

  (
    g176_p,
    g175_p_spl_,
    g142_n_spl_
  );


  or

  (
    g176_n,
    g175_n_spl_,
    g142_p_spl_
  );


  and

  (
    g177_p,
    g175_n_spl_,
    g142_p_spl_
  );


  or

  (
    g177_n,
    g175_p_spl_,
    g142_n_spl_
  );


  and

  (
    g178_p,
    g177_n,
    g176_n_spl_
  );


  or

  (
    g178_n,
    g177_p,
    g176_p_spl_
  );


  and

  (
    g179_p,
    g178_p_spl_,
    g141_n_spl_
  );


  or

  (
    g179_n,
    g178_n_spl_,
    g141_p_spl_
  );


  and

  (
    g180_p,
    g178_n_spl_,
    g141_p_spl_
  );


  or

  (
    g180_n,
    g178_p_spl_,
    g141_n_spl_
  );


  and

  (
    g181_p,
    g180_n,
    g179_n_spl_
  );


  or

  (
    g181_n,
    g180_p,
    g179_p_spl_
  );


  and

  (
    g182_p,
    g181_p,
    g140_n
  );


  or

  (
    g182_n,
    g181_n_spl_,
    g140_p_spl_
  );


  and

  (
    g183_p,
    g181_n_spl_,
    g140_p_spl_
  );


  or

  (
    g184_n,
    g183_p,
    g182_p_spl_
  );


  and

  (
    g185_p,
    G24_p_spl_000,
    G1_p_spl_011
  );


  or

  (
    g185_n,
    G24_n_spl_000,
    G1_n_spl_011
  );


  and

  (
    g186_p,
    g182_n,
    g179_n_spl_
  );


  or

  (
    g186_n,
    g182_p_spl_,
    g179_p_spl_
  );


  and

  (
    g187_p,
    G23_p_spl_000,
    G2_p_spl_011
  );


  or

  (
    g187_n,
    G23_n_spl_000,
    G2_n_spl_011
  );


  and

  (
    g188_p,
    g176_n_spl_,
    g173_n_spl_
  );


  or

  (
    g188_n,
    g176_p_spl_,
    g173_p_spl_
  );


  and

  (
    g189_p,
    G22_p_spl_001,
    G3_p_spl_010
  );


  or

  (
    g189_n,
    G22_n_spl_001,
    G3_n_spl_010
  );


  and

  (
    g190_p,
    g170_n_spl_,
    g167_n_spl_
  );


  or

  (
    g190_n,
    g170_p_spl_,
    g167_p_spl_
  );


  and

  (
    g191_p,
    G21_p_spl_001,
    G4_p_spl_010
  );


  or

  (
    g191_n,
    G21_n_spl_001,
    G4_n_spl_010
  );


  and

  (
    g192_p,
    g164_n_spl_,
    g161_n_spl_
  );


  or

  (
    g192_n,
    g164_p_spl_,
    g161_p_spl_
  );


  and

  (
    g193_p,
    G20_p_spl_010,
    G5_p_spl_001
  );


  or

  (
    g193_n,
    G20_n_spl_010,
    G5_n_spl_001
  );


  and

  (
    g194_p,
    g158_n_spl_,
    g155_n_spl_
  );


  or

  (
    g194_n,
    g158_p_spl_,
    g155_p_spl_
  );


  and

  (
    g195_p,
    G19_p_spl_010,
    G6_p_spl_001
  );


  or

  (
    g195_n,
    G19_n_spl_010,
    G6_n_spl_001
  );


  and

  (
    g196_p,
    G17_p_spl_011,
    G8_p_spl_000
  );


  or

  (
    g196_n,
    G17_n_spl_011,
    G8_n_spl_000
  );


  and

  (
    g197_p,
    G18_p_spl_011,
    G7_p_spl_000
  );


  or

  (
    g197_n,
    G18_n_spl_011,
    G7_n_spl_000
  );


  and

  (
    g198_p,
    g197_n_spl_,
    g196_p_spl_
  );


  or

  (
    g198_n,
    g197_p_spl_,
    g196_n_spl_
  );


  and

  (
    g199_p,
    g198_n_spl_,
    g196_p_spl_
  );


  or

  (
    g199_n,
    g198_p_spl_,
    g196_n_spl_
  );


  and

  (
    g200_p,
    g198_n_spl_,
    g197_n_spl_
  );


  or

  (
    g200_n,
    g198_p_spl_,
    g197_p_spl_
  );


  and

  (
    g201_p,
    g200_n,
    g199_n_spl_0
  );


  or

  (
    g201_n,
    g200_p,
    g199_p_spl_0
  );


  and

  (
    g202_p,
    g201_n_spl_,
    g152_n_spl_0
  );


  or

  (
    g202_n,
    g201_p_spl_,
    g152_p_spl_0
  );


  and

  (
    g203_p,
    g201_p_spl_,
    g152_p_spl_
  );


  or

  (
    g203_n,
    g201_n_spl_,
    g152_n_spl_
  );


  and

  (
    g204_p,
    g203_n,
    g202_n_spl_
  );


  or

  (
    g204_n,
    g203_p,
    g202_p_spl_
  );


  and

  (
    g205_p,
    g204_p_spl_,
    g195_n_spl_
  );


  or

  (
    g205_n,
    g204_n_spl_,
    g195_p_spl_
  );


  and

  (
    g206_p,
    g204_n_spl_,
    g195_p_spl_
  );


  or

  (
    g206_n,
    g204_p_spl_,
    g195_n_spl_
  );


  and

  (
    g207_p,
    g206_n,
    g205_n_spl_
  );


  or

  (
    g207_n,
    g206_p,
    g205_p_spl_
  );


  and

  (
    g208_p,
    g207_p_spl_,
    g194_n_spl_
  );


  or

  (
    g208_n,
    g207_n_spl_,
    g194_p_spl_
  );


  and

  (
    g209_p,
    g207_n_spl_,
    g194_p_spl_
  );


  or

  (
    g209_n,
    g207_p_spl_,
    g194_n_spl_
  );


  and

  (
    g210_p,
    g209_n,
    g208_n_spl_
  );


  or

  (
    g210_n,
    g209_p,
    g208_p_spl_
  );


  and

  (
    g211_p,
    g210_p_spl_,
    g193_n_spl_
  );


  or

  (
    g211_n,
    g210_n_spl_,
    g193_p_spl_
  );


  and

  (
    g212_p,
    g210_n_spl_,
    g193_p_spl_
  );


  or

  (
    g212_n,
    g210_p_spl_,
    g193_n_spl_
  );


  and

  (
    g213_p,
    g212_n,
    g211_n_spl_
  );


  or

  (
    g213_n,
    g212_p,
    g211_p_spl_
  );


  and

  (
    g214_p,
    g213_p_spl_,
    g192_n_spl_
  );


  or

  (
    g214_n,
    g213_n_spl_,
    g192_p_spl_
  );


  and

  (
    g215_p,
    g213_n_spl_,
    g192_p_spl_
  );


  or

  (
    g215_n,
    g213_p_spl_,
    g192_n_spl_
  );


  and

  (
    g216_p,
    g215_n,
    g214_n_spl_
  );


  or

  (
    g216_n,
    g215_p,
    g214_p_spl_
  );


  and

  (
    g217_p,
    g216_p_spl_,
    g191_n_spl_
  );


  or

  (
    g217_n,
    g216_n_spl_,
    g191_p_spl_
  );


  and

  (
    g218_p,
    g216_n_spl_,
    g191_p_spl_
  );


  or

  (
    g218_n,
    g216_p_spl_,
    g191_n_spl_
  );


  and

  (
    g219_p,
    g218_n,
    g217_n_spl_
  );


  or

  (
    g219_n,
    g218_p,
    g217_p_spl_
  );


  and

  (
    g220_p,
    g219_p_spl_,
    g190_n_spl_
  );


  or

  (
    g220_n,
    g219_n_spl_,
    g190_p_spl_
  );


  and

  (
    g221_p,
    g219_n_spl_,
    g190_p_spl_
  );


  or

  (
    g221_n,
    g219_p_spl_,
    g190_n_spl_
  );


  and

  (
    g222_p,
    g221_n,
    g220_n_spl_
  );


  or

  (
    g222_n,
    g221_p,
    g220_p_spl_
  );


  and

  (
    g223_p,
    g222_p_spl_,
    g189_n_spl_
  );


  or

  (
    g223_n,
    g222_n_spl_,
    g189_p_spl_
  );


  and

  (
    g224_p,
    g222_n_spl_,
    g189_p_spl_
  );


  or

  (
    g224_n,
    g222_p_spl_,
    g189_n_spl_
  );


  and

  (
    g225_p,
    g224_n,
    g223_n_spl_
  );


  or

  (
    g225_n,
    g224_p,
    g223_p_spl_
  );


  and

  (
    g226_p,
    g225_p_spl_,
    g188_n_spl_
  );


  or

  (
    g226_n,
    g225_n_spl_,
    g188_p_spl_
  );


  and

  (
    g227_p,
    g225_n_spl_,
    g188_p_spl_
  );


  or

  (
    g227_n,
    g225_p_spl_,
    g188_n_spl_
  );


  and

  (
    g228_p,
    g227_n,
    g226_n_spl_
  );


  or

  (
    g228_n,
    g227_p,
    g226_p_spl_
  );


  and

  (
    g229_p,
    g228_p_spl_,
    g187_n_spl_
  );


  or

  (
    g229_n,
    g228_n_spl_,
    g187_p_spl_
  );


  and

  (
    g230_p,
    g228_n_spl_,
    g187_p_spl_
  );


  or

  (
    g230_n,
    g228_p_spl_,
    g187_n_spl_
  );


  and

  (
    g231_p,
    g230_n,
    g229_n_spl_
  );


  or

  (
    g231_n,
    g230_p,
    g229_p_spl_
  );


  and

  (
    g232_p,
    g231_p_spl_,
    g186_n_spl_
  );


  or

  (
    g232_n,
    g231_n_spl_,
    g186_p_spl_
  );


  and

  (
    g233_p,
    g231_n_spl_,
    g186_p_spl_
  );


  or

  (
    g233_n,
    g231_p_spl_,
    g186_n_spl_
  );


  and

  (
    g234_p,
    g233_n,
    g232_n_spl_
  );


  or

  (
    g234_n,
    g233_p,
    g232_p_spl_
  );


  and

  (
    g235_p,
    g234_p,
    g185_n
  );


  or

  (
    g235_n,
    g234_n_spl_,
    g185_p_spl_
  );


  and

  (
    g236_p,
    g234_n_spl_,
    g185_p_spl_
  );


  or

  (
    g237_n,
    g236_p,
    g235_p_spl_
  );


  and

  (
    g238_p,
    G25_p_spl_000,
    G1_p_spl_100
  );


  or

  (
    g238_n,
    G25_n_spl_000,
    G1_n_spl_011
  );


  and

  (
    g239_p,
    g235_n,
    g232_n_spl_
  );


  or

  (
    g239_n,
    g235_p_spl_,
    g232_p_spl_
  );


  and

  (
    g240_p,
    G24_p_spl_000,
    G2_p_spl_011
  );


  or

  (
    g240_n,
    G24_n_spl_000,
    G2_n_spl_011
  );


  and

  (
    g241_p,
    g229_n_spl_,
    g226_n_spl_
  );


  or

  (
    g241_n,
    g229_p_spl_,
    g226_p_spl_
  );


  and

  (
    g242_p,
    G23_p_spl_001,
    G3_p_spl_011
  );


  or

  (
    g242_n,
    G23_n_spl_001,
    G3_n_spl_011
  );


  and

  (
    g243_p,
    g223_n_spl_,
    g220_n_spl_
  );


  or

  (
    g243_n,
    g223_p_spl_,
    g220_p_spl_
  );


  and

  (
    g244_p,
    G22_p_spl_001,
    G4_p_spl_010
  );


  or

  (
    g244_n,
    G22_n_spl_001,
    G4_n_spl_010
  );


  and

  (
    g245_p,
    g217_n_spl_,
    g214_n_spl_
  );


  or

  (
    g245_n,
    g217_p_spl_,
    g214_p_spl_
  );


  and

  (
    g246_p,
    G21_p_spl_010,
    G5_p_spl_010
  );


  or

  (
    g246_n,
    G21_n_spl_010,
    G5_n_spl_010
  );


  and

  (
    g247_p,
    g211_n_spl_,
    g208_n_spl_
  );


  or

  (
    g247_n,
    g211_p_spl_,
    g208_p_spl_
  );


  and

  (
    g248_p,
    G20_p_spl_010,
    G6_p_spl_001
  );


  or

  (
    g248_n,
    G20_n_spl_010,
    G6_n_spl_001
  );


  and

  (
    g249_p,
    g205_n_spl_,
    g202_n_spl_
  );


  or

  (
    g249_n,
    g205_p_spl_,
    g202_p_spl_
  );


  and

  (
    g250_p,
    G19_p_spl_011,
    G7_p_spl_001
  );


  or

  (
    g250_n,
    G19_n_spl_011,
    G7_n_spl_001
  );


  and

  (
    g251_p,
    G17_p_spl_100,
    G9_p_spl_000
  );


  or

  (
    g251_n,
    G17_n_spl_011,
    G9_n_spl_000
  );


  and

  (
    g252_p,
    G18_p_spl_011,
    G8_p_spl_000
  );


  or

  (
    g252_n,
    G18_n_spl_011,
    G8_n_spl_000
  );


  and

  (
    g253_p,
    g252_n_spl_,
    g251_p_spl_
  );


  or

  (
    g253_n,
    g252_p_spl_,
    g251_n_spl_
  );


  and

  (
    g254_p,
    g253_n_spl_,
    g251_p_spl_
  );


  or

  (
    g254_n,
    g253_p_spl_,
    g251_n_spl_
  );


  and

  (
    g255_p,
    g253_n_spl_,
    g252_n_spl_
  );


  or

  (
    g255_n,
    g253_p_spl_,
    g252_p_spl_
  );


  and

  (
    g256_p,
    g255_n,
    g254_n_spl_0
  );


  or

  (
    g256_n,
    g255_p,
    g254_p_spl_0
  );


  and

  (
    g257_p,
    g256_n_spl_,
    g199_n_spl_0
  );


  or

  (
    g257_n,
    g256_p_spl_,
    g199_p_spl_0
  );


  and

  (
    g258_p,
    g256_p_spl_,
    g199_p_spl_
  );


  or

  (
    g258_n,
    g256_n_spl_,
    g199_n_spl_
  );


  and

  (
    g259_p,
    g258_n,
    g257_n_spl_
  );


  or

  (
    g259_n,
    g258_p,
    g257_p_spl_
  );


  and

  (
    g260_p,
    g259_p_spl_,
    g250_n_spl_
  );


  or

  (
    g260_n,
    g259_n_spl_,
    g250_p_spl_
  );


  and

  (
    g261_p,
    g259_n_spl_,
    g250_p_spl_
  );


  or

  (
    g261_n,
    g259_p_spl_,
    g250_n_spl_
  );


  and

  (
    g262_p,
    g261_n,
    g260_n_spl_
  );


  or

  (
    g262_n,
    g261_p,
    g260_p_spl_
  );


  and

  (
    g263_p,
    g262_p_spl_,
    g249_n_spl_
  );


  or

  (
    g263_n,
    g262_n_spl_,
    g249_p_spl_
  );


  and

  (
    g264_p,
    g262_n_spl_,
    g249_p_spl_
  );


  or

  (
    g264_n,
    g262_p_spl_,
    g249_n_spl_
  );


  and

  (
    g265_p,
    g264_n,
    g263_n_spl_
  );


  or

  (
    g265_n,
    g264_p,
    g263_p_spl_
  );


  and

  (
    g266_p,
    g265_p_spl_,
    g248_n_spl_
  );


  or

  (
    g266_n,
    g265_n_spl_,
    g248_p_spl_
  );


  and

  (
    g267_p,
    g265_n_spl_,
    g248_p_spl_
  );


  or

  (
    g267_n,
    g265_p_spl_,
    g248_n_spl_
  );


  and

  (
    g268_p,
    g267_n,
    g266_n_spl_
  );


  or

  (
    g268_n,
    g267_p,
    g266_p_spl_
  );


  and

  (
    g269_p,
    g268_p_spl_,
    g247_n_spl_
  );


  or

  (
    g269_n,
    g268_n_spl_,
    g247_p_spl_
  );


  and

  (
    g270_p,
    g268_n_spl_,
    g247_p_spl_
  );


  or

  (
    g270_n,
    g268_p_spl_,
    g247_n_spl_
  );


  and

  (
    g271_p,
    g270_n,
    g269_n_spl_
  );


  or

  (
    g271_n,
    g270_p,
    g269_p_spl_
  );


  and

  (
    g272_p,
    g271_p_spl_,
    g246_n_spl_
  );


  or

  (
    g272_n,
    g271_n_spl_,
    g246_p_spl_
  );


  and

  (
    g273_p,
    g271_n_spl_,
    g246_p_spl_
  );


  or

  (
    g273_n,
    g271_p_spl_,
    g246_n_spl_
  );


  and

  (
    g274_p,
    g273_n,
    g272_n_spl_
  );


  or

  (
    g274_n,
    g273_p,
    g272_p_spl_
  );


  and

  (
    g275_p,
    g274_p_spl_,
    g245_n_spl_
  );


  or

  (
    g275_n,
    g274_n_spl_,
    g245_p_spl_
  );


  and

  (
    g276_p,
    g274_n_spl_,
    g245_p_spl_
  );


  or

  (
    g276_n,
    g274_p_spl_,
    g245_n_spl_
  );


  and

  (
    g277_p,
    g276_n,
    g275_n_spl_
  );


  or

  (
    g277_n,
    g276_p,
    g275_p_spl_
  );


  and

  (
    g278_p,
    g277_p_spl_,
    g244_n_spl_
  );


  or

  (
    g278_n,
    g277_n_spl_,
    g244_p_spl_
  );


  and

  (
    g279_p,
    g277_n_spl_,
    g244_p_spl_
  );


  or

  (
    g279_n,
    g277_p_spl_,
    g244_n_spl_
  );


  and

  (
    g280_p,
    g279_n,
    g278_n_spl_
  );


  or

  (
    g280_n,
    g279_p,
    g278_p_spl_
  );


  and

  (
    g281_p,
    g280_p_spl_,
    g243_n_spl_
  );


  or

  (
    g281_n,
    g280_n_spl_,
    g243_p_spl_
  );


  and

  (
    g282_p,
    g280_n_spl_,
    g243_p_spl_
  );


  or

  (
    g282_n,
    g280_p_spl_,
    g243_n_spl_
  );


  and

  (
    g283_p,
    g282_n,
    g281_n_spl_
  );


  or

  (
    g283_n,
    g282_p,
    g281_p_spl_
  );


  and

  (
    g284_p,
    g283_p_spl_,
    g242_n_spl_
  );


  or

  (
    g284_n,
    g283_n_spl_,
    g242_p_spl_
  );


  and

  (
    g285_p,
    g283_n_spl_,
    g242_p_spl_
  );


  or

  (
    g285_n,
    g283_p_spl_,
    g242_n_spl_
  );


  and

  (
    g286_p,
    g285_n,
    g284_n_spl_
  );


  or

  (
    g286_n,
    g285_p,
    g284_p_spl_
  );


  and

  (
    g287_p,
    g286_p_spl_,
    g241_n_spl_
  );


  or

  (
    g287_n,
    g286_n_spl_,
    g241_p_spl_
  );


  and

  (
    g288_p,
    g286_n_spl_,
    g241_p_spl_
  );


  or

  (
    g288_n,
    g286_p_spl_,
    g241_n_spl_
  );


  and

  (
    g289_p,
    g288_n,
    g287_n_spl_
  );


  or

  (
    g289_n,
    g288_p,
    g287_p_spl_
  );


  and

  (
    g290_p,
    g289_p_spl_,
    g240_n_spl_
  );


  or

  (
    g290_n,
    g289_n_spl_,
    g240_p_spl_
  );


  and

  (
    g291_p,
    g289_n_spl_,
    g240_p_spl_
  );


  or

  (
    g291_n,
    g289_p_spl_,
    g240_n_spl_
  );


  and

  (
    g292_p,
    g291_n,
    g290_n_spl_
  );


  or

  (
    g292_n,
    g291_p,
    g290_p_spl_
  );


  and

  (
    g293_p,
    g292_p_spl_,
    g239_n_spl_
  );


  or

  (
    g293_n,
    g292_n_spl_,
    g239_p_spl_
  );


  and

  (
    g294_p,
    g292_n_spl_,
    g239_p_spl_
  );


  or

  (
    g294_n,
    g292_p_spl_,
    g239_n_spl_
  );


  and

  (
    g295_p,
    g294_n,
    g293_n_spl_
  );


  or

  (
    g295_n,
    g294_p,
    g293_p_spl_
  );


  and

  (
    g296_p,
    g295_p,
    g238_n
  );


  or

  (
    g296_n,
    g295_n_spl_,
    g238_p_spl_
  );


  and

  (
    g297_p,
    g295_n_spl_,
    g238_p_spl_
  );


  or

  (
    g298_n,
    g297_p,
    g296_p_spl_
  );


  and

  (
    g299_p,
    G26_p_spl_000,
    G1_p_spl_100
  );


  or

  (
    g299_n,
    G26_n_spl_000,
    G1_n_spl_100
  );


  and

  (
    g300_p,
    g296_n,
    g293_n_spl_
  );


  or

  (
    g300_n,
    g296_p_spl_,
    g293_p_spl_
  );


  and

  (
    g301_p,
    G25_p_spl_000,
    G2_p_spl_100
  );


  or

  (
    g301_n,
    G25_n_spl_000,
    G2_n_spl_100
  );


  and

  (
    g302_p,
    g290_n_spl_,
    g287_n_spl_
  );


  or

  (
    g302_n,
    g290_p_spl_,
    g287_p_spl_
  );


  and

  (
    g303_p,
    G24_p_spl_001,
    G3_p_spl_011
  );


  or

  (
    g303_n,
    G24_n_spl_001,
    G3_n_spl_011
  );


  and

  (
    g304_p,
    g284_n_spl_,
    g281_n_spl_
  );


  or

  (
    g304_n,
    g284_p_spl_,
    g281_p_spl_
  );


  and

  (
    g305_p,
    G23_p_spl_001,
    G4_p_spl_011
  );


  or

  (
    g305_n,
    G23_n_spl_001,
    G4_n_spl_011
  );


  and

  (
    g306_p,
    g278_n_spl_,
    g275_n_spl_
  );


  or

  (
    g306_n,
    g278_p_spl_,
    g275_p_spl_
  );


  and

  (
    g307_p,
    G22_p_spl_010,
    G5_p_spl_010
  );


  or

  (
    g307_n,
    G22_n_spl_010,
    G5_n_spl_010
  );


  and

  (
    g308_p,
    g272_n_spl_,
    g269_n_spl_
  );


  or

  (
    g308_n,
    g272_p_spl_,
    g269_p_spl_
  );


  and

  (
    g309_p,
    G21_p_spl_010,
    G6_p_spl_010
  );


  or

  (
    g309_n,
    G21_n_spl_010,
    G6_n_spl_010
  );


  and

  (
    g310_p,
    g266_n_spl_,
    g263_n_spl_
  );


  or

  (
    g310_n,
    g266_p_spl_,
    g263_p_spl_
  );


  and

  (
    g311_p,
    G20_p_spl_011,
    G7_p_spl_001
  );


  or

  (
    g311_n,
    G20_n_spl_011,
    G7_n_spl_001
  );


  and

  (
    g312_p,
    g260_n_spl_,
    g257_n_spl_
  );


  or

  (
    g312_n,
    g260_p_spl_,
    g257_p_spl_
  );


  and

  (
    g313_p,
    G19_p_spl_011,
    G8_p_spl_001
  );


  or

  (
    g313_n,
    G19_n_spl_011,
    G8_n_spl_001
  );


  and

  (
    g314_p,
    G17_p_spl_100,
    G10_p_spl_000
  );


  or

  (
    g314_n,
    G17_n_spl_100,
    G10_n_spl_000
  );


  and

  (
    g315_p,
    G18_p_spl_100,
    G9_p_spl_000
  );


  or

  (
    g315_n,
    G18_n_spl_100,
    G9_n_spl_000
  );


  and

  (
    g316_p,
    g315_n_spl_,
    g314_p_spl_
  );


  or

  (
    g316_n,
    g315_p_spl_,
    g314_n_spl_
  );


  and

  (
    g317_p,
    g316_n_spl_,
    g314_p_spl_
  );


  or

  (
    g317_n,
    g316_p_spl_,
    g314_n_spl_
  );


  and

  (
    g318_p,
    g316_n_spl_,
    g315_n_spl_
  );


  or

  (
    g318_n,
    g316_p_spl_,
    g315_p_spl_
  );


  and

  (
    g319_p,
    g318_n,
    g317_n_spl_0
  );


  or

  (
    g319_n,
    g318_p,
    g317_p_spl_0
  );


  and

  (
    g320_p,
    g319_n_spl_,
    g254_n_spl_0
  );


  or

  (
    g320_n,
    g319_p_spl_,
    g254_p_spl_0
  );


  and

  (
    g321_p,
    g319_p_spl_,
    g254_p_spl_
  );


  or

  (
    g321_n,
    g319_n_spl_,
    g254_n_spl_
  );


  and

  (
    g322_p,
    g321_n,
    g320_n_spl_
  );


  or

  (
    g322_n,
    g321_p,
    g320_p_spl_
  );


  and

  (
    g323_p,
    g322_p_spl_,
    g313_n_spl_
  );


  or

  (
    g323_n,
    g322_n_spl_,
    g313_p_spl_
  );


  and

  (
    g324_p,
    g322_n_spl_,
    g313_p_spl_
  );


  or

  (
    g324_n,
    g322_p_spl_,
    g313_n_spl_
  );


  and

  (
    g325_p,
    g324_n,
    g323_n_spl_
  );


  or

  (
    g325_n,
    g324_p,
    g323_p_spl_
  );


  and

  (
    g326_p,
    g325_p_spl_,
    g312_n_spl_
  );


  or

  (
    g326_n,
    g325_n_spl_,
    g312_p_spl_
  );


  and

  (
    g327_p,
    g325_n_spl_,
    g312_p_spl_
  );


  or

  (
    g327_n,
    g325_p_spl_,
    g312_n_spl_
  );


  and

  (
    g328_p,
    g327_n,
    g326_n_spl_
  );


  or

  (
    g328_n,
    g327_p,
    g326_p_spl_
  );


  and

  (
    g329_p,
    g328_p_spl_,
    g311_n_spl_
  );


  or

  (
    g329_n,
    g328_n_spl_,
    g311_p_spl_
  );


  and

  (
    g330_p,
    g328_n_spl_,
    g311_p_spl_
  );


  or

  (
    g330_n,
    g328_p_spl_,
    g311_n_spl_
  );


  and

  (
    g331_p,
    g330_n,
    g329_n_spl_
  );


  or

  (
    g331_n,
    g330_p,
    g329_p_spl_
  );


  and

  (
    g332_p,
    g331_p_spl_,
    g310_n_spl_
  );


  or

  (
    g332_n,
    g331_n_spl_,
    g310_p_spl_
  );


  and

  (
    g333_p,
    g331_n_spl_,
    g310_p_spl_
  );


  or

  (
    g333_n,
    g331_p_spl_,
    g310_n_spl_
  );


  and

  (
    g334_p,
    g333_n,
    g332_n_spl_
  );


  or

  (
    g334_n,
    g333_p,
    g332_p_spl_
  );


  and

  (
    g335_p,
    g334_p_spl_,
    g309_n_spl_
  );


  or

  (
    g335_n,
    g334_n_spl_,
    g309_p_spl_
  );


  and

  (
    g336_p,
    g334_n_spl_,
    g309_p_spl_
  );


  or

  (
    g336_n,
    g334_p_spl_,
    g309_n_spl_
  );


  and

  (
    g337_p,
    g336_n,
    g335_n_spl_
  );


  or

  (
    g337_n,
    g336_p,
    g335_p_spl_
  );


  and

  (
    g338_p,
    g337_p_spl_,
    g308_n_spl_
  );


  or

  (
    g338_n,
    g337_n_spl_,
    g308_p_spl_
  );


  and

  (
    g339_p,
    g337_n_spl_,
    g308_p_spl_
  );


  or

  (
    g339_n,
    g337_p_spl_,
    g308_n_spl_
  );


  and

  (
    g340_p,
    g339_n,
    g338_n_spl_
  );


  or

  (
    g340_n,
    g339_p,
    g338_p_spl_
  );


  and

  (
    g341_p,
    g340_p_spl_,
    g307_n_spl_
  );


  or

  (
    g341_n,
    g340_n_spl_,
    g307_p_spl_
  );


  and

  (
    g342_p,
    g340_n_spl_,
    g307_p_spl_
  );


  or

  (
    g342_n,
    g340_p_spl_,
    g307_n_spl_
  );


  and

  (
    g343_p,
    g342_n,
    g341_n_spl_
  );


  or

  (
    g343_n,
    g342_p,
    g341_p_spl_
  );


  and

  (
    g344_p,
    g343_p_spl_,
    g306_n_spl_
  );


  or

  (
    g344_n,
    g343_n_spl_,
    g306_p_spl_
  );


  and

  (
    g345_p,
    g343_n_spl_,
    g306_p_spl_
  );


  or

  (
    g345_n,
    g343_p_spl_,
    g306_n_spl_
  );


  and

  (
    g346_p,
    g345_n,
    g344_n_spl_
  );


  or

  (
    g346_n,
    g345_p,
    g344_p_spl_
  );


  and

  (
    g347_p,
    g346_p_spl_,
    g305_n_spl_
  );


  or

  (
    g347_n,
    g346_n_spl_,
    g305_p_spl_
  );


  and

  (
    g348_p,
    g346_n_spl_,
    g305_p_spl_
  );


  or

  (
    g348_n,
    g346_p_spl_,
    g305_n_spl_
  );


  and

  (
    g349_p,
    g348_n,
    g347_n_spl_
  );


  or

  (
    g349_n,
    g348_p,
    g347_p_spl_
  );


  and

  (
    g350_p,
    g349_p_spl_,
    g304_n_spl_
  );


  or

  (
    g350_n,
    g349_n_spl_,
    g304_p_spl_
  );


  and

  (
    g351_p,
    g349_n_spl_,
    g304_p_spl_
  );


  or

  (
    g351_n,
    g349_p_spl_,
    g304_n_spl_
  );


  and

  (
    g352_p,
    g351_n,
    g350_n_spl_
  );


  or

  (
    g352_n,
    g351_p,
    g350_p_spl_
  );


  and

  (
    g353_p,
    g352_p_spl_,
    g303_n_spl_
  );


  or

  (
    g353_n,
    g352_n_spl_,
    g303_p_spl_
  );


  and

  (
    g354_p,
    g352_n_spl_,
    g303_p_spl_
  );


  or

  (
    g354_n,
    g352_p_spl_,
    g303_n_spl_
  );


  and

  (
    g355_p,
    g354_n,
    g353_n_spl_
  );


  or

  (
    g355_n,
    g354_p,
    g353_p_spl_
  );


  and

  (
    g356_p,
    g355_p_spl_,
    g302_n_spl_
  );


  or

  (
    g356_n,
    g355_n_spl_,
    g302_p_spl_
  );


  and

  (
    g357_p,
    g355_n_spl_,
    g302_p_spl_
  );


  or

  (
    g357_n,
    g355_p_spl_,
    g302_n_spl_
  );


  and

  (
    g358_p,
    g357_n,
    g356_n_spl_
  );


  or

  (
    g358_n,
    g357_p,
    g356_p_spl_
  );


  and

  (
    g359_p,
    g358_p_spl_,
    g301_n_spl_
  );


  or

  (
    g359_n,
    g358_n_spl_,
    g301_p_spl_
  );


  and

  (
    g360_p,
    g358_n_spl_,
    g301_p_spl_
  );


  or

  (
    g360_n,
    g358_p_spl_,
    g301_n_spl_
  );


  and

  (
    g361_p,
    g360_n,
    g359_n_spl_
  );


  or

  (
    g361_n,
    g360_p,
    g359_p_spl_
  );


  and

  (
    g362_p,
    g361_p_spl_,
    g300_n_spl_
  );


  or

  (
    g362_n,
    g361_n_spl_,
    g300_p_spl_
  );


  and

  (
    g363_p,
    g361_n_spl_,
    g300_p_spl_
  );


  or

  (
    g363_n,
    g361_p_spl_,
    g300_n_spl_
  );


  and

  (
    g364_p,
    g363_n,
    g362_n_spl_
  );


  or

  (
    g364_n,
    g363_p,
    g362_p_spl_
  );


  and

  (
    g365_p,
    g364_p,
    g299_n
  );


  or

  (
    g365_n,
    g364_n_spl_,
    g299_p_spl_
  );


  and

  (
    g366_p,
    g364_n_spl_,
    g299_p_spl_
  );


  or

  (
    g367_n,
    g366_p,
    g365_p_spl_
  );


  and

  (
    g368_p,
    G27_p_spl_000,
    G1_p_spl_101
  );


  or

  (
    g368_n,
    G27_n_spl_000,
    G1_n_spl_100
  );


  and

  (
    g369_p,
    g365_n,
    g362_n_spl_
  );


  or

  (
    g369_n,
    g365_p_spl_,
    g362_p_spl_
  );


  and

  (
    g370_p,
    G26_p_spl_000,
    G2_p_spl_100
  );


  or

  (
    g370_n,
    G26_n_spl_000,
    G2_n_spl_100
  );


  and

  (
    g371_p,
    g359_n_spl_,
    g356_n_spl_
  );


  or

  (
    g371_n,
    g359_p_spl_,
    g356_p_spl_
  );


  and

  (
    g372_p,
    G25_p_spl_001,
    G3_p_spl_100
  );


  or

  (
    g372_n,
    G25_n_spl_001,
    G3_n_spl_100
  );


  and

  (
    g373_p,
    g353_n_spl_,
    g350_n_spl_
  );


  or

  (
    g373_n,
    g353_p_spl_,
    g350_p_spl_
  );


  and

  (
    g374_p,
    G24_p_spl_001,
    G4_p_spl_011
  );


  or

  (
    g374_n,
    G24_n_spl_001,
    G4_n_spl_011
  );


  and

  (
    g375_p,
    g347_n_spl_,
    g344_n_spl_
  );


  or

  (
    g375_n,
    g347_p_spl_,
    g344_p_spl_
  );


  and

  (
    g376_p,
    G23_p_spl_010,
    G5_p_spl_011
  );


  or

  (
    g376_n,
    G23_n_spl_010,
    G5_n_spl_011
  );


  and

  (
    g377_p,
    g341_n_spl_,
    g338_n_spl_
  );


  or

  (
    g377_n,
    g341_p_spl_,
    g338_p_spl_
  );


  and

  (
    g378_p,
    G22_p_spl_010,
    G6_p_spl_010
  );


  or

  (
    g378_n,
    G22_n_spl_010,
    G6_n_spl_010
  );


  and

  (
    g379_p,
    g335_n_spl_,
    g332_n_spl_
  );


  or

  (
    g379_n,
    g335_p_spl_,
    g332_p_spl_
  );


  and

  (
    g380_p,
    G21_p_spl_011,
    G7_p_spl_010
  );


  or

  (
    g380_n,
    G21_n_spl_011,
    G7_n_spl_010
  );


  and

  (
    g381_p,
    g329_n_spl_,
    g326_n_spl_
  );


  or

  (
    g381_n,
    g329_p_spl_,
    g326_p_spl_
  );


  and

  (
    g382_p,
    G20_p_spl_011,
    G8_p_spl_001
  );


  or

  (
    g382_n,
    G20_n_spl_011,
    G8_n_spl_001
  );


  and

  (
    g383_p,
    g323_n_spl_,
    g320_n_spl_
  );


  or

  (
    g383_n,
    g323_p_spl_,
    g320_p_spl_
  );


  and

  (
    g384_p,
    G19_p_spl_100,
    G9_p_spl_001
  );


  or

  (
    g384_n,
    G19_n_spl_100,
    G9_n_spl_001
  );


  and

  (
    g385_p,
    G17_p_spl_101,
    G11_p_spl_000
  );


  or

  (
    g385_n,
    G17_n_spl_100,
    G11_n_spl_000
  );


  and

  (
    g386_p,
    G18_p_spl_100,
    G10_p_spl_000
  );


  or

  (
    g386_n,
    G18_n_spl_100,
    G10_n_spl_000
  );


  and

  (
    g387_p,
    g386_n_spl_,
    g385_p_spl_
  );


  or

  (
    g387_n,
    g386_p_spl_,
    g385_n_spl_
  );


  and

  (
    g388_p,
    g387_n_spl_,
    g385_p_spl_
  );


  or

  (
    g388_n,
    g387_p_spl_,
    g385_n_spl_
  );


  and

  (
    g389_p,
    g387_n_spl_,
    g386_n_spl_
  );


  or

  (
    g389_n,
    g387_p_spl_,
    g386_p_spl_
  );


  and

  (
    g390_p,
    g389_n,
    g388_n_spl_0
  );


  or

  (
    g390_n,
    g389_p,
    g388_p_spl_0
  );


  and

  (
    g391_p,
    g390_n_spl_,
    g317_n_spl_0
  );


  or

  (
    g391_n,
    g390_p_spl_,
    g317_p_spl_0
  );


  and

  (
    g392_p,
    g390_p_spl_,
    g317_p_spl_
  );


  or

  (
    g392_n,
    g390_n_spl_,
    g317_n_spl_
  );


  and

  (
    g393_p,
    g392_n,
    g391_n_spl_
  );


  or

  (
    g393_n,
    g392_p,
    g391_p_spl_
  );


  and

  (
    g394_p,
    g393_p_spl_,
    g384_n_spl_
  );


  or

  (
    g394_n,
    g393_n_spl_,
    g384_p_spl_
  );


  and

  (
    g395_p,
    g393_n_spl_,
    g384_p_spl_
  );


  or

  (
    g395_n,
    g393_p_spl_,
    g384_n_spl_
  );


  and

  (
    g396_p,
    g395_n,
    g394_n_spl_
  );


  or

  (
    g396_n,
    g395_p,
    g394_p_spl_
  );


  and

  (
    g397_p,
    g396_p_spl_,
    g383_n_spl_
  );


  or

  (
    g397_n,
    g396_n_spl_,
    g383_p_spl_
  );


  and

  (
    g398_p,
    g396_n_spl_,
    g383_p_spl_
  );


  or

  (
    g398_n,
    g396_p_spl_,
    g383_n_spl_
  );


  and

  (
    g399_p,
    g398_n,
    g397_n_spl_
  );


  or

  (
    g399_n,
    g398_p,
    g397_p_spl_
  );


  and

  (
    g400_p,
    g399_p_spl_,
    g382_n_spl_
  );


  or

  (
    g400_n,
    g399_n_spl_,
    g382_p_spl_
  );


  and

  (
    g401_p,
    g399_n_spl_,
    g382_p_spl_
  );


  or

  (
    g401_n,
    g399_p_spl_,
    g382_n_spl_
  );


  and

  (
    g402_p,
    g401_n,
    g400_n_spl_
  );


  or

  (
    g402_n,
    g401_p,
    g400_p_spl_
  );


  and

  (
    g403_p,
    g402_p_spl_,
    g381_n_spl_
  );


  or

  (
    g403_n,
    g402_n_spl_,
    g381_p_spl_
  );


  and

  (
    g404_p,
    g402_n_spl_,
    g381_p_spl_
  );


  or

  (
    g404_n,
    g402_p_spl_,
    g381_n_spl_
  );


  and

  (
    g405_p,
    g404_n,
    g403_n_spl_
  );


  or

  (
    g405_n,
    g404_p,
    g403_p_spl_
  );


  and

  (
    g406_p,
    g405_p_spl_,
    g380_n_spl_
  );


  or

  (
    g406_n,
    g405_n_spl_,
    g380_p_spl_
  );


  and

  (
    g407_p,
    g405_n_spl_,
    g380_p_spl_
  );


  or

  (
    g407_n,
    g405_p_spl_,
    g380_n_spl_
  );


  and

  (
    g408_p,
    g407_n,
    g406_n_spl_
  );


  or

  (
    g408_n,
    g407_p,
    g406_p_spl_
  );


  and

  (
    g409_p,
    g408_p_spl_,
    g379_n_spl_
  );


  or

  (
    g409_n,
    g408_n_spl_,
    g379_p_spl_
  );


  and

  (
    g410_p,
    g408_n_spl_,
    g379_p_spl_
  );


  or

  (
    g410_n,
    g408_p_spl_,
    g379_n_spl_
  );


  and

  (
    g411_p,
    g410_n,
    g409_n_spl_
  );


  or

  (
    g411_n,
    g410_p,
    g409_p_spl_
  );


  and

  (
    g412_p,
    g411_p_spl_,
    g378_n_spl_
  );


  or

  (
    g412_n,
    g411_n_spl_,
    g378_p_spl_
  );


  and

  (
    g413_p,
    g411_n_spl_,
    g378_p_spl_
  );


  or

  (
    g413_n,
    g411_p_spl_,
    g378_n_spl_
  );


  and

  (
    g414_p,
    g413_n,
    g412_n_spl_
  );


  or

  (
    g414_n,
    g413_p,
    g412_p_spl_
  );


  and

  (
    g415_p,
    g414_p_spl_,
    g377_n_spl_
  );


  or

  (
    g415_n,
    g414_n_spl_,
    g377_p_spl_
  );


  and

  (
    g416_p,
    g414_n_spl_,
    g377_p_spl_
  );


  or

  (
    g416_n,
    g414_p_spl_,
    g377_n_spl_
  );


  and

  (
    g417_p,
    g416_n,
    g415_n_spl_
  );


  or

  (
    g417_n,
    g416_p,
    g415_p_spl_
  );


  and

  (
    g418_p,
    g417_p_spl_,
    g376_n_spl_
  );


  or

  (
    g418_n,
    g417_n_spl_,
    g376_p_spl_
  );


  and

  (
    g419_p,
    g417_n_spl_,
    g376_p_spl_
  );


  or

  (
    g419_n,
    g417_p_spl_,
    g376_n_spl_
  );


  and

  (
    g420_p,
    g419_n,
    g418_n_spl_
  );


  or

  (
    g420_n,
    g419_p,
    g418_p_spl_
  );


  and

  (
    g421_p,
    g420_p_spl_,
    g375_n_spl_
  );


  or

  (
    g421_n,
    g420_n_spl_,
    g375_p_spl_
  );


  and

  (
    g422_p,
    g420_n_spl_,
    g375_p_spl_
  );


  or

  (
    g422_n,
    g420_p_spl_,
    g375_n_spl_
  );


  and

  (
    g423_p,
    g422_n,
    g421_n_spl_
  );


  or

  (
    g423_n,
    g422_p,
    g421_p_spl_
  );


  and

  (
    g424_p,
    g423_p_spl_,
    g374_n_spl_
  );


  or

  (
    g424_n,
    g423_n_spl_,
    g374_p_spl_
  );


  and

  (
    g425_p,
    g423_n_spl_,
    g374_p_spl_
  );


  or

  (
    g425_n,
    g423_p_spl_,
    g374_n_spl_
  );


  and

  (
    g426_p,
    g425_n,
    g424_n_spl_
  );


  or

  (
    g426_n,
    g425_p,
    g424_p_spl_
  );


  and

  (
    g427_p,
    g426_p_spl_,
    g373_n_spl_
  );


  or

  (
    g427_n,
    g426_n_spl_,
    g373_p_spl_
  );


  and

  (
    g428_p,
    g426_n_spl_,
    g373_p_spl_
  );


  or

  (
    g428_n,
    g426_p_spl_,
    g373_n_spl_
  );


  and

  (
    g429_p,
    g428_n,
    g427_n_spl_
  );


  or

  (
    g429_n,
    g428_p,
    g427_p_spl_
  );


  and

  (
    g430_p,
    g429_p_spl_,
    g372_n_spl_
  );


  or

  (
    g430_n,
    g429_n_spl_,
    g372_p_spl_
  );


  and

  (
    g431_p,
    g429_n_spl_,
    g372_p_spl_
  );


  or

  (
    g431_n,
    g429_p_spl_,
    g372_n_spl_
  );


  and

  (
    g432_p,
    g431_n,
    g430_n_spl_
  );


  or

  (
    g432_n,
    g431_p,
    g430_p_spl_
  );


  and

  (
    g433_p,
    g432_p_spl_,
    g371_n_spl_
  );


  or

  (
    g433_n,
    g432_n_spl_,
    g371_p_spl_
  );


  and

  (
    g434_p,
    g432_n_spl_,
    g371_p_spl_
  );


  or

  (
    g434_n,
    g432_p_spl_,
    g371_n_spl_
  );


  and

  (
    g435_p,
    g434_n,
    g433_n_spl_
  );


  or

  (
    g435_n,
    g434_p,
    g433_p_spl_
  );


  and

  (
    g436_p,
    g435_p_spl_,
    g370_n_spl_
  );


  or

  (
    g436_n,
    g435_n_spl_,
    g370_p_spl_
  );


  and

  (
    g437_p,
    g435_n_spl_,
    g370_p_spl_
  );


  or

  (
    g437_n,
    g435_p_spl_,
    g370_n_spl_
  );


  and

  (
    g438_p,
    g437_n,
    g436_n_spl_
  );


  or

  (
    g438_n,
    g437_p,
    g436_p_spl_
  );


  and

  (
    g439_p,
    g438_p_spl_,
    g369_n_spl_
  );


  or

  (
    g439_n,
    g438_n_spl_,
    g369_p_spl_
  );


  and

  (
    g440_p,
    g438_n_spl_,
    g369_p_spl_
  );


  or

  (
    g440_n,
    g438_p_spl_,
    g369_n_spl_
  );


  and

  (
    g441_p,
    g440_n,
    g439_n_spl_
  );


  or

  (
    g441_n,
    g440_p,
    g439_p_spl_
  );


  and

  (
    g442_p,
    g441_p,
    g368_n
  );


  or

  (
    g442_n,
    g441_n_spl_,
    g368_p_spl_
  );


  and

  (
    g443_p,
    g441_n_spl_,
    g368_p_spl_
  );


  or

  (
    g444_n,
    g443_p,
    g442_p_spl_
  );


  and

  (
    g445_p,
    G28_p_spl_000,
    G1_p_spl_101
  );


  or

  (
    g445_n,
    G28_n_spl_000,
    G1_n_spl_101
  );


  and

  (
    g446_p,
    g442_n,
    g439_n_spl_
  );


  or

  (
    g446_n,
    g442_p_spl_,
    g439_p_spl_
  );


  and

  (
    g447_p,
    G27_p_spl_000,
    G2_p_spl_101
  );


  or

  (
    g447_n,
    G27_n_spl_000,
    G2_n_spl_101
  );


  and

  (
    g448_p,
    g436_n_spl_,
    g433_n_spl_
  );


  or

  (
    g448_n,
    g436_p_spl_,
    g433_p_spl_
  );


  and

  (
    g449_p,
    G26_p_spl_001,
    G3_p_spl_100
  );


  or

  (
    g449_n,
    G26_n_spl_001,
    G3_n_spl_100
  );


  and

  (
    g450_p,
    g430_n_spl_,
    g427_n_spl_
  );


  or

  (
    g450_n,
    g430_p_spl_,
    g427_p_spl_
  );


  and

  (
    g451_p,
    G25_p_spl_001,
    G4_p_spl_100
  );


  or

  (
    g451_n,
    G25_n_spl_001,
    G4_n_spl_100
  );


  and

  (
    g452_p,
    g424_n_spl_,
    g421_n_spl_
  );


  or

  (
    g452_n,
    g424_p_spl_,
    g421_p_spl_
  );


  and

  (
    g453_p,
    G24_p_spl_010,
    G5_p_spl_011
  );


  or

  (
    g453_n,
    G24_n_spl_010,
    G5_n_spl_011
  );


  and

  (
    g454_p,
    g418_n_spl_,
    g415_n_spl_
  );


  or

  (
    g454_n,
    g418_p_spl_,
    g415_p_spl_
  );


  and

  (
    g455_p,
    G23_p_spl_010,
    G6_p_spl_011
  );


  or

  (
    g455_n,
    G23_n_spl_010,
    G6_n_spl_011
  );


  and

  (
    g456_p,
    g412_n_spl_,
    g409_n_spl_
  );


  or

  (
    g456_n,
    g412_p_spl_,
    g409_p_spl_
  );


  and

  (
    g457_p,
    G22_p_spl_011,
    G7_p_spl_010
  );


  or

  (
    g457_n,
    G22_n_spl_011,
    G7_n_spl_010
  );


  and

  (
    g458_p,
    g406_n_spl_,
    g403_n_spl_
  );


  or

  (
    g458_n,
    g406_p_spl_,
    g403_p_spl_
  );


  and

  (
    g459_p,
    G21_p_spl_011,
    G8_p_spl_010
  );


  or

  (
    g459_n,
    G21_n_spl_011,
    G8_n_spl_010
  );


  and

  (
    g460_p,
    g400_n_spl_,
    g397_n_spl_
  );


  or

  (
    g460_n,
    g400_p_spl_,
    g397_p_spl_
  );


  and

  (
    g461_p,
    G20_p_spl_100,
    G9_p_spl_001
  );


  or

  (
    g461_n,
    G20_n_spl_100,
    G9_n_spl_001
  );


  and

  (
    g462_p,
    g394_n_spl_,
    g391_n_spl_
  );


  or

  (
    g462_n,
    g394_p_spl_,
    g391_p_spl_
  );


  and

  (
    g463_p,
    G19_p_spl_100,
    G10_p_spl_001
  );


  or

  (
    g463_n,
    G19_n_spl_100,
    G10_n_spl_001
  );


  and

  (
    g464_p,
    G17_p_spl_101,
    G12_p_spl_000
  );


  or

  (
    g464_n,
    G17_n_spl_101,
    G12_n_spl_000
  );


  and

  (
    g465_p,
    G18_p_spl_101,
    G11_p_spl_000
  );


  or

  (
    g465_n,
    G18_n_spl_101,
    G11_n_spl_000
  );


  and

  (
    g466_p,
    g465_n_spl_,
    g464_p_spl_
  );


  or

  (
    g466_n,
    g465_p_spl_,
    g464_n_spl_
  );


  and

  (
    g467_p,
    g466_n_spl_,
    g464_p_spl_
  );


  or

  (
    g467_n,
    g466_p_spl_,
    g464_n_spl_
  );


  and

  (
    g468_p,
    g466_n_spl_,
    g465_n_spl_
  );


  or

  (
    g468_n,
    g466_p_spl_,
    g465_p_spl_
  );


  and

  (
    g469_p,
    g468_n,
    g467_n_spl_0
  );


  or

  (
    g469_n,
    g468_p,
    g467_p_spl_0
  );


  and

  (
    g470_p,
    g469_n_spl_,
    g388_n_spl_0
  );


  or

  (
    g470_n,
    g469_p_spl_,
    g388_p_spl_0
  );


  and

  (
    g471_p,
    g469_p_spl_,
    g388_p_spl_
  );


  or

  (
    g471_n,
    g469_n_spl_,
    g388_n_spl_
  );


  and

  (
    g472_p,
    g471_n,
    g470_n_spl_
  );


  or

  (
    g472_n,
    g471_p,
    g470_p_spl_
  );


  and

  (
    g473_p,
    g472_p_spl_,
    g463_n_spl_
  );


  or

  (
    g473_n,
    g472_n_spl_,
    g463_p_spl_
  );


  and

  (
    g474_p,
    g472_n_spl_,
    g463_p_spl_
  );


  or

  (
    g474_n,
    g472_p_spl_,
    g463_n_spl_
  );


  and

  (
    g475_p,
    g474_n,
    g473_n_spl_
  );


  or

  (
    g475_n,
    g474_p,
    g473_p_spl_
  );


  and

  (
    g476_p,
    g475_p_spl_,
    g462_n_spl_
  );


  or

  (
    g476_n,
    g475_n_spl_,
    g462_p_spl_
  );


  and

  (
    g477_p,
    g475_n_spl_,
    g462_p_spl_
  );


  or

  (
    g477_n,
    g475_p_spl_,
    g462_n_spl_
  );


  and

  (
    g478_p,
    g477_n,
    g476_n_spl_
  );


  or

  (
    g478_n,
    g477_p,
    g476_p_spl_
  );


  and

  (
    g479_p,
    g478_p_spl_,
    g461_n_spl_
  );


  or

  (
    g479_n,
    g478_n_spl_,
    g461_p_spl_
  );


  and

  (
    g480_p,
    g478_n_spl_,
    g461_p_spl_
  );


  or

  (
    g480_n,
    g478_p_spl_,
    g461_n_spl_
  );


  and

  (
    g481_p,
    g480_n,
    g479_n_spl_
  );


  or

  (
    g481_n,
    g480_p,
    g479_p_spl_
  );


  and

  (
    g482_p,
    g481_p_spl_,
    g460_n_spl_
  );


  or

  (
    g482_n,
    g481_n_spl_,
    g460_p_spl_
  );


  and

  (
    g483_p,
    g481_n_spl_,
    g460_p_spl_
  );


  or

  (
    g483_n,
    g481_p_spl_,
    g460_n_spl_
  );


  and

  (
    g484_p,
    g483_n,
    g482_n_spl_
  );


  or

  (
    g484_n,
    g483_p,
    g482_p_spl_
  );


  and

  (
    g485_p,
    g484_p_spl_,
    g459_n_spl_
  );


  or

  (
    g485_n,
    g484_n_spl_,
    g459_p_spl_
  );


  and

  (
    g486_p,
    g484_n_spl_,
    g459_p_spl_
  );


  or

  (
    g486_n,
    g484_p_spl_,
    g459_n_spl_
  );


  and

  (
    g487_p,
    g486_n,
    g485_n_spl_
  );


  or

  (
    g487_n,
    g486_p,
    g485_p_spl_
  );


  and

  (
    g488_p,
    g487_p_spl_,
    g458_n_spl_
  );


  or

  (
    g488_n,
    g487_n_spl_,
    g458_p_spl_
  );


  and

  (
    g489_p,
    g487_n_spl_,
    g458_p_spl_
  );


  or

  (
    g489_n,
    g487_p_spl_,
    g458_n_spl_
  );


  and

  (
    g490_p,
    g489_n,
    g488_n_spl_
  );


  or

  (
    g490_n,
    g489_p,
    g488_p_spl_
  );


  and

  (
    g491_p,
    g490_p_spl_,
    g457_n_spl_
  );


  or

  (
    g491_n,
    g490_n_spl_,
    g457_p_spl_
  );


  and

  (
    g492_p,
    g490_n_spl_,
    g457_p_spl_
  );


  or

  (
    g492_n,
    g490_p_spl_,
    g457_n_spl_
  );


  and

  (
    g493_p,
    g492_n,
    g491_n_spl_
  );


  or

  (
    g493_n,
    g492_p,
    g491_p_spl_
  );


  and

  (
    g494_p,
    g493_p_spl_,
    g456_n_spl_
  );


  or

  (
    g494_n,
    g493_n_spl_,
    g456_p_spl_
  );


  and

  (
    g495_p,
    g493_n_spl_,
    g456_p_spl_
  );


  or

  (
    g495_n,
    g493_p_spl_,
    g456_n_spl_
  );


  and

  (
    g496_p,
    g495_n,
    g494_n_spl_
  );


  or

  (
    g496_n,
    g495_p,
    g494_p_spl_
  );


  and

  (
    g497_p,
    g496_p_spl_,
    g455_n_spl_
  );


  or

  (
    g497_n,
    g496_n_spl_,
    g455_p_spl_
  );


  and

  (
    g498_p,
    g496_n_spl_,
    g455_p_spl_
  );


  or

  (
    g498_n,
    g496_p_spl_,
    g455_n_spl_
  );


  and

  (
    g499_p,
    g498_n,
    g497_n_spl_
  );


  or

  (
    g499_n,
    g498_p,
    g497_p_spl_
  );


  and

  (
    g500_p,
    g499_p_spl_,
    g454_n_spl_
  );


  or

  (
    g500_n,
    g499_n_spl_,
    g454_p_spl_
  );


  and

  (
    g501_p,
    g499_n_spl_,
    g454_p_spl_
  );


  or

  (
    g501_n,
    g499_p_spl_,
    g454_n_spl_
  );


  and

  (
    g502_p,
    g501_n,
    g500_n_spl_
  );


  or

  (
    g502_n,
    g501_p,
    g500_p_spl_
  );


  and

  (
    g503_p,
    g502_p_spl_,
    g453_n_spl_
  );


  or

  (
    g503_n,
    g502_n_spl_,
    g453_p_spl_
  );


  and

  (
    g504_p,
    g502_n_spl_,
    g453_p_spl_
  );


  or

  (
    g504_n,
    g502_p_spl_,
    g453_n_spl_
  );


  and

  (
    g505_p,
    g504_n,
    g503_n_spl_
  );


  or

  (
    g505_n,
    g504_p,
    g503_p_spl_
  );


  and

  (
    g506_p,
    g505_p_spl_,
    g452_n_spl_
  );


  or

  (
    g506_n,
    g505_n_spl_,
    g452_p_spl_
  );


  and

  (
    g507_p,
    g505_n_spl_,
    g452_p_spl_
  );


  or

  (
    g507_n,
    g505_p_spl_,
    g452_n_spl_
  );


  and

  (
    g508_p,
    g507_n,
    g506_n_spl_
  );


  or

  (
    g508_n,
    g507_p,
    g506_p_spl_
  );


  and

  (
    g509_p,
    g508_p_spl_,
    g451_n_spl_
  );


  or

  (
    g509_n,
    g508_n_spl_,
    g451_p_spl_
  );


  and

  (
    g510_p,
    g508_n_spl_,
    g451_p_spl_
  );


  or

  (
    g510_n,
    g508_p_spl_,
    g451_n_spl_
  );


  and

  (
    g511_p,
    g510_n,
    g509_n_spl_
  );


  or

  (
    g511_n,
    g510_p,
    g509_p_spl_
  );


  and

  (
    g512_p,
    g511_p_spl_,
    g450_n_spl_
  );


  or

  (
    g512_n,
    g511_n_spl_,
    g450_p_spl_
  );


  and

  (
    g513_p,
    g511_n_spl_,
    g450_p_spl_
  );


  or

  (
    g513_n,
    g511_p_spl_,
    g450_n_spl_
  );


  and

  (
    g514_p,
    g513_n,
    g512_n_spl_
  );


  or

  (
    g514_n,
    g513_p,
    g512_p_spl_
  );


  and

  (
    g515_p,
    g514_p_spl_,
    g449_n_spl_
  );


  or

  (
    g515_n,
    g514_n_spl_,
    g449_p_spl_
  );


  and

  (
    g516_p,
    g514_n_spl_,
    g449_p_spl_
  );


  or

  (
    g516_n,
    g514_p_spl_,
    g449_n_spl_
  );


  and

  (
    g517_p,
    g516_n,
    g515_n_spl_
  );


  or

  (
    g517_n,
    g516_p,
    g515_p_spl_
  );


  and

  (
    g518_p,
    g517_p_spl_,
    g448_n_spl_
  );


  or

  (
    g518_n,
    g517_n_spl_,
    g448_p_spl_
  );


  and

  (
    g519_p,
    g517_n_spl_,
    g448_p_spl_
  );


  or

  (
    g519_n,
    g517_p_spl_,
    g448_n_spl_
  );


  and

  (
    g520_p,
    g519_n,
    g518_n_spl_
  );


  or

  (
    g520_n,
    g519_p,
    g518_p_spl_
  );


  and

  (
    g521_p,
    g520_p_spl_,
    g447_n_spl_
  );


  or

  (
    g521_n,
    g520_n_spl_,
    g447_p_spl_
  );


  and

  (
    g522_p,
    g520_n_spl_,
    g447_p_spl_
  );


  or

  (
    g522_n,
    g520_p_spl_,
    g447_n_spl_
  );


  and

  (
    g523_p,
    g522_n,
    g521_n_spl_
  );


  or

  (
    g523_n,
    g522_p,
    g521_p_spl_
  );


  and

  (
    g524_p,
    g523_p_spl_,
    g446_n_spl_
  );


  or

  (
    g524_n,
    g523_n_spl_,
    g446_p_spl_
  );


  and

  (
    g525_p,
    g523_n_spl_,
    g446_p_spl_
  );


  or

  (
    g525_n,
    g523_p_spl_,
    g446_n_spl_
  );


  and

  (
    g526_p,
    g525_n,
    g524_n_spl_
  );


  or

  (
    g526_n,
    g525_p,
    g524_p_spl_
  );


  and

  (
    g527_p,
    g526_p,
    g445_n
  );


  or

  (
    g527_n,
    g526_n_spl_,
    g445_p_spl_
  );


  and

  (
    g528_p,
    g526_n_spl_,
    g445_p_spl_
  );


  or

  (
    g529_n,
    g528_p,
    g527_p_spl_
  );


  and

  (
    g530_p,
    G29_p_spl_000,
    G1_p_spl_110
  );


  or

  (
    g530_n,
    G29_n_spl_000,
    G1_n_spl_101
  );


  and

  (
    g531_p,
    g527_n,
    g524_n_spl_
  );


  or

  (
    g531_n,
    g527_p_spl_,
    g524_p_spl_
  );


  and

  (
    g532_p,
    G28_p_spl_000,
    G2_p_spl_101
  );


  or

  (
    g532_n,
    G28_n_spl_000,
    G2_n_spl_101
  );


  and

  (
    g533_p,
    g521_n_spl_,
    g518_n_spl_
  );


  or

  (
    g533_n,
    g521_p_spl_,
    g518_p_spl_
  );


  and

  (
    g534_p,
    G27_p_spl_001,
    G3_p_spl_101
  );


  or

  (
    g534_n,
    G27_n_spl_001,
    G3_n_spl_101
  );


  and

  (
    g535_p,
    g515_n_spl_,
    g512_n_spl_
  );


  or

  (
    g535_n,
    g515_p_spl_,
    g512_p_spl_
  );


  and

  (
    g536_p,
    G26_p_spl_001,
    G4_p_spl_100
  );


  or

  (
    g536_n,
    G26_n_spl_001,
    G4_n_spl_100
  );


  and

  (
    g537_p,
    g509_n_spl_,
    g506_n_spl_
  );


  or

  (
    g537_n,
    g509_p_spl_,
    g506_p_spl_
  );


  and

  (
    g538_p,
    G25_p_spl_010,
    G5_p_spl_100
  );


  or

  (
    g538_n,
    G25_n_spl_010,
    G5_n_spl_100
  );


  and

  (
    g539_p,
    g503_n_spl_,
    g500_n_spl_
  );


  or

  (
    g539_n,
    g503_p_spl_,
    g500_p_spl_
  );


  and

  (
    g540_p,
    G24_p_spl_010,
    G6_p_spl_011
  );


  or

  (
    g540_n,
    G24_n_spl_010,
    G6_n_spl_011
  );


  and

  (
    g541_p,
    g497_n_spl_,
    g494_n_spl_
  );


  or

  (
    g541_n,
    g497_p_spl_,
    g494_p_spl_
  );


  and

  (
    g542_p,
    G23_p_spl_011,
    G7_p_spl_011
  );


  or

  (
    g542_n,
    G23_n_spl_011,
    G7_n_spl_011
  );


  and

  (
    g543_p,
    g491_n_spl_,
    g488_n_spl_
  );


  or

  (
    g543_n,
    g491_p_spl_,
    g488_p_spl_
  );


  and

  (
    g544_p,
    G22_p_spl_011,
    G8_p_spl_010
  );


  or

  (
    g544_n,
    G22_n_spl_011,
    G8_n_spl_010
  );


  and

  (
    g545_p,
    g485_n_spl_,
    g482_n_spl_
  );


  or

  (
    g545_n,
    g485_p_spl_,
    g482_p_spl_
  );


  and

  (
    g546_p,
    G21_p_spl_100,
    G9_p_spl_010
  );


  or

  (
    g546_n,
    G21_n_spl_100,
    G9_n_spl_010
  );


  and

  (
    g547_p,
    g479_n_spl_,
    g476_n_spl_
  );


  or

  (
    g547_n,
    g479_p_spl_,
    g476_p_spl_
  );


  and

  (
    g548_p,
    G20_p_spl_100,
    G10_p_spl_001
  );


  or

  (
    g548_n,
    G20_n_spl_100,
    G10_n_spl_001
  );


  and

  (
    g549_p,
    g473_n_spl_,
    g470_n_spl_
  );


  or

  (
    g549_n,
    g473_p_spl_,
    g470_p_spl_
  );


  and

  (
    g550_p,
    G19_p_spl_101,
    G11_p_spl_001
  );


  or

  (
    g550_n,
    G19_n_spl_101,
    G11_n_spl_001
  );


  and

  (
    g551_p,
    G17_p_spl_110,
    G13_p_spl_000
  );


  or

  (
    g551_n,
    G17_n_spl_101,
    G13_n_spl_000
  );


  and

  (
    g552_p,
    G18_p_spl_101,
    G12_p_spl_000
  );


  or

  (
    g552_n,
    G18_n_spl_101,
    G12_n_spl_000
  );


  and

  (
    g553_p,
    g552_n_spl_,
    g551_p_spl_
  );


  or

  (
    g553_n,
    g552_p_spl_,
    g551_n_spl_
  );


  and

  (
    g554_p,
    g553_n_spl_,
    g551_p_spl_
  );


  or

  (
    g554_n,
    g553_p_spl_,
    g551_n_spl_
  );


  and

  (
    g555_p,
    g553_n_spl_,
    g552_n_spl_
  );


  or

  (
    g555_n,
    g553_p_spl_,
    g552_p_spl_
  );


  and

  (
    g556_p,
    g555_n,
    g554_n_spl_0
  );


  or

  (
    g556_n,
    g555_p,
    g554_p_spl_0
  );


  and

  (
    g557_p,
    g556_n_spl_,
    g467_n_spl_0
  );


  or

  (
    g557_n,
    g556_p_spl_,
    g467_p_spl_0
  );


  and

  (
    g558_p,
    g556_p_spl_,
    g467_p_spl_
  );


  or

  (
    g558_n,
    g556_n_spl_,
    g467_n_spl_
  );


  and

  (
    g559_p,
    g558_n,
    g557_n_spl_
  );


  or

  (
    g559_n,
    g558_p,
    g557_p_spl_
  );


  and

  (
    g560_p,
    g559_p_spl_,
    g550_n_spl_
  );


  or

  (
    g560_n,
    g559_n_spl_,
    g550_p_spl_
  );


  and

  (
    g561_p,
    g559_n_spl_,
    g550_p_spl_
  );


  or

  (
    g561_n,
    g559_p_spl_,
    g550_n_spl_
  );


  and

  (
    g562_p,
    g561_n,
    g560_n_spl_
  );


  or

  (
    g562_n,
    g561_p,
    g560_p_spl_
  );


  and

  (
    g563_p,
    g562_p_spl_,
    g549_n_spl_
  );


  or

  (
    g563_n,
    g562_n_spl_,
    g549_p_spl_
  );


  and

  (
    g564_p,
    g562_n_spl_,
    g549_p_spl_
  );


  or

  (
    g564_n,
    g562_p_spl_,
    g549_n_spl_
  );


  and

  (
    g565_p,
    g564_n,
    g563_n_spl_
  );


  or

  (
    g565_n,
    g564_p,
    g563_p_spl_
  );


  and

  (
    g566_p,
    g565_p_spl_,
    g548_n_spl_
  );


  or

  (
    g566_n,
    g565_n_spl_,
    g548_p_spl_
  );


  and

  (
    g567_p,
    g565_n_spl_,
    g548_p_spl_
  );


  or

  (
    g567_n,
    g565_p_spl_,
    g548_n_spl_
  );


  and

  (
    g568_p,
    g567_n,
    g566_n_spl_
  );


  or

  (
    g568_n,
    g567_p,
    g566_p_spl_
  );


  and

  (
    g569_p,
    g568_p_spl_,
    g547_n_spl_
  );


  or

  (
    g569_n,
    g568_n_spl_,
    g547_p_spl_
  );


  and

  (
    g570_p,
    g568_n_spl_,
    g547_p_spl_
  );


  or

  (
    g570_n,
    g568_p_spl_,
    g547_n_spl_
  );


  and

  (
    g571_p,
    g570_n,
    g569_n_spl_
  );


  or

  (
    g571_n,
    g570_p,
    g569_p_spl_
  );


  and

  (
    g572_p,
    g571_p_spl_,
    g546_n_spl_
  );


  or

  (
    g572_n,
    g571_n_spl_,
    g546_p_spl_
  );


  and

  (
    g573_p,
    g571_n_spl_,
    g546_p_spl_
  );


  or

  (
    g573_n,
    g571_p_spl_,
    g546_n_spl_
  );


  and

  (
    g574_p,
    g573_n,
    g572_n_spl_
  );


  or

  (
    g574_n,
    g573_p,
    g572_p_spl_
  );


  and

  (
    g575_p,
    g574_p_spl_,
    g545_n_spl_
  );


  or

  (
    g575_n,
    g574_n_spl_,
    g545_p_spl_
  );


  and

  (
    g576_p,
    g574_n_spl_,
    g545_p_spl_
  );


  or

  (
    g576_n,
    g574_p_spl_,
    g545_n_spl_
  );


  and

  (
    g577_p,
    g576_n,
    g575_n_spl_
  );


  or

  (
    g577_n,
    g576_p,
    g575_p_spl_
  );


  and

  (
    g578_p,
    g577_p_spl_,
    g544_n_spl_
  );


  or

  (
    g578_n,
    g577_n_spl_,
    g544_p_spl_
  );


  and

  (
    g579_p,
    g577_n_spl_,
    g544_p_spl_
  );


  or

  (
    g579_n,
    g577_p_spl_,
    g544_n_spl_
  );


  and

  (
    g580_p,
    g579_n,
    g578_n_spl_
  );


  or

  (
    g580_n,
    g579_p,
    g578_p_spl_
  );


  and

  (
    g581_p,
    g580_p_spl_,
    g543_n_spl_
  );


  or

  (
    g581_n,
    g580_n_spl_,
    g543_p_spl_
  );


  and

  (
    g582_p,
    g580_n_spl_,
    g543_p_spl_
  );


  or

  (
    g582_n,
    g580_p_spl_,
    g543_n_spl_
  );


  and

  (
    g583_p,
    g582_n,
    g581_n_spl_
  );


  or

  (
    g583_n,
    g582_p,
    g581_p_spl_
  );


  and

  (
    g584_p,
    g583_p_spl_,
    g542_n_spl_
  );


  or

  (
    g584_n,
    g583_n_spl_,
    g542_p_spl_
  );


  and

  (
    g585_p,
    g583_n_spl_,
    g542_p_spl_
  );


  or

  (
    g585_n,
    g583_p_spl_,
    g542_n_spl_
  );


  and

  (
    g586_p,
    g585_n,
    g584_n_spl_
  );


  or

  (
    g586_n,
    g585_p,
    g584_p_spl_
  );


  and

  (
    g587_p,
    g586_p_spl_,
    g541_n_spl_
  );


  or

  (
    g587_n,
    g586_n_spl_,
    g541_p_spl_
  );


  and

  (
    g588_p,
    g586_n_spl_,
    g541_p_spl_
  );


  or

  (
    g588_n,
    g586_p_spl_,
    g541_n_spl_
  );


  and

  (
    g589_p,
    g588_n,
    g587_n_spl_
  );


  or

  (
    g589_n,
    g588_p,
    g587_p_spl_
  );


  and

  (
    g590_p,
    g589_p_spl_,
    g540_n_spl_
  );


  or

  (
    g590_n,
    g589_n_spl_,
    g540_p_spl_
  );


  and

  (
    g591_p,
    g589_n_spl_,
    g540_p_spl_
  );


  or

  (
    g591_n,
    g589_p_spl_,
    g540_n_spl_
  );


  and

  (
    g592_p,
    g591_n,
    g590_n_spl_
  );


  or

  (
    g592_n,
    g591_p,
    g590_p_spl_
  );


  and

  (
    g593_p,
    g592_p_spl_,
    g539_n_spl_
  );


  or

  (
    g593_n,
    g592_n_spl_,
    g539_p_spl_
  );


  and

  (
    g594_p,
    g592_n_spl_,
    g539_p_spl_
  );


  or

  (
    g594_n,
    g592_p_spl_,
    g539_n_spl_
  );


  and

  (
    g595_p,
    g594_n,
    g593_n_spl_
  );


  or

  (
    g595_n,
    g594_p,
    g593_p_spl_
  );


  and

  (
    g596_p,
    g595_p_spl_,
    g538_n_spl_
  );


  or

  (
    g596_n,
    g595_n_spl_,
    g538_p_spl_
  );


  and

  (
    g597_p,
    g595_n_spl_,
    g538_p_spl_
  );


  or

  (
    g597_n,
    g595_p_spl_,
    g538_n_spl_
  );


  and

  (
    g598_p,
    g597_n,
    g596_n_spl_
  );


  or

  (
    g598_n,
    g597_p,
    g596_p_spl_
  );


  and

  (
    g599_p,
    g598_p_spl_,
    g537_n_spl_
  );


  or

  (
    g599_n,
    g598_n_spl_,
    g537_p_spl_
  );


  and

  (
    g600_p,
    g598_n_spl_,
    g537_p_spl_
  );


  or

  (
    g600_n,
    g598_p_spl_,
    g537_n_spl_
  );


  and

  (
    g601_p,
    g600_n,
    g599_n_spl_
  );


  or

  (
    g601_n,
    g600_p,
    g599_p_spl_
  );


  and

  (
    g602_p,
    g601_p_spl_,
    g536_n_spl_
  );


  or

  (
    g602_n,
    g601_n_spl_,
    g536_p_spl_
  );


  and

  (
    g603_p,
    g601_n_spl_,
    g536_p_spl_
  );


  or

  (
    g603_n,
    g601_p_spl_,
    g536_n_spl_
  );


  and

  (
    g604_p,
    g603_n,
    g602_n_spl_
  );


  or

  (
    g604_n,
    g603_p,
    g602_p_spl_
  );


  and

  (
    g605_p,
    g604_p_spl_,
    g535_n_spl_
  );


  or

  (
    g605_n,
    g604_n_spl_,
    g535_p_spl_
  );


  and

  (
    g606_p,
    g604_n_spl_,
    g535_p_spl_
  );


  or

  (
    g606_n,
    g604_p_spl_,
    g535_n_spl_
  );


  and

  (
    g607_p,
    g606_n,
    g605_n_spl_
  );


  or

  (
    g607_n,
    g606_p,
    g605_p_spl_
  );


  and

  (
    g608_p,
    g607_p_spl_,
    g534_n_spl_
  );


  or

  (
    g608_n,
    g607_n_spl_,
    g534_p_spl_
  );


  and

  (
    g609_p,
    g607_n_spl_,
    g534_p_spl_
  );


  or

  (
    g609_n,
    g607_p_spl_,
    g534_n_spl_
  );


  and

  (
    g610_p,
    g609_n,
    g608_n_spl_
  );


  or

  (
    g610_n,
    g609_p,
    g608_p_spl_
  );


  and

  (
    g611_p,
    g610_p_spl_,
    g533_n_spl_
  );


  or

  (
    g611_n,
    g610_n_spl_,
    g533_p_spl_
  );


  and

  (
    g612_p,
    g610_n_spl_,
    g533_p_spl_
  );


  or

  (
    g612_n,
    g610_p_spl_,
    g533_n_spl_
  );


  and

  (
    g613_p,
    g612_n,
    g611_n_spl_
  );


  or

  (
    g613_n,
    g612_p,
    g611_p_spl_
  );


  and

  (
    g614_p,
    g613_p_spl_,
    g532_n_spl_
  );


  or

  (
    g614_n,
    g613_n_spl_,
    g532_p_spl_
  );


  and

  (
    g615_p,
    g613_n_spl_,
    g532_p_spl_
  );


  or

  (
    g615_n,
    g613_p_spl_,
    g532_n_spl_
  );


  and

  (
    g616_p,
    g615_n,
    g614_n_spl_
  );


  or

  (
    g616_n,
    g615_p,
    g614_p_spl_
  );


  and

  (
    g617_p,
    g616_p_spl_,
    g531_n_spl_
  );


  or

  (
    g617_n,
    g616_n_spl_,
    g531_p_spl_
  );


  and

  (
    g618_p,
    g616_n_spl_,
    g531_p_spl_
  );


  or

  (
    g618_n,
    g616_p_spl_,
    g531_n_spl_
  );


  and

  (
    g619_p,
    g618_n,
    g617_n_spl_
  );


  or

  (
    g619_n,
    g618_p,
    g617_p_spl_
  );


  and

  (
    g620_p,
    g619_p,
    g530_n
  );


  or

  (
    g620_n,
    g619_n_spl_,
    g530_p_spl_
  );


  and

  (
    g621_p,
    g619_n_spl_,
    g530_p_spl_
  );


  or

  (
    g622_n,
    g621_p,
    g620_p_spl_
  );


  and

  (
    g623_p,
    G30_p_spl_000,
    G1_p_spl_110
  );


  or

  (
    g623_n,
    G30_n_spl_000,
    G1_n_spl_110
  );


  and

  (
    g624_p,
    g620_n,
    g617_n_spl_
  );


  or

  (
    g624_n,
    g620_p_spl_,
    g617_p_spl_
  );


  and

  (
    g625_p,
    G29_p_spl_000,
    G2_p_spl_110
  );


  or

  (
    g625_n,
    G29_n_spl_000,
    G2_n_spl_110
  );


  and

  (
    g626_p,
    g614_n_spl_,
    g611_n_spl_
  );


  or

  (
    g626_n,
    g614_p_spl_,
    g611_p_spl_
  );


  and

  (
    g627_p,
    G28_p_spl_001,
    G3_p_spl_101
  );


  or

  (
    g627_n,
    G28_n_spl_001,
    G3_n_spl_101
  );


  and

  (
    g628_p,
    g608_n_spl_,
    g605_n_spl_
  );


  or

  (
    g628_n,
    g608_p_spl_,
    g605_p_spl_
  );


  and

  (
    g629_p,
    G27_p_spl_001,
    G4_p_spl_101
  );


  or

  (
    g629_n,
    G27_n_spl_001,
    G4_n_spl_101
  );


  and

  (
    g630_p,
    g602_n_spl_,
    g599_n_spl_
  );


  or

  (
    g630_n,
    g602_p_spl_,
    g599_p_spl_
  );


  and

  (
    g631_p,
    G26_p_spl_010,
    G5_p_spl_100
  );


  or

  (
    g631_n,
    G26_n_spl_010,
    G5_n_spl_100
  );


  and

  (
    g632_p,
    g596_n_spl_,
    g593_n_spl_
  );


  or

  (
    g632_n,
    g596_p_spl_,
    g593_p_spl_
  );


  and

  (
    g633_p,
    G25_p_spl_010,
    G6_p_spl_100
  );


  or

  (
    g633_n,
    G25_n_spl_010,
    G6_n_spl_100
  );


  and

  (
    g634_p,
    g590_n_spl_,
    g587_n_spl_
  );


  or

  (
    g634_n,
    g590_p_spl_,
    g587_p_spl_
  );


  and

  (
    g635_p,
    G24_p_spl_011,
    G7_p_spl_011
  );


  or

  (
    g635_n,
    G24_n_spl_011,
    G7_n_spl_011
  );


  and

  (
    g636_p,
    g584_n_spl_,
    g581_n_spl_
  );


  or

  (
    g636_n,
    g584_p_spl_,
    g581_p_spl_
  );


  and

  (
    g637_p,
    G23_p_spl_011,
    G8_p_spl_011
  );


  or

  (
    g637_n,
    G23_n_spl_011,
    G8_n_spl_011
  );


  and

  (
    g638_p,
    g578_n_spl_,
    g575_n_spl_
  );


  or

  (
    g638_n,
    g578_p_spl_,
    g575_p_spl_
  );


  and

  (
    g639_p,
    G22_p_spl_100,
    G9_p_spl_010
  );


  or

  (
    g639_n,
    G22_n_spl_100,
    G9_n_spl_010
  );


  and

  (
    g640_p,
    g572_n_spl_,
    g569_n_spl_
  );


  or

  (
    g640_n,
    g572_p_spl_,
    g569_p_spl_
  );


  and

  (
    g641_p,
    G21_p_spl_100,
    G10_p_spl_010
  );


  or

  (
    g641_n,
    G21_n_spl_100,
    G10_n_spl_010
  );


  and

  (
    g642_p,
    g566_n_spl_,
    g563_n_spl_
  );


  or

  (
    g642_n,
    g566_p_spl_,
    g563_p_spl_
  );


  and

  (
    g643_p,
    G20_p_spl_101,
    G11_p_spl_001
  );


  or

  (
    g643_n,
    G20_n_spl_101,
    G11_n_spl_001
  );


  and

  (
    g644_p,
    g560_n_spl_,
    g557_n_spl_
  );


  or

  (
    g644_n,
    g560_p_spl_,
    g557_p_spl_
  );


  and

  (
    g645_p,
    G19_p_spl_101,
    G12_p_spl_001
  );


  or

  (
    g645_n,
    G19_n_spl_101,
    G12_n_spl_001
  );


  and

  (
    g646_p,
    G17_p_spl_110,
    G14_p_spl_000
  );


  or

  (
    g646_n,
    G17_n_spl_110,
    G14_n_spl_000
  );


  and

  (
    g647_p,
    G18_p_spl_110,
    G13_p_spl_000
  );


  or

  (
    g647_n,
    G18_n_spl_110,
    G13_n_spl_000
  );


  and

  (
    g648_p,
    g647_n_spl_,
    g646_p_spl_
  );


  or

  (
    g648_n,
    g647_p_spl_,
    g646_n_spl_
  );


  and

  (
    g649_p,
    g648_n_spl_,
    g646_p_spl_
  );


  or

  (
    g649_n,
    g648_p_spl_,
    g646_n_spl_
  );


  and

  (
    g650_p,
    g648_n_spl_,
    g647_n_spl_
  );


  or

  (
    g650_n,
    g648_p_spl_,
    g647_p_spl_
  );


  and

  (
    g651_p,
    g650_n,
    g649_n_spl_0
  );


  or

  (
    g651_n,
    g650_p,
    g649_p_spl_0
  );


  and

  (
    g652_p,
    g651_n_spl_,
    g554_n_spl_0
  );


  or

  (
    g652_n,
    g651_p_spl_,
    g554_p_spl_0
  );


  and

  (
    g653_p,
    g651_p_spl_,
    g554_p_spl_
  );


  or

  (
    g653_n,
    g651_n_spl_,
    g554_n_spl_
  );


  and

  (
    g654_p,
    g653_n,
    g652_n_spl_
  );


  or

  (
    g654_n,
    g653_p,
    g652_p_spl_
  );


  and

  (
    g655_p,
    g654_p_spl_,
    g645_n_spl_
  );


  or

  (
    g655_n,
    g654_n_spl_,
    g645_p_spl_
  );


  and

  (
    g656_p,
    g654_n_spl_,
    g645_p_spl_
  );


  or

  (
    g656_n,
    g654_p_spl_,
    g645_n_spl_
  );


  and

  (
    g657_p,
    g656_n,
    g655_n_spl_
  );


  or

  (
    g657_n,
    g656_p,
    g655_p_spl_
  );


  and

  (
    g658_p,
    g657_p_spl_,
    g644_n_spl_
  );


  or

  (
    g658_n,
    g657_n_spl_,
    g644_p_spl_
  );


  and

  (
    g659_p,
    g657_n_spl_,
    g644_p_spl_
  );


  or

  (
    g659_n,
    g657_p_spl_,
    g644_n_spl_
  );


  and

  (
    g660_p,
    g659_n,
    g658_n_spl_
  );


  or

  (
    g660_n,
    g659_p,
    g658_p_spl_
  );


  and

  (
    g661_p,
    g660_p_spl_,
    g643_n_spl_
  );


  or

  (
    g661_n,
    g660_n_spl_,
    g643_p_spl_
  );


  and

  (
    g662_p,
    g660_n_spl_,
    g643_p_spl_
  );


  or

  (
    g662_n,
    g660_p_spl_,
    g643_n_spl_
  );


  and

  (
    g663_p,
    g662_n,
    g661_n_spl_
  );


  or

  (
    g663_n,
    g662_p,
    g661_p_spl_
  );


  and

  (
    g664_p,
    g663_p_spl_,
    g642_n_spl_
  );


  or

  (
    g664_n,
    g663_n_spl_,
    g642_p_spl_
  );


  and

  (
    g665_p,
    g663_n_spl_,
    g642_p_spl_
  );


  or

  (
    g665_n,
    g663_p_spl_,
    g642_n_spl_
  );


  and

  (
    g666_p,
    g665_n,
    g664_n_spl_
  );


  or

  (
    g666_n,
    g665_p,
    g664_p_spl_
  );


  and

  (
    g667_p,
    g666_p_spl_,
    g641_n_spl_
  );


  or

  (
    g667_n,
    g666_n_spl_,
    g641_p_spl_
  );


  and

  (
    g668_p,
    g666_n_spl_,
    g641_p_spl_
  );


  or

  (
    g668_n,
    g666_p_spl_,
    g641_n_spl_
  );


  and

  (
    g669_p,
    g668_n,
    g667_n_spl_
  );


  or

  (
    g669_n,
    g668_p,
    g667_p_spl_
  );


  and

  (
    g670_p,
    g669_p_spl_,
    g640_n_spl_
  );


  or

  (
    g670_n,
    g669_n_spl_,
    g640_p_spl_
  );


  and

  (
    g671_p,
    g669_n_spl_,
    g640_p_spl_
  );


  or

  (
    g671_n,
    g669_p_spl_,
    g640_n_spl_
  );


  and

  (
    g672_p,
    g671_n,
    g670_n_spl_
  );


  or

  (
    g672_n,
    g671_p,
    g670_p_spl_
  );


  and

  (
    g673_p,
    g672_p_spl_,
    g639_n_spl_
  );


  or

  (
    g673_n,
    g672_n_spl_,
    g639_p_spl_
  );


  and

  (
    g674_p,
    g672_n_spl_,
    g639_p_spl_
  );


  or

  (
    g674_n,
    g672_p_spl_,
    g639_n_spl_
  );


  and

  (
    g675_p,
    g674_n,
    g673_n_spl_
  );


  or

  (
    g675_n,
    g674_p,
    g673_p_spl_
  );


  and

  (
    g676_p,
    g675_p_spl_,
    g638_n_spl_
  );


  or

  (
    g676_n,
    g675_n_spl_,
    g638_p_spl_
  );


  and

  (
    g677_p,
    g675_n_spl_,
    g638_p_spl_
  );


  or

  (
    g677_n,
    g675_p_spl_,
    g638_n_spl_
  );


  and

  (
    g678_p,
    g677_n,
    g676_n_spl_
  );


  or

  (
    g678_n,
    g677_p,
    g676_p_spl_
  );


  and

  (
    g679_p,
    g678_p_spl_,
    g637_n_spl_
  );


  or

  (
    g679_n,
    g678_n_spl_,
    g637_p_spl_
  );


  and

  (
    g680_p,
    g678_n_spl_,
    g637_p_spl_
  );


  or

  (
    g680_n,
    g678_p_spl_,
    g637_n_spl_
  );


  and

  (
    g681_p,
    g680_n,
    g679_n_spl_
  );


  or

  (
    g681_n,
    g680_p,
    g679_p_spl_
  );


  and

  (
    g682_p,
    g681_p_spl_,
    g636_n_spl_
  );


  or

  (
    g682_n,
    g681_n_spl_,
    g636_p_spl_
  );


  and

  (
    g683_p,
    g681_n_spl_,
    g636_p_spl_
  );


  or

  (
    g683_n,
    g681_p_spl_,
    g636_n_spl_
  );


  and

  (
    g684_p,
    g683_n,
    g682_n_spl_
  );


  or

  (
    g684_n,
    g683_p,
    g682_p_spl_
  );


  and

  (
    g685_p,
    g684_p_spl_,
    g635_n_spl_
  );


  or

  (
    g685_n,
    g684_n_spl_,
    g635_p_spl_
  );


  and

  (
    g686_p,
    g684_n_spl_,
    g635_p_spl_
  );


  or

  (
    g686_n,
    g684_p_spl_,
    g635_n_spl_
  );


  and

  (
    g687_p,
    g686_n,
    g685_n_spl_
  );


  or

  (
    g687_n,
    g686_p,
    g685_p_spl_
  );


  and

  (
    g688_p,
    g687_p_spl_,
    g634_n_spl_
  );


  or

  (
    g688_n,
    g687_n_spl_,
    g634_p_spl_
  );


  and

  (
    g689_p,
    g687_n_spl_,
    g634_p_spl_
  );


  or

  (
    g689_n,
    g687_p_spl_,
    g634_n_spl_
  );


  and

  (
    g690_p,
    g689_n,
    g688_n_spl_
  );


  or

  (
    g690_n,
    g689_p,
    g688_p_spl_
  );


  and

  (
    g691_p,
    g690_p_spl_,
    g633_n_spl_
  );


  or

  (
    g691_n,
    g690_n_spl_,
    g633_p_spl_
  );


  and

  (
    g692_p,
    g690_n_spl_,
    g633_p_spl_
  );


  or

  (
    g692_n,
    g690_p_spl_,
    g633_n_spl_
  );


  and

  (
    g693_p,
    g692_n,
    g691_n_spl_
  );


  or

  (
    g693_n,
    g692_p,
    g691_p_spl_
  );


  and

  (
    g694_p,
    g693_p_spl_,
    g632_n_spl_
  );


  or

  (
    g694_n,
    g693_n_spl_,
    g632_p_spl_
  );


  and

  (
    g695_p,
    g693_n_spl_,
    g632_p_spl_
  );


  or

  (
    g695_n,
    g693_p_spl_,
    g632_n_spl_
  );


  and

  (
    g696_p,
    g695_n,
    g694_n_spl_
  );


  or

  (
    g696_n,
    g695_p,
    g694_p_spl_
  );


  and

  (
    g697_p,
    g696_p_spl_,
    g631_n_spl_
  );


  or

  (
    g697_n,
    g696_n_spl_,
    g631_p_spl_
  );


  and

  (
    g698_p,
    g696_n_spl_,
    g631_p_spl_
  );


  or

  (
    g698_n,
    g696_p_spl_,
    g631_n_spl_
  );


  and

  (
    g699_p,
    g698_n,
    g697_n_spl_
  );


  or

  (
    g699_n,
    g698_p,
    g697_p_spl_
  );


  and

  (
    g700_p,
    g699_p_spl_,
    g630_n_spl_
  );


  or

  (
    g700_n,
    g699_n_spl_,
    g630_p_spl_
  );


  and

  (
    g701_p,
    g699_n_spl_,
    g630_p_spl_
  );


  or

  (
    g701_n,
    g699_p_spl_,
    g630_n_spl_
  );


  and

  (
    g702_p,
    g701_n,
    g700_n_spl_
  );


  or

  (
    g702_n,
    g701_p,
    g700_p_spl_
  );


  and

  (
    g703_p,
    g702_p_spl_,
    g629_n_spl_
  );


  or

  (
    g703_n,
    g702_n_spl_,
    g629_p_spl_
  );


  and

  (
    g704_p,
    g702_n_spl_,
    g629_p_spl_
  );


  or

  (
    g704_n,
    g702_p_spl_,
    g629_n_spl_
  );


  and

  (
    g705_p,
    g704_n,
    g703_n_spl_
  );


  or

  (
    g705_n,
    g704_p,
    g703_p_spl_
  );


  and

  (
    g706_p,
    g705_p_spl_,
    g628_n_spl_
  );


  or

  (
    g706_n,
    g705_n_spl_,
    g628_p_spl_
  );


  and

  (
    g707_p,
    g705_n_spl_,
    g628_p_spl_
  );


  or

  (
    g707_n,
    g705_p_spl_,
    g628_n_spl_
  );


  and

  (
    g708_p,
    g707_n,
    g706_n_spl_
  );


  or

  (
    g708_n,
    g707_p,
    g706_p_spl_
  );


  and

  (
    g709_p,
    g708_p_spl_,
    g627_n_spl_
  );


  or

  (
    g709_n,
    g708_n_spl_,
    g627_p_spl_
  );


  and

  (
    g710_p,
    g708_n_spl_,
    g627_p_spl_
  );


  or

  (
    g710_n,
    g708_p_spl_,
    g627_n_spl_
  );


  and

  (
    g711_p,
    g710_n,
    g709_n_spl_
  );


  or

  (
    g711_n,
    g710_p,
    g709_p_spl_
  );


  and

  (
    g712_p,
    g711_p_spl_,
    g626_n_spl_
  );


  or

  (
    g712_n,
    g711_n_spl_,
    g626_p_spl_
  );


  and

  (
    g713_p,
    g711_n_spl_,
    g626_p_spl_
  );


  or

  (
    g713_n,
    g711_p_spl_,
    g626_n_spl_
  );


  and

  (
    g714_p,
    g713_n,
    g712_n_spl_
  );


  or

  (
    g714_n,
    g713_p,
    g712_p_spl_
  );


  and

  (
    g715_p,
    g714_p_spl_,
    g625_n_spl_
  );


  or

  (
    g715_n,
    g714_n_spl_,
    g625_p_spl_
  );


  and

  (
    g716_p,
    g714_n_spl_,
    g625_p_spl_
  );


  or

  (
    g716_n,
    g714_p_spl_,
    g625_n_spl_
  );


  and

  (
    g717_p,
    g716_n,
    g715_n_spl_
  );


  or

  (
    g717_n,
    g716_p,
    g715_p_spl_
  );


  and

  (
    g718_p,
    g717_p_spl_,
    g624_n_spl_
  );


  or

  (
    g718_n,
    g717_n_spl_,
    g624_p_spl_
  );


  and

  (
    g719_p,
    g717_n_spl_,
    g624_p_spl_
  );


  or

  (
    g719_n,
    g717_p_spl_,
    g624_n_spl_
  );


  and

  (
    g720_p,
    g719_n,
    g718_n_spl_
  );


  or

  (
    g720_n,
    g719_p,
    g718_p_spl_
  );


  and

  (
    g721_p,
    g720_p,
    g623_n
  );


  or

  (
    g721_n,
    g720_n_spl_,
    g623_p_spl_
  );


  and

  (
    g722_p,
    g720_n_spl_,
    g623_p_spl_
  );


  or

  (
    g723_n,
    g722_p,
    g721_p_spl_
  );


  and

  (
    g724_p,
    G31_p_spl_000,
    G1_p_spl_111
  );


  or

  (
    g724_n,
    G31_n_spl_000,
    G1_n_spl_110
  );


  and

  (
    g725_p,
    g721_n,
    g718_n_spl_
  );


  or

  (
    g725_n,
    g721_p_spl_,
    g718_p_spl_
  );


  and

  (
    g726_p,
    G30_p_spl_000,
    G2_p_spl_110
  );


  or

  (
    g726_n,
    G30_n_spl_000,
    G2_n_spl_110
  );


  and

  (
    g727_p,
    g715_n_spl_,
    g712_n_spl_
  );


  or

  (
    g727_n,
    g715_p_spl_,
    g712_p_spl_
  );


  and

  (
    g728_p,
    G29_p_spl_001,
    G3_p_spl_110
  );


  or

  (
    g728_n,
    G29_n_spl_001,
    G3_n_spl_110
  );


  and

  (
    g729_p,
    g709_n_spl_,
    g706_n_spl_
  );


  or

  (
    g729_n,
    g709_p_spl_,
    g706_p_spl_
  );


  and

  (
    g730_p,
    G28_p_spl_001,
    G4_p_spl_101
  );


  or

  (
    g730_n,
    G28_n_spl_001,
    G4_n_spl_101
  );


  and

  (
    g731_p,
    g703_n_spl_,
    g700_n_spl_
  );


  or

  (
    g731_n,
    g703_p_spl_,
    g700_p_spl_
  );


  and

  (
    g732_p,
    G27_p_spl_010,
    G5_p_spl_101
  );


  or

  (
    g732_n,
    G27_n_spl_010,
    G5_n_spl_101
  );


  and

  (
    g733_p,
    g697_n_spl_,
    g694_n_spl_
  );


  or

  (
    g733_n,
    g697_p_spl_,
    g694_p_spl_
  );


  and

  (
    g734_p,
    G26_p_spl_010,
    G6_p_spl_100
  );


  or

  (
    g734_n,
    G26_n_spl_010,
    G6_n_spl_100
  );


  and

  (
    g735_p,
    g691_n_spl_,
    g688_n_spl_
  );


  or

  (
    g735_n,
    g691_p_spl_,
    g688_p_spl_
  );


  and

  (
    g736_p,
    G25_p_spl_011,
    G7_p_spl_100
  );


  or

  (
    g736_n,
    G25_n_spl_011,
    G7_n_spl_100
  );


  and

  (
    g737_p,
    g685_n_spl_,
    g682_n_spl_
  );


  or

  (
    g737_n,
    g685_p_spl_,
    g682_p_spl_
  );


  and

  (
    g738_p,
    G24_p_spl_011,
    G8_p_spl_011
  );


  or

  (
    g738_n,
    G24_n_spl_011,
    G8_n_spl_011
  );


  and

  (
    g739_p,
    g679_n_spl_,
    g676_n_spl_
  );


  or

  (
    g739_n,
    g679_p_spl_,
    g676_p_spl_
  );


  and

  (
    g740_p,
    G23_p_spl_100,
    G9_p_spl_011
  );


  or

  (
    g740_n,
    G23_n_spl_100,
    G9_n_spl_011
  );


  and

  (
    g741_p,
    g673_n_spl_,
    g670_n_spl_
  );


  or

  (
    g741_n,
    g673_p_spl_,
    g670_p_spl_
  );


  and

  (
    g742_p,
    G22_p_spl_100,
    G10_p_spl_010
  );


  or

  (
    g742_n,
    G22_n_spl_100,
    G10_n_spl_010
  );


  and

  (
    g743_p,
    g667_n_spl_,
    g664_n_spl_
  );


  or

  (
    g743_n,
    g667_p_spl_,
    g664_p_spl_
  );


  and

  (
    g744_p,
    G21_p_spl_101,
    G11_p_spl_010
  );


  or

  (
    g744_n,
    G21_n_spl_101,
    G11_n_spl_010
  );


  and

  (
    g745_p,
    g661_n_spl_,
    g658_n_spl_
  );


  or

  (
    g745_n,
    g661_p_spl_,
    g658_p_spl_
  );


  and

  (
    g746_p,
    G20_p_spl_101,
    G12_p_spl_001
  );


  or

  (
    g746_n,
    G20_n_spl_101,
    G12_n_spl_001
  );


  and

  (
    g747_p,
    g655_n_spl_,
    g652_n_spl_
  );


  or

  (
    g747_n,
    g655_p_spl_,
    g652_p_spl_
  );


  and

  (
    g748_p,
    G19_p_spl_110,
    G13_p_spl_001
  );


  or

  (
    g748_n,
    G19_n_spl_110,
    G13_n_spl_001
  );


  and

  (
    g749_p,
    G17_p_spl_111,
    G15_p_spl_000
  );


  or

  (
    g749_n,
    G17_n_spl_110,
    G15_n_spl_000
  );


  and

  (
    g750_p,
    G18_p_spl_110,
    G14_p_spl_000
  );


  or

  (
    g750_n,
    G18_n_spl_110,
    G14_n_spl_000
  );


  and

  (
    g751_p,
    g750_n_spl_,
    g749_p_spl_
  );


  or

  (
    g751_n,
    g750_p_spl_,
    g749_n_spl_
  );


  and

  (
    g752_p,
    g751_n_spl_,
    g749_p_spl_
  );


  or

  (
    g752_n,
    g751_p_spl_,
    g749_n_spl_
  );


  and

  (
    g753_p,
    g751_n_spl_,
    g750_n_spl_
  );


  or

  (
    g753_n,
    g751_p_spl_,
    g750_p_spl_
  );


  and

  (
    g754_p,
    g753_n,
    g752_n_spl_0
  );


  or

  (
    g754_n,
    g753_p,
    g752_p_spl_0
  );


  and

  (
    g755_p,
    g754_n_spl_,
    g649_n_spl_0
  );


  or

  (
    g755_n,
    g754_p_spl_,
    g649_p_spl_0
  );


  and

  (
    g756_p,
    g754_p_spl_,
    g649_p_spl_
  );


  or

  (
    g756_n,
    g754_n_spl_,
    g649_n_spl_
  );


  and

  (
    g757_p,
    g756_n,
    g755_n_spl_
  );


  or

  (
    g757_n,
    g756_p,
    g755_p_spl_
  );


  and

  (
    g758_p,
    g757_p_spl_,
    g748_n_spl_
  );


  or

  (
    g758_n,
    g757_n_spl_,
    g748_p_spl_
  );


  and

  (
    g759_p,
    g757_n_spl_,
    g748_p_spl_
  );


  or

  (
    g759_n,
    g757_p_spl_,
    g748_n_spl_
  );


  and

  (
    g760_p,
    g759_n,
    g758_n_spl_
  );


  or

  (
    g760_n,
    g759_p,
    g758_p_spl_
  );


  and

  (
    g761_p,
    g760_p_spl_,
    g747_n_spl_
  );


  or

  (
    g761_n,
    g760_n_spl_,
    g747_p_spl_
  );


  and

  (
    g762_p,
    g760_n_spl_,
    g747_p_spl_
  );


  or

  (
    g762_n,
    g760_p_spl_,
    g747_n_spl_
  );


  and

  (
    g763_p,
    g762_n,
    g761_n_spl_
  );


  or

  (
    g763_n,
    g762_p,
    g761_p_spl_
  );


  and

  (
    g764_p,
    g763_p_spl_,
    g746_n_spl_
  );


  or

  (
    g764_n,
    g763_n_spl_,
    g746_p_spl_
  );


  and

  (
    g765_p,
    g763_n_spl_,
    g746_p_spl_
  );


  or

  (
    g765_n,
    g763_p_spl_,
    g746_n_spl_
  );


  and

  (
    g766_p,
    g765_n,
    g764_n_spl_
  );


  or

  (
    g766_n,
    g765_p,
    g764_p_spl_
  );


  and

  (
    g767_p,
    g766_p_spl_,
    g745_n_spl_
  );


  or

  (
    g767_n,
    g766_n_spl_,
    g745_p_spl_
  );


  and

  (
    g768_p,
    g766_n_spl_,
    g745_p_spl_
  );


  or

  (
    g768_n,
    g766_p_spl_,
    g745_n_spl_
  );


  and

  (
    g769_p,
    g768_n,
    g767_n_spl_
  );


  or

  (
    g769_n,
    g768_p,
    g767_p_spl_
  );


  and

  (
    g770_p,
    g769_p_spl_,
    g744_n_spl_
  );


  or

  (
    g770_n,
    g769_n_spl_,
    g744_p_spl_
  );


  and

  (
    g771_p,
    g769_n_spl_,
    g744_p_spl_
  );


  or

  (
    g771_n,
    g769_p_spl_,
    g744_n_spl_
  );


  and

  (
    g772_p,
    g771_n,
    g770_n_spl_
  );


  or

  (
    g772_n,
    g771_p,
    g770_p_spl_
  );


  and

  (
    g773_p,
    g772_p_spl_,
    g743_n_spl_
  );


  or

  (
    g773_n,
    g772_n_spl_,
    g743_p_spl_
  );


  and

  (
    g774_p,
    g772_n_spl_,
    g743_p_spl_
  );


  or

  (
    g774_n,
    g772_p_spl_,
    g743_n_spl_
  );


  and

  (
    g775_p,
    g774_n,
    g773_n_spl_
  );


  or

  (
    g775_n,
    g774_p,
    g773_p_spl_
  );


  and

  (
    g776_p,
    g775_p_spl_,
    g742_n_spl_
  );


  or

  (
    g776_n,
    g775_n_spl_,
    g742_p_spl_
  );


  and

  (
    g777_p,
    g775_n_spl_,
    g742_p_spl_
  );


  or

  (
    g777_n,
    g775_p_spl_,
    g742_n_spl_
  );


  and

  (
    g778_p,
    g777_n,
    g776_n_spl_
  );


  or

  (
    g778_n,
    g777_p,
    g776_p_spl_
  );


  and

  (
    g779_p,
    g778_p_spl_,
    g741_n_spl_
  );


  or

  (
    g779_n,
    g778_n_spl_,
    g741_p_spl_
  );


  and

  (
    g780_p,
    g778_n_spl_,
    g741_p_spl_
  );


  or

  (
    g780_n,
    g778_p_spl_,
    g741_n_spl_
  );


  and

  (
    g781_p,
    g780_n,
    g779_n_spl_
  );


  or

  (
    g781_n,
    g780_p,
    g779_p_spl_
  );


  and

  (
    g782_p,
    g781_p_spl_,
    g740_n_spl_
  );


  or

  (
    g782_n,
    g781_n_spl_,
    g740_p_spl_
  );


  and

  (
    g783_p,
    g781_n_spl_,
    g740_p_spl_
  );


  or

  (
    g783_n,
    g781_p_spl_,
    g740_n_spl_
  );


  and

  (
    g784_p,
    g783_n,
    g782_n_spl_
  );


  or

  (
    g784_n,
    g783_p,
    g782_p_spl_
  );


  and

  (
    g785_p,
    g784_p_spl_,
    g739_n_spl_
  );


  or

  (
    g785_n,
    g784_n_spl_,
    g739_p_spl_
  );


  and

  (
    g786_p,
    g784_n_spl_,
    g739_p_spl_
  );


  or

  (
    g786_n,
    g784_p_spl_,
    g739_n_spl_
  );


  and

  (
    g787_p,
    g786_n,
    g785_n_spl_
  );


  or

  (
    g787_n,
    g786_p,
    g785_p_spl_
  );


  and

  (
    g788_p,
    g787_p_spl_,
    g738_n_spl_
  );


  or

  (
    g788_n,
    g787_n_spl_,
    g738_p_spl_
  );


  and

  (
    g789_p,
    g787_n_spl_,
    g738_p_spl_
  );


  or

  (
    g789_n,
    g787_p_spl_,
    g738_n_spl_
  );


  and

  (
    g790_p,
    g789_n,
    g788_n_spl_
  );


  or

  (
    g790_n,
    g789_p,
    g788_p_spl_
  );


  and

  (
    g791_p,
    g790_p_spl_,
    g737_n_spl_
  );


  or

  (
    g791_n,
    g790_n_spl_,
    g737_p_spl_
  );


  and

  (
    g792_p,
    g790_n_spl_,
    g737_p_spl_
  );


  or

  (
    g792_n,
    g790_p_spl_,
    g737_n_spl_
  );


  and

  (
    g793_p,
    g792_n,
    g791_n_spl_
  );


  or

  (
    g793_n,
    g792_p,
    g791_p_spl_
  );


  and

  (
    g794_p,
    g793_p_spl_,
    g736_n_spl_
  );


  or

  (
    g794_n,
    g793_n_spl_,
    g736_p_spl_
  );


  and

  (
    g795_p,
    g793_n_spl_,
    g736_p_spl_
  );


  or

  (
    g795_n,
    g793_p_spl_,
    g736_n_spl_
  );


  and

  (
    g796_p,
    g795_n,
    g794_n_spl_
  );


  or

  (
    g796_n,
    g795_p,
    g794_p_spl_
  );


  and

  (
    g797_p,
    g796_p_spl_,
    g735_n_spl_
  );


  or

  (
    g797_n,
    g796_n_spl_,
    g735_p_spl_
  );


  and

  (
    g798_p,
    g796_n_spl_,
    g735_p_spl_
  );


  or

  (
    g798_n,
    g796_p_spl_,
    g735_n_spl_
  );


  and

  (
    g799_p,
    g798_n,
    g797_n_spl_
  );


  or

  (
    g799_n,
    g798_p,
    g797_p_spl_
  );


  and

  (
    g800_p,
    g799_p_spl_,
    g734_n_spl_
  );


  or

  (
    g800_n,
    g799_n_spl_,
    g734_p_spl_
  );


  and

  (
    g801_p,
    g799_n_spl_,
    g734_p_spl_
  );


  or

  (
    g801_n,
    g799_p_spl_,
    g734_n_spl_
  );


  and

  (
    g802_p,
    g801_n,
    g800_n_spl_
  );


  or

  (
    g802_n,
    g801_p,
    g800_p_spl_
  );


  and

  (
    g803_p,
    g802_p_spl_,
    g733_n_spl_
  );


  or

  (
    g803_n,
    g802_n_spl_,
    g733_p_spl_
  );


  and

  (
    g804_p,
    g802_n_spl_,
    g733_p_spl_
  );


  or

  (
    g804_n,
    g802_p_spl_,
    g733_n_spl_
  );


  and

  (
    g805_p,
    g804_n,
    g803_n_spl_
  );


  or

  (
    g805_n,
    g804_p,
    g803_p_spl_
  );


  and

  (
    g806_p,
    g805_p_spl_,
    g732_n_spl_
  );


  or

  (
    g806_n,
    g805_n_spl_,
    g732_p_spl_
  );


  and

  (
    g807_p,
    g805_n_spl_,
    g732_p_spl_
  );


  or

  (
    g807_n,
    g805_p_spl_,
    g732_n_spl_
  );


  and

  (
    g808_p,
    g807_n,
    g806_n_spl_
  );


  or

  (
    g808_n,
    g807_p,
    g806_p_spl_
  );


  and

  (
    g809_p,
    g808_p_spl_,
    g731_n_spl_
  );


  or

  (
    g809_n,
    g808_n_spl_,
    g731_p_spl_
  );


  and

  (
    g810_p,
    g808_n_spl_,
    g731_p_spl_
  );


  or

  (
    g810_n,
    g808_p_spl_,
    g731_n_spl_
  );


  and

  (
    g811_p,
    g810_n,
    g809_n_spl_
  );


  or

  (
    g811_n,
    g810_p,
    g809_p_spl_
  );


  and

  (
    g812_p,
    g811_p_spl_,
    g730_n_spl_
  );


  or

  (
    g812_n,
    g811_n_spl_,
    g730_p_spl_
  );


  and

  (
    g813_p,
    g811_n_spl_,
    g730_p_spl_
  );


  or

  (
    g813_n,
    g811_p_spl_,
    g730_n_spl_
  );


  and

  (
    g814_p,
    g813_n,
    g812_n_spl_
  );


  or

  (
    g814_n,
    g813_p,
    g812_p_spl_
  );


  and

  (
    g815_p,
    g814_p_spl_,
    g729_n_spl_
  );


  or

  (
    g815_n,
    g814_n_spl_,
    g729_p_spl_
  );


  and

  (
    g816_p,
    g814_n_spl_,
    g729_p_spl_
  );


  or

  (
    g816_n,
    g814_p_spl_,
    g729_n_spl_
  );


  and

  (
    g817_p,
    g816_n,
    g815_n_spl_
  );


  or

  (
    g817_n,
    g816_p,
    g815_p_spl_
  );


  and

  (
    g818_p,
    g817_p_spl_,
    g728_n_spl_
  );


  or

  (
    g818_n,
    g817_n_spl_,
    g728_p_spl_
  );


  and

  (
    g819_p,
    g817_n_spl_,
    g728_p_spl_
  );


  or

  (
    g819_n,
    g817_p_spl_,
    g728_n_spl_
  );


  and

  (
    g820_p,
    g819_n,
    g818_n_spl_
  );


  or

  (
    g820_n,
    g819_p,
    g818_p_spl_
  );


  and

  (
    g821_p,
    g820_p_spl_,
    g727_n_spl_
  );


  or

  (
    g821_n,
    g820_n_spl_,
    g727_p_spl_
  );


  and

  (
    g822_p,
    g820_n_spl_,
    g727_p_spl_
  );


  or

  (
    g822_n,
    g820_p_spl_,
    g727_n_spl_
  );


  and

  (
    g823_p,
    g822_n,
    g821_n_spl_
  );


  or

  (
    g823_n,
    g822_p,
    g821_p_spl_
  );


  and

  (
    g824_p,
    g823_p_spl_,
    g726_n_spl_
  );


  or

  (
    g824_n,
    g823_n_spl_,
    g726_p_spl_
  );


  and

  (
    g825_p,
    g823_n_spl_,
    g726_p_spl_
  );


  or

  (
    g825_n,
    g823_p_spl_,
    g726_n_spl_
  );


  and

  (
    g826_p,
    g825_n,
    g824_n_spl_
  );


  or

  (
    g826_n,
    g825_p,
    g824_p_spl_
  );


  and

  (
    g827_p,
    g826_p_spl_,
    g725_n_spl_
  );


  or

  (
    g827_n,
    g826_n_spl_,
    g725_p_spl_
  );


  and

  (
    g828_p,
    g826_n_spl_,
    g725_p_spl_
  );


  or

  (
    g828_n,
    g826_p_spl_,
    g725_n_spl_
  );


  and

  (
    g829_p,
    g828_n,
    g827_n_spl_
  );


  or

  (
    g829_n,
    g828_p,
    g827_p_spl_
  );


  and

  (
    g830_p,
    g829_p,
    g724_n
  );


  or

  (
    g830_n,
    g829_n_spl_,
    g724_p_spl_
  );


  and

  (
    g831_p,
    g829_n_spl_,
    g724_p_spl_
  );


  or

  (
    g832_n,
    g831_p,
    g830_p_spl_
  );


  and

  (
    g833_p,
    G32_p_spl_000,
    G1_p_spl_111
  );


  or

  (
    g833_n,
    G32_n_spl_000,
    G1_n_spl_11
  );


  and

  (
    g834_p,
    g830_n,
    g827_n_spl_
  );


  or

  (
    g834_n,
    g830_p_spl_,
    g827_p_spl_
  );


  and

  (
    g835_p,
    G31_p_spl_000,
    G2_p_spl_111
  );


  or

  (
    g835_n,
    G31_n_spl_000,
    G2_n_spl_111
  );


  and

  (
    g836_p,
    g824_n_spl_,
    g821_n_spl_
  );


  or

  (
    g836_n,
    g824_p_spl_,
    g821_p_spl_
  );


  and

  (
    g837_p,
    G30_p_spl_001,
    G3_p_spl_110
  );


  or

  (
    g837_n,
    G30_n_spl_001,
    G3_n_spl_110
  );


  and

  (
    g838_p,
    g818_n_spl_,
    g815_n_spl_
  );


  or

  (
    g838_n,
    g818_p_spl_,
    g815_p_spl_
  );


  and

  (
    g839_p,
    G29_p_spl_001,
    G4_p_spl_110
  );


  or

  (
    g839_n,
    G29_n_spl_001,
    G4_n_spl_110
  );


  and

  (
    g840_p,
    g812_n_spl_,
    g809_n_spl_
  );


  or

  (
    g840_n,
    g812_p_spl_,
    g809_p_spl_
  );


  and

  (
    g841_p,
    G28_p_spl_010,
    G5_p_spl_101
  );


  or

  (
    g841_n,
    G28_n_spl_010,
    G5_n_spl_101
  );


  and

  (
    g842_p,
    g806_n_spl_,
    g803_n_spl_
  );


  or

  (
    g842_n,
    g806_p_spl_,
    g803_p_spl_
  );


  and

  (
    g843_p,
    G27_p_spl_010,
    G6_p_spl_101
  );


  or

  (
    g843_n,
    G27_n_spl_010,
    G6_n_spl_101
  );


  and

  (
    g844_p,
    g800_n_spl_,
    g797_n_spl_
  );


  or

  (
    g844_n,
    g800_p_spl_,
    g797_p_spl_
  );


  and

  (
    g845_p,
    G26_p_spl_011,
    G7_p_spl_100
  );


  or

  (
    g845_n,
    G26_n_spl_011,
    G7_n_spl_100
  );


  and

  (
    g846_p,
    g794_n_spl_,
    g791_n_spl_
  );


  or

  (
    g846_n,
    g794_p_spl_,
    g791_p_spl_
  );


  and

  (
    g847_p,
    G25_p_spl_011,
    G8_p_spl_100
  );


  or

  (
    g847_n,
    G25_n_spl_011,
    G8_n_spl_100
  );


  and

  (
    g848_p,
    g788_n_spl_,
    g785_n_spl_
  );


  or

  (
    g848_n,
    g788_p_spl_,
    g785_p_spl_
  );


  and

  (
    g849_p,
    G24_p_spl_100,
    G9_p_spl_011
  );


  or

  (
    g849_n,
    G24_n_spl_100,
    G9_n_spl_011
  );


  and

  (
    g850_p,
    g782_n_spl_,
    g779_n_spl_
  );


  or

  (
    g850_n,
    g782_p_spl_,
    g779_p_spl_
  );


  and

  (
    g851_p,
    G23_p_spl_100,
    G10_p_spl_011
  );


  or

  (
    g851_n,
    G23_n_spl_100,
    G10_n_spl_011
  );


  and

  (
    g852_p,
    g776_n_spl_,
    g773_n_spl_
  );


  or

  (
    g852_n,
    g776_p_spl_,
    g773_p_spl_
  );


  and

  (
    g853_p,
    G22_p_spl_101,
    G11_p_spl_010
  );


  or

  (
    g853_n,
    G22_n_spl_101,
    G11_n_spl_010
  );


  and

  (
    g854_p,
    g770_n_spl_,
    g767_n_spl_
  );


  or

  (
    g854_n,
    g770_p_spl_,
    g767_p_spl_
  );


  and

  (
    g855_p,
    G21_p_spl_101,
    G12_p_spl_010
  );


  or

  (
    g855_n,
    G21_n_spl_101,
    G12_n_spl_010
  );


  and

  (
    g856_p,
    g764_n_spl_,
    g761_n_spl_
  );


  or

  (
    g856_n,
    g764_p_spl_,
    g761_p_spl_
  );


  and

  (
    g857_p,
    G20_p_spl_110,
    G13_p_spl_001
  );


  or

  (
    g857_n,
    G20_n_spl_110,
    G13_n_spl_001
  );


  and

  (
    g858_p,
    g758_n_spl_,
    g755_n_spl_
  );


  or

  (
    g858_n,
    g758_p_spl_,
    g755_p_spl_
  );


  and

  (
    g859_p,
    G19_p_spl_110,
    G14_p_spl_001
  );


  or

  (
    g859_n,
    G19_n_spl_110,
    G14_n_spl_001
  );


  and

  (
    g860_p,
    G17_p_spl_111,
    G16_p_spl_000
  );


  or

  (
    g860_n,
    G17_n_spl_11,
    G16_n_spl_000
  );


  and

  (
    g861_p,
    G18_p_spl_111,
    G15_p_spl_000
  );


  or

  (
    g861_n,
    G18_n_spl_111,
    G15_n_spl_000
  );


  and

  (
    g862_p,
    g861_n_spl_,
    g860_p_spl_
  );


  or

  (
    g862_n,
    g861_p_spl_,
    g860_n_spl_
  );


  and

  (
    g863_p,
    g862_n_spl_,
    g860_p_spl_
  );


  or

  (
    g863_n,
    g862_p_spl_,
    g860_n_spl_
  );


  and

  (
    g864_p,
    g862_n_spl_,
    g861_n_spl_
  );


  or

  (
    g864_n,
    g862_p_spl_,
    g861_p_spl_
  );


  and

  (
    g865_p,
    g864_n,
    g863_n_spl_
  );


  or

  (
    g865_n,
    g864_p,
    g863_p_spl_
  );


  and

  (
    g866_p,
    g865_n_spl_,
    g752_n_spl_0
  );


  or

  (
    g866_n,
    g865_p_spl_,
    g752_p_spl_0
  );


  and

  (
    g867_p,
    g865_p_spl_,
    g752_p_spl_
  );


  or

  (
    g867_n,
    g865_n_spl_,
    g752_n_spl_
  );


  and

  (
    g868_p,
    g867_n,
    g866_n_spl_
  );


  or

  (
    g868_n,
    g867_p,
    g866_p_spl_
  );


  and

  (
    g869_p,
    g868_p_spl_,
    g859_n_spl_
  );


  or

  (
    g869_n,
    g868_n_spl_,
    g859_p_spl_
  );


  and

  (
    g870_p,
    g868_n_spl_,
    g859_p_spl_
  );


  or

  (
    g870_n,
    g868_p_spl_,
    g859_n_spl_
  );


  and

  (
    g871_p,
    g870_n,
    g869_n_spl_
  );


  or

  (
    g871_n,
    g870_p,
    g869_p_spl_
  );


  and

  (
    g872_p,
    g871_p_spl_,
    g858_n_spl_
  );


  or

  (
    g872_n,
    g871_n_spl_,
    g858_p_spl_
  );


  and

  (
    g873_p,
    g871_n_spl_,
    g858_p_spl_
  );


  or

  (
    g873_n,
    g871_p_spl_,
    g858_n_spl_
  );


  and

  (
    g874_p,
    g873_n,
    g872_n_spl_
  );


  or

  (
    g874_n,
    g873_p,
    g872_p_spl_
  );


  and

  (
    g875_p,
    g874_p_spl_,
    g857_n_spl_
  );


  or

  (
    g875_n,
    g874_n_spl_,
    g857_p_spl_
  );


  and

  (
    g876_p,
    g874_n_spl_,
    g857_p_spl_
  );


  or

  (
    g876_n,
    g874_p_spl_,
    g857_n_spl_
  );


  and

  (
    g877_p,
    g876_n,
    g875_n_spl_
  );


  or

  (
    g877_n,
    g876_p,
    g875_p_spl_
  );


  and

  (
    g878_p,
    g877_p_spl_,
    g856_n_spl_
  );


  or

  (
    g878_n,
    g877_n_spl_,
    g856_p_spl_
  );


  and

  (
    g879_p,
    g877_n_spl_,
    g856_p_spl_
  );


  or

  (
    g879_n,
    g877_p_spl_,
    g856_n_spl_
  );


  and

  (
    g880_p,
    g879_n,
    g878_n_spl_
  );


  or

  (
    g880_n,
    g879_p,
    g878_p_spl_
  );


  and

  (
    g881_p,
    g880_p_spl_,
    g855_n_spl_
  );


  or

  (
    g881_n,
    g880_n_spl_,
    g855_p_spl_
  );


  and

  (
    g882_p,
    g880_n_spl_,
    g855_p_spl_
  );


  or

  (
    g882_n,
    g880_p_spl_,
    g855_n_spl_
  );


  and

  (
    g883_p,
    g882_n,
    g881_n_spl_
  );


  or

  (
    g883_n,
    g882_p,
    g881_p_spl_
  );


  and

  (
    g884_p,
    g883_p_spl_,
    g854_n_spl_
  );


  or

  (
    g884_n,
    g883_n_spl_,
    g854_p_spl_
  );


  and

  (
    g885_p,
    g883_n_spl_,
    g854_p_spl_
  );


  or

  (
    g885_n,
    g883_p_spl_,
    g854_n_spl_
  );


  and

  (
    g886_p,
    g885_n,
    g884_n_spl_
  );


  or

  (
    g886_n,
    g885_p,
    g884_p_spl_
  );


  and

  (
    g887_p,
    g886_p_spl_,
    g853_n_spl_
  );


  or

  (
    g887_n,
    g886_n_spl_,
    g853_p_spl_
  );


  and

  (
    g888_p,
    g886_n_spl_,
    g853_p_spl_
  );


  or

  (
    g888_n,
    g886_p_spl_,
    g853_n_spl_
  );


  and

  (
    g889_p,
    g888_n,
    g887_n_spl_
  );


  or

  (
    g889_n,
    g888_p,
    g887_p_spl_
  );


  and

  (
    g890_p,
    g889_p_spl_,
    g852_n_spl_
  );


  or

  (
    g890_n,
    g889_n_spl_,
    g852_p_spl_
  );


  and

  (
    g891_p,
    g889_n_spl_,
    g852_p_spl_
  );


  or

  (
    g891_n,
    g889_p_spl_,
    g852_n_spl_
  );


  and

  (
    g892_p,
    g891_n,
    g890_n_spl_
  );


  or

  (
    g892_n,
    g891_p,
    g890_p_spl_
  );


  and

  (
    g893_p,
    g892_p_spl_,
    g851_n_spl_
  );


  or

  (
    g893_n,
    g892_n_spl_,
    g851_p_spl_
  );


  and

  (
    g894_p,
    g892_n_spl_,
    g851_p_spl_
  );


  or

  (
    g894_n,
    g892_p_spl_,
    g851_n_spl_
  );


  and

  (
    g895_p,
    g894_n,
    g893_n_spl_
  );


  or

  (
    g895_n,
    g894_p,
    g893_p_spl_
  );


  and

  (
    g896_p,
    g895_p_spl_,
    g850_n_spl_
  );


  or

  (
    g896_n,
    g895_n_spl_,
    g850_p_spl_
  );


  and

  (
    g897_p,
    g895_n_spl_,
    g850_p_spl_
  );


  or

  (
    g897_n,
    g895_p_spl_,
    g850_n_spl_
  );


  and

  (
    g898_p,
    g897_n,
    g896_n_spl_
  );


  or

  (
    g898_n,
    g897_p,
    g896_p_spl_
  );


  and

  (
    g899_p,
    g898_p_spl_,
    g849_n_spl_
  );


  or

  (
    g899_n,
    g898_n_spl_,
    g849_p_spl_
  );


  and

  (
    g900_p,
    g898_n_spl_,
    g849_p_spl_
  );


  or

  (
    g900_n,
    g898_p_spl_,
    g849_n_spl_
  );


  and

  (
    g901_p,
    g900_n,
    g899_n_spl_
  );


  or

  (
    g901_n,
    g900_p,
    g899_p_spl_
  );


  and

  (
    g902_p,
    g901_p_spl_,
    g848_n_spl_
  );


  or

  (
    g902_n,
    g901_n_spl_,
    g848_p_spl_
  );


  and

  (
    g903_p,
    g901_n_spl_,
    g848_p_spl_
  );


  or

  (
    g903_n,
    g901_p_spl_,
    g848_n_spl_
  );


  and

  (
    g904_p,
    g903_n,
    g902_n_spl_
  );


  or

  (
    g904_n,
    g903_p,
    g902_p_spl_
  );


  and

  (
    g905_p,
    g904_p_spl_,
    g847_n_spl_
  );


  or

  (
    g905_n,
    g904_n_spl_,
    g847_p_spl_
  );


  and

  (
    g906_p,
    g904_n_spl_,
    g847_p_spl_
  );


  or

  (
    g906_n,
    g904_p_spl_,
    g847_n_spl_
  );


  and

  (
    g907_p,
    g906_n,
    g905_n_spl_
  );


  or

  (
    g907_n,
    g906_p,
    g905_p_spl_
  );


  and

  (
    g908_p,
    g907_p_spl_,
    g846_n_spl_
  );


  or

  (
    g908_n,
    g907_n_spl_,
    g846_p_spl_
  );


  and

  (
    g909_p,
    g907_n_spl_,
    g846_p_spl_
  );


  or

  (
    g909_n,
    g907_p_spl_,
    g846_n_spl_
  );


  and

  (
    g910_p,
    g909_n,
    g908_n_spl_
  );


  or

  (
    g910_n,
    g909_p,
    g908_p_spl_
  );


  and

  (
    g911_p,
    g910_p_spl_,
    g845_n_spl_
  );


  or

  (
    g911_n,
    g910_n_spl_,
    g845_p_spl_
  );


  and

  (
    g912_p,
    g910_n_spl_,
    g845_p_spl_
  );


  or

  (
    g912_n,
    g910_p_spl_,
    g845_n_spl_
  );


  and

  (
    g913_p,
    g912_n,
    g911_n_spl_
  );


  or

  (
    g913_n,
    g912_p,
    g911_p_spl_
  );


  and

  (
    g914_p,
    g913_p_spl_,
    g844_n_spl_
  );


  or

  (
    g914_n,
    g913_n_spl_,
    g844_p_spl_
  );


  and

  (
    g915_p,
    g913_n_spl_,
    g844_p_spl_
  );


  or

  (
    g915_n,
    g913_p_spl_,
    g844_n_spl_
  );


  and

  (
    g916_p,
    g915_n,
    g914_n_spl_
  );


  or

  (
    g916_n,
    g915_p,
    g914_p_spl_
  );


  and

  (
    g917_p,
    g916_p_spl_,
    g843_n_spl_
  );


  or

  (
    g917_n,
    g916_n_spl_,
    g843_p_spl_
  );


  and

  (
    g918_p,
    g916_n_spl_,
    g843_p_spl_
  );


  or

  (
    g918_n,
    g916_p_spl_,
    g843_n_spl_
  );


  and

  (
    g919_p,
    g918_n,
    g917_n_spl_
  );


  or

  (
    g919_n,
    g918_p,
    g917_p_spl_
  );


  and

  (
    g920_p,
    g919_p_spl_,
    g842_n_spl_
  );


  or

  (
    g920_n,
    g919_n_spl_,
    g842_p_spl_
  );


  and

  (
    g921_p,
    g919_n_spl_,
    g842_p_spl_
  );


  or

  (
    g921_n,
    g919_p_spl_,
    g842_n_spl_
  );


  and

  (
    g922_p,
    g921_n,
    g920_n_spl_
  );


  or

  (
    g922_n,
    g921_p,
    g920_p_spl_
  );


  and

  (
    g923_p,
    g922_p_spl_,
    g841_n_spl_
  );


  or

  (
    g923_n,
    g922_n_spl_,
    g841_p_spl_
  );


  and

  (
    g924_p,
    g922_n_spl_,
    g841_p_spl_
  );


  or

  (
    g924_n,
    g922_p_spl_,
    g841_n_spl_
  );


  and

  (
    g925_p,
    g924_n,
    g923_n_spl_
  );


  or

  (
    g925_n,
    g924_p,
    g923_p_spl_
  );


  and

  (
    g926_p,
    g925_p_spl_,
    g840_n_spl_
  );


  or

  (
    g926_n,
    g925_n_spl_,
    g840_p_spl_
  );


  and

  (
    g927_p,
    g925_n_spl_,
    g840_p_spl_
  );


  or

  (
    g927_n,
    g925_p_spl_,
    g840_n_spl_
  );


  and

  (
    g928_p,
    g927_n,
    g926_n_spl_
  );


  or

  (
    g928_n,
    g927_p,
    g926_p_spl_
  );


  and

  (
    g929_p,
    g928_p_spl_,
    g839_n_spl_
  );


  or

  (
    g929_n,
    g928_n_spl_,
    g839_p_spl_
  );


  and

  (
    g930_p,
    g928_n_spl_,
    g839_p_spl_
  );


  or

  (
    g930_n,
    g928_p_spl_,
    g839_n_spl_
  );


  and

  (
    g931_p,
    g930_n,
    g929_n_spl_
  );


  or

  (
    g931_n,
    g930_p,
    g929_p_spl_
  );


  and

  (
    g932_p,
    g931_p_spl_,
    g838_n_spl_
  );


  or

  (
    g932_n,
    g931_n_spl_,
    g838_p_spl_
  );


  and

  (
    g933_p,
    g931_n_spl_,
    g838_p_spl_
  );


  or

  (
    g933_n,
    g931_p_spl_,
    g838_n_spl_
  );


  and

  (
    g934_p,
    g933_n,
    g932_n_spl_
  );


  or

  (
    g934_n,
    g933_p,
    g932_p_spl_
  );


  and

  (
    g935_p,
    g934_p_spl_,
    g837_n_spl_
  );


  or

  (
    g935_n,
    g934_n_spl_,
    g837_p_spl_
  );


  and

  (
    g936_p,
    g934_n_spl_,
    g837_p_spl_
  );


  or

  (
    g936_n,
    g934_p_spl_,
    g837_n_spl_
  );


  and

  (
    g937_p,
    g936_n,
    g935_n_spl_
  );


  or

  (
    g937_n,
    g936_p,
    g935_p_spl_
  );


  and

  (
    g938_p,
    g937_p_spl_,
    g836_n_spl_
  );


  or

  (
    g938_n,
    g937_n_spl_,
    g836_p_spl_
  );


  and

  (
    g939_p,
    g937_n_spl_,
    g836_p_spl_
  );


  or

  (
    g939_n,
    g937_p_spl_,
    g836_n_spl_
  );


  and

  (
    g940_p,
    g939_n,
    g938_n_spl_
  );


  or

  (
    g940_n,
    g939_p,
    g938_p_spl_
  );


  and

  (
    g941_p,
    g940_p_spl_,
    g835_n_spl_
  );


  or

  (
    g941_n,
    g940_n_spl_,
    g835_p_spl_
  );


  and

  (
    g942_p,
    g940_n_spl_,
    g835_p_spl_
  );


  or

  (
    g942_n,
    g940_p_spl_,
    g835_n_spl_
  );


  and

  (
    g943_p,
    g942_n,
    g941_n_spl_
  );


  or

  (
    g943_n,
    g942_p,
    g941_p_spl_
  );


  and

  (
    g944_p,
    g943_p_spl_,
    g834_n_spl_
  );


  or

  (
    g944_n,
    g943_n_spl_,
    g834_p_spl_
  );


  and

  (
    g945_p,
    g943_n_spl_,
    g834_p_spl_
  );


  or

  (
    g945_n,
    g943_p_spl_,
    g834_n_spl_
  );


  and

  (
    g946_p,
    g945_n,
    g944_n_spl_
  );


  or

  (
    g946_n,
    g945_p,
    g944_p_spl_
  );


  and

  (
    g947_p,
    g946_p,
    g833_n
  );


  or

  (
    g947_n,
    g946_n_spl_,
    g833_p_spl_
  );


  and

  (
    g948_p,
    g946_n_spl_,
    g833_p_spl_
  );


  or

  (
    g949_n,
    g948_p,
    g947_p_spl_
  );


  and

  (
    g950_p,
    g947_n,
    g944_n_spl_
  );


  or

  (
    g950_n,
    g947_p_spl_,
    g944_p_spl_
  );


  and

  (
    g951_p,
    G32_p_spl_000,
    G2_p_spl_111
  );


  or

  (
    g951_n,
    G32_n_spl_000,
    G2_n_spl_111
  );


  and

  (
    g952_p,
    g941_n_spl_,
    g938_n_spl_
  );


  or

  (
    g952_n,
    g941_p_spl_,
    g938_p_spl_
  );


  and

  (
    g953_p,
    G31_p_spl_001,
    G3_p_spl_111
  );


  or

  (
    g953_n,
    G31_n_spl_001,
    G3_n_spl_111
  );


  and

  (
    g954_p,
    g935_n_spl_,
    g932_n_spl_
  );


  or

  (
    g954_n,
    g935_p_spl_,
    g932_p_spl_
  );


  and

  (
    g955_p,
    G30_p_spl_001,
    G4_p_spl_110
  );


  or

  (
    g955_n,
    G30_n_spl_001,
    G4_n_spl_110
  );


  and

  (
    g956_p,
    g929_n_spl_,
    g926_n_spl_
  );


  or

  (
    g956_n,
    g929_p_spl_,
    g926_p_spl_
  );


  and

  (
    g957_p,
    G29_p_spl_010,
    G5_p_spl_110
  );


  or

  (
    g957_n,
    G29_n_spl_010,
    G5_n_spl_110
  );


  and

  (
    g958_p,
    g923_n_spl_,
    g920_n_spl_
  );


  or

  (
    g958_n,
    g923_p_spl_,
    g920_p_spl_
  );


  and

  (
    g959_p,
    G28_p_spl_010,
    G6_p_spl_101
  );


  or

  (
    g959_n,
    G28_n_spl_010,
    G6_n_spl_101
  );


  and

  (
    g960_p,
    g917_n_spl_,
    g914_n_spl_
  );


  or

  (
    g960_n,
    g917_p_spl_,
    g914_p_spl_
  );


  and

  (
    g961_p,
    G27_p_spl_011,
    G7_p_spl_101
  );


  or

  (
    g961_n,
    G27_n_spl_011,
    G7_n_spl_101
  );


  and

  (
    g962_p,
    g911_n_spl_,
    g908_n_spl_
  );


  or

  (
    g962_n,
    g911_p_spl_,
    g908_p_spl_
  );


  and

  (
    g963_p,
    G26_p_spl_011,
    G8_p_spl_100
  );


  or

  (
    g963_n,
    G26_n_spl_011,
    G8_n_spl_100
  );


  and

  (
    g964_p,
    g905_n_spl_,
    g902_n_spl_
  );


  or

  (
    g964_n,
    g905_p_spl_,
    g902_p_spl_
  );


  and

  (
    g965_p,
    G25_p_spl_100,
    G9_p_spl_100
  );


  or

  (
    g965_n,
    G25_n_spl_100,
    G9_n_spl_100
  );


  and

  (
    g966_p,
    g899_n_spl_,
    g896_n_spl_
  );


  or

  (
    g966_n,
    g899_p_spl_,
    g896_p_spl_
  );


  and

  (
    g967_p,
    G24_p_spl_100,
    G10_p_spl_011
  );


  or

  (
    g967_n,
    G24_n_spl_100,
    G10_n_spl_011
  );


  and

  (
    g968_p,
    g893_n_spl_,
    g890_n_spl_
  );


  or

  (
    g968_n,
    g893_p_spl_,
    g890_p_spl_
  );


  and

  (
    g969_p,
    G23_p_spl_101,
    G11_p_spl_011
  );


  or

  (
    g969_n,
    G23_n_spl_101,
    G11_n_spl_011
  );


  and

  (
    g970_p,
    g887_n_spl_,
    g884_n_spl_
  );


  or

  (
    g970_n,
    g887_p_spl_,
    g884_p_spl_
  );


  and

  (
    g971_p,
    G22_p_spl_101,
    G12_p_spl_010
  );


  or

  (
    g971_n,
    G22_n_spl_101,
    G12_n_spl_010
  );


  and

  (
    g972_p,
    g881_n_spl_,
    g878_n_spl_
  );


  or

  (
    g972_n,
    g881_p_spl_,
    g878_p_spl_
  );


  and

  (
    g973_p,
    G21_p_spl_110,
    G13_p_spl_010
  );


  or

  (
    g973_n,
    G21_n_spl_110,
    G13_n_spl_010
  );


  and

  (
    g974_p,
    g875_n_spl_,
    g872_n_spl_
  );


  or

  (
    g974_n,
    g875_p_spl_,
    g872_p_spl_
  );


  and

  (
    g975_p,
    G20_p_spl_110,
    G14_p_spl_001
  );


  or

  (
    g975_n,
    G20_n_spl_110,
    G14_n_spl_001
  );


  and

  (
    g976_p,
    g869_n_spl_,
    g866_n_spl_
  );


  or

  (
    g976_n,
    g869_p_spl_,
    g866_p_spl_
  );


  and

  (
    g977_p,
    G18_p_spl_111,
    G16_p_spl_000
  );


  or

  (
    g977_n,
    G18_n_spl_111,
    G16_n_spl_000
  );


  and

  (
    g978_p,
    g977_p_spl_,
    g863_n_spl_
  );


  or

  (
    g978_n,
    g977_n_spl_,
    g863_p_spl_
  );


  and

  (
    g979_p,
    G19_p_spl_111,
    G15_p_spl_001
  );


  or

  (
    g979_n,
    G19_n_spl_111,
    G15_n_spl_001
  );


  and

  (
    g980_p,
    g979_n_spl_,
    g978_p_spl_
  );


  or

  (
    g980_n,
    g979_p_spl_,
    g978_n_spl_
  );


  and

  (
    g981_p,
    g979_p_spl_,
    g978_n_spl_
  );


  or

  (
    g981_n,
    g979_n_spl_,
    g978_p_spl_
  );


  and

  (
    g982_p,
    g981_n,
    g980_n_spl_
  );


  or

  (
    g982_n,
    g981_p,
    g980_p_spl_
  );


  and

  (
    g983_p,
    g982_p_spl_,
    g976_n_spl_
  );


  or

  (
    g983_n,
    g982_n_spl_,
    g976_p_spl_
  );


  and

  (
    g984_p,
    g982_n_spl_,
    g976_p_spl_
  );


  or

  (
    g984_n,
    g982_p_spl_,
    g976_n_spl_
  );


  and

  (
    g985_p,
    g984_n,
    g983_n_spl_
  );


  or

  (
    g985_n,
    g984_p,
    g983_p_spl_
  );


  and

  (
    g986_p,
    g985_p_spl_,
    g975_n_spl_
  );


  or

  (
    g986_n,
    g985_n_spl_,
    g975_p_spl_
  );


  and

  (
    g987_p,
    g985_n_spl_,
    g975_p_spl_
  );


  or

  (
    g987_n,
    g985_p_spl_,
    g975_n_spl_
  );


  and

  (
    g988_p,
    g987_n,
    g986_n_spl_
  );


  or

  (
    g988_n,
    g987_p,
    g986_p_spl_
  );


  and

  (
    g989_p,
    g988_p_spl_,
    g974_n_spl_
  );


  or

  (
    g989_n,
    g988_n_spl_,
    g974_p_spl_
  );


  and

  (
    g990_p,
    g988_n_spl_,
    g974_p_spl_
  );


  or

  (
    g990_n,
    g988_p_spl_,
    g974_n_spl_
  );


  and

  (
    g991_p,
    g990_n,
    g989_n_spl_
  );


  or

  (
    g991_n,
    g990_p,
    g989_p_spl_
  );


  and

  (
    g992_p,
    g991_p_spl_,
    g973_n_spl_
  );


  or

  (
    g992_n,
    g991_n_spl_,
    g973_p_spl_
  );


  and

  (
    g993_p,
    g991_n_spl_,
    g973_p_spl_
  );


  or

  (
    g993_n,
    g991_p_spl_,
    g973_n_spl_
  );


  and

  (
    g994_p,
    g993_n,
    g992_n_spl_
  );


  or

  (
    g994_n,
    g993_p,
    g992_p_spl_
  );


  and

  (
    g995_p,
    g994_p_spl_,
    g972_n_spl_
  );


  or

  (
    g995_n,
    g994_n_spl_,
    g972_p_spl_
  );


  and

  (
    g996_p,
    g994_n_spl_,
    g972_p_spl_
  );


  or

  (
    g996_n,
    g994_p_spl_,
    g972_n_spl_
  );


  and

  (
    g997_p,
    g996_n,
    g995_n_spl_
  );


  or

  (
    g997_n,
    g996_p,
    g995_p_spl_
  );


  and

  (
    g998_p,
    g997_p_spl_,
    g971_n_spl_
  );


  or

  (
    g998_n,
    g997_n_spl_,
    g971_p_spl_
  );


  and

  (
    g999_p,
    g997_n_spl_,
    g971_p_spl_
  );


  or

  (
    g999_n,
    g997_p_spl_,
    g971_n_spl_
  );


  and

  (
    g1000_p,
    g999_n,
    g998_n_spl_
  );


  or

  (
    g1000_n,
    g999_p,
    g998_p_spl_
  );


  and

  (
    g1001_p,
    g1000_p_spl_,
    g970_n_spl_
  );


  or

  (
    g1001_n,
    g1000_n_spl_,
    g970_p_spl_
  );


  and

  (
    g1002_p,
    g1000_n_spl_,
    g970_p_spl_
  );


  or

  (
    g1002_n,
    g1000_p_spl_,
    g970_n_spl_
  );


  and

  (
    g1003_p,
    g1002_n,
    g1001_n_spl_
  );


  or

  (
    g1003_n,
    g1002_p,
    g1001_p_spl_
  );


  and

  (
    g1004_p,
    g1003_p_spl_,
    g969_n_spl_
  );


  or

  (
    g1004_n,
    g1003_n_spl_,
    g969_p_spl_
  );


  and

  (
    g1005_p,
    g1003_n_spl_,
    g969_p_spl_
  );


  or

  (
    g1005_n,
    g1003_p_spl_,
    g969_n_spl_
  );


  and

  (
    g1006_p,
    g1005_n,
    g1004_n_spl_
  );


  or

  (
    g1006_n,
    g1005_p,
    g1004_p_spl_
  );


  and

  (
    g1007_p,
    g1006_p_spl_,
    g968_n_spl_
  );


  or

  (
    g1007_n,
    g1006_n_spl_,
    g968_p_spl_
  );


  and

  (
    g1008_p,
    g1006_n_spl_,
    g968_p_spl_
  );


  or

  (
    g1008_n,
    g1006_p_spl_,
    g968_n_spl_
  );


  and

  (
    g1009_p,
    g1008_n,
    g1007_n_spl_
  );


  or

  (
    g1009_n,
    g1008_p,
    g1007_p_spl_
  );


  and

  (
    g1010_p,
    g1009_p_spl_,
    g967_n_spl_
  );


  or

  (
    g1010_n,
    g1009_n_spl_,
    g967_p_spl_
  );


  and

  (
    g1011_p,
    g1009_n_spl_,
    g967_p_spl_
  );


  or

  (
    g1011_n,
    g1009_p_spl_,
    g967_n_spl_
  );


  and

  (
    g1012_p,
    g1011_n,
    g1010_n_spl_
  );


  or

  (
    g1012_n,
    g1011_p,
    g1010_p_spl_
  );


  and

  (
    g1013_p,
    g1012_p_spl_,
    g966_n_spl_
  );


  or

  (
    g1013_n,
    g1012_n_spl_,
    g966_p_spl_
  );


  and

  (
    g1014_p,
    g1012_n_spl_,
    g966_p_spl_
  );


  or

  (
    g1014_n,
    g1012_p_spl_,
    g966_n_spl_
  );


  and

  (
    g1015_p,
    g1014_n,
    g1013_n_spl_
  );


  or

  (
    g1015_n,
    g1014_p,
    g1013_p_spl_
  );


  and

  (
    g1016_p,
    g1015_p_spl_,
    g965_n_spl_
  );


  or

  (
    g1016_n,
    g1015_n_spl_,
    g965_p_spl_
  );


  and

  (
    g1017_p,
    g1015_n_spl_,
    g965_p_spl_
  );


  or

  (
    g1017_n,
    g1015_p_spl_,
    g965_n_spl_
  );


  and

  (
    g1018_p,
    g1017_n,
    g1016_n_spl_
  );


  or

  (
    g1018_n,
    g1017_p,
    g1016_p_spl_
  );


  and

  (
    g1019_p,
    g1018_p_spl_,
    g964_n_spl_
  );


  or

  (
    g1019_n,
    g1018_n_spl_,
    g964_p_spl_
  );


  and

  (
    g1020_p,
    g1018_n_spl_,
    g964_p_spl_
  );


  or

  (
    g1020_n,
    g1018_p_spl_,
    g964_n_spl_
  );


  and

  (
    g1021_p,
    g1020_n,
    g1019_n_spl_
  );


  or

  (
    g1021_n,
    g1020_p,
    g1019_p_spl_
  );


  and

  (
    g1022_p,
    g1021_p_spl_,
    g963_n_spl_
  );


  or

  (
    g1022_n,
    g1021_n_spl_,
    g963_p_spl_
  );


  and

  (
    g1023_p,
    g1021_n_spl_,
    g963_p_spl_
  );


  or

  (
    g1023_n,
    g1021_p_spl_,
    g963_n_spl_
  );


  and

  (
    g1024_p,
    g1023_n,
    g1022_n_spl_
  );


  or

  (
    g1024_n,
    g1023_p,
    g1022_p_spl_
  );


  and

  (
    g1025_p,
    g1024_p_spl_,
    g962_n_spl_
  );


  or

  (
    g1025_n,
    g1024_n_spl_,
    g962_p_spl_
  );


  and

  (
    g1026_p,
    g1024_n_spl_,
    g962_p_spl_
  );


  or

  (
    g1026_n,
    g1024_p_spl_,
    g962_n_spl_
  );


  and

  (
    g1027_p,
    g1026_n,
    g1025_n_spl_
  );


  or

  (
    g1027_n,
    g1026_p,
    g1025_p_spl_
  );


  and

  (
    g1028_p,
    g1027_p_spl_,
    g961_n_spl_
  );


  or

  (
    g1028_n,
    g1027_n_spl_,
    g961_p_spl_
  );


  and

  (
    g1029_p,
    g1027_n_spl_,
    g961_p_spl_
  );


  or

  (
    g1029_n,
    g1027_p_spl_,
    g961_n_spl_
  );


  and

  (
    g1030_p,
    g1029_n,
    g1028_n_spl_
  );


  or

  (
    g1030_n,
    g1029_p,
    g1028_p_spl_
  );


  and

  (
    g1031_p,
    g1030_p_spl_,
    g960_n_spl_
  );


  or

  (
    g1031_n,
    g1030_n_spl_,
    g960_p_spl_
  );


  and

  (
    g1032_p,
    g1030_n_spl_,
    g960_p_spl_
  );


  or

  (
    g1032_n,
    g1030_p_spl_,
    g960_n_spl_
  );


  and

  (
    g1033_p,
    g1032_n,
    g1031_n_spl_
  );


  or

  (
    g1033_n,
    g1032_p,
    g1031_p_spl_
  );


  and

  (
    g1034_p,
    g1033_p_spl_,
    g959_n_spl_
  );


  or

  (
    g1034_n,
    g1033_n_spl_,
    g959_p_spl_
  );


  and

  (
    g1035_p,
    g1033_n_spl_,
    g959_p_spl_
  );


  or

  (
    g1035_n,
    g1033_p_spl_,
    g959_n_spl_
  );


  and

  (
    g1036_p,
    g1035_n,
    g1034_n_spl_
  );


  or

  (
    g1036_n,
    g1035_p,
    g1034_p_spl_
  );


  and

  (
    g1037_p,
    g1036_p_spl_,
    g958_n_spl_
  );


  or

  (
    g1037_n,
    g1036_n_spl_,
    g958_p_spl_
  );


  and

  (
    g1038_p,
    g1036_n_spl_,
    g958_p_spl_
  );


  or

  (
    g1038_n,
    g1036_p_spl_,
    g958_n_spl_
  );


  and

  (
    g1039_p,
    g1038_n,
    g1037_n_spl_
  );


  or

  (
    g1039_n,
    g1038_p,
    g1037_p_spl_
  );


  and

  (
    g1040_p,
    g1039_p_spl_,
    g957_n_spl_
  );


  or

  (
    g1040_n,
    g1039_n_spl_,
    g957_p_spl_
  );


  and

  (
    g1041_p,
    g1039_n_spl_,
    g957_p_spl_
  );


  or

  (
    g1041_n,
    g1039_p_spl_,
    g957_n_spl_
  );


  and

  (
    g1042_p,
    g1041_n,
    g1040_n_spl_
  );


  or

  (
    g1042_n,
    g1041_p,
    g1040_p_spl_
  );


  and

  (
    g1043_p,
    g1042_p_spl_,
    g956_n_spl_
  );


  or

  (
    g1043_n,
    g1042_n_spl_,
    g956_p_spl_
  );


  and

  (
    g1044_p,
    g1042_n_spl_,
    g956_p_spl_
  );


  or

  (
    g1044_n,
    g1042_p_spl_,
    g956_n_spl_
  );


  and

  (
    g1045_p,
    g1044_n,
    g1043_n_spl_
  );


  or

  (
    g1045_n,
    g1044_p,
    g1043_p_spl_
  );


  and

  (
    g1046_p,
    g1045_p_spl_,
    g955_n_spl_
  );


  or

  (
    g1046_n,
    g1045_n_spl_,
    g955_p_spl_
  );


  and

  (
    g1047_p,
    g1045_n_spl_,
    g955_p_spl_
  );


  or

  (
    g1047_n,
    g1045_p_spl_,
    g955_n_spl_
  );


  and

  (
    g1048_p,
    g1047_n,
    g1046_n_spl_
  );


  or

  (
    g1048_n,
    g1047_p,
    g1046_p_spl_
  );


  and

  (
    g1049_p,
    g1048_p_spl_,
    g954_n_spl_
  );


  or

  (
    g1049_n,
    g1048_n_spl_,
    g954_p_spl_
  );


  and

  (
    g1050_p,
    g1048_n_spl_,
    g954_p_spl_
  );


  or

  (
    g1050_n,
    g1048_p_spl_,
    g954_n_spl_
  );


  and

  (
    g1051_p,
    g1050_n,
    g1049_n_spl_
  );


  or

  (
    g1051_n,
    g1050_p,
    g1049_p_spl_
  );


  and

  (
    g1052_p,
    g1051_p_spl_,
    g953_n_spl_
  );


  or

  (
    g1052_n,
    g1051_n_spl_,
    g953_p_spl_
  );


  and

  (
    g1053_p,
    g1051_n_spl_,
    g953_p_spl_
  );


  or

  (
    g1053_n,
    g1051_p_spl_,
    g953_n_spl_
  );


  and

  (
    g1054_p,
    g1053_n,
    g1052_n_spl_
  );


  or

  (
    g1054_n,
    g1053_p,
    g1052_p_spl_
  );


  and

  (
    g1055_p,
    g1054_p_spl_,
    g952_n_spl_
  );


  or

  (
    g1055_n,
    g1054_n_spl_,
    g952_p_spl_
  );


  and

  (
    g1056_p,
    g1054_n_spl_,
    g952_p_spl_
  );


  or

  (
    g1056_n,
    g1054_p_spl_,
    g952_n_spl_
  );


  and

  (
    g1057_p,
    g1056_n,
    g1055_n_spl_
  );


  or

  (
    g1057_n,
    g1056_p,
    g1055_p_spl_
  );


  and

  (
    g1058_p,
    g1057_p_spl_,
    g951_n_spl_
  );


  or

  (
    g1058_n,
    g1057_n_spl_,
    g951_p_spl_
  );


  and

  (
    g1059_p,
    g1057_n_spl_,
    g951_p_spl_
  );


  or

  (
    g1059_n,
    g1057_p_spl_,
    g951_n_spl_
  );


  and

  (
    g1060_p,
    g1059_n,
    g1058_n_spl_
  );


  or

  (
    g1060_n,
    g1059_p,
    g1058_p_spl_
  );


  or

  (
    g1061_n,
    g1060_n_spl_,
    g950_p_spl_
  );


  and

  (
    g1062_p,
    g1060_n_spl_,
    g950_p_spl_
  );


  or

  (
    g1062_n,
    g1060_p,
    g950_n
  );


  and

  (
    g1063_p,
    g1062_n_spl_,
    g1061_n
  );


  and

  (
    g1064_p,
    g1058_n_spl_,
    g1055_n_spl_
  );


  or

  (
    g1064_n,
    g1058_p_spl_,
    g1055_p_spl_
  );


  and

  (
    g1065_p,
    G32_p_spl_001,
    G3_p_spl_111
  );


  or

  (
    g1065_n,
    G32_n_spl_001,
    G3_n_spl_111
  );


  and

  (
    g1066_p,
    g1052_n_spl_,
    g1049_n_spl_
  );


  or

  (
    g1066_n,
    g1052_p_spl_,
    g1049_p_spl_
  );


  and

  (
    g1067_p,
    G31_p_spl_001,
    G4_p_spl_111
  );


  or

  (
    g1067_n,
    G31_n_spl_001,
    G4_n_spl_111
  );


  and

  (
    g1068_p,
    g1046_n_spl_,
    g1043_n_spl_
  );


  or

  (
    g1068_n,
    g1046_p_spl_,
    g1043_p_spl_
  );


  and

  (
    g1069_p,
    G30_p_spl_010,
    G5_p_spl_110
  );


  or

  (
    g1069_n,
    G30_n_spl_010,
    G5_n_spl_110
  );


  and

  (
    g1070_p,
    g1040_n_spl_,
    g1037_n_spl_
  );


  or

  (
    g1070_n,
    g1040_p_spl_,
    g1037_p_spl_
  );


  and

  (
    g1071_p,
    G29_p_spl_010,
    G6_p_spl_110
  );


  or

  (
    g1071_n,
    G29_n_spl_010,
    G6_n_spl_110
  );


  and

  (
    g1072_p,
    g1034_n_spl_,
    g1031_n_spl_
  );


  or

  (
    g1072_n,
    g1034_p_spl_,
    g1031_p_spl_
  );


  and

  (
    g1073_p,
    G28_p_spl_011,
    G7_p_spl_101
  );


  or

  (
    g1073_n,
    G28_n_spl_011,
    G7_n_spl_101
  );


  and

  (
    g1074_p,
    g1028_n_spl_,
    g1025_n_spl_
  );


  or

  (
    g1074_n,
    g1028_p_spl_,
    g1025_p_spl_
  );


  and

  (
    g1075_p,
    G27_p_spl_011,
    G8_p_spl_101
  );


  or

  (
    g1075_n,
    G27_n_spl_011,
    G8_n_spl_101
  );


  and

  (
    g1076_p,
    g1022_n_spl_,
    g1019_n_spl_
  );


  or

  (
    g1076_n,
    g1022_p_spl_,
    g1019_p_spl_
  );


  and

  (
    g1077_p,
    G26_p_spl_100,
    G9_p_spl_100
  );


  or

  (
    g1077_n,
    G26_n_spl_100,
    G9_n_spl_100
  );


  and

  (
    g1078_p,
    g1016_n_spl_,
    g1013_n_spl_
  );


  or

  (
    g1078_n,
    g1016_p_spl_,
    g1013_p_spl_
  );


  and

  (
    g1079_p,
    G25_p_spl_100,
    G10_p_spl_100
  );


  or

  (
    g1079_n,
    G25_n_spl_100,
    G10_n_spl_100
  );


  and

  (
    g1080_p,
    g1010_n_spl_,
    g1007_n_spl_
  );


  or

  (
    g1080_n,
    g1010_p_spl_,
    g1007_p_spl_
  );


  and

  (
    g1081_p,
    G24_p_spl_101,
    G11_p_spl_011
  );


  or

  (
    g1081_n,
    G24_n_spl_101,
    G11_n_spl_011
  );


  and

  (
    g1082_p,
    g1004_n_spl_,
    g1001_n_spl_
  );


  or

  (
    g1082_n,
    g1004_p_spl_,
    g1001_p_spl_
  );


  and

  (
    g1083_p,
    G23_p_spl_101,
    G12_p_spl_011
  );


  or

  (
    g1083_n,
    G23_n_spl_101,
    G12_n_spl_011
  );


  and

  (
    g1084_p,
    g998_n_spl_,
    g995_n_spl_
  );


  or

  (
    g1084_n,
    g998_p_spl_,
    g995_p_spl_
  );


  and

  (
    g1085_p,
    G22_p_spl_110,
    G13_p_spl_010
  );


  or

  (
    g1085_n,
    G22_n_spl_110,
    G13_n_spl_010
  );


  and

  (
    g1086_p,
    g992_n_spl_,
    g989_n_spl_
  );


  or

  (
    g1086_n,
    g992_p_spl_,
    g989_p_spl_
  );


  and

  (
    g1087_p,
    G21_p_spl_110,
    G14_p_spl_010
  );


  or

  (
    g1087_n,
    G21_n_spl_110,
    G14_n_spl_010
  );


  and

  (
    g1088_p,
    g986_n_spl_,
    g983_n_spl_
  );


  or

  (
    g1088_n,
    g986_p_spl_,
    g983_p_spl_
  );


  and

  (
    g1089_p,
    G20_p_spl_111,
    G15_p_spl_001
  );


  or

  (
    g1089_n,
    G20_n_spl_111,
    G15_n_spl_001
  );


  and

  (
    g1090_p,
    G19_p_spl_111,
    G16_p_spl_001
  );


  or

  (
    g1090_n,
    G19_n_spl_111,
    G16_n_spl_001
  );


  and

  (
    g1091_p,
    g980_n_spl_,
    g977_p_spl_
  );


  or

  (
    g1091_n,
    g980_p_spl_,
    g977_n_spl_
  );


  and

  (
    g1092_p,
    g1091_n_spl_,
    g1090_n_spl_
  );


  or

  (
    g1092_n,
    g1091_p_spl_,
    g1090_p_spl_
  );


  and

  (
    g1093_p,
    g1091_p_spl_,
    g1090_p_spl_
  );


  or

  (
    g1093_n,
    g1091_n_spl_,
    g1090_n_spl_
  );


  and

  (
    g1094_p,
    g1093_n,
    g1092_n_spl_
  );


  or

  (
    g1094_n,
    g1093_p,
    g1092_p_spl_
  );


  and

  (
    g1095_p,
    g1094_p_spl_,
    g1089_n_spl_
  );


  or

  (
    g1095_n,
    g1094_n_spl_,
    g1089_p_spl_
  );


  and

  (
    g1096_p,
    g1094_n_spl_,
    g1089_p_spl_
  );


  or

  (
    g1096_n,
    g1094_p_spl_,
    g1089_n_spl_
  );


  and

  (
    g1097_p,
    g1096_n,
    g1095_n_spl_
  );


  or

  (
    g1097_n,
    g1096_p,
    g1095_p_spl_
  );


  and

  (
    g1098_p,
    g1097_p_spl_,
    g1088_n_spl_
  );


  or

  (
    g1098_n,
    g1097_n_spl_,
    g1088_p_spl_
  );


  and

  (
    g1099_p,
    g1097_n_spl_,
    g1088_p_spl_
  );


  or

  (
    g1099_n,
    g1097_p_spl_,
    g1088_n_spl_
  );


  and

  (
    g1100_p,
    g1099_n,
    g1098_n_spl_
  );


  or

  (
    g1100_n,
    g1099_p,
    g1098_p_spl_
  );


  and

  (
    g1101_p,
    g1100_p_spl_,
    g1087_n_spl_
  );


  or

  (
    g1101_n,
    g1100_n_spl_,
    g1087_p_spl_
  );


  and

  (
    g1102_p,
    g1100_n_spl_,
    g1087_p_spl_
  );


  or

  (
    g1102_n,
    g1100_p_spl_,
    g1087_n_spl_
  );


  and

  (
    g1103_p,
    g1102_n,
    g1101_n_spl_
  );


  or

  (
    g1103_n,
    g1102_p,
    g1101_p_spl_
  );


  and

  (
    g1104_p,
    g1103_p_spl_,
    g1086_n_spl_
  );


  or

  (
    g1104_n,
    g1103_n_spl_,
    g1086_p_spl_
  );


  and

  (
    g1105_p,
    g1103_n_spl_,
    g1086_p_spl_
  );


  or

  (
    g1105_n,
    g1103_p_spl_,
    g1086_n_spl_
  );


  and

  (
    g1106_p,
    g1105_n,
    g1104_n_spl_
  );


  or

  (
    g1106_n,
    g1105_p,
    g1104_p_spl_
  );


  and

  (
    g1107_p,
    g1106_p_spl_,
    g1085_n_spl_
  );


  or

  (
    g1107_n,
    g1106_n_spl_,
    g1085_p_spl_
  );


  and

  (
    g1108_p,
    g1106_n_spl_,
    g1085_p_spl_
  );


  or

  (
    g1108_n,
    g1106_p_spl_,
    g1085_n_spl_
  );


  and

  (
    g1109_p,
    g1108_n,
    g1107_n_spl_
  );


  or

  (
    g1109_n,
    g1108_p,
    g1107_p_spl_
  );


  and

  (
    g1110_p,
    g1109_p_spl_,
    g1084_n_spl_
  );


  or

  (
    g1110_n,
    g1109_n_spl_,
    g1084_p_spl_
  );


  and

  (
    g1111_p,
    g1109_n_spl_,
    g1084_p_spl_
  );


  or

  (
    g1111_n,
    g1109_p_spl_,
    g1084_n_spl_
  );


  and

  (
    g1112_p,
    g1111_n,
    g1110_n_spl_
  );


  or

  (
    g1112_n,
    g1111_p,
    g1110_p_spl_
  );


  and

  (
    g1113_p,
    g1112_p_spl_,
    g1083_n_spl_
  );


  or

  (
    g1113_n,
    g1112_n_spl_,
    g1083_p_spl_
  );


  and

  (
    g1114_p,
    g1112_n_spl_,
    g1083_p_spl_
  );


  or

  (
    g1114_n,
    g1112_p_spl_,
    g1083_n_spl_
  );


  and

  (
    g1115_p,
    g1114_n,
    g1113_n_spl_
  );


  or

  (
    g1115_n,
    g1114_p,
    g1113_p_spl_
  );


  and

  (
    g1116_p,
    g1115_p_spl_,
    g1082_n_spl_
  );


  or

  (
    g1116_n,
    g1115_n_spl_,
    g1082_p_spl_
  );


  and

  (
    g1117_p,
    g1115_n_spl_,
    g1082_p_spl_
  );


  or

  (
    g1117_n,
    g1115_p_spl_,
    g1082_n_spl_
  );


  and

  (
    g1118_p,
    g1117_n,
    g1116_n_spl_
  );


  or

  (
    g1118_n,
    g1117_p,
    g1116_p_spl_
  );


  and

  (
    g1119_p,
    g1118_p_spl_,
    g1081_n_spl_
  );


  or

  (
    g1119_n,
    g1118_n_spl_,
    g1081_p_spl_
  );


  and

  (
    g1120_p,
    g1118_n_spl_,
    g1081_p_spl_
  );


  or

  (
    g1120_n,
    g1118_p_spl_,
    g1081_n_spl_
  );


  and

  (
    g1121_p,
    g1120_n,
    g1119_n_spl_
  );


  or

  (
    g1121_n,
    g1120_p,
    g1119_p_spl_
  );


  and

  (
    g1122_p,
    g1121_p_spl_,
    g1080_n_spl_
  );


  or

  (
    g1122_n,
    g1121_n_spl_,
    g1080_p_spl_
  );


  and

  (
    g1123_p,
    g1121_n_spl_,
    g1080_p_spl_
  );


  or

  (
    g1123_n,
    g1121_p_spl_,
    g1080_n_spl_
  );


  and

  (
    g1124_p,
    g1123_n,
    g1122_n_spl_
  );


  or

  (
    g1124_n,
    g1123_p,
    g1122_p_spl_
  );


  and

  (
    g1125_p,
    g1124_p_spl_,
    g1079_n_spl_
  );


  or

  (
    g1125_n,
    g1124_n_spl_,
    g1079_p_spl_
  );


  and

  (
    g1126_p,
    g1124_n_spl_,
    g1079_p_spl_
  );


  or

  (
    g1126_n,
    g1124_p_spl_,
    g1079_n_spl_
  );


  and

  (
    g1127_p,
    g1126_n,
    g1125_n_spl_
  );


  or

  (
    g1127_n,
    g1126_p,
    g1125_p_spl_
  );


  and

  (
    g1128_p,
    g1127_p_spl_,
    g1078_n_spl_
  );


  or

  (
    g1128_n,
    g1127_n_spl_,
    g1078_p_spl_
  );


  and

  (
    g1129_p,
    g1127_n_spl_,
    g1078_p_spl_
  );


  or

  (
    g1129_n,
    g1127_p_spl_,
    g1078_n_spl_
  );


  and

  (
    g1130_p,
    g1129_n,
    g1128_n_spl_
  );


  or

  (
    g1130_n,
    g1129_p,
    g1128_p_spl_
  );


  and

  (
    g1131_p,
    g1130_p_spl_,
    g1077_n_spl_
  );


  or

  (
    g1131_n,
    g1130_n_spl_,
    g1077_p_spl_
  );


  and

  (
    g1132_p,
    g1130_n_spl_,
    g1077_p_spl_
  );


  or

  (
    g1132_n,
    g1130_p_spl_,
    g1077_n_spl_
  );


  and

  (
    g1133_p,
    g1132_n,
    g1131_n_spl_
  );


  or

  (
    g1133_n,
    g1132_p,
    g1131_p_spl_
  );


  and

  (
    g1134_p,
    g1133_p_spl_,
    g1076_n_spl_
  );


  or

  (
    g1134_n,
    g1133_n_spl_,
    g1076_p_spl_
  );


  and

  (
    g1135_p,
    g1133_n_spl_,
    g1076_p_spl_
  );


  or

  (
    g1135_n,
    g1133_p_spl_,
    g1076_n_spl_
  );


  and

  (
    g1136_p,
    g1135_n,
    g1134_n_spl_
  );


  or

  (
    g1136_n,
    g1135_p,
    g1134_p_spl_
  );


  and

  (
    g1137_p,
    g1136_p_spl_,
    g1075_n_spl_
  );


  or

  (
    g1137_n,
    g1136_n_spl_,
    g1075_p_spl_
  );


  and

  (
    g1138_p,
    g1136_n_spl_,
    g1075_p_spl_
  );


  or

  (
    g1138_n,
    g1136_p_spl_,
    g1075_n_spl_
  );


  and

  (
    g1139_p,
    g1138_n,
    g1137_n_spl_
  );


  or

  (
    g1139_n,
    g1138_p,
    g1137_p_spl_
  );


  and

  (
    g1140_p,
    g1139_p_spl_,
    g1074_n_spl_
  );


  or

  (
    g1140_n,
    g1139_n_spl_,
    g1074_p_spl_
  );


  and

  (
    g1141_p,
    g1139_n_spl_,
    g1074_p_spl_
  );


  or

  (
    g1141_n,
    g1139_p_spl_,
    g1074_n_spl_
  );


  and

  (
    g1142_p,
    g1141_n,
    g1140_n_spl_
  );


  or

  (
    g1142_n,
    g1141_p,
    g1140_p_spl_
  );


  and

  (
    g1143_p,
    g1142_p_spl_,
    g1073_n_spl_
  );


  or

  (
    g1143_n,
    g1142_n_spl_,
    g1073_p_spl_
  );


  and

  (
    g1144_p,
    g1142_n_spl_,
    g1073_p_spl_
  );


  or

  (
    g1144_n,
    g1142_p_spl_,
    g1073_n_spl_
  );


  and

  (
    g1145_p,
    g1144_n,
    g1143_n_spl_
  );


  or

  (
    g1145_n,
    g1144_p,
    g1143_p_spl_
  );


  and

  (
    g1146_p,
    g1145_p_spl_,
    g1072_n_spl_
  );


  or

  (
    g1146_n,
    g1145_n_spl_,
    g1072_p_spl_
  );


  and

  (
    g1147_p,
    g1145_n_spl_,
    g1072_p_spl_
  );


  or

  (
    g1147_n,
    g1145_p_spl_,
    g1072_n_spl_
  );


  and

  (
    g1148_p,
    g1147_n,
    g1146_n_spl_
  );


  or

  (
    g1148_n,
    g1147_p,
    g1146_p_spl_
  );


  and

  (
    g1149_p,
    g1148_p_spl_,
    g1071_n_spl_
  );


  or

  (
    g1149_n,
    g1148_n_spl_,
    g1071_p_spl_
  );


  and

  (
    g1150_p,
    g1148_n_spl_,
    g1071_p_spl_
  );


  or

  (
    g1150_n,
    g1148_p_spl_,
    g1071_n_spl_
  );


  and

  (
    g1151_p,
    g1150_n,
    g1149_n_spl_
  );


  or

  (
    g1151_n,
    g1150_p,
    g1149_p_spl_
  );


  and

  (
    g1152_p,
    g1151_p_spl_,
    g1070_n_spl_
  );


  or

  (
    g1152_n,
    g1151_n_spl_,
    g1070_p_spl_
  );


  and

  (
    g1153_p,
    g1151_n_spl_,
    g1070_p_spl_
  );


  or

  (
    g1153_n,
    g1151_p_spl_,
    g1070_n_spl_
  );


  and

  (
    g1154_p,
    g1153_n,
    g1152_n_spl_
  );


  or

  (
    g1154_n,
    g1153_p,
    g1152_p_spl_
  );


  and

  (
    g1155_p,
    g1154_p_spl_,
    g1069_n_spl_
  );


  or

  (
    g1155_n,
    g1154_n_spl_,
    g1069_p_spl_
  );


  and

  (
    g1156_p,
    g1154_n_spl_,
    g1069_p_spl_
  );


  or

  (
    g1156_n,
    g1154_p_spl_,
    g1069_n_spl_
  );


  and

  (
    g1157_p,
    g1156_n,
    g1155_n_spl_
  );


  or

  (
    g1157_n,
    g1156_p,
    g1155_p_spl_
  );


  and

  (
    g1158_p,
    g1157_p_spl_,
    g1068_n_spl_
  );


  or

  (
    g1158_n,
    g1157_n_spl_,
    g1068_p_spl_
  );


  and

  (
    g1159_p,
    g1157_n_spl_,
    g1068_p_spl_
  );


  or

  (
    g1159_n,
    g1157_p_spl_,
    g1068_n_spl_
  );


  and

  (
    g1160_p,
    g1159_n,
    g1158_n_spl_
  );


  or

  (
    g1160_n,
    g1159_p,
    g1158_p_spl_
  );


  and

  (
    g1161_p,
    g1160_p_spl_,
    g1067_n_spl_
  );


  or

  (
    g1161_n,
    g1160_n_spl_,
    g1067_p_spl_
  );


  and

  (
    g1162_p,
    g1160_n_spl_,
    g1067_p_spl_
  );


  or

  (
    g1162_n,
    g1160_p_spl_,
    g1067_n_spl_
  );


  and

  (
    g1163_p,
    g1162_n,
    g1161_n_spl_
  );


  or

  (
    g1163_n,
    g1162_p,
    g1161_p_spl_
  );


  and

  (
    g1164_p,
    g1163_p_spl_,
    g1066_n_spl_
  );


  or

  (
    g1164_n,
    g1163_n_spl_,
    g1066_p_spl_
  );


  and

  (
    g1165_p,
    g1163_n_spl_,
    g1066_p_spl_
  );


  or

  (
    g1165_n,
    g1163_p_spl_,
    g1066_n_spl_
  );


  and

  (
    g1166_p,
    g1165_n,
    g1164_n_spl_
  );


  or

  (
    g1166_n,
    g1165_p,
    g1164_p_spl_
  );


  and

  (
    g1167_p,
    g1166_p_spl_,
    g1065_n_spl_
  );


  or

  (
    g1167_n,
    g1166_n_spl_,
    g1065_p_spl_
  );


  and

  (
    g1168_p,
    g1166_n_spl_,
    g1065_p_spl_
  );


  or

  (
    g1168_n,
    g1166_p_spl_,
    g1065_n_spl_
  );


  and

  (
    g1169_p,
    g1168_n,
    g1167_n_spl_
  );


  or

  (
    g1169_n,
    g1168_p,
    g1167_p_spl_
  );


  and

  (
    g1170_p,
    g1169_p_spl_,
    g1064_n_spl_
  );


  or

  (
    g1170_n,
    g1169_n_spl_,
    g1064_p_spl_
  );


  and

  (
    g1171_p,
    g1169_n_spl_,
    g1064_p_spl_
  );


  or

  (
    g1171_n,
    g1169_p_spl_,
    g1064_n_spl_
  );


  and

  (
    g1172_p,
    g1171_n,
    g1170_n_spl_
  );


  or

  (
    g1172_n,
    g1171_p,
    g1170_p_spl_
  );


  and

  (
    g1173_p,
    g1172_p,
    g1062_n_spl_
  );


  or

  (
    g1173_n,
    g1172_n_spl_,
    g1062_p_spl_
  );


  and

  (
    g1174_p,
    g1172_n_spl_,
    g1062_p_spl_
  );


  or

  (
    g1175_n,
    g1174_p,
    g1173_p_spl_
  );


  and

  (
    g1176_p,
    g1173_n,
    g1170_n_spl_
  );


  or

  (
    g1176_n,
    g1173_p_spl_,
    g1170_p_spl_
  );


  and

  (
    g1177_p,
    g1167_n_spl_,
    g1164_n_spl_
  );


  or

  (
    g1177_n,
    g1167_p_spl_,
    g1164_p_spl_
  );


  and

  (
    g1178_p,
    G32_p_spl_001,
    G4_p_spl_111
  );


  or

  (
    g1178_n,
    G32_n_spl_001,
    G4_n_spl_111
  );


  and

  (
    g1179_p,
    g1161_n_spl_,
    g1158_n_spl_
  );


  or

  (
    g1179_n,
    g1161_p_spl_,
    g1158_p_spl_
  );


  and

  (
    g1180_p,
    G31_p_spl_010,
    G5_p_spl_111
  );


  or

  (
    g1180_n,
    G31_n_spl_010,
    G5_n_spl_111
  );


  and

  (
    g1181_p,
    g1155_n_spl_,
    g1152_n_spl_
  );


  or

  (
    g1181_n,
    g1155_p_spl_,
    g1152_p_spl_
  );


  and

  (
    g1182_p,
    G30_p_spl_010,
    G6_p_spl_110
  );


  or

  (
    g1182_n,
    G30_n_spl_010,
    G6_n_spl_110
  );


  and

  (
    g1183_p,
    g1149_n_spl_,
    g1146_n_spl_
  );


  or

  (
    g1183_n,
    g1149_p_spl_,
    g1146_p_spl_
  );


  and

  (
    g1184_p,
    G29_p_spl_011,
    G7_p_spl_110
  );


  or

  (
    g1184_n,
    G29_n_spl_011,
    G7_n_spl_110
  );


  and

  (
    g1185_p,
    g1143_n_spl_,
    g1140_n_spl_
  );


  or

  (
    g1185_n,
    g1143_p_spl_,
    g1140_p_spl_
  );


  and

  (
    g1186_p,
    G28_p_spl_011,
    G8_p_spl_101
  );


  or

  (
    g1186_n,
    G28_n_spl_011,
    G8_n_spl_101
  );


  and

  (
    g1187_p,
    g1137_n_spl_,
    g1134_n_spl_
  );


  or

  (
    g1187_n,
    g1137_p_spl_,
    g1134_p_spl_
  );


  and

  (
    g1188_p,
    G27_p_spl_100,
    G9_p_spl_101
  );


  or

  (
    g1188_n,
    G27_n_spl_100,
    G9_n_spl_101
  );


  and

  (
    g1189_p,
    g1131_n_spl_,
    g1128_n_spl_
  );


  or

  (
    g1189_n,
    g1131_p_spl_,
    g1128_p_spl_
  );


  and

  (
    g1190_p,
    G26_p_spl_100,
    G10_p_spl_100
  );


  or

  (
    g1190_n,
    G26_n_spl_100,
    G10_n_spl_100
  );


  and

  (
    g1191_p,
    g1125_n_spl_,
    g1122_n_spl_
  );


  or

  (
    g1191_n,
    g1125_p_spl_,
    g1122_p_spl_
  );


  and

  (
    g1192_p,
    G25_p_spl_101,
    G11_p_spl_100
  );


  or

  (
    g1192_n,
    G25_n_spl_101,
    G11_n_spl_100
  );


  and

  (
    g1193_p,
    g1119_n_spl_,
    g1116_n_spl_
  );


  or

  (
    g1193_n,
    g1119_p_spl_,
    g1116_p_spl_
  );


  and

  (
    g1194_p,
    G24_p_spl_101,
    G12_p_spl_011
  );


  or

  (
    g1194_n,
    G24_n_spl_101,
    G12_n_spl_011
  );


  and

  (
    g1195_p,
    g1113_n_spl_,
    g1110_n_spl_
  );


  or

  (
    g1195_n,
    g1113_p_spl_,
    g1110_p_spl_
  );


  and

  (
    g1196_p,
    G23_p_spl_110,
    G13_p_spl_011
  );


  or

  (
    g1196_n,
    G23_n_spl_110,
    G13_n_spl_011
  );


  and

  (
    g1197_p,
    g1107_n_spl_,
    g1104_n_spl_
  );


  or

  (
    g1197_n,
    g1107_p_spl_,
    g1104_p_spl_
  );


  and

  (
    g1198_p,
    G22_p_spl_110,
    G14_p_spl_010
  );


  or

  (
    g1198_n,
    G22_n_spl_110,
    G14_n_spl_010
  );


  and

  (
    g1199_p,
    g1101_n_spl_,
    g1098_n_spl_
  );


  or

  (
    g1199_n,
    g1101_p_spl_,
    g1098_p_spl_
  );


  and

  (
    g1200_p,
    G21_p_spl_111,
    G15_p_spl_010
  );


  or

  (
    g1200_n,
    G21_n_spl_111,
    G15_n_spl_010
  );


  and

  (
    g1201_p,
    G20_p_spl_111,
    G16_p_spl_001
  );


  or

  (
    g1201_n,
    G20_n_spl_111,
    G16_n_spl_001
  );


  and

  (
    g1202_p,
    g1095_n_spl_,
    g1092_n_spl_
  );


  or

  (
    g1202_n,
    g1095_p_spl_,
    g1092_p_spl_
  );


  and

  (
    g1203_p,
    g1202_n_spl_,
    g1201_n_spl_
  );


  or

  (
    g1203_n,
    g1202_p_spl_,
    g1201_p_spl_
  );


  and

  (
    g1204_p,
    g1202_p_spl_,
    g1201_p_spl_
  );


  or

  (
    g1204_n,
    g1202_n_spl_,
    g1201_n_spl_
  );


  and

  (
    g1205_p,
    g1204_n,
    g1203_n_spl_
  );


  or

  (
    g1205_n,
    g1204_p,
    g1203_p_spl_
  );


  and

  (
    g1206_p,
    g1205_p_spl_,
    g1200_n_spl_
  );


  or

  (
    g1206_n,
    g1205_n_spl_,
    g1200_p_spl_
  );


  and

  (
    g1207_p,
    g1205_n_spl_,
    g1200_p_spl_
  );


  or

  (
    g1207_n,
    g1205_p_spl_,
    g1200_n_spl_
  );


  and

  (
    g1208_p,
    g1207_n,
    g1206_n_spl_
  );


  or

  (
    g1208_n,
    g1207_p,
    g1206_p_spl_
  );


  and

  (
    g1209_p,
    g1208_p_spl_,
    g1199_n_spl_
  );


  or

  (
    g1209_n,
    g1208_n_spl_,
    g1199_p_spl_
  );


  and

  (
    g1210_p,
    g1208_n_spl_,
    g1199_p_spl_
  );


  or

  (
    g1210_n,
    g1208_p_spl_,
    g1199_n_spl_
  );


  and

  (
    g1211_p,
    g1210_n,
    g1209_n_spl_
  );


  or

  (
    g1211_n,
    g1210_p,
    g1209_p_spl_
  );


  and

  (
    g1212_p,
    g1211_p_spl_,
    g1198_n_spl_
  );


  or

  (
    g1212_n,
    g1211_n_spl_,
    g1198_p_spl_
  );


  and

  (
    g1213_p,
    g1211_n_spl_,
    g1198_p_spl_
  );


  or

  (
    g1213_n,
    g1211_p_spl_,
    g1198_n_spl_
  );


  and

  (
    g1214_p,
    g1213_n,
    g1212_n_spl_
  );


  or

  (
    g1214_n,
    g1213_p,
    g1212_p_spl_
  );


  and

  (
    g1215_p,
    g1214_p_spl_,
    g1197_n_spl_
  );


  or

  (
    g1215_n,
    g1214_n_spl_,
    g1197_p_spl_
  );


  and

  (
    g1216_p,
    g1214_n_spl_,
    g1197_p_spl_
  );


  or

  (
    g1216_n,
    g1214_p_spl_,
    g1197_n_spl_
  );


  and

  (
    g1217_p,
    g1216_n,
    g1215_n_spl_
  );


  or

  (
    g1217_n,
    g1216_p,
    g1215_p_spl_
  );


  and

  (
    g1218_p,
    g1217_p_spl_,
    g1196_n_spl_
  );


  or

  (
    g1218_n,
    g1217_n_spl_,
    g1196_p_spl_
  );


  and

  (
    g1219_p,
    g1217_n_spl_,
    g1196_p_spl_
  );


  or

  (
    g1219_n,
    g1217_p_spl_,
    g1196_n_spl_
  );


  and

  (
    g1220_p,
    g1219_n,
    g1218_n_spl_
  );


  or

  (
    g1220_n,
    g1219_p,
    g1218_p_spl_
  );


  and

  (
    g1221_p,
    g1220_p_spl_,
    g1195_n_spl_
  );


  or

  (
    g1221_n,
    g1220_n_spl_,
    g1195_p_spl_
  );


  and

  (
    g1222_p,
    g1220_n_spl_,
    g1195_p_spl_
  );


  or

  (
    g1222_n,
    g1220_p_spl_,
    g1195_n_spl_
  );


  and

  (
    g1223_p,
    g1222_n,
    g1221_n_spl_
  );


  or

  (
    g1223_n,
    g1222_p,
    g1221_p_spl_
  );


  and

  (
    g1224_p,
    g1223_p_spl_,
    g1194_n_spl_
  );


  or

  (
    g1224_n,
    g1223_n_spl_,
    g1194_p_spl_
  );


  and

  (
    g1225_p,
    g1223_n_spl_,
    g1194_p_spl_
  );


  or

  (
    g1225_n,
    g1223_p_spl_,
    g1194_n_spl_
  );


  and

  (
    g1226_p,
    g1225_n,
    g1224_n_spl_
  );


  or

  (
    g1226_n,
    g1225_p,
    g1224_p_spl_
  );


  and

  (
    g1227_p,
    g1226_p_spl_,
    g1193_n_spl_
  );


  or

  (
    g1227_n,
    g1226_n_spl_,
    g1193_p_spl_
  );


  and

  (
    g1228_p,
    g1226_n_spl_,
    g1193_p_spl_
  );


  or

  (
    g1228_n,
    g1226_p_spl_,
    g1193_n_spl_
  );


  and

  (
    g1229_p,
    g1228_n,
    g1227_n_spl_
  );


  or

  (
    g1229_n,
    g1228_p,
    g1227_p_spl_
  );


  and

  (
    g1230_p,
    g1229_p_spl_,
    g1192_n_spl_
  );


  or

  (
    g1230_n,
    g1229_n_spl_,
    g1192_p_spl_
  );


  and

  (
    g1231_p,
    g1229_n_spl_,
    g1192_p_spl_
  );


  or

  (
    g1231_n,
    g1229_p_spl_,
    g1192_n_spl_
  );


  and

  (
    g1232_p,
    g1231_n,
    g1230_n_spl_
  );


  or

  (
    g1232_n,
    g1231_p,
    g1230_p_spl_
  );


  and

  (
    g1233_p,
    g1232_p_spl_,
    g1191_n_spl_
  );


  or

  (
    g1233_n,
    g1232_n_spl_,
    g1191_p_spl_
  );


  and

  (
    g1234_p,
    g1232_n_spl_,
    g1191_p_spl_
  );


  or

  (
    g1234_n,
    g1232_p_spl_,
    g1191_n_spl_
  );


  and

  (
    g1235_p,
    g1234_n,
    g1233_n_spl_
  );


  or

  (
    g1235_n,
    g1234_p,
    g1233_p_spl_
  );


  and

  (
    g1236_p,
    g1235_p_spl_,
    g1190_n_spl_
  );


  or

  (
    g1236_n,
    g1235_n_spl_,
    g1190_p_spl_
  );


  and

  (
    g1237_p,
    g1235_n_spl_,
    g1190_p_spl_
  );


  or

  (
    g1237_n,
    g1235_p_spl_,
    g1190_n_spl_
  );


  and

  (
    g1238_p,
    g1237_n,
    g1236_n_spl_
  );


  or

  (
    g1238_n,
    g1237_p,
    g1236_p_spl_
  );


  and

  (
    g1239_p,
    g1238_p_spl_,
    g1189_n_spl_
  );


  or

  (
    g1239_n,
    g1238_n_spl_,
    g1189_p_spl_
  );


  and

  (
    g1240_p,
    g1238_n_spl_,
    g1189_p_spl_
  );


  or

  (
    g1240_n,
    g1238_p_spl_,
    g1189_n_spl_
  );


  and

  (
    g1241_p,
    g1240_n,
    g1239_n_spl_
  );


  or

  (
    g1241_n,
    g1240_p,
    g1239_p_spl_
  );


  and

  (
    g1242_p,
    g1241_p_spl_,
    g1188_n_spl_
  );


  or

  (
    g1242_n,
    g1241_n_spl_,
    g1188_p_spl_
  );


  and

  (
    g1243_p,
    g1241_n_spl_,
    g1188_p_spl_
  );


  or

  (
    g1243_n,
    g1241_p_spl_,
    g1188_n_spl_
  );


  and

  (
    g1244_p,
    g1243_n,
    g1242_n_spl_
  );


  or

  (
    g1244_n,
    g1243_p,
    g1242_p_spl_
  );


  and

  (
    g1245_p,
    g1244_p_spl_,
    g1187_n_spl_
  );


  or

  (
    g1245_n,
    g1244_n_spl_,
    g1187_p_spl_
  );


  and

  (
    g1246_p,
    g1244_n_spl_,
    g1187_p_spl_
  );


  or

  (
    g1246_n,
    g1244_p_spl_,
    g1187_n_spl_
  );


  and

  (
    g1247_p,
    g1246_n,
    g1245_n_spl_
  );


  or

  (
    g1247_n,
    g1246_p,
    g1245_p_spl_
  );


  and

  (
    g1248_p,
    g1247_p_spl_,
    g1186_n_spl_
  );


  or

  (
    g1248_n,
    g1247_n_spl_,
    g1186_p_spl_
  );


  and

  (
    g1249_p,
    g1247_n_spl_,
    g1186_p_spl_
  );


  or

  (
    g1249_n,
    g1247_p_spl_,
    g1186_n_spl_
  );


  and

  (
    g1250_p,
    g1249_n,
    g1248_n_spl_
  );


  or

  (
    g1250_n,
    g1249_p,
    g1248_p_spl_
  );


  and

  (
    g1251_p,
    g1250_p_spl_,
    g1185_n_spl_
  );


  or

  (
    g1251_n,
    g1250_n_spl_,
    g1185_p_spl_
  );


  and

  (
    g1252_p,
    g1250_n_spl_,
    g1185_p_spl_
  );


  or

  (
    g1252_n,
    g1250_p_spl_,
    g1185_n_spl_
  );


  and

  (
    g1253_p,
    g1252_n,
    g1251_n_spl_
  );


  or

  (
    g1253_n,
    g1252_p,
    g1251_p_spl_
  );


  and

  (
    g1254_p,
    g1253_p_spl_,
    g1184_n_spl_
  );


  or

  (
    g1254_n,
    g1253_n_spl_,
    g1184_p_spl_
  );


  and

  (
    g1255_p,
    g1253_n_spl_,
    g1184_p_spl_
  );


  or

  (
    g1255_n,
    g1253_p_spl_,
    g1184_n_spl_
  );


  and

  (
    g1256_p,
    g1255_n,
    g1254_n_spl_
  );


  or

  (
    g1256_n,
    g1255_p,
    g1254_p_spl_
  );


  and

  (
    g1257_p,
    g1256_p_spl_,
    g1183_n_spl_
  );


  or

  (
    g1257_n,
    g1256_n_spl_,
    g1183_p_spl_
  );


  and

  (
    g1258_p,
    g1256_n_spl_,
    g1183_p_spl_
  );


  or

  (
    g1258_n,
    g1256_p_spl_,
    g1183_n_spl_
  );


  and

  (
    g1259_p,
    g1258_n,
    g1257_n_spl_
  );


  or

  (
    g1259_n,
    g1258_p,
    g1257_p_spl_
  );


  and

  (
    g1260_p,
    g1259_p_spl_,
    g1182_n_spl_
  );


  or

  (
    g1260_n,
    g1259_n_spl_,
    g1182_p_spl_
  );


  and

  (
    g1261_p,
    g1259_n_spl_,
    g1182_p_spl_
  );


  or

  (
    g1261_n,
    g1259_p_spl_,
    g1182_n_spl_
  );


  and

  (
    g1262_p,
    g1261_n,
    g1260_n_spl_
  );


  or

  (
    g1262_n,
    g1261_p,
    g1260_p_spl_
  );


  and

  (
    g1263_p,
    g1262_p_spl_,
    g1181_n_spl_
  );


  or

  (
    g1263_n,
    g1262_n_spl_,
    g1181_p_spl_
  );


  and

  (
    g1264_p,
    g1262_n_spl_,
    g1181_p_spl_
  );


  or

  (
    g1264_n,
    g1262_p_spl_,
    g1181_n_spl_
  );


  and

  (
    g1265_p,
    g1264_n,
    g1263_n_spl_
  );


  or

  (
    g1265_n,
    g1264_p,
    g1263_p_spl_
  );


  and

  (
    g1266_p,
    g1265_p_spl_,
    g1180_n_spl_
  );


  or

  (
    g1266_n,
    g1265_n_spl_,
    g1180_p_spl_
  );


  and

  (
    g1267_p,
    g1265_n_spl_,
    g1180_p_spl_
  );


  or

  (
    g1267_n,
    g1265_p_spl_,
    g1180_n_spl_
  );


  and

  (
    g1268_p,
    g1267_n,
    g1266_n_spl_
  );


  or

  (
    g1268_n,
    g1267_p,
    g1266_p_spl_
  );


  and

  (
    g1269_p,
    g1268_p_spl_,
    g1179_n_spl_
  );


  or

  (
    g1269_n,
    g1268_n_spl_,
    g1179_p_spl_
  );


  and

  (
    g1270_p,
    g1268_n_spl_,
    g1179_p_spl_
  );


  or

  (
    g1270_n,
    g1268_p_spl_,
    g1179_n_spl_
  );


  and

  (
    g1271_p,
    g1270_n,
    g1269_n_spl_
  );


  or

  (
    g1271_n,
    g1270_p,
    g1269_p_spl_
  );


  and

  (
    g1272_p,
    g1271_p_spl_,
    g1178_n_spl_
  );


  or

  (
    g1272_n,
    g1271_n_spl_,
    g1178_p_spl_
  );


  and

  (
    g1273_p,
    g1271_n_spl_,
    g1178_p_spl_
  );


  or

  (
    g1273_n,
    g1271_p_spl_,
    g1178_n_spl_
  );


  and

  (
    g1274_p,
    g1273_n,
    g1272_n_spl_
  );


  or

  (
    g1274_n,
    g1273_p,
    g1272_p_spl_
  );


  and

  (
    g1275_p,
    g1274_p_spl_,
    g1177_n_spl_
  );


  or

  (
    g1275_n,
    g1274_n_spl_,
    g1177_p_spl_
  );


  and

  (
    g1276_p,
    g1274_n_spl_,
    g1177_p_spl_
  );


  or

  (
    g1276_n,
    g1274_p_spl_,
    g1177_n_spl_
  );


  and

  (
    g1277_p,
    g1276_n,
    g1275_n_spl_
  );


  or

  (
    g1277_n,
    g1276_p,
    g1275_p_spl_
  );


  and

  (
    g1278_p,
    g1277_p,
    g1176_n
  );


  or

  (
    g1278_n,
    g1277_n_spl_,
    g1176_p_spl_
  );


  and

  (
    g1279_p,
    g1277_n_spl_,
    g1176_p_spl_
  );


  or

  (
    g1280_n,
    g1279_p,
    g1278_p_spl_
  );


  and

  (
    g1281_p,
    g1278_n,
    g1275_n_spl_
  );


  or

  (
    g1281_n,
    g1278_p_spl_,
    g1275_p_spl_
  );


  and

  (
    g1282_p,
    g1272_n_spl_,
    g1269_n_spl_
  );


  or

  (
    g1282_n,
    g1272_p_spl_,
    g1269_p_spl_
  );


  and

  (
    g1283_p,
    G32_p_spl_010,
    G5_p_spl_111
  );


  or

  (
    g1283_n,
    G32_n_spl_010,
    G5_n_spl_111
  );


  and

  (
    g1284_p,
    g1266_n_spl_,
    g1263_n_spl_
  );


  or

  (
    g1284_n,
    g1266_p_spl_,
    g1263_p_spl_
  );


  and

  (
    g1285_p,
    G31_p_spl_010,
    G6_p_spl_111
  );


  or

  (
    g1285_n,
    G31_n_spl_010,
    G6_n_spl_111
  );


  and

  (
    g1286_p,
    g1260_n_spl_,
    g1257_n_spl_
  );


  or

  (
    g1286_n,
    g1260_p_spl_,
    g1257_p_spl_
  );


  and

  (
    g1287_p,
    G30_p_spl_011,
    G7_p_spl_110
  );


  or

  (
    g1287_n,
    G30_n_spl_011,
    G7_n_spl_110
  );


  and

  (
    g1288_p,
    g1254_n_spl_,
    g1251_n_spl_
  );


  or

  (
    g1288_n,
    g1254_p_spl_,
    g1251_p_spl_
  );


  and

  (
    g1289_p,
    G29_p_spl_011,
    G8_p_spl_110
  );


  or

  (
    g1289_n,
    G29_n_spl_011,
    G8_n_spl_110
  );


  and

  (
    g1290_p,
    g1248_n_spl_,
    g1245_n_spl_
  );


  or

  (
    g1290_n,
    g1248_p_spl_,
    g1245_p_spl_
  );


  and

  (
    g1291_p,
    G28_p_spl_100,
    G9_p_spl_101
  );


  or

  (
    g1291_n,
    G28_n_spl_100,
    G9_n_spl_101
  );


  and

  (
    g1292_p,
    g1242_n_spl_,
    g1239_n_spl_
  );


  or

  (
    g1292_n,
    g1242_p_spl_,
    g1239_p_spl_
  );


  and

  (
    g1293_p,
    G27_p_spl_100,
    G10_p_spl_101
  );


  or

  (
    g1293_n,
    G27_n_spl_100,
    G10_n_spl_101
  );


  and

  (
    g1294_p,
    g1236_n_spl_,
    g1233_n_spl_
  );


  or

  (
    g1294_n,
    g1236_p_spl_,
    g1233_p_spl_
  );


  and

  (
    g1295_p,
    G26_p_spl_101,
    G11_p_spl_100
  );


  or

  (
    g1295_n,
    G26_n_spl_101,
    G11_n_spl_100
  );


  and

  (
    g1296_p,
    g1230_n_spl_,
    g1227_n_spl_
  );


  or

  (
    g1296_n,
    g1230_p_spl_,
    g1227_p_spl_
  );


  and

  (
    g1297_p,
    G25_p_spl_101,
    G12_p_spl_100
  );


  or

  (
    g1297_n,
    G25_n_spl_101,
    G12_n_spl_100
  );


  and

  (
    g1298_p,
    g1224_n_spl_,
    g1221_n_spl_
  );


  or

  (
    g1298_n,
    g1224_p_spl_,
    g1221_p_spl_
  );


  and

  (
    g1299_p,
    G24_p_spl_110,
    G13_p_spl_011
  );


  or

  (
    g1299_n,
    G24_n_spl_110,
    G13_n_spl_011
  );


  and

  (
    g1300_p,
    g1218_n_spl_,
    g1215_n_spl_
  );


  or

  (
    g1300_n,
    g1218_p_spl_,
    g1215_p_spl_
  );


  and

  (
    g1301_p,
    G23_p_spl_110,
    G14_p_spl_011
  );


  or

  (
    g1301_n,
    G23_n_spl_110,
    G14_n_spl_011
  );


  and

  (
    g1302_p,
    g1212_n_spl_,
    g1209_n_spl_
  );


  or

  (
    g1302_n,
    g1212_p_spl_,
    g1209_p_spl_
  );


  and

  (
    g1303_p,
    G22_p_spl_111,
    G15_p_spl_010
  );


  or

  (
    g1303_n,
    G22_n_spl_111,
    G15_n_spl_010
  );


  and

  (
    g1304_p,
    G21_p_spl_111,
    G16_p_spl_010
  );


  or

  (
    g1304_n,
    G21_n_spl_111,
    G16_n_spl_010
  );


  and

  (
    g1305_p,
    g1206_n_spl_,
    g1203_n_spl_
  );


  or

  (
    g1305_n,
    g1206_p_spl_,
    g1203_p_spl_
  );


  and

  (
    g1306_p,
    g1305_n_spl_,
    g1304_n_spl_
  );


  or

  (
    g1306_n,
    g1305_p_spl_,
    g1304_p_spl_
  );


  and

  (
    g1307_p,
    g1305_p_spl_,
    g1304_p_spl_
  );


  or

  (
    g1307_n,
    g1305_n_spl_,
    g1304_n_spl_
  );


  and

  (
    g1308_p,
    g1307_n,
    g1306_n_spl_
  );


  or

  (
    g1308_n,
    g1307_p,
    g1306_p_spl_
  );


  and

  (
    g1309_p,
    g1308_p_spl_,
    g1303_n_spl_
  );


  or

  (
    g1309_n,
    g1308_n_spl_,
    g1303_p_spl_
  );


  and

  (
    g1310_p,
    g1308_n_spl_,
    g1303_p_spl_
  );


  or

  (
    g1310_n,
    g1308_p_spl_,
    g1303_n_spl_
  );


  and

  (
    g1311_p,
    g1310_n,
    g1309_n_spl_
  );


  or

  (
    g1311_n,
    g1310_p,
    g1309_p_spl_
  );


  and

  (
    g1312_p,
    g1311_p_spl_,
    g1302_n_spl_
  );


  or

  (
    g1312_n,
    g1311_n_spl_,
    g1302_p_spl_
  );


  and

  (
    g1313_p,
    g1311_n_spl_,
    g1302_p_spl_
  );


  or

  (
    g1313_n,
    g1311_p_spl_,
    g1302_n_spl_
  );


  and

  (
    g1314_p,
    g1313_n,
    g1312_n_spl_
  );


  or

  (
    g1314_n,
    g1313_p,
    g1312_p_spl_
  );


  and

  (
    g1315_p,
    g1314_p_spl_,
    g1301_n_spl_
  );


  or

  (
    g1315_n,
    g1314_n_spl_,
    g1301_p_spl_
  );


  and

  (
    g1316_p,
    g1314_n_spl_,
    g1301_p_spl_
  );


  or

  (
    g1316_n,
    g1314_p_spl_,
    g1301_n_spl_
  );


  and

  (
    g1317_p,
    g1316_n,
    g1315_n_spl_
  );


  or

  (
    g1317_n,
    g1316_p,
    g1315_p_spl_
  );


  and

  (
    g1318_p,
    g1317_p_spl_,
    g1300_n_spl_
  );


  or

  (
    g1318_n,
    g1317_n_spl_,
    g1300_p_spl_
  );


  and

  (
    g1319_p,
    g1317_n_spl_,
    g1300_p_spl_
  );


  or

  (
    g1319_n,
    g1317_p_spl_,
    g1300_n_spl_
  );


  and

  (
    g1320_p,
    g1319_n,
    g1318_n_spl_
  );


  or

  (
    g1320_n,
    g1319_p,
    g1318_p_spl_
  );


  and

  (
    g1321_p,
    g1320_p_spl_,
    g1299_n_spl_
  );


  or

  (
    g1321_n,
    g1320_n_spl_,
    g1299_p_spl_
  );


  and

  (
    g1322_p,
    g1320_n_spl_,
    g1299_p_spl_
  );


  or

  (
    g1322_n,
    g1320_p_spl_,
    g1299_n_spl_
  );


  and

  (
    g1323_p,
    g1322_n,
    g1321_n_spl_
  );


  or

  (
    g1323_n,
    g1322_p,
    g1321_p_spl_
  );


  and

  (
    g1324_p,
    g1323_p_spl_,
    g1298_n_spl_
  );


  or

  (
    g1324_n,
    g1323_n_spl_,
    g1298_p_spl_
  );


  and

  (
    g1325_p,
    g1323_n_spl_,
    g1298_p_spl_
  );


  or

  (
    g1325_n,
    g1323_p_spl_,
    g1298_n_spl_
  );


  and

  (
    g1326_p,
    g1325_n,
    g1324_n_spl_
  );


  or

  (
    g1326_n,
    g1325_p,
    g1324_p_spl_
  );


  and

  (
    g1327_p,
    g1326_p_spl_,
    g1297_n_spl_
  );


  or

  (
    g1327_n,
    g1326_n_spl_,
    g1297_p_spl_
  );


  and

  (
    g1328_p,
    g1326_n_spl_,
    g1297_p_spl_
  );


  or

  (
    g1328_n,
    g1326_p_spl_,
    g1297_n_spl_
  );


  and

  (
    g1329_p,
    g1328_n,
    g1327_n_spl_
  );


  or

  (
    g1329_n,
    g1328_p,
    g1327_p_spl_
  );


  and

  (
    g1330_p,
    g1329_p_spl_,
    g1296_n_spl_
  );


  or

  (
    g1330_n,
    g1329_n_spl_,
    g1296_p_spl_
  );


  and

  (
    g1331_p,
    g1329_n_spl_,
    g1296_p_spl_
  );


  or

  (
    g1331_n,
    g1329_p_spl_,
    g1296_n_spl_
  );


  and

  (
    g1332_p,
    g1331_n,
    g1330_n_spl_
  );


  or

  (
    g1332_n,
    g1331_p,
    g1330_p_spl_
  );


  and

  (
    g1333_p,
    g1332_p_spl_,
    g1295_n_spl_
  );


  or

  (
    g1333_n,
    g1332_n_spl_,
    g1295_p_spl_
  );


  and

  (
    g1334_p,
    g1332_n_spl_,
    g1295_p_spl_
  );


  or

  (
    g1334_n,
    g1332_p_spl_,
    g1295_n_spl_
  );


  and

  (
    g1335_p,
    g1334_n,
    g1333_n_spl_
  );


  or

  (
    g1335_n,
    g1334_p,
    g1333_p_spl_
  );


  and

  (
    g1336_p,
    g1335_p_spl_,
    g1294_n_spl_
  );


  or

  (
    g1336_n,
    g1335_n_spl_,
    g1294_p_spl_
  );


  and

  (
    g1337_p,
    g1335_n_spl_,
    g1294_p_spl_
  );


  or

  (
    g1337_n,
    g1335_p_spl_,
    g1294_n_spl_
  );


  and

  (
    g1338_p,
    g1337_n,
    g1336_n_spl_
  );


  or

  (
    g1338_n,
    g1337_p,
    g1336_p_spl_
  );


  and

  (
    g1339_p,
    g1338_p_spl_,
    g1293_n_spl_
  );


  or

  (
    g1339_n,
    g1338_n_spl_,
    g1293_p_spl_
  );


  and

  (
    g1340_p,
    g1338_n_spl_,
    g1293_p_spl_
  );


  or

  (
    g1340_n,
    g1338_p_spl_,
    g1293_n_spl_
  );


  and

  (
    g1341_p,
    g1340_n,
    g1339_n_spl_
  );


  or

  (
    g1341_n,
    g1340_p,
    g1339_p_spl_
  );


  and

  (
    g1342_p,
    g1341_p_spl_,
    g1292_n_spl_
  );


  or

  (
    g1342_n,
    g1341_n_spl_,
    g1292_p_spl_
  );


  and

  (
    g1343_p,
    g1341_n_spl_,
    g1292_p_spl_
  );


  or

  (
    g1343_n,
    g1341_p_spl_,
    g1292_n_spl_
  );


  and

  (
    g1344_p,
    g1343_n,
    g1342_n_spl_
  );


  or

  (
    g1344_n,
    g1343_p,
    g1342_p_spl_
  );


  and

  (
    g1345_p,
    g1344_p_spl_,
    g1291_n_spl_
  );


  or

  (
    g1345_n,
    g1344_n_spl_,
    g1291_p_spl_
  );


  and

  (
    g1346_p,
    g1344_n_spl_,
    g1291_p_spl_
  );


  or

  (
    g1346_n,
    g1344_p_spl_,
    g1291_n_spl_
  );


  and

  (
    g1347_p,
    g1346_n,
    g1345_n_spl_
  );


  or

  (
    g1347_n,
    g1346_p,
    g1345_p_spl_
  );


  and

  (
    g1348_p,
    g1347_p_spl_,
    g1290_n_spl_
  );


  or

  (
    g1348_n,
    g1347_n_spl_,
    g1290_p_spl_
  );


  and

  (
    g1349_p,
    g1347_n_spl_,
    g1290_p_spl_
  );


  or

  (
    g1349_n,
    g1347_p_spl_,
    g1290_n_spl_
  );


  and

  (
    g1350_p,
    g1349_n,
    g1348_n_spl_
  );


  or

  (
    g1350_n,
    g1349_p,
    g1348_p_spl_
  );


  and

  (
    g1351_p,
    g1350_p_spl_,
    g1289_n_spl_
  );


  or

  (
    g1351_n,
    g1350_n_spl_,
    g1289_p_spl_
  );


  and

  (
    g1352_p,
    g1350_n_spl_,
    g1289_p_spl_
  );


  or

  (
    g1352_n,
    g1350_p_spl_,
    g1289_n_spl_
  );


  and

  (
    g1353_p,
    g1352_n,
    g1351_n_spl_
  );


  or

  (
    g1353_n,
    g1352_p,
    g1351_p_spl_
  );


  and

  (
    g1354_p,
    g1353_p_spl_,
    g1288_n_spl_
  );


  or

  (
    g1354_n,
    g1353_n_spl_,
    g1288_p_spl_
  );


  and

  (
    g1355_p,
    g1353_n_spl_,
    g1288_p_spl_
  );


  or

  (
    g1355_n,
    g1353_p_spl_,
    g1288_n_spl_
  );


  and

  (
    g1356_p,
    g1355_n,
    g1354_n_spl_
  );


  or

  (
    g1356_n,
    g1355_p,
    g1354_p_spl_
  );


  and

  (
    g1357_p,
    g1356_p_spl_,
    g1287_n_spl_
  );


  or

  (
    g1357_n,
    g1356_n_spl_,
    g1287_p_spl_
  );


  and

  (
    g1358_p,
    g1356_n_spl_,
    g1287_p_spl_
  );


  or

  (
    g1358_n,
    g1356_p_spl_,
    g1287_n_spl_
  );


  and

  (
    g1359_p,
    g1358_n,
    g1357_n_spl_
  );


  or

  (
    g1359_n,
    g1358_p,
    g1357_p_spl_
  );


  and

  (
    g1360_p,
    g1359_p_spl_,
    g1286_n_spl_
  );


  or

  (
    g1360_n,
    g1359_n_spl_,
    g1286_p_spl_
  );


  and

  (
    g1361_p,
    g1359_n_spl_,
    g1286_p_spl_
  );


  or

  (
    g1361_n,
    g1359_p_spl_,
    g1286_n_spl_
  );


  and

  (
    g1362_p,
    g1361_n,
    g1360_n_spl_
  );


  or

  (
    g1362_n,
    g1361_p,
    g1360_p_spl_
  );


  and

  (
    g1363_p,
    g1362_p_spl_,
    g1285_n_spl_
  );


  or

  (
    g1363_n,
    g1362_n_spl_,
    g1285_p_spl_
  );


  and

  (
    g1364_p,
    g1362_n_spl_,
    g1285_p_spl_
  );


  or

  (
    g1364_n,
    g1362_p_spl_,
    g1285_n_spl_
  );


  and

  (
    g1365_p,
    g1364_n,
    g1363_n_spl_
  );


  or

  (
    g1365_n,
    g1364_p,
    g1363_p_spl_
  );


  and

  (
    g1366_p,
    g1365_p_spl_,
    g1284_n_spl_
  );


  or

  (
    g1366_n,
    g1365_n_spl_,
    g1284_p_spl_
  );


  and

  (
    g1367_p,
    g1365_n_spl_,
    g1284_p_spl_
  );


  or

  (
    g1367_n,
    g1365_p_spl_,
    g1284_n_spl_
  );


  and

  (
    g1368_p,
    g1367_n,
    g1366_n_spl_
  );


  or

  (
    g1368_n,
    g1367_p,
    g1366_p_spl_
  );


  and

  (
    g1369_p,
    g1368_p_spl_,
    g1283_n_spl_
  );


  or

  (
    g1369_n,
    g1368_n_spl_,
    g1283_p_spl_
  );


  and

  (
    g1370_p,
    g1368_n_spl_,
    g1283_p_spl_
  );


  or

  (
    g1370_n,
    g1368_p_spl_,
    g1283_n_spl_
  );


  and

  (
    g1371_p,
    g1370_n,
    g1369_n_spl_
  );


  or

  (
    g1371_n,
    g1370_p,
    g1369_p_spl_
  );


  and

  (
    g1372_p,
    g1371_p_spl_,
    g1282_n_spl_
  );


  or

  (
    g1372_n,
    g1371_n_spl_,
    g1282_p_spl_
  );


  and

  (
    g1373_p,
    g1371_n_spl_,
    g1282_p_spl_
  );


  or

  (
    g1373_n,
    g1371_p_spl_,
    g1282_n_spl_
  );


  and

  (
    g1374_p,
    g1373_n,
    g1372_n_spl_
  );


  or

  (
    g1374_n,
    g1373_p,
    g1372_p_spl_
  );


  and

  (
    g1375_p,
    g1374_p,
    g1281_n
  );


  or

  (
    g1375_n,
    g1374_n_spl_,
    g1281_p_spl_
  );


  and

  (
    g1376_p,
    g1374_n_spl_,
    g1281_p_spl_
  );


  or

  (
    g1377_n,
    g1376_p,
    g1375_p_spl_
  );


  and

  (
    g1378_p,
    g1375_n,
    g1372_n_spl_
  );


  or

  (
    g1378_n,
    g1375_p_spl_,
    g1372_p_spl_
  );


  and

  (
    g1379_p,
    g1369_n_spl_,
    g1366_n_spl_
  );


  or

  (
    g1379_n,
    g1369_p_spl_,
    g1366_p_spl_
  );


  and

  (
    g1380_p,
    G32_p_spl_010,
    G6_p_spl_111
  );


  or

  (
    g1380_n,
    G32_n_spl_010,
    G6_n_spl_111
  );


  and

  (
    g1381_p,
    g1363_n_spl_,
    g1360_n_spl_
  );


  or

  (
    g1381_n,
    g1363_p_spl_,
    g1360_p_spl_
  );


  and

  (
    g1382_p,
    G31_p_spl_011,
    G7_p_spl_111
  );


  or

  (
    g1382_n,
    G31_n_spl_011,
    G7_n_spl_111
  );


  and

  (
    g1383_p,
    g1357_n_spl_,
    g1354_n_spl_
  );


  or

  (
    g1383_n,
    g1357_p_spl_,
    g1354_p_spl_
  );


  and

  (
    g1384_p,
    G30_p_spl_011,
    G8_p_spl_110
  );


  or

  (
    g1384_n,
    G30_n_spl_011,
    G8_n_spl_110
  );


  and

  (
    g1385_p,
    g1351_n_spl_,
    g1348_n_spl_
  );


  or

  (
    g1385_n,
    g1351_p_spl_,
    g1348_p_spl_
  );


  and

  (
    g1386_p,
    G29_p_spl_100,
    G9_p_spl_110
  );


  or

  (
    g1386_n,
    G29_n_spl_100,
    G9_n_spl_110
  );


  and

  (
    g1387_p,
    g1345_n_spl_,
    g1342_n_spl_
  );


  or

  (
    g1387_n,
    g1345_p_spl_,
    g1342_p_spl_
  );


  and

  (
    g1388_p,
    G28_p_spl_100,
    G10_p_spl_101
  );


  or

  (
    g1388_n,
    G28_n_spl_100,
    G10_n_spl_101
  );


  and

  (
    g1389_p,
    g1339_n_spl_,
    g1336_n_spl_
  );


  or

  (
    g1389_n,
    g1339_p_spl_,
    g1336_p_spl_
  );


  and

  (
    g1390_p,
    G27_p_spl_101,
    G11_p_spl_101
  );


  or

  (
    g1390_n,
    G27_n_spl_101,
    G11_n_spl_101
  );


  and

  (
    g1391_p,
    g1333_n_spl_,
    g1330_n_spl_
  );


  or

  (
    g1391_n,
    g1333_p_spl_,
    g1330_p_spl_
  );


  and

  (
    g1392_p,
    G26_p_spl_101,
    G12_p_spl_100
  );


  or

  (
    g1392_n,
    G26_n_spl_101,
    G12_n_spl_100
  );


  and

  (
    g1393_p,
    g1327_n_spl_,
    g1324_n_spl_
  );


  or

  (
    g1393_n,
    g1327_p_spl_,
    g1324_p_spl_
  );


  and

  (
    g1394_p,
    G25_p_spl_110,
    G13_p_spl_100
  );


  or

  (
    g1394_n,
    G25_n_spl_110,
    G13_n_spl_100
  );


  and

  (
    g1395_p,
    g1321_n_spl_,
    g1318_n_spl_
  );


  or

  (
    g1395_n,
    g1321_p_spl_,
    g1318_p_spl_
  );


  and

  (
    g1396_p,
    G24_p_spl_110,
    G14_p_spl_011
  );


  or

  (
    g1396_n,
    G24_n_spl_110,
    G14_n_spl_011
  );


  and

  (
    g1397_p,
    g1315_n_spl_,
    g1312_n_spl_
  );


  or

  (
    g1397_n,
    g1315_p_spl_,
    g1312_p_spl_
  );


  and

  (
    g1398_p,
    G23_p_spl_111,
    G15_p_spl_011
  );


  or

  (
    g1398_n,
    G23_n_spl_111,
    G15_n_spl_011
  );


  and

  (
    g1399_p,
    G22_p_spl_111,
    G16_p_spl_010
  );


  or

  (
    g1399_n,
    G22_n_spl_111,
    G16_n_spl_010
  );


  and

  (
    g1400_p,
    g1309_n_spl_,
    g1306_n_spl_
  );


  or

  (
    g1400_n,
    g1309_p_spl_,
    g1306_p_spl_
  );


  and

  (
    g1401_p,
    g1400_n_spl_,
    g1399_n_spl_
  );


  or

  (
    g1401_n,
    g1400_p_spl_,
    g1399_p_spl_
  );


  and

  (
    g1402_p,
    g1400_p_spl_,
    g1399_p_spl_
  );


  or

  (
    g1402_n,
    g1400_n_spl_,
    g1399_n_spl_
  );


  and

  (
    g1403_p,
    g1402_n,
    g1401_n_spl_
  );


  or

  (
    g1403_n,
    g1402_p,
    g1401_p_spl_
  );


  and

  (
    g1404_p,
    g1403_p_spl_,
    g1398_n_spl_
  );


  or

  (
    g1404_n,
    g1403_n_spl_,
    g1398_p_spl_
  );


  and

  (
    g1405_p,
    g1403_n_spl_,
    g1398_p_spl_
  );


  or

  (
    g1405_n,
    g1403_p_spl_,
    g1398_n_spl_
  );


  and

  (
    g1406_p,
    g1405_n,
    g1404_n_spl_
  );


  or

  (
    g1406_n,
    g1405_p,
    g1404_p_spl_
  );


  and

  (
    g1407_p,
    g1406_p_spl_,
    g1397_n_spl_
  );


  or

  (
    g1407_n,
    g1406_n_spl_,
    g1397_p_spl_
  );


  and

  (
    g1408_p,
    g1406_n_spl_,
    g1397_p_spl_
  );


  or

  (
    g1408_n,
    g1406_p_spl_,
    g1397_n_spl_
  );


  and

  (
    g1409_p,
    g1408_n,
    g1407_n_spl_
  );


  or

  (
    g1409_n,
    g1408_p,
    g1407_p_spl_
  );


  and

  (
    g1410_p,
    g1409_p_spl_,
    g1396_n_spl_
  );


  or

  (
    g1410_n,
    g1409_n_spl_,
    g1396_p_spl_
  );


  and

  (
    g1411_p,
    g1409_n_spl_,
    g1396_p_spl_
  );


  or

  (
    g1411_n,
    g1409_p_spl_,
    g1396_n_spl_
  );


  and

  (
    g1412_p,
    g1411_n,
    g1410_n_spl_
  );


  or

  (
    g1412_n,
    g1411_p,
    g1410_p_spl_
  );


  and

  (
    g1413_p,
    g1412_p_spl_,
    g1395_n_spl_
  );


  or

  (
    g1413_n,
    g1412_n_spl_,
    g1395_p_spl_
  );


  and

  (
    g1414_p,
    g1412_n_spl_,
    g1395_p_spl_
  );


  or

  (
    g1414_n,
    g1412_p_spl_,
    g1395_n_spl_
  );


  and

  (
    g1415_p,
    g1414_n,
    g1413_n_spl_
  );


  or

  (
    g1415_n,
    g1414_p,
    g1413_p_spl_
  );


  and

  (
    g1416_p,
    g1415_p_spl_,
    g1394_n_spl_
  );


  or

  (
    g1416_n,
    g1415_n_spl_,
    g1394_p_spl_
  );


  and

  (
    g1417_p,
    g1415_n_spl_,
    g1394_p_spl_
  );


  or

  (
    g1417_n,
    g1415_p_spl_,
    g1394_n_spl_
  );


  and

  (
    g1418_p,
    g1417_n,
    g1416_n_spl_
  );


  or

  (
    g1418_n,
    g1417_p,
    g1416_p_spl_
  );


  and

  (
    g1419_p,
    g1418_p_spl_,
    g1393_n_spl_
  );


  or

  (
    g1419_n,
    g1418_n_spl_,
    g1393_p_spl_
  );


  and

  (
    g1420_p,
    g1418_n_spl_,
    g1393_p_spl_
  );


  or

  (
    g1420_n,
    g1418_p_spl_,
    g1393_n_spl_
  );


  and

  (
    g1421_p,
    g1420_n,
    g1419_n_spl_
  );


  or

  (
    g1421_n,
    g1420_p,
    g1419_p_spl_
  );


  and

  (
    g1422_p,
    g1421_p_spl_,
    g1392_n_spl_
  );


  or

  (
    g1422_n,
    g1421_n_spl_,
    g1392_p_spl_
  );


  and

  (
    g1423_p,
    g1421_n_spl_,
    g1392_p_spl_
  );


  or

  (
    g1423_n,
    g1421_p_spl_,
    g1392_n_spl_
  );


  and

  (
    g1424_p,
    g1423_n,
    g1422_n_spl_
  );


  or

  (
    g1424_n,
    g1423_p,
    g1422_p_spl_
  );


  and

  (
    g1425_p,
    g1424_p_spl_,
    g1391_n_spl_
  );


  or

  (
    g1425_n,
    g1424_n_spl_,
    g1391_p_spl_
  );


  and

  (
    g1426_p,
    g1424_n_spl_,
    g1391_p_spl_
  );


  or

  (
    g1426_n,
    g1424_p_spl_,
    g1391_n_spl_
  );


  and

  (
    g1427_p,
    g1426_n,
    g1425_n_spl_
  );


  or

  (
    g1427_n,
    g1426_p,
    g1425_p_spl_
  );


  and

  (
    g1428_p,
    g1427_p_spl_,
    g1390_n_spl_
  );


  or

  (
    g1428_n,
    g1427_n_spl_,
    g1390_p_spl_
  );


  and

  (
    g1429_p,
    g1427_n_spl_,
    g1390_p_spl_
  );


  or

  (
    g1429_n,
    g1427_p_spl_,
    g1390_n_spl_
  );


  and

  (
    g1430_p,
    g1429_n,
    g1428_n_spl_
  );


  or

  (
    g1430_n,
    g1429_p,
    g1428_p_spl_
  );


  and

  (
    g1431_p,
    g1430_p_spl_,
    g1389_n_spl_
  );


  or

  (
    g1431_n,
    g1430_n_spl_,
    g1389_p_spl_
  );


  and

  (
    g1432_p,
    g1430_n_spl_,
    g1389_p_spl_
  );


  or

  (
    g1432_n,
    g1430_p_spl_,
    g1389_n_spl_
  );


  and

  (
    g1433_p,
    g1432_n,
    g1431_n_spl_
  );


  or

  (
    g1433_n,
    g1432_p,
    g1431_p_spl_
  );


  and

  (
    g1434_p,
    g1433_p_spl_,
    g1388_n_spl_
  );


  or

  (
    g1434_n,
    g1433_n_spl_,
    g1388_p_spl_
  );


  and

  (
    g1435_p,
    g1433_n_spl_,
    g1388_p_spl_
  );


  or

  (
    g1435_n,
    g1433_p_spl_,
    g1388_n_spl_
  );


  and

  (
    g1436_p,
    g1435_n,
    g1434_n_spl_
  );


  or

  (
    g1436_n,
    g1435_p,
    g1434_p_spl_
  );


  and

  (
    g1437_p,
    g1436_p_spl_,
    g1387_n_spl_
  );


  or

  (
    g1437_n,
    g1436_n_spl_,
    g1387_p_spl_
  );


  and

  (
    g1438_p,
    g1436_n_spl_,
    g1387_p_spl_
  );


  or

  (
    g1438_n,
    g1436_p_spl_,
    g1387_n_spl_
  );


  and

  (
    g1439_p,
    g1438_n,
    g1437_n_spl_
  );


  or

  (
    g1439_n,
    g1438_p,
    g1437_p_spl_
  );


  and

  (
    g1440_p,
    g1439_p_spl_,
    g1386_n_spl_
  );


  or

  (
    g1440_n,
    g1439_n_spl_,
    g1386_p_spl_
  );


  and

  (
    g1441_p,
    g1439_n_spl_,
    g1386_p_spl_
  );


  or

  (
    g1441_n,
    g1439_p_spl_,
    g1386_n_spl_
  );


  and

  (
    g1442_p,
    g1441_n,
    g1440_n_spl_
  );


  or

  (
    g1442_n,
    g1441_p,
    g1440_p_spl_
  );


  and

  (
    g1443_p,
    g1442_p_spl_,
    g1385_n_spl_
  );


  or

  (
    g1443_n,
    g1442_n_spl_,
    g1385_p_spl_
  );


  and

  (
    g1444_p,
    g1442_n_spl_,
    g1385_p_spl_
  );


  or

  (
    g1444_n,
    g1442_p_spl_,
    g1385_n_spl_
  );


  and

  (
    g1445_p,
    g1444_n,
    g1443_n_spl_
  );


  or

  (
    g1445_n,
    g1444_p,
    g1443_p_spl_
  );


  and

  (
    g1446_p,
    g1445_p_spl_,
    g1384_n_spl_
  );


  or

  (
    g1446_n,
    g1445_n_spl_,
    g1384_p_spl_
  );


  and

  (
    g1447_p,
    g1445_n_spl_,
    g1384_p_spl_
  );


  or

  (
    g1447_n,
    g1445_p_spl_,
    g1384_n_spl_
  );


  and

  (
    g1448_p,
    g1447_n,
    g1446_n_spl_
  );


  or

  (
    g1448_n,
    g1447_p,
    g1446_p_spl_
  );


  and

  (
    g1449_p,
    g1448_p_spl_,
    g1383_n_spl_
  );


  or

  (
    g1449_n,
    g1448_n_spl_,
    g1383_p_spl_
  );


  and

  (
    g1450_p,
    g1448_n_spl_,
    g1383_p_spl_
  );


  or

  (
    g1450_n,
    g1448_p_spl_,
    g1383_n_spl_
  );


  and

  (
    g1451_p,
    g1450_n,
    g1449_n_spl_
  );


  or

  (
    g1451_n,
    g1450_p,
    g1449_p_spl_
  );


  and

  (
    g1452_p,
    g1451_p_spl_,
    g1382_n_spl_
  );


  or

  (
    g1452_n,
    g1451_n_spl_,
    g1382_p_spl_
  );


  and

  (
    g1453_p,
    g1451_n_spl_,
    g1382_p_spl_
  );


  or

  (
    g1453_n,
    g1451_p_spl_,
    g1382_n_spl_
  );


  and

  (
    g1454_p,
    g1453_n,
    g1452_n_spl_
  );


  or

  (
    g1454_n,
    g1453_p,
    g1452_p_spl_
  );


  and

  (
    g1455_p,
    g1454_p_spl_,
    g1381_n_spl_
  );


  or

  (
    g1455_n,
    g1454_n_spl_,
    g1381_p_spl_
  );


  and

  (
    g1456_p,
    g1454_n_spl_,
    g1381_p_spl_
  );


  or

  (
    g1456_n,
    g1454_p_spl_,
    g1381_n_spl_
  );


  and

  (
    g1457_p,
    g1456_n,
    g1455_n_spl_
  );


  or

  (
    g1457_n,
    g1456_p,
    g1455_p_spl_
  );


  and

  (
    g1458_p,
    g1457_p_spl_,
    g1380_n_spl_
  );


  or

  (
    g1458_n,
    g1457_n_spl_,
    g1380_p_spl_
  );


  and

  (
    g1459_p,
    g1457_n_spl_,
    g1380_p_spl_
  );


  or

  (
    g1459_n,
    g1457_p_spl_,
    g1380_n_spl_
  );


  and

  (
    g1460_p,
    g1459_n,
    g1458_n_spl_
  );


  or

  (
    g1460_n,
    g1459_p,
    g1458_p_spl_
  );


  and

  (
    g1461_p,
    g1460_p_spl_,
    g1379_n_spl_
  );


  or

  (
    g1461_n,
    g1460_n_spl_,
    g1379_p_spl_
  );


  and

  (
    g1462_p,
    g1460_n_spl_,
    g1379_p_spl_
  );


  or

  (
    g1462_n,
    g1460_p_spl_,
    g1379_n_spl_
  );


  and

  (
    g1463_p,
    g1462_n,
    g1461_n_spl_
  );


  or

  (
    g1463_n,
    g1462_p,
    g1461_p_spl_
  );


  and

  (
    g1464_p,
    g1463_p,
    g1378_n
  );


  or

  (
    g1464_n,
    g1463_n_spl_,
    g1378_p_spl_
  );


  and

  (
    g1465_p,
    g1463_n_spl_,
    g1378_p_spl_
  );


  or

  (
    g1466_n,
    g1465_p,
    g1464_p_spl_
  );


  and

  (
    g1467_p,
    g1464_n,
    g1461_n_spl_
  );


  or

  (
    g1467_n,
    g1464_p_spl_,
    g1461_p_spl_
  );


  and

  (
    g1468_p,
    g1458_n_spl_,
    g1455_n_spl_
  );


  or

  (
    g1468_n,
    g1458_p_spl_,
    g1455_p_spl_
  );


  and

  (
    g1469_p,
    G32_p_spl_011,
    G7_p_spl_111
  );


  or

  (
    g1469_n,
    G32_n_spl_011,
    G7_n_spl_111
  );


  and

  (
    g1470_p,
    g1452_n_spl_,
    g1449_n_spl_
  );


  or

  (
    g1470_n,
    g1452_p_spl_,
    g1449_p_spl_
  );


  and

  (
    g1471_p,
    G31_p_spl_011,
    G8_p_spl_111
  );


  or

  (
    g1471_n,
    G31_n_spl_011,
    G8_n_spl_111
  );


  and

  (
    g1472_p,
    g1446_n_spl_,
    g1443_n_spl_
  );


  or

  (
    g1472_n,
    g1446_p_spl_,
    g1443_p_spl_
  );


  and

  (
    g1473_p,
    G30_p_spl_100,
    G9_p_spl_110
  );


  or

  (
    g1473_n,
    G30_n_spl_100,
    G9_n_spl_110
  );


  and

  (
    g1474_p,
    g1440_n_spl_,
    g1437_n_spl_
  );


  or

  (
    g1474_n,
    g1440_p_spl_,
    g1437_p_spl_
  );


  and

  (
    g1475_p,
    G29_p_spl_100,
    G10_p_spl_110
  );


  or

  (
    g1475_n,
    G29_n_spl_100,
    G10_n_spl_110
  );


  and

  (
    g1476_p,
    g1434_n_spl_,
    g1431_n_spl_
  );


  or

  (
    g1476_n,
    g1434_p_spl_,
    g1431_p_spl_
  );


  and

  (
    g1477_p,
    G28_p_spl_101,
    G11_p_spl_101
  );


  or

  (
    g1477_n,
    G28_n_spl_101,
    G11_n_spl_101
  );


  and

  (
    g1478_p,
    g1428_n_spl_,
    g1425_n_spl_
  );


  or

  (
    g1478_n,
    g1428_p_spl_,
    g1425_p_spl_
  );


  and

  (
    g1479_p,
    G27_p_spl_101,
    G12_p_spl_101
  );


  or

  (
    g1479_n,
    G27_n_spl_101,
    G12_n_spl_101
  );


  and

  (
    g1480_p,
    g1422_n_spl_,
    g1419_n_spl_
  );


  or

  (
    g1480_n,
    g1422_p_spl_,
    g1419_p_spl_
  );


  and

  (
    g1481_p,
    G26_p_spl_110,
    G13_p_spl_100
  );


  or

  (
    g1481_n,
    G26_n_spl_110,
    G13_n_spl_100
  );


  and

  (
    g1482_p,
    g1416_n_spl_,
    g1413_n_spl_
  );


  or

  (
    g1482_n,
    g1416_p_spl_,
    g1413_p_spl_
  );


  and

  (
    g1483_p,
    G25_p_spl_110,
    G14_p_spl_100
  );


  or

  (
    g1483_n,
    G25_n_spl_110,
    G14_n_spl_100
  );


  and

  (
    g1484_p,
    g1410_n_spl_,
    g1407_n_spl_
  );


  or

  (
    g1484_n,
    g1410_p_spl_,
    g1407_p_spl_
  );


  and

  (
    g1485_p,
    G24_p_spl_111,
    G15_p_spl_011
  );


  or

  (
    g1485_n,
    G24_n_spl_111,
    G15_n_spl_011
  );


  and

  (
    g1486_p,
    G23_p_spl_111,
    G16_p_spl_011
  );


  or

  (
    g1486_n,
    G23_n_spl_111,
    G16_n_spl_011
  );


  and

  (
    g1487_p,
    g1404_n_spl_,
    g1401_n_spl_
  );


  or

  (
    g1487_n,
    g1404_p_spl_,
    g1401_p_spl_
  );


  and

  (
    g1488_p,
    g1487_n_spl_,
    g1486_n_spl_
  );


  or

  (
    g1488_n,
    g1487_p_spl_,
    g1486_p_spl_
  );


  and

  (
    g1489_p,
    g1487_p_spl_,
    g1486_p_spl_
  );


  or

  (
    g1489_n,
    g1487_n_spl_,
    g1486_n_spl_
  );


  and

  (
    g1490_p,
    g1489_n,
    g1488_n_spl_
  );


  or

  (
    g1490_n,
    g1489_p,
    g1488_p_spl_
  );


  and

  (
    g1491_p,
    g1490_p_spl_,
    g1485_n_spl_
  );


  or

  (
    g1491_n,
    g1490_n_spl_,
    g1485_p_spl_
  );


  and

  (
    g1492_p,
    g1490_n_spl_,
    g1485_p_spl_
  );


  or

  (
    g1492_n,
    g1490_p_spl_,
    g1485_n_spl_
  );


  and

  (
    g1493_p,
    g1492_n,
    g1491_n_spl_
  );


  or

  (
    g1493_n,
    g1492_p,
    g1491_p_spl_
  );


  and

  (
    g1494_p,
    g1493_p_spl_,
    g1484_n_spl_
  );


  or

  (
    g1494_n,
    g1493_n_spl_,
    g1484_p_spl_
  );


  and

  (
    g1495_p,
    g1493_n_spl_,
    g1484_p_spl_
  );


  or

  (
    g1495_n,
    g1493_p_spl_,
    g1484_n_spl_
  );


  and

  (
    g1496_p,
    g1495_n,
    g1494_n_spl_
  );


  or

  (
    g1496_n,
    g1495_p,
    g1494_p_spl_
  );


  and

  (
    g1497_p,
    g1496_p_spl_,
    g1483_n_spl_
  );


  or

  (
    g1497_n,
    g1496_n_spl_,
    g1483_p_spl_
  );


  and

  (
    g1498_p,
    g1496_n_spl_,
    g1483_p_spl_
  );


  or

  (
    g1498_n,
    g1496_p_spl_,
    g1483_n_spl_
  );


  and

  (
    g1499_p,
    g1498_n,
    g1497_n_spl_
  );


  or

  (
    g1499_n,
    g1498_p,
    g1497_p_spl_
  );


  and

  (
    g1500_p,
    g1499_p_spl_,
    g1482_n_spl_
  );


  or

  (
    g1500_n,
    g1499_n_spl_,
    g1482_p_spl_
  );


  and

  (
    g1501_p,
    g1499_n_spl_,
    g1482_p_spl_
  );


  or

  (
    g1501_n,
    g1499_p_spl_,
    g1482_n_spl_
  );


  and

  (
    g1502_p,
    g1501_n,
    g1500_n_spl_
  );


  or

  (
    g1502_n,
    g1501_p,
    g1500_p_spl_
  );


  and

  (
    g1503_p,
    g1502_p_spl_,
    g1481_n_spl_
  );


  or

  (
    g1503_n,
    g1502_n_spl_,
    g1481_p_spl_
  );


  and

  (
    g1504_p,
    g1502_n_spl_,
    g1481_p_spl_
  );


  or

  (
    g1504_n,
    g1502_p_spl_,
    g1481_n_spl_
  );


  and

  (
    g1505_p,
    g1504_n,
    g1503_n_spl_
  );


  or

  (
    g1505_n,
    g1504_p,
    g1503_p_spl_
  );


  and

  (
    g1506_p,
    g1505_p_spl_,
    g1480_n_spl_
  );


  or

  (
    g1506_n,
    g1505_n_spl_,
    g1480_p_spl_
  );


  and

  (
    g1507_p,
    g1505_n_spl_,
    g1480_p_spl_
  );


  or

  (
    g1507_n,
    g1505_p_spl_,
    g1480_n_spl_
  );


  and

  (
    g1508_p,
    g1507_n,
    g1506_n_spl_
  );


  or

  (
    g1508_n,
    g1507_p,
    g1506_p_spl_
  );


  and

  (
    g1509_p,
    g1508_p_spl_,
    g1479_n_spl_
  );


  or

  (
    g1509_n,
    g1508_n_spl_,
    g1479_p_spl_
  );


  and

  (
    g1510_p,
    g1508_n_spl_,
    g1479_p_spl_
  );


  or

  (
    g1510_n,
    g1508_p_spl_,
    g1479_n_spl_
  );


  and

  (
    g1511_p,
    g1510_n,
    g1509_n_spl_
  );


  or

  (
    g1511_n,
    g1510_p,
    g1509_p_spl_
  );


  and

  (
    g1512_p,
    g1511_p_spl_,
    g1478_n_spl_
  );


  or

  (
    g1512_n,
    g1511_n_spl_,
    g1478_p_spl_
  );


  and

  (
    g1513_p,
    g1511_n_spl_,
    g1478_p_spl_
  );


  or

  (
    g1513_n,
    g1511_p_spl_,
    g1478_n_spl_
  );


  and

  (
    g1514_p,
    g1513_n,
    g1512_n_spl_
  );


  or

  (
    g1514_n,
    g1513_p,
    g1512_p_spl_
  );


  and

  (
    g1515_p,
    g1514_p_spl_,
    g1477_n_spl_
  );


  or

  (
    g1515_n,
    g1514_n_spl_,
    g1477_p_spl_
  );


  and

  (
    g1516_p,
    g1514_n_spl_,
    g1477_p_spl_
  );


  or

  (
    g1516_n,
    g1514_p_spl_,
    g1477_n_spl_
  );


  and

  (
    g1517_p,
    g1516_n,
    g1515_n_spl_
  );


  or

  (
    g1517_n,
    g1516_p,
    g1515_p_spl_
  );


  and

  (
    g1518_p,
    g1517_p_spl_,
    g1476_n_spl_
  );


  or

  (
    g1518_n,
    g1517_n_spl_,
    g1476_p_spl_
  );


  and

  (
    g1519_p,
    g1517_n_spl_,
    g1476_p_spl_
  );


  or

  (
    g1519_n,
    g1517_p_spl_,
    g1476_n_spl_
  );


  and

  (
    g1520_p,
    g1519_n,
    g1518_n_spl_
  );


  or

  (
    g1520_n,
    g1519_p,
    g1518_p_spl_
  );


  and

  (
    g1521_p,
    g1520_p_spl_,
    g1475_n_spl_
  );


  or

  (
    g1521_n,
    g1520_n_spl_,
    g1475_p_spl_
  );


  and

  (
    g1522_p,
    g1520_n_spl_,
    g1475_p_spl_
  );


  or

  (
    g1522_n,
    g1520_p_spl_,
    g1475_n_spl_
  );


  and

  (
    g1523_p,
    g1522_n,
    g1521_n_spl_
  );


  or

  (
    g1523_n,
    g1522_p,
    g1521_p_spl_
  );


  and

  (
    g1524_p,
    g1523_p_spl_,
    g1474_n_spl_
  );


  or

  (
    g1524_n,
    g1523_n_spl_,
    g1474_p_spl_
  );


  and

  (
    g1525_p,
    g1523_n_spl_,
    g1474_p_spl_
  );


  or

  (
    g1525_n,
    g1523_p_spl_,
    g1474_n_spl_
  );


  and

  (
    g1526_p,
    g1525_n,
    g1524_n_spl_
  );


  or

  (
    g1526_n,
    g1525_p,
    g1524_p_spl_
  );


  and

  (
    g1527_p,
    g1526_p_spl_,
    g1473_n_spl_
  );


  or

  (
    g1527_n,
    g1526_n_spl_,
    g1473_p_spl_
  );


  and

  (
    g1528_p,
    g1526_n_spl_,
    g1473_p_spl_
  );


  or

  (
    g1528_n,
    g1526_p_spl_,
    g1473_n_spl_
  );


  and

  (
    g1529_p,
    g1528_n,
    g1527_n_spl_
  );


  or

  (
    g1529_n,
    g1528_p,
    g1527_p_spl_
  );


  and

  (
    g1530_p,
    g1529_p_spl_,
    g1472_n_spl_
  );


  or

  (
    g1530_n,
    g1529_n_spl_,
    g1472_p_spl_
  );


  and

  (
    g1531_p,
    g1529_n_spl_,
    g1472_p_spl_
  );


  or

  (
    g1531_n,
    g1529_p_spl_,
    g1472_n_spl_
  );


  and

  (
    g1532_p,
    g1531_n,
    g1530_n_spl_
  );


  or

  (
    g1532_n,
    g1531_p,
    g1530_p_spl_
  );


  and

  (
    g1533_p,
    g1532_p_spl_,
    g1471_n_spl_
  );


  or

  (
    g1533_n,
    g1532_n_spl_,
    g1471_p_spl_
  );


  and

  (
    g1534_p,
    g1532_n_spl_,
    g1471_p_spl_
  );


  or

  (
    g1534_n,
    g1532_p_spl_,
    g1471_n_spl_
  );


  and

  (
    g1535_p,
    g1534_n,
    g1533_n_spl_
  );


  or

  (
    g1535_n,
    g1534_p,
    g1533_p_spl_
  );


  and

  (
    g1536_p,
    g1535_p_spl_,
    g1470_n_spl_
  );


  or

  (
    g1536_n,
    g1535_n_spl_,
    g1470_p_spl_
  );


  and

  (
    g1537_p,
    g1535_n_spl_,
    g1470_p_spl_
  );


  or

  (
    g1537_n,
    g1535_p_spl_,
    g1470_n_spl_
  );


  and

  (
    g1538_p,
    g1537_n,
    g1536_n_spl_
  );


  or

  (
    g1538_n,
    g1537_p,
    g1536_p_spl_
  );


  and

  (
    g1539_p,
    g1538_p_spl_,
    g1469_n_spl_
  );


  or

  (
    g1539_n,
    g1538_n_spl_,
    g1469_p_spl_
  );


  and

  (
    g1540_p,
    g1538_n_spl_,
    g1469_p_spl_
  );


  or

  (
    g1540_n,
    g1538_p_spl_,
    g1469_n_spl_
  );


  and

  (
    g1541_p,
    g1540_n,
    g1539_n_spl_
  );


  or

  (
    g1541_n,
    g1540_p,
    g1539_p_spl_
  );


  and

  (
    g1542_p,
    g1541_p_spl_,
    g1468_n_spl_
  );


  or

  (
    g1542_n,
    g1541_n_spl_,
    g1468_p_spl_
  );


  and

  (
    g1543_p,
    g1541_n_spl_,
    g1468_p_spl_
  );


  or

  (
    g1543_n,
    g1541_p_spl_,
    g1468_n_spl_
  );


  and

  (
    g1544_p,
    g1543_n,
    g1542_n_spl_
  );


  or

  (
    g1544_n,
    g1543_p,
    g1542_p_spl_
  );


  and

  (
    g1545_p,
    g1544_p,
    g1467_n
  );


  or

  (
    g1545_n,
    g1544_n_spl_,
    g1467_p_spl_
  );


  and

  (
    g1546_p,
    g1544_n_spl_,
    g1467_p_spl_
  );


  or

  (
    g1547_n,
    g1546_p,
    g1545_p_spl_
  );


  and

  (
    g1548_p,
    g1545_n,
    g1542_n_spl_
  );


  or

  (
    g1548_n,
    g1545_p_spl_,
    g1542_p_spl_
  );


  and

  (
    g1549_p,
    g1539_n_spl_,
    g1536_n_spl_
  );


  or

  (
    g1549_n,
    g1539_p_spl_,
    g1536_p_spl_
  );


  and

  (
    g1550_p,
    G32_p_spl_011,
    G8_p_spl_111
  );


  or

  (
    g1550_n,
    G32_n_spl_011,
    G8_n_spl_111
  );


  and

  (
    g1551_p,
    g1533_n_spl_,
    g1530_n_spl_
  );


  or

  (
    g1551_n,
    g1533_p_spl_,
    g1530_p_spl_
  );


  and

  (
    g1552_p,
    G31_p_spl_100,
    G9_p_spl_111
  );


  or

  (
    g1552_n,
    G31_n_spl_100,
    G9_n_spl_111
  );


  and

  (
    g1553_p,
    g1527_n_spl_,
    g1524_n_spl_
  );


  or

  (
    g1553_n,
    g1527_p_spl_,
    g1524_p_spl_
  );


  and

  (
    g1554_p,
    G30_p_spl_100,
    G10_p_spl_110
  );


  or

  (
    g1554_n,
    G30_n_spl_100,
    G10_n_spl_110
  );


  and

  (
    g1555_p,
    g1521_n_spl_,
    g1518_n_spl_
  );


  or

  (
    g1555_n,
    g1521_p_spl_,
    g1518_p_spl_
  );


  and

  (
    g1556_p,
    G29_p_spl_101,
    G11_p_spl_110
  );


  or

  (
    g1556_n,
    G29_n_spl_101,
    G11_n_spl_110
  );


  and

  (
    g1557_p,
    g1515_n_spl_,
    g1512_n_spl_
  );


  or

  (
    g1557_n,
    g1515_p_spl_,
    g1512_p_spl_
  );


  and

  (
    g1558_p,
    G28_p_spl_101,
    G12_p_spl_101
  );


  or

  (
    g1558_n,
    G28_n_spl_101,
    G12_n_spl_101
  );


  and

  (
    g1559_p,
    g1509_n_spl_,
    g1506_n_spl_
  );


  or

  (
    g1559_n,
    g1509_p_spl_,
    g1506_p_spl_
  );


  and

  (
    g1560_p,
    G27_p_spl_110,
    G13_p_spl_101
  );


  or

  (
    g1560_n,
    G27_n_spl_110,
    G13_n_spl_101
  );


  and

  (
    g1561_p,
    g1503_n_spl_,
    g1500_n_spl_
  );


  or

  (
    g1561_n,
    g1503_p_spl_,
    g1500_p_spl_
  );


  and

  (
    g1562_p,
    G26_p_spl_110,
    G14_p_spl_100
  );


  or

  (
    g1562_n,
    G26_n_spl_110,
    G14_n_spl_100
  );


  and

  (
    g1563_p,
    g1497_n_spl_,
    g1494_n_spl_
  );


  or

  (
    g1563_n,
    g1497_p_spl_,
    g1494_p_spl_
  );


  and

  (
    g1564_p,
    G25_p_spl_111,
    G15_p_spl_100
  );


  or

  (
    g1564_n,
    G25_n_spl_111,
    G15_n_spl_100
  );


  and

  (
    g1565_p,
    G24_p_spl_111,
    G16_p_spl_011
  );


  or

  (
    g1565_n,
    G24_n_spl_111,
    G16_n_spl_011
  );


  and

  (
    g1566_p,
    g1491_n_spl_,
    g1488_n_spl_
  );


  or

  (
    g1566_n,
    g1491_p_spl_,
    g1488_p_spl_
  );


  and

  (
    g1567_p,
    g1566_n_spl_,
    g1565_n_spl_
  );


  or

  (
    g1567_n,
    g1566_p_spl_,
    g1565_p_spl_
  );


  and

  (
    g1568_p,
    g1566_p_spl_,
    g1565_p_spl_
  );


  or

  (
    g1568_n,
    g1566_n_spl_,
    g1565_n_spl_
  );


  and

  (
    g1569_p,
    g1568_n,
    g1567_n_spl_
  );


  or

  (
    g1569_n,
    g1568_p,
    g1567_p_spl_
  );


  and

  (
    g1570_p,
    g1569_p_spl_,
    g1564_n_spl_
  );


  or

  (
    g1570_n,
    g1569_n_spl_,
    g1564_p_spl_
  );


  and

  (
    g1571_p,
    g1569_n_spl_,
    g1564_p_spl_
  );


  or

  (
    g1571_n,
    g1569_p_spl_,
    g1564_n_spl_
  );


  and

  (
    g1572_p,
    g1571_n,
    g1570_n_spl_
  );


  or

  (
    g1572_n,
    g1571_p,
    g1570_p_spl_
  );


  and

  (
    g1573_p,
    g1572_p_spl_,
    g1563_n_spl_
  );


  or

  (
    g1573_n,
    g1572_n_spl_,
    g1563_p_spl_
  );


  and

  (
    g1574_p,
    g1572_n_spl_,
    g1563_p_spl_
  );


  or

  (
    g1574_n,
    g1572_p_spl_,
    g1563_n_spl_
  );


  and

  (
    g1575_p,
    g1574_n,
    g1573_n_spl_
  );


  or

  (
    g1575_n,
    g1574_p,
    g1573_p_spl_
  );


  and

  (
    g1576_p,
    g1575_p_spl_,
    g1562_n_spl_
  );


  or

  (
    g1576_n,
    g1575_n_spl_,
    g1562_p_spl_
  );


  and

  (
    g1577_p,
    g1575_n_spl_,
    g1562_p_spl_
  );


  or

  (
    g1577_n,
    g1575_p_spl_,
    g1562_n_spl_
  );


  and

  (
    g1578_p,
    g1577_n,
    g1576_n_spl_
  );


  or

  (
    g1578_n,
    g1577_p,
    g1576_p_spl_
  );


  and

  (
    g1579_p,
    g1578_p_spl_,
    g1561_n_spl_
  );


  or

  (
    g1579_n,
    g1578_n_spl_,
    g1561_p_spl_
  );


  and

  (
    g1580_p,
    g1578_n_spl_,
    g1561_p_spl_
  );


  or

  (
    g1580_n,
    g1578_p_spl_,
    g1561_n_spl_
  );


  and

  (
    g1581_p,
    g1580_n,
    g1579_n_spl_
  );


  or

  (
    g1581_n,
    g1580_p,
    g1579_p_spl_
  );


  and

  (
    g1582_p,
    g1581_p_spl_,
    g1560_n_spl_
  );


  or

  (
    g1582_n,
    g1581_n_spl_,
    g1560_p_spl_
  );


  and

  (
    g1583_p,
    g1581_n_spl_,
    g1560_p_spl_
  );


  or

  (
    g1583_n,
    g1581_p_spl_,
    g1560_n_spl_
  );


  and

  (
    g1584_p,
    g1583_n,
    g1582_n_spl_
  );


  or

  (
    g1584_n,
    g1583_p,
    g1582_p_spl_
  );


  and

  (
    g1585_p,
    g1584_p_spl_,
    g1559_n_spl_
  );


  or

  (
    g1585_n,
    g1584_n_spl_,
    g1559_p_spl_
  );


  and

  (
    g1586_p,
    g1584_n_spl_,
    g1559_p_spl_
  );


  or

  (
    g1586_n,
    g1584_p_spl_,
    g1559_n_spl_
  );


  and

  (
    g1587_p,
    g1586_n,
    g1585_n_spl_
  );


  or

  (
    g1587_n,
    g1586_p,
    g1585_p_spl_
  );


  and

  (
    g1588_p,
    g1587_p_spl_,
    g1558_n_spl_
  );


  or

  (
    g1588_n,
    g1587_n_spl_,
    g1558_p_spl_
  );


  and

  (
    g1589_p,
    g1587_n_spl_,
    g1558_p_spl_
  );


  or

  (
    g1589_n,
    g1587_p_spl_,
    g1558_n_spl_
  );


  and

  (
    g1590_p,
    g1589_n,
    g1588_n_spl_
  );


  or

  (
    g1590_n,
    g1589_p,
    g1588_p_spl_
  );


  and

  (
    g1591_p,
    g1590_p_spl_,
    g1557_n_spl_
  );


  or

  (
    g1591_n,
    g1590_n_spl_,
    g1557_p_spl_
  );


  and

  (
    g1592_p,
    g1590_n_spl_,
    g1557_p_spl_
  );


  or

  (
    g1592_n,
    g1590_p_spl_,
    g1557_n_spl_
  );


  and

  (
    g1593_p,
    g1592_n,
    g1591_n_spl_
  );


  or

  (
    g1593_n,
    g1592_p,
    g1591_p_spl_
  );


  and

  (
    g1594_p,
    g1593_p_spl_,
    g1556_n_spl_
  );


  or

  (
    g1594_n,
    g1593_n_spl_,
    g1556_p_spl_
  );


  and

  (
    g1595_p,
    g1593_n_spl_,
    g1556_p_spl_
  );


  or

  (
    g1595_n,
    g1593_p_spl_,
    g1556_n_spl_
  );


  and

  (
    g1596_p,
    g1595_n,
    g1594_n_spl_
  );


  or

  (
    g1596_n,
    g1595_p,
    g1594_p_spl_
  );


  and

  (
    g1597_p,
    g1596_p_spl_,
    g1555_n_spl_
  );


  or

  (
    g1597_n,
    g1596_n_spl_,
    g1555_p_spl_
  );


  and

  (
    g1598_p,
    g1596_n_spl_,
    g1555_p_spl_
  );


  or

  (
    g1598_n,
    g1596_p_spl_,
    g1555_n_spl_
  );


  and

  (
    g1599_p,
    g1598_n,
    g1597_n_spl_
  );


  or

  (
    g1599_n,
    g1598_p,
    g1597_p_spl_
  );


  and

  (
    g1600_p,
    g1599_p_spl_,
    g1554_n_spl_
  );


  or

  (
    g1600_n,
    g1599_n_spl_,
    g1554_p_spl_
  );


  and

  (
    g1601_p,
    g1599_n_spl_,
    g1554_p_spl_
  );


  or

  (
    g1601_n,
    g1599_p_spl_,
    g1554_n_spl_
  );


  and

  (
    g1602_p,
    g1601_n,
    g1600_n_spl_
  );


  or

  (
    g1602_n,
    g1601_p,
    g1600_p_spl_
  );


  and

  (
    g1603_p,
    g1602_p_spl_,
    g1553_n_spl_
  );


  or

  (
    g1603_n,
    g1602_n_spl_,
    g1553_p_spl_
  );


  and

  (
    g1604_p,
    g1602_n_spl_,
    g1553_p_spl_
  );


  or

  (
    g1604_n,
    g1602_p_spl_,
    g1553_n_spl_
  );


  and

  (
    g1605_p,
    g1604_n,
    g1603_n_spl_
  );


  or

  (
    g1605_n,
    g1604_p,
    g1603_p_spl_
  );


  and

  (
    g1606_p,
    g1605_p_spl_,
    g1552_n_spl_
  );


  or

  (
    g1606_n,
    g1605_n_spl_,
    g1552_p_spl_
  );


  and

  (
    g1607_p,
    g1605_n_spl_,
    g1552_p_spl_
  );


  or

  (
    g1607_n,
    g1605_p_spl_,
    g1552_n_spl_
  );


  and

  (
    g1608_p,
    g1607_n,
    g1606_n_spl_
  );


  or

  (
    g1608_n,
    g1607_p,
    g1606_p_spl_
  );


  and

  (
    g1609_p,
    g1608_p_spl_,
    g1551_n_spl_
  );


  or

  (
    g1609_n,
    g1608_n_spl_,
    g1551_p_spl_
  );


  and

  (
    g1610_p,
    g1608_n_spl_,
    g1551_p_spl_
  );


  or

  (
    g1610_n,
    g1608_p_spl_,
    g1551_n_spl_
  );


  and

  (
    g1611_p,
    g1610_n,
    g1609_n_spl_
  );


  or

  (
    g1611_n,
    g1610_p,
    g1609_p_spl_
  );


  and

  (
    g1612_p,
    g1611_p_spl_,
    g1550_n_spl_
  );


  or

  (
    g1612_n,
    g1611_n_spl_,
    g1550_p_spl_
  );


  and

  (
    g1613_p,
    g1611_n_spl_,
    g1550_p_spl_
  );


  or

  (
    g1613_n,
    g1611_p_spl_,
    g1550_n_spl_
  );


  and

  (
    g1614_p,
    g1613_n,
    g1612_n_spl_
  );


  or

  (
    g1614_n,
    g1613_p,
    g1612_p_spl_
  );


  and

  (
    g1615_p,
    g1614_p_spl_,
    g1549_n_spl_
  );


  or

  (
    g1615_n,
    g1614_n_spl_,
    g1549_p_spl_
  );


  and

  (
    g1616_p,
    g1614_n_spl_,
    g1549_p_spl_
  );


  or

  (
    g1616_n,
    g1614_p_spl_,
    g1549_n_spl_
  );


  and

  (
    g1617_p,
    g1616_n,
    g1615_n_spl_
  );


  or

  (
    g1617_n,
    g1616_p,
    g1615_p_spl_
  );


  and

  (
    g1618_p,
    g1617_p,
    g1548_n
  );


  or

  (
    g1618_n,
    g1617_n_spl_,
    g1548_p_spl_
  );


  and

  (
    g1619_p,
    g1617_n_spl_,
    g1548_p_spl_
  );


  or

  (
    g1620_n,
    g1619_p,
    g1618_p_spl_
  );


  and

  (
    g1621_p,
    g1618_n,
    g1615_n_spl_
  );


  or

  (
    g1621_n,
    g1618_p_spl_,
    g1615_p_spl_
  );


  and

  (
    g1622_p,
    g1612_n_spl_,
    g1609_n_spl_
  );


  or

  (
    g1622_n,
    g1612_p_spl_,
    g1609_p_spl_
  );


  and

  (
    g1623_p,
    G32_p_spl_100,
    G9_p_spl_111
  );


  or

  (
    g1623_n,
    G32_n_spl_100,
    G9_n_spl_111
  );


  and

  (
    g1624_p,
    g1606_n_spl_,
    g1603_n_spl_
  );


  or

  (
    g1624_n,
    g1606_p_spl_,
    g1603_p_spl_
  );


  and

  (
    g1625_p,
    G31_p_spl_100,
    G10_p_spl_111
  );


  or

  (
    g1625_n,
    G31_n_spl_100,
    G10_n_spl_111
  );


  and

  (
    g1626_p,
    g1600_n_spl_,
    g1597_n_spl_
  );


  or

  (
    g1626_n,
    g1600_p_spl_,
    g1597_p_spl_
  );


  and

  (
    g1627_p,
    G30_p_spl_101,
    G11_p_spl_110
  );


  or

  (
    g1627_n,
    G30_n_spl_101,
    G11_n_spl_110
  );


  and

  (
    g1628_p,
    g1594_n_spl_,
    g1591_n_spl_
  );


  or

  (
    g1628_n,
    g1594_p_spl_,
    g1591_p_spl_
  );


  and

  (
    g1629_p,
    G29_p_spl_101,
    G12_p_spl_110
  );


  or

  (
    g1629_n,
    G29_n_spl_101,
    G12_n_spl_110
  );


  and

  (
    g1630_p,
    g1588_n_spl_,
    g1585_n_spl_
  );


  or

  (
    g1630_n,
    g1588_p_spl_,
    g1585_p_spl_
  );


  and

  (
    g1631_p,
    G28_p_spl_110,
    G13_p_spl_101
  );


  or

  (
    g1631_n,
    G28_n_spl_110,
    G13_n_spl_101
  );


  and

  (
    g1632_p,
    g1582_n_spl_,
    g1579_n_spl_
  );


  or

  (
    g1632_n,
    g1582_p_spl_,
    g1579_p_spl_
  );


  and

  (
    g1633_p,
    G27_p_spl_110,
    G14_p_spl_101
  );


  or

  (
    g1633_n,
    G27_n_spl_110,
    G14_n_spl_101
  );


  and

  (
    g1634_p,
    g1576_n_spl_,
    g1573_n_spl_
  );


  or

  (
    g1634_n,
    g1576_p_spl_,
    g1573_p_spl_
  );


  and

  (
    g1635_p,
    G26_p_spl_111,
    G15_p_spl_100
  );


  or

  (
    g1635_n,
    G26_n_spl_111,
    G15_n_spl_100
  );


  and

  (
    g1636_p,
    G25_p_spl_111,
    G16_p_spl_100
  );


  or

  (
    g1636_n,
    G25_n_spl_111,
    G16_n_spl_100
  );


  and

  (
    g1637_p,
    g1570_n_spl_,
    g1567_n_spl_
  );


  or

  (
    g1637_n,
    g1570_p_spl_,
    g1567_p_spl_
  );


  and

  (
    g1638_p,
    g1637_n_spl_,
    g1636_n_spl_
  );


  or

  (
    g1638_n,
    g1637_p_spl_,
    g1636_p_spl_
  );


  and

  (
    g1639_p,
    g1637_p_spl_,
    g1636_p_spl_
  );


  or

  (
    g1639_n,
    g1637_n_spl_,
    g1636_n_spl_
  );


  and

  (
    g1640_p,
    g1639_n,
    g1638_n_spl_
  );


  or

  (
    g1640_n,
    g1639_p,
    g1638_p_spl_
  );


  and

  (
    g1641_p,
    g1640_p_spl_,
    g1635_n_spl_
  );


  or

  (
    g1641_n,
    g1640_n_spl_,
    g1635_p_spl_
  );


  and

  (
    g1642_p,
    g1640_n_spl_,
    g1635_p_spl_
  );


  or

  (
    g1642_n,
    g1640_p_spl_,
    g1635_n_spl_
  );


  and

  (
    g1643_p,
    g1642_n,
    g1641_n_spl_
  );


  or

  (
    g1643_n,
    g1642_p,
    g1641_p_spl_
  );


  and

  (
    g1644_p,
    g1643_p_spl_,
    g1634_n_spl_
  );


  or

  (
    g1644_n,
    g1643_n_spl_,
    g1634_p_spl_
  );


  and

  (
    g1645_p,
    g1643_n_spl_,
    g1634_p_spl_
  );


  or

  (
    g1645_n,
    g1643_p_spl_,
    g1634_n_spl_
  );


  and

  (
    g1646_p,
    g1645_n,
    g1644_n_spl_
  );


  or

  (
    g1646_n,
    g1645_p,
    g1644_p_spl_
  );


  and

  (
    g1647_p,
    g1646_p_spl_,
    g1633_n_spl_
  );


  or

  (
    g1647_n,
    g1646_n_spl_,
    g1633_p_spl_
  );


  and

  (
    g1648_p,
    g1646_n_spl_,
    g1633_p_spl_
  );


  or

  (
    g1648_n,
    g1646_p_spl_,
    g1633_n_spl_
  );


  and

  (
    g1649_p,
    g1648_n,
    g1647_n_spl_
  );


  or

  (
    g1649_n,
    g1648_p,
    g1647_p_spl_
  );


  and

  (
    g1650_p,
    g1649_p_spl_,
    g1632_n_spl_
  );


  or

  (
    g1650_n,
    g1649_n_spl_,
    g1632_p_spl_
  );


  and

  (
    g1651_p,
    g1649_n_spl_,
    g1632_p_spl_
  );


  or

  (
    g1651_n,
    g1649_p_spl_,
    g1632_n_spl_
  );


  and

  (
    g1652_p,
    g1651_n,
    g1650_n_spl_
  );


  or

  (
    g1652_n,
    g1651_p,
    g1650_p_spl_
  );


  and

  (
    g1653_p,
    g1652_p_spl_,
    g1631_n_spl_
  );


  or

  (
    g1653_n,
    g1652_n_spl_,
    g1631_p_spl_
  );


  and

  (
    g1654_p,
    g1652_n_spl_,
    g1631_p_spl_
  );


  or

  (
    g1654_n,
    g1652_p_spl_,
    g1631_n_spl_
  );


  and

  (
    g1655_p,
    g1654_n,
    g1653_n_spl_
  );


  or

  (
    g1655_n,
    g1654_p,
    g1653_p_spl_
  );


  and

  (
    g1656_p,
    g1655_p_spl_,
    g1630_n_spl_
  );


  or

  (
    g1656_n,
    g1655_n_spl_,
    g1630_p_spl_
  );


  and

  (
    g1657_p,
    g1655_n_spl_,
    g1630_p_spl_
  );


  or

  (
    g1657_n,
    g1655_p_spl_,
    g1630_n_spl_
  );


  and

  (
    g1658_p,
    g1657_n,
    g1656_n_spl_
  );


  or

  (
    g1658_n,
    g1657_p,
    g1656_p_spl_
  );


  and

  (
    g1659_p,
    g1658_p_spl_,
    g1629_n_spl_
  );


  or

  (
    g1659_n,
    g1658_n_spl_,
    g1629_p_spl_
  );


  and

  (
    g1660_p,
    g1658_n_spl_,
    g1629_p_spl_
  );


  or

  (
    g1660_n,
    g1658_p_spl_,
    g1629_n_spl_
  );


  and

  (
    g1661_p,
    g1660_n,
    g1659_n_spl_
  );


  or

  (
    g1661_n,
    g1660_p,
    g1659_p_spl_
  );


  and

  (
    g1662_p,
    g1661_p_spl_,
    g1628_n_spl_
  );


  or

  (
    g1662_n,
    g1661_n_spl_,
    g1628_p_spl_
  );


  and

  (
    g1663_p,
    g1661_n_spl_,
    g1628_p_spl_
  );


  or

  (
    g1663_n,
    g1661_p_spl_,
    g1628_n_spl_
  );


  and

  (
    g1664_p,
    g1663_n,
    g1662_n_spl_
  );


  or

  (
    g1664_n,
    g1663_p,
    g1662_p_spl_
  );


  and

  (
    g1665_p,
    g1664_p_spl_,
    g1627_n_spl_
  );


  or

  (
    g1665_n,
    g1664_n_spl_,
    g1627_p_spl_
  );


  and

  (
    g1666_p,
    g1664_n_spl_,
    g1627_p_spl_
  );


  or

  (
    g1666_n,
    g1664_p_spl_,
    g1627_n_spl_
  );


  and

  (
    g1667_p,
    g1666_n,
    g1665_n_spl_
  );


  or

  (
    g1667_n,
    g1666_p,
    g1665_p_spl_
  );


  and

  (
    g1668_p,
    g1667_p_spl_,
    g1626_n_spl_
  );


  or

  (
    g1668_n,
    g1667_n_spl_,
    g1626_p_spl_
  );


  and

  (
    g1669_p,
    g1667_n_spl_,
    g1626_p_spl_
  );


  or

  (
    g1669_n,
    g1667_p_spl_,
    g1626_n_spl_
  );


  and

  (
    g1670_p,
    g1669_n,
    g1668_n_spl_
  );


  or

  (
    g1670_n,
    g1669_p,
    g1668_p_spl_
  );


  and

  (
    g1671_p,
    g1670_p_spl_,
    g1625_n_spl_
  );


  or

  (
    g1671_n,
    g1670_n_spl_,
    g1625_p_spl_
  );


  and

  (
    g1672_p,
    g1670_n_spl_,
    g1625_p_spl_
  );


  or

  (
    g1672_n,
    g1670_p_spl_,
    g1625_n_spl_
  );


  and

  (
    g1673_p,
    g1672_n,
    g1671_n_spl_
  );


  or

  (
    g1673_n,
    g1672_p,
    g1671_p_spl_
  );


  and

  (
    g1674_p,
    g1673_p_spl_,
    g1624_n_spl_
  );


  or

  (
    g1674_n,
    g1673_n_spl_,
    g1624_p_spl_
  );


  and

  (
    g1675_p,
    g1673_n_spl_,
    g1624_p_spl_
  );


  or

  (
    g1675_n,
    g1673_p_spl_,
    g1624_n_spl_
  );


  and

  (
    g1676_p,
    g1675_n,
    g1674_n_spl_
  );


  or

  (
    g1676_n,
    g1675_p,
    g1674_p_spl_
  );


  and

  (
    g1677_p,
    g1676_p_spl_,
    g1623_n_spl_
  );


  or

  (
    g1677_n,
    g1676_n_spl_,
    g1623_p_spl_
  );


  and

  (
    g1678_p,
    g1676_n_spl_,
    g1623_p_spl_
  );


  or

  (
    g1678_n,
    g1676_p_spl_,
    g1623_n_spl_
  );


  and

  (
    g1679_p,
    g1678_n,
    g1677_n_spl_
  );


  or

  (
    g1679_n,
    g1678_p,
    g1677_p_spl_
  );


  and

  (
    g1680_p,
    g1679_p_spl_,
    g1622_n_spl_
  );


  or

  (
    g1680_n,
    g1679_n_spl_,
    g1622_p_spl_
  );


  and

  (
    g1681_p,
    g1679_n_spl_,
    g1622_p_spl_
  );


  or

  (
    g1681_n,
    g1679_p_spl_,
    g1622_n_spl_
  );


  and

  (
    g1682_p,
    g1681_n,
    g1680_n_spl_
  );


  or

  (
    g1682_n,
    g1681_p,
    g1680_p_spl_
  );


  and

  (
    g1683_p,
    g1682_p,
    g1621_n
  );


  or

  (
    g1683_n,
    g1682_n_spl_,
    g1621_p_spl_
  );


  and

  (
    g1684_p,
    g1682_n_spl_,
    g1621_p_spl_
  );


  or

  (
    g1685_n,
    g1684_p,
    g1683_p_spl_
  );


  and

  (
    g1686_p,
    g1683_n,
    g1680_n_spl_
  );


  or

  (
    g1686_n,
    g1683_p_spl_,
    g1680_p_spl_
  );


  and

  (
    g1687_p,
    g1677_n_spl_,
    g1674_n_spl_
  );


  or

  (
    g1687_n,
    g1677_p_spl_,
    g1674_p_spl_
  );


  and

  (
    g1688_p,
    G32_p_spl_100,
    G10_p_spl_111
  );


  or

  (
    g1688_n,
    G32_n_spl_100,
    G10_n_spl_111
  );


  and

  (
    g1689_p,
    g1671_n_spl_,
    g1668_n_spl_
  );


  or

  (
    g1689_n,
    g1671_p_spl_,
    g1668_p_spl_
  );


  and

  (
    g1690_p,
    G31_p_spl_101,
    G11_p_spl_111
  );


  or

  (
    g1690_n,
    G31_n_spl_101,
    G11_n_spl_111
  );


  and

  (
    g1691_p,
    g1665_n_spl_,
    g1662_n_spl_
  );


  or

  (
    g1691_n,
    g1665_p_spl_,
    g1662_p_spl_
  );


  and

  (
    g1692_p,
    G30_p_spl_101,
    G12_p_spl_110
  );


  or

  (
    g1692_n,
    G30_n_spl_101,
    G12_n_spl_110
  );


  and

  (
    g1693_p,
    g1659_n_spl_,
    g1656_n_spl_
  );


  or

  (
    g1693_n,
    g1659_p_spl_,
    g1656_p_spl_
  );


  and

  (
    g1694_p,
    G29_p_spl_110,
    G13_p_spl_110
  );


  or

  (
    g1694_n,
    G29_n_spl_110,
    G13_n_spl_110
  );


  and

  (
    g1695_p,
    g1653_n_spl_,
    g1650_n_spl_
  );


  or

  (
    g1695_n,
    g1653_p_spl_,
    g1650_p_spl_
  );


  and

  (
    g1696_p,
    G28_p_spl_110,
    G14_p_spl_101
  );


  or

  (
    g1696_n,
    G28_n_spl_110,
    G14_n_spl_101
  );


  and

  (
    g1697_p,
    g1647_n_spl_,
    g1644_n_spl_
  );


  or

  (
    g1697_n,
    g1647_p_spl_,
    g1644_p_spl_
  );


  and

  (
    g1698_p,
    G27_p_spl_111,
    G15_p_spl_101
  );


  or

  (
    g1698_n,
    G27_n_spl_111,
    G15_n_spl_101
  );


  and

  (
    g1699_p,
    G26_p_spl_111,
    G16_p_spl_100
  );


  or

  (
    g1699_n,
    G26_n_spl_111,
    G16_n_spl_100
  );


  and

  (
    g1700_p,
    g1641_n_spl_,
    g1638_n_spl_
  );


  or

  (
    g1700_n,
    g1641_p_spl_,
    g1638_p_spl_
  );


  and

  (
    g1701_p,
    g1700_n_spl_,
    g1699_n_spl_
  );


  or

  (
    g1701_n,
    g1700_p_spl_,
    g1699_p_spl_
  );


  and

  (
    g1702_p,
    g1700_p_spl_,
    g1699_p_spl_
  );


  or

  (
    g1702_n,
    g1700_n_spl_,
    g1699_n_spl_
  );


  and

  (
    g1703_p,
    g1702_n,
    g1701_n_spl_
  );


  or

  (
    g1703_n,
    g1702_p,
    g1701_p_spl_
  );


  and

  (
    g1704_p,
    g1703_p_spl_,
    g1698_n_spl_
  );


  or

  (
    g1704_n,
    g1703_n_spl_,
    g1698_p_spl_
  );


  and

  (
    g1705_p,
    g1703_n_spl_,
    g1698_p_spl_
  );


  or

  (
    g1705_n,
    g1703_p_spl_,
    g1698_n_spl_
  );


  and

  (
    g1706_p,
    g1705_n,
    g1704_n_spl_
  );


  or

  (
    g1706_n,
    g1705_p,
    g1704_p_spl_
  );


  and

  (
    g1707_p,
    g1706_p_spl_,
    g1697_n_spl_
  );


  or

  (
    g1707_n,
    g1706_n_spl_,
    g1697_p_spl_
  );


  and

  (
    g1708_p,
    g1706_n_spl_,
    g1697_p_spl_
  );


  or

  (
    g1708_n,
    g1706_p_spl_,
    g1697_n_spl_
  );


  and

  (
    g1709_p,
    g1708_n,
    g1707_n_spl_
  );


  or

  (
    g1709_n,
    g1708_p,
    g1707_p_spl_
  );


  and

  (
    g1710_p,
    g1709_p_spl_,
    g1696_n_spl_
  );


  or

  (
    g1710_n,
    g1709_n_spl_,
    g1696_p_spl_
  );


  and

  (
    g1711_p,
    g1709_n_spl_,
    g1696_p_spl_
  );


  or

  (
    g1711_n,
    g1709_p_spl_,
    g1696_n_spl_
  );


  and

  (
    g1712_p,
    g1711_n,
    g1710_n_spl_
  );


  or

  (
    g1712_n,
    g1711_p,
    g1710_p_spl_
  );


  and

  (
    g1713_p,
    g1712_p_spl_,
    g1695_n_spl_
  );


  or

  (
    g1713_n,
    g1712_n_spl_,
    g1695_p_spl_
  );


  and

  (
    g1714_p,
    g1712_n_spl_,
    g1695_p_spl_
  );


  or

  (
    g1714_n,
    g1712_p_spl_,
    g1695_n_spl_
  );


  and

  (
    g1715_p,
    g1714_n,
    g1713_n_spl_
  );


  or

  (
    g1715_n,
    g1714_p,
    g1713_p_spl_
  );


  and

  (
    g1716_p,
    g1715_p_spl_,
    g1694_n_spl_
  );


  or

  (
    g1716_n,
    g1715_n_spl_,
    g1694_p_spl_
  );


  and

  (
    g1717_p,
    g1715_n_spl_,
    g1694_p_spl_
  );


  or

  (
    g1717_n,
    g1715_p_spl_,
    g1694_n_spl_
  );


  and

  (
    g1718_p,
    g1717_n,
    g1716_n_spl_
  );


  or

  (
    g1718_n,
    g1717_p,
    g1716_p_spl_
  );


  and

  (
    g1719_p,
    g1718_p_spl_,
    g1693_n_spl_
  );


  or

  (
    g1719_n,
    g1718_n_spl_,
    g1693_p_spl_
  );


  and

  (
    g1720_p,
    g1718_n_spl_,
    g1693_p_spl_
  );


  or

  (
    g1720_n,
    g1718_p_spl_,
    g1693_n_spl_
  );


  and

  (
    g1721_p,
    g1720_n,
    g1719_n_spl_
  );


  or

  (
    g1721_n,
    g1720_p,
    g1719_p_spl_
  );


  and

  (
    g1722_p,
    g1721_p_spl_,
    g1692_n_spl_
  );


  or

  (
    g1722_n,
    g1721_n_spl_,
    g1692_p_spl_
  );


  and

  (
    g1723_p,
    g1721_n_spl_,
    g1692_p_spl_
  );


  or

  (
    g1723_n,
    g1721_p_spl_,
    g1692_n_spl_
  );


  and

  (
    g1724_p,
    g1723_n,
    g1722_n_spl_
  );


  or

  (
    g1724_n,
    g1723_p,
    g1722_p_spl_
  );


  and

  (
    g1725_p,
    g1724_p_spl_,
    g1691_n_spl_
  );


  or

  (
    g1725_n,
    g1724_n_spl_,
    g1691_p_spl_
  );


  and

  (
    g1726_p,
    g1724_n_spl_,
    g1691_p_spl_
  );


  or

  (
    g1726_n,
    g1724_p_spl_,
    g1691_n_spl_
  );


  and

  (
    g1727_p,
    g1726_n,
    g1725_n_spl_
  );


  or

  (
    g1727_n,
    g1726_p,
    g1725_p_spl_
  );


  and

  (
    g1728_p,
    g1727_p_spl_,
    g1690_n_spl_
  );


  or

  (
    g1728_n,
    g1727_n_spl_,
    g1690_p_spl_
  );


  and

  (
    g1729_p,
    g1727_n_spl_,
    g1690_p_spl_
  );


  or

  (
    g1729_n,
    g1727_p_spl_,
    g1690_n_spl_
  );


  and

  (
    g1730_p,
    g1729_n,
    g1728_n_spl_
  );


  or

  (
    g1730_n,
    g1729_p,
    g1728_p_spl_
  );


  and

  (
    g1731_p,
    g1730_p_spl_,
    g1689_n_spl_
  );


  or

  (
    g1731_n,
    g1730_n_spl_,
    g1689_p_spl_
  );


  and

  (
    g1732_p,
    g1730_n_spl_,
    g1689_p_spl_
  );


  or

  (
    g1732_n,
    g1730_p_spl_,
    g1689_n_spl_
  );


  and

  (
    g1733_p,
    g1732_n,
    g1731_n_spl_
  );


  or

  (
    g1733_n,
    g1732_p,
    g1731_p_spl_
  );


  and

  (
    g1734_p,
    g1733_p_spl_,
    g1688_n_spl_
  );


  or

  (
    g1734_n,
    g1733_n_spl_,
    g1688_p_spl_
  );


  and

  (
    g1735_p,
    g1733_n_spl_,
    g1688_p_spl_
  );


  or

  (
    g1735_n,
    g1733_p_spl_,
    g1688_n_spl_
  );


  and

  (
    g1736_p,
    g1735_n,
    g1734_n_spl_
  );


  or

  (
    g1736_n,
    g1735_p,
    g1734_p_spl_
  );


  and

  (
    g1737_p,
    g1736_p_spl_,
    g1687_n_spl_
  );


  or

  (
    g1737_n,
    g1736_n_spl_,
    g1687_p_spl_
  );


  and

  (
    g1738_p,
    g1736_n_spl_,
    g1687_p_spl_
  );


  or

  (
    g1738_n,
    g1736_p_spl_,
    g1687_n_spl_
  );


  and

  (
    g1739_p,
    g1738_n,
    g1737_n_spl_
  );


  or

  (
    g1739_n,
    g1738_p,
    g1737_p_spl_
  );


  and

  (
    g1740_p,
    g1739_p,
    g1686_n
  );


  or

  (
    g1740_n,
    g1739_n_spl_,
    g1686_p_spl_
  );


  and

  (
    g1741_p,
    g1739_n_spl_,
    g1686_p_spl_
  );


  or

  (
    g1742_n,
    g1741_p,
    g1740_p_spl_
  );


  and

  (
    g1743_p,
    g1740_n,
    g1737_n_spl_
  );


  or

  (
    g1743_n,
    g1740_p_spl_,
    g1737_p_spl_
  );


  and

  (
    g1744_p,
    g1734_n_spl_,
    g1731_n_spl_
  );


  or

  (
    g1744_n,
    g1734_p_spl_,
    g1731_p_spl_
  );


  and

  (
    g1745_p,
    G32_p_spl_101,
    G11_p_spl_111
  );


  or

  (
    g1745_n,
    G32_n_spl_101,
    G11_n_spl_111
  );


  and

  (
    g1746_p,
    g1728_n_spl_,
    g1725_n_spl_
  );


  or

  (
    g1746_n,
    g1728_p_spl_,
    g1725_p_spl_
  );


  and

  (
    g1747_p,
    G31_p_spl_101,
    G12_p_spl_111
  );


  or

  (
    g1747_n,
    G31_n_spl_101,
    G12_n_spl_111
  );


  and

  (
    g1748_p,
    g1722_n_spl_,
    g1719_n_spl_
  );


  or

  (
    g1748_n,
    g1722_p_spl_,
    g1719_p_spl_
  );


  and

  (
    g1749_p,
    G30_p_spl_110,
    G13_p_spl_110
  );


  or

  (
    g1749_n,
    G30_n_spl_110,
    G13_n_spl_110
  );


  and

  (
    g1750_p,
    g1716_n_spl_,
    g1713_n_spl_
  );


  or

  (
    g1750_n,
    g1716_p_spl_,
    g1713_p_spl_
  );


  and

  (
    g1751_p,
    G29_p_spl_110,
    G14_p_spl_110
  );


  or

  (
    g1751_n,
    G29_n_spl_110,
    G14_n_spl_110
  );


  and

  (
    g1752_p,
    g1710_n_spl_,
    g1707_n_spl_
  );


  or

  (
    g1752_n,
    g1710_p_spl_,
    g1707_p_spl_
  );


  and

  (
    g1753_p,
    G28_p_spl_111,
    G15_p_spl_101
  );


  or

  (
    g1753_n,
    G28_n_spl_111,
    G15_n_spl_101
  );


  and

  (
    g1754_p,
    G27_p_spl_111,
    G16_p_spl_101
  );


  or

  (
    g1754_n,
    G27_n_spl_111,
    G16_n_spl_101
  );


  and

  (
    g1755_p,
    g1704_n_spl_,
    g1701_n_spl_
  );


  or

  (
    g1755_n,
    g1704_p_spl_,
    g1701_p_spl_
  );


  and

  (
    g1756_p,
    g1755_n_spl_,
    g1754_n_spl_
  );


  or

  (
    g1756_n,
    g1755_p_spl_,
    g1754_p_spl_
  );


  and

  (
    g1757_p,
    g1755_p_spl_,
    g1754_p_spl_
  );


  or

  (
    g1757_n,
    g1755_n_spl_,
    g1754_n_spl_
  );


  and

  (
    g1758_p,
    g1757_n,
    g1756_n_spl_
  );


  or

  (
    g1758_n,
    g1757_p,
    g1756_p_spl_
  );


  and

  (
    g1759_p,
    g1758_p_spl_,
    g1753_n_spl_
  );


  or

  (
    g1759_n,
    g1758_n_spl_,
    g1753_p_spl_
  );


  and

  (
    g1760_p,
    g1758_n_spl_,
    g1753_p_spl_
  );


  or

  (
    g1760_n,
    g1758_p_spl_,
    g1753_n_spl_
  );


  and

  (
    g1761_p,
    g1760_n,
    g1759_n_spl_
  );


  or

  (
    g1761_n,
    g1760_p,
    g1759_p_spl_
  );


  and

  (
    g1762_p,
    g1761_p_spl_,
    g1752_n_spl_
  );


  or

  (
    g1762_n,
    g1761_n_spl_,
    g1752_p_spl_
  );


  and

  (
    g1763_p,
    g1761_n_spl_,
    g1752_p_spl_
  );


  or

  (
    g1763_n,
    g1761_p_spl_,
    g1752_n_spl_
  );


  and

  (
    g1764_p,
    g1763_n,
    g1762_n_spl_
  );


  or

  (
    g1764_n,
    g1763_p,
    g1762_p_spl_
  );


  and

  (
    g1765_p,
    g1764_p_spl_,
    g1751_n_spl_
  );


  or

  (
    g1765_n,
    g1764_n_spl_,
    g1751_p_spl_
  );


  and

  (
    g1766_p,
    g1764_n_spl_,
    g1751_p_spl_
  );


  or

  (
    g1766_n,
    g1764_p_spl_,
    g1751_n_spl_
  );


  and

  (
    g1767_p,
    g1766_n,
    g1765_n_spl_
  );


  or

  (
    g1767_n,
    g1766_p,
    g1765_p_spl_
  );


  and

  (
    g1768_p,
    g1767_p_spl_,
    g1750_n_spl_
  );


  or

  (
    g1768_n,
    g1767_n_spl_,
    g1750_p_spl_
  );


  and

  (
    g1769_p,
    g1767_n_spl_,
    g1750_p_spl_
  );


  or

  (
    g1769_n,
    g1767_p_spl_,
    g1750_n_spl_
  );


  and

  (
    g1770_p,
    g1769_n,
    g1768_n_spl_
  );


  or

  (
    g1770_n,
    g1769_p,
    g1768_p_spl_
  );


  and

  (
    g1771_p,
    g1770_p_spl_,
    g1749_n_spl_
  );


  or

  (
    g1771_n,
    g1770_n_spl_,
    g1749_p_spl_
  );


  and

  (
    g1772_p,
    g1770_n_spl_,
    g1749_p_spl_
  );


  or

  (
    g1772_n,
    g1770_p_spl_,
    g1749_n_spl_
  );


  and

  (
    g1773_p,
    g1772_n,
    g1771_n_spl_
  );


  or

  (
    g1773_n,
    g1772_p,
    g1771_p_spl_
  );


  and

  (
    g1774_p,
    g1773_p_spl_,
    g1748_n_spl_
  );


  or

  (
    g1774_n,
    g1773_n_spl_,
    g1748_p_spl_
  );


  and

  (
    g1775_p,
    g1773_n_spl_,
    g1748_p_spl_
  );


  or

  (
    g1775_n,
    g1773_p_spl_,
    g1748_n_spl_
  );


  and

  (
    g1776_p,
    g1775_n,
    g1774_n_spl_
  );


  or

  (
    g1776_n,
    g1775_p,
    g1774_p_spl_
  );


  and

  (
    g1777_p,
    g1776_p_spl_,
    g1747_n_spl_
  );


  or

  (
    g1777_n,
    g1776_n_spl_,
    g1747_p_spl_
  );


  and

  (
    g1778_p,
    g1776_n_spl_,
    g1747_p_spl_
  );


  or

  (
    g1778_n,
    g1776_p_spl_,
    g1747_n_spl_
  );


  and

  (
    g1779_p,
    g1778_n,
    g1777_n_spl_
  );


  or

  (
    g1779_n,
    g1778_p,
    g1777_p_spl_
  );


  and

  (
    g1780_p,
    g1779_p_spl_,
    g1746_n_spl_
  );


  or

  (
    g1780_n,
    g1779_n_spl_,
    g1746_p_spl_
  );


  and

  (
    g1781_p,
    g1779_n_spl_,
    g1746_p_spl_
  );


  or

  (
    g1781_n,
    g1779_p_spl_,
    g1746_n_spl_
  );


  and

  (
    g1782_p,
    g1781_n,
    g1780_n_spl_
  );


  or

  (
    g1782_n,
    g1781_p,
    g1780_p_spl_
  );


  and

  (
    g1783_p,
    g1782_p_spl_,
    g1745_n_spl_
  );


  or

  (
    g1783_n,
    g1782_n_spl_,
    g1745_p_spl_
  );


  and

  (
    g1784_p,
    g1782_n_spl_,
    g1745_p_spl_
  );


  or

  (
    g1784_n,
    g1782_p_spl_,
    g1745_n_spl_
  );


  and

  (
    g1785_p,
    g1784_n,
    g1783_n_spl_
  );


  or

  (
    g1785_n,
    g1784_p,
    g1783_p_spl_
  );


  and

  (
    g1786_p,
    g1785_p_spl_,
    g1744_n_spl_
  );


  or

  (
    g1786_n,
    g1785_n_spl_,
    g1744_p_spl_
  );


  and

  (
    g1787_p,
    g1785_n_spl_,
    g1744_p_spl_
  );


  or

  (
    g1787_n,
    g1785_p_spl_,
    g1744_n_spl_
  );


  and

  (
    g1788_p,
    g1787_n,
    g1786_n_spl_
  );


  or

  (
    g1788_n,
    g1787_p,
    g1786_p_spl_
  );


  and

  (
    g1789_p,
    g1788_p,
    g1743_n
  );


  or

  (
    g1789_n,
    g1788_n_spl_,
    g1743_p_spl_
  );


  and

  (
    g1790_p,
    g1788_n_spl_,
    g1743_p_spl_
  );


  or

  (
    g1791_n,
    g1790_p,
    g1789_p_spl_
  );


  and

  (
    g1792_p,
    g1789_n,
    g1786_n_spl_
  );


  or

  (
    g1792_n,
    g1789_p_spl_,
    g1786_p_spl_
  );


  and

  (
    g1793_p,
    g1783_n_spl_,
    g1780_n_spl_
  );


  or

  (
    g1793_n,
    g1783_p_spl_,
    g1780_p_spl_
  );


  and

  (
    g1794_p,
    G32_p_spl_101,
    G12_p_spl_111
  );


  or

  (
    g1794_n,
    G32_n_spl_101,
    G12_n_spl_111
  );


  and

  (
    g1795_p,
    g1777_n_spl_,
    g1774_n_spl_
  );


  or

  (
    g1795_n,
    g1777_p_spl_,
    g1774_p_spl_
  );


  and

  (
    g1796_p,
    G31_p_spl_110,
    G13_p_spl_111
  );


  or

  (
    g1796_n,
    G31_n_spl_110,
    G13_n_spl_111
  );


  and

  (
    g1797_p,
    g1771_n_spl_,
    g1768_n_spl_
  );


  or

  (
    g1797_n,
    g1771_p_spl_,
    g1768_p_spl_
  );


  and

  (
    g1798_p,
    G30_p_spl_110,
    G14_p_spl_110
  );


  or

  (
    g1798_n,
    G30_n_spl_110,
    G14_n_spl_110
  );


  and

  (
    g1799_p,
    g1765_n_spl_,
    g1762_n_spl_
  );


  or

  (
    g1799_n,
    g1765_p_spl_,
    g1762_p_spl_
  );


  and

  (
    g1800_p,
    G29_p_spl_111,
    G15_p_spl_110
  );


  or

  (
    g1800_n,
    G29_n_spl_111,
    G15_n_spl_110
  );


  and

  (
    g1801_p,
    G28_p_spl_111,
    G16_p_spl_101
  );


  or

  (
    g1801_n,
    G28_n_spl_111,
    G16_n_spl_101
  );


  and

  (
    g1802_p,
    g1759_n_spl_,
    g1756_n_spl_
  );


  or

  (
    g1802_n,
    g1759_p_spl_,
    g1756_p_spl_
  );


  and

  (
    g1803_p,
    g1802_n_spl_,
    g1801_n_spl_
  );


  or

  (
    g1803_n,
    g1802_p_spl_,
    g1801_p_spl_
  );


  and

  (
    g1804_p,
    g1802_p_spl_,
    g1801_p_spl_
  );


  or

  (
    g1804_n,
    g1802_n_spl_,
    g1801_n_spl_
  );


  and

  (
    g1805_p,
    g1804_n,
    g1803_n_spl_
  );


  or

  (
    g1805_n,
    g1804_p,
    g1803_p_spl_
  );


  and

  (
    g1806_p,
    g1805_p_spl_,
    g1800_n_spl_
  );


  or

  (
    g1806_n,
    g1805_n_spl_,
    g1800_p_spl_
  );


  and

  (
    g1807_p,
    g1805_n_spl_,
    g1800_p_spl_
  );


  or

  (
    g1807_n,
    g1805_p_spl_,
    g1800_n_spl_
  );


  and

  (
    g1808_p,
    g1807_n,
    g1806_n_spl_
  );


  or

  (
    g1808_n,
    g1807_p,
    g1806_p_spl_
  );


  and

  (
    g1809_p,
    g1808_p_spl_,
    g1799_n_spl_
  );


  or

  (
    g1809_n,
    g1808_n_spl_,
    g1799_p_spl_
  );


  and

  (
    g1810_p,
    g1808_n_spl_,
    g1799_p_spl_
  );


  or

  (
    g1810_n,
    g1808_p_spl_,
    g1799_n_spl_
  );


  and

  (
    g1811_p,
    g1810_n,
    g1809_n_spl_
  );


  or

  (
    g1811_n,
    g1810_p,
    g1809_p_spl_
  );


  and

  (
    g1812_p,
    g1811_p_spl_,
    g1798_n_spl_
  );


  or

  (
    g1812_n,
    g1811_n_spl_,
    g1798_p_spl_
  );


  and

  (
    g1813_p,
    g1811_n_spl_,
    g1798_p_spl_
  );


  or

  (
    g1813_n,
    g1811_p_spl_,
    g1798_n_spl_
  );


  and

  (
    g1814_p,
    g1813_n,
    g1812_n_spl_
  );


  or

  (
    g1814_n,
    g1813_p,
    g1812_p_spl_
  );


  and

  (
    g1815_p,
    g1814_p_spl_,
    g1797_n_spl_
  );


  or

  (
    g1815_n,
    g1814_n_spl_,
    g1797_p_spl_
  );


  and

  (
    g1816_p,
    g1814_n_spl_,
    g1797_p_spl_
  );


  or

  (
    g1816_n,
    g1814_p_spl_,
    g1797_n_spl_
  );


  and

  (
    g1817_p,
    g1816_n,
    g1815_n_spl_
  );


  or

  (
    g1817_n,
    g1816_p,
    g1815_p_spl_
  );


  and

  (
    g1818_p,
    g1817_p_spl_,
    g1796_n_spl_
  );


  or

  (
    g1818_n,
    g1817_n_spl_,
    g1796_p_spl_
  );


  and

  (
    g1819_p,
    g1817_n_spl_,
    g1796_p_spl_
  );


  or

  (
    g1819_n,
    g1817_p_spl_,
    g1796_n_spl_
  );


  and

  (
    g1820_p,
    g1819_n,
    g1818_n_spl_
  );


  or

  (
    g1820_n,
    g1819_p,
    g1818_p_spl_
  );


  and

  (
    g1821_p,
    g1820_p_spl_,
    g1795_n_spl_
  );


  or

  (
    g1821_n,
    g1820_n_spl_,
    g1795_p_spl_
  );


  and

  (
    g1822_p,
    g1820_n_spl_,
    g1795_p_spl_
  );


  or

  (
    g1822_n,
    g1820_p_spl_,
    g1795_n_spl_
  );


  and

  (
    g1823_p,
    g1822_n,
    g1821_n_spl_
  );


  or

  (
    g1823_n,
    g1822_p,
    g1821_p_spl_
  );


  and

  (
    g1824_p,
    g1823_p_spl_,
    g1794_n_spl_
  );


  or

  (
    g1824_n,
    g1823_n_spl_,
    g1794_p_spl_
  );


  and

  (
    g1825_p,
    g1823_n_spl_,
    g1794_p_spl_
  );


  or

  (
    g1825_n,
    g1823_p_spl_,
    g1794_n_spl_
  );


  and

  (
    g1826_p,
    g1825_n,
    g1824_n_spl_
  );


  or

  (
    g1826_n,
    g1825_p,
    g1824_p_spl_
  );


  and

  (
    g1827_p,
    g1826_p_spl_,
    g1793_n_spl_
  );


  or

  (
    g1827_n,
    g1826_n_spl_,
    g1793_p_spl_
  );


  and

  (
    g1828_p,
    g1826_n_spl_,
    g1793_p_spl_
  );


  or

  (
    g1828_n,
    g1826_p_spl_,
    g1793_n_spl_
  );


  and

  (
    g1829_p,
    g1828_n,
    g1827_n_spl_
  );


  or

  (
    g1829_n,
    g1828_p,
    g1827_p_spl_
  );


  and

  (
    g1830_p,
    g1829_p,
    g1792_n
  );


  or

  (
    g1830_n,
    g1829_n_spl_,
    g1792_p_spl_
  );


  and

  (
    g1831_p,
    g1829_n_spl_,
    g1792_p_spl_
  );


  or

  (
    g1832_n,
    g1831_p,
    g1830_p_spl_
  );


  and

  (
    g1833_p,
    g1830_n,
    g1827_n_spl_
  );


  or

  (
    g1833_n,
    g1830_p_spl_,
    g1827_p_spl_
  );


  and

  (
    g1834_p,
    g1824_n_spl_,
    g1821_n_spl_
  );


  or

  (
    g1834_n,
    g1824_p_spl_,
    g1821_p_spl_
  );


  and

  (
    g1835_p,
    G32_p_spl_110,
    G13_p_spl_111
  );


  or

  (
    g1835_n,
    G32_n_spl_110,
    G13_n_spl_111
  );


  and

  (
    g1836_p,
    g1818_n_spl_,
    g1815_n_spl_
  );


  or

  (
    g1836_n,
    g1818_p_spl_,
    g1815_p_spl_
  );


  and

  (
    g1837_p,
    G31_p_spl_110,
    G14_p_spl_111
  );


  or

  (
    g1837_n,
    G31_n_spl_110,
    G14_n_spl_111
  );


  and

  (
    g1838_p,
    g1812_n_spl_,
    g1809_n_spl_
  );


  or

  (
    g1838_n,
    g1812_p_spl_,
    g1809_p_spl_
  );


  and

  (
    g1839_p,
    G30_p_spl_111,
    G15_p_spl_110
  );


  or

  (
    g1839_n,
    G30_n_spl_111,
    G15_n_spl_110
  );


  and

  (
    g1840_p,
    G29_p_spl_111,
    G16_p_spl_110
  );


  or

  (
    g1840_n,
    G29_n_spl_111,
    G16_n_spl_110
  );


  and

  (
    g1841_p,
    g1806_n_spl_,
    g1803_n_spl_
  );


  or

  (
    g1841_n,
    g1806_p_spl_,
    g1803_p_spl_
  );


  and

  (
    g1842_p,
    g1841_n_spl_,
    g1840_n_spl_
  );


  or

  (
    g1842_n,
    g1841_p_spl_,
    g1840_p_spl_
  );


  and

  (
    g1843_p,
    g1841_p_spl_,
    g1840_p_spl_
  );


  or

  (
    g1843_n,
    g1841_n_spl_,
    g1840_n_spl_
  );


  and

  (
    g1844_p,
    g1843_n,
    g1842_n_spl_
  );


  or

  (
    g1844_n,
    g1843_p,
    g1842_p_spl_
  );


  and

  (
    g1845_p,
    g1844_p_spl_,
    g1839_n_spl_
  );


  or

  (
    g1845_n,
    g1844_n_spl_,
    g1839_p_spl_
  );


  and

  (
    g1846_p,
    g1844_n_spl_,
    g1839_p_spl_
  );


  or

  (
    g1846_n,
    g1844_p_spl_,
    g1839_n_spl_
  );


  and

  (
    g1847_p,
    g1846_n,
    g1845_n_spl_
  );


  or

  (
    g1847_n,
    g1846_p,
    g1845_p_spl_
  );


  and

  (
    g1848_p,
    g1847_p_spl_,
    g1838_n_spl_
  );


  or

  (
    g1848_n,
    g1847_n_spl_,
    g1838_p_spl_
  );


  and

  (
    g1849_p,
    g1847_n_spl_,
    g1838_p_spl_
  );


  or

  (
    g1849_n,
    g1847_p_spl_,
    g1838_n_spl_
  );


  and

  (
    g1850_p,
    g1849_n,
    g1848_n_spl_
  );


  or

  (
    g1850_n,
    g1849_p,
    g1848_p_spl_
  );


  and

  (
    g1851_p,
    g1850_p_spl_,
    g1837_n_spl_
  );


  or

  (
    g1851_n,
    g1850_n_spl_,
    g1837_p_spl_
  );


  and

  (
    g1852_p,
    g1850_n_spl_,
    g1837_p_spl_
  );


  or

  (
    g1852_n,
    g1850_p_spl_,
    g1837_n_spl_
  );


  and

  (
    g1853_p,
    g1852_n,
    g1851_n_spl_
  );


  or

  (
    g1853_n,
    g1852_p,
    g1851_p_spl_
  );


  and

  (
    g1854_p,
    g1853_p_spl_,
    g1836_n_spl_
  );


  or

  (
    g1854_n,
    g1853_n_spl_,
    g1836_p_spl_
  );


  and

  (
    g1855_p,
    g1853_n_spl_,
    g1836_p_spl_
  );


  or

  (
    g1855_n,
    g1853_p_spl_,
    g1836_n_spl_
  );


  and

  (
    g1856_p,
    g1855_n,
    g1854_n_spl_
  );


  or

  (
    g1856_n,
    g1855_p,
    g1854_p_spl_
  );


  and

  (
    g1857_p,
    g1856_p_spl_,
    g1835_n_spl_
  );


  or

  (
    g1857_n,
    g1856_n_spl_,
    g1835_p_spl_
  );


  and

  (
    g1858_p,
    g1856_n_spl_,
    g1835_p_spl_
  );


  or

  (
    g1858_n,
    g1856_p_spl_,
    g1835_n_spl_
  );


  and

  (
    g1859_p,
    g1858_n,
    g1857_n_spl_
  );


  or

  (
    g1859_n,
    g1858_p,
    g1857_p_spl_
  );


  and

  (
    g1860_p,
    g1859_p_spl_,
    g1834_n_spl_
  );


  or

  (
    g1860_n,
    g1859_n_spl_,
    g1834_p_spl_
  );


  and

  (
    g1861_p,
    g1859_n_spl_,
    g1834_p_spl_
  );


  or

  (
    g1861_n,
    g1859_p_spl_,
    g1834_n_spl_
  );


  and

  (
    g1862_p,
    g1861_n,
    g1860_n_spl_
  );


  or

  (
    g1862_n,
    g1861_p,
    g1860_p_spl_
  );


  and

  (
    g1863_p,
    g1862_p,
    g1833_n
  );


  or

  (
    g1863_n,
    g1862_n_spl_,
    g1833_p_spl_
  );


  and

  (
    g1864_p,
    g1862_n_spl_,
    g1833_p_spl_
  );


  or

  (
    g1865_n,
    g1864_p,
    g1863_p_spl_
  );


  and

  (
    g1866_p,
    g1863_n,
    g1860_n_spl_
  );


  or

  (
    g1866_n,
    g1863_p_spl_,
    g1860_p_spl_
  );


  and

  (
    g1867_p,
    g1857_n_spl_,
    g1854_n_spl_
  );


  or

  (
    g1867_n,
    g1857_p_spl_,
    g1854_p_spl_
  );


  and

  (
    g1868_p,
    G32_p_spl_110,
    G14_p_spl_111
  );


  or

  (
    g1868_n,
    G32_n_spl_110,
    G14_n_spl_111
  );


  and

  (
    g1869_p,
    g1851_n_spl_,
    g1848_n_spl_
  );


  or

  (
    g1869_n,
    g1851_p_spl_,
    g1848_p_spl_
  );


  and

  (
    g1870_p,
    G31_p_spl_111,
    G15_p_spl_111
  );


  or

  (
    g1870_n,
    G31_n_spl_111,
    G15_n_spl_111
  );


  and

  (
    g1871_p,
    G30_p_spl_111,
    G16_p_spl_110
  );


  or

  (
    g1871_n,
    G30_n_spl_111,
    G16_n_spl_110
  );


  and

  (
    g1872_p,
    g1845_n_spl_,
    g1842_n_spl_
  );


  or

  (
    g1872_n,
    g1845_p_spl_,
    g1842_p_spl_
  );


  and

  (
    g1873_p,
    g1872_n_spl_,
    g1871_n_spl_
  );


  or

  (
    g1873_n,
    g1872_p_spl_,
    g1871_p_spl_
  );


  and

  (
    g1874_p,
    g1872_p_spl_,
    g1871_p_spl_
  );


  or

  (
    g1874_n,
    g1872_n_spl_,
    g1871_n_spl_
  );


  and

  (
    g1875_p,
    g1874_n,
    g1873_n_spl_
  );


  or

  (
    g1875_n,
    g1874_p,
    g1873_p_spl_
  );


  and

  (
    g1876_p,
    g1875_p_spl_,
    g1870_n_spl_
  );


  or

  (
    g1876_n,
    g1875_n_spl_,
    g1870_p_spl_
  );


  and

  (
    g1877_p,
    g1875_n_spl_,
    g1870_p_spl_
  );


  or

  (
    g1877_n,
    g1875_p_spl_,
    g1870_n_spl_
  );


  and

  (
    g1878_p,
    g1877_n,
    g1876_n_spl_
  );


  or

  (
    g1878_n,
    g1877_p,
    g1876_p_spl_
  );


  and

  (
    g1879_p,
    g1878_p_spl_,
    g1869_n_spl_
  );


  or

  (
    g1879_n,
    g1878_n_spl_,
    g1869_p_spl_
  );


  and

  (
    g1880_p,
    g1878_n_spl_,
    g1869_p_spl_
  );


  or

  (
    g1880_n,
    g1878_p_spl_,
    g1869_n_spl_
  );


  and

  (
    g1881_p,
    g1880_n,
    g1879_n_spl_
  );


  or

  (
    g1881_n,
    g1880_p,
    g1879_p_spl_
  );


  and

  (
    g1882_p,
    g1881_p_spl_,
    g1868_n_spl_
  );


  or

  (
    g1882_n,
    g1881_n_spl_,
    g1868_p_spl_
  );


  and

  (
    g1883_p,
    g1881_n_spl_,
    g1868_p_spl_
  );


  or

  (
    g1883_n,
    g1881_p_spl_,
    g1868_n_spl_
  );


  and

  (
    g1884_p,
    g1883_n,
    g1882_n_spl_
  );


  or

  (
    g1884_n,
    g1883_p,
    g1882_p_spl_
  );


  and

  (
    g1885_p,
    g1884_p_spl_,
    g1867_n_spl_
  );


  or

  (
    g1885_n,
    g1884_n_spl_,
    g1867_p_spl_
  );


  and

  (
    g1886_p,
    g1884_n_spl_,
    g1867_p_spl_
  );


  or

  (
    g1886_n,
    g1884_p_spl_,
    g1867_n_spl_
  );


  and

  (
    g1887_p,
    g1886_n,
    g1885_n_spl_
  );


  or

  (
    g1887_n,
    g1886_p,
    g1885_p_spl_
  );


  and

  (
    g1888_p,
    g1887_p,
    g1866_n
  );


  or

  (
    g1888_n,
    g1887_n_spl_,
    g1866_p_spl_
  );


  and

  (
    g1889_p,
    g1887_n_spl_,
    g1866_p_spl_
  );


  or

  (
    g1890_n,
    g1889_p,
    g1888_p_spl_
  );


  and

  (
    g1891_p,
    g1888_n,
    g1885_n_spl_
  );


  or

  (
    g1891_n,
    g1888_p_spl_,
    g1885_p_spl_
  );


  and

  (
    g1892_p,
    g1882_n_spl_,
    g1879_n_spl_
  );


  or

  (
    g1892_n,
    g1882_p_spl_,
    g1879_p_spl_
  );


  and

  (
    g1893_p,
    G32_p_spl_111,
    G15_p_spl_111
  );


  or

  (
    g1893_n,
    G32_n_spl_111,
    G15_n_spl_111
  );


  and

  (
    g1894_p,
    G31_p_spl_111,
    G16_p_spl_111
  );


  or

  (
    g1894_n,
    G31_n_spl_111,
    G16_n_spl_111
  );


  and

  (
    g1895_p,
    g1876_n_spl_,
    g1873_n_spl_
  );


  or

  (
    g1895_n,
    g1876_p_spl_,
    g1873_p_spl_
  );


  and

  (
    g1896_p,
    g1895_n_spl_,
    g1894_n_spl_
  );


  or

  (
    g1896_n,
    g1895_p_spl_,
    g1894_p_spl_
  );


  and

  (
    g1897_p,
    g1895_p_spl_,
    g1894_p_spl_
  );


  or

  (
    g1897_n,
    g1895_n_spl_,
    g1894_n_spl_
  );


  and

  (
    g1898_p,
    g1897_n,
    g1896_n_spl_
  );


  or

  (
    g1898_n,
    g1897_p,
    g1896_p_spl_
  );


  and

  (
    g1899_p,
    g1898_p_spl_,
    g1893_n_spl_
  );


  or

  (
    g1899_n,
    g1898_n_spl_,
    g1893_p_spl_
  );


  and

  (
    g1900_p,
    g1898_n_spl_,
    g1893_p_spl_
  );


  or

  (
    g1900_n,
    g1898_p_spl_,
    g1893_n_spl_
  );


  and

  (
    g1901_p,
    g1900_n,
    g1899_n_spl_
  );


  or

  (
    g1901_n,
    g1900_p,
    g1899_p_spl_
  );


  and

  (
    g1902_p,
    g1901_p_spl_,
    g1892_n_spl_
  );


  or

  (
    g1902_n,
    g1901_n_spl_,
    g1892_p_spl_
  );


  and

  (
    g1903_p,
    g1901_n_spl_,
    g1892_p_spl_
  );


  or

  (
    g1903_n,
    g1901_p_spl_,
    g1892_n_spl_
  );


  and

  (
    g1904_p,
    g1903_n,
    g1902_n_spl_
  );


  or

  (
    g1904_n,
    g1903_p,
    g1902_p_spl_
  );


  and

  (
    g1905_p,
    g1904_p,
    g1891_n
  );


  or

  (
    g1905_n,
    g1904_n_spl_,
    g1891_p_spl_
  );


  and

  (
    g1906_p,
    g1904_n_spl_,
    g1891_p_spl_
  );


  or

  (
    g1907_n,
    g1906_p,
    g1905_p_spl_
  );


  and

  (
    g1908_p,
    G32_p_spl_111,
    G16_p_spl_111
  );


  or

  (
    g1908_n,
    G32_n_spl_111,
    G16_n_spl_111
  );


  and

  (
    g1909_p,
    g1899_n_spl_,
    g1896_n_spl_
  );


  or

  (
    g1909_n,
    g1899_p_spl_,
    g1896_p_spl_
  );


  and

  (
    g1910_p,
    g1909_n_spl_,
    g1908_n_spl_
  );


  or

  (
    g1910_n,
    g1909_p_spl_,
    g1908_p_spl_
  );


  and

  (
    g1911_p,
    g1905_n,
    g1902_n_spl_
  );


  or

  (
    g1911_n,
    g1905_p_spl_,
    g1902_p_spl_
  );


  and

  (
    g1912_p,
    g1909_p_spl_,
    g1908_p_spl_
  );


  or

  (
    g1912_n,
    g1909_n_spl_,
    g1908_n_spl_
  );


  and

  (
    g1913_p,
    g1912_n,
    g1910_n_spl_
  );


  or

  (
    g1913_n,
    g1912_p,
    g1910_p
  );


  or

  (
    g1914_n,
    g1913_n,
    g1911_p
  );


  and

  (
    g1915_p,
    g1914_n_spl_,
    g1910_n_spl_
  );


  or

  (
    g1916_n,
    g1913_p,
    g1911_n
  );


  and

  (
    g1917_p,
    g1916_n,
    g1914_n_spl_
  );


  buf

  (
    G6257,
    g33_p
  );


  buf

  (
    G6258,
    g39_p
  );


  buf

  (
    G6259,
    g52_n
  );


  buf

  (
    G6260,
    g73_n
  );


  buf

  (
    G6261,
    g102_n
  );


  buf

  (
    G6262,
    g139_n
  );


  buf

  (
    G6263,
    g184_n
  );


  buf

  (
    G6264,
    g237_n
  );


  buf

  (
    G6265,
    g298_n
  );


  buf

  (
    G6266,
    g367_n
  );


  buf

  (
    G6267,
    g444_n
  );


  buf

  (
    G6268,
    g529_n
  );


  buf

  (
    G6269,
    g622_n
  );


  buf

  (
    G6270,
    g723_n
  );


  buf

  (
    G6271,
    g832_n
  );


  buf

  (
    G6272,
    g949_n
  );


  buf

  (
    G6273,
    g1063_p
  );


  buf

  (
    G6274,
    g1175_n
  );


  buf

  (
    G6275,
    g1280_n
  );


  buf

  (
    G6276,
    g1377_n
  );


  buf

  (
    G6277,
    g1466_n
  );


  buf

  (
    G6278,
    g1547_n
  );


  buf

  (
    G6279,
    g1620_n
  );


  buf

  (
    G6280,
    g1685_n
  );


  buf

  (
    G6281,
    g1742_n
  );


  buf

  (
    G6282,
    g1791_n
  );


  buf

  (
    G6283,
    g1832_n
  );


  buf

  (
    G6284,
    g1865_n
  );


  buf

  (
    G6285,
    g1890_n
  );


  buf

  (
    G6286,
    g1907_n
  );


  buf

  (
    G6287,
    g1915_p
  );


  not

  (
    G6288,
    g1917_p
  );


  buf

  (
    G17_p_spl_,
    G17_p
  );


  buf

  (
    G17_p_spl_0,
    G17_p_spl_
  );


  buf

  (
    G17_p_spl_00,
    G17_p_spl_0
  );


  buf

  (
    G17_p_spl_000,
    G17_p_spl_00
  );


  buf

  (
    G17_p_spl_001,
    G17_p_spl_00
  );


  buf

  (
    G17_p_spl_01,
    G17_p_spl_0
  );


  buf

  (
    G17_p_spl_010,
    G17_p_spl_01
  );


  buf

  (
    G17_p_spl_011,
    G17_p_spl_01
  );


  buf

  (
    G17_p_spl_1,
    G17_p_spl_
  );


  buf

  (
    G17_p_spl_10,
    G17_p_spl_1
  );


  buf

  (
    G17_p_spl_100,
    G17_p_spl_10
  );


  buf

  (
    G17_p_spl_101,
    G17_p_spl_10
  );


  buf

  (
    G17_p_spl_11,
    G17_p_spl_1
  );


  buf

  (
    G17_p_spl_110,
    G17_p_spl_11
  );


  buf

  (
    G17_p_spl_111,
    G17_p_spl_11
  );


  buf

  (
    G1_p_spl_,
    G1_p
  );


  buf

  (
    G1_p_spl_0,
    G1_p_spl_
  );


  buf

  (
    G1_p_spl_00,
    G1_p_spl_0
  );


  buf

  (
    G1_p_spl_000,
    G1_p_spl_00
  );


  buf

  (
    G1_p_spl_001,
    G1_p_spl_00
  );


  buf

  (
    G1_p_spl_01,
    G1_p_spl_0
  );


  buf

  (
    G1_p_spl_010,
    G1_p_spl_01
  );


  buf

  (
    G1_p_spl_011,
    G1_p_spl_01
  );


  buf

  (
    G1_p_spl_1,
    G1_p_spl_
  );


  buf

  (
    G1_p_spl_10,
    G1_p_spl_1
  );


  buf

  (
    G1_p_spl_100,
    G1_p_spl_10
  );


  buf

  (
    G1_p_spl_101,
    G1_p_spl_10
  );


  buf

  (
    G1_p_spl_11,
    G1_p_spl_1
  );


  buf

  (
    G1_p_spl_110,
    G1_p_spl_11
  );


  buf

  (
    G1_p_spl_111,
    G1_p_spl_11
  );


  buf

  (
    G2_p_spl_,
    G2_p
  );


  buf

  (
    G2_p_spl_0,
    G2_p_spl_
  );


  buf

  (
    G2_p_spl_00,
    G2_p_spl_0
  );


  buf

  (
    G2_p_spl_000,
    G2_p_spl_00
  );


  buf

  (
    G2_p_spl_001,
    G2_p_spl_00
  );


  buf

  (
    G2_p_spl_01,
    G2_p_spl_0
  );


  buf

  (
    G2_p_spl_010,
    G2_p_spl_01
  );


  buf

  (
    G2_p_spl_011,
    G2_p_spl_01
  );


  buf

  (
    G2_p_spl_1,
    G2_p_spl_
  );


  buf

  (
    G2_p_spl_10,
    G2_p_spl_1
  );


  buf

  (
    G2_p_spl_100,
    G2_p_spl_10
  );


  buf

  (
    G2_p_spl_101,
    G2_p_spl_10
  );


  buf

  (
    G2_p_spl_11,
    G2_p_spl_1
  );


  buf

  (
    G2_p_spl_110,
    G2_p_spl_11
  );


  buf

  (
    G2_p_spl_111,
    G2_p_spl_11
  );


  buf

  (
    G17_n_spl_,
    G17_n
  );


  buf

  (
    G17_n_spl_0,
    G17_n_spl_
  );


  buf

  (
    G17_n_spl_00,
    G17_n_spl_0
  );


  buf

  (
    G17_n_spl_000,
    G17_n_spl_00
  );


  buf

  (
    G17_n_spl_001,
    G17_n_spl_00
  );


  buf

  (
    G17_n_spl_01,
    G17_n_spl_0
  );


  buf

  (
    G17_n_spl_010,
    G17_n_spl_01
  );


  buf

  (
    G17_n_spl_011,
    G17_n_spl_01
  );


  buf

  (
    G17_n_spl_1,
    G17_n_spl_
  );


  buf

  (
    G17_n_spl_10,
    G17_n_spl_1
  );


  buf

  (
    G17_n_spl_100,
    G17_n_spl_10
  );


  buf

  (
    G17_n_spl_101,
    G17_n_spl_10
  );


  buf

  (
    G17_n_spl_11,
    G17_n_spl_1
  );


  buf

  (
    G17_n_spl_110,
    G17_n_spl_11
  );


  buf

  (
    G2_n_spl_,
    G2_n
  );


  buf

  (
    G2_n_spl_0,
    G2_n_spl_
  );


  buf

  (
    G2_n_spl_00,
    G2_n_spl_0
  );


  buf

  (
    G2_n_spl_000,
    G2_n_spl_00
  );


  buf

  (
    G2_n_spl_001,
    G2_n_spl_00
  );


  buf

  (
    G2_n_spl_01,
    G2_n_spl_0
  );


  buf

  (
    G2_n_spl_010,
    G2_n_spl_01
  );


  buf

  (
    G2_n_spl_011,
    G2_n_spl_01
  );


  buf

  (
    G2_n_spl_1,
    G2_n_spl_
  );


  buf

  (
    G2_n_spl_10,
    G2_n_spl_1
  );


  buf

  (
    G2_n_spl_100,
    G2_n_spl_10
  );


  buf

  (
    G2_n_spl_101,
    G2_n_spl_10
  );


  buf

  (
    G2_n_spl_11,
    G2_n_spl_1
  );


  buf

  (
    G2_n_spl_110,
    G2_n_spl_11
  );


  buf

  (
    G2_n_spl_111,
    G2_n_spl_11
  );


  buf

  (
    G18_p_spl_,
    G18_p
  );


  buf

  (
    G18_p_spl_0,
    G18_p_spl_
  );


  buf

  (
    G18_p_spl_00,
    G18_p_spl_0
  );


  buf

  (
    G18_p_spl_000,
    G18_p_spl_00
  );


  buf

  (
    G18_p_spl_001,
    G18_p_spl_00
  );


  buf

  (
    G18_p_spl_01,
    G18_p_spl_0
  );


  buf

  (
    G18_p_spl_010,
    G18_p_spl_01
  );


  buf

  (
    G18_p_spl_011,
    G18_p_spl_01
  );


  buf

  (
    G18_p_spl_1,
    G18_p_spl_
  );


  buf

  (
    G18_p_spl_10,
    G18_p_spl_1
  );


  buf

  (
    G18_p_spl_100,
    G18_p_spl_10
  );


  buf

  (
    G18_p_spl_101,
    G18_p_spl_10
  );


  buf

  (
    G18_p_spl_11,
    G18_p_spl_1
  );


  buf

  (
    G18_p_spl_110,
    G18_p_spl_11
  );


  buf

  (
    G18_p_spl_111,
    G18_p_spl_11
  );


  buf

  (
    G18_n_spl_,
    G18_n
  );


  buf

  (
    G18_n_spl_0,
    G18_n_spl_
  );


  buf

  (
    G18_n_spl_00,
    G18_n_spl_0
  );


  buf

  (
    G18_n_spl_000,
    G18_n_spl_00
  );


  buf

  (
    G18_n_spl_001,
    G18_n_spl_00
  );


  buf

  (
    G18_n_spl_01,
    G18_n_spl_0
  );


  buf

  (
    G18_n_spl_010,
    G18_n_spl_01
  );


  buf

  (
    G18_n_spl_011,
    G18_n_spl_01
  );


  buf

  (
    G18_n_spl_1,
    G18_n_spl_
  );


  buf

  (
    G18_n_spl_10,
    G18_n_spl_1
  );


  buf

  (
    G18_n_spl_100,
    G18_n_spl_10
  );


  buf

  (
    G18_n_spl_101,
    G18_n_spl_10
  );


  buf

  (
    G18_n_spl_11,
    G18_n_spl_1
  );


  buf

  (
    G18_n_spl_110,
    G18_n_spl_11
  );


  buf

  (
    G18_n_spl_111,
    G18_n_spl_11
  );


  buf

  (
    G1_n_spl_,
    G1_n
  );


  buf

  (
    G1_n_spl_0,
    G1_n_spl_
  );


  buf

  (
    G1_n_spl_00,
    G1_n_spl_0
  );


  buf

  (
    G1_n_spl_000,
    G1_n_spl_00
  );


  buf

  (
    G1_n_spl_001,
    G1_n_spl_00
  );


  buf

  (
    G1_n_spl_01,
    G1_n_spl_0
  );


  buf

  (
    G1_n_spl_010,
    G1_n_spl_01
  );


  buf

  (
    G1_n_spl_011,
    G1_n_spl_01
  );


  buf

  (
    G1_n_spl_1,
    G1_n_spl_
  );


  buf

  (
    G1_n_spl_10,
    G1_n_spl_1
  );


  buf

  (
    G1_n_spl_100,
    G1_n_spl_10
  );


  buf

  (
    G1_n_spl_101,
    G1_n_spl_10
  );


  buf

  (
    G1_n_spl_11,
    G1_n_spl_1
  );


  buf

  (
    G1_n_spl_110,
    G1_n_spl_11
  );


  buf

  (
    g34_p_spl_,
    g34_p
  );


  buf

  (
    g35_p_spl_,
    g35_p
  );


  buf

  (
    g34_n_spl_,
    g34_n
  );


  buf

  (
    g36_p_spl_,
    g36_p
  );


  buf

  (
    g37_n_spl_,
    g37_n
  );


  buf

  (
    g37_n_spl_0,
    g37_n_spl_
  );


  buf

  (
    G19_p_spl_,
    G19_p
  );


  buf

  (
    G19_p_spl_0,
    G19_p_spl_
  );


  buf

  (
    G19_p_spl_00,
    G19_p_spl_0
  );


  buf

  (
    G19_p_spl_000,
    G19_p_spl_00
  );


  buf

  (
    G19_p_spl_001,
    G19_p_spl_00
  );


  buf

  (
    G19_p_spl_01,
    G19_p_spl_0
  );


  buf

  (
    G19_p_spl_010,
    G19_p_spl_01
  );


  buf

  (
    G19_p_spl_011,
    G19_p_spl_01
  );


  buf

  (
    G19_p_spl_1,
    G19_p_spl_
  );


  buf

  (
    G19_p_spl_10,
    G19_p_spl_1
  );


  buf

  (
    G19_p_spl_100,
    G19_p_spl_10
  );


  buf

  (
    G19_p_spl_101,
    G19_p_spl_10
  );


  buf

  (
    G19_p_spl_11,
    G19_p_spl_1
  );


  buf

  (
    G19_p_spl_110,
    G19_p_spl_11
  );


  buf

  (
    G19_p_spl_111,
    G19_p_spl_11
  );


  buf

  (
    G19_n_spl_,
    G19_n
  );


  buf

  (
    G19_n_spl_0,
    G19_n_spl_
  );


  buf

  (
    G19_n_spl_00,
    G19_n_spl_0
  );


  buf

  (
    G19_n_spl_000,
    G19_n_spl_00
  );


  buf

  (
    G19_n_spl_001,
    G19_n_spl_00
  );


  buf

  (
    G19_n_spl_01,
    G19_n_spl_0
  );


  buf

  (
    G19_n_spl_010,
    G19_n_spl_01
  );


  buf

  (
    G19_n_spl_011,
    G19_n_spl_01
  );


  buf

  (
    G19_n_spl_1,
    G19_n_spl_
  );


  buf

  (
    G19_n_spl_10,
    G19_n_spl_1
  );


  buf

  (
    G19_n_spl_100,
    G19_n_spl_10
  );


  buf

  (
    G19_n_spl_101,
    G19_n_spl_10
  );


  buf

  (
    G19_n_spl_11,
    G19_n_spl_1
  );


  buf

  (
    G19_n_spl_110,
    G19_n_spl_11
  );


  buf

  (
    G19_n_spl_111,
    G19_n_spl_11
  );


  buf

  (
    G3_p_spl_,
    G3_p
  );


  buf

  (
    G3_p_spl_0,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_00,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_000,
    G3_p_spl_00
  );


  buf

  (
    G3_p_spl_001,
    G3_p_spl_00
  );


  buf

  (
    G3_p_spl_01,
    G3_p_spl_0
  );


  buf

  (
    G3_p_spl_010,
    G3_p_spl_01
  );


  buf

  (
    G3_p_spl_011,
    G3_p_spl_01
  );


  buf

  (
    G3_p_spl_1,
    G3_p_spl_
  );


  buf

  (
    G3_p_spl_10,
    G3_p_spl_1
  );


  buf

  (
    G3_p_spl_100,
    G3_p_spl_10
  );


  buf

  (
    G3_p_spl_101,
    G3_p_spl_10
  );


  buf

  (
    G3_p_spl_11,
    G3_p_spl_1
  );


  buf

  (
    G3_p_spl_110,
    G3_p_spl_11
  );


  buf

  (
    G3_p_spl_111,
    G3_p_spl_11
  );


  buf

  (
    G3_n_spl_,
    G3_n
  );


  buf

  (
    G3_n_spl_0,
    G3_n_spl_
  );


  buf

  (
    G3_n_spl_00,
    G3_n_spl_0
  );


  buf

  (
    G3_n_spl_000,
    G3_n_spl_00
  );


  buf

  (
    G3_n_spl_001,
    G3_n_spl_00
  );


  buf

  (
    G3_n_spl_01,
    G3_n_spl_0
  );


  buf

  (
    G3_n_spl_010,
    G3_n_spl_01
  );


  buf

  (
    G3_n_spl_011,
    G3_n_spl_01
  );


  buf

  (
    G3_n_spl_1,
    G3_n_spl_
  );


  buf

  (
    G3_n_spl_10,
    G3_n_spl_1
  );


  buf

  (
    G3_n_spl_100,
    G3_n_spl_10
  );


  buf

  (
    G3_n_spl_101,
    G3_n_spl_10
  );


  buf

  (
    G3_n_spl_11,
    G3_n_spl_1
  );


  buf

  (
    G3_n_spl_110,
    G3_n_spl_11
  );


  buf

  (
    G3_n_spl_111,
    G3_n_spl_11
  );


  buf

  (
    g42_n_spl_,
    g42_n
  );


  buf

  (
    g41_p_spl_,
    g41_p
  );


  buf

  (
    g42_p_spl_,
    g42_p
  );


  buf

  (
    g41_n_spl_,
    g41_n
  );


  buf

  (
    g43_n_spl_,
    g43_n
  );


  buf

  (
    g43_p_spl_,
    g43_p
  );


  buf

  (
    g44_n_spl_,
    g44_n
  );


  buf

  (
    g44_n_spl_0,
    g44_n_spl_
  );


  buf

  (
    g44_p_spl_,
    g44_p
  );


  buf

  (
    g44_p_spl_0,
    g44_p_spl_
  );


  buf

  (
    g46_n_spl_,
    g46_n
  );


  buf

  (
    g46_p_spl_,
    g46_p
  );


  buf

  (
    g37_p_spl_,
    g37_p
  );


  buf

  (
    g47_n_spl_,
    g47_n
  );


  buf

  (
    g47_p_spl_,
    g47_p
  );


  buf

  (
    g49_n_spl_,
    g49_n
  );


  buf

  (
    g40_p_spl_,
    g40_p
  );


  buf

  (
    g50_p_spl_,
    g50_p
  );


  buf

  (
    G20_p_spl_,
    G20_p
  );


  buf

  (
    G20_p_spl_0,
    G20_p_spl_
  );


  buf

  (
    G20_p_spl_00,
    G20_p_spl_0
  );


  buf

  (
    G20_p_spl_000,
    G20_p_spl_00
  );


  buf

  (
    G20_p_spl_001,
    G20_p_spl_00
  );


  buf

  (
    G20_p_spl_01,
    G20_p_spl_0
  );


  buf

  (
    G20_p_spl_010,
    G20_p_spl_01
  );


  buf

  (
    G20_p_spl_011,
    G20_p_spl_01
  );


  buf

  (
    G20_p_spl_1,
    G20_p_spl_
  );


  buf

  (
    G20_p_spl_10,
    G20_p_spl_1
  );


  buf

  (
    G20_p_spl_100,
    G20_p_spl_10
  );


  buf

  (
    G20_p_spl_101,
    G20_p_spl_10
  );


  buf

  (
    G20_p_spl_11,
    G20_p_spl_1
  );


  buf

  (
    G20_p_spl_110,
    G20_p_spl_11
  );


  buf

  (
    G20_p_spl_111,
    G20_p_spl_11
  );


  buf

  (
    G20_n_spl_,
    G20_n
  );


  buf

  (
    G20_n_spl_0,
    G20_n_spl_
  );


  buf

  (
    G20_n_spl_00,
    G20_n_spl_0
  );


  buf

  (
    G20_n_spl_000,
    G20_n_spl_00
  );


  buf

  (
    G20_n_spl_001,
    G20_n_spl_00
  );


  buf

  (
    G20_n_spl_01,
    G20_n_spl_0
  );


  buf

  (
    G20_n_spl_010,
    G20_n_spl_01
  );


  buf

  (
    G20_n_spl_011,
    G20_n_spl_01
  );


  buf

  (
    G20_n_spl_1,
    G20_n_spl_
  );


  buf

  (
    G20_n_spl_10,
    G20_n_spl_1
  );


  buf

  (
    G20_n_spl_100,
    G20_n_spl_10
  );


  buf

  (
    G20_n_spl_101,
    G20_n_spl_10
  );


  buf

  (
    G20_n_spl_11,
    G20_n_spl_1
  );


  buf

  (
    G20_n_spl_110,
    G20_n_spl_11
  );


  buf

  (
    G20_n_spl_111,
    G20_n_spl_11
  );


  buf

  (
    G4_p_spl_,
    G4_p
  );


  buf

  (
    G4_p_spl_0,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_00,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_000,
    G4_p_spl_00
  );


  buf

  (
    G4_p_spl_001,
    G4_p_spl_00
  );


  buf

  (
    G4_p_spl_01,
    G4_p_spl_0
  );


  buf

  (
    G4_p_spl_010,
    G4_p_spl_01
  );


  buf

  (
    G4_p_spl_011,
    G4_p_spl_01
  );


  buf

  (
    G4_p_spl_1,
    G4_p_spl_
  );


  buf

  (
    G4_p_spl_10,
    G4_p_spl_1
  );


  buf

  (
    G4_p_spl_100,
    G4_p_spl_10
  );


  buf

  (
    G4_p_spl_101,
    G4_p_spl_10
  );


  buf

  (
    G4_p_spl_11,
    G4_p_spl_1
  );


  buf

  (
    G4_p_spl_110,
    G4_p_spl_11
  );


  buf

  (
    G4_p_spl_111,
    G4_p_spl_11
  );


  buf

  (
    G4_n_spl_,
    G4_n
  );


  buf

  (
    G4_n_spl_0,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_00,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_000,
    G4_n_spl_00
  );


  buf

  (
    G4_n_spl_001,
    G4_n_spl_00
  );


  buf

  (
    G4_n_spl_01,
    G4_n_spl_0
  );


  buf

  (
    G4_n_spl_010,
    G4_n_spl_01
  );


  buf

  (
    G4_n_spl_011,
    G4_n_spl_01
  );


  buf

  (
    G4_n_spl_1,
    G4_n_spl_
  );


  buf

  (
    G4_n_spl_10,
    G4_n_spl_1
  );


  buf

  (
    G4_n_spl_100,
    G4_n_spl_10
  );


  buf

  (
    G4_n_spl_101,
    G4_n_spl_10
  );


  buf

  (
    G4_n_spl_11,
    G4_n_spl_1
  );


  buf

  (
    G4_n_spl_110,
    G4_n_spl_11
  );


  buf

  (
    G4_n_spl_111,
    G4_n_spl_11
  );


  buf

  (
    g57_n_spl_,
    g57_n
  );


  buf

  (
    g56_p_spl_,
    g56_p
  );


  buf

  (
    g57_p_spl_,
    g57_p
  );


  buf

  (
    g56_n_spl_,
    g56_n
  );


  buf

  (
    g58_n_spl_,
    g58_n
  );


  buf

  (
    g58_p_spl_,
    g58_p
  );


  buf

  (
    g59_n_spl_,
    g59_n
  );


  buf

  (
    g59_n_spl_0,
    g59_n_spl_
  );


  buf

  (
    g59_p_spl_,
    g59_p
  );


  buf

  (
    g59_p_spl_0,
    g59_p_spl_
  );


  buf

  (
    g61_n_spl_,
    g61_n
  );


  buf

  (
    g61_p_spl_,
    g61_p
  );


  buf

  (
    g62_n_spl_,
    g62_n
  );


  buf

  (
    g62_p_spl_,
    g62_p
  );


  buf

  (
    g64_p_spl_,
    g64_p
  );


  buf

  (
    g55_n_spl_,
    g55_n
  );


  buf

  (
    g64_n_spl_,
    g64_n
  );


  buf

  (
    g55_p_spl_,
    g55_p
  );


  buf

  (
    g65_n_spl_,
    g65_n
  );


  buf

  (
    g65_p_spl_,
    g65_p
  );


  buf

  (
    g67_p_spl_,
    g67_p
  );


  buf

  (
    g54_n_spl_,
    g54_n
  );


  buf

  (
    g67_n_spl_,
    g67_n
  );


  buf

  (
    g54_p_spl_,
    g54_p
  );


  buf

  (
    g68_n_spl_,
    g68_n
  );


  buf

  (
    g68_p_spl_,
    g68_p
  );


  buf

  (
    g70_n_spl_,
    g70_n
  );


  buf

  (
    g53_p_spl_,
    g53_p
  );


  buf

  (
    g71_p_spl_,
    g71_p
  );


  buf

  (
    G21_p_spl_,
    G21_p
  );


  buf

  (
    G21_p_spl_0,
    G21_p_spl_
  );


  buf

  (
    G21_p_spl_00,
    G21_p_spl_0
  );


  buf

  (
    G21_p_spl_000,
    G21_p_spl_00
  );


  buf

  (
    G21_p_spl_001,
    G21_p_spl_00
  );


  buf

  (
    G21_p_spl_01,
    G21_p_spl_0
  );


  buf

  (
    G21_p_spl_010,
    G21_p_spl_01
  );


  buf

  (
    G21_p_spl_011,
    G21_p_spl_01
  );


  buf

  (
    G21_p_spl_1,
    G21_p_spl_
  );


  buf

  (
    G21_p_spl_10,
    G21_p_spl_1
  );


  buf

  (
    G21_p_spl_100,
    G21_p_spl_10
  );


  buf

  (
    G21_p_spl_101,
    G21_p_spl_10
  );


  buf

  (
    G21_p_spl_11,
    G21_p_spl_1
  );


  buf

  (
    G21_p_spl_110,
    G21_p_spl_11
  );


  buf

  (
    G21_p_spl_111,
    G21_p_spl_11
  );


  buf

  (
    G21_n_spl_,
    G21_n
  );


  buf

  (
    G21_n_spl_0,
    G21_n_spl_
  );


  buf

  (
    G21_n_spl_00,
    G21_n_spl_0
  );


  buf

  (
    G21_n_spl_000,
    G21_n_spl_00
  );


  buf

  (
    G21_n_spl_001,
    G21_n_spl_00
  );


  buf

  (
    G21_n_spl_01,
    G21_n_spl_0
  );


  buf

  (
    G21_n_spl_010,
    G21_n_spl_01
  );


  buf

  (
    G21_n_spl_011,
    G21_n_spl_01
  );


  buf

  (
    G21_n_spl_1,
    G21_n_spl_
  );


  buf

  (
    G21_n_spl_10,
    G21_n_spl_1
  );


  buf

  (
    G21_n_spl_100,
    G21_n_spl_10
  );


  buf

  (
    G21_n_spl_101,
    G21_n_spl_10
  );


  buf

  (
    G21_n_spl_11,
    G21_n_spl_1
  );


  buf

  (
    G21_n_spl_110,
    G21_n_spl_11
  );


  buf

  (
    G21_n_spl_111,
    G21_n_spl_11
  );


  buf

  (
    G5_p_spl_,
    G5_p
  );


  buf

  (
    G5_p_spl_0,
    G5_p_spl_
  );


  buf

  (
    G5_p_spl_00,
    G5_p_spl_0
  );


  buf

  (
    G5_p_spl_000,
    G5_p_spl_00
  );


  buf

  (
    G5_p_spl_001,
    G5_p_spl_00
  );


  buf

  (
    G5_p_spl_01,
    G5_p_spl_0
  );


  buf

  (
    G5_p_spl_010,
    G5_p_spl_01
  );


  buf

  (
    G5_p_spl_011,
    G5_p_spl_01
  );


  buf

  (
    G5_p_spl_1,
    G5_p_spl_
  );


  buf

  (
    G5_p_spl_10,
    G5_p_spl_1
  );


  buf

  (
    G5_p_spl_100,
    G5_p_spl_10
  );


  buf

  (
    G5_p_spl_101,
    G5_p_spl_10
  );


  buf

  (
    G5_p_spl_11,
    G5_p_spl_1
  );


  buf

  (
    G5_p_spl_110,
    G5_p_spl_11
  );


  buf

  (
    G5_p_spl_111,
    G5_p_spl_11
  );


  buf

  (
    G5_n_spl_,
    G5_n
  );


  buf

  (
    G5_n_spl_0,
    G5_n_spl_
  );


  buf

  (
    G5_n_spl_00,
    G5_n_spl_0
  );


  buf

  (
    G5_n_spl_000,
    G5_n_spl_00
  );


  buf

  (
    G5_n_spl_001,
    G5_n_spl_00
  );


  buf

  (
    G5_n_spl_01,
    G5_n_spl_0
  );


  buf

  (
    G5_n_spl_010,
    G5_n_spl_01
  );


  buf

  (
    G5_n_spl_011,
    G5_n_spl_01
  );


  buf

  (
    G5_n_spl_1,
    G5_n_spl_
  );


  buf

  (
    G5_n_spl_10,
    G5_n_spl_1
  );


  buf

  (
    G5_n_spl_100,
    G5_n_spl_10
  );


  buf

  (
    G5_n_spl_101,
    G5_n_spl_10
  );


  buf

  (
    G5_n_spl_11,
    G5_n_spl_1
  );


  buf

  (
    G5_n_spl_110,
    G5_n_spl_11
  );


  buf

  (
    G5_n_spl_111,
    G5_n_spl_11
  );


  buf

  (
    g80_n_spl_,
    g80_n
  );


  buf

  (
    g79_p_spl_,
    g79_p
  );


  buf

  (
    g80_p_spl_,
    g80_p
  );


  buf

  (
    g79_n_spl_,
    g79_n
  );


  buf

  (
    g81_n_spl_,
    g81_n
  );


  buf

  (
    g81_p_spl_,
    g81_p
  );


  buf

  (
    g82_n_spl_,
    g82_n
  );


  buf

  (
    g82_n_spl_0,
    g82_n_spl_
  );


  buf

  (
    g82_p_spl_,
    g82_p
  );


  buf

  (
    g82_p_spl_0,
    g82_p_spl_
  );


  buf

  (
    g84_n_spl_,
    g84_n
  );


  buf

  (
    g84_p_spl_,
    g84_p
  );


  buf

  (
    g85_n_spl_,
    g85_n
  );


  buf

  (
    g85_p_spl_,
    g85_p
  );


  buf

  (
    g87_p_spl_,
    g87_p
  );


  buf

  (
    g78_n_spl_,
    g78_n
  );


  buf

  (
    g87_n_spl_,
    g87_n
  );


  buf

  (
    g78_p_spl_,
    g78_p
  );


  buf

  (
    g88_n_spl_,
    g88_n
  );


  buf

  (
    g88_p_spl_,
    g88_p
  );


  buf

  (
    g90_p_spl_,
    g90_p
  );


  buf

  (
    g77_n_spl_,
    g77_n
  );


  buf

  (
    g90_n_spl_,
    g90_n
  );


  buf

  (
    g77_p_spl_,
    g77_p
  );


  buf

  (
    g91_n_spl_,
    g91_n
  );


  buf

  (
    g91_p_spl_,
    g91_p
  );


  buf

  (
    g93_p_spl_,
    g93_p
  );


  buf

  (
    g76_n_spl_,
    g76_n
  );


  buf

  (
    g93_n_spl_,
    g93_n
  );


  buf

  (
    g76_p_spl_,
    g76_p
  );


  buf

  (
    g94_n_spl_,
    g94_n
  );


  buf

  (
    g94_p_spl_,
    g94_p
  );


  buf

  (
    g96_p_spl_,
    g96_p
  );


  buf

  (
    g75_n_spl_,
    g75_n
  );


  buf

  (
    g96_n_spl_,
    g96_n
  );


  buf

  (
    g75_p_spl_,
    g75_p
  );


  buf

  (
    g97_n_spl_,
    g97_n
  );


  buf

  (
    g97_p_spl_,
    g97_p
  );


  buf

  (
    g99_n_spl_,
    g99_n
  );


  buf

  (
    g74_p_spl_,
    g74_p
  );


  buf

  (
    g100_p_spl_,
    g100_p
  );


  buf

  (
    G22_p_spl_,
    G22_p
  );


  buf

  (
    G22_p_spl_0,
    G22_p_spl_
  );


  buf

  (
    G22_p_spl_00,
    G22_p_spl_0
  );


  buf

  (
    G22_p_spl_000,
    G22_p_spl_00
  );


  buf

  (
    G22_p_spl_001,
    G22_p_spl_00
  );


  buf

  (
    G22_p_spl_01,
    G22_p_spl_0
  );


  buf

  (
    G22_p_spl_010,
    G22_p_spl_01
  );


  buf

  (
    G22_p_spl_011,
    G22_p_spl_01
  );


  buf

  (
    G22_p_spl_1,
    G22_p_spl_
  );


  buf

  (
    G22_p_spl_10,
    G22_p_spl_1
  );


  buf

  (
    G22_p_spl_100,
    G22_p_spl_10
  );


  buf

  (
    G22_p_spl_101,
    G22_p_spl_10
  );


  buf

  (
    G22_p_spl_11,
    G22_p_spl_1
  );


  buf

  (
    G22_p_spl_110,
    G22_p_spl_11
  );


  buf

  (
    G22_p_spl_111,
    G22_p_spl_11
  );


  buf

  (
    G22_n_spl_,
    G22_n
  );


  buf

  (
    G22_n_spl_0,
    G22_n_spl_
  );


  buf

  (
    G22_n_spl_00,
    G22_n_spl_0
  );


  buf

  (
    G22_n_spl_000,
    G22_n_spl_00
  );


  buf

  (
    G22_n_spl_001,
    G22_n_spl_00
  );


  buf

  (
    G22_n_spl_01,
    G22_n_spl_0
  );


  buf

  (
    G22_n_spl_010,
    G22_n_spl_01
  );


  buf

  (
    G22_n_spl_011,
    G22_n_spl_01
  );


  buf

  (
    G22_n_spl_1,
    G22_n_spl_
  );


  buf

  (
    G22_n_spl_10,
    G22_n_spl_1
  );


  buf

  (
    G22_n_spl_100,
    G22_n_spl_10
  );


  buf

  (
    G22_n_spl_101,
    G22_n_spl_10
  );


  buf

  (
    G22_n_spl_11,
    G22_n_spl_1
  );


  buf

  (
    G22_n_spl_110,
    G22_n_spl_11
  );


  buf

  (
    G22_n_spl_111,
    G22_n_spl_11
  );


  buf

  (
    G6_p_spl_,
    G6_p
  );


  buf

  (
    G6_p_spl_0,
    G6_p_spl_
  );


  buf

  (
    G6_p_spl_00,
    G6_p_spl_0
  );


  buf

  (
    G6_p_spl_000,
    G6_p_spl_00
  );


  buf

  (
    G6_p_spl_001,
    G6_p_spl_00
  );


  buf

  (
    G6_p_spl_01,
    G6_p_spl_0
  );


  buf

  (
    G6_p_spl_010,
    G6_p_spl_01
  );


  buf

  (
    G6_p_spl_011,
    G6_p_spl_01
  );


  buf

  (
    G6_p_spl_1,
    G6_p_spl_
  );


  buf

  (
    G6_p_spl_10,
    G6_p_spl_1
  );


  buf

  (
    G6_p_spl_100,
    G6_p_spl_10
  );


  buf

  (
    G6_p_spl_101,
    G6_p_spl_10
  );


  buf

  (
    G6_p_spl_11,
    G6_p_spl_1
  );


  buf

  (
    G6_p_spl_110,
    G6_p_spl_11
  );


  buf

  (
    G6_p_spl_111,
    G6_p_spl_11
  );


  buf

  (
    G6_n_spl_,
    G6_n
  );


  buf

  (
    G6_n_spl_0,
    G6_n_spl_
  );


  buf

  (
    G6_n_spl_00,
    G6_n_spl_0
  );


  buf

  (
    G6_n_spl_000,
    G6_n_spl_00
  );


  buf

  (
    G6_n_spl_001,
    G6_n_spl_00
  );


  buf

  (
    G6_n_spl_01,
    G6_n_spl_0
  );


  buf

  (
    G6_n_spl_010,
    G6_n_spl_01
  );


  buf

  (
    G6_n_spl_011,
    G6_n_spl_01
  );


  buf

  (
    G6_n_spl_1,
    G6_n_spl_
  );


  buf

  (
    G6_n_spl_10,
    G6_n_spl_1
  );


  buf

  (
    G6_n_spl_100,
    G6_n_spl_10
  );


  buf

  (
    G6_n_spl_101,
    G6_n_spl_10
  );


  buf

  (
    G6_n_spl_11,
    G6_n_spl_1
  );


  buf

  (
    G6_n_spl_110,
    G6_n_spl_11
  );


  buf

  (
    G6_n_spl_111,
    G6_n_spl_11
  );


  buf

  (
    g111_n_spl_,
    g111_n
  );


  buf

  (
    g110_p_spl_,
    g110_p
  );


  buf

  (
    g111_p_spl_,
    g111_p
  );


  buf

  (
    g110_n_spl_,
    g110_n
  );


  buf

  (
    g112_n_spl_,
    g112_n
  );


  buf

  (
    g112_p_spl_,
    g112_p
  );


  buf

  (
    g113_n_spl_,
    g113_n
  );


  buf

  (
    g113_n_spl_0,
    g113_n_spl_
  );


  buf

  (
    g113_p_spl_,
    g113_p
  );


  buf

  (
    g113_p_spl_0,
    g113_p_spl_
  );


  buf

  (
    g115_n_spl_,
    g115_n
  );


  buf

  (
    g115_p_spl_,
    g115_p
  );


  buf

  (
    g116_n_spl_,
    g116_n
  );


  buf

  (
    g116_p_spl_,
    g116_p
  );


  buf

  (
    g118_p_spl_,
    g118_p
  );


  buf

  (
    g109_n_spl_,
    g109_n
  );


  buf

  (
    g118_n_spl_,
    g118_n
  );


  buf

  (
    g109_p_spl_,
    g109_p
  );


  buf

  (
    g119_n_spl_,
    g119_n
  );


  buf

  (
    g119_p_spl_,
    g119_p
  );


  buf

  (
    g121_p_spl_,
    g121_p
  );


  buf

  (
    g108_n_spl_,
    g108_n
  );


  buf

  (
    g121_n_spl_,
    g121_n
  );


  buf

  (
    g108_p_spl_,
    g108_p
  );


  buf

  (
    g122_n_spl_,
    g122_n
  );


  buf

  (
    g122_p_spl_,
    g122_p
  );


  buf

  (
    g124_p_spl_,
    g124_p
  );


  buf

  (
    g107_n_spl_,
    g107_n
  );


  buf

  (
    g124_n_spl_,
    g124_n
  );


  buf

  (
    g107_p_spl_,
    g107_p
  );


  buf

  (
    g125_n_spl_,
    g125_n
  );


  buf

  (
    g125_p_spl_,
    g125_p
  );


  buf

  (
    g127_p_spl_,
    g127_p
  );


  buf

  (
    g106_n_spl_,
    g106_n
  );


  buf

  (
    g127_n_spl_,
    g127_n
  );


  buf

  (
    g106_p_spl_,
    g106_p
  );


  buf

  (
    g128_n_spl_,
    g128_n
  );


  buf

  (
    g128_p_spl_,
    g128_p
  );


  buf

  (
    g130_p_spl_,
    g130_p
  );


  buf

  (
    g105_n_spl_,
    g105_n
  );


  buf

  (
    g130_n_spl_,
    g130_n
  );


  buf

  (
    g105_p_spl_,
    g105_p
  );


  buf

  (
    g131_n_spl_,
    g131_n
  );


  buf

  (
    g131_p_spl_,
    g131_p
  );


  buf

  (
    g133_p_spl_,
    g133_p
  );


  buf

  (
    g104_n_spl_,
    g104_n
  );


  buf

  (
    g133_n_spl_,
    g133_n
  );


  buf

  (
    g104_p_spl_,
    g104_p
  );


  buf

  (
    g134_n_spl_,
    g134_n
  );


  buf

  (
    g134_p_spl_,
    g134_p
  );


  buf

  (
    g136_n_spl_,
    g136_n
  );


  buf

  (
    g103_p_spl_,
    g103_p
  );


  buf

  (
    g137_p_spl_,
    g137_p
  );


  buf

  (
    G23_p_spl_,
    G23_p
  );


  buf

  (
    G23_p_spl_0,
    G23_p_spl_
  );


  buf

  (
    G23_p_spl_00,
    G23_p_spl_0
  );


  buf

  (
    G23_p_spl_000,
    G23_p_spl_00
  );


  buf

  (
    G23_p_spl_001,
    G23_p_spl_00
  );


  buf

  (
    G23_p_spl_01,
    G23_p_spl_0
  );


  buf

  (
    G23_p_spl_010,
    G23_p_spl_01
  );


  buf

  (
    G23_p_spl_011,
    G23_p_spl_01
  );


  buf

  (
    G23_p_spl_1,
    G23_p_spl_
  );


  buf

  (
    G23_p_spl_10,
    G23_p_spl_1
  );


  buf

  (
    G23_p_spl_100,
    G23_p_spl_10
  );


  buf

  (
    G23_p_spl_101,
    G23_p_spl_10
  );


  buf

  (
    G23_p_spl_11,
    G23_p_spl_1
  );


  buf

  (
    G23_p_spl_110,
    G23_p_spl_11
  );


  buf

  (
    G23_p_spl_111,
    G23_p_spl_11
  );


  buf

  (
    G23_n_spl_,
    G23_n
  );


  buf

  (
    G23_n_spl_0,
    G23_n_spl_
  );


  buf

  (
    G23_n_spl_00,
    G23_n_spl_0
  );


  buf

  (
    G23_n_spl_000,
    G23_n_spl_00
  );


  buf

  (
    G23_n_spl_001,
    G23_n_spl_00
  );


  buf

  (
    G23_n_spl_01,
    G23_n_spl_0
  );


  buf

  (
    G23_n_spl_010,
    G23_n_spl_01
  );


  buf

  (
    G23_n_spl_011,
    G23_n_spl_01
  );


  buf

  (
    G23_n_spl_1,
    G23_n_spl_
  );


  buf

  (
    G23_n_spl_10,
    G23_n_spl_1
  );


  buf

  (
    G23_n_spl_100,
    G23_n_spl_10
  );


  buf

  (
    G23_n_spl_101,
    G23_n_spl_10
  );


  buf

  (
    G23_n_spl_11,
    G23_n_spl_1
  );


  buf

  (
    G23_n_spl_110,
    G23_n_spl_11
  );


  buf

  (
    G23_n_spl_111,
    G23_n_spl_11
  );


  buf

  (
    G7_p_spl_,
    G7_p
  );


  buf

  (
    G7_p_spl_0,
    G7_p_spl_
  );


  buf

  (
    G7_p_spl_00,
    G7_p_spl_0
  );


  buf

  (
    G7_p_spl_000,
    G7_p_spl_00
  );


  buf

  (
    G7_p_spl_001,
    G7_p_spl_00
  );


  buf

  (
    G7_p_spl_01,
    G7_p_spl_0
  );


  buf

  (
    G7_p_spl_010,
    G7_p_spl_01
  );


  buf

  (
    G7_p_spl_011,
    G7_p_spl_01
  );


  buf

  (
    G7_p_spl_1,
    G7_p_spl_
  );


  buf

  (
    G7_p_spl_10,
    G7_p_spl_1
  );


  buf

  (
    G7_p_spl_100,
    G7_p_spl_10
  );


  buf

  (
    G7_p_spl_101,
    G7_p_spl_10
  );


  buf

  (
    G7_p_spl_11,
    G7_p_spl_1
  );


  buf

  (
    G7_p_spl_110,
    G7_p_spl_11
  );


  buf

  (
    G7_p_spl_111,
    G7_p_spl_11
  );


  buf

  (
    G7_n_spl_,
    G7_n
  );


  buf

  (
    G7_n_spl_0,
    G7_n_spl_
  );


  buf

  (
    G7_n_spl_00,
    G7_n_spl_0
  );


  buf

  (
    G7_n_spl_000,
    G7_n_spl_00
  );


  buf

  (
    G7_n_spl_001,
    G7_n_spl_00
  );


  buf

  (
    G7_n_spl_01,
    G7_n_spl_0
  );


  buf

  (
    G7_n_spl_010,
    G7_n_spl_01
  );


  buf

  (
    G7_n_spl_011,
    G7_n_spl_01
  );


  buf

  (
    G7_n_spl_1,
    G7_n_spl_
  );


  buf

  (
    G7_n_spl_10,
    G7_n_spl_1
  );


  buf

  (
    G7_n_spl_100,
    G7_n_spl_10
  );


  buf

  (
    G7_n_spl_101,
    G7_n_spl_10
  );


  buf

  (
    G7_n_spl_11,
    G7_n_spl_1
  );


  buf

  (
    G7_n_spl_110,
    G7_n_spl_11
  );


  buf

  (
    G7_n_spl_111,
    G7_n_spl_11
  );


  buf

  (
    g150_n_spl_,
    g150_n
  );


  buf

  (
    g149_p_spl_,
    g149_p
  );


  buf

  (
    g150_p_spl_,
    g150_p
  );


  buf

  (
    g149_n_spl_,
    g149_n
  );


  buf

  (
    g151_n_spl_,
    g151_n
  );


  buf

  (
    g151_p_spl_,
    g151_p
  );


  buf

  (
    g152_n_spl_,
    g152_n
  );


  buf

  (
    g152_n_spl_0,
    g152_n_spl_
  );


  buf

  (
    g152_p_spl_,
    g152_p
  );


  buf

  (
    g152_p_spl_0,
    g152_p_spl_
  );


  buf

  (
    g154_n_spl_,
    g154_n
  );


  buf

  (
    g154_p_spl_,
    g154_p
  );


  buf

  (
    g155_n_spl_,
    g155_n
  );


  buf

  (
    g155_p_spl_,
    g155_p
  );


  buf

  (
    g157_p_spl_,
    g157_p
  );


  buf

  (
    g148_n_spl_,
    g148_n
  );


  buf

  (
    g157_n_spl_,
    g157_n
  );


  buf

  (
    g148_p_spl_,
    g148_p
  );


  buf

  (
    g158_n_spl_,
    g158_n
  );


  buf

  (
    g158_p_spl_,
    g158_p
  );


  buf

  (
    g160_p_spl_,
    g160_p
  );


  buf

  (
    g147_n_spl_,
    g147_n
  );


  buf

  (
    g160_n_spl_,
    g160_n
  );


  buf

  (
    g147_p_spl_,
    g147_p
  );


  buf

  (
    g161_n_spl_,
    g161_n
  );


  buf

  (
    g161_p_spl_,
    g161_p
  );


  buf

  (
    g163_p_spl_,
    g163_p
  );


  buf

  (
    g146_n_spl_,
    g146_n
  );


  buf

  (
    g163_n_spl_,
    g163_n
  );


  buf

  (
    g146_p_spl_,
    g146_p
  );


  buf

  (
    g164_n_spl_,
    g164_n
  );


  buf

  (
    g164_p_spl_,
    g164_p
  );


  buf

  (
    g166_p_spl_,
    g166_p
  );


  buf

  (
    g145_n_spl_,
    g145_n
  );


  buf

  (
    g166_n_spl_,
    g166_n
  );


  buf

  (
    g145_p_spl_,
    g145_p
  );


  buf

  (
    g167_n_spl_,
    g167_n
  );


  buf

  (
    g167_p_spl_,
    g167_p
  );


  buf

  (
    g169_p_spl_,
    g169_p
  );


  buf

  (
    g144_n_spl_,
    g144_n
  );


  buf

  (
    g169_n_spl_,
    g169_n
  );


  buf

  (
    g144_p_spl_,
    g144_p
  );


  buf

  (
    g170_n_spl_,
    g170_n
  );


  buf

  (
    g170_p_spl_,
    g170_p
  );


  buf

  (
    g172_p_spl_,
    g172_p
  );


  buf

  (
    g143_n_spl_,
    g143_n
  );


  buf

  (
    g172_n_spl_,
    g172_n
  );


  buf

  (
    g143_p_spl_,
    g143_p
  );


  buf

  (
    g173_n_spl_,
    g173_n
  );


  buf

  (
    g173_p_spl_,
    g173_p
  );


  buf

  (
    g175_p_spl_,
    g175_p
  );


  buf

  (
    g142_n_spl_,
    g142_n
  );


  buf

  (
    g175_n_spl_,
    g175_n
  );


  buf

  (
    g142_p_spl_,
    g142_p
  );


  buf

  (
    g176_n_spl_,
    g176_n
  );


  buf

  (
    g176_p_spl_,
    g176_p
  );


  buf

  (
    g178_p_spl_,
    g178_p
  );


  buf

  (
    g141_n_spl_,
    g141_n
  );


  buf

  (
    g178_n_spl_,
    g178_n
  );


  buf

  (
    g141_p_spl_,
    g141_p
  );


  buf

  (
    g179_n_spl_,
    g179_n
  );


  buf

  (
    g179_p_spl_,
    g179_p
  );


  buf

  (
    g181_n_spl_,
    g181_n
  );


  buf

  (
    g140_p_spl_,
    g140_p
  );


  buf

  (
    g182_p_spl_,
    g182_p
  );


  buf

  (
    G24_p_spl_,
    G24_p
  );


  buf

  (
    G24_p_spl_0,
    G24_p_spl_
  );


  buf

  (
    G24_p_spl_00,
    G24_p_spl_0
  );


  buf

  (
    G24_p_spl_000,
    G24_p_spl_00
  );


  buf

  (
    G24_p_spl_001,
    G24_p_spl_00
  );


  buf

  (
    G24_p_spl_01,
    G24_p_spl_0
  );


  buf

  (
    G24_p_spl_010,
    G24_p_spl_01
  );


  buf

  (
    G24_p_spl_011,
    G24_p_spl_01
  );


  buf

  (
    G24_p_spl_1,
    G24_p_spl_
  );


  buf

  (
    G24_p_spl_10,
    G24_p_spl_1
  );


  buf

  (
    G24_p_spl_100,
    G24_p_spl_10
  );


  buf

  (
    G24_p_spl_101,
    G24_p_spl_10
  );


  buf

  (
    G24_p_spl_11,
    G24_p_spl_1
  );


  buf

  (
    G24_p_spl_110,
    G24_p_spl_11
  );


  buf

  (
    G24_p_spl_111,
    G24_p_spl_11
  );


  buf

  (
    G24_n_spl_,
    G24_n
  );


  buf

  (
    G24_n_spl_0,
    G24_n_spl_
  );


  buf

  (
    G24_n_spl_00,
    G24_n_spl_0
  );


  buf

  (
    G24_n_spl_000,
    G24_n_spl_00
  );


  buf

  (
    G24_n_spl_001,
    G24_n_spl_00
  );


  buf

  (
    G24_n_spl_01,
    G24_n_spl_0
  );


  buf

  (
    G24_n_spl_010,
    G24_n_spl_01
  );


  buf

  (
    G24_n_spl_011,
    G24_n_spl_01
  );


  buf

  (
    G24_n_spl_1,
    G24_n_spl_
  );


  buf

  (
    G24_n_spl_10,
    G24_n_spl_1
  );


  buf

  (
    G24_n_spl_100,
    G24_n_spl_10
  );


  buf

  (
    G24_n_spl_101,
    G24_n_spl_10
  );


  buf

  (
    G24_n_spl_11,
    G24_n_spl_1
  );


  buf

  (
    G24_n_spl_110,
    G24_n_spl_11
  );


  buf

  (
    G24_n_spl_111,
    G24_n_spl_11
  );


  buf

  (
    G8_p_spl_,
    G8_p
  );


  buf

  (
    G8_p_spl_0,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_00,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_000,
    G8_p_spl_00
  );


  buf

  (
    G8_p_spl_001,
    G8_p_spl_00
  );


  buf

  (
    G8_p_spl_01,
    G8_p_spl_0
  );


  buf

  (
    G8_p_spl_010,
    G8_p_spl_01
  );


  buf

  (
    G8_p_spl_011,
    G8_p_spl_01
  );


  buf

  (
    G8_p_spl_1,
    G8_p_spl_
  );


  buf

  (
    G8_p_spl_10,
    G8_p_spl_1
  );


  buf

  (
    G8_p_spl_100,
    G8_p_spl_10
  );


  buf

  (
    G8_p_spl_101,
    G8_p_spl_10
  );


  buf

  (
    G8_p_spl_11,
    G8_p_spl_1
  );


  buf

  (
    G8_p_spl_110,
    G8_p_spl_11
  );


  buf

  (
    G8_p_spl_111,
    G8_p_spl_11
  );


  buf

  (
    G8_n_spl_,
    G8_n
  );


  buf

  (
    G8_n_spl_0,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_00,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_000,
    G8_n_spl_00
  );


  buf

  (
    G8_n_spl_001,
    G8_n_spl_00
  );


  buf

  (
    G8_n_spl_01,
    G8_n_spl_0
  );


  buf

  (
    G8_n_spl_010,
    G8_n_spl_01
  );


  buf

  (
    G8_n_spl_011,
    G8_n_spl_01
  );


  buf

  (
    G8_n_spl_1,
    G8_n_spl_
  );


  buf

  (
    G8_n_spl_10,
    G8_n_spl_1
  );


  buf

  (
    G8_n_spl_100,
    G8_n_spl_10
  );


  buf

  (
    G8_n_spl_101,
    G8_n_spl_10
  );


  buf

  (
    G8_n_spl_11,
    G8_n_spl_1
  );


  buf

  (
    G8_n_spl_110,
    G8_n_spl_11
  );


  buf

  (
    G8_n_spl_111,
    G8_n_spl_11
  );


  buf

  (
    g197_n_spl_,
    g197_n
  );


  buf

  (
    g196_p_spl_,
    g196_p
  );


  buf

  (
    g197_p_spl_,
    g197_p
  );


  buf

  (
    g196_n_spl_,
    g196_n
  );


  buf

  (
    g198_n_spl_,
    g198_n
  );


  buf

  (
    g198_p_spl_,
    g198_p
  );


  buf

  (
    g199_n_spl_,
    g199_n
  );


  buf

  (
    g199_n_spl_0,
    g199_n_spl_
  );


  buf

  (
    g199_p_spl_,
    g199_p
  );


  buf

  (
    g199_p_spl_0,
    g199_p_spl_
  );


  buf

  (
    g201_n_spl_,
    g201_n
  );


  buf

  (
    g201_p_spl_,
    g201_p
  );


  buf

  (
    g202_n_spl_,
    g202_n
  );


  buf

  (
    g202_p_spl_,
    g202_p
  );


  buf

  (
    g204_p_spl_,
    g204_p
  );


  buf

  (
    g195_n_spl_,
    g195_n
  );


  buf

  (
    g204_n_spl_,
    g204_n
  );


  buf

  (
    g195_p_spl_,
    g195_p
  );


  buf

  (
    g205_n_spl_,
    g205_n
  );


  buf

  (
    g205_p_spl_,
    g205_p
  );


  buf

  (
    g207_p_spl_,
    g207_p
  );


  buf

  (
    g194_n_spl_,
    g194_n
  );


  buf

  (
    g207_n_spl_,
    g207_n
  );


  buf

  (
    g194_p_spl_,
    g194_p
  );


  buf

  (
    g208_n_spl_,
    g208_n
  );


  buf

  (
    g208_p_spl_,
    g208_p
  );


  buf

  (
    g210_p_spl_,
    g210_p
  );


  buf

  (
    g193_n_spl_,
    g193_n
  );


  buf

  (
    g210_n_spl_,
    g210_n
  );


  buf

  (
    g193_p_spl_,
    g193_p
  );


  buf

  (
    g211_n_spl_,
    g211_n
  );


  buf

  (
    g211_p_spl_,
    g211_p
  );


  buf

  (
    g213_p_spl_,
    g213_p
  );


  buf

  (
    g192_n_spl_,
    g192_n
  );


  buf

  (
    g213_n_spl_,
    g213_n
  );


  buf

  (
    g192_p_spl_,
    g192_p
  );


  buf

  (
    g214_n_spl_,
    g214_n
  );


  buf

  (
    g214_p_spl_,
    g214_p
  );


  buf

  (
    g216_p_spl_,
    g216_p
  );


  buf

  (
    g191_n_spl_,
    g191_n
  );


  buf

  (
    g216_n_spl_,
    g216_n
  );


  buf

  (
    g191_p_spl_,
    g191_p
  );


  buf

  (
    g217_n_spl_,
    g217_n
  );


  buf

  (
    g217_p_spl_,
    g217_p
  );


  buf

  (
    g219_p_spl_,
    g219_p
  );


  buf

  (
    g190_n_spl_,
    g190_n
  );


  buf

  (
    g219_n_spl_,
    g219_n
  );


  buf

  (
    g190_p_spl_,
    g190_p
  );


  buf

  (
    g220_n_spl_,
    g220_n
  );


  buf

  (
    g220_p_spl_,
    g220_p
  );


  buf

  (
    g222_p_spl_,
    g222_p
  );


  buf

  (
    g189_n_spl_,
    g189_n
  );


  buf

  (
    g222_n_spl_,
    g222_n
  );


  buf

  (
    g189_p_spl_,
    g189_p
  );


  buf

  (
    g223_n_spl_,
    g223_n
  );


  buf

  (
    g223_p_spl_,
    g223_p
  );


  buf

  (
    g225_p_spl_,
    g225_p
  );


  buf

  (
    g188_n_spl_,
    g188_n
  );


  buf

  (
    g225_n_spl_,
    g225_n
  );


  buf

  (
    g188_p_spl_,
    g188_p
  );


  buf

  (
    g226_n_spl_,
    g226_n
  );


  buf

  (
    g226_p_spl_,
    g226_p
  );


  buf

  (
    g228_p_spl_,
    g228_p
  );


  buf

  (
    g187_n_spl_,
    g187_n
  );


  buf

  (
    g228_n_spl_,
    g228_n
  );


  buf

  (
    g187_p_spl_,
    g187_p
  );


  buf

  (
    g229_n_spl_,
    g229_n
  );


  buf

  (
    g229_p_spl_,
    g229_p
  );


  buf

  (
    g231_p_spl_,
    g231_p
  );


  buf

  (
    g186_n_spl_,
    g186_n
  );


  buf

  (
    g231_n_spl_,
    g231_n
  );


  buf

  (
    g186_p_spl_,
    g186_p
  );


  buf

  (
    g232_n_spl_,
    g232_n
  );


  buf

  (
    g232_p_spl_,
    g232_p
  );


  buf

  (
    g234_n_spl_,
    g234_n
  );


  buf

  (
    g185_p_spl_,
    g185_p
  );


  buf

  (
    g235_p_spl_,
    g235_p
  );


  buf

  (
    G25_p_spl_,
    G25_p
  );


  buf

  (
    G25_p_spl_0,
    G25_p_spl_
  );


  buf

  (
    G25_p_spl_00,
    G25_p_spl_0
  );


  buf

  (
    G25_p_spl_000,
    G25_p_spl_00
  );


  buf

  (
    G25_p_spl_001,
    G25_p_spl_00
  );


  buf

  (
    G25_p_spl_01,
    G25_p_spl_0
  );


  buf

  (
    G25_p_spl_010,
    G25_p_spl_01
  );


  buf

  (
    G25_p_spl_011,
    G25_p_spl_01
  );


  buf

  (
    G25_p_spl_1,
    G25_p_spl_
  );


  buf

  (
    G25_p_spl_10,
    G25_p_spl_1
  );


  buf

  (
    G25_p_spl_100,
    G25_p_spl_10
  );


  buf

  (
    G25_p_spl_101,
    G25_p_spl_10
  );


  buf

  (
    G25_p_spl_11,
    G25_p_spl_1
  );


  buf

  (
    G25_p_spl_110,
    G25_p_spl_11
  );


  buf

  (
    G25_p_spl_111,
    G25_p_spl_11
  );


  buf

  (
    G25_n_spl_,
    G25_n
  );


  buf

  (
    G25_n_spl_0,
    G25_n_spl_
  );


  buf

  (
    G25_n_spl_00,
    G25_n_spl_0
  );


  buf

  (
    G25_n_spl_000,
    G25_n_spl_00
  );


  buf

  (
    G25_n_spl_001,
    G25_n_spl_00
  );


  buf

  (
    G25_n_spl_01,
    G25_n_spl_0
  );


  buf

  (
    G25_n_spl_010,
    G25_n_spl_01
  );


  buf

  (
    G25_n_spl_011,
    G25_n_spl_01
  );


  buf

  (
    G25_n_spl_1,
    G25_n_spl_
  );


  buf

  (
    G25_n_spl_10,
    G25_n_spl_1
  );


  buf

  (
    G25_n_spl_100,
    G25_n_spl_10
  );


  buf

  (
    G25_n_spl_101,
    G25_n_spl_10
  );


  buf

  (
    G25_n_spl_11,
    G25_n_spl_1
  );


  buf

  (
    G25_n_spl_110,
    G25_n_spl_11
  );


  buf

  (
    G25_n_spl_111,
    G25_n_spl_11
  );


  buf

  (
    G9_p_spl_,
    G9_p
  );


  buf

  (
    G9_p_spl_0,
    G9_p_spl_
  );


  buf

  (
    G9_p_spl_00,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_000,
    G9_p_spl_00
  );


  buf

  (
    G9_p_spl_001,
    G9_p_spl_00
  );


  buf

  (
    G9_p_spl_01,
    G9_p_spl_0
  );


  buf

  (
    G9_p_spl_010,
    G9_p_spl_01
  );


  buf

  (
    G9_p_spl_011,
    G9_p_spl_01
  );


  buf

  (
    G9_p_spl_1,
    G9_p_spl_
  );


  buf

  (
    G9_p_spl_10,
    G9_p_spl_1
  );


  buf

  (
    G9_p_spl_100,
    G9_p_spl_10
  );


  buf

  (
    G9_p_spl_101,
    G9_p_spl_10
  );


  buf

  (
    G9_p_spl_11,
    G9_p_spl_1
  );


  buf

  (
    G9_p_spl_110,
    G9_p_spl_11
  );


  buf

  (
    G9_p_spl_111,
    G9_p_spl_11
  );


  buf

  (
    G9_n_spl_,
    G9_n
  );


  buf

  (
    G9_n_spl_0,
    G9_n_spl_
  );


  buf

  (
    G9_n_spl_00,
    G9_n_spl_0
  );


  buf

  (
    G9_n_spl_000,
    G9_n_spl_00
  );


  buf

  (
    G9_n_spl_001,
    G9_n_spl_00
  );


  buf

  (
    G9_n_spl_01,
    G9_n_spl_0
  );


  buf

  (
    G9_n_spl_010,
    G9_n_spl_01
  );


  buf

  (
    G9_n_spl_011,
    G9_n_spl_01
  );


  buf

  (
    G9_n_spl_1,
    G9_n_spl_
  );


  buf

  (
    G9_n_spl_10,
    G9_n_spl_1
  );


  buf

  (
    G9_n_spl_100,
    G9_n_spl_10
  );


  buf

  (
    G9_n_spl_101,
    G9_n_spl_10
  );


  buf

  (
    G9_n_spl_11,
    G9_n_spl_1
  );


  buf

  (
    G9_n_spl_110,
    G9_n_spl_11
  );


  buf

  (
    G9_n_spl_111,
    G9_n_spl_11
  );


  buf

  (
    g252_n_spl_,
    g252_n
  );


  buf

  (
    g251_p_spl_,
    g251_p
  );


  buf

  (
    g252_p_spl_,
    g252_p
  );


  buf

  (
    g251_n_spl_,
    g251_n
  );


  buf

  (
    g253_n_spl_,
    g253_n
  );


  buf

  (
    g253_p_spl_,
    g253_p
  );


  buf

  (
    g254_n_spl_,
    g254_n
  );


  buf

  (
    g254_n_spl_0,
    g254_n_spl_
  );


  buf

  (
    g254_p_spl_,
    g254_p
  );


  buf

  (
    g254_p_spl_0,
    g254_p_spl_
  );


  buf

  (
    g256_n_spl_,
    g256_n
  );


  buf

  (
    g256_p_spl_,
    g256_p
  );


  buf

  (
    g257_n_spl_,
    g257_n
  );


  buf

  (
    g257_p_spl_,
    g257_p
  );


  buf

  (
    g259_p_spl_,
    g259_p
  );


  buf

  (
    g250_n_spl_,
    g250_n
  );


  buf

  (
    g259_n_spl_,
    g259_n
  );


  buf

  (
    g250_p_spl_,
    g250_p
  );


  buf

  (
    g260_n_spl_,
    g260_n
  );


  buf

  (
    g260_p_spl_,
    g260_p
  );


  buf

  (
    g262_p_spl_,
    g262_p
  );


  buf

  (
    g249_n_spl_,
    g249_n
  );


  buf

  (
    g262_n_spl_,
    g262_n
  );


  buf

  (
    g249_p_spl_,
    g249_p
  );


  buf

  (
    g263_n_spl_,
    g263_n
  );


  buf

  (
    g263_p_spl_,
    g263_p
  );


  buf

  (
    g265_p_spl_,
    g265_p
  );


  buf

  (
    g248_n_spl_,
    g248_n
  );


  buf

  (
    g265_n_spl_,
    g265_n
  );


  buf

  (
    g248_p_spl_,
    g248_p
  );


  buf

  (
    g266_n_spl_,
    g266_n
  );


  buf

  (
    g266_p_spl_,
    g266_p
  );


  buf

  (
    g268_p_spl_,
    g268_p
  );


  buf

  (
    g247_n_spl_,
    g247_n
  );


  buf

  (
    g268_n_spl_,
    g268_n
  );


  buf

  (
    g247_p_spl_,
    g247_p
  );


  buf

  (
    g269_n_spl_,
    g269_n
  );


  buf

  (
    g269_p_spl_,
    g269_p
  );


  buf

  (
    g271_p_spl_,
    g271_p
  );


  buf

  (
    g246_n_spl_,
    g246_n
  );


  buf

  (
    g271_n_spl_,
    g271_n
  );


  buf

  (
    g246_p_spl_,
    g246_p
  );


  buf

  (
    g272_n_spl_,
    g272_n
  );


  buf

  (
    g272_p_spl_,
    g272_p
  );


  buf

  (
    g274_p_spl_,
    g274_p
  );


  buf

  (
    g245_n_spl_,
    g245_n
  );


  buf

  (
    g274_n_spl_,
    g274_n
  );


  buf

  (
    g245_p_spl_,
    g245_p
  );


  buf

  (
    g275_n_spl_,
    g275_n
  );


  buf

  (
    g275_p_spl_,
    g275_p
  );


  buf

  (
    g277_p_spl_,
    g277_p
  );


  buf

  (
    g244_n_spl_,
    g244_n
  );


  buf

  (
    g277_n_spl_,
    g277_n
  );


  buf

  (
    g244_p_spl_,
    g244_p
  );


  buf

  (
    g278_n_spl_,
    g278_n
  );


  buf

  (
    g278_p_spl_,
    g278_p
  );


  buf

  (
    g280_p_spl_,
    g280_p
  );


  buf

  (
    g243_n_spl_,
    g243_n
  );


  buf

  (
    g280_n_spl_,
    g280_n
  );


  buf

  (
    g243_p_spl_,
    g243_p
  );


  buf

  (
    g281_n_spl_,
    g281_n
  );


  buf

  (
    g281_p_spl_,
    g281_p
  );


  buf

  (
    g283_p_spl_,
    g283_p
  );


  buf

  (
    g242_n_spl_,
    g242_n
  );


  buf

  (
    g283_n_spl_,
    g283_n
  );


  buf

  (
    g242_p_spl_,
    g242_p
  );


  buf

  (
    g284_n_spl_,
    g284_n
  );


  buf

  (
    g284_p_spl_,
    g284_p
  );


  buf

  (
    g286_p_spl_,
    g286_p
  );


  buf

  (
    g241_n_spl_,
    g241_n
  );


  buf

  (
    g286_n_spl_,
    g286_n
  );


  buf

  (
    g241_p_spl_,
    g241_p
  );


  buf

  (
    g287_n_spl_,
    g287_n
  );


  buf

  (
    g287_p_spl_,
    g287_p
  );


  buf

  (
    g289_p_spl_,
    g289_p
  );


  buf

  (
    g240_n_spl_,
    g240_n
  );


  buf

  (
    g289_n_spl_,
    g289_n
  );


  buf

  (
    g240_p_spl_,
    g240_p
  );


  buf

  (
    g290_n_spl_,
    g290_n
  );


  buf

  (
    g290_p_spl_,
    g290_p
  );


  buf

  (
    g292_p_spl_,
    g292_p
  );


  buf

  (
    g239_n_spl_,
    g239_n
  );


  buf

  (
    g292_n_spl_,
    g292_n
  );


  buf

  (
    g239_p_spl_,
    g239_p
  );


  buf

  (
    g293_n_spl_,
    g293_n
  );


  buf

  (
    g293_p_spl_,
    g293_p
  );


  buf

  (
    g295_n_spl_,
    g295_n
  );


  buf

  (
    g238_p_spl_,
    g238_p
  );


  buf

  (
    g296_p_spl_,
    g296_p
  );


  buf

  (
    G26_p_spl_,
    G26_p
  );


  buf

  (
    G26_p_spl_0,
    G26_p_spl_
  );


  buf

  (
    G26_p_spl_00,
    G26_p_spl_0
  );


  buf

  (
    G26_p_spl_000,
    G26_p_spl_00
  );


  buf

  (
    G26_p_spl_001,
    G26_p_spl_00
  );


  buf

  (
    G26_p_spl_01,
    G26_p_spl_0
  );


  buf

  (
    G26_p_spl_010,
    G26_p_spl_01
  );


  buf

  (
    G26_p_spl_011,
    G26_p_spl_01
  );


  buf

  (
    G26_p_spl_1,
    G26_p_spl_
  );


  buf

  (
    G26_p_spl_10,
    G26_p_spl_1
  );


  buf

  (
    G26_p_spl_100,
    G26_p_spl_10
  );


  buf

  (
    G26_p_spl_101,
    G26_p_spl_10
  );


  buf

  (
    G26_p_spl_11,
    G26_p_spl_1
  );


  buf

  (
    G26_p_spl_110,
    G26_p_spl_11
  );


  buf

  (
    G26_p_spl_111,
    G26_p_spl_11
  );


  buf

  (
    G26_n_spl_,
    G26_n
  );


  buf

  (
    G26_n_spl_0,
    G26_n_spl_
  );


  buf

  (
    G26_n_spl_00,
    G26_n_spl_0
  );


  buf

  (
    G26_n_spl_000,
    G26_n_spl_00
  );


  buf

  (
    G26_n_spl_001,
    G26_n_spl_00
  );


  buf

  (
    G26_n_spl_01,
    G26_n_spl_0
  );


  buf

  (
    G26_n_spl_010,
    G26_n_spl_01
  );


  buf

  (
    G26_n_spl_011,
    G26_n_spl_01
  );


  buf

  (
    G26_n_spl_1,
    G26_n_spl_
  );


  buf

  (
    G26_n_spl_10,
    G26_n_spl_1
  );


  buf

  (
    G26_n_spl_100,
    G26_n_spl_10
  );


  buf

  (
    G26_n_spl_101,
    G26_n_spl_10
  );


  buf

  (
    G26_n_spl_11,
    G26_n_spl_1
  );


  buf

  (
    G26_n_spl_110,
    G26_n_spl_11
  );


  buf

  (
    G26_n_spl_111,
    G26_n_spl_11
  );


  buf

  (
    G10_p_spl_,
    G10_p
  );


  buf

  (
    G10_p_spl_0,
    G10_p_spl_
  );


  buf

  (
    G10_p_spl_00,
    G10_p_spl_0
  );


  buf

  (
    G10_p_spl_000,
    G10_p_spl_00
  );


  buf

  (
    G10_p_spl_001,
    G10_p_spl_00
  );


  buf

  (
    G10_p_spl_01,
    G10_p_spl_0
  );


  buf

  (
    G10_p_spl_010,
    G10_p_spl_01
  );


  buf

  (
    G10_p_spl_011,
    G10_p_spl_01
  );


  buf

  (
    G10_p_spl_1,
    G10_p_spl_
  );


  buf

  (
    G10_p_spl_10,
    G10_p_spl_1
  );


  buf

  (
    G10_p_spl_100,
    G10_p_spl_10
  );


  buf

  (
    G10_p_spl_101,
    G10_p_spl_10
  );


  buf

  (
    G10_p_spl_11,
    G10_p_spl_1
  );


  buf

  (
    G10_p_spl_110,
    G10_p_spl_11
  );


  buf

  (
    G10_p_spl_111,
    G10_p_spl_11
  );


  buf

  (
    G10_n_spl_,
    G10_n
  );


  buf

  (
    G10_n_spl_0,
    G10_n_spl_
  );


  buf

  (
    G10_n_spl_00,
    G10_n_spl_0
  );


  buf

  (
    G10_n_spl_000,
    G10_n_spl_00
  );


  buf

  (
    G10_n_spl_001,
    G10_n_spl_00
  );


  buf

  (
    G10_n_spl_01,
    G10_n_spl_0
  );


  buf

  (
    G10_n_spl_010,
    G10_n_spl_01
  );


  buf

  (
    G10_n_spl_011,
    G10_n_spl_01
  );


  buf

  (
    G10_n_spl_1,
    G10_n_spl_
  );


  buf

  (
    G10_n_spl_10,
    G10_n_spl_1
  );


  buf

  (
    G10_n_spl_100,
    G10_n_spl_10
  );


  buf

  (
    G10_n_spl_101,
    G10_n_spl_10
  );


  buf

  (
    G10_n_spl_11,
    G10_n_spl_1
  );


  buf

  (
    G10_n_spl_110,
    G10_n_spl_11
  );


  buf

  (
    G10_n_spl_111,
    G10_n_spl_11
  );


  buf

  (
    g315_n_spl_,
    g315_n
  );


  buf

  (
    g314_p_spl_,
    g314_p
  );


  buf

  (
    g315_p_spl_,
    g315_p
  );


  buf

  (
    g314_n_spl_,
    g314_n
  );


  buf

  (
    g316_n_spl_,
    g316_n
  );


  buf

  (
    g316_p_spl_,
    g316_p
  );


  buf

  (
    g317_n_spl_,
    g317_n
  );


  buf

  (
    g317_n_spl_0,
    g317_n_spl_
  );


  buf

  (
    g317_p_spl_,
    g317_p
  );


  buf

  (
    g317_p_spl_0,
    g317_p_spl_
  );


  buf

  (
    g319_n_spl_,
    g319_n
  );


  buf

  (
    g319_p_spl_,
    g319_p
  );


  buf

  (
    g320_n_spl_,
    g320_n
  );


  buf

  (
    g320_p_spl_,
    g320_p
  );


  buf

  (
    g322_p_spl_,
    g322_p
  );


  buf

  (
    g313_n_spl_,
    g313_n
  );


  buf

  (
    g322_n_spl_,
    g322_n
  );


  buf

  (
    g313_p_spl_,
    g313_p
  );


  buf

  (
    g323_n_spl_,
    g323_n
  );


  buf

  (
    g323_p_spl_,
    g323_p
  );


  buf

  (
    g325_p_spl_,
    g325_p
  );


  buf

  (
    g312_n_spl_,
    g312_n
  );


  buf

  (
    g325_n_spl_,
    g325_n
  );


  buf

  (
    g312_p_spl_,
    g312_p
  );


  buf

  (
    g326_n_spl_,
    g326_n
  );


  buf

  (
    g326_p_spl_,
    g326_p
  );


  buf

  (
    g328_p_spl_,
    g328_p
  );


  buf

  (
    g311_n_spl_,
    g311_n
  );


  buf

  (
    g328_n_spl_,
    g328_n
  );


  buf

  (
    g311_p_spl_,
    g311_p
  );


  buf

  (
    g329_n_spl_,
    g329_n
  );


  buf

  (
    g329_p_spl_,
    g329_p
  );


  buf

  (
    g331_p_spl_,
    g331_p
  );


  buf

  (
    g310_n_spl_,
    g310_n
  );


  buf

  (
    g331_n_spl_,
    g331_n
  );


  buf

  (
    g310_p_spl_,
    g310_p
  );


  buf

  (
    g332_n_spl_,
    g332_n
  );


  buf

  (
    g332_p_spl_,
    g332_p
  );


  buf

  (
    g334_p_spl_,
    g334_p
  );


  buf

  (
    g309_n_spl_,
    g309_n
  );


  buf

  (
    g334_n_spl_,
    g334_n
  );


  buf

  (
    g309_p_spl_,
    g309_p
  );


  buf

  (
    g335_n_spl_,
    g335_n
  );


  buf

  (
    g335_p_spl_,
    g335_p
  );


  buf

  (
    g337_p_spl_,
    g337_p
  );


  buf

  (
    g308_n_spl_,
    g308_n
  );


  buf

  (
    g337_n_spl_,
    g337_n
  );


  buf

  (
    g308_p_spl_,
    g308_p
  );


  buf

  (
    g338_n_spl_,
    g338_n
  );


  buf

  (
    g338_p_spl_,
    g338_p
  );


  buf

  (
    g340_p_spl_,
    g340_p
  );


  buf

  (
    g307_n_spl_,
    g307_n
  );


  buf

  (
    g340_n_spl_,
    g340_n
  );


  buf

  (
    g307_p_spl_,
    g307_p
  );


  buf

  (
    g341_n_spl_,
    g341_n
  );


  buf

  (
    g341_p_spl_,
    g341_p
  );


  buf

  (
    g343_p_spl_,
    g343_p
  );


  buf

  (
    g306_n_spl_,
    g306_n
  );


  buf

  (
    g343_n_spl_,
    g343_n
  );


  buf

  (
    g306_p_spl_,
    g306_p
  );


  buf

  (
    g344_n_spl_,
    g344_n
  );


  buf

  (
    g344_p_spl_,
    g344_p
  );


  buf

  (
    g346_p_spl_,
    g346_p
  );


  buf

  (
    g305_n_spl_,
    g305_n
  );


  buf

  (
    g346_n_spl_,
    g346_n
  );


  buf

  (
    g305_p_spl_,
    g305_p
  );


  buf

  (
    g347_n_spl_,
    g347_n
  );


  buf

  (
    g347_p_spl_,
    g347_p
  );


  buf

  (
    g349_p_spl_,
    g349_p
  );


  buf

  (
    g304_n_spl_,
    g304_n
  );


  buf

  (
    g349_n_spl_,
    g349_n
  );


  buf

  (
    g304_p_spl_,
    g304_p
  );


  buf

  (
    g350_n_spl_,
    g350_n
  );


  buf

  (
    g350_p_spl_,
    g350_p
  );


  buf

  (
    g352_p_spl_,
    g352_p
  );


  buf

  (
    g303_n_spl_,
    g303_n
  );


  buf

  (
    g352_n_spl_,
    g352_n
  );


  buf

  (
    g303_p_spl_,
    g303_p
  );


  buf

  (
    g353_n_spl_,
    g353_n
  );


  buf

  (
    g353_p_spl_,
    g353_p
  );


  buf

  (
    g355_p_spl_,
    g355_p
  );


  buf

  (
    g302_n_spl_,
    g302_n
  );


  buf

  (
    g355_n_spl_,
    g355_n
  );


  buf

  (
    g302_p_spl_,
    g302_p
  );


  buf

  (
    g356_n_spl_,
    g356_n
  );


  buf

  (
    g356_p_spl_,
    g356_p
  );


  buf

  (
    g358_p_spl_,
    g358_p
  );


  buf

  (
    g301_n_spl_,
    g301_n
  );


  buf

  (
    g358_n_spl_,
    g358_n
  );


  buf

  (
    g301_p_spl_,
    g301_p
  );


  buf

  (
    g359_n_spl_,
    g359_n
  );


  buf

  (
    g359_p_spl_,
    g359_p
  );


  buf

  (
    g361_p_spl_,
    g361_p
  );


  buf

  (
    g300_n_spl_,
    g300_n
  );


  buf

  (
    g361_n_spl_,
    g361_n
  );


  buf

  (
    g300_p_spl_,
    g300_p
  );


  buf

  (
    g362_n_spl_,
    g362_n
  );


  buf

  (
    g362_p_spl_,
    g362_p
  );


  buf

  (
    g364_n_spl_,
    g364_n
  );


  buf

  (
    g299_p_spl_,
    g299_p
  );


  buf

  (
    g365_p_spl_,
    g365_p
  );


  buf

  (
    G27_p_spl_,
    G27_p
  );


  buf

  (
    G27_p_spl_0,
    G27_p_spl_
  );


  buf

  (
    G27_p_spl_00,
    G27_p_spl_0
  );


  buf

  (
    G27_p_spl_000,
    G27_p_spl_00
  );


  buf

  (
    G27_p_spl_001,
    G27_p_spl_00
  );


  buf

  (
    G27_p_spl_01,
    G27_p_spl_0
  );


  buf

  (
    G27_p_spl_010,
    G27_p_spl_01
  );


  buf

  (
    G27_p_spl_011,
    G27_p_spl_01
  );


  buf

  (
    G27_p_spl_1,
    G27_p_spl_
  );


  buf

  (
    G27_p_spl_10,
    G27_p_spl_1
  );


  buf

  (
    G27_p_spl_100,
    G27_p_spl_10
  );


  buf

  (
    G27_p_spl_101,
    G27_p_spl_10
  );


  buf

  (
    G27_p_spl_11,
    G27_p_spl_1
  );


  buf

  (
    G27_p_spl_110,
    G27_p_spl_11
  );


  buf

  (
    G27_p_spl_111,
    G27_p_spl_11
  );


  buf

  (
    G27_n_spl_,
    G27_n
  );


  buf

  (
    G27_n_spl_0,
    G27_n_spl_
  );


  buf

  (
    G27_n_spl_00,
    G27_n_spl_0
  );


  buf

  (
    G27_n_spl_000,
    G27_n_spl_00
  );


  buf

  (
    G27_n_spl_001,
    G27_n_spl_00
  );


  buf

  (
    G27_n_spl_01,
    G27_n_spl_0
  );


  buf

  (
    G27_n_spl_010,
    G27_n_spl_01
  );


  buf

  (
    G27_n_spl_011,
    G27_n_spl_01
  );


  buf

  (
    G27_n_spl_1,
    G27_n_spl_
  );


  buf

  (
    G27_n_spl_10,
    G27_n_spl_1
  );


  buf

  (
    G27_n_spl_100,
    G27_n_spl_10
  );


  buf

  (
    G27_n_spl_101,
    G27_n_spl_10
  );


  buf

  (
    G27_n_spl_11,
    G27_n_spl_1
  );


  buf

  (
    G27_n_spl_110,
    G27_n_spl_11
  );


  buf

  (
    G27_n_spl_111,
    G27_n_spl_11
  );


  buf

  (
    G11_p_spl_,
    G11_p
  );


  buf

  (
    G11_p_spl_0,
    G11_p_spl_
  );


  buf

  (
    G11_p_spl_00,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_000,
    G11_p_spl_00
  );


  buf

  (
    G11_p_spl_001,
    G11_p_spl_00
  );


  buf

  (
    G11_p_spl_01,
    G11_p_spl_0
  );


  buf

  (
    G11_p_spl_010,
    G11_p_spl_01
  );


  buf

  (
    G11_p_spl_011,
    G11_p_spl_01
  );


  buf

  (
    G11_p_spl_1,
    G11_p_spl_
  );


  buf

  (
    G11_p_spl_10,
    G11_p_spl_1
  );


  buf

  (
    G11_p_spl_100,
    G11_p_spl_10
  );


  buf

  (
    G11_p_spl_101,
    G11_p_spl_10
  );


  buf

  (
    G11_p_spl_11,
    G11_p_spl_1
  );


  buf

  (
    G11_p_spl_110,
    G11_p_spl_11
  );


  buf

  (
    G11_p_spl_111,
    G11_p_spl_11
  );


  buf

  (
    G11_n_spl_,
    G11_n
  );


  buf

  (
    G11_n_spl_0,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_00,
    G11_n_spl_0
  );


  buf

  (
    G11_n_spl_000,
    G11_n_spl_00
  );


  buf

  (
    G11_n_spl_001,
    G11_n_spl_00
  );


  buf

  (
    G11_n_spl_01,
    G11_n_spl_0
  );


  buf

  (
    G11_n_spl_010,
    G11_n_spl_01
  );


  buf

  (
    G11_n_spl_011,
    G11_n_spl_01
  );


  buf

  (
    G11_n_spl_1,
    G11_n_spl_
  );


  buf

  (
    G11_n_spl_10,
    G11_n_spl_1
  );


  buf

  (
    G11_n_spl_100,
    G11_n_spl_10
  );


  buf

  (
    G11_n_spl_101,
    G11_n_spl_10
  );


  buf

  (
    G11_n_spl_11,
    G11_n_spl_1
  );


  buf

  (
    G11_n_spl_110,
    G11_n_spl_11
  );


  buf

  (
    G11_n_spl_111,
    G11_n_spl_11
  );


  buf

  (
    g386_n_spl_,
    g386_n
  );


  buf

  (
    g385_p_spl_,
    g385_p
  );


  buf

  (
    g386_p_spl_,
    g386_p
  );


  buf

  (
    g385_n_spl_,
    g385_n
  );


  buf

  (
    g387_n_spl_,
    g387_n
  );


  buf

  (
    g387_p_spl_,
    g387_p
  );


  buf

  (
    g388_n_spl_,
    g388_n
  );


  buf

  (
    g388_n_spl_0,
    g388_n_spl_
  );


  buf

  (
    g388_p_spl_,
    g388_p
  );


  buf

  (
    g388_p_spl_0,
    g388_p_spl_
  );


  buf

  (
    g390_n_spl_,
    g390_n
  );


  buf

  (
    g390_p_spl_,
    g390_p
  );


  buf

  (
    g391_n_spl_,
    g391_n
  );


  buf

  (
    g391_p_spl_,
    g391_p
  );


  buf

  (
    g393_p_spl_,
    g393_p
  );


  buf

  (
    g384_n_spl_,
    g384_n
  );


  buf

  (
    g393_n_spl_,
    g393_n
  );


  buf

  (
    g384_p_spl_,
    g384_p
  );


  buf

  (
    g394_n_spl_,
    g394_n
  );


  buf

  (
    g394_p_spl_,
    g394_p
  );


  buf

  (
    g396_p_spl_,
    g396_p
  );


  buf

  (
    g383_n_spl_,
    g383_n
  );


  buf

  (
    g396_n_spl_,
    g396_n
  );


  buf

  (
    g383_p_spl_,
    g383_p
  );


  buf

  (
    g397_n_spl_,
    g397_n
  );


  buf

  (
    g397_p_spl_,
    g397_p
  );


  buf

  (
    g399_p_spl_,
    g399_p
  );


  buf

  (
    g382_n_spl_,
    g382_n
  );


  buf

  (
    g399_n_spl_,
    g399_n
  );


  buf

  (
    g382_p_spl_,
    g382_p
  );


  buf

  (
    g400_n_spl_,
    g400_n
  );


  buf

  (
    g400_p_spl_,
    g400_p
  );


  buf

  (
    g402_p_spl_,
    g402_p
  );


  buf

  (
    g381_n_spl_,
    g381_n
  );


  buf

  (
    g402_n_spl_,
    g402_n
  );


  buf

  (
    g381_p_spl_,
    g381_p
  );


  buf

  (
    g403_n_spl_,
    g403_n
  );


  buf

  (
    g403_p_spl_,
    g403_p
  );


  buf

  (
    g405_p_spl_,
    g405_p
  );


  buf

  (
    g380_n_spl_,
    g380_n
  );


  buf

  (
    g405_n_spl_,
    g405_n
  );


  buf

  (
    g380_p_spl_,
    g380_p
  );


  buf

  (
    g406_n_spl_,
    g406_n
  );


  buf

  (
    g406_p_spl_,
    g406_p
  );


  buf

  (
    g408_p_spl_,
    g408_p
  );


  buf

  (
    g379_n_spl_,
    g379_n
  );


  buf

  (
    g408_n_spl_,
    g408_n
  );


  buf

  (
    g379_p_spl_,
    g379_p
  );


  buf

  (
    g409_n_spl_,
    g409_n
  );


  buf

  (
    g409_p_spl_,
    g409_p
  );


  buf

  (
    g411_p_spl_,
    g411_p
  );


  buf

  (
    g378_n_spl_,
    g378_n
  );


  buf

  (
    g411_n_spl_,
    g411_n
  );


  buf

  (
    g378_p_spl_,
    g378_p
  );


  buf

  (
    g412_n_spl_,
    g412_n
  );


  buf

  (
    g412_p_spl_,
    g412_p
  );


  buf

  (
    g414_p_spl_,
    g414_p
  );


  buf

  (
    g377_n_spl_,
    g377_n
  );


  buf

  (
    g414_n_spl_,
    g414_n
  );


  buf

  (
    g377_p_spl_,
    g377_p
  );


  buf

  (
    g415_n_spl_,
    g415_n
  );


  buf

  (
    g415_p_spl_,
    g415_p
  );


  buf

  (
    g417_p_spl_,
    g417_p
  );


  buf

  (
    g376_n_spl_,
    g376_n
  );


  buf

  (
    g417_n_spl_,
    g417_n
  );


  buf

  (
    g376_p_spl_,
    g376_p
  );


  buf

  (
    g418_n_spl_,
    g418_n
  );


  buf

  (
    g418_p_spl_,
    g418_p
  );


  buf

  (
    g420_p_spl_,
    g420_p
  );


  buf

  (
    g375_n_spl_,
    g375_n
  );


  buf

  (
    g420_n_spl_,
    g420_n
  );


  buf

  (
    g375_p_spl_,
    g375_p
  );


  buf

  (
    g421_n_spl_,
    g421_n
  );


  buf

  (
    g421_p_spl_,
    g421_p
  );


  buf

  (
    g423_p_spl_,
    g423_p
  );


  buf

  (
    g374_n_spl_,
    g374_n
  );


  buf

  (
    g423_n_spl_,
    g423_n
  );


  buf

  (
    g374_p_spl_,
    g374_p
  );


  buf

  (
    g424_n_spl_,
    g424_n
  );


  buf

  (
    g424_p_spl_,
    g424_p
  );


  buf

  (
    g426_p_spl_,
    g426_p
  );


  buf

  (
    g373_n_spl_,
    g373_n
  );


  buf

  (
    g426_n_spl_,
    g426_n
  );


  buf

  (
    g373_p_spl_,
    g373_p
  );


  buf

  (
    g427_n_spl_,
    g427_n
  );


  buf

  (
    g427_p_spl_,
    g427_p
  );


  buf

  (
    g429_p_spl_,
    g429_p
  );


  buf

  (
    g372_n_spl_,
    g372_n
  );


  buf

  (
    g429_n_spl_,
    g429_n
  );


  buf

  (
    g372_p_spl_,
    g372_p
  );


  buf

  (
    g430_n_spl_,
    g430_n
  );


  buf

  (
    g430_p_spl_,
    g430_p
  );


  buf

  (
    g432_p_spl_,
    g432_p
  );


  buf

  (
    g371_n_spl_,
    g371_n
  );


  buf

  (
    g432_n_spl_,
    g432_n
  );


  buf

  (
    g371_p_spl_,
    g371_p
  );


  buf

  (
    g433_n_spl_,
    g433_n
  );


  buf

  (
    g433_p_spl_,
    g433_p
  );


  buf

  (
    g435_p_spl_,
    g435_p
  );


  buf

  (
    g370_n_spl_,
    g370_n
  );


  buf

  (
    g435_n_spl_,
    g435_n
  );


  buf

  (
    g370_p_spl_,
    g370_p
  );


  buf

  (
    g436_n_spl_,
    g436_n
  );


  buf

  (
    g436_p_spl_,
    g436_p
  );


  buf

  (
    g438_p_spl_,
    g438_p
  );


  buf

  (
    g369_n_spl_,
    g369_n
  );


  buf

  (
    g438_n_spl_,
    g438_n
  );


  buf

  (
    g369_p_spl_,
    g369_p
  );


  buf

  (
    g439_n_spl_,
    g439_n
  );


  buf

  (
    g439_p_spl_,
    g439_p
  );


  buf

  (
    g441_n_spl_,
    g441_n
  );


  buf

  (
    g368_p_spl_,
    g368_p
  );


  buf

  (
    g442_p_spl_,
    g442_p
  );


  buf

  (
    G28_p_spl_,
    G28_p
  );


  buf

  (
    G28_p_spl_0,
    G28_p_spl_
  );


  buf

  (
    G28_p_spl_00,
    G28_p_spl_0
  );


  buf

  (
    G28_p_spl_000,
    G28_p_spl_00
  );


  buf

  (
    G28_p_spl_001,
    G28_p_spl_00
  );


  buf

  (
    G28_p_spl_01,
    G28_p_spl_0
  );


  buf

  (
    G28_p_spl_010,
    G28_p_spl_01
  );


  buf

  (
    G28_p_spl_011,
    G28_p_spl_01
  );


  buf

  (
    G28_p_spl_1,
    G28_p_spl_
  );


  buf

  (
    G28_p_spl_10,
    G28_p_spl_1
  );


  buf

  (
    G28_p_spl_100,
    G28_p_spl_10
  );


  buf

  (
    G28_p_spl_101,
    G28_p_spl_10
  );


  buf

  (
    G28_p_spl_11,
    G28_p_spl_1
  );


  buf

  (
    G28_p_spl_110,
    G28_p_spl_11
  );


  buf

  (
    G28_p_spl_111,
    G28_p_spl_11
  );


  buf

  (
    G28_n_spl_,
    G28_n
  );


  buf

  (
    G28_n_spl_0,
    G28_n_spl_
  );


  buf

  (
    G28_n_spl_00,
    G28_n_spl_0
  );


  buf

  (
    G28_n_spl_000,
    G28_n_spl_00
  );


  buf

  (
    G28_n_spl_001,
    G28_n_spl_00
  );


  buf

  (
    G28_n_spl_01,
    G28_n_spl_0
  );


  buf

  (
    G28_n_spl_010,
    G28_n_spl_01
  );


  buf

  (
    G28_n_spl_011,
    G28_n_spl_01
  );


  buf

  (
    G28_n_spl_1,
    G28_n_spl_
  );


  buf

  (
    G28_n_spl_10,
    G28_n_spl_1
  );


  buf

  (
    G28_n_spl_100,
    G28_n_spl_10
  );


  buf

  (
    G28_n_spl_101,
    G28_n_spl_10
  );


  buf

  (
    G28_n_spl_11,
    G28_n_spl_1
  );


  buf

  (
    G28_n_spl_110,
    G28_n_spl_11
  );


  buf

  (
    G28_n_spl_111,
    G28_n_spl_11
  );


  buf

  (
    G12_p_spl_,
    G12_p
  );


  buf

  (
    G12_p_spl_0,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_00,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_000,
    G12_p_spl_00
  );


  buf

  (
    G12_p_spl_001,
    G12_p_spl_00
  );


  buf

  (
    G12_p_spl_01,
    G12_p_spl_0
  );


  buf

  (
    G12_p_spl_010,
    G12_p_spl_01
  );


  buf

  (
    G12_p_spl_011,
    G12_p_spl_01
  );


  buf

  (
    G12_p_spl_1,
    G12_p_spl_
  );


  buf

  (
    G12_p_spl_10,
    G12_p_spl_1
  );


  buf

  (
    G12_p_spl_100,
    G12_p_spl_10
  );


  buf

  (
    G12_p_spl_101,
    G12_p_spl_10
  );


  buf

  (
    G12_p_spl_11,
    G12_p_spl_1
  );


  buf

  (
    G12_p_spl_110,
    G12_p_spl_11
  );


  buf

  (
    G12_p_spl_111,
    G12_p_spl_11
  );


  buf

  (
    G12_n_spl_,
    G12_n
  );


  buf

  (
    G12_n_spl_0,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_00,
    G12_n_spl_0
  );


  buf

  (
    G12_n_spl_000,
    G12_n_spl_00
  );


  buf

  (
    G12_n_spl_001,
    G12_n_spl_00
  );


  buf

  (
    G12_n_spl_01,
    G12_n_spl_0
  );


  buf

  (
    G12_n_spl_010,
    G12_n_spl_01
  );


  buf

  (
    G12_n_spl_011,
    G12_n_spl_01
  );


  buf

  (
    G12_n_spl_1,
    G12_n_spl_
  );


  buf

  (
    G12_n_spl_10,
    G12_n_spl_1
  );


  buf

  (
    G12_n_spl_100,
    G12_n_spl_10
  );


  buf

  (
    G12_n_spl_101,
    G12_n_spl_10
  );


  buf

  (
    G12_n_spl_11,
    G12_n_spl_1
  );


  buf

  (
    G12_n_spl_110,
    G12_n_spl_11
  );


  buf

  (
    G12_n_spl_111,
    G12_n_spl_11
  );


  buf

  (
    g465_n_spl_,
    g465_n
  );


  buf

  (
    g464_p_spl_,
    g464_p
  );


  buf

  (
    g465_p_spl_,
    g465_p
  );


  buf

  (
    g464_n_spl_,
    g464_n
  );


  buf

  (
    g466_n_spl_,
    g466_n
  );


  buf

  (
    g466_p_spl_,
    g466_p
  );


  buf

  (
    g467_n_spl_,
    g467_n
  );


  buf

  (
    g467_n_spl_0,
    g467_n_spl_
  );


  buf

  (
    g467_p_spl_,
    g467_p
  );


  buf

  (
    g467_p_spl_0,
    g467_p_spl_
  );


  buf

  (
    g469_n_spl_,
    g469_n
  );


  buf

  (
    g469_p_spl_,
    g469_p
  );


  buf

  (
    g470_n_spl_,
    g470_n
  );


  buf

  (
    g470_p_spl_,
    g470_p
  );


  buf

  (
    g472_p_spl_,
    g472_p
  );


  buf

  (
    g463_n_spl_,
    g463_n
  );


  buf

  (
    g472_n_spl_,
    g472_n
  );


  buf

  (
    g463_p_spl_,
    g463_p
  );


  buf

  (
    g473_n_spl_,
    g473_n
  );


  buf

  (
    g473_p_spl_,
    g473_p
  );


  buf

  (
    g475_p_spl_,
    g475_p
  );


  buf

  (
    g462_n_spl_,
    g462_n
  );


  buf

  (
    g475_n_spl_,
    g475_n
  );


  buf

  (
    g462_p_spl_,
    g462_p
  );


  buf

  (
    g476_n_spl_,
    g476_n
  );


  buf

  (
    g476_p_spl_,
    g476_p
  );


  buf

  (
    g478_p_spl_,
    g478_p
  );


  buf

  (
    g461_n_spl_,
    g461_n
  );


  buf

  (
    g478_n_spl_,
    g478_n
  );


  buf

  (
    g461_p_spl_,
    g461_p
  );


  buf

  (
    g479_n_spl_,
    g479_n
  );


  buf

  (
    g479_p_spl_,
    g479_p
  );


  buf

  (
    g481_p_spl_,
    g481_p
  );


  buf

  (
    g460_n_spl_,
    g460_n
  );


  buf

  (
    g481_n_spl_,
    g481_n
  );


  buf

  (
    g460_p_spl_,
    g460_p
  );


  buf

  (
    g482_n_spl_,
    g482_n
  );


  buf

  (
    g482_p_spl_,
    g482_p
  );


  buf

  (
    g484_p_spl_,
    g484_p
  );


  buf

  (
    g459_n_spl_,
    g459_n
  );


  buf

  (
    g484_n_spl_,
    g484_n
  );


  buf

  (
    g459_p_spl_,
    g459_p
  );


  buf

  (
    g485_n_spl_,
    g485_n
  );


  buf

  (
    g485_p_spl_,
    g485_p
  );


  buf

  (
    g487_p_spl_,
    g487_p
  );


  buf

  (
    g458_n_spl_,
    g458_n
  );


  buf

  (
    g487_n_spl_,
    g487_n
  );


  buf

  (
    g458_p_spl_,
    g458_p
  );


  buf

  (
    g488_n_spl_,
    g488_n
  );


  buf

  (
    g488_p_spl_,
    g488_p
  );


  buf

  (
    g490_p_spl_,
    g490_p
  );


  buf

  (
    g457_n_spl_,
    g457_n
  );


  buf

  (
    g490_n_spl_,
    g490_n
  );


  buf

  (
    g457_p_spl_,
    g457_p
  );


  buf

  (
    g491_n_spl_,
    g491_n
  );


  buf

  (
    g491_p_spl_,
    g491_p
  );


  buf

  (
    g493_p_spl_,
    g493_p
  );


  buf

  (
    g456_n_spl_,
    g456_n
  );


  buf

  (
    g493_n_spl_,
    g493_n
  );


  buf

  (
    g456_p_spl_,
    g456_p
  );


  buf

  (
    g494_n_spl_,
    g494_n
  );


  buf

  (
    g494_p_spl_,
    g494_p
  );


  buf

  (
    g496_p_spl_,
    g496_p
  );


  buf

  (
    g455_n_spl_,
    g455_n
  );


  buf

  (
    g496_n_spl_,
    g496_n
  );


  buf

  (
    g455_p_spl_,
    g455_p
  );


  buf

  (
    g497_n_spl_,
    g497_n
  );


  buf

  (
    g497_p_spl_,
    g497_p
  );


  buf

  (
    g499_p_spl_,
    g499_p
  );


  buf

  (
    g454_n_spl_,
    g454_n
  );


  buf

  (
    g499_n_spl_,
    g499_n
  );


  buf

  (
    g454_p_spl_,
    g454_p
  );


  buf

  (
    g500_n_spl_,
    g500_n
  );


  buf

  (
    g500_p_spl_,
    g500_p
  );


  buf

  (
    g502_p_spl_,
    g502_p
  );


  buf

  (
    g453_n_spl_,
    g453_n
  );


  buf

  (
    g502_n_spl_,
    g502_n
  );


  buf

  (
    g453_p_spl_,
    g453_p
  );


  buf

  (
    g503_n_spl_,
    g503_n
  );


  buf

  (
    g503_p_spl_,
    g503_p
  );


  buf

  (
    g505_p_spl_,
    g505_p
  );


  buf

  (
    g452_n_spl_,
    g452_n
  );


  buf

  (
    g505_n_spl_,
    g505_n
  );


  buf

  (
    g452_p_spl_,
    g452_p
  );


  buf

  (
    g506_n_spl_,
    g506_n
  );


  buf

  (
    g506_p_spl_,
    g506_p
  );


  buf

  (
    g508_p_spl_,
    g508_p
  );


  buf

  (
    g451_n_spl_,
    g451_n
  );


  buf

  (
    g508_n_spl_,
    g508_n
  );


  buf

  (
    g451_p_spl_,
    g451_p
  );


  buf

  (
    g509_n_spl_,
    g509_n
  );


  buf

  (
    g509_p_spl_,
    g509_p
  );


  buf

  (
    g511_p_spl_,
    g511_p
  );


  buf

  (
    g450_n_spl_,
    g450_n
  );


  buf

  (
    g511_n_spl_,
    g511_n
  );


  buf

  (
    g450_p_spl_,
    g450_p
  );


  buf

  (
    g512_n_spl_,
    g512_n
  );


  buf

  (
    g512_p_spl_,
    g512_p
  );


  buf

  (
    g514_p_spl_,
    g514_p
  );


  buf

  (
    g449_n_spl_,
    g449_n
  );


  buf

  (
    g514_n_spl_,
    g514_n
  );


  buf

  (
    g449_p_spl_,
    g449_p
  );


  buf

  (
    g515_n_spl_,
    g515_n
  );


  buf

  (
    g515_p_spl_,
    g515_p
  );


  buf

  (
    g517_p_spl_,
    g517_p
  );


  buf

  (
    g448_n_spl_,
    g448_n
  );


  buf

  (
    g517_n_spl_,
    g517_n
  );


  buf

  (
    g448_p_spl_,
    g448_p
  );


  buf

  (
    g518_n_spl_,
    g518_n
  );


  buf

  (
    g518_p_spl_,
    g518_p
  );


  buf

  (
    g520_p_spl_,
    g520_p
  );


  buf

  (
    g447_n_spl_,
    g447_n
  );


  buf

  (
    g520_n_spl_,
    g520_n
  );


  buf

  (
    g447_p_spl_,
    g447_p
  );


  buf

  (
    g521_n_spl_,
    g521_n
  );


  buf

  (
    g521_p_spl_,
    g521_p
  );


  buf

  (
    g523_p_spl_,
    g523_p
  );


  buf

  (
    g446_n_spl_,
    g446_n
  );


  buf

  (
    g523_n_spl_,
    g523_n
  );


  buf

  (
    g446_p_spl_,
    g446_p
  );


  buf

  (
    g524_n_spl_,
    g524_n
  );


  buf

  (
    g524_p_spl_,
    g524_p
  );


  buf

  (
    g526_n_spl_,
    g526_n
  );


  buf

  (
    g445_p_spl_,
    g445_p
  );


  buf

  (
    g527_p_spl_,
    g527_p
  );


  buf

  (
    G29_p_spl_,
    G29_p
  );


  buf

  (
    G29_p_spl_0,
    G29_p_spl_
  );


  buf

  (
    G29_p_spl_00,
    G29_p_spl_0
  );


  buf

  (
    G29_p_spl_000,
    G29_p_spl_00
  );


  buf

  (
    G29_p_spl_001,
    G29_p_spl_00
  );


  buf

  (
    G29_p_spl_01,
    G29_p_spl_0
  );


  buf

  (
    G29_p_spl_010,
    G29_p_spl_01
  );


  buf

  (
    G29_p_spl_011,
    G29_p_spl_01
  );


  buf

  (
    G29_p_spl_1,
    G29_p_spl_
  );


  buf

  (
    G29_p_spl_10,
    G29_p_spl_1
  );


  buf

  (
    G29_p_spl_100,
    G29_p_spl_10
  );


  buf

  (
    G29_p_spl_101,
    G29_p_spl_10
  );


  buf

  (
    G29_p_spl_11,
    G29_p_spl_1
  );


  buf

  (
    G29_p_spl_110,
    G29_p_spl_11
  );


  buf

  (
    G29_p_spl_111,
    G29_p_spl_11
  );


  buf

  (
    G29_n_spl_,
    G29_n
  );


  buf

  (
    G29_n_spl_0,
    G29_n_spl_
  );


  buf

  (
    G29_n_spl_00,
    G29_n_spl_0
  );


  buf

  (
    G29_n_spl_000,
    G29_n_spl_00
  );


  buf

  (
    G29_n_spl_001,
    G29_n_spl_00
  );


  buf

  (
    G29_n_spl_01,
    G29_n_spl_0
  );


  buf

  (
    G29_n_spl_010,
    G29_n_spl_01
  );


  buf

  (
    G29_n_spl_011,
    G29_n_spl_01
  );


  buf

  (
    G29_n_spl_1,
    G29_n_spl_
  );


  buf

  (
    G29_n_spl_10,
    G29_n_spl_1
  );


  buf

  (
    G29_n_spl_100,
    G29_n_spl_10
  );


  buf

  (
    G29_n_spl_101,
    G29_n_spl_10
  );


  buf

  (
    G29_n_spl_11,
    G29_n_spl_1
  );


  buf

  (
    G29_n_spl_110,
    G29_n_spl_11
  );


  buf

  (
    G29_n_spl_111,
    G29_n_spl_11
  );


  buf

  (
    G13_p_spl_,
    G13_p
  );


  buf

  (
    G13_p_spl_0,
    G13_p_spl_
  );


  buf

  (
    G13_p_spl_00,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_000,
    G13_p_spl_00
  );


  buf

  (
    G13_p_spl_001,
    G13_p_spl_00
  );


  buf

  (
    G13_p_spl_01,
    G13_p_spl_0
  );


  buf

  (
    G13_p_spl_010,
    G13_p_spl_01
  );


  buf

  (
    G13_p_spl_011,
    G13_p_spl_01
  );


  buf

  (
    G13_p_spl_1,
    G13_p_spl_
  );


  buf

  (
    G13_p_spl_10,
    G13_p_spl_1
  );


  buf

  (
    G13_p_spl_100,
    G13_p_spl_10
  );


  buf

  (
    G13_p_spl_101,
    G13_p_spl_10
  );


  buf

  (
    G13_p_spl_11,
    G13_p_spl_1
  );


  buf

  (
    G13_p_spl_110,
    G13_p_spl_11
  );


  buf

  (
    G13_p_spl_111,
    G13_p_spl_11
  );


  buf

  (
    G13_n_spl_,
    G13_n
  );


  buf

  (
    G13_n_spl_0,
    G13_n_spl_
  );


  buf

  (
    G13_n_spl_00,
    G13_n_spl_0
  );


  buf

  (
    G13_n_spl_000,
    G13_n_spl_00
  );


  buf

  (
    G13_n_spl_001,
    G13_n_spl_00
  );


  buf

  (
    G13_n_spl_01,
    G13_n_spl_0
  );


  buf

  (
    G13_n_spl_010,
    G13_n_spl_01
  );


  buf

  (
    G13_n_spl_011,
    G13_n_spl_01
  );


  buf

  (
    G13_n_spl_1,
    G13_n_spl_
  );


  buf

  (
    G13_n_spl_10,
    G13_n_spl_1
  );


  buf

  (
    G13_n_spl_100,
    G13_n_spl_10
  );


  buf

  (
    G13_n_spl_101,
    G13_n_spl_10
  );


  buf

  (
    G13_n_spl_11,
    G13_n_spl_1
  );


  buf

  (
    G13_n_spl_110,
    G13_n_spl_11
  );


  buf

  (
    G13_n_spl_111,
    G13_n_spl_11
  );


  buf

  (
    g552_n_spl_,
    g552_n
  );


  buf

  (
    g551_p_spl_,
    g551_p
  );


  buf

  (
    g552_p_spl_,
    g552_p
  );


  buf

  (
    g551_n_spl_,
    g551_n
  );


  buf

  (
    g553_n_spl_,
    g553_n
  );


  buf

  (
    g553_p_spl_,
    g553_p
  );


  buf

  (
    g554_n_spl_,
    g554_n
  );


  buf

  (
    g554_n_spl_0,
    g554_n_spl_
  );


  buf

  (
    g554_p_spl_,
    g554_p
  );


  buf

  (
    g554_p_spl_0,
    g554_p_spl_
  );


  buf

  (
    g556_n_spl_,
    g556_n
  );


  buf

  (
    g556_p_spl_,
    g556_p
  );


  buf

  (
    g557_n_spl_,
    g557_n
  );


  buf

  (
    g557_p_spl_,
    g557_p
  );


  buf

  (
    g559_p_spl_,
    g559_p
  );


  buf

  (
    g550_n_spl_,
    g550_n
  );


  buf

  (
    g559_n_spl_,
    g559_n
  );


  buf

  (
    g550_p_spl_,
    g550_p
  );


  buf

  (
    g560_n_spl_,
    g560_n
  );


  buf

  (
    g560_p_spl_,
    g560_p
  );


  buf

  (
    g562_p_spl_,
    g562_p
  );


  buf

  (
    g549_n_spl_,
    g549_n
  );


  buf

  (
    g562_n_spl_,
    g562_n
  );


  buf

  (
    g549_p_spl_,
    g549_p
  );


  buf

  (
    g563_n_spl_,
    g563_n
  );


  buf

  (
    g563_p_spl_,
    g563_p
  );


  buf

  (
    g565_p_spl_,
    g565_p
  );


  buf

  (
    g548_n_spl_,
    g548_n
  );


  buf

  (
    g565_n_spl_,
    g565_n
  );


  buf

  (
    g548_p_spl_,
    g548_p
  );


  buf

  (
    g566_n_spl_,
    g566_n
  );


  buf

  (
    g566_p_spl_,
    g566_p
  );


  buf

  (
    g568_p_spl_,
    g568_p
  );


  buf

  (
    g547_n_spl_,
    g547_n
  );


  buf

  (
    g568_n_spl_,
    g568_n
  );


  buf

  (
    g547_p_spl_,
    g547_p
  );


  buf

  (
    g569_n_spl_,
    g569_n
  );


  buf

  (
    g569_p_spl_,
    g569_p
  );


  buf

  (
    g571_p_spl_,
    g571_p
  );


  buf

  (
    g546_n_spl_,
    g546_n
  );


  buf

  (
    g571_n_spl_,
    g571_n
  );


  buf

  (
    g546_p_spl_,
    g546_p
  );


  buf

  (
    g572_n_spl_,
    g572_n
  );


  buf

  (
    g572_p_spl_,
    g572_p
  );


  buf

  (
    g574_p_spl_,
    g574_p
  );


  buf

  (
    g545_n_spl_,
    g545_n
  );


  buf

  (
    g574_n_spl_,
    g574_n
  );


  buf

  (
    g545_p_spl_,
    g545_p
  );


  buf

  (
    g575_n_spl_,
    g575_n
  );


  buf

  (
    g575_p_spl_,
    g575_p
  );


  buf

  (
    g577_p_spl_,
    g577_p
  );


  buf

  (
    g544_n_spl_,
    g544_n
  );


  buf

  (
    g577_n_spl_,
    g577_n
  );


  buf

  (
    g544_p_spl_,
    g544_p
  );


  buf

  (
    g578_n_spl_,
    g578_n
  );


  buf

  (
    g578_p_spl_,
    g578_p
  );


  buf

  (
    g580_p_spl_,
    g580_p
  );


  buf

  (
    g543_n_spl_,
    g543_n
  );


  buf

  (
    g580_n_spl_,
    g580_n
  );


  buf

  (
    g543_p_spl_,
    g543_p
  );


  buf

  (
    g581_n_spl_,
    g581_n
  );


  buf

  (
    g581_p_spl_,
    g581_p
  );


  buf

  (
    g583_p_spl_,
    g583_p
  );


  buf

  (
    g542_n_spl_,
    g542_n
  );


  buf

  (
    g583_n_spl_,
    g583_n
  );


  buf

  (
    g542_p_spl_,
    g542_p
  );


  buf

  (
    g584_n_spl_,
    g584_n
  );


  buf

  (
    g584_p_spl_,
    g584_p
  );


  buf

  (
    g586_p_spl_,
    g586_p
  );


  buf

  (
    g541_n_spl_,
    g541_n
  );


  buf

  (
    g586_n_spl_,
    g586_n
  );


  buf

  (
    g541_p_spl_,
    g541_p
  );


  buf

  (
    g587_n_spl_,
    g587_n
  );


  buf

  (
    g587_p_spl_,
    g587_p
  );


  buf

  (
    g589_p_spl_,
    g589_p
  );


  buf

  (
    g540_n_spl_,
    g540_n
  );


  buf

  (
    g589_n_spl_,
    g589_n
  );


  buf

  (
    g540_p_spl_,
    g540_p
  );


  buf

  (
    g590_n_spl_,
    g590_n
  );


  buf

  (
    g590_p_spl_,
    g590_p
  );


  buf

  (
    g592_p_spl_,
    g592_p
  );


  buf

  (
    g539_n_spl_,
    g539_n
  );


  buf

  (
    g592_n_spl_,
    g592_n
  );


  buf

  (
    g539_p_spl_,
    g539_p
  );


  buf

  (
    g593_n_spl_,
    g593_n
  );


  buf

  (
    g593_p_spl_,
    g593_p
  );


  buf

  (
    g595_p_spl_,
    g595_p
  );


  buf

  (
    g538_n_spl_,
    g538_n
  );


  buf

  (
    g595_n_spl_,
    g595_n
  );


  buf

  (
    g538_p_spl_,
    g538_p
  );


  buf

  (
    g596_n_spl_,
    g596_n
  );


  buf

  (
    g596_p_spl_,
    g596_p
  );


  buf

  (
    g598_p_spl_,
    g598_p
  );


  buf

  (
    g537_n_spl_,
    g537_n
  );


  buf

  (
    g598_n_spl_,
    g598_n
  );


  buf

  (
    g537_p_spl_,
    g537_p
  );


  buf

  (
    g599_n_spl_,
    g599_n
  );


  buf

  (
    g599_p_spl_,
    g599_p
  );


  buf

  (
    g601_p_spl_,
    g601_p
  );


  buf

  (
    g536_n_spl_,
    g536_n
  );


  buf

  (
    g601_n_spl_,
    g601_n
  );


  buf

  (
    g536_p_spl_,
    g536_p
  );


  buf

  (
    g602_n_spl_,
    g602_n
  );


  buf

  (
    g602_p_spl_,
    g602_p
  );


  buf

  (
    g604_p_spl_,
    g604_p
  );


  buf

  (
    g535_n_spl_,
    g535_n
  );


  buf

  (
    g604_n_spl_,
    g604_n
  );


  buf

  (
    g535_p_spl_,
    g535_p
  );


  buf

  (
    g605_n_spl_,
    g605_n
  );


  buf

  (
    g605_p_spl_,
    g605_p
  );


  buf

  (
    g607_p_spl_,
    g607_p
  );


  buf

  (
    g534_n_spl_,
    g534_n
  );


  buf

  (
    g607_n_spl_,
    g607_n
  );


  buf

  (
    g534_p_spl_,
    g534_p
  );


  buf

  (
    g608_n_spl_,
    g608_n
  );


  buf

  (
    g608_p_spl_,
    g608_p
  );


  buf

  (
    g610_p_spl_,
    g610_p
  );


  buf

  (
    g533_n_spl_,
    g533_n
  );


  buf

  (
    g610_n_spl_,
    g610_n
  );


  buf

  (
    g533_p_spl_,
    g533_p
  );


  buf

  (
    g611_n_spl_,
    g611_n
  );


  buf

  (
    g611_p_spl_,
    g611_p
  );


  buf

  (
    g613_p_spl_,
    g613_p
  );


  buf

  (
    g532_n_spl_,
    g532_n
  );


  buf

  (
    g613_n_spl_,
    g613_n
  );


  buf

  (
    g532_p_spl_,
    g532_p
  );


  buf

  (
    g614_n_spl_,
    g614_n
  );


  buf

  (
    g614_p_spl_,
    g614_p
  );


  buf

  (
    g616_p_spl_,
    g616_p
  );


  buf

  (
    g531_n_spl_,
    g531_n
  );


  buf

  (
    g616_n_spl_,
    g616_n
  );


  buf

  (
    g531_p_spl_,
    g531_p
  );


  buf

  (
    g617_n_spl_,
    g617_n
  );


  buf

  (
    g617_p_spl_,
    g617_p
  );


  buf

  (
    g619_n_spl_,
    g619_n
  );


  buf

  (
    g530_p_spl_,
    g530_p
  );


  buf

  (
    g620_p_spl_,
    g620_p
  );


  buf

  (
    G30_p_spl_,
    G30_p
  );


  buf

  (
    G30_p_spl_0,
    G30_p_spl_
  );


  buf

  (
    G30_p_spl_00,
    G30_p_spl_0
  );


  buf

  (
    G30_p_spl_000,
    G30_p_spl_00
  );


  buf

  (
    G30_p_spl_001,
    G30_p_spl_00
  );


  buf

  (
    G30_p_spl_01,
    G30_p_spl_0
  );


  buf

  (
    G30_p_spl_010,
    G30_p_spl_01
  );


  buf

  (
    G30_p_spl_011,
    G30_p_spl_01
  );


  buf

  (
    G30_p_spl_1,
    G30_p_spl_
  );


  buf

  (
    G30_p_spl_10,
    G30_p_spl_1
  );


  buf

  (
    G30_p_spl_100,
    G30_p_spl_10
  );


  buf

  (
    G30_p_spl_101,
    G30_p_spl_10
  );


  buf

  (
    G30_p_spl_11,
    G30_p_spl_1
  );


  buf

  (
    G30_p_spl_110,
    G30_p_spl_11
  );


  buf

  (
    G30_p_spl_111,
    G30_p_spl_11
  );


  buf

  (
    G30_n_spl_,
    G30_n
  );


  buf

  (
    G30_n_spl_0,
    G30_n_spl_
  );


  buf

  (
    G30_n_spl_00,
    G30_n_spl_0
  );


  buf

  (
    G30_n_spl_000,
    G30_n_spl_00
  );


  buf

  (
    G30_n_spl_001,
    G30_n_spl_00
  );


  buf

  (
    G30_n_spl_01,
    G30_n_spl_0
  );


  buf

  (
    G30_n_spl_010,
    G30_n_spl_01
  );


  buf

  (
    G30_n_spl_011,
    G30_n_spl_01
  );


  buf

  (
    G30_n_spl_1,
    G30_n_spl_
  );


  buf

  (
    G30_n_spl_10,
    G30_n_spl_1
  );


  buf

  (
    G30_n_spl_100,
    G30_n_spl_10
  );


  buf

  (
    G30_n_spl_101,
    G30_n_spl_10
  );


  buf

  (
    G30_n_spl_11,
    G30_n_spl_1
  );


  buf

  (
    G30_n_spl_110,
    G30_n_spl_11
  );


  buf

  (
    G30_n_spl_111,
    G30_n_spl_11
  );


  buf

  (
    G14_p_spl_,
    G14_p
  );


  buf

  (
    G14_p_spl_0,
    G14_p_spl_
  );


  buf

  (
    G14_p_spl_00,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_000,
    G14_p_spl_00
  );


  buf

  (
    G14_p_spl_001,
    G14_p_spl_00
  );


  buf

  (
    G14_p_spl_01,
    G14_p_spl_0
  );


  buf

  (
    G14_p_spl_010,
    G14_p_spl_01
  );


  buf

  (
    G14_p_spl_011,
    G14_p_spl_01
  );


  buf

  (
    G14_p_spl_1,
    G14_p_spl_
  );


  buf

  (
    G14_p_spl_10,
    G14_p_spl_1
  );


  buf

  (
    G14_p_spl_100,
    G14_p_spl_10
  );


  buf

  (
    G14_p_spl_101,
    G14_p_spl_10
  );


  buf

  (
    G14_p_spl_11,
    G14_p_spl_1
  );


  buf

  (
    G14_p_spl_110,
    G14_p_spl_11
  );


  buf

  (
    G14_p_spl_111,
    G14_p_spl_11
  );


  buf

  (
    G14_n_spl_,
    G14_n
  );


  buf

  (
    G14_n_spl_0,
    G14_n_spl_
  );


  buf

  (
    G14_n_spl_00,
    G14_n_spl_0
  );


  buf

  (
    G14_n_spl_000,
    G14_n_spl_00
  );


  buf

  (
    G14_n_spl_001,
    G14_n_spl_00
  );


  buf

  (
    G14_n_spl_01,
    G14_n_spl_0
  );


  buf

  (
    G14_n_spl_010,
    G14_n_spl_01
  );


  buf

  (
    G14_n_spl_011,
    G14_n_spl_01
  );


  buf

  (
    G14_n_spl_1,
    G14_n_spl_
  );


  buf

  (
    G14_n_spl_10,
    G14_n_spl_1
  );


  buf

  (
    G14_n_spl_100,
    G14_n_spl_10
  );


  buf

  (
    G14_n_spl_101,
    G14_n_spl_10
  );


  buf

  (
    G14_n_spl_11,
    G14_n_spl_1
  );


  buf

  (
    G14_n_spl_110,
    G14_n_spl_11
  );


  buf

  (
    G14_n_spl_111,
    G14_n_spl_11
  );


  buf

  (
    g647_n_spl_,
    g647_n
  );


  buf

  (
    g646_p_spl_,
    g646_p
  );


  buf

  (
    g647_p_spl_,
    g647_p
  );


  buf

  (
    g646_n_spl_,
    g646_n
  );


  buf

  (
    g648_n_spl_,
    g648_n
  );


  buf

  (
    g648_p_spl_,
    g648_p
  );


  buf

  (
    g649_n_spl_,
    g649_n
  );


  buf

  (
    g649_n_spl_0,
    g649_n_spl_
  );


  buf

  (
    g649_p_spl_,
    g649_p
  );


  buf

  (
    g649_p_spl_0,
    g649_p_spl_
  );


  buf

  (
    g651_n_spl_,
    g651_n
  );


  buf

  (
    g651_p_spl_,
    g651_p
  );


  buf

  (
    g652_n_spl_,
    g652_n
  );


  buf

  (
    g652_p_spl_,
    g652_p
  );


  buf

  (
    g654_p_spl_,
    g654_p
  );


  buf

  (
    g645_n_spl_,
    g645_n
  );


  buf

  (
    g654_n_spl_,
    g654_n
  );


  buf

  (
    g645_p_spl_,
    g645_p
  );


  buf

  (
    g655_n_spl_,
    g655_n
  );


  buf

  (
    g655_p_spl_,
    g655_p
  );


  buf

  (
    g657_p_spl_,
    g657_p
  );


  buf

  (
    g644_n_spl_,
    g644_n
  );


  buf

  (
    g657_n_spl_,
    g657_n
  );


  buf

  (
    g644_p_spl_,
    g644_p
  );


  buf

  (
    g658_n_spl_,
    g658_n
  );


  buf

  (
    g658_p_spl_,
    g658_p
  );


  buf

  (
    g660_p_spl_,
    g660_p
  );


  buf

  (
    g643_n_spl_,
    g643_n
  );


  buf

  (
    g660_n_spl_,
    g660_n
  );


  buf

  (
    g643_p_spl_,
    g643_p
  );


  buf

  (
    g661_n_spl_,
    g661_n
  );


  buf

  (
    g661_p_spl_,
    g661_p
  );


  buf

  (
    g663_p_spl_,
    g663_p
  );


  buf

  (
    g642_n_spl_,
    g642_n
  );


  buf

  (
    g663_n_spl_,
    g663_n
  );


  buf

  (
    g642_p_spl_,
    g642_p
  );


  buf

  (
    g664_n_spl_,
    g664_n
  );


  buf

  (
    g664_p_spl_,
    g664_p
  );


  buf

  (
    g666_p_spl_,
    g666_p
  );


  buf

  (
    g641_n_spl_,
    g641_n
  );


  buf

  (
    g666_n_spl_,
    g666_n
  );


  buf

  (
    g641_p_spl_,
    g641_p
  );


  buf

  (
    g667_n_spl_,
    g667_n
  );


  buf

  (
    g667_p_spl_,
    g667_p
  );


  buf

  (
    g669_p_spl_,
    g669_p
  );


  buf

  (
    g640_n_spl_,
    g640_n
  );


  buf

  (
    g669_n_spl_,
    g669_n
  );


  buf

  (
    g640_p_spl_,
    g640_p
  );


  buf

  (
    g670_n_spl_,
    g670_n
  );


  buf

  (
    g670_p_spl_,
    g670_p
  );


  buf

  (
    g672_p_spl_,
    g672_p
  );


  buf

  (
    g639_n_spl_,
    g639_n
  );


  buf

  (
    g672_n_spl_,
    g672_n
  );


  buf

  (
    g639_p_spl_,
    g639_p
  );


  buf

  (
    g673_n_spl_,
    g673_n
  );


  buf

  (
    g673_p_spl_,
    g673_p
  );


  buf

  (
    g675_p_spl_,
    g675_p
  );


  buf

  (
    g638_n_spl_,
    g638_n
  );


  buf

  (
    g675_n_spl_,
    g675_n
  );


  buf

  (
    g638_p_spl_,
    g638_p
  );


  buf

  (
    g676_n_spl_,
    g676_n
  );


  buf

  (
    g676_p_spl_,
    g676_p
  );


  buf

  (
    g678_p_spl_,
    g678_p
  );


  buf

  (
    g637_n_spl_,
    g637_n
  );


  buf

  (
    g678_n_spl_,
    g678_n
  );


  buf

  (
    g637_p_spl_,
    g637_p
  );


  buf

  (
    g679_n_spl_,
    g679_n
  );


  buf

  (
    g679_p_spl_,
    g679_p
  );


  buf

  (
    g681_p_spl_,
    g681_p
  );


  buf

  (
    g636_n_spl_,
    g636_n
  );


  buf

  (
    g681_n_spl_,
    g681_n
  );


  buf

  (
    g636_p_spl_,
    g636_p
  );


  buf

  (
    g682_n_spl_,
    g682_n
  );


  buf

  (
    g682_p_spl_,
    g682_p
  );


  buf

  (
    g684_p_spl_,
    g684_p
  );


  buf

  (
    g635_n_spl_,
    g635_n
  );


  buf

  (
    g684_n_spl_,
    g684_n
  );


  buf

  (
    g635_p_spl_,
    g635_p
  );


  buf

  (
    g685_n_spl_,
    g685_n
  );


  buf

  (
    g685_p_spl_,
    g685_p
  );


  buf

  (
    g687_p_spl_,
    g687_p
  );


  buf

  (
    g634_n_spl_,
    g634_n
  );


  buf

  (
    g687_n_spl_,
    g687_n
  );


  buf

  (
    g634_p_spl_,
    g634_p
  );


  buf

  (
    g688_n_spl_,
    g688_n
  );


  buf

  (
    g688_p_spl_,
    g688_p
  );


  buf

  (
    g690_p_spl_,
    g690_p
  );


  buf

  (
    g633_n_spl_,
    g633_n
  );


  buf

  (
    g690_n_spl_,
    g690_n
  );


  buf

  (
    g633_p_spl_,
    g633_p
  );


  buf

  (
    g691_n_spl_,
    g691_n
  );


  buf

  (
    g691_p_spl_,
    g691_p
  );


  buf

  (
    g693_p_spl_,
    g693_p
  );


  buf

  (
    g632_n_spl_,
    g632_n
  );


  buf

  (
    g693_n_spl_,
    g693_n
  );


  buf

  (
    g632_p_spl_,
    g632_p
  );


  buf

  (
    g694_n_spl_,
    g694_n
  );


  buf

  (
    g694_p_spl_,
    g694_p
  );


  buf

  (
    g696_p_spl_,
    g696_p
  );


  buf

  (
    g631_n_spl_,
    g631_n
  );


  buf

  (
    g696_n_spl_,
    g696_n
  );


  buf

  (
    g631_p_spl_,
    g631_p
  );


  buf

  (
    g697_n_spl_,
    g697_n
  );


  buf

  (
    g697_p_spl_,
    g697_p
  );


  buf

  (
    g699_p_spl_,
    g699_p
  );


  buf

  (
    g630_n_spl_,
    g630_n
  );


  buf

  (
    g699_n_spl_,
    g699_n
  );


  buf

  (
    g630_p_spl_,
    g630_p
  );


  buf

  (
    g700_n_spl_,
    g700_n
  );


  buf

  (
    g700_p_spl_,
    g700_p
  );


  buf

  (
    g702_p_spl_,
    g702_p
  );


  buf

  (
    g629_n_spl_,
    g629_n
  );


  buf

  (
    g702_n_spl_,
    g702_n
  );


  buf

  (
    g629_p_spl_,
    g629_p
  );


  buf

  (
    g703_n_spl_,
    g703_n
  );


  buf

  (
    g703_p_spl_,
    g703_p
  );


  buf

  (
    g705_p_spl_,
    g705_p
  );


  buf

  (
    g628_n_spl_,
    g628_n
  );


  buf

  (
    g705_n_spl_,
    g705_n
  );


  buf

  (
    g628_p_spl_,
    g628_p
  );


  buf

  (
    g706_n_spl_,
    g706_n
  );


  buf

  (
    g706_p_spl_,
    g706_p
  );


  buf

  (
    g708_p_spl_,
    g708_p
  );


  buf

  (
    g627_n_spl_,
    g627_n
  );


  buf

  (
    g708_n_spl_,
    g708_n
  );


  buf

  (
    g627_p_spl_,
    g627_p
  );


  buf

  (
    g709_n_spl_,
    g709_n
  );


  buf

  (
    g709_p_spl_,
    g709_p
  );


  buf

  (
    g711_p_spl_,
    g711_p
  );


  buf

  (
    g626_n_spl_,
    g626_n
  );


  buf

  (
    g711_n_spl_,
    g711_n
  );


  buf

  (
    g626_p_spl_,
    g626_p
  );


  buf

  (
    g712_n_spl_,
    g712_n
  );


  buf

  (
    g712_p_spl_,
    g712_p
  );


  buf

  (
    g714_p_spl_,
    g714_p
  );


  buf

  (
    g625_n_spl_,
    g625_n
  );


  buf

  (
    g714_n_spl_,
    g714_n
  );


  buf

  (
    g625_p_spl_,
    g625_p
  );


  buf

  (
    g715_n_spl_,
    g715_n
  );


  buf

  (
    g715_p_spl_,
    g715_p
  );


  buf

  (
    g717_p_spl_,
    g717_p
  );


  buf

  (
    g624_n_spl_,
    g624_n
  );


  buf

  (
    g717_n_spl_,
    g717_n
  );


  buf

  (
    g624_p_spl_,
    g624_p
  );


  buf

  (
    g718_n_spl_,
    g718_n
  );


  buf

  (
    g718_p_spl_,
    g718_p
  );


  buf

  (
    g720_n_spl_,
    g720_n
  );


  buf

  (
    g623_p_spl_,
    g623_p
  );


  buf

  (
    g721_p_spl_,
    g721_p
  );


  buf

  (
    G31_p_spl_,
    G31_p
  );


  buf

  (
    G31_p_spl_0,
    G31_p_spl_
  );


  buf

  (
    G31_p_spl_00,
    G31_p_spl_0
  );


  buf

  (
    G31_p_spl_000,
    G31_p_spl_00
  );


  buf

  (
    G31_p_spl_001,
    G31_p_spl_00
  );


  buf

  (
    G31_p_spl_01,
    G31_p_spl_0
  );


  buf

  (
    G31_p_spl_010,
    G31_p_spl_01
  );


  buf

  (
    G31_p_spl_011,
    G31_p_spl_01
  );


  buf

  (
    G31_p_spl_1,
    G31_p_spl_
  );


  buf

  (
    G31_p_spl_10,
    G31_p_spl_1
  );


  buf

  (
    G31_p_spl_100,
    G31_p_spl_10
  );


  buf

  (
    G31_p_spl_101,
    G31_p_spl_10
  );


  buf

  (
    G31_p_spl_11,
    G31_p_spl_1
  );


  buf

  (
    G31_p_spl_110,
    G31_p_spl_11
  );


  buf

  (
    G31_p_spl_111,
    G31_p_spl_11
  );


  buf

  (
    G31_n_spl_,
    G31_n
  );


  buf

  (
    G31_n_spl_0,
    G31_n_spl_
  );


  buf

  (
    G31_n_spl_00,
    G31_n_spl_0
  );


  buf

  (
    G31_n_spl_000,
    G31_n_spl_00
  );


  buf

  (
    G31_n_spl_001,
    G31_n_spl_00
  );


  buf

  (
    G31_n_spl_01,
    G31_n_spl_0
  );


  buf

  (
    G31_n_spl_010,
    G31_n_spl_01
  );


  buf

  (
    G31_n_spl_011,
    G31_n_spl_01
  );


  buf

  (
    G31_n_spl_1,
    G31_n_spl_
  );


  buf

  (
    G31_n_spl_10,
    G31_n_spl_1
  );


  buf

  (
    G31_n_spl_100,
    G31_n_spl_10
  );


  buf

  (
    G31_n_spl_101,
    G31_n_spl_10
  );


  buf

  (
    G31_n_spl_11,
    G31_n_spl_1
  );


  buf

  (
    G31_n_spl_110,
    G31_n_spl_11
  );


  buf

  (
    G31_n_spl_111,
    G31_n_spl_11
  );


  buf

  (
    G15_p_spl_,
    G15_p
  );


  buf

  (
    G15_p_spl_0,
    G15_p_spl_
  );


  buf

  (
    G15_p_spl_00,
    G15_p_spl_0
  );


  buf

  (
    G15_p_spl_000,
    G15_p_spl_00
  );


  buf

  (
    G15_p_spl_001,
    G15_p_spl_00
  );


  buf

  (
    G15_p_spl_01,
    G15_p_spl_0
  );


  buf

  (
    G15_p_spl_010,
    G15_p_spl_01
  );


  buf

  (
    G15_p_spl_011,
    G15_p_spl_01
  );


  buf

  (
    G15_p_spl_1,
    G15_p_spl_
  );


  buf

  (
    G15_p_spl_10,
    G15_p_spl_1
  );


  buf

  (
    G15_p_spl_100,
    G15_p_spl_10
  );


  buf

  (
    G15_p_spl_101,
    G15_p_spl_10
  );


  buf

  (
    G15_p_spl_11,
    G15_p_spl_1
  );


  buf

  (
    G15_p_spl_110,
    G15_p_spl_11
  );


  buf

  (
    G15_p_spl_111,
    G15_p_spl_11
  );


  buf

  (
    G15_n_spl_,
    G15_n
  );


  buf

  (
    G15_n_spl_0,
    G15_n_spl_
  );


  buf

  (
    G15_n_spl_00,
    G15_n_spl_0
  );


  buf

  (
    G15_n_spl_000,
    G15_n_spl_00
  );


  buf

  (
    G15_n_spl_001,
    G15_n_spl_00
  );


  buf

  (
    G15_n_spl_01,
    G15_n_spl_0
  );


  buf

  (
    G15_n_spl_010,
    G15_n_spl_01
  );


  buf

  (
    G15_n_spl_011,
    G15_n_spl_01
  );


  buf

  (
    G15_n_spl_1,
    G15_n_spl_
  );


  buf

  (
    G15_n_spl_10,
    G15_n_spl_1
  );


  buf

  (
    G15_n_spl_100,
    G15_n_spl_10
  );


  buf

  (
    G15_n_spl_101,
    G15_n_spl_10
  );


  buf

  (
    G15_n_spl_11,
    G15_n_spl_1
  );


  buf

  (
    G15_n_spl_110,
    G15_n_spl_11
  );


  buf

  (
    G15_n_spl_111,
    G15_n_spl_11
  );


  buf

  (
    g750_n_spl_,
    g750_n
  );


  buf

  (
    g749_p_spl_,
    g749_p
  );


  buf

  (
    g750_p_spl_,
    g750_p
  );


  buf

  (
    g749_n_spl_,
    g749_n
  );


  buf

  (
    g751_n_spl_,
    g751_n
  );


  buf

  (
    g751_p_spl_,
    g751_p
  );


  buf

  (
    g752_n_spl_,
    g752_n
  );


  buf

  (
    g752_n_spl_0,
    g752_n_spl_
  );


  buf

  (
    g752_p_spl_,
    g752_p
  );


  buf

  (
    g752_p_spl_0,
    g752_p_spl_
  );


  buf

  (
    g754_n_spl_,
    g754_n
  );


  buf

  (
    g754_p_spl_,
    g754_p
  );


  buf

  (
    g755_n_spl_,
    g755_n
  );


  buf

  (
    g755_p_spl_,
    g755_p
  );


  buf

  (
    g757_p_spl_,
    g757_p
  );


  buf

  (
    g748_n_spl_,
    g748_n
  );


  buf

  (
    g757_n_spl_,
    g757_n
  );


  buf

  (
    g748_p_spl_,
    g748_p
  );


  buf

  (
    g758_n_spl_,
    g758_n
  );


  buf

  (
    g758_p_spl_,
    g758_p
  );


  buf

  (
    g760_p_spl_,
    g760_p
  );


  buf

  (
    g747_n_spl_,
    g747_n
  );


  buf

  (
    g760_n_spl_,
    g760_n
  );


  buf

  (
    g747_p_spl_,
    g747_p
  );


  buf

  (
    g761_n_spl_,
    g761_n
  );


  buf

  (
    g761_p_spl_,
    g761_p
  );


  buf

  (
    g763_p_spl_,
    g763_p
  );


  buf

  (
    g746_n_spl_,
    g746_n
  );


  buf

  (
    g763_n_spl_,
    g763_n
  );


  buf

  (
    g746_p_spl_,
    g746_p
  );


  buf

  (
    g764_n_spl_,
    g764_n
  );


  buf

  (
    g764_p_spl_,
    g764_p
  );


  buf

  (
    g766_p_spl_,
    g766_p
  );


  buf

  (
    g745_n_spl_,
    g745_n
  );


  buf

  (
    g766_n_spl_,
    g766_n
  );


  buf

  (
    g745_p_spl_,
    g745_p
  );


  buf

  (
    g767_n_spl_,
    g767_n
  );


  buf

  (
    g767_p_spl_,
    g767_p
  );


  buf

  (
    g769_p_spl_,
    g769_p
  );


  buf

  (
    g744_n_spl_,
    g744_n
  );


  buf

  (
    g769_n_spl_,
    g769_n
  );


  buf

  (
    g744_p_spl_,
    g744_p
  );


  buf

  (
    g770_n_spl_,
    g770_n
  );


  buf

  (
    g770_p_spl_,
    g770_p
  );


  buf

  (
    g772_p_spl_,
    g772_p
  );


  buf

  (
    g743_n_spl_,
    g743_n
  );


  buf

  (
    g772_n_spl_,
    g772_n
  );


  buf

  (
    g743_p_spl_,
    g743_p
  );


  buf

  (
    g773_n_spl_,
    g773_n
  );


  buf

  (
    g773_p_spl_,
    g773_p
  );


  buf

  (
    g775_p_spl_,
    g775_p
  );


  buf

  (
    g742_n_spl_,
    g742_n
  );


  buf

  (
    g775_n_spl_,
    g775_n
  );


  buf

  (
    g742_p_spl_,
    g742_p
  );


  buf

  (
    g776_n_spl_,
    g776_n
  );


  buf

  (
    g776_p_spl_,
    g776_p
  );


  buf

  (
    g778_p_spl_,
    g778_p
  );


  buf

  (
    g741_n_spl_,
    g741_n
  );


  buf

  (
    g778_n_spl_,
    g778_n
  );


  buf

  (
    g741_p_spl_,
    g741_p
  );


  buf

  (
    g779_n_spl_,
    g779_n
  );


  buf

  (
    g779_p_spl_,
    g779_p
  );


  buf

  (
    g781_p_spl_,
    g781_p
  );


  buf

  (
    g740_n_spl_,
    g740_n
  );


  buf

  (
    g781_n_spl_,
    g781_n
  );


  buf

  (
    g740_p_spl_,
    g740_p
  );


  buf

  (
    g782_n_spl_,
    g782_n
  );


  buf

  (
    g782_p_spl_,
    g782_p
  );


  buf

  (
    g784_p_spl_,
    g784_p
  );


  buf

  (
    g739_n_spl_,
    g739_n
  );


  buf

  (
    g784_n_spl_,
    g784_n
  );


  buf

  (
    g739_p_spl_,
    g739_p
  );


  buf

  (
    g785_n_spl_,
    g785_n
  );


  buf

  (
    g785_p_spl_,
    g785_p
  );


  buf

  (
    g787_p_spl_,
    g787_p
  );


  buf

  (
    g738_n_spl_,
    g738_n
  );


  buf

  (
    g787_n_spl_,
    g787_n
  );


  buf

  (
    g738_p_spl_,
    g738_p
  );


  buf

  (
    g788_n_spl_,
    g788_n
  );


  buf

  (
    g788_p_spl_,
    g788_p
  );


  buf

  (
    g790_p_spl_,
    g790_p
  );


  buf

  (
    g737_n_spl_,
    g737_n
  );


  buf

  (
    g790_n_spl_,
    g790_n
  );


  buf

  (
    g737_p_spl_,
    g737_p
  );


  buf

  (
    g791_n_spl_,
    g791_n
  );


  buf

  (
    g791_p_spl_,
    g791_p
  );


  buf

  (
    g793_p_spl_,
    g793_p
  );


  buf

  (
    g736_n_spl_,
    g736_n
  );


  buf

  (
    g793_n_spl_,
    g793_n
  );


  buf

  (
    g736_p_spl_,
    g736_p
  );


  buf

  (
    g794_n_spl_,
    g794_n
  );


  buf

  (
    g794_p_spl_,
    g794_p
  );


  buf

  (
    g796_p_spl_,
    g796_p
  );


  buf

  (
    g735_n_spl_,
    g735_n
  );


  buf

  (
    g796_n_spl_,
    g796_n
  );


  buf

  (
    g735_p_spl_,
    g735_p
  );


  buf

  (
    g797_n_spl_,
    g797_n
  );


  buf

  (
    g797_p_spl_,
    g797_p
  );


  buf

  (
    g799_p_spl_,
    g799_p
  );


  buf

  (
    g734_n_spl_,
    g734_n
  );


  buf

  (
    g799_n_spl_,
    g799_n
  );


  buf

  (
    g734_p_spl_,
    g734_p
  );


  buf

  (
    g800_n_spl_,
    g800_n
  );


  buf

  (
    g800_p_spl_,
    g800_p
  );


  buf

  (
    g802_p_spl_,
    g802_p
  );


  buf

  (
    g733_n_spl_,
    g733_n
  );


  buf

  (
    g802_n_spl_,
    g802_n
  );


  buf

  (
    g733_p_spl_,
    g733_p
  );


  buf

  (
    g803_n_spl_,
    g803_n
  );


  buf

  (
    g803_p_spl_,
    g803_p
  );


  buf

  (
    g805_p_spl_,
    g805_p
  );


  buf

  (
    g732_n_spl_,
    g732_n
  );


  buf

  (
    g805_n_spl_,
    g805_n
  );


  buf

  (
    g732_p_spl_,
    g732_p
  );


  buf

  (
    g806_n_spl_,
    g806_n
  );


  buf

  (
    g806_p_spl_,
    g806_p
  );


  buf

  (
    g808_p_spl_,
    g808_p
  );


  buf

  (
    g731_n_spl_,
    g731_n
  );


  buf

  (
    g808_n_spl_,
    g808_n
  );


  buf

  (
    g731_p_spl_,
    g731_p
  );


  buf

  (
    g809_n_spl_,
    g809_n
  );


  buf

  (
    g809_p_spl_,
    g809_p
  );


  buf

  (
    g811_p_spl_,
    g811_p
  );


  buf

  (
    g730_n_spl_,
    g730_n
  );


  buf

  (
    g811_n_spl_,
    g811_n
  );


  buf

  (
    g730_p_spl_,
    g730_p
  );


  buf

  (
    g812_n_spl_,
    g812_n
  );


  buf

  (
    g812_p_spl_,
    g812_p
  );


  buf

  (
    g814_p_spl_,
    g814_p
  );


  buf

  (
    g729_n_spl_,
    g729_n
  );


  buf

  (
    g814_n_spl_,
    g814_n
  );


  buf

  (
    g729_p_spl_,
    g729_p
  );


  buf

  (
    g815_n_spl_,
    g815_n
  );


  buf

  (
    g815_p_spl_,
    g815_p
  );


  buf

  (
    g817_p_spl_,
    g817_p
  );


  buf

  (
    g728_n_spl_,
    g728_n
  );


  buf

  (
    g817_n_spl_,
    g817_n
  );


  buf

  (
    g728_p_spl_,
    g728_p
  );


  buf

  (
    g818_n_spl_,
    g818_n
  );


  buf

  (
    g818_p_spl_,
    g818_p
  );


  buf

  (
    g820_p_spl_,
    g820_p
  );


  buf

  (
    g727_n_spl_,
    g727_n
  );


  buf

  (
    g820_n_spl_,
    g820_n
  );


  buf

  (
    g727_p_spl_,
    g727_p
  );


  buf

  (
    g821_n_spl_,
    g821_n
  );


  buf

  (
    g821_p_spl_,
    g821_p
  );


  buf

  (
    g823_p_spl_,
    g823_p
  );


  buf

  (
    g726_n_spl_,
    g726_n
  );


  buf

  (
    g823_n_spl_,
    g823_n
  );


  buf

  (
    g726_p_spl_,
    g726_p
  );


  buf

  (
    g824_n_spl_,
    g824_n
  );


  buf

  (
    g824_p_spl_,
    g824_p
  );


  buf

  (
    g826_p_spl_,
    g826_p
  );


  buf

  (
    g725_n_spl_,
    g725_n
  );


  buf

  (
    g826_n_spl_,
    g826_n
  );


  buf

  (
    g725_p_spl_,
    g725_p
  );


  buf

  (
    g827_n_spl_,
    g827_n
  );


  buf

  (
    g827_p_spl_,
    g827_p
  );


  buf

  (
    g829_n_spl_,
    g829_n
  );


  buf

  (
    g724_p_spl_,
    g724_p
  );


  buf

  (
    g830_p_spl_,
    g830_p
  );


  buf

  (
    G32_p_spl_,
    G32_p
  );


  buf

  (
    G32_p_spl_0,
    G32_p_spl_
  );


  buf

  (
    G32_p_spl_00,
    G32_p_spl_0
  );


  buf

  (
    G32_p_spl_000,
    G32_p_spl_00
  );


  buf

  (
    G32_p_spl_001,
    G32_p_spl_00
  );


  buf

  (
    G32_p_spl_01,
    G32_p_spl_0
  );


  buf

  (
    G32_p_spl_010,
    G32_p_spl_01
  );


  buf

  (
    G32_p_spl_011,
    G32_p_spl_01
  );


  buf

  (
    G32_p_spl_1,
    G32_p_spl_
  );


  buf

  (
    G32_p_spl_10,
    G32_p_spl_1
  );


  buf

  (
    G32_p_spl_100,
    G32_p_spl_10
  );


  buf

  (
    G32_p_spl_101,
    G32_p_spl_10
  );


  buf

  (
    G32_p_spl_11,
    G32_p_spl_1
  );


  buf

  (
    G32_p_spl_110,
    G32_p_spl_11
  );


  buf

  (
    G32_p_spl_111,
    G32_p_spl_11
  );


  buf

  (
    G32_n_spl_,
    G32_n
  );


  buf

  (
    G32_n_spl_0,
    G32_n_spl_
  );


  buf

  (
    G32_n_spl_00,
    G32_n_spl_0
  );


  buf

  (
    G32_n_spl_000,
    G32_n_spl_00
  );


  buf

  (
    G32_n_spl_001,
    G32_n_spl_00
  );


  buf

  (
    G32_n_spl_01,
    G32_n_spl_0
  );


  buf

  (
    G32_n_spl_010,
    G32_n_spl_01
  );


  buf

  (
    G32_n_spl_011,
    G32_n_spl_01
  );


  buf

  (
    G32_n_spl_1,
    G32_n_spl_
  );


  buf

  (
    G32_n_spl_10,
    G32_n_spl_1
  );


  buf

  (
    G32_n_spl_100,
    G32_n_spl_10
  );


  buf

  (
    G32_n_spl_101,
    G32_n_spl_10
  );


  buf

  (
    G32_n_spl_11,
    G32_n_spl_1
  );


  buf

  (
    G32_n_spl_110,
    G32_n_spl_11
  );


  buf

  (
    G32_n_spl_111,
    G32_n_spl_11
  );


  buf

  (
    G16_p_spl_,
    G16_p
  );


  buf

  (
    G16_p_spl_0,
    G16_p_spl_
  );


  buf

  (
    G16_p_spl_00,
    G16_p_spl_0
  );


  buf

  (
    G16_p_spl_000,
    G16_p_spl_00
  );


  buf

  (
    G16_p_spl_001,
    G16_p_spl_00
  );


  buf

  (
    G16_p_spl_01,
    G16_p_spl_0
  );


  buf

  (
    G16_p_spl_010,
    G16_p_spl_01
  );


  buf

  (
    G16_p_spl_011,
    G16_p_spl_01
  );


  buf

  (
    G16_p_spl_1,
    G16_p_spl_
  );


  buf

  (
    G16_p_spl_10,
    G16_p_spl_1
  );


  buf

  (
    G16_p_spl_100,
    G16_p_spl_10
  );


  buf

  (
    G16_p_spl_101,
    G16_p_spl_10
  );


  buf

  (
    G16_p_spl_11,
    G16_p_spl_1
  );


  buf

  (
    G16_p_spl_110,
    G16_p_spl_11
  );


  buf

  (
    G16_p_spl_111,
    G16_p_spl_11
  );


  buf

  (
    G16_n_spl_,
    G16_n
  );


  buf

  (
    G16_n_spl_0,
    G16_n_spl_
  );


  buf

  (
    G16_n_spl_00,
    G16_n_spl_0
  );


  buf

  (
    G16_n_spl_000,
    G16_n_spl_00
  );


  buf

  (
    G16_n_spl_001,
    G16_n_spl_00
  );


  buf

  (
    G16_n_spl_01,
    G16_n_spl_0
  );


  buf

  (
    G16_n_spl_010,
    G16_n_spl_01
  );


  buf

  (
    G16_n_spl_011,
    G16_n_spl_01
  );


  buf

  (
    G16_n_spl_1,
    G16_n_spl_
  );


  buf

  (
    G16_n_spl_10,
    G16_n_spl_1
  );


  buf

  (
    G16_n_spl_100,
    G16_n_spl_10
  );


  buf

  (
    G16_n_spl_101,
    G16_n_spl_10
  );


  buf

  (
    G16_n_spl_11,
    G16_n_spl_1
  );


  buf

  (
    G16_n_spl_110,
    G16_n_spl_11
  );


  buf

  (
    G16_n_spl_111,
    G16_n_spl_11
  );


  buf

  (
    g861_n_spl_,
    g861_n
  );


  buf

  (
    g860_p_spl_,
    g860_p
  );


  buf

  (
    g861_p_spl_,
    g861_p
  );


  buf

  (
    g860_n_spl_,
    g860_n
  );


  buf

  (
    g862_n_spl_,
    g862_n
  );


  buf

  (
    g862_p_spl_,
    g862_p
  );


  buf

  (
    g863_n_spl_,
    g863_n
  );


  buf

  (
    g863_p_spl_,
    g863_p
  );


  buf

  (
    g865_n_spl_,
    g865_n
  );


  buf

  (
    g865_p_spl_,
    g865_p
  );


  buf

  (
    g866_n_spl_,
    g866_n
  );


  buf

  (
    g866_p_spl_,
    g866_p
  );


  buf

  (
    g868_p_spl_,
    g868_p
  );


  buf

  (
    g859_n_spl_,
    g859_n
  );


  buf

  (
    g868_n_spl_,
    g868_n
  );


  buf

  (
    g859_p_spl_,
    g859_p
  );


  buf

  (
    g869_n_spl_,
    g869_n
  );


  buf

  (
    g869_p_spl_,
    g869_p
  );


  buf

  (
    g871_p_spl_,
    g871_p
  );


  buf

  (
    g858_n_spl_,
    g858_n
  );


  buf

  (
    g871_n_spl_,
    g871_n
  );


  buf

  (
    g858_p_spl_,
    g858_p
  );


  buf

  (
    g872_n_spl_,
    g872_n
  );


  buf

  (
    g872_p_spl_,
    g872_p
  );


  buf

  (
    g874_p_spl_,
    g874_p
  );


  buf

  (
    g857_n_spl_,
    g857_n
  );


  buf

  (
    g874_n_spl_,
    g874_n
  );


  buf

  (
    g857_p_spl_,
    g857_p
  );


  buf

  (
    g875_n_spl_,
    g875_n
  );


  buf

  (
    g875_p_spl_,
    g875_p
  );


  buf

  (
    g877_p_spl_,
    g877_p
  );


  buf

  (
    g856_n_spl_,
    g856_n
  );


  buf

  (
    g877_n_spl_,
    g877_n
  );


  buf

  (
    g856_p_spl_,
    g856_p
  );


  buf

  (
    g878_n_spl_,
    g878_n
  );


  buf

  (
    g878_p_spl_,
    g878_p
  );


  buf

  (
    g880_p_spl_,
    g880_p
  );


  buf

  (
    g855_n_spl_,
    g855_n
  );


  buf

  (
    g880_n_spl_,
    g880_n
  );


  buf

  (
    g855_p_spl_,
    g855_p
  );


  buf

  (
    g881_n_spl_,
    g881_n
  );


  buf

  (
    g881_p_spl_,
    g881_p
  );


  buf

  (
    g883_p_spl_,
    g883_p
  );


  buf

  (
    g854_n_spl_,
    g854_n
  );


  buf

  (
    g883_n_spl_,
    g883_n
  );


  buf

  (
    g854_p_spl_,
    g854_p
  );


  buf

  (
    g884_n_spl_,
    g884_n
  );


  buf

  (
    g884_p_spl_,
    g884_p
  );


  buf

  (
    g886_p_spl_,
    g886_p
  );


  buf

  (
    g853_n_spl_,
    g853_n
  );


  buf

  (
    g886_n_spl_,
    g886_n
  );


  buf

  (
    g853_p_spl_,
    g853_p
  );


  buf

  (
    g887_n_spl_,
    g887_n
  );


  buf

  (
    g887_p_spl_,
    g887_p
  );


  buf

  (
    g889_p_spl_,
    g889_p
  );


  buf

  (
    g852_n_spl_,
    g852_n
  );


  buf

  (
    g889_n_spl_,
    g889_n
  );


  buf

  (
    g852_p_spl_,
    g852_p
  );


  buf

  (
    g890_n_spl_,
    g890_n
  );


  buf

  (
    g890_p_spl_,
    g890_p
  );


  buf

  (
    g892_p_spl_,
    g892_p
  );


  buf

  (
    g851_n_spl_,
    g851_n
  );


  buf

  (
    g892_n_spl_,
    g892_n
  );


  buf

  (
    g851_p_spl_,
    g851_p
  );


  buf

  (
    g893_n_spl_,
    g893_n
  );


  buf

  (
    g893_p_spl_,
    g893_p
  );


  buf

  (
    g895_p_spl_,
    g895_p
  );


  buf

  (
    g850_n_spl_,
    g850_n
  );


  buf

  (
    g895_n_spl_,
    g895_n
  );


  buf

  (
    g850_p_spl_,
    g850_p
  );


  buf

  (
    g896_n_spl_,
    g896_n
  );


  buf

  (
    g896_p_spl_,
    g896_p
  );


  buf

  (
    g898_p_spl_,
    g898_p
  );


  buf

  (
    g849_n_spl_,
    g849_n
  );


  buf

  (
    g898_n_spl_,
    g898_n
  );


  buf

  (
    g849_p_spl_,
    g849_p
  );


  buf

  (
    g899_n_spl_,
    g899_n
  );


  buf

  (
    g899_p_spl_,
    g899_p
  );


  buf

  (
    g901_p_spl_,
    g901_p
  );


  buf

  (
    g848_n_spl_,
    g848_n
  );


  buf

  (
    g901_n_spl_,
    g901_n
  );


  buf

  (
    g848_p_spl_,
    g848_p
  );


  buf

  (
    g902_n_spl_,
    g902_n
  );


  buf

  (
    g902_p_spl_,
    g902_p
  );


  buf

  (
    g904_p_spl_,
    g904_p
  );


  buf

  (
    g847_n_spl_,
    g847_n
  );


  buf

  (
    g904_n_spl_,
    g904_n
  );


  buf

  (
    g847_p_spl_,
    g847_p
  );


  buf

  (
    g905_n_spl_,
    g905_n
  );


  buf

  (
    g905_p_spl_,
    g905_p
  );


  buf

  (
    g907_p_spl_,
    g907_p
  );


  buf

  (
    g846_n_spl_,
    g846_n
  );


  buf

  (
    g907_n_spl_,
    g907_n
  );


  buf

  (
    g846_p_spl_,
    g846_p
  );


  buf

  (
    g908_n_spl_,
    g908_n
  );


  buf

  (
    g908_p_spl_,
    g908_p
  );


  buf

  (
    g910_p_spl_,
    g910_p
  );


  buf

  (
    g845_n_spl_,
    g845_n
  );


  buf

  (
    g910_n_spl_,
    g910_n
  );


  buf

  (
    g845_p_spl_,
    g845_p
  );


  buf

  (
    g911_n_spl_,
    g911_n
  );


  buf

  (
    g911_p_spl_,
    g911_p
  );


  buf

  (
    g913_p_spl_,
    g913_p
  );


  buf

  (
    g844_n_spl_,
    g844_n
  );


  buf

  (
    g913_n_spl_,
    g913_n
  );


  buf

  (
    g844_p_spl_,
    g844_p
  );


  buf

  (
    g914_n_spl_,
    g914_n
  );


  buf

  (
    g914_p_spl_,
    g914_p
  );


  buf

  (
    g916_p_spl_,
    g916_p
  );


  buf

  (
    g843_n_spl_,
    g843_n
  );


  buf

  (
    g916_n_spl_,
    g916_n
  );


  buf

  (
    g843_p_spl_,
    g843_p
  );


  buf

  (
    g917_n_spl_,
    g917_n
  );


  buf

  (
    g917_p_spl_,
    g917_p
  );


  buf

  (
    g919_p_spl_,
    g919_p
  );


  buf

  (
    g842_n_spl_,
    g842_n
  );


  buf

  (
    g919_n_spl_,
    g919_n
  );


  buf

  (
    g842_p_spl_,
    g842_p
  );


  buf

  (
    g920_n_spl_,
    g920_n
  );


  buf

  (
    g920_p_spl_,
    g920_p
  );


  buf

  (
    g922_p_spl_,
    g922_p
  );


  buf

  (
    g841_n_spl_,
    g841_n
  );


  buf

  (
    g922_n_spl_,
    g922_n
  );


  buf

  (
    g841_p_spl_,
    g841_p
  );


  buf

  (
    g923_n_spl_,
    g923_n
  );


  buf

  (
    g923_p_spl_,
    g923_p
  );


  buf

  (
    g925_p_spl_,
    g925_p
  );


  buf

  (
    g840_n_spl_,
    g840_n
  );


  buf

  (
    g925_n_spl_,
    g925_n
  );


  buf

  (
    g840_p_spl_,
    g840_p
  );


  buf

  (
    g926_n_spl_,
    g926_n
  );


  buf

  (
    g926_p_spl_,
    g926_p
  );


  buf

  (
    g928_p_spl_,
    g928_p
  );


  buf

  (
    g839_n_spl_,
    g839_n
  );


  buf

  (
    g928_n_spl_,
    g928_n
  );


  buf

  (
    g839_p_spl_,
    g839_p
  );


  buf

  (
    g929_n_spl_,
    g929_n
  );


  buf

  (
    g929_p_spl_,
    g929_p
  );


  buf

  (
    g931_p_spl_,
    g931_p
  );


  buf

  (
    g838_n_spl_,
    g838_n
  );


  buf

  (
    g931_n_spl_,
    g931_n
  );


  buf

  (
    g838_p_spl_,
    g838_p
  );


  buf

  (
    g932_n_spl_,
    g932_n
  );


  buf

  (
    g932_p_spl_,
    g932_p
  );


  buf

  (
    g934_p_spl_,
    g934_p
  );


  buf

  (
    g837_n_spl_,
    g837_n
  );


  buf

  (
    g934_n_spl_,
    g934_n
  );


  buf

  (
    g837_p_spl_,
    g837_p
  );


  buf

  (
    g935_n_spl_,
    g935_n
  );


  buf

  (
    g935_p_spl_,
    g935_p
  );


  buf

  (
    g937_p_spl_,
    g937_p
  );


  buf

  (
    g836_n_spl_,
    g836_n
  );


  buf

  (
    g937_n_spl_,
    g937_n
  );


  buf

  (
    g836_p_spl_,
    g836_p
  );


  buf

  (
    g938_n_spl_,
    g938_n
  );


  buf

  (
    g938_p_spl_,
    g938_p
  );


  buf

  (
    g940_p_spl_,
    g940_p
  );


  buf

  (
    g835_n_spl_,
    g835_n
  );


  buf

  (
    g940_n_spl_,
    g940_n
  );


  buf

  (
    g835_p_spl_,
    g835_p
  );


  buf

  (
    g941_n_spl_,
    g941_n
  );


  buf

  (
    g941_p_spl_,
    g941_p
  );


  buf

  (
    g943_p_spl_,
    g943_p
  );


  buf

  (
    g834_n_spl_,
    g834_n
  );


  buf

  (
    g943_n_spl_,
    g943_n
  );


  buf

  (
    g834_p_spl_,
    g834_p
  );


  buf

  (
    g944_n_spl_,
    g944_n
  );


  buf

  (
    g944_p_spl_,
    g944_p
  );


  buf

  (
    g946_n_spl_,
    g946_n
  );


  buf

  (
    g833_p_spl_,
    g833_p
  );


  buf

  (
    g947_p_spl_,
    g947_p
  );


  buf

  (
    g977_p_spl_,
    g977_p
  );


  buf

  (
    g977_n_spl_,
    g977_n
  );


  buf

  (
    g979_n_spl_,
    g979_n
  );


  buf

  (
    g978_p_spl_,
    g978_p
  );


  buf

  (
    g979_p_spl_,
    g979_p
  );


  buf

  (
    g978_n_spl_,
    g978_n
  );


  buf

  (
    g980_n_spl_,
    g980_n
  );


  buf

  (
    g980_p_spl_,
    g980_p
  );


  buf

  (
    g982_p_spl_,
    g982_p
  );


  buf

  (
    g976_n_spl_,
    g976_n
  );


  buf

  (
    g982_n_spl_,
    g982_n
  );


  buf

  (
    g976_p_spl_,
    g976_p
  );


  buf

  (
    g983_n_spl_,
    g983_n
  );


  buf

  (
    g983_p_spl_,
    g983_p
  );


  buf

  (
    g985_p_spl_,
    g985_p
  );


  buf

  (
    g975_n_spl_,
    g975_n
  );


  buf

  (
    g985_n_spl_,
    g985_n
  );


  buf

  (
    g975_p_spl_,
    g975_p
  );


  buf

  (
    g986_n_spl_,
    g986_n
  );


  buf

  (
    g986_p_spl_,
    g986_p
  );


  buf

  (
    g988_p_spl_,
    g988_p
  );


  buf

  (
    g974_n_spl_,
    g974_n
  );


  buf

  (
    g988_n_spl_,
    g988_n
  );


  buf

  (
    g974_p_spl_,
    g974_p
  );


  buf

  (
    g989_n_spl_,
    g989_n
  );


  buf

  (
    g989_p_spl_,
    g989_p
  );


  buf

  (
    g991_p_spl_,
    g991_p
  );


  buf

  (
    g973_n_spl_,
    g973_n
  );


  buf

  (
    g991_n_spl_,
    g991_n
  );


  buf

  (
    g973_p_spl_,
    g973_p
  );


  buf

  (
    g992_n_spl_,
    g992_n
  );


  buf

  (
    g992_p_spl_,
    g992_p
  );


  buf

  (
    g994_p_spl_,
    g994_p
  );


  buf

  (
    g972_n_spl_,
    g972_n
  );


  buf

  (
    g994_n_spl_,
    g994_n
  );


  buf

  (
    g972_p_spl_,
    g972_p
  );


  buf

  (
    g995_n_spl_,
    g995_n
  );


  buf

  (
    g995_p_spl_,
    g995_p
  );


  buf

  (
    g997_p_spl_,
    g997_p
  );


  buf

  (
    g971_n_spl_,
    g971_n
  );


  buf

  (
    g997_n_spl_,
    g997_n
  );


  buf

  (
    g971_p_spl_,
    g971_p
  );


  buf

  (
    g998_n_spl_,
    g998_n
  );


  buf

  (
    g998_p_spl_,
    g998_p
  );


  buf

  (
    g1000_p_spl_,
    g1000_p
  );


  buf

  (
    g970_n_spl_,
    g970_n
  );


  buf

  (
    g1000_n_spl_,
    g1000_n
  );


  buf

  (
    g970_p_spl_,
    g970_p
  );


  buf

  (
    g1001_n_spl_,
    g1001_n
  );


  buf

  (
    g1001_p_spl_,
    g1001_p
  );


  buf

  (
    g1003_p_spl_,
    g1003_p
  );


  buf

  (
    g969_n_spl_,
    g969_n
  );


  buf

  (
    g1003_n_spl_,
    g1003_n
  );


  buf

  (
    g969_p_spl_,
    g969_p
  );


  buf

  (
    g1004_n_spl_,
    g1004_n
  );


  buf

  (
    g1004_p_spl_,
    g1004_p
  );


  buf

  (
    g1006_p_spl_,
    g1006_p
  );


  buf

  (
    g968_n_spl_,
    g968_n
  );


  buf

  (
    g1006_n_spl_,
    g1006_n
  );


  buf

  (
    g968_p_spl_,
    g968_p
  );


  buf

  (
    g1007_n_spl_,
    g1007_n
  );


  buf

  (
    g1007_p_spl_,
    g1007_p
  );


  buf

  (
    g1009_p_spl_,
    g1009_p
  );


  buf

  (
    g967_n_spl_,
    g967_n
  );


  buf

  (
    g1009_n_spl_,
    g1009_n
  );


  buf

  (
    g967_p_spl_,
    g967_p
  );


  buf

  (
    g1010_n_spl_,
    g1010_n
  );


  buf

  (
    g1010_p_spl_,
    g1010_p
  );


  buf

  (
    g1012_p_spl_,
    g1012_p
  );


  buf

  (
    g966_n_spl_,
    g966_n
  );


  buf

  (
    g1012_n_spl_,
    g1012_n
  );


  buf

  (
    g966_p_spl_,
    g966_p
  );


  buf

  (
    g1013_n_spl_,
    g1013_n
  );


  buf

  (
    g1013_p_spl_,
    g1013_p
  );


  buf

  (
    g1015_p_spl_,
    g1015_p
  );


  buf

  (
    g965_n_spl_,
    g965_n
  );


  buf

  (
    g1015_n_spl_,
    g1015_n
  );


  buf

  (
    g965_p_spl_,
    g965_p
  );


  buf

  (
    g1016_n_spl_,
    g1016_n
  );


  buf

  (
    g1016_p_spl_,
    g1016_p
  );


  buf

  (
    g1018_p_spl_,
    g1018_p
  );


  buf

  (
    g964_n_spl_,
    g964_n
  );


  buf

  (
    g1018_n_spl_,
    g1018_n
  );


  buf

  (
    g964_p_spl_,
    g964_p
  );


  buf

  (
    g1019_n_spl_,
    g1019_n
  );


  buf

  (
    g1019_p_spl_,
    g1019_p
  );


  buf

  (
    g1021_p_spl_,
    g1021_p
  );


  buf

  (
    g963_n_spl_,
    g963_n
  );


  buf

  (
    g1021_n_spl_,
    g1021_n
  );


  buf

  (
    g963_p_spl_,
    g963_p
  );


  buf

  (
    g1022_n_spl_,
    g1022_n
  );


  buf

  (
    g1022_p_spl_,
    g1022_p
  );


  buf

  (
    g1024_p_spl_,
    g1024_p
  );


  buf

  (
    g962_n_spl_,
    g962_n
  );


  buf

  (
    g1024_n_spl_,
    g1024_n
  );


  buf

  (
    g962_p_spl_,
    g962_p
  );


  buf

  (
    g1025_n_spl_,
    g1025_n
  );


  buf

  (
    g1025_p_spl_,
    g1025_p
  );


  buf

  (
    g1027_p_spl_,
    g1027_p
  );


  buf

  (
    g961_n_spl_,
    g961_n
  );


  buf

  (
    g1027_n_spl_,
    g1027_n
  );


  buf

  (
    g961_p_spl_,
    g961_p
  );


  buf

  (
    g1028_n_spl_,
    g1028_n
  );


  buf

  (
    g1028_p_spl_,
    g1028_p
  );


  buf

  (
    g1030_p_spl_,
    g1030_p
  );


  buf

  (
    g960_n_spl_,
    g960_n
  );


  buf

  (
    g1030_n_spl_,
    g1030_n
  );


  buf

  (
    g960_p_spl_,
    g960_p
  );


  buf

  (
    g1031_n_spl_,
    g1031_n
  );


  buf

  (
    g1031_p_spl_,
    g1031_p
  );


  buf

  (
    g1033_p_spl_,
    g1033_p
  );


  buf

  (
    g959_n_spl_,
    g959_n
  );


  buf

  (
    g1033_n_spl_,
    g1033_n
  );


  buf

  (
    g959_p_spl_,
    g959_p
  );


  buf

  (
    g1034_n_spl_,
    g1034_n
  );


  buf

  (
    g1034_p_spl_,
    g1034_p
  );


  buf

  (
    g1036_p_spl_,
    g1036_p
  );


  buf

  (
    g958_n_spl_,
    g958_n
  );


  buf

  (
    g1036_n_spl_,
    g1036_n
  );


  buf

  (
    g958_p_spl_,
    g958_p
  );


  buf

  (
    g1037_n_spl_,
    g1037_n
  );


  buf

  (
    g1037_p_spl_,
    g1037_p
  );


  buf

  (
    g1039_p_spl_,
    g1039_p
  );


  buf

  (
    g957_n_spl_,
    g957_n
  );


  buf

  (
    g1039_n_spl_,
    g1039_n
  );


  buf

  (
    g957_p_spl_,
    g957_p
  );


  buf

  (
    g1040_n_spl_,
    g1040_n
  );


  buf

  (
    g1040_p_spl_,
    g1040_p
  );


  buf

  (
    g1042_p_spl_,
    g1042_p
  );


  buf

  (
    g956_n_spl_,
    g956_n
  );


  buf

  (
    g1042_n_spl_,
    g1042_n
  );


  buf

  (
    g956_p_spl_,
    g956_p
  );


  buf

  (
    g1043_n_spl_,
    g1043_n
  );


  buf

  (
    g1043_p_spl_,
    g1043_p
  );


  buf

  (
    g1045_p_spl_,
    g1045_p
  );


  buf

  (
    g955_n_spl_,
    g955_n
  );


  buf

  (
    g1045_n_spl_,
    g1045_n
  );


  buf

  (
    g955_p_spl_,
    g955_p
  );


  buf

  (
    g1046_n_spl_,
    g1046_n
  );


  buf

  (
    g1046_p_spl_,
    g1046_p
  );


  buf

  (
    g1048_p_spl_,
    g1048_p
  );


  buf

  (
    g954_n_spl_,
    g954_n
  );


  buf

  (
    g1048_n_spl_,
    g1048_n
  );


  buf

  (
    g954_p_spl_,
    g954_p
  );


  buf

  (
    g1049_n_spl_,
    g1049_n
  );


  buf

  (
    g1049_p_spl_,
    g1049_p
  );


  buf

  (
    g1051_p_spl_,
    g1051_p
  );


  buf

  (
    g953_n_spl_,
    g953_n
  );


  buf

  (
    g1051_n_spl_,
    g1051_n
  );


  buf

  (
    g953_p_spl_,
    g953_p
  );


  buf

  (
    g1052_n_spl_,
    g1052_n
  );


  buf

  (
    g1052_p_spl_,
    g1052_p
  );


  buf

  (
    g1054_p_spl_,
    g1054_p
  );


  buf

  (
    g952_n_spl_,
    g952_n
  );


  buf

  (
    g1054_n_spl_,
    g1054_n
  );


  buf

  (
    g952_p_spl_,
    g952_p
  );


  buf

  (
    g1055_n_spl_,
    g1055_n
  );


  buf

  (
    g1055_p_spl_,
    g1055_p
  );


  buf

  (
    g1057_p_spl_,
    g1057_p
  );


  buf

  (
    g951_n_spl_,
    g951_n
  );


  buf

  (
    g1057_n_spl_,
    g1057_n
  );


  buf

  (
    g951_p_spl_,
    g951_p
  );


  buf

  (
    g1058_n_spl_,
    g1058_n
  );


  buf

  (
    g1058_p_spl_,
    g1058_p
  );


  buf

  (
    g1060_n_spl_,
    g1060_n
  );


  buf

  (
    g950_p_spl_,
    g950_p
  );


  buf

  (
    g1062_n_spl_,
    g1062_n
  );


  buf

  (
    g1091_n_spl_,
    g1091_n
  );


  buf

  (
    g1090_n_spl_,
    g1090_n
  );


  buf

  (
    g1091_p_spl_,
    g1091_p
  );


  buf

  (
    g1090_p_spl_,
    g1090_p
  );


  buf

  (
    g1092_n_spl_,
    g1092_n
  );


  buf

  (
    g1092_p_spl_,
    g1092_p
  );


  buf

  (
    g1094_p_spl_,
    g1094_p
  );


  buf

  (
    g1089_n_spl_,
    g1089_n
  );


  buf

  (
    g1094_n_spl_,
    g1094_n
  );


  buf

  (
    g1089_p_spl_,
    g1089_p
  );


  buf

  (
    g1095_n_spl_,
    g1095_n
  );


  buf

  (
    g1095_p_spl_,
    g1095_p
  );


  buf

  (
    g1097_p_spl_,
    g1097_p
  );


  buf

  (
    g1088_n_spl_,
    g1088_n
  );


  buf

  (
    g1097_n_spl_,
    g1097_n
  );


  buf

  (
    g1088_p_spl_,
    g1088_p
  );


  buf

  (
    g1098_n_spl_,
    g1098_n
  );


  buf

  (
    g1098_p_spl_,
    g1098_p
  );


  buf

  (
    g1100_p_spl_,
    g1100_p
  );


  buf

  (
    g1087_n_spl_,
    g1087_n
  );


  buf

  (
    g1100_n_spl_,
    g1100_n
  );


  buf

  (
    g1087_p_spl_,
    g1087_p
  );


  buf

  (
    g1101_n_spl_,
    g1101_n
  );


  buf

  (
    g1101_p_spl_,
    g1101_p
  );


  buf

  (
    g1103_p_spl_,
    g1103_p
  );


  buf

  (
    g1086_n_spl_,
    g1086_n
  );


  buf

  (
    g1103_n_spl_,
    g1103_n
  );


  buf

  (
    g1086_p_spl_,
    g1086_p
  );


  buf

  (
    g1104_n_spl_,
    g1104_n
  );


  buf

  (
    g1104_p_spl_,
    g1104_p
  );


  buf

  (
    g1106_p_spl_,
    g1106_p
  );


  buf

  (
    g1085_n_spl_,
    g1085_n
  );


  buf

  (
    g1106_n_spl_,
    g1106_n
  );


  buf

  (
    g1085_p_spl_,
    g1085_p
  );


  buf

  (
    g1107_n_spl_,
    g1107_n
  );


  buf

  (
    g1107_p_spl_,
    g1107_p
  );


  buf

  (
    g1109_p_spl_,
    g1109_p
  );


  buf

  (
    g1084_n_spl_,
    g1084_n
  );


  buf

  (
    g1109_n_spl_,
    g1109_n
  );


  buf

  (
    g1084_p_spl_,
    g1084_p
  );


  buf

  (
    g1110_n_spl_,
    g1110_n
  );


  buf

  (
    g1110_p_spl_,
    g1110_p
  );


  buf

  (
    g1112_p_spl_,
    g1112_p
  );


  buf

  (
    g1083_n_spl_,
    g1083_n
  );


  buf

  (
    g1112_n_spl_,
    g1112_n
  );


  buf

  (
    g1083_p_spl_,
    g1083_p
  );


  buf

  (
    g1113_n_spl_,
    g1113_n
  );


  buf

  (
    g1113_p_spl_,
    g1113_p
  );


  buf

  (
    g1115_p_spl_,
    g1115_p
  );


  buf

  (
    g1082_n_spl_,
    g1082_n
  );


  buf

  (
    g1115_n_spl_,
    g1115_n
  );


  buf

  (
    g1082_p_spl_,
    g1082_p
  );


  buf

  (
    g1116_n_spl_,
    g1116_n
  );


  buf

  (
    g1116_p_spl_,
    g1116_p
  );


  buf

  (
    g1118_p_spl_,
    g1118_p
  );


  buf

  (
    g1081_n_spl_,
    g1081_n
  );


  buf

  (
    g1118_n_spl_,
    g1118_n
  );


  buf

  (
    g1081_p_spl_,
    g1081_p
  );


  buf

  (
    g1119_n_spl_,
    g1119_n
  );


  buf

  (
    g1119_p_spl_,
    g1119_p
  );


  buf

  (
    g1121_p_spl_,
    g1121_p
  );


  buf

  (
    g1080_n_spl_,
    g1080_n
  );


  buf

  (
    g1121_n_spl_,
    g1121_n
  );


  buf

  (
    g1080_p_spl_,
    g1080_p
  );


  buf

  (
    g1122_n_spl_,
    g1122_n
  );


  buf

  (
    g1122_p_spl_,
    g1122_p
  );


  buf

  (
    g1124_p_spl_,
    g1124_p
  );


  buf

  (
    g1079_n_spl_,
    g1079_n
  );


  buf

  (
    g1124_n_spl_,
    g1124_n
  );


  buf

  (
    g1079_p_spl_,
    g1079_p
  );


  buf

  (
    g1125_n_spl_,
    g1125_n
  );


  buf

  (
    g1125_p_spl_,
    g1125_p
  );


  buf

  (
    g1127_p_spl_,
    g1127_p
  );


  buf

  (
    g1078_n_spl_,
    g1078_n
  );


  buf

  (
    g1127_n_spl_,
    g1127_n
  );


  buf

  (
    g1078_p_spl_,
    g1078_p
  );


  buf

  (
    g1128_n_spl_,
    g1128_n
  );


  buf

  (
    g1128_p_spl_,
    g1128_p
  );


  buf

  (
    g1130_p_spl_,
    g1130_p
  );


  buf

  (
    g1077_n_spl_,
    g1077_n
  );


  buf

  (
    g1130_n_spl_,
    g1130_n
  );


  buf

  (
    g1077_p_spl_,
    g1077_p
  );


  buf

  (
    g1131_n_spl_,
    g1131_n
  );


  buf

  (
    g1131_p_spl_,
    g1131_p
  );


  buf

  (
    g1133_p_spl_,
    g1133_p
  );


  buf

  (
    g1076_n_spl_,
    g1076_n
  );


  buf

  (
    g1133_n_spl_,
    g1133_n
  );


  buf

  (
    g1076_p_spl_,
    g1076_p
  );


  buf

  (
    g1134_n_spl_,
    g1134_n
  );


  buf

  (
    g1134_p_spl_,
    g1134_p
  );


  buf

  (
    g1136_p_spl_,
    g1136_p
  );


  buf

  (
    g1075_n_spl_,
    g1075_n
  );


  buf

  (
    g1136_n_spl_,
    g1136_n
  );


  buf

  (
    g1075_p_spl_,
    g1075_p
  );


  buf

  (
    g1137_n_spl_,
    g1137_n
  );


  buf

  (
    g1137_p_spl_,
    g1137_p
  );


  buf

  (
    g1139_p_spl_,
    g1139_p
  );


  buf

  (
    g1074_n_spl_,
    g1074_n
  );


  buf

  (
    g1139_n_spl_,
    g1139_n
  );


  buf

  (
    g1074_p_spl_,
    g1074_p
  );


  buf

  (
    g1140_n_spl_,
    g1140_n
  );


  buf

  (
    g1140_p_spl_,
    g1140_p
  );


  buf

  (
    g1142_p_spl_,
    g1142_p
  );


  buf

  (
    g1073_n_spl_,
    g1073_n
  );


  buf

  (
    g1142_n_spl_,
    g1142_n
  );


  buf

  (
    g1073_p_spl_,
    g1073_p
  );


  buf

  (
    g1143_n_spl_,
    g1143_n
  );


  buf

  (
    g1143_p_spl_,
    g1143_p
  );


  buf

  (
    g1145_p_spl_,
    g1145_p
  );


  buf

  (
    g1072_n_spl_,
    g1072_n
  );


  buf

  (
    g1145_n_spl_,
    g1145_n
  );


  buf

  (
    g1072_p_spl_,
    g1072_p
  );


  buf

  (
    g1146_n_spl_,
    g1146_n
  );


  buf

  (
    g1146_p_spl_,
    g1146_p
  );


  buf

  (
    g1148_p_spl_,
    g1148_p
  );


  buf

  (
    g1071_n_spl_,
    g1071_n
  );


  buf

  (
    g1148_n_spl_,
    g1148_n
  );


  buf

  (
    g1071_p_spl_,
    g1071_p
  );


  buf

  (
    g1149_n_spl_,
    g1149_n
  );


  buf

  (
    g1149_p_spl_,
    g1149_p
  );


  buf

  (
    g1151_p_spl_,
    g1151_p
  );


  buf

  (
    g1070_n_spl_,
    g1070_n
  );


  buf

  (
    g1151_n_spl_,
    g1151_n
  );


  buf

  (
    g1070_p_spl_,
    g1070_p
  );


  buf

  (
    g1152_n_spl_,
    g1152_n
  );


  buf

  (
    g1152_p_spl_,
    g1152_p
  );


  buf

  (
    g1154_p_spl_,
    g1154_p
  );


  buf

  (
    g1069_n_spl_,
    g1069_n
  );


  buf

  (
    g1154_n_spl_,
    g1154_n
  );


  buf

  (
    g1069_p_spl_,
    g1069_p
  );


  buf

  (
    g1155_n_spl_,
    g1155_n
  );


  buf

  (
    g1155_p_spl_,
    g1155_p
  );


  buf

  (
    g1157_p_spl_,
    g1157_p
  );


  buf

  (
    g1068_n_spl_,
    g1068_n
  );


  buf

  (
    g1157_n_spl_,
    g1157_n
  );


  buf

  (
    g1068_p_spl_,
    g1068_p
  );


  buf

  (
    g1158_n_spl_,
    g1158_n
  );


  buf

  (
    g1158_p_spl_,
    g1158_p
  );


  buf

  (
    g1160_p_spl_,
    g1160_p
  );


  buf

  (
    g1067_n_spl_,
    g1067_n
  );


  buf

  (
    g1160_n_spl_,
    g1160_n
  );


  buf

  (
    g1067_p_spl_,
    g1067_p
  );


  buf

  (
    g1161_n_spl_,
    g1161_n
  );


  buf

  (
    g1161_p_spl_,
    g1161_p
  );


  buf

  (
    g1163_p_spl_,
    g1163_p
  );


  buf

  (
    g1066_n_spl_,
    g1066_n
  );


  buf

  (
    g1163_n_spl_,
    g1163_n
  );


  buf

  (
    g1066_p_spl_,
    g1066_p
  );


  buf

  (
    g1164_n_spl_,
    g1164_n
  );


  buf

  (
    g1164_p_spl_,
    g1164_p
  );


  buf

  (
    g1166_p_spl_,
    g1166_p
  );


  buf

  (
    g1065_n_spl_,
    g1065_n
  );


  buf

  (
    g1166_n_spl_,
    g1166_n
  );


  buf

  (
    g1065_p_spl_,
    g1065_p
  );


  buf

  (
    g1167_n_spl_,
    g1167_n
  );


  buf

  (
    g1167_p_spl_,
    g1167_p
  );


  buf

  (
    g1169_p_spl_,
    g1169_p
  );


  buf

  (
    g1064_n_spl_,
    g1064_n
  );


  buf

  (
    g1169_n_spl_,
    g1169_n
  );


  buf

  (
    g1064_p_spl_,
    g1064_p
  );


  buf

  (
    g1170_n_spl_,
    g1170_n
  );


  buf

  (
    g1170_p_spl_,
    g1170_p
  );


  buf

  (
    g1172_n_spl_,
    g1172_n
  );


  buf

  (
    g1062_p_spl_,
    g1062_p
  );


  buf

  (
    g1173_p_spl_,
    g1173_p
  );


  buf

  (
    g1202_n_spl_,
    g1202_n
  );


  buf

  (
    g1201_n_spl_,
    g1201_n
  );


  buf

  (
    g1202_p_spl_,
    g1202_p
  );


  buf

  (
    g1201_p_spl_,
    g1201_p
  );


  buf

  (
    g1203_n_spl_,
    g1203_n
  );


  buf

  (
    g1203_p_spl_,
    g1203_p
  );


  buf

  (
    g1205_p_spl_,
    g1205_p
  );


  buf

  (
    g1200_n_spl_,
    g1200_n
  );


  buf

  (
    g1205_n_spl_,
    g1205_n
  );


  buf

  (
    g1200_p_spl_,
    g1200_p
  );


  buf

  (
    g1206_n_spl_,
    g1206_n
  );


  buf

  (
    g1206_p_spl_,
    g1206_p
  );


  buf

  (
    g1208_p_spl_,
    g1208_p
  );


  buf

  (
    g1199_n_spl_,
    g1199_n
  );


  buf

  (
    g1208_n_spl_,
    g1208_n
  );


  buf

  (
    g1199_p_spl_,
    g1199_p
  );


  buf

  (
    g1209_n_spl_,
    g1209_n
  );


  buf

  (
    g1209_p_spl_,
    g1209_p
  );


  buf

  (
    g1211_p_spl_,
    g1211_p
  );


  buf

  (
    g1198_n_spl_,
    g1198_n
  );


  buf

  (
    g1211_n_spl_,
    g1211_n
  );


  buf

  (
    g1198_p_spl_,
    g1198_p
  );


  buf

  (
    g1212_n_spl_,
    g1212_n
  );


  buf

  (
    g1212_p_spl_,
    g1212_p
  );


  buf

  (
    g1214_p_spl_,
    g1214_p
  );


  buf

  (
    g1197_n_spl_,
    g1197_n
  );


  buf

  (
    g1214_n_spl_,
    g1214_n
  );


  buf

  (
    g1197_p_spl_,
    g1197_p
  );


  buf

  (
    g1215_n_spl_,
    g1215_n
  );


  buf

  (
    g1215_p_spl_,
    g1215_p
  );


  buf

  (
    g1217_p_spl_,
    g1217_p
  );


  buf

  (
    g1196_n_spl_,
    g1196_n
  );


  buf

  (
    g1217_n_spl_,
    g1217_n
  );


  buf

  (
    g1196_p_spl_,
    g1196_p
  );


  buf

  (
    g1218_n_spl_,
    g1218_n
  );


  buf

  (
    g1218_p_spl_,
    g1218_p
  );


  buf

  (
    g1220_p_spl_,
    g1220_p
  );


  buf

  (
    g1195_n_spl_,
    g1195_n
  );


  buf

  (
    g1220_n_spl_,
    g1220_n
  );


  buf

  (
    g1195_p_spl_,
    g1195_p
  );


  buf

  (
    g1221_n_spl_,
    g1221_n
  );


  buf

  (
    g1221_p_spl_,
    g1221_p
  );


  buf

  (
    g1223_p_spl_,
    g1223_p
  );


  buf

  (
    g1194_n_spl_,
    g1194_n
  );


  buf

  (
    g1223_n_spl_,
    g1223_n
  );


  buf

  (
    g1194_p_spl_,
    g1194_p
  );


  buf

  (
    g1224_n_spl_,
    g1224_n
  );


  buf

  (
    g1224_p_spl_,
    g1224_p
  );


  buf

  (
    g1226_p_spl_,
    g1226_p
  );


  buf

  (
    g1193_n_spl_,
    g1193_n
  );


  buf

  (
    g1226_n_spl_,
    g1226_n
  );


  buf

  (
    g1193_p_spl_,
    g1193_p
  );


  buf

  (
    g1227_n_spl_,
    g1227_n
  );


  buf

  (
    g1227_p_spl_,
    g1227_p
  );


  buf

  (
    g1229_p_spl_,
    g1229_p
  );


  buf

  (
    g1192_n_spl_,
    g1192_n
  );


  buf

  (
    g1229_n_spl_,
    g1229_n
  );


  buf

  (
    g1192_p_spl_,
    g1192_p
  );


  buf

  (
    g1230_n_spl_,
    g1230_n
  );


  buf

  (
    g1230_p_spl_,
    g1230_p
  );


  buf

  (
    g1232_p_spl_,
    g1232_p
  );


  buf

  (
    g1191_n_spl_,
    g1191_n
  );


  buf

  (
    g1232_n_spl_,
    g1232_n
  );


  buf

  (
    g1191_p_spl_,
    g1191_p
  );


  buf

  (
    g1233_n_spl_,
    g1233_n
  );


  buf

  (
    g1233_p_spl_,
    g1233_p
  );


  buf

  (
    g1235_p_spl_,
    g1235_p
  );


  buf

  (
    g1190_n_spl_,
    g1190_n
  );


  buf

  (
    g1235_n_spl_,
    g1235_n
  );


  buf

  (
    g1190_p_spl_,
    g1190_p
  );


  buf

  (
    g1236_n_spl_,
    g1236_n
  );


  buf

  (
    g1236_p_spl_,
    g1236_p
  );


  buf

  (
    g1238_p_spl_,
    g1238_p
  );


  buf

  (
    g1189_n_spl_,
    g1189_n
  );


  buf

  (
    g1238_n_spl_,
    g1238_n
  );


  buf

  (
    g1189_p_spl_,
    g1189_p
  );


  buf

  (
    g1239_n_spl_,
    g1239_n
  );


  buf

  (
    g1239_p_spl_,
    g1239_p
  );


  buf

  (
    g1241_p_spl_,
    g1241_p
  );


  buf

  (
    g1188_n_spl_,
    g1188_n
  );


  buf

  (
    g1241_n_spl_,
    g1241_n
  );


  buf

  (
    g1188_p_spl_,
    g1188_p
  );


  buf

  (
    g1242_n_spl_,
    g1242_n
  );


  buf

  (
    g1242_p_spl_,
    g1242_p
  );


  buf

  (
    g1244_p_spl_,
    g1244_p
  );


  buf

  (
    g1187_n_spl_,
    g1187_n
  );


  buf

  (
    g1244_n_spl_,
    g1244_n
  );


  buf

  (
    g1187_p_spl_,
    g1187_p
  );


  buf

  (
    g1245_n_spl_,
    g1245_n
  );


  buf

  (
    g1245_p_spl_,
    g1245_p
  );


  buf

  (
    g1247_p_spl_,
    g1247_p
  );


  buf

  (
    g1186_n_spl_,
    g1186_n
  );


  buf

  (
    g1247_n_spl_,
    g1247_n
  );


  buf

  (
    g1186_p_spl_,
    g1186_p
  );


  buf

  (
    g1248_n_spl_,
    g1248_n
  );


  buf

  (
    g1248_p_spl_,
    g1248_p
  );


  buf

  (
    g1250_p_spl_,
    g1250_p
  );


  buf

  (
    g1185_n_spl_,
    g1185_n
  );


  buf

  (
    g1250_n_spl_,
    g1250_n
  );


  buf

  (
    g1185_p_spl_,
    g1185_p
  );


  buf

  (
    g1251_n_spl_,
    g1251_n
  );


  buf

  (
    g1251_p_spl_,
    g1251_p
  );


  buf

  (
    g1253_p_spl_,
    g1253_p
  );


  buf

  (
    g1184_n_spl_,
    g1184_n
  );


  buf

  (
    g1253_n_spl_,
    g1253_n
  );


  buf

  (
    g1184_p_spl_,
    g1184_p
  );


  buf

  (
    g1254_n_spl_,
    g1254_n
  );


  buf

  (
    g1254_p_spl_,
    g1254_p
  );


  buf

  (
    g1256_p_spl_,
    g1256_p
  );


  buf

  (
    g1183_n_spl_,
    g1183_n
  );


  buf

  (
    g1256_n_spl_,
    g1256_n
  );


  buf

  (
    g1183_p_spl_,
    g1183_p
  );


  buf

  (
    g1257_n_spl_,
    g1257_n
  );


  buf

  (
    g1257_p_spl_,
    g1257_p
  );


  buf

  (
    g1259_p_spl_,
    g1259_p
  );


  buf

  (
    g1182_n_spl_,
    g1182_n
  );


  buf

  (
    g1259_n_spl_,
    g1259_n
  );


  buf

  (
    g1182_p_spl_,
    g1182_p
  );


  buf

  (
    g1260_n_spl_,
    g1260_n
  );


  buf

  (
    g1260_p_spl_,
    g1260_p
  );


  buf

  (
    g1262_p_spl_,
    g1262_p
  );


  buf

  (
    g1181_n_spl_,
    g1181_n
  );


  buf

  (
    g1262_n_spl_,
    g1262_n
  );


  buf

  (
    g1181_p_spl_,
    g1181_p
  );


  buf

  (
    g1263_n_spl_,
    g1263_n
  );


  buf

  (
    g1263_p_spl_,
    g1263_p
  );


  buf

  (
    g1265_p_spl_,
    g1265_p
  );


  buf

  (
    g1180_n_spl_,
    g1180_n
  );


  buf

  (
    g1265_n_spl_,
    g1265_n
  );


  buf

  (
    g1180_p_spl_,
    g1180_p
  );


  buf

  (
    g1266_n_spl_,
    g1266_n
  );


  buf

  (
    g1266_p_spl_,
    g1266_p
  );


  buf

  (
    g1268_p_spl_,
    g1268_p
  );


  buf

  (
    g1179_n_spl_,
    g1179_n
  );


  buf

  (
    g1268_n_spl_,
    g1268_n
  );


  buf

  (
    g1179_p_spl_,
    g1179_p
  );


  buf

  (
    g1269_n_spl_,
    g1269_n
  );


  buf

  (
    g1269_p_spl_,
    g1269_p
  );


  buf

  (
    g1271_p_spl_,
    g1271_p
  );


  buf

  (
    g1178_n_spl_,
    g1178_n
  );


  buf

  (
    g1271_n_spl_,
    g1271_n
  );


  buf

  (
    g1178_p_spl_,
    g1178_p
  );


  buf

  (
    g1272_n_spl_,
    g1272_n
  );


  buf

  (
    g1272_p_spl_,
    g1272_p
  );


  buf

  (
    g1274_p_spl_,
    g1274_p
  );


  buf

  (
    g1177_n_spl_,
    g1177_n
  );


  buf

  (
    g1274_n_spl_,
    g1274_n
  );


  buf

  (
    g1177_p_spl_,
    g1177_p
  );


  buf

  (
    g1275_n_spl_,
    g1275_n
  );


  buf

  (
    g1275_p_spl_,
    g1275_p
  );


  buf

  (
    g1277_n_spl_,
    g1277_n
  );


  buf

  (
    g1176_p_spl_,
    g1176_p
  );


  buf

  (
    g1278_p_spl_,
    g1278_p
  );


  buf

  (
    g1305_n_spl_,
    g1305_n
  );


  buf

  (
    g1304_n_spl_,
    g1304_n
  );


  buf

  (
    g1305_p_spl_,
    g1305_p
  );


  buf

  (
    g1304_p_spl_,
    g1304_p
  );


  buf

  (
    g1306_n_spl_,
    g1306_n
  );


  buf

  (
    g1306_p_spl_,
    g1306_p
  );


  buf

  (
    g1308_p_spl_,
    g1308_p
  );


  buf

  (
    g1303_n_spl_,
    g1303_n
  );


  buf

  (
    g1308_n_spl_,
    g1308_n
  );


  buf

  (
    g1303_p_spl_,
    g1303_p
  );


  buf

  (
    g1309_n_spl_,
    g1309_n
  );


  buf

  (
    g1309_p_spl_,
    g1309_p
  );


  buf

  (
    g1311_p_spl_,
    g1311_p
  );


  buf

  (
    g1302_n_spl_,
    g1302_n
  );


  buf

  (
    g1311_n_spl_,
    g1311_n
  );


  buf

  (
    g1302_p_spl_,
    g1302_p
  );


  buf

  (
    g1312_n_spl_,
    g1312_n
  );


  buf

  (
    g1312_p_spl_,
    g1312_p
  );


  buf

  (
    g1314_p_spl_,
    g1314_p
  );


  buf

  (
    g1301_n_spl_,
    g1301_n
  );


  buf

  (
    g1314_n_spl_,
    g1314_n
  );


  buf

  (
    g1301_p_spl_,
    g1301_p
  );


  buf

  (
    g1315_n_spl_,
    g1315_n
  );


  buf

  (
    g1315_p_spl_,
    g1315_p
  );


  buf

  (
    g1317_p_spl_,
    g1317_p
  );


  buf

  (
    g1300_n_spl_,
    g1300_n
  );


  buf

  (
    g1317_n_spl_,
    g1317_n
  );


  buf

  (
    g1300_p_spl_,
    g1300_p
  );


  buf

  (
    g1318_n_spl_,
    g1318_n
  );


  buf

  (
    g1318_p_spl_,
    g1318_p
  );


  buf

  (
    g1320_p_spl_,
    g1320_p
  );


  buf

  (
    g1299_n_spl_,
    g1299_n
  );


  buf

  (
    g1320_n_spl_,
    g1320_n
  );


  buf

  (
    g1299_p_spl_,
    g1299_p
  );


  buf

  (
    g1321_n_spl_,
    g1321_n
  );


  buf

  (
    g1321_p_spl_,
    g1321_p
  );


  buf

  (
    g1323_p_spl_,
    g1323_p
  );


  buf

  (
    g1298_n_spl_,
    g1298_n
  );


  buf

  (
    g1323_n_spl_,
    g1323_n
  );


  buf

  (
    g1298_p_spl_,
    g1298_p
  );


  buf

  (
    g1324_n_spl_,
    g1324_n
  );


  buf

  (
    g1324_p_spl_,
    g1324_p
  );


  buf

  (
    g1326_p_spl_,
    g1326_p
  );


  buf

  (
    g1297_n_spl_,
    g1297_n
  );


  buf

  (
    g1326_n_spl_,
    g1326_n
  );


  buf

  (
    g1297_p_spl_,
    g1297_p
  );


  buf

  (
    g1327_n_spl_,
    g1327_n
  );


  buf

  (
    g1327_p_spl_,
    g1327_p
  );


  buf

  (
    g1329_p_spl_,
    g1329_p
  );


  buf

  (
    g1296_n_spl_,
    g1296_n
  );


  buf

  (
    g1329_n_spl_,
    g1329_n
  );


  buf

  (
    g1296_p_spl_,
    g1296_p
  );


  buf

  (
    g1330_n_spl_,
    g1330_n
  );


  buf

  (
    g1330_p_spl_,
    g1330_p
  );


  buf

  (
    g1332_p_spl_,
    g1332_p
  );


  buf

  (
    g1295_n_spl_,
    g1295_n
  );


  buf

  (
    g1332_n_spl_,
    g1332_n
  );


  buf

  (
    g1295_p_spl_,
    g1295_p
  );


  buf

  (
    g1333_n_spl_,
    g1333_n
  );


  buf

  (
    g1333_p_spl_,
    g1333_p
  );


  buf

  (
    g1335_p_spl_,
    g1335_p
  );


  buf

  (
    g1294_n_spl_,
    g1294_n
  );


  buf

  (
    g1335_n_spl_,
    g1335_n
  );


  buf

  (
    g1294_p_spl_,
    g1294_p
  );


  buf

  (
    g1336_n_spl_,
    g1336_n
  );


  buf

  (
    g1336_p_spl_,
    g1336_p
  );


  buf

  (
    g1338_p_spl_,
    g1338_p
  );


  buf

  (
    g1293_n_spl_,
    g1293_n
  );


  buf

  (
    g1338_n_spl_,
    g1338_n
  );


  buf

  (
    g1293_p_spl_,
    g1293_p
  );


  buf

  (
    g1339_n_spl_,
    g1339_n
  );


  buf

  (
    g1339_p_spl_,
    g1339_p
  );


  buf

  (
    g1341_p_spl_,
    g1341_p
  );


  buf

  (
    g1292_n_spl_,
    g1292_n
  );


  buf

  (
    g1341_n_spl_,
    g1341_n
  );


  buf

  (
    g1292_p_spl_,
    g1292_p
  );


  buf

  (
    g1342_n_spl_,
    g1342_n
  );


  buf

  (
    g1342_p_spl_,
    g1342_p
  );


  buf

  (
    g1344_p_spl_,
    g1344_p
  );


  buf

  (
    g1291_n_spl_,
    g1291_n
  );


  buf

  (
    g1344_n_spl_,
    g1344_n
  );


  buf

  (
    g1291_p_spl_,
    g1291_p
  );


  buf

  (
    g1345_n_spl_,
    g1345_n
  );


  buf

  (
    g1345_p_spl_,
    g1345_p
  );


  buf

  (
    g1347_p_spl_,
    g1347_p
  );


  buf

  (
    g1290_n_spl_,
    g1290_n
  );


  buf

  (
    g1347_n_spl_,
    g1347_n
  );


  buf

  (
    g1290_p_spl_,
    g1290_p
  );


  buf

  (
    g1348_n_spl_,
    g1348_n
  );


  buf

  (
    g1348_p_spl_,
    g1348_p
  );


  buf

  (
    g1350_p_spl_,
    g1350_p
  );


  buf

  (
    g1289_n_spl_,
    g1289_n
  );


  buf

  (
    g1350_n_spl_,
    g1350_n
  );


  buf

  (
    g1289_p_spl_,
    g1289_p
  );


  buf

  (
    g1351_n_spl_,
    g1351_n
  );


  buf

  (
    g1351_p_spl_,
    g1351_p
  );


  buf

  (
    g1353_p_spl_,
    g1353_p
  );


  buf

  (
    g1288_n_spl_,
    g1288_n
  );


  buf

  (
    g1353_n_spl_,
    g1353_n
  );


  buf

  (
    g1288_p_spl_,
    g1288_p
  );


  buf

  (
    g1354_n_spl_,
    g1354_n
  );


  buf

  (
    g1354_p_spl_,
    g1354_p
  );


  buf

  (
    g1356_p_spl_,
    g1356_p
  );


  buf

  (
    g1287_n_spl_,
    g1287_n
  );


  buf

  (
    g1356_n_spl_,
    g1356_n
  );


  buf

  (
    g1287_p_spl_,
    g1287_p
  );


  buf

  (
    g1357_n_spl_,
    g1357_n
  );


  buf

  (
    g1357_p_spl_,
    g1357_p
  );


  buf

  (
    g1359_p_spl_,
    g1359_p
  );


  buf

  (
    g1286_n_spl_,
    g1286_n
  );


  buf

  (
    g1359_n_spl_,
    g1359_n
  );


  buf

  (
    g1286_p_spl_,
    g1286_p
  );


  buf

  (
    g1360_n_spl_,
    g1360_n
  );


  buf

  (
    g1360_p_spl_,
    g1360_p
  );


  buf

  (
    g1362_p_spl_,
    g1362_p
  );


  buf

  (
    g1285_n_spl_,
    g1285_n
  );


  buf

  (
    g1362_n_spl_,
    g1362_n
  );


  buf

  (
    g1285_p_spl_,
    g1285_p
  );


  buf

  (
    g1363_n_spl_,
    g1363_n
  );


  buf

  (
    g1363_p_spl_,
    g1363_p
  );


  buf

  (
    g1365_p_spl_,
    g1365_p
  );


  buf

  (
    g1284_n_spl_,
    g1284_n
  );


  buf

  (
    g1365_n_spl_,
    g1365_n
  );


  buf

  (
    g1284_p_spl_,
    g1284_p
  );


  buf

  (
    g1366_n_spl_,
    g1366_n
  );


  buf

  (
    g1366_p_spl_,
    g1366_p
  );


  buf

  (
    g1368_p_spl_,
    g1368_p
  );


  buf

  (
    g1283_n_spl_,
    g1283_n
  );


  buf

  (
    g1368_n_spl_,
    g1368_n
  );


  buf

  (
    g1283_p_spl_,
    g1283_p
  );


  buf

  (
    g1369_n_spl_,
    g1369_n
  );


  buf

  (
    g1369_p_spl_,
    g1369_p
  );


  buf

  (
    g1371_p_spl_,
    g1371_p
  );


  buf

  (
    g1282_n_spl_,
    g1282_n
  );


  buf

  (
    g1371_n_spl_,
    g1371_n
  );


  buf

  (
    g1282_p_spl_,
    g1282_p
  );


  buf

  (
    g1372_n_spl_,
    g1372_n
  );


  buf

  (
    g1372_p_spl_,
    g1372_p
  );


  buf

  (
    g1374_n_spl_,
    g1374_n
  );


  buf

  (
    g1281_p_spl_,
    g1281_p
  );


  buf

  (
    g1375_p_spl_,
    g1375_p
  );


  buf

  (
    g1400_n_spl_,
    g1400_n
  );


  buf

  (
    g1399_n_spl_,
    g1399_n
  );


  buf

  (
    g1400_p_spl_,
    g1400_p
  );


  buf

  (
    g1399_p_spl_,
    g1399_p
  );


  buf

  (
    g1401_n_spl_,
    g1401_n
  );


  buf

  (
    g1401_p_spl_,
    g1401_p
  );


  buf

  (
    g1403_p_spl_,
    g1403_p
  );


  buf

  (
    g1398_n_spl_,
    g1398_n
  );


  buf

  (
    g1403_n_spl_,
    g1403_n
  );


  buf

  (
    g1398_p_spl_,
    g1398_p
  );


  buf

  (
    g1404_n_spl_,
    g1404_n
  );


  buf

  (
    g1404_p_spl_,
    g1404_p
  );


  buf

  (
    g1406_p_spl_,
    g1406_p
  );


  buf

  (
    g1397_n_spl_,
    g1397_n
  );


  buf

  (
    g1406_n_spl_,
    g1406_n
  );


  buf

  (
    g1397_p_spl_,
    g1397_p
  );


  buf

  (
    g1407_n_spl_,
    g1407_n
  );


  buf

  (
    g1407_p_spl_,
    g1407_p
  );


  buf

  (
    g1409_p_spl_,
    g1409_p
  );


  buf

  (
    g1396_n_spl_,
    g1396_n
  );


  buf

  (
    g1409_n_spl_,
    g1409_n
  );


  buf

  (
    g1396_p_spl_,
    g1396_p
  );


  buf

  (
    g1410_n_spl_,
    g1410_n
  );


  buf

  (
    g1410_p_spl_,
    g1410_p
  );


  buf

  (
    g1412_p_spl_,
    g1412_p
  );


  buf

  (
    g1395_n_spl_,
    g1395_n
  );


  buf

  (
    g1412_n_spl_,
    g1412_n
  );


  buf

  (
    g1395_p_spl_,
    g1395_p
  );


  buf

  (
    g1413_n_spl_,
    g1413_n
  );


  buf

  (
    g1413_p_spl_,
    g1413_p
  );


  buf

  (
    g1415_p_spl_,
    g1415_p
  );


  buf

  (
    g1394_n_spl_,
    g1394_n
  );


  buf

  (
    g1415_n_spl_,
    g1415_n
  );


  buf

  (
    g1394_p_spl_,
    g1394_p
  );


  buf

  (
    g1416_n_spl_,
    g1416_n
  );


  buf

  (
    g1416_p_spl_,
    g1416_p
  );


  buf

  (
    g1418_p_spl_,
    g1418_p
  );


  buf

  (
    g1393_n_spl_,
    g1393_n
  );


  buf

  (
    g1418_n_spl_,
    g1418_n
  );


  buf

  (
    g1393_p_spl_,
    g1393_p
  );


  buf

  (
    g1419_n_spl_,
    g1419_n
  );


  buf

  (
    g1419_p_spl_,
    g1419_p
  );


  buf

  (
    g1421_p_spl_,
    g1421_p
  );


  buf

  (
    g1392_n_spl_,
    g1392_n
  );


  buf

  (
    g1421_n_spl_,
    g1421_n
  );


  buf

  (
    g1392_p_spl_,
    g1392_p
  );


  buf

  (
    g1422_n_spl_,
    g1422_n
  );


  buf

  (
    g1422_p_spl_,
    g1422_p
  );


  buf

  (
    g1424_p_spl_,
    g1424_p
  );


  buf

  (
    g1391_n_spl_,
    g1391_n
  );


  buf

  (
    g1424_n_spl_,
    g1424_n
  );


  buf

  (
    g1391_p_spl_,
    g1391_p
  );


  buf

  (
    g1425_n_spl_,
    g1425_n
  );


  buf

  (
    g1425_p_spl_,
    g1425_p
  );


  buf

  (
    g1427_p_spl_,
    g1427_p
  );


  buf

  (
    g1390_n_spl_,
    g1390_n
  );


  buf

  (
    g1427_n_spl_,
    g1427_n
  );


  buf

  (
    g1390_p_spl_,
    g1390_p
  );


  buf

  (
    g1428_n_spl_,
    g1428_n
  );


  buf

  (
    g1428_p_spl_,
    g1428_p
  );


  buf

  (
    g1430_p_spl_,
    g1430_p
  );


  buf

  (
    g1389_n_spl_,
    g1389_n
  );


  buf

  (
    g1430_n_spl_,
    g1430_n
  );


  buf

  (
    g1389_p_spl_,
    g1389_p
  );


  buf

  (
    g1431_n_spl_,
    g1431_n
  );


  buf

  (
    g1431_p_spl_,
    g1431_p
  );


  buf

  (
    g1433_p_spl_,
    g1433_p
  );


  buf

  (
    g1388_n_spl_,
    g1388_n
  );


  buf

  (
    g1433_n_spl_,
    g1433_n
  );


  buf

  (
    g1388_p_spl_,
    g1388_p
  );


  buf

  (
    g1434_n_spl_,
    g1434_n
  );


  buf

  (
    g1434_p_spl_,
    g1434_p
  );


  buf

  (
    g1436_p_spl_,
    g1436_p
  );


  buf

  (
    g1387_n_spl_,
    g1387_n
  );


  buf

  (
    g1436_n_spl_,
    g1436_n
  );


  buf

  (
    g1387_p_spl_,
    g1387_p
  );


  buf

  (
    g1437_n_spl_,
    g1437_n
  );


  buf

  (
    g1437_p_spl_,
    g1437_p
  );


  buf

  (
    g1439_p_spl_,
    g1439_p
  );


  buf

  (
    g1386_n_spl_,
    g1386_n
  );


  buf

  (
    g1439_n_spl_,
    g1439_n
  );


  buf

  (
    g1386_p_spl_,
    g1386_p
  );


  buf

  (
    g1440_n_spl_,
    g1440_n
  );


  buf

  (
    g1440_p_spl_,
    g1440_p
  );


  buf

  (
    g1442_p_spl_,
    g1442_p
  );


  buf

  (
    g1385_n_spl_,
    g1385_n
  );


  buf

  (
    g1442_n_spl_,
    g1442_n
  );


  buf

  (
    g1385_p_spl_,
    g1385_p
  );


  buf

  (
    g1443_n_spl_,
    g1443_n
  );


  buf

  (
    g1443_p_spl_,
    g1443_p
  );


  buf

  (
    g1445_p_spl_,
    g1445_p
  );


  buf

  (
    g1384_n_spl_,
    g1384_n
  );


  buf

  (
    g1445_n_spl_,
    g1445_n
  );


  buf

  (
    g1384_p_spl_,
    g1384_p
  );


  buf

  (
    g1446_n_spl_,
    g1446_n
  );


  buf

  (
    g1446_p_spl_,
    g1446_p
  );


  buf

  (
    g1448_p_spl_,
    g1448_p
  );


  buf

  (
    g1383_n_spl_,
    g1383_n
  );


  buf

  (
    g1448_n_spl_,
    g1448_n
  );


  buf

  (
    g1383_p_spl_,
    g1383_p
  );


  buf

  (
    g1449_n_spl_,
    g1449_n
  );


  buf

  (
    g1449_p_spl_,
    g1449_p
  );


  buf

  (
    g1451_p_spl_,
    g1451_p
  );


  buf

  (
    g1382_n_spl_,
    g1382_n
  );


  buf

  (
    g1451_n_spl_,
    g1451_n
  );


  buf

  (
    g1382_p_spl_,
    g1382_p
  );


  buf

  (
    g1452_n_spl_,
    g1452_n
  );


  buf

  (
    g1452_p_spl_,
    g1452_p
  );


  buf

  (
    g1454_p_spl_,
    g1454_p
  );


  buf

  (
    g1381_n_spl_,
    g1381_n
  );


  buf

  (
    g1454_n_spl_,
    g1454_n
  );


  buf

  (
    g1381_p_spl_,
    g1381_p
  );


  buf

  (
    g1455_n_spl_,
    g1455_n
  );


  buf

  (
    g1455_p_spl_,
    g1455_p
  );


  buf

  (
    g1457_p_spl_,
    g1457_p
  );


  buf

  (
    g1380_n_spl_,
    g1380_n
  );


  buf

  (
    g1457_n_spl_,
    g1457_n
  );


  buf

  (
    g1380_p_spl_,
    g1380_p
  );


  buf

  (
    g1458_n_spl_,
    g1458_n
  );


  buf

  (
    g1458_p_spl_,
    g1458_p
  );


  buf

  (
    g1460_p_spl_,
    g1460_p
  );


  buf

  (
    g1379_n_spl_,
    g1379_n
  );


  buf

  (
    g1460_n_spl_,
    g1460_n
  );


  buf

  (
    g1379_p_spl_,
    g1379_p
  );


  buf

  (
    g1461_n_spl_,
    g1461_n
  );


  buf

  (
    g1461_p_spl_,
    g1461_p
  );


  buf

  (
    g1463_n_spl_,
    g1463_n
  );


  buf

  (
    g1378_p_spl_,
    g1378_p
  );


  buf

  (
    g1464_p_spl_,
    g1464_p
  );


  buf

  (
    g1487_n_spl_,
    g1487_n
  );


  buf

  (
    g1486_n_spl_,
    g1486_n
  );


  buf

  (
    g1487_p_spl_,
    g1487_p
  );


  buf

  (
    g1486_p_spl_,
    g1486_p
  );


  buf

  (
    g1488_n_spl_,
    g1488_n
  );


  buf

  (
    g1488_p_spl_,
    g1488_p
  );


  buf

  (
    g1490_p_spl_,
    g1490_p
  );


  buf

  (
    g1485_n_spl_,
    g1485_n
  );


  buf

  (
    g1490_n_spl_,
    g1490_n
  );


  buf

  (
    g1485_p_spl_,
    g1485_p
  );


  buf

  (
    g1491_n_spl_,
    g1491_n
  );


  buf

  (
    g1491_p_spl_,
    g1491_p
  );


  buf

  (
    g1493_p_spl_,
    g1493_p
  );


  buf

  (
    g1484_n_spl_,
    g1484_n
  );


  buf

  (
    g1493_n_spl_,
    g1493_n
  );


  buf

  (
    g1484_p_spl_,
    g1484_p
  );


  buf

  (
    g1494_n_spl_,
    g1494_n
  );


  buf

  (
    g1494_p_spl_,
    g1494_p
  );


  buf

  (
    g1496_p_spl_,
    g1496_p
  );


  buf

  (
    g1483_n_spl_,
    g1483_n
  );


  buf

  (
    g1496_n_spl_,
    g1496_n
  );


  buf

  (
    g1483_p_spl_,
    g1483_p
  );


  buf

  (
    g1497_n_spl_,
    g1497_n
  );


  buf

  (
    g1497_p_spl_,
    g1497_p
  );


  buf

  (
    g1499_p_spl_,
    g1499_p
  );


  buf

  (
    g1482_n_spl_,
    g1482_n
  );


  buf

  (
    g1499_n_spl_,
    g1499_n
  );


  buf

  (
    g1482_p_spl_,
    g1482_p
  );


  buf

  (
    g1500_n_spl_,
    g1500_n
  );


  buf

  (
    g1500_p_spl_,
    g1500_p
  );


  buf

  (
    g1502_p_spl_,
    g1502_p
  );


  buf

  (
    g1481_n_spl_,
    g1481_n
  );


  buf

  (
    g1502_n_spl_,
    g1502_n
  );


  buf

  (
    g1481_p_spl_,
    g1481_p
  );


  buf

  (
    g1503_n_spl_,
    g1503_n
  );


  buf

  (
    g1503_p_spl_,
    g1503_p
  );


  buf

  (
    g1505_p_spl_,
    g1505_p
  );


  buf

  (
    g1480_n_spl_,
    g1480_n
  );


  buf

  (
    g1505_n_spl_,
    g1505_n
  );


  buf

  (
    g1480_p_spl_,
    g1480_p
  );


  buf

  (
    g1506_n_spl_,
    g1506_n
  );


  buf

  (
    g1506_p_spl_,
    g1506_p
  );


  buf

  (
    g1508_p_spl_,
    g1508_p
  );


  buf

  (
    g1479_n_spl_,
    g1479_n
  );


  buf

  (
    g1508_n_spl_,
    g1508_n
  );


  buf

  (
    g1479_p_spl_,
    g1479_p
  );


  buf

  (
    g1509_n_spl_,
    g1509_n
  );


  buf

  (
    g1509_p_spl_,
    g1509_p
  );


  buf

  (
    g1511_p_spl_,
    g1511_p
  );


  buf

  (
    g1478_n_spl_,
    g1478_n
  );


  buf

  (
    g1511_n_spl_,
    g1511_n
  );


  buf

  (
    g1478_p_spl_,
    g1478_p
  );


  buf

  (
    g1512_n_spl_,
    g1512_n
  );


  buf

  (
    g1512_p_spl_,
    g1512_p
  );


  buf

  (
    g1514_p_spl_,
    g1514_p
  );


  buf

  (
    g1477_n_spl_,
    g1477_n
  );


  buf

  (
    g1514_n_spl_,
    g1514_n
  );


  buf

  (
    g1477_p_spl_,
    g1477_p
  );


  buf

  (
    g1515_n_spl_,
    g1515_n
  );


  buf

  (
    g1515_p_spl_,
    g1515_p
  );


  buf

  (
    g1517_p_spl_,
    g1517_p
  );


  buf

  (
    g1476_n_spl_,
    g1476_n
  );


  buf

  (
    g1517_n_spl_,
    g1517_n
  );


  buf

  (
    g1476_p_spl_,
    g1476_p
  );


  buf

  (
    g1518_n_spl_,
    g1518_n
  );


  buf

  (
    g1518_p_spl_,
    g1518_p
  );


  buf

  (
    g1520_p_spl_,
    g1520_p
  );


  buf

  (
    g1475_n_spl_,
    g1475_n
  );


  buf

  (
    g1520_n_spl_,
    g1520_n
  );


  buf

  (
    g1475_p_spl_,
    g1475_p
  );


  buf

  (
    g1521_n_spl_,
    g1521_n
  );


  buf

  (
    g1521_p_spl_,
    g1521_p
  );


  buf

  (
    g1523_p_spl_,
    g1523_p
  );


  buf

  (
    g1474_n_spl_,
    g1474_n
  );


  buf

  (
    g1523_n_spl_,
    g1523_n
  );


  buf

  (
    g1474_p_spl_,
    g1474_p
  );


  buf

  (
    g1524_n_spl_,
    g1524_n
  );


  buf

  (
    g1524_p_spl_,
    g1524_p
  );


  buf

  (
    g1526_p_spl_,
    g1526_p
  );


  buf

  (
    g1473_n_spl_,
    g1473_n
  );


  buf

  (
    g1526_n_spl_,
    g1526_n
  );


  buf

  (
    g1473_p_spl_,
    g1473_p
  );


  buf

  (
    g1527_n_spl_,
    g1527_n
  );


  buf

  (
    g1527_p_spl_,
    g1527_p
  );


  buf

  (
    g1529_p_spl_,
    g1529_p
  );


  buf

  (
    g1472_n_spl_,
    g1472_n
  );


  buf

  (
    g1529_n_spl_,
    g1529_n
  );


  buf

  (
    g1472_p_spl_,
    g1472_p
  );


  buf

  (
    g1530_n_spl_,
    g1530_n
  );


  buf

  (
    g1530_p_spl_,
    g1530_p
  );


  buf

  (
    g1532_p_spl_,
    g1532_p
  );


  buf

  (
    g1471_n_spl_,
    g1471_n
  );


  buf

  (
    g1532_n_spl_,
    g1532_n
  );


  buf

  (
    g1471_p_spl_,
    g1471_p
  );


  buf

  (
    g1533_n_spl_,
    g1533_n
  );


  buf

  (
    g1533_p_spl_,
    g1533_p
  );


  buf

  (
    g1535_p_spl_,
    g1535_p
  );


  buf

  (
    g1470_n_spl_,
    g1470_n
  );


  buf

  (
    g1535_n_spl_,
    g1535_n
  );


  buf

  (
    g1470_p_spl_,
    g1470_p
  );


  buf

  (
    g1536_n_spl_,
    g1536_n
  );


  buf

  (
    g1536_p_spl_,
    g1536_p
  );


  buf

  (
    g1538_p_spl_,
    g1538_p
  );


  buf

  (
    g1469_n_spl_,
    g1469_n
  );


  buf

  (
    g1538_n_spl_,
    g1538_n
  );


  buf

  (
    g1469_p_spl_,
    g1469_p
  );


  buf

  (
    g1539_n_spl_,
    g1539_n
  );


  buf

  (
    g1539_p_spl_,
    g1539_p
  );


  buf

  (
    g1541_p_spl_,
    g1541_p
  );


  buf

  (
    g1468_n_spl_,
    g1468_n
  );


  buf

  (
    g1541_n_spl_,
    g1541_n
  );


  buf

  (
    g1468_p_spl_,
    g1468_p
  );


  buf

  (
    g1542_n_spl_,
    g1542_n
  );


  buf

  (
    g1542_p_spl_,
    g1542_p
  );


  buf

  (
    g1544_n_spl_,
    g1544_n
  );


  buf

  (
    g1467_p_spl_,
    g1467_p
  );


  buf

  (
    g1545_p_spl_,
    g1545_p
  );


  buf

  (
    g1566_n_spl_,
    g1566_n
  );


  buf

  (
    g1565_n_spl_,
    g1565_n
  );


  buf

  (
    g1566_p_spl_,
    g1566_p
  );


  buf

  (
    g1565_p_spl_,
    g1565_p
  );


  buf

  (
    g1567_n_spl_,
    g1567_n
  );


  buf

  (
    g1567_p_spl_,
    g1567_p
  );


  buf

  (
    g1569_p_spl_,
    g1569_p
  );


  buf

  (
    g1564_n_spl_,
    g1564_n
  );


  buf

  (
    g1569_n_spl_,
    g1569_n
  );


  buf

  (
    g1564_p_spl_,
    g1564_p
  );


  buf

  (
    g1570_n_spl_,
    g1570_n
  );


  buf

  (
    g1570_p_spl_,
    g1570_p
  );


  buf

  (
    g1572_p_spl_,
    g1572_p
  );


  buf

  (
    g1563_n_spl_,
    g1563_n
  );


  buf

  (
    g1572_n_spl_,
    g1572_n
  );


  buf

  (
    g1563_p_spl_,
    g1563_p
  );


  buf

  (
    g1573_n_spl_,
    g1573_n
  );


  buf

  (
    g1573_p_spl_,
    g1573_p
  );


  buf

  (
    g1575_p_spl_,
    g1575_p
  );


  buf

  (
    g1562_n_spl_,
    g1562_n
  );


  buf

  (
    g1575_n_spl_,
    g1575_n
  );


  buf

  (
    g1562_p_spl_,
    g1562_p
  );


  buf

  (
    g1576_n_spl_,
    g1576_n
  );


  buf

  (
    g1576_p_spl_,
    g1576_p
  );


  buf

  (
    g1578_p_spl_,
    g1578_p
  );


  buf

  (
    g1561_n_spl_,
    g1561_n
  );


  buf

  (
    g1578_n_spl_,
    g1578_n
  );


  buf

  (
    g1561_p_spl_,
    g1561_p
  );


  buf

  (
    g1579_n_spl_,
    g1579_n
  );


  buf

  (
    g1579_p_spl_,
    g1579_p
  );


  buf

  (
    g1581_p_spl_,
    g1581_p
  );


  buf

  (
    g1560_n_spl_,
    g1560_n
  );


  buf

  (
    g1581_n_spl_,
    g1581_n
  );


  buf

  (
    g1560_p_spl_,
    g1560_p
  );


  buf

  (
    g1582_n_spl_,
    g1582_n
  );


  buf

  (
    g1582_p_spl_,
    g1582_p
  );


  buf

  (
    g1584_p_spl_,
    g1584_p
  );


  buf

  (
    g1559_n_spl_,
    g1559_n
  );


  buf

  (
    g1584_n_spl_,
    g1584_n
  );


  buf

  (
    g1559_p_spl_,
    g1559_p
  );


  buf

  (
    g1585_n_spl_,
    g1585_n
  );


  buf

  (
    g1585_p_spl_,
    g1585_p
  );


  buf

  (
    g1587_p_spl_,
    g1587_p
  );


  buf

  (
    g1558_n_spl_,
    g1558_n
  );


  buf

  (
    g1587_n_spl_,
    g1587_n
  );


  buf

  (
    g1558_p_spl_,
    g1558_p
  );


  buf

  (
    g1588_n_spl_,
    g1588_n
  );


  buf

  (
    g1588_p_spl_,
    g1588_p
  );


  buf

  (
    g1590_p_spl_,
    g1590_p
  );


  buf

  (
    g1557_n_spl_,
    g1557_n
  );


  buf

  (
    g1590_n_spl_,
    g1590_n
  );


  buf

  (
    g1557_p_spl_,
    g1557_p
  );


  buf

  (
    g1591_n_spl_,
    g1591_n
  );


  buf

  (
    g1591_p_spl_,
    g1591_p
  );


  buf

  (
    g1593_p_spl_,
    g1593_p
  );


  buf

  (
    g1556_n_spl_,
    g1556_n
  );


  buf

  (
    g1593_n_spl_,
    g1593_n
  );


  buf

  (
    g1556_p_spl_,
    g1556_p
  );


  buf

  (
    g1594_n_spl_,
    g1594_n
  );


  buf

  (
    g1594_p_spl_,
    g1594_p
  );


  buf

  (
    g1596_p_spl_,
    g1596_p
  );


  buf

  (
    g1555_n_spl_,
    g1555_n
  );


  buf

  (
    g1596_n_spl_,
    g1596_n
  );


  buf

  (
    g1555_p_spl_,
    g1555_p
  );


  buf

  (
    g1597_n_spl_,
    g1597_n
  );


  buf

  (
    g1597_p_spl_,
    g1597_p
  );


  buf

  (
    g1599_p_spl_,
    g1599_p
  );


  buf

  (
    g1554_n_spl_,
    g1554_n
  );


  buf

  (
    g1599_n_spl_,
    g1599_n
  );


  buf

  (
    g1554_p_spl_,
    g1554_p
  );


  buf

  (
    g1600_n_spl_,
    g1600_n
  );


  buf

  (
    g1600_p_spl_,
    g1600_p
  );


  buf

  (
    g1602_p_spl_,
    g1602_p
  );


  buf

  (
    g1553_n_spl_,
    g1553_n
  );


  buf

  (
    g1602_n_spl_,
    g1602_n
  );


  buf

  (
    g1553_p_spl_,
    g1553_p
  );


  buf

  (
    g1603_n_spl_,
    g1603_n
  );


  buf

  (
    g1603_p_spl_,
    g1603_p
  );


  buf

  (
    g1605_p_spl_,
    g1605_p
  );


  buf

  (
    g1552_n_spl_,
    g1552_n
  );


  buf

  (
    g1605_n_spl_,
    g1605_n
  );


  buf

  (
    g1552_p_spl_,
    g1552_p
  );


  buf

  (
    g1606_n_spl_,
    g1606_n
  );


  buf

  (
    g1606_p_spl_,
    g1606_p
  );


  buf

  (
    g1608_p_spl_,
    g1608_p
  );


  buf

  (
    g1551_n_spl_,
    g1551_n
  );


  buf

  (
    g1608_n_spl_,
    g1608_n
  );


  buf

  (
    g1551_p_spl_,
    g1551_p
  );


  buf

  (
    g1609_n_spl_,
    g1609_n
  );


  buf

  (
    g1609_p_spl_,
    g1609_p
  );


  buf

  (
    g1611_p_spl_,
    g1611_p
  );


  buf

  (
    g1550_n_spl_,
    g1550_n
  );


  buf

  (
    g1611_n_spl_,
    g1611_n
  );


  buf

  (
    g1550_p_spl_,
    g1550_p
  );


  buf

  (
    g1612_n_spl_,
    g1612_n
  );


  buf

  (
    g1612_p_spl_,
    g1612_p
  );


  buf

  (
    g1614_p_spl_,
    g1614_p
  );


  buf

  (
    g1549_n_spl_,
    g1549_n
  );


  buf

  (
    g1614_n_spl_,
    g1614_n
  );


  buf

  (
    g1549_p_spl_,
    g1549_p
  );


  buf

  (
    g1615_n_spl_,
    g1615_n
  );


  buf

  (
    g1615_p_spl_,
    g1615_p
  );


  buf

  (
    g1617_n_spl_,
    g1617_n
  );


  buf

  (
    g1548_p_spl_,
    g1548_p
  );


  buf

  (
    g1618_p_spl_,
    g1618_p
  );


  buf

  (
    g1637_n_spl_,
    g1637_n
  );


  buf

  (
    g1636_n_spl_,
    g1636_n
  );


  buf

  (
    g1637_p_spl_,
    g1637_p
  );


  buf

  (
    g1636_p_spl_,
    g1636_p
  );


  buf

  (
    g1638_n_spl_,
    g1638_n
  );


  buf

  (
    g1638_p_spl_,
    g1638_p
  );


  buf

  (
    g1640_p_spl_,
    g1640_p
  );


  buf

  (
    g1635_n_spl_,
    g1635_n
  );


  buf

  (
    g1640_n_spl_,
    g1640_n
  );


  buf

  (
    g1635_p_spl_,
    g1635_p
  );


  buf

  (
    g1641_n_spl_,
    g1641_n
  );


  buf

  (
    g1641_p_spl_,
    g1641_p
  );


  buf

  (
    g1643_p_spl_,
    g1643_p
  );


  buf

  (
    g1634_n_spl_,
    g1634_n
  );


  buf

  (
    g1643_n_spl_,
    g1643_n
  );


  buf

  (
    g1634_p_spl_,
    g1634_p
  );


  buf

  (
    g1644_n_spl_,
    g1644_n
  );


  buf

  (
    g1644_p_spl_,
    g1644_p
  );


  buf

  (
    g1646_p_spl_,
    g1646_p
  );


  buf

  (
    g1633_n_spl_,
    g1633_n
  );


  buf

  (
    g1646_n_spl_,
    g1646_n
  );


  buf

  (
    g1633_p_spl_,
    g1633_p
  );


  buf

  (
    g1647_n_spl_,
    g1647_n
  );


  buf

  (
    g1647_p_spl_,
    g1647_p
  );


  buf

  (
    g1649_p_spl_,
    g1649_p
  );


  buf

  (
    g1632_n_spl_,
    g1632_n
  );


  buf

  (
    g1649_n_spl_,
    g1649_n
  );


  buf

  (
    g1632_p_spl_,
    g1632_p
  );


  buf

  (
    g1650_n_spl_,
    g1650_n
  );


  buf

  (
    g1650_p_spl_,
    g1650_p
  );


  buf

  (
    g1652_p_spl_,
    g1652_p
  );


  buf

  (
    g1631_n_spl_,
    g1631_n
  );


  buf

  (
    g1652_n_spl_,
    g1652_n
  );


  buf

  (
    g1631_p_spl_,
    g1631_p
  );


  buf

  (
    g1653_n_spl_,
    g1653_n
  );


  buf

  (
    g1653_p_spl_,
    g1653_p
  );


  buf

  (
    g1655_p_spl_,
    g1655_p
  );


  buf

  (
    g1630_n_spl_,
    g1630_n
  );


  buf

  (
    g1655_n_spl_,
    g1655_n
  );


  buf

  (
    g1630_p_spl_,
    g1630_p
  );


  buf

  (
    g1656_n_spl_,
    g1656_n
  );


  buf

  (
    g1656_p_spl_,
    g1656_p
  );


  buf

  (
    g1658_p_spl_,
    g1658_p
  );


  buf

  (
    g1629_n_spl_,
    g1629_n
  );


  buf

  (
    g1658_n_spl_,
    g1658_n
  );


  buf

  (
    g1629_p_spl_,
    g1629_p
  );


  buf

  (
    g1659_n_spl_,
    g1659_n
  );


  buf

  (
    g1659_p_spl_,
    g1659_p
  );


  buf

  (
    g1661_p_spl_,
    g1661_p
  );


  buf

  (
    g1628_n_spl_,
    g1628_n
  );


  buf

  (
    g1661_n_spl_,
    g1661_n
  );


  buf

  (
    g1628_p_spl_,
    g1628_p
  );


  buf

  (
    g1662_n_spl_,
    g1662_n
  );


  buf

  (
    g1662_p_spl_,
    g1662_p
  );


  buf

  (
    g1664_p_spl_,
    g1664_p
  );


  buf

  (
    g1627_n_spl_,
    g1627_n
  );


  buf

  (
    g1664_n_spl_,
    g1664_n
  );


  buf

  (
    g1627_p_spl_,
    g1627_p
  );


  buf

  (
    g1665_n_spl_,
    g1665_n
  );


  buf

  (
    g1665_p_spl_,
    g1665_p
  );


  buf

  (
    g1667_p_spl_,
    g1667_p
  );


  buf

  (
    g1626_n_spl_,
    g1626_n
  );


  buf

  (
    g1667_n_spl_,
    g1667_n
  );


  buf

  (
    g1626_p_spl_,
    g1626_p
  );


  buf

  (
    g1668_n_spl_,
    g1668_n
  );


  buf

  (
    g1668_p_spl_,
    g1668_p
  );


  buf

  (
    g1670_p_spl_,
    g1670_p
  );


  buf

  (
    g1625_n_spl_,
    g1625_n
  );


  buf

  (
    g1670_n_spl_,
    g1670_n
  );


  buf

  (
    g1625_p_spl_,
    g1625_p
  );


  buf

  (
    g1671_n_spl_,
    g1671_n
  );


  buf

  (
    g1671_p_spl_,
    g1671_p
  );


  buf

  (
    g1673_p_spl_,
    g1673_p
  );


  buf

  (
    g1624_n_spl_,
    g1624_n
  );


  buf

  (
    g1673_n_spl_,
    g1673_n
  );


  buf

  (
    g1624_p_spl_,
    g1624_p
  );


  buf

  (
    g1674_n_spl_,
    g1674_n
  );


  buf

  (
    g1674_p_spl_,
    g1674_p
  );


  buf

  (
    g1676_p_spl_,
    g1676_p
  );


  buf

  (
    g1623_n_spl_,
    g1623_n
  );


  buf

  (
    g1676_n_spl_,
    g1676_n
  );


  buf

  (
    g1623_p_spl_,
    g1623_p
  );


  buf

  (
    g1677_n_spl_,
    g1677_n
  );


  buf

  (
    g1677_p_spl_,
    g1677_p
  );


  buf

  (
    g1679_p_spl_,
    g1679_p
  );


  buf

  (
    g1622_n_spl_,
    g1622_n
  );


  buf

  (
    g1679_n_spl_,
    g1679_n
  );


  buf

  (
    g1622_p_spl_,
    g1622_p
  );


  buf

  (
    g1680_n_spl_,
    g1680_n
  );


  buf

  (
    g1680_p_spl_,
    g1680_p
  );


  buf

  (
    g1682_n_spl_,
    g1682_n
  );


  buf

  (
    g1621_p_spl_,
    g1621_p
  );


  buf

  (
    g1683_p_spl_,
    g1683_p
  );


  buf

  (
    g1700_n_spl_,
    g1700_n
  );


  buf

  (
    g1699_n_spl_,
    g1699_n
  );


  buf

  (
    g1700_p_spl_,
    g1700_p
  );


  buf

  (
    g1699_p_spl_,
    g1699_p
  );


  buf

  (
    g1701_n_spl_,
    g1701_n
  );


  buf

  (
    g1701_p_spl_,
    g1701_p
  );


  buf

  (
    g1703_p_spl_,
    g1703_p
  );


  buf

  (
    g1698_n_spl_,
    g1698_n
  );


  buf

  (
    g1703_n_spl_,
    g1703_n
  );


  buf

  (
    g1698_p_spl_,
    g1698_p
  );


  buf

  (
    g1704_n_spl_,
    g1704_n
  );


  buf

  (
    g1704_p_spl_,
    g1704_p
  );


  buf

  (
    g1706_p_spl_,
    g1706_p
  );


  buf

  (
    g1697_n_spl_,
    g1697_n
  );


  buf

  (
    g1706_n_spl_,
    g1706_n
  );


  buf

  (
    g1697_p_spl_,
    g1697_p
  );


  buf

  (
    g1707_n_spl_,
    g1707_n
  );


  buf

  (
    g1707_p_spl_,
    g1707_p
  );


  buf

  (
    g1709_p_spl_,
    g1709_p
  );


  buf

  (
    g1696_n_spl_,
    g1696_n
  );


  buf

  (
    g1709_n_spl_,
    g1709_n
  );


  buf

  (
    g1696_p_spl_,
    g1696_p
  );


  buf

  (
    g1710_n_spl_,
    g1710_n
  );


  buf

  (
    g1710_p_spl_,
    g1710_p
  );


  buf

  (
    g1712_p_spl_,
    g1712_p
  );


  buf

  (
    g1695_n_spl_,
    g1695_n
  );


  buf

  (
    g1712_n_spl_,
    g1712_n
  );


  buf

  (
    g1695_p_spl_,
    g1695_p
  );


  buf

  (
    g1713_n_spl_,
    g1713_n
  );


  buf

  (
    g1713_p_spl_,
    g1713_p
  );


  buf

  (
    g1715_p_spl_,
    g1715_p
  );


  buf

  (
    g1694_n_spl_,
    g1694_n
  );


  buf

  (
    g1715_n_spl_,
    g1715_n
  );


  buf

  (
    g1694_p_spl_,
    g1694_p
  );


  buf

  (
    g1716_n_spl_,
    g1716_n
  );


  buf

  (
    g1716_p_spl_,
    g1716_p
  );


  buf

  (
    g1718_p_spl_,
    g1718_p
  );


  buf

  (
    g1693_n_spl_,
    g1693_n
  );


  buf

  (
    g1718_n_spl_,
    g1718_n
  );


  buf

  (
    g1693_p_spl_,
    g1693_p
  );


  buf

  (
    g1719_n_spl_,
    g1719_n
  );


  buf

  (
    g1719_p_spl_,
    g1719_p
  );


  buf

  (
    g1721_p_spl_,
    g1721_p
  );


  buf

  (
    g1692_n_spl_,
    g1692_n
  );


  buf

  (
    g1721_n_spl_,
    g1721_n
  );


  buf

  (
    g1692_p_spl_,
    g1692_p
  );


  buf

  (
    g1722_n_spl_,
    g1722_n
  );


  buf

  (
    g1722_p_spl_,
    g1722_p
  );


  buf

  (
    g1724_p_spl_,
    g1724_p
  );


  buf

  (
    g1691_n_spl_,
    g1691_n
  );


  buf

  (
    g1724_n_spl_,
    g1724_n
  );


  buf

  (
    g1691_p_spl_,
    g1691_p
  );


  buf

  (
    g1725_n_spl_,
    g1725_n
  );


  buf

  (
    g1725_p_spl_,
    g1725_p
  );


  buf

  (
    g1727_p_spl_,
    g1727_p
  );


  buf

  (
    g1690_n_spl_,
    g1690_n
  );


  buf

  (
    g1727_n_spl_,
    g1727_n
  );


  buf

  (
    g1690_p_spl_,
    g1690_p
  );


  buf

  (
    g1728_n_spl_,
    g1728_n
  );


  buf

  (
    g1728_p_spl_,
    g1728_p
  );


  buf

  (
    g1730_p_spl_,
    g1730_p
  );


  buf

  (
    g1689_n_spl_,
    g1689_n
  );


  buf

  (
    g1730_n_spl_,
    g1730_n
  );


  buf

  (
    g1689_p_spl_,
    g1689_p
  );


  buf

  (
    g1731_n_spl_,
    g1731_n
  );


  buf

  (
    g1731_p_spl_,
    g1731_p
  );


  buf

  (
    g1733_p_spl_,
    g1733_p
  );


  buf

  (
    g1688_n_spl_,
    g1688_n
  );


  buf

  (
    g1733_n_spl_,
    g1733_n
  );


  buf

  (
    g1688_p_spl_,
    g1688_p
  );


  buf

  (
    g1734_n_spl_,
    g1734_n
  );


  buf

  (
    g1734_p_spl_,
    g1734_p
  );


  buf

  (
    g1736_p_spl_,
    g1736_p
  );


  buf

  (
    g1687_n_spl_,
    g1687_n
  );


  buf

  (
    g1736_n_spl_,
    g1736_n
  );


  buf

  (
    g1687_p_spl_,
    g1687_p
  );


  buf

  (
    g1737_n_spl_,
    g1737_n
  );


  buf

  (
    g1737_p_spl_,
    g1737_p
  );


  buf

  (
    g1739_n_spl_,
    g1739_n
  );


  buf

  (
    g1686_p_spl_,
    g1686_p
  );


  buf

  (
    g1740_p_spl_,
    g1740_p
  );


  buf

  (
    g1755_n_spl_,
    g1755_n
  );


  buf

  (
    g1754_n_spl_,
    g1754_n
  );


  buf

  (
    g1755_p_spl_,
    g1755_p
  );


  buf

  (
    g1754_p_spl_,
    g1754_p
  );


  buf

  (
    g1756_n_spl_,
    g1756_n
  );


  buf

  (
    g1756_p_spl_,
    g1756_p
  );


  buf

  (
    g1758_p_spl_,
    g1758_p
  );


  buf

  (
    g1753_n_spl_,
    g1753_n
  );


  buf

  (
    g1758_n_spl_,
    g1758_n
  );


  buf

  (
    g1753_p_spl_,
    g1753_p
  );


  buf

  (
    g1759_n_spl_,
    g1759_n
  );


  buf

  (
    g1759_p_spl_,
    g1759_p
  );


  buf

  (
    g1761_p_spl_,
    g1761_p
  );


  buf

  (
    g1752_n_spl_,
    g1752_n
  );


  buf

  (
    g1761_n_spl_,
    g1761_n
  );


  buf

  (
    g1752_p_spl_,
    g1752_p
  );


  buf

  (
    g1762_n_spl_,
    g1762_n
  );


  buf

  (
    g1762_p_spl_,
    g1762_p
  );


  buf

  (
    g1764_p_spl_,
    g1764_p
  );


  buf

  (
    g1751_n_spl_,
    g1751_n
  );


  buf

  (
    g1764_n_spl_,
    g1764_n
  );


  buf

  (
    g1751_p_spl_,
    g1751_p
  );


  buf

  (
    g1765_n_spl_,
    g1765_n
  );


  buf

  (
    g1765_p_spl_,
    g1765_p
  );


  buf

  (
    g1767_p_spl_,
    g1767_p
  );


  buf

  (
    g1750_n_spl_,
    g1750_n
  );


  buf

  (
    g1767_n_spl_,
    g1767_n
  );


  buf

  (
    g1750_p_spl_,
    g1750_p
  );


  buf

  (
    g1768_n_spl_,
    g1768_n
  );


  buf

  (
    g1768_p_spl_,
    g1768_p
  );


  buf

  (
    g1770_p_spl_,
    g1770_p
  );


  buf

  (
    g1749_n_spl_,
    g1749_n
  );


  buf

  (
    g1770_n_spl_,
    g1770_n
  );


  buf

  (
    g1749_p_spl_,
    g1749_p
  );


  buf

  (
    g1771_n_spl_,
    g1771_n
  );


  buf

  (
    g1771_p_spl_,
    g1771_p
  );


  buf

  (
    g1773_p_spl_,
    g1773_p
  );


  buf

  (
    g1748_n_spl_,
    g1748_n
  );


  buf

  (
    g1773_n_spl_,
    g1773_n
  );


  buf

  (
    g1748_p_spl_,
    g1748_p
  );


  buf

  (
    g1774_n_spl_,
    g1774_n
  );


  buf

  (
    g1774_p_spl_,
    g1774_p
  );


  buf

  (
    g1776_p_spl_,
    g1776_p
  );


  buf

  (
    g1747_n_spl_,
    g1747_n
  );


  buf

  (
    g1776_n_spl_,
    g1776_n
  );


  buf

  (
    g1747_p_spl_,
    g1747_p
  );


  buf

  (
    g1777_n_spl_,
    g1777_n
  );


  buf

  (
    g1777_p_spl_,
    g1777_p
  );


  buf

  (
    g1779_p_spl_,
    g1779_p
  );


  buf

  (
    g1746_n_spl_,
    g1746_n
  );


  buf

  (
    g1779_n_spl_,
    g1779_n
  );


  buf

  (
    g1746_p_spl_,
    g1746_p
  );


  buf

  (
    g1780_n_spl_,
    g1780_n
  );


  buf

  (
    g1780_p_spl_,
    g1780_p
  );


  buf

  (
    g1782_p_spl_,
    g1782_p
  );


  buf

  (
    g1745_n_spl_,
    g1745_n
  );


  buf

  (
    g1782_n_spl_,
    g1782_n
  );


  buf

  (
    g1745_p_spl_,
    g1745_p
  );


  buf

  (
    g1783_n_spl_,
    g1783_n
  );


  buf

  (
    g1783_p_spl_,
    g1783_p
  );


  buf

  (
    g1785_p_spl_,
    g1785_p
  );


  buf

  (
    g1744_n_spl_,
    g1744_n
  );


  buf

  (
    g1785_n_spl_,
    g1785_n
  );


  buf

  (
    g1744_p_spl_,
    g1744_p
  );


  buf

  (
    g1786_n_spl_,
    g1786_n
  );


  buf

  (
    g1786_p_spl_,
    g1786_p
  );


  buf

  (
    g1788_n_spl_,
    g1788_n
  );


  buf

  (
    g1743_p_spl_,
    g1743_p
  );


  buf

  (
    g1789_p_spl_,
    g1789_p
  );


  buf

  (
    g1802_n_spl_,
    g1802_n
  );


  buf

  (
    g1801_n_spl_,
    g1801_n
  );


  buf

  (
    g1802_p_spl_,
    g1802_p
  );


  buf

  (
    g1801_p_spl_,
    g1801_p
  );


  buf

  (
    g1803_n_spl_,
    g1803_n
  );


  buf

  (
    g1803_p_spl_,
    g1803_p
  );


  buf

  (
    g1805_p_spl_,
    g1805_p
  );


  buf

  (
    g1800_n_spl_,
    g1800_n
  );


  buf

  (
    g1805_n_spl_,
    g1805_n
  );


  buf

  (
    g1800_p_spl_,
    g1800_p
  );


  buf

  (
    g1806_n_spl_,
    g1806_n
  );


  buf

  (
    g1806_p_spl_,
    g1806_p
  );


  buf

  (
    g1808_p_spl_,
    g1808_p
  );


  buf

  (
    g1799_n_spl_,
    g1799_n
  );


  buf

  (
    g1808_n_spl_,
    g1808_n
  );


  buf

  (
    g1799_p_spl_,
    g1799_p
  );


  buf

  (
    g1809_n_spl_,
    g1809_n
  );


  buf

  (
    g1809_p_spl_,
    g1809_p
  );


  buf

  (
    g1811_p_spl_,
    g1811_p
  );


  buf

  (
    g1798_n_spl_,
    g1798_n
  );


  buf

  (
    g1811_n_spl_,
    g1811_n
  );


  buf

  (
    g1798_p_spl_,
    g1798_p
  );


  buf

  (
    g1812_n_spl_,
    g1812_n
  );


  buf

  (
    g1812_p_spl_,
    g1812_p
  );


  buf

  (
    g1814_p_spl_,
    g1814_p
  );


  buf

  (
    g1797_n_spl_,
    g1797_n
  );


  buf

  (
    g1814_n_spl_,
    g1814_n
  );


  buf

  (
    g1797_p_spl_,
    g1797_p
  );


  buf

  (
    g1815_n_spl_,
    g1815_n
  );


  buf

  (
    g1815_p_spl_,
    g1815_p
  );


  buf

  (
    g1817_p_spl_,
    g1817_p
  );


  buf

  (
    g1796_n_spl_,
    g1796_n
  );


  buf

  (
    g1817_n_spl_,
    g1817_n
  );


  buf

  (
    g1796_p_spl_,
    g1796_p
  );


  buf

  (
    g1818_n_spl_,
    g1818_n
  );


  buf

  (
    g1818_p_spl_,
    g1818_p
  );


  buf

  (
    g1820_p_spl_,
    g1820_p
  );


  buf

  (
    g1795_n_spl_,
    g1795_n
  );


  buf

  (
    g1820_n_spl_,
    g1820_n
  );


  buf

  (
    g1795_p_spl_,
    g1795_p
  );


  buf

  (
    g1821_n_spl_,
    g1821_n
  );


  buf

  (
    g1821_p_spl_,
    g1821_p
  );


  buf

  (
    g1823_p_spl_,
    g1823_p
  );


  buf

  (
    g1794_n_spl_,
    g1794_n
  );


  buf

  (
    g1823_n_spl_,
    g1823_n
  );


  buf

  (
    g1794_p_spl_,
    g1794_p
  );


  buf

  (
    g1824_n_spl_,
    g1824_n
  );


  buf

  (
    g1824_p_spl_,
    g1824_p
  );


  buf

  (
    g1826_p_spl_,
    g1826_p
  );


  buf

  (
    g1793_n_spl_,
    g1793_n
  );


  buf

  (
    g1826_n_spl_,
    g1826_n
  );


  buf

  (
    g1793_p_spl_,
    g1793_p
  );


  buf

  (
    g1827_n_spl_,
    g1827_n
  );


  buf

  (
    g1827_p_spl_,
    g1827_p
  );


  buf

  (
    g1829_n_spl_,
    g1829_n
  );


  buf

  (
    g1792_p_spl_,
    g1792_p
  );


  buf

  (
    g1830_p_spl_,
    g1830_p
  );


  buf

  (
    g1841_n_spl_,
    g1841_n
  );


  buf

  (
    g1840_n_spl_,
    g1840_n
  );


  buf

  (
    g1841_p_spl_,
    g1841_p
  );


  buf

  (
    g1840_p_spl_,
    g1840_p
  );


  buf

  (
    g1842_n_spl_,
    g1842_n
  );


  buf

  (
    g1842_p_spl_,
    g1842_p
  );


  buf

  (
    g1844_p_spl_,
    g1844_p
  );


  buf

  (
    g1839_n_spl_,
    g1839_n
  );


  buf

  (
    g1844_n_spl_,
    g1844_n
  );


  buf

  (
    g1839_p_spl_,
    g1839_p
  );


  buf

  (
    g1845_n_spl_,
    g1845_n
  );


  buf

  (
    g1845_p_spl_,
    g1845_p
  );


  buf

  (
    g1847_p_spl_,
    g1847_p
  );


  buf

  (
    g1838_n_spl_,
    g1838_n
  );


  buf

  (
    g1847_n_spl_,
    g1847_n
  );


  buf

  (
    g1838_p_spl_,
    g1838_p
  );


  buf

  (
    g1848_n_spl_,
    g1848_n
  );


  buf

  (
    g1848_p_spl_,
    g1848_p
  );


  buf

  (
    g1850_p_spl_,
    g1850_p
  );


  buf

  (
    g1837_n_spl_,
    g1837_n
  );


  buf

  (
    g1850_n_spl_,
    g1850_n
  );


  buf

  (
    g1837_p_spl_,
    g1837_p
  );


  buf

  (
    g1851_n_spl_,
    g1851_n
  );


  buf

  (
    g1851_p_spl_,
    g1851_p
  );


  buf

  (
    g1853_p_spl_,
    g1853_p
  );


  buf

  (
    g1836_n_spl_,
    g1836_n
  );


  buf

  (
    g1853_n_spl_,
    g1853_n
  );


  buf

  (
    g1836_p_spl_,
    g1836_p
  );


  buf

  (
    g1854_n_spl_,
    g1854_n
  );


  buf

  (
    g1854_p_spl_,
    g1854_p
  );


  buf

  (
    g1856_p_spl_,
    g1856_p
  );


  buf

  (
    g1835_n_spl_,
    g1835_n
  );


  buf

  (
    g1856_n_spl_,
    g1856_n
  );


  buf

  (
    g1835_p_spl_,
    g1835_p
  );


  buf

  (
    g1857_n_spl_,
    g1857_n
  );


  buf

  (
    g1857_p_spl_,
    g1857_p
  );


  buf

  (
    g1859_p_spl_,
    g1859_p
  );


  buf

  (
    g1834_n_spl_,
    g1834_n
  );


  buf

  (
    g1859_n_spl_,
    g1859_n
  );


  buf

  (
    g1834_p_spl_,
    g1834_p
  );


  buf

  (
    g1860_n_spl_,
    g1860_n
  );


  buf

  (
    g1860_p_spl_,
    g1860_p
  );


  buf

  (
    g1862_n_spl_,
    g1862_n
  );


  buf

  (
    g1833_p_spl_,
    g1833_p
  );


  buf

  (
    g1863_p_spl_,
    g1863_p
  );


  buf

  (
    g1872_n_spl_,
    g1872_n
  );


  buf

  (
    g1871_n_spl_,
    g1871_n
  );


  buf

  (
    g1872_p_spl_,
    g1872_p
  );


  buf

  (
    g1871_p_spl_,
    g1871_p
  );


  buf

  (
    g1873_n_spl_,
    g1873_n
  );


  buf

  (
    g1873_p_spl_,
    g1873_p
  );


  buf

  (
    g1875_p_spl_,
    g1875_p
  );


  buf

  (
    g1870_n_spl_,
    g1870_n
  );


  buf

  (
    g1875_n_spl_,
    g1875_n
  );


  buf

  (
    g1870_p_spl_,
    g1870_p
  );


  buf

  (
    g1876_n_spl_,
    g1876_n
  );


  buf

  (
    g1876_p_spl_,
    g1876_p
  );


  buf

  (
    g1878_p_spl_,
    g1878_p
  );


  buf

  (
    g1869_n_spl_,
    g1869_n
  );


  buf

  (
    g1878_n_spl_,
    g1878_n
  );


  buf

  (
    g1869_p_spl_,
    g1869_p
  );


  buf

  (
    g1879_n_spl_,
    g1879_n
  );


  buf

  (
    g1879_p_spl_,
    g1879_p
  );


  buf

  (
    g1881_p_spl_,
    g1881_p
  );


  buf

  (
    g1868_n_spl_,
    g1868_n
  );


  buf

  (
    g1881_n_spl_,
    g1881_n
  );


  buf

  (
    g1868_p_spl_,
    g1868_p
  );


  buf

  (
    g1882_n_spl_,
    g1882_n
  );


  buf

  (
    g1882_p_spl_,
    g1882_p
  );


  buf

  (
    g1884_p_spl_,
    g1884_p
  );


  buf

  (
    g1867_n_spl_,
    g1867_n
  );


  buf

  (
    g1884_n_spl_,
    g1884_n
  );


  buf

  (
    g1867_p_spl_,
    g1867_p
  );


  buf

  (
    g1885_n_spl_,
    g1885_n
  );


  buf

  (
    g1885_p_spl_,
    g1885_p
  );


  buf

  (
    g1887_n_spl_,
    g1887_n
  );


  buf

  (
    g1866_p_spl_,
    g1866_p
  );


  buf

  (
    g1888_p_spl_,
    g1888_p
  );


  buf

  (
    g1895_n_spl_,
    g1895_n
  );


  buf

  (
    g1894_n_spl_,
    g1894_n
  );


  buf

  (
    g1895_p_spl_,
    g1895_p
  );


  buf

  (
    g1894_p_spl_,
    g1894_p
  );


  buf

  (
    g1896_n_spl_,
    g1896_n
  );


  buf

  (
    g1896_p_spl_,
    g1896_p
  );


  buf

  (
    g1898_p_spl_,
    g1898_p
  );


  buf

  (
    g1893_n_spl_,
    g1893_n
  );


  buf

  (
    g1898_n_spl_,
    g1898_n
  );


  buf

  (
    g1893_p_spl_,
    g1893_p
  );


  buf

  (
    g1899_n_spl_,
    g1899_n
  );


  buf

  (
    g1899_p_spl_,
    g1899_p
  );


  buf

  (
    g1901_p_spl_,
    g1901_p
  );


  buf

  (
    g1892_n_spl_,
    g1892_n
  );


  buf

  (
    g1901_n_spl_,
    g1901_n
  );


  buf

  (
    g1892_p_spl_,
    g1892_p
  );


  buf

  (
    g1902_n_spl_,
    g1902_n
  );


  buf

  (
    g1902_p_spl_,
    g1902_p
  );


  buf

  (
    g1904_n_spl_,
    g1904_n
  );


  buf

  (
    g1891_p_spl_,
    g1891_p
  );


  buf

  (
    g1905_p_spl_,
    g1905_p
  );


  buf

  (
    g1909_n_spl_,
    g1909_n
  );


  buf

  (
    g1908_n_spl_,
    g1908_n
  );


  buf

  (
    g1909_p_spl_,
    g1909_p
  );


  buf

  (
    g1908_p_spl_,
    g1908_p
  );


  buf

  (
    g1910_n_spl_,
    g1910_n
  );


  buf

  (
    g1914_n_spl_,
    g1914_n
  );


endmodule
